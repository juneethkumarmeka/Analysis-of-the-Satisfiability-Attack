module basic_3000_30000_3500_25_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1788,In_2063);
xor U1 (N_1,In_859,In_1552);
xor U2 (N_2,In_1020,In_580);
or U3 (N_3,In_17,In_542);
nand U4 (N_4,In_2007,In_1783);
nor U5 (N_5,In_109,In_2796);
and U6 (N_6,In_443,In_2346);
nand U7 (N_7,In_1104,In_1118);
nand U8 (N_8,In_1094,In_1393);
nor U9 (N_9,In_2638,In_236);
or U10 (N_10,In_931,In_1259);
xor U11 (N_11,In_1097,In_792);
nand U12 (N_12,In_82,In_1798);
or U13 (N_13,In_2992,In_295);
or U14 (N_14,In_1958,In_1970);
nand U15 (N_15,In_1821,In_1446);
and U16 (N_16,In_2042,In_427);
nand U17 (N_17,In_664,In_861);
xnor U18 (N_18,In_838,In_763);
or U19 (N_19,In_690,In_1190);
or U20 (N_20,In_34,In_318);
or U21 (N_21,In_1575,In_2197);
and U22 (N_22,In_2429,In_194);
or U23 (N_23,In_1102,In_578);
nand U24 (N_24,In_216,In_2993);
and U25 (N_25,In_2045,In_2385);
nor U26 (N_26,In_1536,In_633);
and U27 (N_27,In_1306,In_1749);
or U28 (N_28,In_459,In_1315);
and U29 (N_29,In_758,In_2118);
or U30 (N_30,In_2859,In_2359);
nand U31 (N_31,In_2129,In_2682);
or U32 (N_32,In_2616,In_2089);
xnor U33 (N_33,In_2282,In_1171);
nor U34 (N_34,In_1903,In_2231);
or U35 (N_35,In_396,In_1321);
nor U36 (N_36,In_2391,In_2493);
xnor U37 (N_37,In_935,In_663);
nor U38 (N_38,In_239,In_2111);
nor U39 (N_39,In_1207,In_1916);
nor U40 (N_40,In_2749,In_48);
nand U41 (N_41,In_1281,In_1506);
and U42 (N_42,In_1981,In_2910);
xnor U43 (N_43,In_441,In_399);
or U44 (N_44,In_1373,In_2750);
nand U45 (N_45,In_1319,In_1408);
xor U46 (N_46,In_1496,In_2753);
nand U47 (N_47,In_1482,In_915);
nand U48 (N_48,In_937,In_2087);
nor U49 (N_49,In_1612,In_1467);
and U50 (N_50,In_285,In_1900);
nand U51 (N_51,In_195,In_1947);
or U52 (N_52,In_2527,In_1353);
xnor U53 (N_53,In_417,In_2785);
and U54 (N_54,In_2081,In_2286);
xnor U55 (N_55,In_52,In_1126);
nor U56 (N_56,In_848,In_1110);
or U57 (N_57,In_615,In_1567);
nand U58 (N_58,In_2053,In_1234);
nor U59 (N_59,In_1061,In_631);
and U60 (N_60,In_976,In_899);
nand U61 (N_61,In_1818,In_1803);
and U62 (N_62,In_984,In_1809);
and U63 (N_63,In_2412,In_1731);
xnor U64 (N_64,In_761,In_769);
and U65 (N_65,In_795,In_1713);
xnor U66 (N_66,In_928,In_1462);
nor U67 (N_67,In_1883,In_469);
and U68 (N_68,In_1638,In_1745);
nand U69 (N_69,In_1372,In_2787);
nor U70 (N_70,In_1115,In_423);
nor U71 (N_71,In_1577,In_2091);
nor U72 (N_72,In_2159,In_2948);
xor U73 (N_73,In_61,In_2372);
nand U74 (N_74,In_864,In_748);
nor U75 (N_75,In_2510,In_1652);
xor U76 (N_76,In_2699,In_2764);
and U77 (N_77,In_394,In_37);
and U78 (N_78,In_275,In_1295);
or U79 (N_79,In_193,In_1822);
nor U80 (N_80,In_1195,In_2812);
nand U81 (N_81,In_2839,In_1868);
nand U82 (N_82,In_1837,In_2138);
nand U83 (N_83,In_2647,In_1855);
nand U84 (N_84,In_2702,In_682);
nand U85 (N_85,In_1682,In_2117);
nand U86 (N_86,In_865,In_2605);
nor U87 (N_87,In_666,In_2675);
nor U88 (N_88,In_1833,In_1009);
nand U89 (N_89,In_632,In_1323);
and U90 (N_90,In_1326,In_463);
nand U91 (N_91,In_1170,In_719);
nor U92 (N_92,In_2137,In_1193);
xnor U93 (N_93,In_823,In_760);
and U94 (N_94,In_97,In_860);
and U95 (N_95,In_2641,In_780);
or U96 (N_96,In_729,In_2399);
or U97 (N_97,In_1334,In_1874);
and U98 (N_98,In_1298,In_139);
xor U99 (N_99,In_913,In_2665);
nand U100 (N_100,In_552,In_608);
nand U101 (N_101,In_2206,In_2108);
and U102 (N_102,In_1687,In_2590);
nand U103 (N_103,In_2247,In_957);
or U104 (N_104,In_2301,In_2440);
or U105 (N_105,In_1896,In_1166);
xor U106 (N_106,In_969,In_2719);
nand U107 (N_107,In_2496,In_1099);
nand U108 (N_108,In_2736,In_2691);
nand U109 (N_109,In_1367,In_562);
xnor U110 (N_110,In_618,In_809);
nand U111 (N_111,In_28,In_1401);
and U112 (N_112,In_1180,In_508);
and U113 (N_113,In_1699,In_1673);
or U114 (N_114,In_66,In_14);
and U115 (N_115,In_2002,In_359);
and U116 (N_116,In_2959,In_2791);
xnor U117 (N_117,In_468,In_2587);
and U118 (N_118,In_456,In_107);
and U119 (N_119,In_834,In_1279);
or U120 (N_120,In_2656,In_2082);
or U121 (N_121,In_2446,In_223);
or U122 (N_122,In_1152,In_1263);
nand U123 (N_123,In_870,In_1483);
xor U124 (N_124,In_2283,In_2645);
and U125 (N_125,In_1389,In_1379);
nor U126 (N_126,In_2744,In_1332);
xor U127 (N_127,In_1028,In_1480);
nor U128 (N_128,In_2631,In_2908);
nor U129 (N_129,In_1459,In_1975);
nor U130 (N_130,In_660,In_1225);
nand U131 (N_131,In_772,In_1430);
nand U132 (N_132,In_1014,In_1677);
nor U133 (N_133,In_651,In_2407);
xor U134 (N_134,In_171,In_500);
or U135 (N_135,In_2882,In_2986);
or U136 (N_136,In_2507,In_577);
and U137 (N_137,In_739,In_1562);
and U138 (N_138,In_627,In_148);
or U139 (N_139,In_2909,In_251);
nand U140 (N_140,In_2141,In_2975);
and U141 (N_141,In_324,In_2798);
nand U142 (N_142,In_2029,In_2503);
xor U143 (N_143,In_1895,In_1156);
nand U144 (N_144,In_2545,In_1787);
and U145 (N_145,In_1280,In_1831);
xor U146 (N_146,In_455,In_2660);
nor U147 (N_147,In_1993,In_1678);
and U148 (N_148,In_1985,In_2852);
nand U149 (N_149,In_1850,In_1651);
nand U150 (N_150,In_115,In_1712);
and U151 (N_151,In_2763,In_2394);
and U152 (N_152,In_2725,In_2062);
or U153 (N_153,In_2735,In_1558);
or U154 (N_154,In_551,In_2776);
xnor U155 (N_155,In_2274,In_319);
and U156 (N_156,In_829,In_2835);
nor U157 (N_157,In_2047,In_704);
xnor U158 (N_158,In_953,In_141);
nand U159 (N_159,In_2020,In_2658);
nand U160 (N_160,In_2293,In_2436);
nand U161 (N_161,In_1842,In_1365);
xor U162 (N_162,In_1992,In_661);
nor U163 (N_163,In_1939,In_1845);
xnor U164 (N_164,In_1595,In_2522);
nand U165 (N_165,In_2542,In_1364);
nor U166 (N_166,In_2547,In_181);
xnor U167 (N_167,In_1953,In_1262);
nor U168 (N_168,In_2677,In_717);
or U169 (N_169,In_2561,In_2668);
nor U170 (N_170,In_1666,In_2426);
xor U171 (N_171,In_2096,In_84);
or U172 (N_172,In_2718,In_225);
or U173 (N_173,In_231,In_1490);
nor U174 (N_174,In_1972,In_825);
and U175 (N_175,In_305,In_2410);
nor U176 (N_176,In_1721,In_2632);
nand U177 (N_177,In_2300,In_1576);
xor U178 (N_178,In_2949,In_2166);
nand U179 (N_179,In_2758,In_411);
xor U180 (N_180,In_596,In_1318);
nor U181 (N_181,In_2194,In_2099);
nand U182 (N_182,In_1986,In_985);
or U183 (N_183,In_862,In_2661);
or U184 (N_184,In_791,In_198);
or U185 (N_185,In_1314,In_1605);
and U186 (N_186,In_1534,In_1275);
nand U187 (N_187,In_385,In_1320);
or U188 (N_188,In_2075,In_1479);
nand U189 (N_189,In_2983,In_1136);
nor U190 (N_190,In_1924,In_1418);
xnor U191 (N_191,In_418,In_124);
or U192 (N_192,In_2145,In_1145);
and U193 (N_193,In_1342,In_624);
xor U194 (N_194,In_1050,In_401);
and U195 (N_195,In_404,In_185);
nor U196 (N_196,In_1265,In_2822);
xnor U197 (N_197,In_1048,In_2652);
or U198 (N_198,In_1226,In_806);
and U199 (N_199,In_308,In_10);
or U200 (N_200,In_894,In_2706);
or U201 (N_201,In_2664,In_2176);
or U202 (N_202,In_179,In_123);
and U203 (N_203,In_2774,In_1182);
nand U204 (N_204,In_1823,In_416);
nor U205 (N_205,In_157,In_2085);
or U206 (N_206,In_1101,In_668);
nor U207 (N_207,In_1722,In_2088);
or U208 (N_208,In_2279,In_1137);
nand U209 (N_209,In_2602,In_966);
and U210 (N_210,In_1002,In_2922);
xor U211 (N_211,In_1424,In_2315);
or U212 (N_212,In_238,In_696);
or U213 (N_213,In_1734,In_801);
nor U214 (N_214,In_1944,In_2729);
nand U215 (N_215,In_1998,In_1689);
and U216 (N_216,In_2343,In_465);
nand U217 (N_217,In_149,In_2460);
xor U218 (N_218,In_869,In_653);
and U219 (N_219,In_1354,In_515);
nor U220 (N_220,In_1602,In_786);
nand U221 (N_221,In_1287,In_510);
or U222 (N_222,In_912,In_778);
nor U223 (N_223,In_453,In_1657);
or U224 (N_224,In_2873,In_1269);
nor U225 (N_225,In_2851,In_2997);
xor U226 (N_226,In_634,In_1840);
nand U227 (N_227,In_1624,In_2926);
nand U228 (N_228,In_2708,In_1071);
nor U229 (N_229,In_911,In_2713);
and U230 (N_230,In_556,In_1214);
or U231 (N_231,In_20,In_1864);
xnor U232 (N_232,In_1766,In_1755);
nand U233 (N_233,In_182,In_1007);
xnor U234 (N_234,In_2698,In_1813);
xnor U235 (N_235,In_2840,In_2532);
nand U236 (N_236,In_1728,In_626);
nor U237 (N_237,In_486,In_1481);
xor U238 (N_238,In_2237,In_2671);
or U239 (N_239,In_2704,In_312);
or U240 (N_240,In_2485,In_1327);
nand U241 (N_241,In_2756,In_18);
nand U242 (N_242,In_481,In_924);
nand U243 (N_243,In_1033,In_1869);
or U244 (N_244,In_1247,In_2953);
or U245 (N_245,In_76,In_1108);
nor U246 (N_246,In_2657,In_2695);
nand U247 (N_247,In_2737,In_2328);
nor U248 (N_248,In_496,In_1244);
nor U249 (N_249,In_232,In_1396);
nand U250 (N_250,In_1839,In_1436);
and U251 (N_251,In_120,In_40);
and U252 (N_252,In_1264,In_1512);
xor U253 (N_253,In_2074,In_1059);
or U254 (N_254,In_371,In_2229);
xnor U255 (N_255,In_887,In_2519);
or U256 (N_256,In_2296,In_363);
and U257 (N_257,In_2620,In_21);
nor U258 (N_258,In_2627,In_2363);
nand U259 (N_259,In_755,In_2662);
nand U260 (N_260,In_1439,In_176);
or U261 (N_261,In_1088,In_991);
xnor U262 (N_262,In_595,In_1935);
nand U263 (N_263,In_958,In_2598);
and U264 (N_264,In_1829,In_2585);
and U265 (N_265,In_1475,In_2498);
or U266 (N_266,In_1410,In_2353);
and U267 (N_267,In_784,In_1290);
nor U268 (N_268,In_1627,In_623);
or U269 (N_269,In_2920,In_2896);
or U270 (N_270,In_513,In_684);
nor U271 (N_271,In_2678,In_871);
nor U272 (N_272,In_2371,In_31);
or U273 (N_273,In_2938,In_906);
and U274 (N_274,In_1750,In_2849);
nand U275 (N_275,In_942,In_846);
and U276 (N_276,In_92,In_307);
nand U277 (N_277,In_1125,In_1163);
nand U278 (N_278,In_2472,In_1824);
or U279 (N_279,In_954,In_614);
xor U280 (N_280,In_1926,In_2700);
or U281 (N_281,In_1511,In_1405);
nor U282 (N_282,In_2850,In_2894);
nand U283 (N_283,In_2649,In_2728);
nor U284 (N_284,In_2794,In_1616);
xnor U285 (N_285,In_1675,In_2222);
xnor U286 (N_286,In_568,In_837);
and U287 (N_287,In_1371,In_221);
nand U288 (N_288,In_2628,In_1715);
nand U289 (N_289,In_983,In_1569);
and U290 (N_290,In_1772,In_734);
xor U291 (N_291,In_2888,In_2960);
nand U292 (N_292,In_125,In_521);
nand U293 (N_293,In_2965,In_706);
nand U294 (N_294,In_810,In_589);
or U295 (N_295,In_1375,In_726);
nand U296 (N_296,In_2866,In_2816);
nor U297 (N_297,In_534,In_75);
nor U298 (N_298,In_2367,In_2098);
or U299 (N_299,In_2956,In_372);
nand U300 (N_300,In_2788,In_582);
nand U301 (N_301,In_2100,In_2513);
nor U302 (N_302,In_2121,In_1211);
or U303 (N_303,In_2619,In_2418);
nand U304 (N_304,In_1044,In_2941);
xnor U305 (N_305,In_1252,In_2720);
and U306 (N_306,In_2258,In_1584);
nand U307 (N_307,In_1685,In_2173);
xnor U308 (N_308,In_2152,In_2443);
and U309 (N_309,In_177,In_1862);
or U310 (N_310,In_1955,In_1267);
nor U311 (N_311,In_1814,In_153);
or U312 (N_312,In_471,In_2964);
xor U313 (N_313,In_524,In_1601);
nor U314 (N_314,In_1764,In_1585);
xnor U315 (N_315,In_197,In_2818);
and U316 (N_316,In_963,In_1168);
or U317 (N_317,In_410,In_2705);
nand U318 (N_318,In_2337,In_271);
xor U319 (N_319,In_2639,In_1425);
or U320 (N_320,In_2734,In_86);
nor U321 (N_321,In_2490,In_1971);
or U322 (N_322,In_2031,In_186);
or U323 (N_323,In_2884,In_2366);
and U324 (N_324,In_424,In_2403);
nand U325 (N_325,In_2504,In_93);
and U326 (N_326,In_1293,In_1502);
nor U327 (N_327,In_607,In_2239);
or U328 (N_328,In_1658,In_2448);
xnor U329 (N_329,In_2685,In_53);
xor U330 (N_330,In_2871,In_2101);
nand U331 (N_331,In_1592,In_2961);
xor U332 (N_332,In_619,In_2921);
nor U333 (N_333,In_27,In_2535);
nand U334 (N_334,In_1856,In_1600);
or U335 (N_335,In_1882,In_2978);
xnor U336 (N_336,In_2825,In_1095);
or U337 (N_337,In_1113,In_635);
and U338 (N_338,In_2287,In_2770);
nor U339 (N_339,In_1802,In_466);
and U340 (N_340,In_2183,In_317);
nand U341 (N_341,In_2548,In_1179);
or U342 (N_342,In_2611,In_322);
or U343 (N_343,In_2663,In_543);
and U344 (N_344,In_1478,In_384);
and U345 (N_345,In_2277,In_1793);
or U346 (N_346,In_155,In_1016);
nor U347 (N_347,In_1487,In_2468);
xnor U348 (N_348,In_167,In_364);
and U349 (N_349,In_1625,In_2876);
or U350 (N_350,In_1236,In_2175);
nor U351 (N_351,In_2955,In_1588);
and U352 (N_352,In_2889,In_2903);
and U353 (N_353,In_178,In_1780);
xor U354 (N_354,In_2610,In_2349);
or U355 (N_355,In_2586,In_896);
xnor U356 (N_356,In_916,In_2752);
or U357 (N_357,In_2241,In_1679);
nor U358 (N_358,In_1646,In_693);
and U359 (N_359,In_669,In_2116);
xnor U360 (N_360,In_2801,In_2743);
or U361 (N_361,In_1027,In_2044);
xor U362 (N_362,In_1172,In_1420);
or U363 (N_363,In_1756,In_2567);
xor U364 (N_364,In_546,In_1284);
nand U365 (N_365,In_1065,In_1617);
or U366 (N_366,In_2717,In_929);
nor U367 (N_367,In_347,In_1933);
or U368 (N_368,In_1383,In_497);
and U369 (N_369,In_2212,In_1196);
nor U370 (N_370,In_2238,In_60);
and U371 (N_371,In_412,In_575);
nor U372 (N_372,In_1786,In_2731);
or U373 (N_373,In_2369,In_2558);
nand U374 (N_374,In_414,In_2898);
xnor U375 (N_375,In_491,In_298);
or U376 (N_376,In_2797,In_1920);
xnor U377 (N_377,In_1526,In_2006);
xnor U378 (N_378,In_930,In_1701);
nor U379 (N_379,In_2957,In_545);
or U380 (N_380,In_1976,In_1520);
or U381 (N_381,In_2267,In_2546);
xnor U382 (N_382,In_494,In_345);
nand U383 (N_383,In_2692,In_286);
xnor U384 (N_384,In_1025,In_1382);
xnor U385 (N_385,In_1181,In_1085);
and U386 (N_386,In_1476,In_2120);
or U387 (N_387,In_2122,In_946);
and U388 (N_388,In_2489,In_827);
and U389 (N_389,In_2807,In_1779);
and U390 (N_390,In_832,In_1243);
or U391 (N_391,In_1254,In_2985);
or U392 (N_392,In_974,In_1455);
and U393 (N_393,In_2273,In_1209);
nor U394 (N_394,In_1134,In_1357);
and U395 (N_395,In_993,In_1504);
xor U396 (N_396,In_343,In_2364);
nor U397 (N_397,In_1827,In_1784);
nand U398 (N_398,In_12,In_1988);
or U399 (N_399,In_1865,In_113);
xor U400 (N_400,In_1544,In_254);
nor U401 (N_401,In_2172,In_1176);
or U402 (N_402,In_750,In_1212);
and U403 (N_403,In_2452,In_977);
and U404 (N_404,In_1630,In_2052);
nand U405 (N_405,In_927,In_87);
xor U406 (N_406,In_2917,In_1497);
xnor U407 (N_407,In_1348,In_1036);
nand U408 (N_408,In_1349,In_1161);
and U409 (N_409,In_1892,In_2179);
or U410 (N_410,In_2265,In_816);
and U411 (N_411,In_527,In_1934);
or U412 (N_412,In_890,In_2009);
or U413 (N_413,In_2018,In_218);
or U414 (N_414,In_722,In_1744);
and U415 (N_415,In_2803,In_2757);
nor U416 (N_416,In_2109,In_2775);
xor U417 (N_417,In_2442,In_2259);
or U418 (N_418,In_678,In_2240);
nand U419 (N_419,In_1537,In_1119);
nand U420 (N_420,In_721,In_77);
or U421 (N_421,In_978,In_1989);
nand U422 (N_422,In_1587,In_292);
xor U423 (N_423,In_1338,In_1051);
and U424 (N_424,In_1811,In_1296);
nor U425 (N_425,In_1256,In_1555);
and U426 (N_426,In_484,In_174);
and U427 (N_427,In_2306,In_2425);
and U428 (N_428,In_970,In_2462);
or U429 (N_429,In_573,In_1308);
or U430 (N_430,In_1457,In_2572);
or U431 (N_431,In_46,In_2565);
xnor U432 (N_432,In_2773,In_2464);
xnor U433 (N_433,In_144,In_2036);
nor U434 (N_434,In_2411,In_2595);
or U435 (N_435,In_1914,In_393);
xnor U436 (N_436,In_1167,In_1727);
nor U437 (N_437,In_2424,In_2827);
xor U438 (N_438,In_2147,In_948);
nand U439 (N_439,In_1019,In_2476);
nor U440 (N_440,In_2936,In_1807);
nor U441 (N_441,In_2626,In_1565);
and U442 (N_442,In_876,In_2174);
xnor U443 (N_443,In_1055,In_1231);
and U444 (N_444,In_2538,In_2612);
nor U445 (N_445,In_2591,In_1192);
and U446 (N_446,In_703,In_517);
and U447 (N_447,In_112,In_2709);
xor U448 (N_448,In_836,In_2479);
nor U449 (N_449,In_2636,In_1162);
and U450 (N_450,In_2039,In_2454);
or U451 (N_451,In_1863,In_2982);
nand U452 (N_452,In_2913,In_1374);
nand U453 (N_453,In_2086,In_600);
xor U454 (N_454,In_821,In_2642);
and U455 (N_455,In_1834,In_22);
or U456 (N_456,In_1003,In_636);
or U457 (N_457,In_2670,In_288);
and U458 (N_458,In_1858,In_1676);
xnor U459 (N_459,In_2979,In_1491);
nor U460 (N_460,In_611,In_897);
or U461 (N_461,In_881,In_1370);
and U462 (N_462,In_73,In_1884);
xor U463 (N_463,In_2326,In_818);
and U464 (N_464,In_1683,In_2083);
and U465 (N_465,In_1164,In_1366);
nor U466 (N_466,In_1517,In_1681);
xor U467 (N_467,In_445,In_1197);
and U468 (N_468,In_41,In_1800);
nor U469 (N_469,In_539,In_741);
nand U470 (N_470,In_504,In_1794);
nand U471 (N_471,In_2484,In_2973);
or U472 (N_472,In_2600,In_938);
or U473 (N_473,In_528,In_1710);
xor U474 (N_474,In_226,In_485);
or U475 (N_475,In_1928,In_1165);
nand U476 (N_476,In_749,In_923);
or U477 (N_477,In_476,In_1859);
and U478 (N_478,In_173,In_1796);
nor U479 (N_479,In_212,In_360);
or U480 (N_480,In_1525,In_2214);
nor U481 (N_481,In_1345,In_857);
and U482 (N_482,In_1335,In_1757);
xnor U483 (N_483,In_2487,In_35);
nor U484 (N_484,In_900,In_2606);
nor U485 (N_485,In_2566,In_557);
nor U486 (N_486,In_1505,In_276);
or U487 (N_487,In_723,In_2581);
and U488 (N_488,In_507,In_1550);
xnor U489 (N_489,In_731,In_169);
or U490 (N_490,In_1980,In_2294);
xnor U491 (N_491,In_2584,In_103);
nor U492 (N_492,In_1203,In_2597);
or U493 (N_493,In_1488,In_440);
nor U494 (N_494,In_1070,In_511);
nor U495 (N_495,In_2723,In_2161);
or U496 (N_496,In_355,In_1999);
xnor U497 (N_497,In_2492,In_189);
nor U498 (N_498,In_1596,In_44);
or U499 (N_499,In_569,In_2946);
or U500 (N_500,In_1128,In_2303);
or U501 (N_501,In_2916,In_2578);
nor U502 (N_502,In_2065,In_2863);
xor U503 (N_503,In_1671,In_2762);
or U504 (N_504,In_2515,In_2525);
nand U505 (N_505,In_1806,In_955);
nand U506 (N_506,In_350,In_1899);
or U507 (N_507,In_2939,In_665);
xnor U508 (N_508,In_1248,In_828);
nor U509 (N_509,In_1400,In_1307);
nor U510 (N_510,In_85,In_2185);
nor U511 (N_511,In_1031,In_2727);
xnor U512 (N_512,In_1921,In_43);
and U513 (N_513,In_242,In_695);
or U514 (N_514,In_531,In_2192);
and U515 (N_515,In_2843,In_2795);
or U516 (N_516,In_671,In_590);
and U517 (N_517,In_1736,In_2090);
xor U518 (N_518,In_2800,In_766);
and U519 (N_519,In_1548,In_1283);
xor U520 (N_520,In_2127,In_1041);
or U521 (N_521,In_567,In_11);
and U522 (N_522,In_1035,In_822);
nand U523 (N_523,In_1634,In_880);
nand U524 (N_524,In_1387,In_248);
and U525 (N_525,In_2115,In_2105);
or U526 (N_526,In_2246,In_2613);
or U527 (N_527,In_426,In_2524);
nor U528 (N_528,In_561,In_776);
nor U529 (N_529,In_130,In_279);
nor U530 (N_530,In_2401,In_2892);
nor U531 (N_531,In_1951,In_2103);
nor U532 (N_532,In_1688,In_775);
or U533 (N_533,In_63,In_968);
xnor U534 (N_534,In_2064,In_1138);
nor U535 (N_535,In_674,In_2205);
nor U536 (N_536,In_785,In_909);
or U537 (N_537,In_2486,In_602);
or U538 (N_538,In_1805,In_1589);
and U539 (N_539,In_2897,In_1741);
nor U540 (N_540,In_2741,In_1904);
and U541 (N_541,In_1540,In_2772);
xor U542 (N_542,In_2316,In_146);
xnor U543 (N_543,In_874,In_609);
and U544 (N_544,In_268,In_431);
nor U545 (N_545,In_2202,In_2434);
xnor U546 (N_546,In_1782,In_2541);
and U547 (N_547,In_2623,In_2517);
nand U548 (N_548,In_2732,In_2022);
nor U549 (N_549,In_2996,In_1978);
nand U550 (N_550,In_247,In_2943);
and U551 (N_551,In_188,In_1228);
nor U552 (N_552,In_2336,In_2124);
and U553 (N_553,In_2135,In_2169);
nand U554 (N_554,In_1608,In_1846);
nor U555 (N_555,In_1919,In_1109);
xor U556 (N_556,In_2748,In_2684);
or U557 (N_557,In_1133,In_571);
xnor U558 (N_558,In_2146,In_2689);
nor U559 (N_559,In_2826,In_1887);
nand U560 (N_560,In_1556,In_32);
nor U561 (N_561,In_2126,In_951);
nand U562 (N_562,In_1274,In_1549);
nand U563 (N_563,In_2270,In_2203);
xnor U564 (N_564,In_961,In_134);
nand U565 (N_565,In_243,In_540);
nand U566 (N_566,In_1022,In_1940);
xnor U567 (N_567,In_2375,In_2551);
nand U568 (N_568,In_840,In_2151);
or U569 (N_569,In_2420,In_1222);
and U570 (N_570,In_914,In_2648);
nor U571 (N_571,In_1123,In_2999);
xnor U572 (N_572,In_116,In_2637);
or U573 (N_573,In_1359,In_2778);
and U574 (N_574,In_340,In_2674);
and U575 (N_575,In_2942,In_203);
nor U576 (N_576,In_1987,In_728);
nor U577 (N_577,In_2019,In_1740);
nor U578 (N_578,In_2059,In_956);
or U579 (N_579,In_2072,In_337);
nand U580 (N_580,In_2416,In_1854);
nand U581 (N_581,In_101,In_2571);
or U582 (N_582,In_1754,In_1268);
nand U583 (N_583,In_2874,In_2837);
nand U584 (N_584,In_652,In_1063);
nand U585 (N_585,In_444,In_2810);
nor U586 (N_586,In_2149,In_38);
nor U587 (N_587,In_1936,In_2004);
nor U588 (N_588,In_2511,In_2128);
nand U589 (N_589,In_2730,In_2322);
or U590 (N_590,In_1983,In_1523);
or U591 (N_591,In_2060,In_1272);
xor U592 (N_592,In_39,In_2374);
nor U593 (N_593,In_1765,In_1594);
or U594 (N_594,In_2102,In_1498);
and U595 (N_595,In_234,In_2745);
nand U596 (N_596,In_1038,In_1294);
or U597 (N_597,In_707,In_1344);
xnor U598 (N_598,In_1224,In_2688);
or U599 (N_599,In_1443,In_2833);
or U600 (N_600,In_686,In_919);
nor U601 (N_601,In_2607,In_1876);
nand U602 (N_602,In_1438,In_192);
or U603 (N_603,In_2995,In_1597);
xor U604 (N_604,In_679,In_2604);
nor U605 (N_605,In_2594,In_505);
and U606 (N_606,In_720,In_1647);
nand U607 (N_607,In_1598,In_629);
xnor U608 (N_608,In_1414,In_2962);
or U609 (N_609,In_1852,In_2861);
nand U610 (N_610,In_2113,In_1718);
nand U611 (N_611,In_2189,In_2932);
or U612 (N_612,In_1461,In_2114);
or U613 (N_613,In_2355,In_1460);
nand U614 (N_614,In_368,In_2272);
nor U615 (N_615,In_137,In_2);
nand U616 (N_616,In_782,In_464);
xnor U617 (N_617,In_1603,In_2123);
or U618 (N_618,In_2164,In_2491);
and U619 (N_619,In_2382,In_1377);
nand U620 (N_620,In_555,In_820);
or U621 (N_621,In_419,In_709);
nand U622 (N_622,In_2805,In_1412);
xnor U623 (N_623,In_2432,In_1711);
nor U624 (N_624,In_506,In_2480);
and U625 (N_625,In_409,In_1907);
and U626 (N_626,In_1698,In_605);
nor U627 (N_627,In_2906,In_2829);
nand U628 (N_628,In_2302,In_1303);
xor U629 (N_629,In_655,In_2919);
xnor U630 (N_630,In_2266,In_1060);
nand U631 (N_631,In_2280,In_1111);
nand U632 (N_632,In_2570,In_1149);
nor U633 (N_633,In_6,In_1289);
xnor U634 (N_634,In_1808,In_1067);
or U635 (N_635,In_2991,In_802);
and U636 (N_636,In_2512,In_2066);
nand U637 (N_637,In_1242,In_2156);
and U638 (N_638,In_425,In_1034);
nor U639 (N_639,In_2003,In_2935);
nand U640 (N_640,In_30,In_2177);
and U641 (N_641,In_483,In_2726);
and U642 (N_642,In_747,In_2806);
or U643 (N_643,In_395,In_2386);
or U644 (N_644,In_1043,In_391);
or U645 (N_645,In_922,In_1774);
and U646 (N_646,In_2621,In_365);
nor U647 (N_647,In_1189,In_1905);
nand U648 (N_648,In_1910,In_1219);
nand U649 (N_649,In_2481,In_299);
nor U650 (N_650,In_430,In_2023);
and U651 (N_651,In_2528,In_2559);
xor U652 (N_652,In_2298,In_1702);
xor U653 (N_653,In_457,In_1522);
nand U654 (N_654,In_1258,In_1730);
and U655 (N_655,In_147,In_458);
or U656 (N_656,In_1751,In_518);
nor U657 (N_657,In_658,In_2579);
or U658 (N_658,In_413,In_2162);
nand U659 (N_659,In_882,In_131);
nand U660 (N_660,In_136,In_235);
nor U661 (N_661,In_280,In_2181);
and U662 (N_662,In_1116,In_1963);
nor U663 (N_663,In_62,In_2421);
nor U664 (N_664,In_904,In_1217);
xnor U665 (N_665,In_550,In_1337);
nor U666 (N_666,In_2439,In_2107);
nor U667 (N_667,In_856,In_200);
nor U668 (N_668,In_2694,In_277);
and U669 (N_669,In_2614,In_1770);
nor U670 (N_670,In_49,In_80);
nand U671 (N_671,In_1435,In_252);
or U672 (N_672,In_1440,In_2010);
and U673 (N_673,In_2815,In_2617);
nor U674 (N_674,In_353,In_1606);
or U675 (N_675,In_438,In_56);
xor U676 (N_676,In_111,In_306);
or U677 (N_677,In_1516,In_2555);
or U678 (N_678,In_2221,In_187);
or U679 (N_679,In_118,In_2877);
and U680 (N_680,In_1300,In_1445);
xor U681 (N_681,In_1157,In_544);
nor U682 (N_682,In_207,In_269);
or U683 (N_683,In_1120,In_1667);
or U684 (N_684,In_811,In_2844);
nand U685 (N_685,In_2881,In_830);
and U686 (N_686,In_2232,In_878);
xor U687 (N_687,In_529,In_2970);
and U688 (N_688,In_2712,In_400);
nor U689 (N_689,In_1716,In_799);
or U690 (N_690,In_2347,In_2733);
or U691 (N_691,In_849,In_926);
nor U692 (N_692,In_2817,In_708);
and U693 (N_693,In_240,In_382);
or U694 (N_694,In_2823,In_1008);
xnor U695 (N_695,In_2860,In_2471);
or U696 (N_696,In_522,In_2325);
xnor U697 (N_697,In_388,In_1297);
and U698 (N_698,In_472,In_478);
nor U699 (N_699,In_1767,In_918);
or U700 (N_700,In_1361,In_1692);
xnor U701 (N_701,In_1819,In_1691);
nor U702 (N_702,In_1129,In_1521);
or U703 (N_703,In_2216,In_1954);
nand U704 (N_704,In_2201,In_932);
and U705 (N_705,In_74,In_2449);
nor U706 (N_706,In_1187,In_547);
nor U707 (N_707,In_1230,In_773);
nor U708 (N_708,In_1100,In_261);
xnor U709 (N_709,In_70,In_884);
nand U710 (N_710,In_2739,In_2501);
xnor U711 (N_711,In_1832,In_2769);
nand U712 (N_712,In_1836,In_2944);
or U713 (N_713,In_2554,In_1559);
nor U714 (N_714,In_1339,In_1964);
nor U715 (N_715,In_1816,In_2428);
and U716 (N_716,In_964,In_519);
xor U717 (N_717,In_2408,In_676);
or U718 (N_718,In_2244,In_208);
xnor U719 (N_719,In_537,In_950);
nor U720 (N_720,In_1959,In_362);
nand U721 (N_721,In_2654,In_1557);
or U722 (N_722,In_868,In_1311);
or U723 (N_723,In_2466,In_1890);
xnor U724 (N_724,In_2969,In_138);
xor U725 (N_725,In_2076,In_2865);
or U726 (N_726,In_1158,In_1251);
nor U727 (N_727,In_889,In_853);
and U728 (N_728,In_357,In_712);
or U729 (N_729,In_1639,In_1591);
xor U730 (N_730,In_990,In_2187);
or U731 (N_731,In_2160,In_616);
nand U732 (N_732,In_2071,In_2208);
nand U733 (N_733,In_2397,In_1227);
and U734 (N_734,In_2721,In_1781);
nand U735 (N_735,In_2024,In_1237);
nand U736 (N_736,In_2278,In_2940);
nand U737 (N_737,In_2878,In_563);
xnor U738 (N_738,In_2344,In_2134);
and U739 (N_739,In_26,In_592);
nor U740 (N_740,In_981,In_523);
nand U741 (N_741,In_2186,In_1737);
nand U742 (N_742,In_905,In_647);
or U743 (N_743,In_858,In_1432);
nor U744 (N_744,In_2857,In_1472);
or U745 (N_745,In_1448,In_449);
nor U746 (N_746,In_2937,In_2872);
and U747 (N_747,In_710,In_2398);
and U748 (N_748,In_1650,In_1330);
nor U749 (N_749,In_2710,In_1341);
or U750 (N_750,In_1618,In_1762);
xor U751 (N_751,In_604,In_1885);
or U752 (N_752,In_1769,In_1994);
xnor U753 (N_753,In_331,In_866);
nor U754 (N_754,In_1937,In_603);
and U755 (N_755,In_2945,In_2793);
and U756 (N_756,In_1422,In_437);
nand U757 (N_757,In_2417,In_439);
and U758 (N_758,In_1142,In_161);
or U759 (N_759,In_516,In_1700);
and U760 (N_760,In_2666,In_1417);
and U761 (N_761,In_1915,In_2320);
xor U762 (N_762,In_320,In_621);
and U763 (N_763,In_1542,In_301);
xnor U764 (N_764,In_1500,In_1208);
nand U765 (N_765,In_274,In_2140);
nor U766 (N_766,In_2582,In_745);
nand U767 (N_767,In_328,In_2026);
and U768 (N_768,In_2886,In_314);
and U769 (N_769,In_151,In_1660);
xor U770 (N_770,In_2080,In_579);
or U771 (N_771,In_790,In_1477);
and U772 (N_772,In_570,In_2473);
nand U773 (N_773,In_1621,In_150);
xor U774 (N_774,In_2041,In_2500);
xor U775 (N_775,In_1112,In_879);
or U776 (N_776,In_2153,In_1356);
nand U777 (N_777,In_2168,In_2972);
or U778 (N_778,In_2925,In_952);
and U779 (N_779,In_106,In_1021);
or U780 (N_780,In_2930,In_2219);
xnor U781 (N_781,In_1723,In_1278);
nand U782 (N_782,In_2574,In_1804);
nand U783 (N_783,In_1743,In_24);
or U784 (N_784,In_2544,In_2669);
nor U785 (N_785,In_1202,In_1573);
nor U786 (N_786,In_2224,In_2924);
nor U787 (N_787,In_672,In_2027);
and U788 (N_788,In_1923,In_1246);
xor U789 (N_789,In_1826,In_622);
nor U790 (N_790,In_2079,In_1081);
xor U791 (N_791,In_1708,In_1066);
and U792 (N_792,In_1395,In_2470);
nand U793 (N_793,In_2196,In_1889);
or U794 (N_794,In_2783,In_2577);
xor U795 (N_795,In_2404,In_327);
or U796 (N_796,In_565,In_2746);
or U797 (N_797,In_237,In_1929);
or U798 (N_798,In_2516,In_1977);
nor U799 (N_799,In_110,In_2106);
xnor U800 (N_800,In_2198,In_2245);
and U801 (N_801,In_1866,In_1039);
xor U802 (N_802,In_1720,In_1042);
nand U803 (N_803,In_1004,In_2459);
nor U804 (N_804,In_886,In_1350);
and U805 (N_805,In_290,In_2904);
or U806 (N_806,In_1891,In_95);
xnor U807 (N_807,In_2078,In_2340);
and U808 (N_808,In_1574,In_163);
nand U809 (N_809,In_2069,In_159);
xor U810 (N_810,In_1029,In_925);
and U811 (N_811,In_2673,In_2057);
xnor U812 (N_812,In_2667,In_711);
nand U813 (N_813,In_996,In_2453);
nor U814 (N_814,In_645,In_461);
nor U815 (N_815,In_2900,In_777);
nand U816 (N_816,In_2771,In_129);
nand U817 (N_817,In_839,In_751);
and U818 (N_818,In_1191,In_1815);
xor U819 (N_819,In_422,In_1670);
nand U820 (N_820,In_1402,In_71);
nor U821 (N_821,In_1539,In_2834);
nand U822 (N_822,In_959,In_1927);
nand U823 (N_823,In_1669,In_872);
nor U824 (N_824,In_2235,In_135);
xnor U825 (N_825,In_2655,In_1201);
xnor U826 (N_826,In_214,In_126);
xor U827 (N_827,In_1114,In_2393);
nor U828 (N_828,In_1735,In_140);
or U829 (N_829,In_1229,In_670);
xnor U830 (N_830,In_2931,In_1995);
nor U831 (N_831,In_2092,In_1271);
xor U832 (N_832,In_2592,In_2281);
xor U833 (N_833,In_610,In_1083);
and U834 (N_834,In_132,In_2220);
or U835 (N_835,In_1363,In_1178);
nor U836 (N_836,In_1260,In_333);
or U837 (N_837,In_1140,In_1261);
nor U838 (N_838,In_1049,In_89);
xor U839 (N_839,In_127,In_1495);
and U840 (N_840,In_289,In_1662);
nor U841 (N_841,In_2650,In_2633);
nand U842 (N_842,In_1979,In_1385);
nor U843 (N_843,In_257,In_2370);
nor U844 (N_844,In_2139,In_548);
xor U845 (N_845,In_100,In_2441);
and U846 (N_846,In_1738,In_381);
xnor U847 (N_847,In_296,In_1930);
nand U848 (N_848,In_16,In_638);
or U849 (N_849,In_2990,In_877);
xnor U850 (N_850,In_2552,In_1580);
or U851 (N_851,In_1820,In_291);
and U852 (N_852,In_183,In_2971);
nand U853 (N_853,In_2643,In_1291);
nor U854 (N_854,In_650,In_1962);
nand U855 (N_855,In_2568,In_1238);
nor U856 (N_856,In_1604,In_2260);
and U857 (N_857,In_284,In_2165);
nor U858 (N_858,In_783,In_206);
and U859 (N_859,In_1340,In_1431);
nor U860 (N_860,In_2864,In_1752);
or U861 (N_861,In_2271,In_1106);
nand U862 (N_862,In_941,In_2508);
or U863 (N_863,In_2557,In_1648);
nand U864 (N_864,In_744,In_1415);
and U865 (N_865,In_2040,In_2868);
nor U866 (N_866,In_253,In_742);
nor U867 (N_867,In_1005,In_1531);
nor U868 (N_868,In_2204,In_2125);
or U869 (N_869,In_503,In_2514);
or U870 (N_870,In_477,In_685);
xor U871 (N_871,In_1040,In_2021);
or U872 (N_872,In_96,In_2914);
nor U873 (N_873,In_688,In_1620);
nor U874 (N_874,In_1773,In_1139);
or U875 (N_875,In_1141,In_117);
or U876 (N_876,In_705,In_1011);
and U877 (N_877,In_1089,In_933);
xnor U878 (N_878,In_2608,In_1997);
xnor U879 (N_879,In_1656,In_1532);
nor U880 (N_880,In_2163,In_1135);
or U881 (N_881,In_2437,In_2596);
nor U882 (N_882,In_1668,In_1077);
xor U883 (N_883,In_727,In_1086);
and U884 (N_884,In_262,In_1000);
xnor U885 (N_885,In_1032,In_344);
xnor U886 (N_886,In_1579,In_2035);
and U887 (N_887,In_1218,In_2148);
or U888 (N_888,In_1894,In_2167);
nor U889 (N_889,In_736,In_1233);
nand U890 (N_890,In_588,In_979);
nor U891 (N_891,In_2305,In_489);
or U892 (N_892,In_813,In_1693);
nor U893 (N_893,In_718,In_1776);
nand U894 (N_894,In_1386,In_1902);
nor U895 (N_895,In_2838,In_2362);
or U896 (N_896,In_1205,In_490);
nor U897 (N_897,In_2494,In_1406);
xnor U898 (N_898,In_2357,In_1056);
or U899 (N_899,In_1464,In_901);
or U900 (N_900,In_2622,In_2215);
and U901 (N_901,In_495,In_1474);
or U902 (N_902,In_1285,In_1543);
xor U903 (N_903,In_2821,In_628);
xnor U904 (N_904,In_1886,In_1148);
xor U905 (N_905,In_166,In_1851);
and U906 (N_906,In_656,In_2414);
or U907 (N_907,In_1768,In_512);
nand U908 (N_908,In_940,In_667);
nor U909 (N_909,In_2784,In_473);
xor U910 (N_910,In_210,In_1838);
nor U911 (N_911,In_2056,In_1632);
or U912 (N_912,In_51,In_2813);
nand U913 (N_913,In_725,In_2766);
or U914 (N_914,In_1922,In_1877);
or U915 (N_915,In_986,In_1861);
nor U916 (N_916,In_1486,In_1938);
and U917 (N_917,In_1317,In_1159);
or U918 (N_918,In_121,In_1763);
nor U919 (N_919,In_1973,In_2575);
or U920 (N_920,In_797,In_574);
and U921 (N_921,In_2885,In_493);
xor U922 (N_922,In_798,In_1725);
nor U923 (N_923,In_841,In_2902);
and U924 (N_924,In_771,In_1967);
xnor U925 (N_925,In_752,In_1913);
xnor U926 (N_926,In_2431,In_1880);
nand U927 (N_927,In_433,In_199);
xor U928 (N_928,In_560,In_1789);
nand U929 (N_929,In_1847,In_788);
and U930 (N_930,In_1322,In_630);
nand U931 (N_931,In_2533,In_903);
xnor U932 (N_932,In_2384,In_273);
nand U933 (N_933,In_2687,In_1599);
nor U934 (N_934,In_1974,In_1130);
nor U935 (N_935,In_1631,In_598);
nor U936 (N_936,In_190,In_1759);
xnor U937 (N_937,In_1447,In_2740);
nor U938 (N_938,In_620,In_779);
or U939 (N_939,In_1949,In_789);
nand U940 (N_940,In_2912,In_1452);
nor U941 (N_941,In_304,In_2780);
and U942 (N_942,In_591,In_143);
or U943 (N_943,In_1982,In_794);
or U944 (N_944,In_2379,In_1908);
or U945 (N_945,In_501,In_302);
xor U946 (N_946,In_259,In_498);
xnor U947 (N_947,In_403,In_2846);
nor U948 (N_948,In_323,In_264);
and U949 (N_949,In_1538,In_2312);
nor U950 (N_950,In_850,In_2963);
or U951 (N_951,In_398,In_448);
nor U952 (N_952,In_2782,In_460);
and U953 (N_953,In_1655,In_2048);
xnor U954 (N_954,In_2351,In_1965);
or U955 (N_955,In_558,In_1945);
and U956 (N_956,In_796,In_2954);
and U957 (N_957,In_2869,In_1232);
nand U958 (N_958,In_1777,In_1853);
nor U959 (N_959,In_354,In_2755);
xor U960 (N_960,In_361,In_738);
nand U961 (N_961,In_2276,In_470);
and U962 (N_962,In_2701,In_2465);
and U963 (N_963,In_2895,In_1324);
and U964 (N_964,In_348,In_2624);
nand U965 (N_965,In_826,In_2505);
xor U966 (N_966,In_341,In_1672);
and U967 (N_967,In_2264,In_2209);
and U968 (N_968,In_1277,In_2352);
nor U969 (N_969,In_2883,In_1572);
nor U970 (N_970,In_694,In_1253);
xnor U971 (N_971,In_691,In_1046);
nor U972 (N_972,In_325,In_1778);
nand U973 (N_973,In_2915,In_54);
nor U974 (N_974,In_1380,In_641);
nand U975 (N_975,In_2423,In_1047);
and U976 (N_976,In_1384,In_2549);
and U977 (N_977,In_451,In_566);
xnor U978 (N_978,In_1090,In_1045);
xor U979 (N_979,In_639,In_492);
and U980 (N_980,In_2461,In_1551);
and U981 (N_981,In_2644,In_2569);
nand U982 (N_982,In_1582,In_104);
nand U983 (N_983,In_1369,In_342);
nor U984 (N_984,In_2094,In_1282);
or U985 (N_985,In_33,In_2862);
and U986 (N_986,In_2309,In_2482);
or U987 (N_987,In_1513,In_2104);
nand U988 (N_988,In_2469,In_1709);
nor U989 (N_989,In_1956,In_1310);
and U990 (N_990,In_2536,In_1493);
or U991 (N_991,In_474,In_2447);
nor U992 (N_992,In_1739,In_2502);
nor U993 (N_993,In_2537,In_1075);
nand U994 (N_994,In_145,In_2768);
nor U995 (N_995,In_2988,In_2899);
nand U996 (N_996,In_2360,In_1010);
or U997 (N_997,In_1062,In_2361);
nor U998 (N_998,In_2038,In_606);
and U999 (N_999,In_408,In_972);
and U1000 (N_1000,In_1442,In_272);
and U1001 (N_1001,In_1316,In_692);
or U1002 (N_1002,In_1155,In_64);
nor U1003 (N_1003,In_1012,In_1437);
and U1004 (N_1004,In_1194,In_735);
xnor U1005 (N_1005,In_730,In_2974);
nand U1006 (N_1006,In_1216,In_1037);
and U1007 (N_1007,In_2025,In_2499);
nand U1008 (N_1008,In_2947,In_2679);
nand U1009 (N_1009,In_2804,In_2262);
and U1010 (N_1010,In_1093,In_1175);
and U1011 (N_1011,In_1058,In_1127);
or U1012 (N_1012,In_845,In_1107);
xor U1013 (N_1013,In_1799,In_2390);
xnor U1014 (N_1014,In_2811,In_2686);
nor U1015 (N_1015,In_1614,In_908);
and U1016 (N_1016,In_2317,In_2583);
nor U1017 (N_1017,In_2218,In_215);
or U1018 (N_1018,In_2433,In_338);
xor U1019 (N_1019,In_309,In_1444);
nor U1020 (N_1020,In_2640,In_714);
xnor U1021 (N_1021,In_1906,In_1663);
nor U1022 (N_1022,In_1875,In_2455);
xnor U1023 (N_1023,In_2288,In_2933);
xor U1024 (N_1024,In_2252,In_2520);
xnor U1025 (N_1025,In_2980,In_746);
xor U1026 (N_1026,In_2483,In_1434);
and U1027 (N_1027,In_1501,In_2368);
and U1028 (N_1028,In_172,In_2348);
and U1029 (N_1029,In_211,In_1013);
and U1030 (N_1030,In_2297,In_94);
xnor U1031 (N_1031,In_1629,In_9);
and U1032 (N_1032,In_1623,In_2477);
nor U1033 (N_1033,In_156,In_2907);
nand U1034 (N_1034,In_2345,In_1223);
nand U1035 (N_1035,In_255,In_2200);
or U1036 (N_1036,In_2435,In_91);
and U1037 (N_1037,In_637,In_356);
xor U1038 (N_1038,In_2680,In_383);
or U1039 (N_1039,In_217,In_1450);
xor U1040 (N_1040,In_2534,In_934);
or U1041 (N_1041,In_2467,In_287);
nor U1042 (N_1042,In_2599,In_2934);
or U1043 (N_1043,In_316,In_1132);
or U1044 (N_1044,In_2051,In_68);
xnor U1045 (N_1045,In_893,In_369);
nand U1046 (N_1046,In_480,In_687);
and U1047 (N_1047,In_154,In_1790);
nand U1048 (N_1048,In_2792,In_2405);
nor U1049 (N_1049,In_196,In_2828);
nor U1050 (N_1050,In_184,In_1961);
or U1051 (N_1051,In_1990,In_1146);
and U1052 (N_1052,In_160,In_1301);
or U1053 (N_1053,In_1390,In_2157);
nand U1054 (N_1054,In_819,In_564);
xor U1055 (N_1055,In_2742,In_2319);
xor U1056 (N_1056,In_1524,In_8);
and U1057 (N_1057,In_1360,In_1533);
nor U1058 (N_1058,In_2445,In_1147);
and U1059 (N_1059,In_2831,In_1266);
nand U1060 (N_1060,In_1991,In_2553);
and U1061 (N_1061,In_370,In_452);
nor U1062 (N_1062,In_2968,In_405);
or U1063 (N_1063,In_1871,In_1932);
nor U1064 (N_1064,In_2765,In_1881);
and U1065 (N_1065,In_1653,In_1105);
or U1066 (N_1066,In_1835,In_2130);
nand U1067 (N_1067,In_2615,In_2715);
xnor U1068 (N_1068,In_891,In_2032);
or U1069 (N_1069,In_0,In_65);
or U1070 (N_1070,In_1153,In_81);
nor U1071 (N_1071,In_2786,In_2269);
xnor U1072 (N_1072,In_1791,In_59);
xnor U1073 (N_1073,In_643,In_2112);
nor U1074 (N_1074,In_1568,In_2790);
nand U1075 (N_1075,In_36,In_1239);
or U1076 (N_1076,In_228,In_2976);
or U1077 (N_1077,In_1697,In_2830);
or U1078 (N_1078,In_1288,In_1547);
nand U1079 (N_1079,In_1686,In_713);
or U1080 (N_1080,In_2180,In_1912);
xnor U1081 (N_1081,In_1404,In_1528);
and U1082 (N_1082,In_201,In_2255);
nor U1083 (N_1083,In_1607,In_1674);
or U1084 (N_1084,In_1857,In_1286);
xnor U1085 (N_1085,In_1649,In_2543);
and U1086 (N_1086,In_1578,In_1704);
xnor U1087 (N_1087,In_2781,In_662);
nand U1088 (N_1088,In_2880,In_675);
and U1089 (N_1089,In_209,In_58);
xor U1090 (N_1090,In_1169,In_2870);
or U1091 (N_1091,In_509,In_2550);
nand U1092 (N_1092,In_743,In_263);
or U1093 (N_1093,In_1848,In_45);
nand U1094 (N_1094,In_657,In_114);
nor U1095 (N_1095,In_2284,In_23);
xnor U1096 (N_1096,In_2358,In_1429);
or U1097 (N_1097,In_3,In_1661);
and U1098 (N_1098,In_479,In_1707);
nand U1099 (N_1099,In_1830,In_1724);
or U1100 (N_1100,In_2950,In_808);
nor U1101 (N_1101,In_2178,In_1423);
and U1102 (N_1102,In_1064,In_1015);
nand U1103 (N_1103,In_219,In_2321);
and U1104 (N_1104,In_817,In_119);
xor U1105 (N_1105,In_793,In_995);
and U1106 (N_1106,In_1068,In_1583);
nand U1107 (N_1107,In_339,In_1968);
nand U1108 (N_1108,In_230,In_1299);
or U1109 (N_1109,In_2225,In_2738);
xnor U1110 (N_1110,In_1684,In_764);
nand U1111 (N_1111,In_1530,In_1659);
nor U1112 (N_1112,In_2377,In_2233);
nand U1113 (N_1113,In_1489,In_888);
nor U1114 (N_1114,In_1017,In_1124);
xor U1115 (N_1115,In_105,In_1742);
nor U1116 (N_1116,In_576,In_554);
nor U1117 (N_1117,In_586,In_1082);
or U1118 (N_1118,In_387,In_1469);
nand U1119 (N_1119,In_683,In_2879);
nand U1120 (N_1120,In_1391,In_2207);
or U1121 (N_1121,In_2143,In_1590);
nor U1122 (N_1122,In_2842,In_50);
nand U1123 (N_1123,In_1801,In_921);
xnor U1124 (N_1124,In_1492,In_2228);
nand U1125 (N_1125,In_133,In_1312);
and U1126 (N_1126,In_867,In_69);
xnor U1127 (N_1127,In_765,In_267);
nand U1128 (N_1128,In_2400,In_572);
or U1129 (N_1129,In_2521,In_804);
nand U1130 (N_1130,In_1593,In_1098);
xor U1131 (N_1131,In_1471,In_1213);
nand U1132 (N_1132,In_1950,In_1581);
and U1133 (N_1133,In_1564,In_1087);
nand U1134 (N_1134,In_2832,In_2927);
nand U1135 (N_1135,In_2967,In_2858);
or U1136 (N_1136,In_233,In_644);
nand U1137 (N_1137,In_389,In_1503);
nor U1138 (N_1138,In_213,In_502);
xor U1139 (N_1139,In_256,In_2017);
nand U1140 (N_1140,In_1331,In_432);
nand U1141 (N_1141,In_724,In_1199);
nor U1142 (N_1142,In_1428,In_2150);
nor U1143 (N_1143,In_1563,In_1001);
nand U1144 (N_1144,In_526,In_807);
and U1145 (N_1145,In_2307,In_2653);
nor U1146 (N_1146,In_2977,In_1362);
nor U1147 (N_1147,In_599,In_2629);
xnor U1148 (N_1148,In_447,In_716);
and U1149 (N_1149,In_2396,In_2084);
nand U1150 (N_1150,In_920,In_2722);
nor U1151 (N_1151,In_768,In_992);
xnor U1152 (N_1152,In_2905,In_1747);
or U1153 (N_1153,In_1257,In_1173);
nor U1154 (N_1154,In_774,In_1053);
nand U1155 (N_1155,In_1996,In_2506);
nor U1156 (N_1156,In_1329,In_2033);
nand U1157 (N_1157,In_1812,In_1566);
nand U1158 (N_1158,In_1514,In_1795);
nor U1159 (N_1159,In_2311,In_67);
or U1160 (N_1160,In_227,In_1388);
or U1161 (N_1161,In_1426,In_2406);
and U1162 (N_1162,In_975,In_392);
or U1163 (N_1163,In_2478,In_949);
nor U1164 (N_1164,In_2354,In_833);
nand U1165 (N_1165,In_2190,In_4);
and U1166 (N_1166,In_1416,In_1072);
nand U1167 (N_1167,In_702,In_835);
or U1168 (N_1168,In_434,In_1381);
nand U1169 (N_1169,In_997,In_88);
xnor U1170 (N_1170,In_2314,In_1515);
and U1171 (N_1171,In_855,In_2808);
xnor U1172 (N_1172,In_960,In_1052);
nor U1173 (N_1173,In_1494,In_162);
nand U1174 (N_1174,In_2329,In_2444);
or U1175 (N_1175,In_1397,In_1844);
and U1176 (N_1176,In_191,In_258);
xnor U1177 (N_1177,In_2073,In_2191);
nand U1178 (N_1178,In_2456,In_597);
and U1179 (N_1179,In_2777,In_2625);
and U1180 (N_1180,In_1427,In_1079);
or U1181 (N_1181,In_99,In_2841);
nand U1182 (N_1182,In_2324,In_1453);
nor U1183 (N_1183,In_2589,In_2008);
nor U1184 (N_1184,In_1690,In_310);
and U1185 (N_1185,In_2250,In_1215);
and U1186 (N_1186,In_2523,In_2356);
or U1187 (N_1187,In_2030,In_2350);
nand U1188 (N_1188,In_1941,In_428);
and U1189 (N_1189,In_875,In_2257);
xnor U1190 (N_1190,In_2142,In_2651);
and U1191 (N_1191,In_2593,In_1873);
or U1192 (N_1192,In_2529,In_2376);
nor U1193 (N_1193,In_982,In_2295);
xnor U1194 (N_1194,In_2292,In_1188);
and U1195 (N_1195,In_2158,In_1771);
or U1196 (N_1196,In_25,In_1636);
nor U1197 (N_1197,In_987,In_847);
and U1198 (N_1198,In_1817,In_2388);
nor U1199 (N_1199,In_1644,In_2217);
and U1200 (N_1200,In_2054,In_1143);
or U1201 (N_1201,In_2918,In_329);
xnor U1202 (N_1202,N_752,N_767);
xnor U1203 (N_1203,In_2242,N_454);
and U1204 (N_1204,N_80,In_1622);
nor U1205 (N_1205,N_535,N_1199);
xor U1206 (N_1206,N_1129,N_671);
xnor U1207 (N_1207,N_1007,N_377);
xnor U1208 (N_1208,In_2155,N_97);
xor U1209 (N_1209,In_2799,N_860);
and U1210 (N_1210,N_229,In_281);
or U1211 (N_1211,In_2630,N_825);
nor U1212 (N_1212,N_904,N_367);
nand U1213 (N_1213,N_762,N_73);
or U1214 (N_1214,N_909,N_159);
or U1215 (N_1215,N_326,N_571);
or U1216 (N_1216,N_1137,N_996);
and U1217 (N_1217,N_414,N_296);
xor U1218 (N_1218,N_255,In_1328);
xnor U1219 (N_1219,N_483,N_288);
xnor U1220 (N_1220,In_2824,N_415);
nor U1221 (N_1221,In_770,In_1160);
or U1222 (N_1222,N_526,In_165);
or U1223 (N_1223,N_176,In_2540);
nor U1224 (N_1224,In_525,N_654);
nand U1225 (N_1225,N_943,N_200);
or U1226 (N_1226,In_1351,N_1093);
or U1227 (N_1227,N_406,N_515);
and U1228 (N_1228,N_1172,In_994);
nand U1229 (N_1229,In_2430,N_647);
nor U1230 (N_1230,In_754,In_102);
xnor U1231 (N_1231,N_625,In_1665);
nand U1232 (N_1232,In_803,In_999);
and U1233 (N_1233,In_1355,N_351);
or U1234 (N_1234,N_811,N_826);
nor U1235 (N_1235,N_1110,N_379);
nor U1236 (N_1236,N_540,N_114);
or U1237 (N_1237,In_57,In_1893);
and U1238 (N_1238,In_373,N_1098);
xor U1239 (N_1239,In_1694,N_452);
and U1240 (N_1240,N_589,N_1049);
and U1241 (N_1241,N_590,N_286);
nand U1242 (N_1242,N_852,N_1009);
or U1243 (N_1243,N_257,N_1083);
nor U1244 (N_1244,N_18,N_431);
and U1245 (N_1245,In_1825,N_47);
xor U1246 (N_1246,N_541,N_471);
and U1247 (N_1247,In_282,In_379);
nand U1248 (N_1248,N_57,N_8);
xnor U1249 (N_1249,N_350,In_1411);
nor U1250 (N_1250,N_1107,N_993);
xnor U1251 (N_1251,N_599,N_256);
nand U1252 (N_1252,N_834,N_906);
nand U1253 (N_1253,N_591,N_1178);
and U1254 (N_1254,N_892,N_472);
and U1255 (N_1255,N_933,In_2335);
nand U1256 (N_1256,N_1136,N_485);
xnor U1257 (N_1257,N_888,N_1025);
and U1258 (N_1258,N_658,N_87);
and U1259 (N_1259,In_374,N_84);
nand U1260 (N_1260,In_2683,In_740);
nand U1261 (N_1261,In_612,In_1018);
xnor U1262 (N_1262,N_1052,In_1069);
or U1263 (N_1263,In_7,N_1169);
xnor U1264 (N_1264,In_1458,In_1943);
nand U1265 (N_1265,In_158,N_10);
or U1266 (N_1266,N_653,N_287);
or U1267 (N_1267,N_500,N_323);
and U1268 (N_1268,N_44,N_468);
or U1269 (N_1269,In_536,N_481);
or U1270 (N_1270,N_167,In_1611);
xnor U1271 (N_1271,In_2923,N_467);
nor U1272 (N_1272,N_1029,N_704);
nand U1273 (N_1273,N_1051,In_2049);
xnor U1274 (N_1274,N_181,N_126);
or U1275 (N_1275,N_853,N_1134);
nor U1276 (N_1276,N_1033,N_355);
or U1277 (N_1277,N_1166,In_844);
nand U1278 (N_1278,N_789,In_1473);
nand U1279 (N_1279,N_558,N_746);
xor U1280 (N_1280,N_724,N_840);
or U1281 (N_1281,N_609,In_1553);
nor U1282 (N_1282,N_979,N_1118);
xor U1283 (N_1283,N_1112,In_1177);
nor U1284 (N_1284,In_1733,N_1053);
xor U1285 (N_1285,N_315,N_461);
and U1286 (N_1286,N_1070,In_2855);
xor U1287 (N_1287,N_1159,N_263);
nor U1288 (N_1288,N_1092,In_1508);
xor U1289 (N_1289,N_1075,N_512);
and U1290 (N_1290,N_645,In_2261);
xnor U1291 (N_1291,In_2304,In_488);
xor U1292 (N_1292,N_1151,In_293);
and U1293 (N_1293,N_771,In_1096);
nand U1294 (N_1294,In_2193,N_196);
and U1295 (N_1295,In_2171,In_175);
xnor U1296 (N_1296,In_988,N_1091);
and U1297 (N_1297,N_808,In_1969);
or U1298 (N_1298,In_601,N_1082);
or U1299 (N_1299,N_82,N_1050);
nand U1300 (N_1300,In_1470,In_378);
or U1301 (N_1301,In_2707,N_1063);
nor U1302 (N_1302,N_968,N_1040);
nor U1303 (N_1303,In_487,N_211);
and U1304 (N_1304,N_534,N_38);
and U1305 (N_1305,In_2395,In_442);
or U1306 (N_1306,N_562,N_1103);
nand U1307 (N_1307,In_1185,N_103);
xor U1308 (N_1308,In_617,N_854);
or U1309 (N_1309,N_513,N_554);
or U1310 (N_1310,N_508,N_498);
and U1311 (N_1311,N_880,N_225);
nand U1312 (N_1312,N_646,N_169);
nor U1313 (N_1313,In_142,N_894);
or U1314 (N_1314,In_351,N_26);
and U1315 (N_1315,N_837,In_659);
xor U1316 (N_1316,N_223,In_2497);
nor U1317 (N_1317,N_958,N_506);
nor U1318 (N_1318,N_172,N_597);
or U1319 (N_1319,N_856,In_1343);
xnor U1320 (N_1320,N_69,N_816);
nor U1321 (N_1321,N_876,N_605);
and U1322 (N_1322,In_1184,N_594);
nand U1323 (N_1323,In_2289,N_191);
or U1324 (N_1324,In_164,In_1198);
nor U1325 (N_1325,N_1068,N_595);
and U1326 (N_1326,N_798,In_965);
and U1327 (N_1327,In_680,N_37);
nand U1328 (N_1328,In_1654,N_676);
xor U1329 (N_1329,N_819,In_1352);
or U1330 (N_1330,N_710,N_313);
nor U1331 (N_1331,N_136,N_1047);
and U1332 (N_1332,In_2014,In_2901);
nor U1333 (N_1333,N_1000,In_2609);
nor U1334 (N_1334,N_733,N_1004);
or U1335 (N_1335,In_2928,In_2681);
xnor U1336 (N_1336,In_1761,In_973);
xor U1337 (N_1337,In_1519,N_1109);
xnor U1338 (N_1338,N_1175,N_316);
nor U1339 (N_1339,In_2989,N_930);
nor U1340 (N_1340,N_320,N_662);
nor U1341 (N_1341,N_375,N_953);
xnor U1342 (N_1342,In_715,N_664);
nor U1343 (N_1343,In_482,In_1333);
or U1344 (N_1344,N_488,N_984);
nor U1345 (N_1345,N_1189,In_812);
xor U1346 (N_1346,N_1141,N_543);
xor U1347 (N_1347,In_2323,In_1753);
nor U1348 (N_1348,In_2210,N_680);
or U1349 (N_1349,N_862,In_244);
and U1350 (N_1350,N_600,N_173);
nor U1351 (N_1351,N_764,N_754);
nand U1352 (N_1352,N_152,N_24);
xor U1353 (N_1353,N_232,In_2248);
and U1354 (N_1354,N_521,In_1076);
and U1355 (N_1355,In_2199,N_6);
and U1356 (N_1356,N_602,N_629);
nand U1357 (N_1357,N_549,N_946);
or U1358 (N_1358,N_1128,In_2392);
or U1359 (N_1359,N_180,N_1061);
nand U1360 (N_1360,In_380,N_245);
and U1361 (N_1361,N_681,In_475);
and U1362 (N_1362,In_767,In_1748);
and U1363 (N_1363,N_584,N_991);
and U1364 (N_1364,N_357,In_407);
xnor U1365 (N_1365,N_1187,N_705);
or U1366 (N_1366,N_519,N_759);
and U1367 (N_1367,N_1184,In_1527);
or U1368 (N_1368,N_130,In_2016);
nor U1369 (N_1369,N_732,N_843);
nor U1370 (N_1370,In_1183,N_858);
nand U1371 (N_1371,N_941,N_944);
nand U1372 (N_1372,In_831,N_969);
nand U1373 (N_1373,N_353,N_766);
and U1374 (N_1374,In_1433,N_966);
nand U1375 (N_1375,In_2802,N_271);
xor U1376 (N_1376,N_348,In_2067);
nor U1377 (N_1377,N_349,N_182);
or U1378 (N_1378,N_456,N_134);
or U1379 (N_1379,In_349,N_687);
nor U1380 (N_1380,N_661,N_812);
nand U1381 (N_1381,In_1898,In_2327);
nand U1382 (N_1382,N_141,N_694);
and U1383 (N_1383,In_377,N_450);
or U1384 (N_1384,N_273,N_20);
nor U1385 (N_1385,In_1151,N_883);
and U1386 (N_1386,In_1878,N_157);
nand U1387 (N_1387,In_640,In_2463);
and U1388 (N_1388,N_921,In_2564);
nand U1389 (N_1389,In_842,N_105);
nand U1390 (N_1390,N_463,N_544);
nand U1391 (N_1391,N_153,N_289);
or U1392 (N_1392,N_1124,N_408);
or U1393 (N_1393,N_612,N_552);
nor U1394 (N_1394,N_846,N_457);
xnor U1395 (N_1395,N_462,N_1146);
xnor U1396 (N_1396,In_1235,N_40);
xnor U1397 (N_1397,N_990,In_1635);
xnor U1398 (N_1398,N_765,In_2474);
or U1399 (N_1399,N_935,N_435);
or U1400 (N_1400,N_305,N_28);
nand U1401 (N_1401,In_2256,In_1696);
and U1402 (N_1402,In_2911,In_1024);
and U1403 (N_1403,N_804,In_1948);
xor U1404 (N_1404,In_1313,In_1309);
xor U1405 (N_1405,In_1560,In_1918);
nand U1406 (N_1406,In_989,In_1121);
or U1407 (N_1407,N_555,In_2856);
nand U1408 (N_1408,In_1586,In_1399);
xor U1409 (N_1409,N_1104,N_494);
nand U1410 (N_1410,N_1085,N_884);
nand U1411 (N_1411,N_529,N_77);
nor U1412 (N_1412,In_265,N_268);
and U1413 (N_1413,N_717,In_397);
and U1414 (N_1414,N_1023,N_301);
xnor U1415 (N_1415,N_486,N_1086);
and U1416 (N_1416,N_567,N_324);
or U1417 (N_1417,In_2427,N_797);
nand U1418 (N_1418,N_306,N_5);
nand U1419 (N_1419,N_685,N_407);
nor U1420 (N_1420,N_748,In_446);
xor U1421 (N_1421,In_222,N_363);
xor U1422 (N_1422,N_618,N_405);
xnor U1423 (N_1423,N_32,In_2365);
or U1424 (N_1424,N_455,N_1008);
nor U1425 (N_1425,N_331,N_234);
or U1426 (N_1426,In_180,N_942);
nor U1427 (N_1427,N_518,N_885);
and U1428 (N_1428,In_386,In_2253);
nand U1429 (N_1429,In_1484,N_859);
or U1430 (N_1430,In_1541,N_1001);
nand U1431 (N_1431,In_967,N_882);
nand U1432 (N_1432,N_818,N_1080);
nand U1433 (N_1433,N_135,N_1044);
xnor U1434 (N_1434,N_1019,N_1142);
xnor U1435 (N_1435,N_311,In_1957);
and U1436 (N_1436,In_654,N_806);
nor U1437 (N_1437,In_249,In_936);
nand U1438 (N_1438,N_249,N_158);
nand U1439 (N_1439,N_31,In_593);
or U1440 (N_1440,N_250,In_15);
xnor U1441 (N_1441,In_1221,N_980);
xnor U1442 (N_1442,N_424,In_2994);
and U1443 (N_1443,N_615,N_436);
xnor U1444 (N_1444,N_835,In_1792);
xor U1445 (N_1445,N_91,N_243);
and U1446 (N_1446,N_445,In_533);
nand U1447 (N_1447,In_311,In_2119);
and U1448 (N_1448,N_1096,N_994);
nand U1449 (N_1449,N_616,N_160);
nor U1450 (N_1450,N_395,N_108);
and U1451 (N_1451,In_1441,In_2751);
xnor U1452 (N_1452,N_439,In_2195);
and U1453 (N_1453,N_235,N_659);
nor U1454 (N_1454,In_205,N_666);
and U1455 (N_1455,N_688,N_538);
and U1456 (N_1456,N_769,N_801);
xor U1457 (N_1457,In_2077,N_546);
nand U1458 (N_1458,In_892,N_224);
or U1459 (N_1459,N_761,N_774);
nor U1460 (N_1460,N_213,N_50);
and U1461 (N_1461,N_723,N_272);
and U1462 (N_1462,N_588,N_1161);
xnor U1463 (N_1463,N_110,N_985);
nand U1464 (N_1464,N_233,N_100);
nand U1465 (N_1465,N_1002,N_66);
nor U1466 (N_1466,N_547,N_1090);
nand U1467 (N_1467,In_1509,N_226);
and U1468 (N_1468,N_1,In_429);
nor U1469 (N_1469,N_497,N_1116);
nor U1470 (N_1470,N_1193,In_2050);
xnor U1471 (N_1471,N_1185,N_112);
nand U1472 (N_1472,N_568,N_1022);
and U1473 (N_1473,In_2334,N_280);
and U1474 (N_1474,N_260,In_260);
nor U1475 (N_1475,N_347,N_115);
or U1476 (N_1476,N_604,N_365);
nand U1477 (N_1477,N_30,In_2275);
nand U1478 (N_1478,N_987,N_218);
and U1479 (N_1479,N_511,N_881);
and U1480 (N_1480,N_490,In_613);
and U1481 (N_1481,N_76,In_2093);
or U1482 (N_1482,N_800,N_45);
or U1483 (N_1483,In_756,N_889);
nand U1484 (N_1484,N_718,N_121);
xnor U1485 (N_1485,N_416,In_535);
nor U1486 (N_1486,In_2211,In_1879);
xnor U1487 (N_1487,N_83,N_1191);
xor U1488 (N_1488,N_330,N_1062);
or U1489 (N_1489,In_2998,N_1084);
nand U1490 (N_1490,N_703,N_274);
or U1491 (N_1491,N_1117,In_1810);
nor U1492 (N_1492,N_848,In_814);
nand U1493 (N_1493,N_709,In_1867);
and U1494 (N_1494,N_502,In_335);
nor U1495 (N_1495,N_212,N_1064);
or U1496 (N_1496,In_1456,In_390);
xor U1497 (N_1497,N_624,In_530);
xnor U1498 (N_1498,In_2299,N_751);
or U1499 (N_1499,In_1518,N_553);
and U1500 (N_1500,N_784,N_504);
nor U1501 (N_1501,N_864,N_1194);
and U1502 (N_1502,In_689,In_1174);
xnor U1503 (N_1503,N_891,N_29);
and U1504 (N_1504,N_517,In_1960);
nand U1505 (N_1505,N_695,N_781);
and U1506 (N_1506,N_36,In_1449);
nand U1507 (N_1507,N_672,In_1122);
nor U1508 (N_1508,In_2373,N_1030);
nand U1509 (N_1509,N_35,N_61);
xor U1510 (N_1510,N_566,N_251);
nor U1511 (N_1511,N_1015,N_865);
xor U1512 (N_1512,N_1190,In_585);
nor U1513 (N_1513,In_2415,In_2563);
or U1514 (N_1514,In_1407,In_1942);
and U1515 (N_1515,In_2696,N_533);
and U1516 (N_1516,N_1171,In_1304);
and U1517 (N_1517,N_787,N_707);
nand U1518 (N_1518,In_2509,N_139);
nand U1519 (N_1519,N_19,N_98);
or U1520 (N_1520,N_220,N_940);
nor U1521 (N_1521,N_1160,N_479);
or U1522 (N_1522,N_841,N_1163);
xnor U1523 (N_1523,N_81,N_1066);
nor U1524 (N_1524,N_537,N_824);
and U1525 (N_1525,N_175,N_815);
and U1526 (N_1526,In_2251,N_39);
nand U1527 (N_1527,In_2747,N_284);
xor U1528 (N_1528,N_404,In_1703);
xor U1529 (N_1529,In_435,N_188);
or U1530 (N_1530,In_1394,In_334);
xor U1531 (N_1531,N_992,N_559);
and U1532 (N_1532,In_2693,N_974);
and U1533 (N_1533,N_146,N_148);
nor U1534 (N_1534,N_1125,In_1398);
and U1535 (N_1535,N_302,N_633);
nand U1536 (N_1536,In_2136,N_934);
and U1537 (N_1537,N_1088,In_1073);
xnor U1538 (N_1538,N_631,In_1546);
xor U1539 (N_1539,In_1870,N_190);
nand U1540 (N_1540,In_300,N_950);
nand U1541 (N_1541,In_1785,N_627);
nor U1542 (N_1542,N_247,In_2068);
or U1543 (N_1543,In_2952,N_1034);
nor U1544 (N_1544,In_2539,N_763);
nor U1545 (N_1545,N_949,In_1637);
or U1546 (N_1546,In_2285,N_434);
nor U1547 (N_1547,In_1336,N_238);
nand U1548 (N_1548,N_677,In_1695);
or U1549 (N_1549,In_420,N_1148);
nor U1550 (N_1550,In_1613,N_899);
or U1551 (N_1551,In_2809,In_2095);
or U1552 (N_1552,N_199,In_1909);
and U1553 (N_1553,N_923,N_667);
and U1554 (N_1554,N_779,In_1664);
xor U1555 (N_1555,In_2789,N_851);
nand U1556 (N_1556,N_453,In_697);
xnor U1557 (N_1557,N_959,In_2226);
nand U1558 (N_1558,In_1302,In_1206);
xnor U1559 (N_1559,N_530,In_2409);
xnor U1560 (N_1560,N_1024,N_592);
xor U1561 (N_1561,In_1403,N_204);
nand U1562 (N_1562,N_374,N_845);
nor U1563 (N_1563,N_768,In_1305);
or U1564 (N_1564,In_2836,N_527);
and U1565 (N_1565,N_509,N_17);
and U1566 (N_1566,In_2618,N_364);
and U1567 (N_1567,In_584,N_722);
nor U1568 (N_1568,N_670,N_161);
xnor U1569 (N_1569,N_1188,N_187);
or U1570 (N_1570,N_371,N_14);
nand U1571 (N_1571,In_2760,N_593);
xor U1572 (N_1572,In_1026,In_313);
or U1573 (N_1573,N_282,In_732);
or U1574 (N_1574,In_278,N_961);
or U1575 (N_1575,N_1017,N_425);
and U1576 (N_1576,In_2711,In_2847);
or U1577 (N_1577,N_397,N_596);
and U1578 (N_1578,In_2383,N_43);
and U1579 (N_1579,In_2634,In_1485);
nand U1580 (N_1580,N_67,In_2530);
xor U1581 (N_1581,In_2556,N_952);
and U1582 (N_1582,In_204,In_1641);
xnor U1583 (N_1583,In_895,In_753);
or U1584 (N_1584,In_2419,N_392);
or U1585 (N_1585,In_1154,In_1378);
nor U1586 (N_1586,N_236,N_1162);
nor U1587 (N_1587,N_1195,In_852);
nand U1588 (N_1588,N_913,N_398);
nor U1589 (N_1589,N_116,In_1273);
xor U1590 (N_1590,N_310,N_258);
xnor U1591 (N_1591,N_897,In_2097);
or U1592 (N_1592,N_409,N_487);
xor U1593 (N_1593,N_1197,N_470);
xor U1594 (N_1594,In_943,In_1643);
or U1595 (N_1595,N_356,N_63);
nand U1596 (N_1596,In_2724,N_1144);
or U1597 (N_1597,N_342,N_531);
xor U1598 (N_1598,In_2243,N_1170);
and U1599 (N_1599,In_358,In_2310);
nand U1600 (N_1600,N_810,N_59);
and U1601 (N_1601,N_747,N_214);
nand U1602 (N_1602,N_607,In_152);
nand U1603 (N_1603,N_563,In_854);
nor U1604 (N_1604,N_154,N_839);
xnor U1605 (N_1605,In_699,N_386);
or U1606 (N_1606,In_246,N_241);
and U1607 (N_1607,N_970,N_396);
and U1608 (N_1608,N_140,N_292);
xor U1609 (N_1609,In_2887,N_118);
xnor U1610 (N_1610,N_739,N_370);
nand U1611 (N_1611,N_278,N_640);
nor U1612 (N_1612,N_684,N_1069);
nor U1613 (N_1613,N_70,In_2603);
xnor U1614 (N_1614,N_283,In_1619);
and U1615 (N_1615,N_64,N_1039);
or U1616 (N_1616,N_651,N_890);
nand U1617 (N_1617,N_432,N_699);
or U1618 (N_1618,In_642,N_520);
nand U1619 (N_1619,In_1276,N_753);
xnor U1620 (N_1620,N_586,N_16);
xnor U1621 (N_1621,N_1005,N_642);
nor U1622 (N_1622,N_964,N_814);
nor U1623 (N_1623,N_623,N_514);
xor U1624 (N_1624,N_1003,N_601);
or U1625 (N_1625,N_21,N_354);
nor U1626 (N_1626,N_649,N_261);
and U1627 (N_1627,In_2984,N_491);
and U1628 (N_1628,In_1421,N_911);
and U1629 (N_1629,N_90,N_579);
nand U1630 (N_1630,In_78,N_72);
xnor U1631 (N_1631,N_185,In_962);
nand U1632 (N_1632,In_1392,N_465);
xnor U1633 (N_1633,In_538,In_2110);
or U1634 (N_1634,N_49,In_321);
nand U1635 (N_1635,N_300,N_828);
or U1636 (N_1636,In_19,In_1984);
nand U1637 (N_1637,N_231,In_375);
or U1638 (N_1638,N_573,N_428);
and U1639 (N_1639,N_79,N_847);
and U1640 (N_1640,N_986,N_878);
nand U1641 (N_1641,In_2518,N_1156);
nand U1642 (N_1642,In_1570,N_252);
xnor U1643 (N_1643,In_939,N_477);
nand U1644 (N_1644,In_907,N_209);
xnor U1645 (N_1645,In_2313,N_113);
xnor U1646 (N_1646,N_696,N_227);
nor U1647 (N_1647,In_1376,N_440);
nand U1648 (N_1648,N_830,N_574);
or U1649 (N_1649,N_850,N_27);
and U1650 (N_1650,N_576,In_2413);
and U1651 (N_1651,In_2154,N_259);
nor U1652 (N_1652,N_708,N_427);
and U1653 (N_1653,In_499,N_9);
or U1654 (N_1654,In_2601,N_1114);
nand U1655 (N_1655,N_606,N_429);
xor U1656 (N_1656,N_1115,In_266);
nand U1657 (N_1657,N_962,N_25);
nand U1658 (N_1658,N_171,N_855);
and U1659 (N_1659,N_603,N_908);
nor U1660 (N_1660,N_99,In_863);
nor U1661 (N_1661,N_1155,In_2697);
xor U1662 (N_1662,N_93,In_2458);
nor U1663 (N_1663,In_587,In_29);
xor U1664 (N_1664,In_2227,In_2037);
xor U1665 (N_1665,In_2318,N_879);
and U1666 (N_1666,N_721,In_1499);
or U1667 (N_1667,In_2182,N_793);
nor U1668 (N_1668,N_101,N_2);
or U1669 (N_1669,In_1074,N_926);
nand U1670 (N_1670,N_734,N_679);
xor U1671 (N_1671,N_86,N_715);
xnor U1672 (N_1672,N_956,In_910);
nor U1673 (N_1673,N_1164,N_23);
nand U1674 (N_1674,In_2475,N_403);
nor U1675 (N_1675,In_2005,In_1255);
and U1676 (N_1676,N_1089,In_2046);
and U1677 (N_1677,N_981,N_332);
xnor U1678 (N_1678,N_307,N_1072);
xor U1679 (N_1679,N_291,N_920);
xor U1680 (N_1680,N_1102,In_2891);
xnor U1681 (N_1681,N_202,In_2754);
nor U1682 (N_1682,N_96,N_189);
xnor U1683 (N_1683,In_2223,N_611);
and U1684 (N_1684,N_372,N_179);
or U1685 (N_1685,N_524,N_277);
xor U1686 (N_1686,N_106,N_270);
xnor U1687 (N_1687,N_637,N_442);
or U1688 (N_1688,N_760,N_413);
and U1689 (N_1689,In_168,In_1468);
xor U1690 (N_1690,N_901,In_2015);
nand U1691 (N_1691,N_1046,In_367);
nor U1692 (N_1692,In_532,N_484);
or U1693 (N_1693,N_720,N_177);
nor U1694 (N_1694,In_520,In_2450);
or U1695 (N_1695,In_2184,N_849);
or U1696 (N_1696,N_780,N_777);
or U1697 (N_1697,In_2001,N_683);
and U1698 (N_1698,In_2588,N_285);
and U1699 (N_1699,N_635,N_237);
nand U1700 (N_1700,N_965,N_207);
or U1701 (N_1701,N_776,In_108);
xor U1702 (N_1702,In_1006,N_1076);
nand U1703 (N_1703,N_458,N_314);
and U1704 (N_1704,N_165,In_2767);
xor U1705 (N_1705,N_129,N_669);
nand U1706 (N_1706,N_874,N_866);
or U1707 (N_1707,In_1150,In_1529);
or U1708 (N_1708,N_560,N_1018);
nand U1709 (N_1709,N_496,In_1640);
and U1710 (N_1710,In_2867,In_762);
nand U1711 (N_1711,In_2893,N_33);
or U1712 (N_1712,In_2331,N_1147);
or U1713 (N_1713,N_1174,In_1952);
nand U1714 (N_1714,N_51,In_1510);
and U1715 (N_1715,N_466,N_937);
xor U1716 (N_1716,N_239,N_652);
or U1717 (N_1717,N_735,N_210);
nand U1718 (N_1718,N_523,N_975);
nor U1719 (N_1719,N_575,N_829);
and U1720 (N_1720,In_681,N_711);
and U1721 (N_1721,In_245,In_2759);
xor U1722 (N_1722,In_1091,In_2402);
nor U1723 (N_1723,N_628,In_1917);
nor U1724 (N_1724,In_2576,N_932);
nand U1725 (N_1725,N_702,In_2845);
nand U1726 (N_1726,In_270,N_1042);
nand U1727 (N_1727,In_2819,N_56);
nand U1728 (N_1728,N_1074,In_2055);
xnor U1729 (N_1729,N_137,N_634);
xor U1730 (N_1730,N_570,N_556);
or U1731 (N_1731,N_580,In_2451);
nor U1732 (N_1732,N_648,N_938);
nor U1733 (N_1733,In_2387,N_755);
nand U1734 (N_1734,N_916,In_1466);
xor U1735 (N_1735,N_75,N_978);
nor U1736 (N_1736,N_464,N_1126);
xnor U1737 (N_1737,In_2848,N_170);
nor U1738 (N_1738,N_308,In_1245);
or U1739 (N_1739,In_2131,N_1127);
nand U1740 (N_1740,N_1054,In_346);
nand U1741 (N_1741,N_786,N_630);
or U1742 (N_1742,N_674,In_13);
or U1743 (N_1743,In_2000,N_905);
and U1744 (N_1744,N_503,N_1183);
nor U1745 (N_1745,In_1615,In_1204);
xnor U1746 (N_1746,In_851,N_896);
and U1747 (N_1747,N_626,N_557);
nor U1748 (N_1748,N_319,In_514);
and U1749 (N_1749,In_2854,In_1465);
nand U1750 (N_1750,N_639,N_322);
and U1751 (N_1751,N_729,In_2703);
or U1752 (N_1752,N_1037,N_474);
and U1753 (N_1753,In_2170,N_820);
nor U1754 (N_1754,N_12,In_757);
and U1755 (N_1755,N_168,In_1241);
and U1756 (N_1756,In_79,N_682);
and U1757 (N_1757,N_418,N_1020);
nand U1758 (N_1758,N_700,In_2562);
xor U1759 (N_1759,N_931,In_1545);
xnor U1760 (N_1760,N_1014,In_898);
nand U1761 (N_1761,N_119,N_632);
and U1762 (N_1762,N_821,In_315);
nand U1763 (N_1763,N_1111,N_873);
nor U1764 (N_1764,N_620,N_727);
nor U1765 (N_1765,N_714,N_657);
xor U1766 (N_1766,N_358,N_936);
and U1767 (N_1767,In_2761,N_736);
or U1768 (N_1768,In_2290,In_98);
or U1769 (N_1769,N_510,In_2676);
xor U1770 (N_1770,In_971,N_1176);
xor U1771 (N_1771,N_1060,N_796);
nor U1772 (N_1772,In_2580,N_336);
nand U1773 (N_1773,N_133,N_731);
nand U1774 (N_1774,N_1071,N_833);
and U1775 (N_1775,N_156,N_262);
xor U1776 (N_1776,N_216,In_1626);
nand U1777 (N_1777,N_893,In_581);
and U1778 (N_1778,N_423,In_1358);
or U1779 (N_1779,N_741,N_802);
or U1780 (N_1780,In_1240,N_1087);
xor U1781 (N_1781,In_1680,In_1746);
xnor U1782 (N_1782,N_836,N_421);
nor U1783 (N_1783,In_998,N_144);
xnor U1784 (N_1784,N_872,N_329);
or U1785 (N_1785,N_1013,N_988);
or U1786 (N_1786,N_823,N_528);
xnor U1787 (N_1787,N_1106,N_143);
nand U1788 (N_1788,N_782,N_373);
nand U1789 (N_1789,In_2987,N_963);
nand U1790 (N_1790,In_1210,In_541);
nor U1791 (N_1791,N_972,N_745);
xor U1792 (N_1792,N_346,N_1135);
or U1793 (N_1793,N_1140,In_2342);
xor U1794 (N_1794,In_1726,N_1152);
and U1795 (N_1795,N_242,N_730);
nor U1796 (N_1796,In_2890,N_857);
nor U1797 (N_1797,N_107,N_1145);
nor U1798 (N_1798,N_132,In_1144);
xor U1799 (N_1799,N_973,N_459);
and U1800 (N_1800,In_2144,In_698);
xor U1801 (N_1801,N_1182,N_297);
or U1802 (N_1802,N_344,N_564);
or U1803 (N_1803,In_1729,In_2034);
or U1804 (N_1804,In_1347,In_2133);
and U1805 (N_1805,N_131,In_1);
and U1806 (N_1806,N_328,N_482);
nor U1807 (N_1807,In_1645,N_875);
xor U1808 (N_1808,N_155,N_1123);
nor U1809 (N_1809,In_1609,N_343);
nand U1810 (N_1810,In_241,N_60);
xnor U1811 (N_1811,N_1073,N_205);
nand U1812 (N_1812,In_583,N_433);
or U1813 (N_1813,N_335,In_1454);
xor U1814 (N_1814,In_2011,In_250);
nor U1815 (N_1815,In_5,N_391);
xor U1816 (N_1816,In_2230,In_402);
nand U1817 (N_1817,N_1045,N_927);
or U1818 (N_1818,In_42,In_2635);
nor U1819 (N_1819,N_345,N_799);
or U1820 (N_1820,N_183,In_883);
xnor U1821 (N_1821,In_2929,In_2339);
and U1822 (N_1822,In_1931,N_411);
nor U1823 (N_1823,N_52,N_473);
xor U1824 (N_1824,N_222,N_192);
and U1825 (N_1825,N_437,In_294);
and U1826 (N_1826,In_2560,In_1719);
and U1827 (N_1827,In_700,N_809);
nand U1828 (N_1828,N_1058,In_467);
or U1829 (N_1829,N_1028,In_55);
nand U1830 (N_1830,N_55,N_844);
xnor U1831 (N_1831,N_295,N_174);
or U1832 (N_1832,In_1535,N_1139);
or U1833 (N_1833,N_831,N_128);
or U1834 (N_1834,In_2716,N_253);
xor U1835 (N_1835,In_2291,N_334);
xnor U1836 (N_1836,N_1010,In_1946);
nor U1837 (N_1837,N_325,N_1158);
and U1838 (N_1838,N_868,N_48);
xnor U1839 (N_1839,In_2438,N_1100);
nor U1840 (N_1840,In_781,N_163);
nor U1841 (N_1841,N_507,In_2820);
nand U1842 (N_1842,N_585,N_898);
xor U1843 (N_1843,N_572,N_417);
xor U1844 (N_1844,N_792,N_1130);
or U1845 (N_1845,N_619,N_1067);
nand U1846 (N_1846,N_378,In_1507);
or U1847 (N_1847,N_53,In_2659);
xnor U1848 (N_1848,N_1027,N_697);
or U1849 (N_1849,N_1043,N_102);
xor U1850 (N_1850,In_2488,N_887);
and U1851 (N_1851,N_565,N_312);
xnor U1852 (N_1852,N_725,In_1797);
and U1853 (N_1853,In_2132,N_561);
nor U1854 (N_1854,N_1036,N_34);
nand U1855 (N_1855,In_2690,N_870);
or U1856 (N_1856,N_917,N_426);
and U1857 (N_1857,N_982,N_240);
nor U1858 (N_1858,N_550,In_815);
nor U1859 (N_1859,N_352,In_1092);
nand U1860 (N_1860,N_74,In_406);
and U1861 (N_1861,In_2958,N_817);
or U1862 (N_1862,N_476,In_646);
nand U1863 (N_1863,N_827,In_843);
nor U1864 (N_1864,N_400,In_2012);
nand U1865 (N_1865,N_967,N_1180);
xnor U1866 (N_1866,N_265,N_900);
xnor U1867 (N_1867,In_283,N_230);
and U1868 (N_1868,N_903,N_402);
nand U1869 (N_1869,N_939,N_85);
and U1870 (N_1870,N_1149,N_338);
nand U1871 (N_1871,In_1325,N_895);
xor U1872 (N_1872,N_376,N_999);
and U1873 (N_1873,N_910,N_955);
or U1874 (N_1874,In_376,In_128);
or U1875 (N_1875,N_660,N_581);
and U1876 (N_1876,N_381,N_867);
and U1877 (N_1877,N_495,N_11);
xnor U1878 (N_1878,In_1292,In_415);
nor U1879 (N_1879,In_947,N_1168);
or U1880 (N_1880,N_945,N_149);
xnor U1881 (N_1881,N_525,N_95);
or U1882 (N_1882,N_120,N_1105);
and U1883 (N_1883,N_692,In_436);
xnor U1884 (N_1884,N_1121,N_62);
nor U1885 (N_1885,N_744,N_778);
and U1886 (N_1886,N_147,N_327);
or U1887 (N_1887,N_803,In_824);
nand U1888 (N_1888,N_1097,N_997);
nand U1889 (N_1889,N_1133,N_478);
xor U1890 (N_1890,N_246,In_1714);
xnor U1891 (N_1891,N_304,In_673);
and U1892 (N_1892,In_2422,N_794);
xnor U1893 (N_1893,In_2389,In_1220);
and U1894 (N_1894,N_1108,In_2531);
and U1895 (N_1895,N_104,In_944);
or U1896 (N_1896,In_885,N_772);
nor U1897 (N_1897,N_361,In_2573);
xnor U1898 (N_1898,N_1143,N_480);
and U1899 (N_1899,N_127,In_2338);
or U1900 (N_1900,N_293,N_1138);
nand U1901 (N_1901,N_545,In_1872);
xor U1902 (N_1902,In_800,In_945);
xnor U1903 (N_1903,In_2779,N_998);
or U1904 (N_1904,N_928,N_922);
nor U1905 (N_1905,N_68,N_492);
nand U1906 (N_1906,N_94,N_1099);
or U1907 (N_1907,N_390,N_644);
xor U1908 (N_1908,N_1065,N_321);
or U1909 (N_1909,N_656,In_1843);
nor U1910 (N_1910,In_1080,In_72);
or U1911 (N_1911,N_92,N_444);
or U1912 (N_1912,N_716,In_1451);
xor U1913 (N_1913,N_151,N_924);
nor U1914 (N_1914,In_202,In_332);
xnor U1915 (N_1915,In_2853,N_617);
and U1916 (N_1916,In_759,N_1055);
nor U1917 (N_1917,N_369,N_832);
nand U1918 (N_1918,In_2526,N_693);
nand U1919 (N_1919,N_221,N_294);
xnor U1920 (N_1920,N_410,N_698);
and U1921 (N_1921,N_290,N_1120);
nor U1922 (N_1922,N_276,N_1113);
and U1923 (N_1923,N_516,N_15);
and U1924 (N_1924,In_1057,N_1079);
nand U1925 (N_1925,N_902,In_2380);
xor U1926 (N_1926,N_493,N_954);
nor U1927 (N_1927,N_983,In_1732);
xor U1928 (N_1928,In_2875,N_548);
nand U1929 (N_1929,N_914,N_719);
xor U1930 (N_1930,N_522,In_2672);
or U1931 (N_1931,N_569,In_1554);
xnor U1932 (N_1932,N_340,N_217);
nor U1933 (N_1933,In_1925,N_675);
nand U1934 (N_1934,In_559,N_1167);
or U1935 (N_1935,N_109,In_1346);
and U1936 (N_1936,N_438,N_598);
nand U1937 (N_1937,N_1181,In_1117);
xnor U1938 (N_1938,N_279,N_614);
and U1939 (N_1939,N_1031,N_58);
and U1940 (N_1940,In_902,N_663);
nand U1941 (N_1941,N_150,N_1132);
and U1942 (N_1942,N_1165,N_389);
or U1943 (N_1943,In_1030,N_248);
nand U1944 (N_1944,N_542,N_795);
nor U1945 (N_1945,N_636,In_980);
nor U1946 (N_1946,In_1633,N_125);
xor U1947 (N_1947,In_733,In_2332);
or U1948 (N_1948,In_2236,N_1006);
or U1949 (N_1949,In_2381,N_42);
xnor U1950 (N_1950,N_366,N_668);
nor U1951 (N_1951,In_1966,N_783);
xor U1952 (N_1952,N_813,N_201);
nor U1953 (N_1953,In_2814,N_267);
xnor U1954 (N_1954,In_805,N_269);
xnor U1955 (N_1955,N_443,N_536);
nor U1956 (N_1956,N_499,N_360);
nand U1957 (N_1957,N_388,N_142);
nand U1958 (N_1958,N_1196,N_384);
xor U1959 (N_1959,N_1048,N_650);
nand U1960 (N_1960,N_441,In_2646);
or U1961 (N_1961,N_918,N_785);
nand U1962 (N_1962,N_728,N_1081);
or U1963 (N_1963,N_807,N_907);
nand U1964 (N_1964,N_842,N_281);
and U1965 (N_1965,N_469,N_1032);
nor U1966 (N_1966,In_2981,In_297);
xor U1967 (N_1967,N_385,N_195);
or U1968 (N_1968,In_1860,N_430);
nor U1969 (N_1969,N_960,In_352);
xnor U1970 (N_1970,N_359,In_1705);
or U1971 (N_1971,In_1706,N_1177);
xnor U1972 (N_1972,N_757,In_1888);
xor U1973 (N_1973,N_919,N_341);
nor U1974 (N_1974,In_1078,N_54);
and U1975 (N_1975,N_610,N_368);
nor U1976 (N_1976,In_1413,In_1103);
xnor U1977 (N_1977,In_83,N_665);
or U1978 (N_1978,N_1150,N_673);
xnor U1979 (N_1979,In_1250,In_326);
nand U1980 (N_1980,N_460,N_71);
and U1981 (N_1981,N_7,In_1084);
or U1982 (N_1982,N_383,N_78);
xor U1983 (N_1983,N_1038,N_539);
nor U1984 (N_1984,N_743,N_1026);
nand U1985 (N_1985,In_1571,In_2028);
or U1986 (N_1986,In_2333,N_138);
and U1987 (N_1987,N_206,N_475);
or U1988 (N_1988,N_582,In_737);
and U1989 (N_1989,N_773,In_2330);
nor U1990 (N_1990,N_449,N_446);
nor U1991 (N_1991,In_2249,N_1012);
or U1992 (N_1992,N_198,N_551);
or U1993 (N_1993,In_2495,N_382);
xor U1994 (N_1994,N_197,In_2268);
nand U1995 (N_1995,N_299,N_215);
and U1996 (N_1996,In_90,In_2263);
and U1997 (N_1997,N_186,In_1897);
and U1998 (N_1998,N_203,N_737);
xor U1999 (N_1999,N_394,In_1775);
xnor U2000 (N_2000,In_917,In_1249);
nand U2001 (N_2001,N_822,In_224);
xnor U2002 (N_2002,N_583,N_1186);
xor U2003 (N_2003,N_244,N_422);
nor U2004 (N_2004,N_3,N_756);
nor U2005 (N_2005,In_229,N_447);
or U2006 (N_2006,In_1758,N_655);
nor U2007 (N_2007,N_1041,N_869);
xor U2008 (N_2008,N_1198,N_995);
xor U2009 (N_2009,N_587,N_578);
nor U2010 (N_2010,N_145,N_401);
or U2011 (N_2011,N_309,N_1173);
nor U2012 (N_2012,N_298,In_303);
nor U2013 (N_2013,N_266,In_594);
or U2014 (N_2014,N_13,N_489);
nand U2015 (N_2015,In_1186,N_947);
nor U2016 (N_2016,N_929,N_228);
or U2017 (N_2017,N_1016,In_873);
nand U2018 (N_2018,N_701,N_1131);
and U2019 (N_2019,N_1057,N_362);
xor U2020 (N_2020,N_1035,N_1192);
nand U2021 (N_2021,N_317,N_164);
and U2022 (N_2022,N_1094,N_219);
nor U2023 (N_2023,In_2070,N_4);
xor U2024 (N_2024,In_1463,In_549);
and U2025 (N_2025,N_117,N_41);
and U2026 (N_2026,In_553,N_532);
nor U2027 (N_2027,In_220,In_122);
or U2028 (N_2028,N_122,N_712);
and U2029 (N_2029,In_454,In_2061);
and U2030 (N_2030,N_451,In_170);
or U2031 (N_2031,N_838,N_303);
and U2032 (N_2032,N_791,In_2951);
nand U2033 (N_2033,In_1610,N_691);
nand U2034 (N_2034,N_577,N_1059);
xnor U2035 (N_2035,N_877,N_643);
or U2036 (N_2036,N_339,N_501);
nor U2037 (N_2037,N_1101,In_2457);
or U2038 (N_2038,N_123,N_505);
or U2039 (N_2039,N_750,N_951);
xnor U2040 (N_2040,N_863,N_0);
and U2041 (N_2041,In_2234,N_775);
xor U2042 (N_2042,N_193,N_1056);
or U2043 (N_2043,In_47,N_871);
nor U2044 (N_2044,N_89,N_1011);
nor U2045 (N_2045,N_1077,N_420);
and U2046 (N_2046,N_726,N_65);
xor U2047 (N_2047,In_2378,N_925);
or U2048 (N_2048,In_1849,N_264);
and U2049 (N_2049,N_387,N_622);
and U2050 (N_2050,N_184,In_2341);
nand U2051 (N_2051,N_638,N_124);
xor U2052 (N_2052,N_111,N_88);
or U2053 (N_2053,In_2043,In_2714);
nand U2054 (N_2054,N_448,In_2308);
and U2055 (N_2055,N_689,In_1054);
xor U2056 (N_2056,N_412,In_1409);
xor U2057 (N_2057,In_1717,In_1200);
nor U2058 (N_2058,N_957,In_2188);
nor U2059 (N_2059,N_976,N_770);
and U2060 (N_2060,In_2254,N_393);
nand U2061 (N_2061,In_1628,In_1642);
xnor U2062 (N_2062,In_1901,N_1119);
nand U2063 (N_2063,In_1760,In_1131);
nand U2064 (N_2064,In_1368,N_678);
and U2065 (N_2065,N_1021,N_758);
nor U2066 (N_2066,N_989,N_166);
nor U2067 (N_2067,In_2013,In_2213);
xor U2068 (N_2068,N_318,N_690);
nor U2069 (N_2069,In_787,N_886);
xor U2070 (N_2070,In_677,N_1179);
nand U2071 (N_2071,In_462,In_648);
xnor U2072 (N_2072,In_421,N_686);
nor U2073 (N_2073,N_162,N_790);
and U2074 (N_2074,N_1122,N_608);
and U2075 (N_2075,In_1828,In_2058);
xor U2076 (N_2076,N_380,In_1841);
or U2077 (N_2077,N_971,N_749);
or U2078 (N_2078,N_1154,In_701);
or U2079 (N_2079,In_330,N_613);
nand U2080 (N_2080,N_641,In_1561);
and U2081 (N_2081,N_178,In_2966);
nand U2082 (N_2082,N_713,In_649);
and U2083 (N_2083,In_1023,N_948);
nor U2084 (N_2084,N_805,N_208);
and U2085 (N_2085,N_621,N_738);
nand U2086 (N_2086,N_1095,N_1153);
nor U2087 (N_2087,N_977,In_625);
or U2088 (N_2088,N_1078,N_788);
and U2089 (N_2089,N_912,N_194);
nor U2090 (N_2090,N_337,N_275);
and U2091 (N_2091,N_333,N_22);
nor U2092 (N_2092,In_1911,N_46);
nand U2093 (N_2093,N_861,N_740);
and U2094 (N_2094,N_1157,In_336);
xnor U2095 (N_2095,In_1419,N_419);
and U2096 (N_2096,In_450,N_742);
xor U2097 (N_2097,N_915,In_366);
and U2098 (N_2098,N_706,In_1270);
nand U2099 (N_2099,N_399,N_254);
and U2100 (N_2100,N_25,N_318);
nor U2101 (N_2101,In_800,N_1190);
nand U2102 (N_2102,N_370,In_2509);
or U2103 (N_2103,In_787,In_514);
or U2104 (N_2104,N_834,In_246);
or U2105 (N_2105,N_1087,N_1047);
nor U2106 (N_2106,In_2256,In_1703);
or U2107 (N_2107,N_1000,In_2005);
and U2108 (N_2108,N_1034,N_71);
xnor U2109 (N_2109,N_842,N_775);
xor U2110 (N_2110,N_751,N_757);
or U2111 (N_2111,N_1010,N_547);
and U2112 (N_2112,In_2043,N_164);
nand U2113 (N_2113,N_239,In_204);
nand U2114 (N_2114,In_1518,N_588);
nand U2115 (N_2115,In_352,In_2848);
nand U2116 (N_2116,N_683,N_294);
and U2117 (N_2117,In_336,In_1714);
nor U2118 (N_2118,N_160,N_705);
and U2119 (N_2119,N_746,N_696);
or U2120 (N_2120,N_953,In_2707);
nor U2121 (N_2121,N_806,In_2387);
and U2122 (N_2122,N_456,N_617);
or U2123 (N_2123,N_1014,N_141);
nor U2124 (N_2124,N_104,N_371);
nand U2125 (N_2125,In_883,In_1328);
and U2126 (N_2126,In_1421,In_1925);
nand U2127 (N_2127,N_137,In_1456);
nor U2128 (N_2128,In_1870,N_131);
xor U2129 (N_2129,N_231,In_844);
and U2130 (N_2130,In_2378,In_336);
xor U2131 (N_2131,N_30,N_567);
nor U2132 (N_2132,N_1105,N_448);
or U2133 (N_2133,In_42,N_591);
xor U2134 (N_2134,N_938,N_787);
and U2135 (N_2135,N_1074,N_16);
nor U2136 (N_2136,N_119,N_1172);
or U2137 (N_2137,N_1136,In_2055);
nand U2138 (N_2138,In_680,In_352);
nor U2139 (N_2139,N_1008,N_1014);
or U2140 (N_2140,N_246,N_142);
and U2141 (N_2141,N_45,In_2054);
xor U2142 (N_2142,N_433,N_631);
and U2143 (N_2143,In_2213,N_985);
xnor U2144 (N_2144,N_666,N_165);
nor U2145 (N_2145,N_324,In_2707);
or U2146 (N_2146,In_1240,In_450);
nand U2147 (N_2147,N_923,N_80);
nand U2148 (N_2148,N_667,N_761);
and U2149 (N_2149,N_471,N_908);
and U2150 (N_2150,N_946,In_442);
xnor U2151 (N_2151,N_1096,N_966);
nor U2152 (N_2152,N_1030,In_689);
nand U2153 (N_2153,N_140,In_442);
or U2154 (N_2154,N_117,N_482);
nand U2155 (N_2155,N_171,N_376);
nand U2156 (N_2156,In_1419,N_805);
nor U2157 (N_2157,In_2365,N_969);
nand U2158 (N_2158,N_360,N_920);
and U2159 (N_2159,In_2767,N_230);
and U2160 (N_2160,N_806,N_1156);
xnor U2161 (N_2161,N_507,N_191);
xor U2162 (N_2162,N_1187,In_72);
and U2163 (N_2163,In_349,N_103);
xnor U2164 (N_2164,N_625,In_2603);
nor U2165 (N_2165,N_946,In_1619);
and U2166 (N_2166,N_393,In_2463);
xor U2167 (N_2167,N_751,In_311);
and U2168 (N_2168,N_1161,In_297);
or U2169 (N_2169,N_1150,In_1560);
nor U2170 (N_2170,N_529,N_442);
xor U2171 (N_2171,N_595,In_2659);
nand U2172 (N_2172,N_954,N_424);
xor U2173 (N_2173,N_842,N_1094);
or U2174 (N_2174,In_2474,N_818);
nand U2175 (N_2175,In_2580,N_484);
and U2176 (N_2176,N_950,N_656);
and U2177 (N_2177,N_612,In_2875);
xnor U2178 (N_2178,N_152,In_936);
xnor U2179 (N_2179,N_801,N_45);
nand U2180 (N_2180,N_155,N_598);
xor U2181 (N_2181,In_378,N_170);
xnor U2182 (N_2182,N_938,N_1071);
or U2183 (N_2183,N_1026,In_1893);
xnor U2184 (N_2184,N_1095,N_453);
and U2185 (N_2185,N_492,In_2526);
nor U2186 (N_2186,N_580,In_467);
nand U2187 (N_2187,N_800,In_2289);
or U2188 (N_2188,N_789,N_83);
or U2189 (N_2189,N_289,N_229);
or U2190 (N_2190,In_781,N_900);
or U2191 (N_2191,N_240,N_11);
nor U2192 (N_2192,N_221,In_397);
xor U2193 (N_2193,N_528,N_937);
nor U2194 (N_2194,N_191,In_907);
or U2195 (N_2195,In_895,In_1313);
nor U2196 (N_2196,N_356,N_329);
nor U2197 (N_2197,In_90,N_588);
xor U2198 (N_2198,N_101,N_400);
or U2199 (N_2199,In_756,N_15);
nor U2200 (N_2200,In_293,N_982);
nor U2201 (N_2201,N_435,N_700);
nand U2202 (N_2202,N_517,In_1074);
xor U2203 (N_2203,N_143,In_152);
nor U2204 (N_2204,N_882,N_56);
xnor U2205 (N_2205,In_2323,N_1087);
or U2206 (N_2206,In_377,N_798);
xnor U2207 (N_2207,In_1347,N_513);
nor U2208 (N_2208,In_1074,In_895);
nand U2209 (N_2209,N_144,N_1184);
nor U2210 (N_2210,In_1403,In_648);
or U2211 (N_2211,N_407,In_475);
nor U2212 (N_2212,N_70,N_954);
nor U2213 (N_2213,N_284,N_645);
and U2214 (N_2214,N_619,In_907);
nand U2215 (N_2215,N_638,N_349);
nor U2216 (N_2216,N_106,N_156);
xnor U2217 (N_2217,N_202,In_2848);
nor U2218 (N_2218,In_2132,N_319);
or U2219 (N_2219,N_316,N_1074);
nor U2220 (N_2220,N_398,In_367);
nand U2221 (N_2221,In_1465,N_319);
nor U2222 (N_2222,In_2195,In_2226);
or U2223 (N_2223,N_1129,N_247);
or U2224 (N_2224,In_2014,In_851);
nand U2225 (N_2225,In_224,N_373);
nand U2226 (N_2226,N_316,N_419);
nor U2227 (N_2227,N_223,N_1011);
nor U2228 (N_2228,In_2814,N_51);
and U2229 (N_2229,In_2450,N_278);
or U2230 (N_2230,N_1015,N_983);
or U2231 (N_2231,N_3,N_417);
xnor U2232 (N_2232,N_445,N_1064);
xnor U2233 (N_2233,In_98,N_117);
and U2234 (N_2234,N_346,N_506);
and U2235 (N_2235,N_70,In_2389);
xnor U2236 (N_2236,In_2714,In_1726);
xnor U2237 (N_2237,In_2724,N_258);
nand U2238 (N_2238,N_699,In_2693);
and U2239 (N_2239,N_575,N_724);
nor U2240 (N_2240,N_309,N_347);
and U2241 (N_2241,In_646,In_973);
and U2242 (N_2242,N_592,N_140);
nor U2243 (N_2243,In_390,In_1917);
and U2244 (N_2244,N_1129,N_1009);
nand U2245 (N_2245,N_1167,In_2767);
nand U2246 (N_2246,N_898,N_821);
nand U2247 (N_2247,N_934,N_260);
nor U2248 (N_2248,In_265,N_1016);
nor U2249 (N_2249,N_481,N_31);
xor U2250 (N_2250,N_438,N_320);
nand U2251 (N_2251,In_164,N_353);
and U2252 (N_2252,In_1610,N_1189);
or U2253 (N_2253,In_2488,In_2697);
and U2254 (N_2254,N_702,N_795);
nor U2255 (N_2255,In_1509,N_297);
and U2256 (N_2256,N_916,N_309);
nor U2257 (N_2257,N_594,N_819);
nand U2258 (N_2258,N_235,In_2067);
nand U2259 (N_2259,N_297,In_13);
nor U2260 (N_2260,N_82,N_95);
or U2261 (N_2261,N_366,N_69);
xnor U2262 (N_2262,N_830,In_1177);
and U2263 (N_2263,In_1733,N_324);
and U2264 (N_2264,N_520,N_919);
xor U2265 (N_2265,N_872,N_1054);
nand U2266 (N_2266,N_762,In_349);
nand U2267 (N_2267,In_947,N_1036);
xor U2268 (N_2268,N_404,N_63);
nand U2269 (N_2269,In_128,N_639);
xnor U2270 (N_2270,N_294,N_1008);
or U2271 (N_2271,N_675,In_2154);
xor U2272 (N_2272,N_226,N_886);
nand U2273 (N_2273,N_178,N_145);
nand U2274 (N_2274,N_904,In_659);
and U2275 (N_2275,N_1,N_624);
nor U2276 (N_2276,N_647,N_1004);
or U2277 (N_2277,N_361,N_1024);
xnor U2278 (N_2278,N_518,In_2820);
xor U2279 (N_2279,In_2226,N_662);
or U2280 (N_2280,N_751,In_1553);
nand U2281 (N_2281,N_539,In_2981);
xnor U2282 (N_2282,N_1114,In_266);
nor U2283 (N_2283,N_50,In_2890);
or U2284 (N_2284,N_982,In_300);
xor U2285 (N_2285,N_235,N_848);
nand U2286 (N_2286,In_800,N_43);
nor U2287 (N_2287,N_975,In_2697);
xnor U2288 (N_2288,N_636,N_1061);
nor U2289 (N_2289,N_144,N_952);
or U2290 (N_2290,N_1067,In_2373);
nand U2291 (N_2291,N_450,In_2630);
or U2292 (N_2292,N_975,N_825);
nor U2293 (N_2293,N_935,In_2263);
nor U2294 (N_2294,In_2310,N_955);
or U2295 (N_2295,N_763,N_154);
and U2296 (N_2296,N_886,N_546);
or U2297 (N_2297,N_626,N_126);
nand U2298 (N_2298,N_1070,In_2268);
nand U2299 (N_2299,N_849,N_756);
xor U2300 (N_2300,In_442,N_778);
and U2301 (N_2301,N_488,N_6);
and U2302 (N_2302,N_566,N_809);
and U2303 (N_2303,N_74,N_741);
or U2304 (N_2304,In_2890,N_25);
or U2305 (N_2305,N_991,N_1028);
xnor U2306 (N_2306,In_737,In_2380);
nor U2307 (N_2307,In_2635,N_45);
xnor U2308 (N_2308,N_932,N_842);
and U2309 (N_2309,N_978,N_702);
nand U2310 (N_2310,N_933,N_45);
nand U2311 (N_2311,N_180,In_1413);
or U2312 (N_2312,N_412,N_401);
and U2313 (N_2313,N_413,N_712);
xor U2314 (N_2314,N_1085,In_2131);
or U2315 (N_2315,N_394,N_175);
xnor U2316 (N_2316,In_1186,N_1113);
nor U2317 (N_2317,N_1103,N_244);
nand U2318 (N_2318,In_907,In_1221);
xor U2319 (N_2319,N_1091,N_278);
nor U2320 (N_2320,N_987,N_628);
xor U2321 (N_2321,In_57,N_536);
nor U2322 (N_2322,N_1006,In_2037);
nor U2323 (N_2323,In_805,N_1074);
and U2324 (N_2324,In_659,N_348);
and U2325 (N_2325,N_929,N_738);
or U2326 (N_2326,N_1011,N_337);
nor U2327 (N_2327,In_1465,N_896);
and U2328 (N_2328,N_914,N_1181);
nand U2329 (N_2329,N_584,In_1096);
nand U2330 (N_2330,N_688,N_139);
or U2331 (N_2331,N_1127,N_11);
and U2332 (N_2332,In_1154,N_157);
nand U2333 (N_2333,In_406,N_898);
nand U2334 (N_2334,N_931,N_31);
or U2335 (N_2335,In_700,N_431);
nor U2336 (N_2336,N_293,N_262);
or U2337 (N_2337,N_452,In_2046);
nor U2338 (N_2338,N_827,N_669);
nor U2339 (N_2339,N_843,In_2275);
xnor U2340 (N_2340,In_2234,N_991);
or U2341 (N_2341,N_1059,N_545);
or U2342 (N_2342,N_738,N_810);
nor U2343 (N_2343,N_499,N_444);
xnor U2344 (N_2344,N_567,In_2304);
and U2345 (N_2345,In_379,N_1103);
nor U2346 (N_2346,N_192,N_78);
or U2347 (N_2347,N_883,In_2387);
nand U2348 (N_2348,N_580,N_969);
nand U2349 (N_2349,In_1753,N_95);
nor U2350 (N_2350,In_1006,N_71);
nor U2351 (N_2351,N_314,N_468);
xnor U2352 (N_2352,N_795,N_907);
xnor U2353 (N_2353,In_1546,In_220);
nand U2354 (N_2354,N_775,In_851);
or U2355 (N_2355,In_2761,N_741);
nand U2356 (N_2356,In_2304,N_158);
nor U2357 (N_2357,N_199,In_2526);
nand U2358 (N_2358,N_584,N_342);
and U2359 (N_2359,In_376,N_764);
xor U2360 (N_2360,N_472,N_792);
and U2361 (N_2361,N_682,N_981);
nand U2362 (N_2362,N_886,In_2951);
and U2363 (N_2363,N_25,In_733);
nand U2364 (N_2364,In_1235,N_841);
and U2365 (N_2365,In_1074,N_1151);
or U2366 (N_2366,N_653,N_140);
or U2367 (N_2367,N_265,N_845);
and U2368 (N_2368,In_2458,N_582);
xnor U2369 (N_2369,N_117,In_2119);
nand U2370 (N_2370,In_1499,N_985);
xnor U2371 (N_2371,In_2848,N_477);
nand U2372 (N_2372,N_300,N_15);
or U2373 (N_2373,N_317,In_205);
xor U2374 (N_2374,N_306,In_648);
or U2375 (N_2375,In_2058,N_753);
nand U2376 (N_2376,N_465,N_972);
xnor U2377 (N_2377,In_202,N_1022);
and U2378 (N_2378,In_346,In_939);
nor U2379 (N_2379,N_1023,N_964);
nand U2380 (N_2380,N_633,N_567);
or U2381 (N_2381,N_742,N_306);
xor U2382 (N_2382,N_348,N_920);
xor U2383 (N_2383,N_88,In_1519);
nor U2384 (N_2384,N_300,N_1199);
and U2385 (N_2385,In_677,N_149);
xor U2386 (N_2386,N_301,N_309);
xnor U2387 (N_2387,N_1077,In_1023);
and U2388 (N_2388,N_396,N_392);
nor U2389 (N_2389,In_1398,N_563);
nand U2390 (N_2390,In_170,N_541);
nand U2391 (N_2391,N_627,In_2911);
xnor U2392 (N_2392,In_229,In_321);
xnor U2393 (N_2393,N_630,N_639);
nand U2394 (N_2394,In_487,N_148);
xnor U2395 (N_2395,N_489,N_735);
and U2396 (N_2396,N_1090,N_649);
nand U2397 (N_2397,N_1176,In_1235);
xnor U2398 (N_2398,In_1643,In_462);
and U2399 (N_2399,N_288,In_2450);
nand U2400 (N_2400,N_1838,N_1416);
or U2401 (N_2401,N_1433,N_2290);
xnor U2402 (N_2402,N_1605,N_1528);
nand U2403 (N_2403,N_2149,N_2366);
xor U2404 (N_2404,N_1606,N_1890);
xnor U2405 (N_2405,N_1389,N_1777);
and U2406 (N_2406,N_2129,N_1685);
nand U2407 (N_2407,N_2318,N_2273);
or U2408 (N_2408,N_1790,N_2211);
nand U2409 (N_2409,N_1537,N_2288);
and U2410 (N_2410,N_2259,N_1627);
and U2411 (N_2411,N_1492,N_2134);
xnor U2412 (N_2412,N_2367,N_1442);
nand U2413 (N_2413,N_2344,N_1424);
nor U2414 (N_2414,N_2039,N_2387);
nand U2415 (N_2415,N_2040,N_2301);
nor U2416 (N_2416,N_2221,N_2314);
xor U2417 (N_2417,N_2078,N_1895);
and U2418 (N_2418,N_1620,N_2092);
and U2419 (N_2419,N_2014,N_1445);
or U2420 (N_2420,N_1354,N_1650);
and U2421 (N_2421,N_1529,N_1574);
xnor U2422 (N_2422,N_1710,N_1258);
or U2423 (N_2423,N_2208,N_2369);
xnor U2424 (N_2424,N_2361,N_1806);
nor U2425 (N_2425,N_1321,N_2026);
nand U2426 (N_2426,N_1207,N_1860);
nand U2427 (N_2427,N_1305,N_1874);
nand U2428 (N_2428,N_1520,N_2325);
nand U2429 (N_2429,N_1669,N_1300);
nor U2430 (N_2430,N_1229,N_1997);
and U2431 (N_2431,N_1314,N_1603);
and U2432 (N_2432,N_2130,N_2010);
nand U2433 (N_2433,N_2021,N_1476);
xnor U2434 (N_2434,N_2048,N_2319);
xnor U2435 (N_2435,N_2277,N_1535);
xor U2436 (N_2436,N_1271,N_1651);
nand U2437 (N_2437,N_1960,N_1660);
or U2438 (N_2438,N_1902,N_2062);
nor U2439 (N_2439,N_1379,N_1430);
and U2440 (N_2440,N_2239,N_2128);
nand U2441 (N_2441,N_2008,N_1940);
nand U2442 (N_2442,N_1532,N_1285);
or U2443 (N_2443,N_1501,N_1594);
nor U2444 (N_2444,N_2107,N_2151);
nand U2445 (N_2445,N_1864,N_1901);
xor U2446 (N_2446,N_1761,N_1545);
nor U2447 (N_2447,N_2087,N_1434);
xor U2448 (N_2448,N_1543,N_2020);
nand U2449 (N_2449,N_1593,N_2046);
nor U2450 (N_2450,N_2090,N_1302);
and U2451 (N_2451,N_2044,N_1971);
and U2452 (N_2452,N_1724,N_1222);
xnor U2453 (N_2453,N_1220,N_2145);
and U2454 (N_2454,N_1201,N_2296);
or U2455 (N_2455,N_2338,N_2225);
nor U2456 (N_2456,N_1250,N_1371);
nand U2457 (N_2457,N_1735,N_1468);
nor U2458 (N_2458,N_1696,N_1580);
nand U2459 (N_2459,N_1984,N_1395);
and U2460 (N_2460,N_1360,N_1571);
or U2461 (N_2461,N_1736,N_1474);
or U2462 (N_2462,N_2279,N_1616);
nand U2463 (N_2463,N_2306,N_1567);
nand U2464 (N_2464,N_2009,N_2043);
nand U2465 (N_2465,N_1401,N_1270);
and U2466 (N_2466,N_1425,N_1772);
nand U2467 (N_2467,N_2059,N_1980);
and U2468 (N_2468,N_1392,N_1586);
nand U2469 (N_2469,N_2381,N_2118);
or U2470 (N_2470,N_1265,N_1942);
nor U2471 (N_2471,N_1269,N_1609);
and U2472 (N_2472,N_2113,N_1415);
and U2473 (N_2473,N_2158,N_1578);
nor U2474 (N_2474,N_2348,N_2322);
or U2475 (N_2475,N_2155,N_1823);
and U2476 (N_2476,N_2389,N_1706);
or U2477 (N_2477,N_2250,N_2198);
nor U2478 (N_2478,N_2212,N_2170);
nand U2479 (N_2479,N_1982,N_1249);
xor U2480 (N_2480,N_2312,N_1503);
or U2481 (N_2481,N_1703,N_2311);
nor U2482 (N_2482,N_1938,N_2127);
nand U2483 (N_2483,N_1753,N_1534);
nand U2484 (N_2484,N_1979,N_1654);
xor U2485 (N_2485,N_1376,N_1555);
xor U2486 (N_2486,N_2206,N_1511);
or U2487 (N_2487,N_2380,N_1732);
or U2488 (N_2488,N_1811,N_2252);
or U2489 (N_2489,N_2308,N_1552);
and U2490 (N_2490,N_1289,N_2139);
or U2491 (N_2491,N_2205,N_1959);
xnor U2492 (N_2492,N_1839,N_1983);
or U2493 (N_2493,N_2335,N_1463);
nand U2494 (N_2494,N_1410,N_1251);
nand U2495 (N_2495,N_2007,N_1284);
xnor U2496 (N_2496,N_1252,N_2375);
nand U2497 (N_2497,N_1438,N_1527);
or U2498 (N_2498,N_1812,N_1619);
xor U2499 (N_2499,N_2353,N_2185);
nor U2500 (N_2500,N_1497,N_2069);
xnor U2501 (N_2501,N_1968,N_2166);
xor U2502 (N_2502,N_1486,N_1862);
or U2503 (N_2503,N_1335,N_1840);
and U2504 (N_2504,N_1319,N_1701);
xnor U2505 (N_2505,N_1718,N_1502);
and U2506 (N_2506,N_2121,N_1469);
or U2507 (N_2507,N_2261,N_1450);
or U2508 (N_2508,N_2359,N_1992);
and U2509 (N_2509,N_2254,N_1693);
or U2510 (N_2510,N_1930,N_1952);
nor U2511 (N_2511,N_1280,N_1741);
xor U2512 (N_2512,N_1523,N_2000);
nand U2513 (N_2513,N_1715,N_1390);
or U2514 (N_2514,N_1244,N_1647);
xnor U2515 (N_2515,N_1372,N_2179);
and U2516 (N_2516,N_1668,N_1883);
nor U2517 (N_2517,N_1870,N_2327);
and U2518 (N_2518,N_1743,N_2349);
nand U2519 (N_2519,N_1924,N_2088);
nand U2520 (N_2520,N_1454,N_1639);
nor U2521 (N_2521,N_1880,N_1751);
or U2522 (N_2522,N_1596,N_1460);
and U2523 (N_2523,N_2214,N_1205);
xor U2524 (N_2524,N_2388,N_1598);
xnor U2525 (N_2525,N_1491,N_1636);
or U2526 (N_2526,N_1867,N_2240);
and U2527 (N_2527,N_2054,N_2159);
nor U2528 (N_2528,N_1807,N_2393);
nor U2529 (N_2529,N_2244,N_1595);
or U2530 (N_2530,N_1334,N_1226);
or U2531 (N_2531,N_1591,N_1509);
and U2532 (N_2532,N_1286,N_2124);
or U2533 (N_2533,N_1353,N_1411);
nor U2534 (N_2534,N_1481,N_1990);
or U2535 (N_2535,N_1394,N_2031);
and U2536 (N_2536,N_2120,N_1246);
xor U2537 (N_2537,N_2309,N_1564);
nor U2538 (N_2538,N_1333,N_1809);
nor U2539 (N_2539,N_1978,N_1854);
and U2540 (N_2540,N_1786,N_1311);
nand U2541 (N_2541,N_1209,N_2017);
and U2542 (N_2542,N_1458,N_1573);
nor U2543 (N_2543,N_1684,N_2077);
nand U2544 (N_2544,N_1602,N_2227);
xnor U2545 (N_2545,N_1652,N_2153);
or U2546 (N_2546,N_2362,N_1256);
nand U2547 (N_2547,N_2099,N_1836);
xor U2548 (N_2548,N_1771,N_2083);
and U2549 (N_2549,N_1780,N_2012);
and U2550 (N_2550,N_1932,N_2045);
nor U2551 (N_2551,N_1871,N_1640);
xor U2552 (N_2552,N_1435,N_2299);
xor U2553 (N_2553,N_1560,N_1259);
nand U2554 (N_2554,N_1533,N_1752);
and U2555 (N_2555,N_2247,N_2142);
xor U2556 (N_2556,N_1775,N_1349);
nand U2557 (N_2557,N_2224,N_1461);
nor U2558 (N_2558,N_1919,N_2372);
xor U2559 (N_2559,N_1202,N_1643);
xor U2560 (N_2560,N_1958,N_1566);
and U2561 (N_2561,N_2096,N_1290);
and U2562 (N_2562,N_1556,N_2167);
or U2563 (N_2563,N_2110,N_2226);
xor U2564 (N_2564,N_2177,N_1500);
and U2565 (N_2565,N_1623,N_1905);
nand U2566 (N_2566,N_2234,N_1318);
and U2567 (N_2567,N_2269,N_1536);
or U2568 (N_2568,N_2154,N_1891);
and U2569 (N_2569,N_2071,N_2233);
and U2570 (N_2570,N_2394,N_1981);
and U2571 (N_2571,N_1826,N_1346);
xnor U2572 (N_2572,N_1581,N_1393);
nand U2573 (N_2573,N_2194,N_1553);
nor U2574 (N_2574,N_1691,N_1236);
xnor U2575 (N_2575,N_2131,N_1549);
or U2576 (N_2576,N_1694,N_1307);
nor U2577 (N_2577,N_1877,N_1316);
and U2578 (N_2578,N_1234,N_1677);
and U2579 (N_2579,N_1784,N_1357);
nand U2580 (N_2580,N_2386,N_1204);
xnor U2581 (N_2581,N_2041,N_1766);
nor U2582 (N_2582,N_1426,N_2392);
and U2583 (N_2583,N_1294,N_1588);
nor U2584 (N_2584,N_1542,N_2085);
and U2585 (N_2585,N_2188,N_1383);
nor U2586 (N_2586,N_1748,N_1687);
nor U2587 (N_2587,N_2333,N_1985);
and U2588 (N_2588,N_1247,N_1713);
and U2589 (N_2589,N_2370,N_2169);
and U2590 (N_2590,N_1667,N_1377);
nand U2591 (N_2591,N_2326,N_1309);
nand U2592 (N_2592,N_1989,N_1245);
nand U2593 (N_2593,N_1731,N_1856);
xor U2594 (N_2594,N_2172,N_1587);
nand U2595 (N_2595,N_2200,N_1576);
xnor U2596 (N_2596,N_1911,N_1261);
or U2597 (N_2597,N_1929,N_1844);
nor U2598 (N_2598,N_2262,N_1853);
and U2599 (N_2599,N_2228,N_2248);
xnor U2600 (N_2600,N_1243,N_1712);
and U2601 (N_2601,N_1274,N_1879);
nand U2602 (N_2602,N_2263,N_2161);
xnor U2603 (N_2603,N_2382,N_1792);
xor U2604 (N_2604,N_1608,N_2339);
and U2605 (N_2605,N_1950,N_2006);
nand U2606 (N_2606,N_1613,N_2191);
and U2607 (N_2607,N_2034,N_1584);
nand U2608 (N_2608,N_2398,N_1373);
nand U2609 (N_2609,N_1459,N_1208);
nor U2610 (N_2610,N_2132,N_2286);
xnor U2611 (N_2611,N_1876,N_1355);
or U2612 (N_2612,N_2255,N_2005);
or U2613 (N_2613,N_1343,N_1657);
or U2614 (N_2614,N_1708,N_1746);
nand U2615 (N_2615,N_1789,N_1575);
nor U2616 (N_2616,N_1530,N_1918);
and U2617 (N_2617,N_1539,N_2303);
or U2618 (N_2618,N_1404,N_1402);
and U2619 (N_2619,N_2049,N_1212);
or U2620 (N_2620,N_2135,N_1881);
nand U2621 (N_2621,N_1628,N_1541);
nand U2622 (N_2622,N_1466,N_1945);
nand U2623 (N_2623,N_1849,N_1916);
nor U2624 (N_2624,N_1625,N_1683);
and U2625 (N_2625,N_2390,N_1794);
xnor U2626 (N_2626,N_1688,N_1827);
nand U2627 (N_2627,N_1730,N_1783);
xor U2628 (N_2628,N_1324,N_1240);
nand U2629 (N_2629,N_1820,N_1336);
and U2630 (N_2630,N_2196,N_1721);
xnor U2631 (N_2631,N_2025,N_2152);
xnor U2632 (N_2632,N_1728,N_1829);
nand U2633 (N_2633,N_1554,N_1590);
and U2634 (N_2634,N_1615,N_1843);
xnor U2635 (N_2635,N_1776,N_2193);
xor U2636 (N_2636,N_1779,N_1462);
xnor U2637 (N_2637,N_2297,N_1592);
and U2638 (N_2638,N_1695,N_2133);
or U2639 (N_2639,N_1634,N_1317);
nor U2640 (N_2640,N_1947,N_2001);
nor U2641 (N_2641,N_1296,N_2105);
or U2642 (N_2642,N_2385,N_1241);
nand U2643 (N_2643,N_2371,N_1493);
or U2644 (N_2644,N_1359,N_1863);
or U2645 (N_2645,N_1365,N_2203);
or U2646 (N_2646,N_1663,N_2190);
or U2647 (N_2647,N_1873,N_1381);
or U2648 (N_2648,N_2317,N_2073);
xnor U2649 (N_2649,N_1561,N_2241);
and U2650 (N_2650,N_1449,N_1488);
nor U2651 (N_2651,N_2374,N_1726);
and U2652 (N_2652,N_1943,N_1907);
or U2653 (N_2653,N_2345,N_1966);
nor U2654 (N_2654,N_2140,N_1690);
or U2655 (N_2655,N_1325,N_1483);
nor U2656 (N_2656,N_2180,N_1750);
or U2657 (N_2657,N_1572,N_2016);
or U2658 (N_2658,N_1577,N_1352);
or U2659 (N_2659,N_1885,N_2164);
xnor U2660 (N_2660,N_2383,N_1366);
xor U2661 (N_2661,N_2209,N_2053);
nand U2662 (N_2662,N_1631,N_2218);
nand U2663 (N_2663,N_2271,N_1646);
and U2664 (N_2664,N_2084,N_1914);
nand U2665 (N_2665,N_1418,N_1872);
and U2666 (N_2666,N_2013,N_1810);
xnor U2667 (N_2667,N_2011,N_1589);
or U2668 (N_2668,N_1364,N_1447);
or U2669 (N_2669,N_2242,N_2186);
and U2670 (N_2670,N_1341,N_1579);
or U2671 (N_2671,N_1740,N_1448);
nand U2672 (N_2672,N_1818,N_2137);
nand U2673 (N_2673,N_1725,N_2215);
nand U2674 (N_2674,N_1729,N_2282);
and U2675 (N_2675,N_2183,N_1283);
xnor U2676 (N_2676,N_2114,N_1799);
xor U2677 (N_2677,N_1275,N_1638);
xor U2678 (N_2678,N_1624,N_2397);
nor U2679 (N_2679,N_2298,N_2079);
or U2680 (N_2680,N_1975,N_1681);
and U2681 (N_2681,N_1697,N_2160);
nor U2682 (N_2682,N_1868,N_1407);
nand U2683 (N_2683,N_1676,N_1742);
nand U2684 (N_2684,N_2094,N_2201);
or U2685 (N_2685,N_1455,N_2258);
and U2686 (N_2686,N_1963,N_1951);
nand U2687 (N_2687,N_1717,N_2341);
or U2688 (N_2688,N_2111,N_1582);
or U2689 (N_2689,N_1745,N_1215);
or U2690 (N_2690,N_1451,N_1206);
xor U2691 (N_2691,N_2336,N_1817);
xor U2692 (N_2692,N_1898,N_1384);
or U2693 (N_2693,N_1999,N_1232);
nand U2694 (N_2694,N_2081,N_1852);
nor U2695 (N_2695,N_2310,N_1765);
or U2696 (N_2696,N_2057,N_1709);
and U2697 (N_2697,N_1887,N_1671);
nand U2698 (N_2698,N_2251,N_1977);
xnor U2699 (N_2699,N_2274,N_2032);
xnor U2700 (N_2700,N_1969,N_2384);
nand U2701 (N_2701,N_1266,N_1964);
nand U2702 (N_2702,N_1457,N_2220);
nand U2703 (N_2703,N_1396,N_1298);
nand U2704 (N_2704,N_2103,N_2080);
xnor U2705 (N_2705,N_2146,N_2123);
nor U2706 (N_2706,N_2267,N_2222);
nor U2707 (N_2707,N_1544,N_1405);
or U2708 (N_2708,N_1716,N_1931);
nor U2709 (N_2709,N_1928,N_2246);
nor U2710 (N_2710,N_1848,N_1387);
nand U2711 (N_2711,N_2323,N_1223);
and U2712 (N_2712,N_1484,N_1277);
xnor U2713 (N_2713,N_1475,N_2056);
and U2714 (N_2714,N_2334,N_2156);
and U2715 (N_2715,N_2238,N_1641);
nand U2716 (N_2716,N_1515,N_1937);
and U2717 (N_2717,N_2192,N_1540);
xor U2718 (N_2718,N_1224,N_1644);
and U2719 (N_2719,N_1795,N_1774);
and U2720 (N_2720,N_1399,N_1443);
and U2721 (N_2721,N_2148,N_1568);
nand U2722 (N_2722,N_2378,N_2015);
or U2723 (N_2723,N_1330,N_2294);
nor U2724 (N_2724,N_1427,N_1673);
or U2725 (N_2725,N_1378,N_2283);
nand U2726 (N_2726,N_2237,N_2376);
nand U2727 (N_2727,N_1478,N_2178);
xor U2728 (N_2728,N_2363,N_1941);
or U2729 (N_2729,N_2230,N_1632);
xor U2730 (N_2730,N_1299,N_1756);
nand U2731 (N_2731,N_1456,N_1257);
xnor U2732 (N_2732,N_1913,N_1920);
or U2733 (N_2733,N_1858,N_1446);
nor U2734 (N_2734,N_2281,N_2302);
nand U2735 (N_2735,N_1367,N_1973);
and U2736 (N_2736,N_1525,N_1522);
nand U2737 (N_2737,N_2061,N_1287);
nor U2738 (N_2738,N_1508,N_1328);
xnor U2739 (N_2739,N_1822,N_1961);
or U2740 (N_2740,N_1626,N_1944);
nor U2741 (N_2741,N_1380,N_1954);
nor U2742 (N_2742,N_1313,N_2285);
nand U2743 (N_2743,N_1218,N_1239);
or U2744 (N_2744,N_2189,N_1308);
xnor U2745 (N_2745,N_2207,N_2102);
and U2746 (N_2746,N_1419,N_1798);
nor U2747 (N_2747,N_2295,N_1906);
xnor U2748 (N_2748,N_1248,N_1819);
nand U2749 (N_2749,N_1842,N_2391);
or U2750 (N_2750,N_1617,N_1692);
and U2751 (N_2751,N_1986,N_1210);
xnor U2752 (N_2752,N_2346,N_2331);
nand U2753 (N_2753,N_1339,N_1368);
or U2754 (N_2754,N_1896,N_1452);
nand U2755 (N_2755,N_1917,N_1227);
nand U2756 (N_2756,N_1847,N_2265);
nand U2757 (N_2757,N_1808,N_2058);
nand U2758 (N_2758,N_2074,N_1583);
xnor U2759 (N_2759,N_2047,N_1213);
nor U2760 (N_2760,N_2066,N_1214);
nor U2761 (N_2761,N_2125,N_2357);
nor U2762 (N_2762,N_1374,N_1825);
nor U2763 (N_2763,N_2027,N_1351);
nand U2764 (N_2764,N_1211,N_1400);
xor U2765 (N_2765,N_1758,N_2068);
nor U2766 (N_2766,N_2275,N_1482);
nand U2767 (N_2767,N_1612,N_1464);
xnor U2768 (N_2768,N_1793,N_2023);
or U2769 (N_2769,N_1796,N_1507);
nor U2770 (N_2770,N_1519,N_2373);
nand U2771 (N_2771,N_2249,N_1859);
nor U2772 (N_2772,N_1948,N_2354);
xor U2773 (N_2773,N_2197,N_2377);
nor U2774 (N_2774,N_1851,N_1225);
nand U2775 (N_2775,N_1835,N_1998);
nand U2776 (N_2776,N_2173,N_1281);
nand U2777 (N_2777,N_1759,N_2210);
nor U2778 (N_2778,N_2030,N_2213);
and U2779 (N_2779,N_2332,N_1782);
nor U2780 (N_2780,N_1955,N_1337);
xnor U2781 (N_2781,N_1888,N_2157);
and U2782 (N_2782,N_2231,N_1679);
nor U2783 (N_2783,N_1788,N_1597);
nand U2784 (N_2784,N_1785,N_1933);
and U2785 (N_2785,N_2024,N_1600);
nor U2786 (N_2786,N_1974,N_1291);
nor U2787 (N_2787,N_1993,N_1487);
nand U2788 (N_2788,N_2202,N_2093);
nor U2789 (N_2789,N_1934,N_1949);
and U2790 (N_2790,N_1326,N_2091);
and U2791 (N_2791,N_2004,N_1505);
nand U2792 (N_2792,N_1734,N_1417);
or U2793 (N_2793,N_2070,N_1604);
or U2794 (N_2794,N_2029,N_2368);
nor U2795 (N_2795,N_1255,N_2313);
nor U2796 (N_2796,N_2199,N_1642);
and U2797 (N_2797,N_1857,N_1967);
xnor U2798 (N_2798,N_1787,N_2300);
nand U2799 (N_2799,N_2101,N_1935);
or U2800 (N_2800,N_1674,N_2337);
nor U2801 (N_2801,N_1322,N_1635);
nor U2802 (N_2802,N_1422,N_2060);
and U2803 (N_2803,N_1340,N_1821);
and U2804 (N_2804,N_1496,N_1962);
xor U2805 (N_2805,N_1976,N_2358);
or U2806 (N_2806,N_1494,N_2284);
nor U2807 (N_2807,N_2355,N_2399);
nand U2808 (N_2808,N_2065,N_2028);
xnor U2809 (N_2809,N_2104,N_2097);
nor U2810 (N_2810,N_2165,N_1420);
nand U2811 (N_2811,N_2082,N_1253);
nor U2812 (N_2812,N_1304,N_2364);
and U2813 (N_2813,N_1513,N_1526);
xnor U2814 (N_2814,N_1614,N_1850);
nand U2815 (N_2815,N_1659,N_1672);
or U2816 (N_2816,N_1665,N_2018);
nor U2817 (N_2817,N_1866,N_1837);
or U2818 (N_2818,N_2136,N_1797);
xnor U2819 (N_2819,N_1661,N_2037);
and U2820 (N_2820,N_2268,N_1760);
xnor U2821 (N_2821,N_1506,N_2064);
and U2822 (N_2822,N_2072,N_1231);
and U2823 (N_2823,N_2181,N_1754);
or U2824 (N_2824,N_1228,N_1331);
or U2825 (N_2825,N_1297,N_1473);
and U2826 (N_2826,N_1987,N_1830);
xnor U2827 (N_2827,N_1953,N_1855);
or U2828 (N_2828,N_1903,N_1722);
or U2829 (N_2829,N_1347,N_1570);
and U2830 (N_2830,N_1510,N_1816);
nand U2831 (N_2831,N_2360,N_2098);
or U2832 (N_2832,N_2195,N_1320);
and U2833 (N_2833,N_1670,N_1832);
or U2834 (N_2834,N_2038,N_2352);
xor U2835 (N_2835,N_1550,N_2050);
xnor U2836 (N_2836,N_1465,N_1517);
xor U2837 (N_2837,N_2042,N_1479);
nand U2838 (N_2838,N_1538,N_2280);
nor U2839 (N_2839,N_1412,N_1845);
or U2840 (N_2840,N_2100,N_1936);
nand U2841 (N_2841,N_1242,N_1350);
nor U2842 (N_2842,N_1899,N_1432);
nor U2843 (N_2843,N_1546,N_1310);
and U2844 (N_2844,N_1909,N_1769);
xnor U2845 (N_2845,N_1388,N_1431);
and U2846 (N_2846,N_1682,N_1733);
xor U2847 (N_2847,N_1908,N_1912);
and U2848 (N_2848,N_1972,N_1348);
nand U2849 (N_2849,N_1700,N_1235);
or U2850 (N_2850,N_1778,N_1861);
and U2851 (N_2851,N_2293,N_1889);
nand U2852 (N_2852,N_1762,N_2075);
or U2853 (N_2853,N_1714,N_2109);
or U2854 (N_2854,N_1421,N_1272);
nor U2855 (N_2855,N_2342,N_2270);
and U2856 (N_2856,N_1805,N_1559);
nor U2857 (N_2857,N_2119,N_1939);
or U2858 (N_2858,N_1894,N_1273);
or U2859 (N_2859,N_1610,N_2147);
and U2860 (N_2860,N_1723,N_1436);
nor U2861 (N_2861,N_1755,N_2055);
and U2862 (N_2862,N_1702,N_1440);
nor U2863 (N_2863,N_1915,N_1927);
nand U2864 (N_2864,N_1391,N_1569);
or U2865 (N_2865,N_1444,N_1707);
or U2866 (N_2866,N_1512,N_2216);
or U2867 (N_2867,N_1956,N_2162);
xor U2868 (N_2868,N_1557,N_1303);
or U2869 (N_2869,N_1994,N_1704);
nor U2870 (N_2870,N_1711,N_1833);
nor U2871 (N_2871,N_1403,N_1869);
nand U2872 (N_2872,N_2106,N_1233);
xor U2873 (N_2873,N_1267,N_1946);
nand U2874 (N_2874,N_1828,N_2347);
xor U2875 (N_2875,N_2033,N_2168);
or U2876 (N_2876,N_2245,N_1524);
nor U2877 (N_2877,N_1649,N_2117);
nor U2878 (N_2878,N_2232,N_1645);
and U2879 (N_2879,N_1264,N_1878);
xor U2880 (N_2880,N_1767,N_1375);
or U2881 (N_2881,N_2150,N_1203);
and U2882 (N_2882,N_2163,N_1648);
or U2883 (N_2883,N_2176,N_1705);
and U2884 (N_2884,N_1922,N_2287);
and U2885 (N_2885,N_1865,N_2063);
or U2886 (N_2886,N_1397,N_1453);
and U2887 (N_2887,N_1306,N_2236);
and U2888 (N_2888,N_1675,N_1770);
xor U2889 (N_2889,N_2115,N_2304);
nand U2890 (N_2890,N_2223,N_2316);
and U2891 (N_2891,N_1925,N_1719);
or U2892 (N_2892,N_1727,N_1926);
nand U2893 (N_2893,N_1477,N_1599);
xor U2894 (N_2894,N_1563,N_1230);
or U2895 (N_2895,N_1621,N_1739);
and U2896 (N_2896,N_1892,N_2138);
nor U2897 (N_2897,N_1803,N_1499);
or U2898 (N_2898,N_1841,N_1262);
or U2899 (N_2899,N_1485,N_1279);
xnor U2900 (N_2900,N_2141,N_1467);
or U2901 (N_2901,N_1565,N_1382);
nor U2902 (N_2902,N_2003,N_1238);
nand U2903 (N_2903,N_2116,N_1791);
xor U2904 (N_2904,N_2019,N_1910);
or U2905 (N_2905,N_1472,N_1370);
nand U2906 (N_2906,N_2219,N_1698);
nand U2907 (N_2907,N_1429,N_1633);
nor U2908 (N_2908,N_1216,N_2076);
and U2909 (N_2909,N_1200,N_2204);
or U2910 (N_2910,N_2253,N_1531);
or U2911 (N_2911,N_2330,N_1813);
nand U2912 (N_2912,N_2112,N_1361);
nand U2913 (N_2913,N_2321,N_1831);
xor U2914 (N_2914,N_1408,N_1680);
nor U2915 (N_2915,N_1622,N_2266);
or U2916 (N_2916,N_1662,N_2343);
nor U2917 (N_2917,N_2052,N_1781);
nor U2918 (N_2918,N_2395,N_2379);
xnor U2919 (N_2919,N_1428,N_1664);
nor U2920 (N_2920,N_1495,N_1471);
nor U2921 (N_2921,N_1923,N_1551);
or U2922 (N_2922,N_1441,N_1585);
and U2923 (N_2923,N_1656,N_1653);
nor U2924 (N_2924,N_1406,N_1607);
and U2925 (N_2925,N_1344,N_2051);
or U2926 (N_2926,N_1921,N_1970);
and U2927 (N_2927,N_1263,N_2171);
or U2928 (N_2928,N_1988,N_1489);
nand U2929 (N_2929,N_1630,N_1884);
xnor U2930 (N_2930,N_1689,N_1498);
nor U2931 (N_2931,N_1414,N_2002);
nand U2932 (N_2932,N_1655,N_1282);
xor U2933 (N_2933,N_1686,N_1678);
and U2934 (N_2934,N_1358,N_2328);
nand U2935 (N_2935,N_1737,N_1332);
xor U2936 (N_2936,N_1768,N_1629);
nand U2937 (N_2937,N_1295,N_1800);
xor U2938 (N_2938,N_1276,N_1260);
nor U2939 (N_2939,N_1409,N_1611);
nand U2940 (N_2940,N_2351,N_1699);
and U2941 (N_2941,N_1504,N_2022);
nor U2942 (N_2942,N_2329,N_2108);
or U2943 (N_2943,N_2340,N_2315);
nor U2944 (N_2944,N_2324,N_1749);
or U2945 (N_2945,N_2126,N_2260);
nand U2946 (N_2946,N_1965,N_1547);
nor U2947 (N_2947,N_2307,N_2305);
and U2948 (N_2948,N_1886,N_1637);
xnor U2949 (N_2949,N_1386,N_2175);
nor U2950 (N_2950,N_1292,N_1312);
or U2951 (N_2951,N_1363,N_2217);
or U2952 (N_2952,N_1897,N_1439);
or U2953 (N_2953,N_1237,N_1562);
nor U2954 (N_2954,N_1757,N_1773);
or U2955 (N_2955,N_1315,N_1470);
nand U2956 (N_2956,N_1369,N_2320);
or U2957 (N_2957,N_1804,N_2257);
and U2958 (N_2958,N_1490,N_1338);
xor U2959 (N_2959,N_1219,N_2174);
and U2960 (N_2960,N_2264,N_2067);
nand U2961 (N_2961,N_1824,N_1516);
nand U2962 (N_2962,N_2272,N_2396);
and U2963 (N_2963,N_2278,N_1763);
xor U2964 (N_2964,N_1658,N_1514);
xnor U2965 (N_2965,N_1846,N_1900);
nor U2966 (N_2966,N_1904,N_1342);
nor U2967 (N_2967,N_2235,N_2365);
and U2968 (N_2968,N_2144,N_1293);
nor U2969 (N_2969,N_2182,N_1764);
and U2970 (N_2970,N_1356,N_1423);
or U2971 (N_2971,N_2256,N_1601);
or U2972 (N_2972,N_1548,N_1995);
nand U2973 (N_2973,N_1217,N_1558);
or U2974 (N_2974,N_2122,N_1815);
or U2975 (N_2975,N_2184,N_1801);
xor U2976 (N_2976,N_1301,N_1278);
and U2977 (N_2977,N_1814,N_2036);
or U2978 (N_2978,N_1323,N_1996);
and U2979 (N_2979,N_1747,N_2292);
nand U2980 (N_2980,N_1882,N_1875);
nor U2981 (N_2981,N_1738,N_2229);
and U2982 (N_2982,N_1618,N_1385);
or U2983 (N_2983,N_2095,N_1893);
nand U2984 (N_2984,N_1744,N_1329);
or U2985 (N_2985,N_2187,N_1834);
nand U2986 (N_2986,N_1666,N_1327);
xor U2987 (N_2987,N_1268,N_2086);
nor U2988 (N_2988,N_1362,N_1957);
or U2989 (N_2989,N_1413,N_2350);
or U2990 (N_2990,N_1254,N_1480);
nor U2991 (N_2991,N_2089,N_1398);
nor U2992 (N_2992,N_2276,N_1221);
or U2993 (N_2993,N_2289,N_2035);
xor U2994 (N_2994,N_2356,N_1518);
or U2995 (N_2995,N_2243,N_1802);
and U2996 (N_2996,N_1521,N_1288);
nor U2997 (N_2997,N_2143,N_2291);
and U2998 (N_2998,N_1991,N_1720);
nor U2999 (N_2999,N_1345,N_1437);
or U3000 (N_3000,N_2052,N_1404);
nor U3001 (N_3001,N_1768,N_1778);
nand U3002 (N_3002,N_1948,N_2088);
nor U3003 (N_3003,N_2332,N_2011);
and U3004 (N_3004,N_2352,N_1238);
xor U3005 (N_3005,N_2195,N_1996);
and U3006 (N_3006,N_2050,N_1853);
or U3007 (N_3007,N_1863,N_1204);
nand U3008 (N_3008,N_2215,N_1666);
xnor U3009 (N_3009,N_1490,N_1624);
xnor U3010 (N_3010,N_1335,N_1446);
xor U3011 (N_3011,N_2061,N_1517);
or U3012 (N_3012,N_1277,N_1287);
nor U3013 (N_3013,N_2006,N_2106);
xor U3014 (N_3014,N_1292,N_1860);
nor U3015 (N_3015,N_1497,N_1440);
nand U3016 (N_3016,N_1277,N_1278);
or U3017 (N_3017,N_1711,N_2239);
xor U3018 (N_3018,N_2034,N_2364);
and U3019 (N_3019,N_2198,N_2066);
nand U3020 (N_3020,N_1464,N_1686);
nand U3021 (N_3021,N_2060,N_2180);
nor U3022 (N_3022,N_1530,N_2269);
xnor U3023 (N_3023,N_1886,N_1883);
nand U3024 (N_3024,N_1643,N_1887);
and U3025 (N_3025,N_1906,N_2350);
nand U3026 (N_3026,N_1613,N_2157);
nand U3027 (N_3027,N_1975,N_2363);
nor U3028 (N_3028,N_2028,N_1908);
or U3029 (N_3029,N_1651,N_1349);
nor U3030 (N_3030,N_2224,N_2055);
or U3031 (N_3031,N_1225,N_1344);
nor U3032 (N_3032,N_1644,N_1939);
xnor U3033 (N_3033,N_1207,N_2373);
nand U3034 (N_3034,N_1430,N_2344);
or U3035 (N_3035,N_1953,N_2175);
xnor U3036 (N_3036,N_1474,N_2319);
and U3037 (N_3037,N_2285,N_1480);
and U3038 (N_3038,N_1938,N_2253);
and U3039 (N_3039,N_2210,N_1905);
nor U3040 (N_3040,N_2025,N_1755);
and U3041 (N_3041,N_1584,N_2032);
or U3042 (N_3042,N_2157,N_1924);
xor U3043 (N_3043,N_2370,N_1945);
xnor U3044 (N_3044,N_1777,N_1538);
and U3045 (N_3045,N_1693,N_1688);
or U3046 (N_3046,N_1737,N_1620);
nand U3047 (N_3047,N_2115,N_1729);
xnor U3048 (N_3048,N_2265,N_1279);
or U3049 (N_3049,N_1831,N_1498);
nand U3050 (N_3050,N_1654,N_1427);
or U3051 (N_3051,N_1292,N_2080);
xor U3052 (N_3052,N_2324,N_1658);
nor U3053 (N_3053,N_1779,N_1265);
xnor U3054 (N_3054,N_1289,N_1824);
nand U3055 (N_3055,N_2139,N_1324);
nand U3056 (N_3056,N_2034,N_1777);
and U3057 (N_3057,N_1598,N_1859);
xnor U3058 (N_3058,N_1654,N_1716);
and U3059 (N_3059,N_2194,N_2270);
nor U3060 (N_3060,N_1216,N_1779);
nand U3061 (N_3061,N_1661,N_1885);
nor U3062 (N_3062,N_1750,N_2388);
nand U3063 (N_3063,N_1487,N_1441);
nand U3064 (N_3064,N_1203,N_1594);
nand U3065 (N_3065,N_1704,N_1625);
nand U3066 (N_3066,N_2305,N_1623);
xnor U3067 (N_3067,N_1329,N_1447);
nor U3068 (N_3068,N_1716,N_1916);
nor U3069 (N_3069,N_1911,N_1550);
xor U3070 (N_3070,N_1960,N_1403);
nor U3071 (N_3071,N_1595,N_2321);
nand U3072 (N_3072,N_1552,N_2128);
nor U3073 (N_3073,N_1995,N_2178);
or U3074 (N_3074,N_2258,N_1553);
nor U3075 (N_3075,N_1625,N_2347);
xnor U3076 (N_3076,N_2207,N_2295);
nand U3077 (N_3077,N_2292,N_2003);
and U3078 (N_3078,N_2291,N_1874);
nor U3079 (N_3079,N_1315,N_2036);
and U3080 (N_3080,N_1849,N_2392);
xnor U3081 (N_3081,N_2334,N_1212);
or U3082 (N_3082,N_1901,N_1207);
nand U3083 (N_3083,N_1802,N_2321);
nand U3084 (N_3084,N_1616,N_1939);
or U3085 (N_3085,N_1238,N_1387);
nand U3086 (N_3086,N_1675,N_2035);
nand U3087 (N_3087,N_1212,N_1765);
and U3088 (N_3088,N_2379,N_1591);
and U3089 (N_3089,N_1764,N_2039);
and U3090 (N_3090,N_1607,N_2118);
nor U3091 (N_3091,N_2344,N_1957);
nand U3092 (N_3092,N_2109,N_1434);
and U3093 (N_3093,N_1459,N_1386);
and U3094 (N_3094,N_2081,N_2170);
and U3095 (N_3095,N_2105,N_1985);
and U3096 (N_3096,N_1383,N_2010);
or U3097 (N_3097,N_1713,N_2140);
xnor U3098 (N_3098,N_1627,N_1789);
xor U3099 (N_3099,N_2007,N_1306);
and U3100 (N_3100,N_1469,N_1263);
nand U3101 (N_3101,N_1358,N_1272);
nand U3102 (N_3102,N_2067,N_1494);
xnor U3103 (N_3103,N_2258,N_2255);
and U3104 (N_3104,N_1763,N_1677);
nand U3105 (N_3105,N_1785,N_1439);
nand U3106 (N_3106,N_2147,N_1655);
and U3107 (N_3107,N_2067,N_1893);
nor U3108 (N_3108,N_1441,N_2214);
and U3109 (N_3109,N_1394,N_2329);
and U3110 (N_3110,N_2251,N_1371);
and U3111 (N_3111,N_1905,N_1468);
or U3112 (N_3112,N_2166,N_1483);
nand U3113 (N_3113,N_1763,N_1424);
or U3114 (N_3114,N_1462,N_2176);
or U3115 (N_3115,N_1351,N_1421);
or U3116 (N_3116,N_2152,N_1433);
and U3117 (N_3117,N_2257,N_1216);
or U3118 (N_3118,N_1733,N_1667);
nor U3119 (N_3119,N_2010,N_2160);
or U3120 (N_3120,N_1526,N_1880);
and U3121 (N_3121,N_1946,N_1488);
nor U3122 (N_3122,N_1586,N_1264);
nor U3123 (N_3123,N_1881,N_1517);
nand U3124 (N_3124,N_2259,N_1226);
or U3125 (N_3125,N_1789,N_1449);
nand U3126 (N_3126,N_1915,N_2206);
nor U3127 (N_3127,N_2093,N_1210);
xor U3128 (N_3128,N_1615,N_2129);
nand U3129 (N_3129,N_1417,N_1563);
nand U3130 (N_3130,N_1553,N_2358);
nor U3131 (N_3131,N_1260,N_1538);
and U3132 (N_3132,N_1917,N_1900);
nor U3133 (N_3133,N_2389,N_1347);
or U3134 (N_3134,N_1354,N_2014);
nor U3135 (N_3135,N_2341,N_2034);
or U3136 (N_3136,N_1367,N_1404);
xnor U3137 (N_3137,N_2077,N_2398);
and U3138 (N_3138,N_1256,N_1237);
or U3139 (N_3139,N_2350,N_1308);
xnor U3140 (N_3140,N_1700,N_1560);
or U3141 (N_3141,N_2108,N_1979);
nand U3142 (N_3142,N_1269,N_1552);
or U3143 (N_3143,N_1754,N_1662);
or U3144 (N_3144,N_2164,N_1646);
xnor U3145 (N_3145,N_1639,N_2282);
xnor U3146 (N_3146,N_1262,N_2297);
nand U3147 (N_3147,N_1837,N_2076);
xnor U3148 (N_3148,N_1447,N_2318);
nor U3149 (N_3149,N_2116,N_1689);
or U3150 (N_3150,N_2218,N_1580);
nand U3151 (N_3151,N_1828,N_2067);
and U3152 (N_3152,N_1419,N_1487);
or U3153 (N_3153,N_1463,N_1704);
nand U3154 (N_3154,N_1871,N_2095);
nor U3155 (N_3155,N_1984,N_1278);
nand U3156 (N_3156,N_2242,N_1305);
xnor U3157 (N_3157,N_1695,N_1376);
nor U3158 (N_3158,N_2278,N_1923);
or U3159 (N_3159,N_2390,N_1838);
nor U3160 (N_3160,N_1276,N_1214);
and U3161 (N_3161,N_2295,N_2385);
xnor U3162 (N_3162,N_2391,N_1305);
and U3163 (N_3163,N_1434,N_2284);
and U3164 (N_3164,N_1797,N_1437);
or U3165 (N_3165,N_1291,N_1640);
nand U3166 (N_3166,N_2131,N_1914);
xor U3167 (N_3167,N_2184,N_2291);
xor U3168 (N_3168,N_1800,N_1783);
nor U3169 (N_3169,N_1531,N_1670);
nor U3170 (N_3170,N_1760,N_1729);
or U3171 (N_3171,N_2184,N_1807);
xnor U3172 (N_3172,N_1802,N_2135);
nand U3173 (N_3173,N_1446,N_2338);
nor U3174 (N_3174,N_1797,N_1218);
nand U3175 (N_3175,N_1923,N_2226);
nand U3176 (N_3176,N_1474,N_2397);
nor U3177 (N_3177,N_1437,N_1843);
and U3178 (N_3178,N_2036,N_2370);
xor U3179 (N_3179,N_2365,N_1822);
or U3180 (N_3180,N_1334,N_1326);
xor U3181 (N_3181,N_1270,N_2152);
or U3182 (N_3182,N_2020,N_2383);
and U3183 (N_3183,N_1691,N_1669);
or U3184 (N_3184,N_2044,N_1346);
or U3185 (N_3185,N_1704,N_1851);
xor U3186 (N_3186,N_1991,N_2176);
nand U3187 (N_3187,N_2249,N_1873);
or U3188 (N_3188,N_1310,N_1799);
nand U3189 (N_3189,N_2057,N_1322);
xor U3190 (N_3190,N_1472,N_1975);
nand U3191 (N_3191,N_1419,N_2321);
nor U3192 (N_3192,N_2196,N_2301);
or U3193 (N_3193,N_1485,N_2249);
and U3194 (N_3194,N_2302,N_2387);
xor U3195 (N_3195,N_2264,N_1315);
or U3196 (N_3196,N_1481,N_1885);
nor U3197 (N_3197,N_1291,N_1825);
and U3198 (N_3198,N_1693,N_1459);
nand U3199 (N_3199,N_1872,N_1457);
nor U3200 (N_3200,N_2378,N_1269);
nor U3201 (N_3201,N_2211,N_1225);
nor U3202 (N_3202,N_1954,N_1362);
or U3203 (N_3203,N_2343,N_1571);
xor U3204 (N_3204,N_1459,N_1474);
xor U3205 (N_3205,N_2241,N_1647);
or U3206 (N_3206,N_1329,N_2262);
xor U3207 (N_3207,N_1500,N_1392);
nand U3208 (N_3208,N_1475,N_1992);
or U3209 (N_3209,N_1857,N_1240);
nand U3210 (N_3210,N_1266,N_2038);
or U3211 (N_3211,N_1581,N_1526);
nand U3212 (N_3212,N_2024,N_2015);
nand U3213 (N_3213,N_2098,N_2012);
nand U3214 (N_3214,N_1763,N_1979);
or U3215 (N_3215,N_1343,N_1355);
and U3216 (N_3216,N_1294,N_1627);
and U3217 (N_3217,N_1539,N_1685);
nor U3218 (N_3218,N_2316,N_1966);
and U3219 (N_3219,N_2264,N_1437);
or U3220 (N_3220,N_1667,N_2255);
xor U3221 (N_3221,N_1554,N_2294);
nor U3222 (N_3222,N_2050,N_1434);
nand U3223 (N_3223,N_1742,N_1460);
or U3224 (N_3224,N_1730,N_2030);
or U3225 (N_3225,N_1209,N_2199);
nand U3226 (N_3226,N_1851,N_2237);
and U3227 (N_3227,N_1610,N_1955);
xor U3228 (N_3228,N_1947,N_1991);
nor U3229 (N_3229,N_2013,N_1417);
or U3230 (N_3230,N_1515,N_1269);
or U3231 (N_3231,N_1438,N_1885);
nand U3232 (N_3232,N_1386,N_1632);
and U3233 (N_3233,N_1341,N_1922);
or U3234 (N_3234,N_2307,N_1896);
or U3235 (N_3235,N_2382,N_1645);
and U3236 (N_3236,N_1395,N_2068);
or U3237 (N_3237,N_1969,N_1688);
xor U3238 (N_3238,N_1884,N_1996);
xor U3239 (N_3239,N_1554,N_1380);
or U3240 (N_3240,N_2003,N_1654);
nand U3241 (N_3241,N_1368,N_2002);
nor U3242 (N_3242,N_1687,N_1587);
nand U3243 (N_3243,N_2360,N_1353);
and U3244 (N_3244,N_1742,N_2297);
nand U3245 (N_3245,N_2371,N_1392);
and U3246 (N_3246,N_1910,N_2203);
nand U3247 (N_3247,N_2008,N_1501);
xnor U3248 (N_3248,N_1720,N_1826);
or U3249 (N_3249,N_2252,N_1257);
nand U3250 (N_3250,N_1989,N_1379);
nand U3251 (N_3251,N_2012,N_1271);
xor U3252 (N_3252,N_2228,N_1707);
nand U3253 (N_3253,N_2392,N_2062);
and U3254 (N_3254,N_1994,N_1684);
or U3255 (N_3255,N_1224,N_1679);
nand U3256 (N_3256,N_1996,N_1292);
xor U3257 (N_3257,N_1793,N_1708);
and U3258 (N_3258,N_1521,N_2005);
nor U3259 (N_3259,N_1509,N_1611);
or U3260 (N_3260,N_1243,N_1436);
and U3261 (N_3261,N_2279,N_2327);
nor U3262 (N_3262,N_1741,N_2232);
nor U3263 (N_3263,N_1682,N_2011);
xor U3264 (N_3264,N_2218,N_1221);
or U3265 (N_3265,N_1333,N_2185);
nor U3266 (N_3266,N_2187,N_1563);
nand U3267 (N_3267,N_1254,N_1921);
or U3268 (N_3268,N_1832,N_1312);
nand U3269 (N_3269,N_2274,N_1950);
and U3270 (N_3270,N_1863,N_2064);
and U3271 (N_3271,N_1770,N_2002);
or U3272 (N_3272,N_2169,N_1931);
xnor U3273 (N_3273,N_1433,N_2112);
nand U3274 (N_3274,N_2214,N_2328);
nand U3275 (N_3275,N_1800,N_1951);
or U3276 (N_3276,N_1775,N_1923);
and U3277 (N_3277,N_2197,N_1790);
nor U3278 (N_3278,N_1944,N_1514);
and U3279 (N_3279,N_2104,N_2023);
nand U3280 (N_3280,N_1502,N_1744);
nor U3281 (N_3281,N_1769,N_1637);
xnor U3282 (N_3282,N_1263,N_2152);
nor U3283 (N_3283,N_1780,N_2288);
nor U3284 (N_3284,N_2233,N_1264);
xnor U3285 (N_3285,N_1842,N_1920);
and U3286 (N_3286,N_1822,N_1533);
nand U3287 (N_3287,N_2216,N_1821);
nand U3288 (N_3288,N_1279,N_1799);
or U3289 (N_3289,N_1683,N_1849);
and U3290 (N_3290,N_1610,N_2356);
or U3291 (N_3291,N_2345,N_1638);
and U3292 (N_3292,N_1304,N_2000);
nor U3293 (N_3293,N_1930,N_1586);
xnor U3294 (N_3294,N_2070,N_1335);
xor U3295 (N_3295,N_1977,N_1257);
nor U3296 (N_3296,N_1516,N_1858);
xor U3297 (N_3297,N_2033,N_1811);
xnor U3298 (N_3298,N_2107,N_1813);
xor U3299 (N_3299,N_1788,N_1449);
xnor U3300 (N_3300,N_2135,N_1514);
and U3301 (N_3301,N_1445,N_1854);
nand U3302 (N_3302,N_1364,N_1453);
and U3303 (N_3303,N_1629,N_2129);
nor U3304 (N_3304,N_1808,N_1681);
nand U3305 (N_3305,N_1354,N_2287);
xor U3306 (N_3306,N_1849,N_1975);
nand U3307 (N_3307,N_1993,N_2057);
nor U3308 (N_3308,N_2180,N_2093);
xnor U3309 (N_3309,N_1381,N_1657);
nand U3310 (N_3310,N_1418,N_2150);
and U3311 (N_3311,N_1462,N_2169);
nand U3312 (N_3312,N_1816,N_1858);
nand U3313 (N_3313,N_2289,N_1736);
xnor U3314 (N_3314,N_1444,N_2302);
nor U3315 (N_3315,N_2236,N_1396);
xnor U3316 (N_3316,N_1712,N_1409);
xnor U3317 (N_3317,N_1638,N_2053);
xor U3318 (N_3318,N_2114,N_1622);
or U3319 (N_3319,N_1219,N_1620);
and U3320 (N_3320,N_1403,N_2329);
nor U3321 (N_3321,N_1999,N_1982);
or U3322 (N_3322,N_1248,N_1411);
or U3323 (N_3323,N_1647,N_1401);
and U3324 (N_3324,N_1916,N_1640);
and U3325 (N_3325,N_1914,N_1899);
and U3326 (N_3326,N_2185,N_1308);
nand U3327 (N_3327,N_1987,N_1985);
and U3328 (N_3328,N_1363,N_2022);
or U3329 (N_3329,N_1710,N_1954);
nor U3330 (N_3330,N_1249,N_1703);
or U3331 (N_3331,N_1210,N_1665);
nand U3332 (N_3332,N_1445,N_1923);
or U3333 (N_3333,N_1595,N_2072);
or U3334 (N_3334,N_1764,N_1897);
and U3335 (N_3335,N_2081,N_2236);
and U3336 (N_3336,N_1852,N_1532);
and U3337 (N_3337,N_1404,N_1354);
and U3338 (N_3338,N_1427,N_1613);
or U3339 (N_3339,N_2224,N_1918);
nor U3340 (N_3340,N_2090,N_1920);
or U3341 (N_3341,N_2215,N_1457);
xnor U3342 (N_3342,N_2031,N_1638);
and U3343 (N_3343,N_2360,N_2125);
and U3344 (N_3344,N_1735,N_2020);
xnor U3345 (N_3345,N_2393,N_2185);
xnor U3346 (N_3346,N_1831,N_2149);
and U3347 (N_3347,N_2234,N_1343);
xor U3348 (N_3348,N_2342,N_1847);
xnor U3349 (N_3349,N_2169,N_1585);
and U3350 (N_3350,N_2213,N_1570);
nand U3351 (N_3351,N_2062,N_2119);
xnor U3352 (N_3352,N_2031,N_1665);
xnor U3353 (N_3353,N_2037,N_1620);
nor U3354 (N_3354,N_2260,N_2181);
xor U3355 (N_3355,N_1836,N_2015);
and U3356 (N_3356,N_2346,N_1434);
xor U3357 (N_3357,N_2229,N_1208);
nor U3358 (N_3358,N_1295,N_1255);
xor U3359 (N_3359,N_1824,N_1823);
and U3360 (N_3360,N_1916,N_1319);
nor U3361 (N_3361,N_1717,N_2181);
or U3362 (N_3362,N_2392,N_1658);
nor U3363 (N_3363,N_1208,N_2319);
nor U3364 (N_3364,N_2180,N_2395);
or U3365 (N_3365,N_1708,N_2166);
nor U3366 (N_3366,N_2067,N_1925);
or U3367 (N_3367,N_1690,N_1718);
nand U3368 (N_3368,N_1912,N_1452);
nand U3369 (N_3369,N_2176,N_1702);
or U3370 (N_3370,N_2205,N_1396);
or U3371 (N_3371,N_2071,N_2027);
nor U3372 (N_3372,N_2391,N_2093);
and U3373 (N_3373,N_1780,N_1526);
nor U3374 (N_3374,N_1356,N_1863);
xnor U3375 (N_3375,N_2219,N_1330);
and U3376 (N_3376,N_2318,N_1602);
nand U3377 (N_3377,N_1963,N_2154);
nand U3378 (N_3378,N_1509,N_1385);
nand U3379 (N_3379,N_2070,N_1976);
nand U3380 (N_3380,N_2146,N_1268);
and U3381 (N_3381,N_1254,N_1922);
and U3382 (N_3382,N_1843,N_1849);
nand U3383 (N_3383,N_1984,N_2069);
and U3384 (N_3384,N_1273,N_2305);
and U3385 (N_3385,N_1538,N_1818);
nand U3386 (N_3386,N_2360,N_1574);
and U3387 (N_3387,N_1612,N_2181);
and U3388 (N_3388,N_1908,N_1446);
and U3389 (N_3389,N_2245,N_1782);
nor U3390 (N_3390,N_1303,N_2153);
or U3391 (N_3391,N_2233,N_1523);
nor U3392 (N_3392,N_2095,N_1343);
and U3393 (N_3393,N_1835,N_2317);
nor U3394 (N_3394,N_2235,N_1848);
and U3395 (N_3395,N_1338,N_1917);
xnor U3396 (N_3396,N_2228,N_1273);
nand U3397 (N_3397,N_1559,N_1467);
nand U3398 (N_3398,N_2234,N_1335);
xor U3399 (N_3399,N_2389,N_1751);
xnor U3400 (N_3400,N_2215,N_1665);
and U3401 (N_3401,N_2393,N_1644);
or U3402 (N_3402,N_2367,N_1714);
or U3403 (N_3403,N_2162,N_1838);
nor U3404 (N_3404,N_1414,N_1485);
nor U3405 (N_3405,N_2041,N_2115);
nor U3406 (N_3406,N_2181,N_1664);
nor U3407 (N_3407,N_1712,N_1496);
or U3408 (N_3408,N_2230,N_1842);
xor U3409 (N_3409,N_1527,N_1329);
xnor U3410 (N_3410,N_1550,N_2010);
nor U3411 (N_3411,N_1901,N_1232);
xor U3412 (N_3412,N_1947,N_1871);
nor U3413 (N_3413,N_2258,N_1309);
nand U3414 (N_3414,N_1322,N_1856);
nor U3415 (N_3415,N_1796,N_2174);
or U3416 (N_3416,N_1403,N_1458);
xor U3417 (N_3417,N_1241,N_1461);
or U3418 (N_3418,N_1868,N_2376);
nand U3419 (N_3419,N_1911,N_1850);
nor U3420 (N_3420,N_1673,N_1711);
nand U3421 (N_3421,N_1921,N_1605);
and U3422 (N_3422,N_2382,N_2364);
nand U3423 (N_3423,N_2395,N_2272);
xor U3424 (N_3424,N_1575,N_1411);
xor U3425 (N_3425,N_1277,N_1641);
nor U3426 (N_3426,N_1502,N_1309);
xnor U3427 (N_3427,N_1256,N_1659);
nor U3428 (N_3428,N_2395,N_2212);
nand U3429 (N_3429,N_2141,N_1563);
or U3430 (N_3430,N_1574,N_1642);
nor U3431 (N_3431,N_1662,N_2207);
or U3432 (N_3432,N_1628,N_1644);
xor U3433 (N_3433,N_1499,N_1331);
xnor U3434 (N_3434,N_2306,N_1890);
or U3435 (N_3435,N_1951,N_1881);
and U3436 (N_3436,N_1555,N_1658);
and U3437 (N_3437,N_2378,N_2184);
and U3438 (N_3438,N_1554,N_2196);
or U3439 (N_3439,N_1348,N_2346);
or U3440 (N_3440,N_1730,N_1787);
nand U3441 (N_3441,N_1484,N_1332);
nand U3442 (N_3442,N_1938,N_1987);
and U3443 (N_3443,N_1575,N_1393);
or U3444 (N_3444,N_1547,N_1379);
xnor U3445 (N_3445,N_1391,N_2310);
xnor U3446 (N_3446,N_1684,N_1243);
nand U3447 (N_3447,N_1280,N_1598);
nor U3448 (N_3448,N_2316,N_1547);
nand U3449 (N_3449,N_2386,N_1402);
nand U3450 (N_3450,N_2088,N_2373);
nor U3451 (N_3451,N_1715,N_2382);
nand U3452 (N_3452,N_1529,N_2372);
nand U3453 (N_3453,N_1934,N_1768);
or U3454 (N_3454,N_2356,N_1858);
nand U3455 (N_3455,N_2331,N_1502);
nor U3456 (N_3456,N_2323,N_1721);
nand U3457 (N_3457,N_1740,N_1767);
xor U3458 (N_3458,N_1397,N_2225);
nor U3459 (N_3459,N_2109,N_1546);
nor U3460 (N_3460,N_1571,N_1608);
nor U3461 (N_3461,N_2207,N_1654);
nand U3462 (N_3462,N_1749,N_1955);
nor U3463 (N_3463,N_1368,N_1993);
nand U3464 (N_3464,N_1714,N_1923);
and U3465 (N_3465,N_1253,N_1232);
nand U3466 (N_3466,N_2099,N_1518);
nand U3467 (N_3467,N_1308,N_1447);
nand U3468 (N_3468,N_1556,N_1729);
nor U3469 (N_3469,N_1260,N_2028);
nor U3470 (N_3470,N_1848,N_1367);
nand U3471 (N_3471,N_1360,N_1827);
nand U3472 (N_3472,N_1291,N_1511);
and U3473 (N_3473,N_1543,N_1572);
and U3474 (N_3474,N_2139,N_2343);
or U3475 (N_3475,N_1696,N_1456);
and U3476 (N_3476,N_2266,N_1956);
or U3477 (N_3477,N_2290,N_1834);
nor U3478 (N_3478,N_1464,N_2264);
and U3479 (N_3479,N_2280,N_1504);
and U3480 (N_3480,N_2210,N_1598);
nand U3481 (N_3481,N_1323,N_1725);
nand U3482 (N_3482,N_1623,N_2396);
nand U3483 (N_3483,N_2130,N_1789);
and U3484 (N_3484,N_1487,N_2302);
nor U3485 (N_3485,N_2158,N_1754);
and U3486 (N_3486,N_1270,N_2305);
or U3487 (N_3487,N_1588,N_1910);
and U3488 (N_3488,N_1982,N_1947);
xor U3489 (N_3489,N_1966,N_2021);
and U3490 (N_3490,N_1336,N_1726);
nand U3491 (N_3491,N_2386,N_1639);
or U3492 (N_3492,N_2243,N_1306);
xor U3493 (N_3493,N_1930,N_1217);
and U3494 (N_3494,N_2045,N_1545);
and U3495 (N_3495,N_1733,N_1599);
nand U3496 (N_3496,N_2093,N_2016);
xnor U3497 (N_3497,N_2240,N_1554);
or U3498 (N_3498,N_1911,N_2347);
and U3499 (N_3499,N_1276,N_1307);
or U3500 (N_3500,N_1644,N_1852);
xnor U3501 (N_3501,N_1661,N_1515);
nand U3502 (N_3502,N_1458,N_1908);
and U3503 (N_3503,N_2331,N_1888);
xor U3504 (N_3504,N_2187,N_1472);
or U3505 (N_3505,N_1924,N_1975);
nand U3506 (N_3506,N_1957,N_1395);
xor U3507 (N_3507,N_2285,N_1226);
and U3508 (N_3508,N_1353,N_1982);
and U3509 (N_3509,N_2052,N_2057);
nand U3510 (N_3510,N_2062,N_1547);
nand U3511 (N_3511,N_2272,N_2286);
or U3512 (N_3512,N_2114,N_2159);
xor U3513 (N_3513,N_2163,N_1550);
and U3514 (N_3514,N_2394,N_1960);
nor U3515 (N_3515,N_1401,N_1989);
or U3516 (N_3516,N_1798,N_1883);
nand U3517 (N_3517,N_2376,N_2277);
and U3518 (N_3518,N_1569,N_1653);
nor U3519 (N_3519,N_1337,N_1342);
or U3520 (N_3520,N_1793,N_2318);
nor U3521 (N_3521,N_1368,N_2192);
or U3522 (N_3522,N_2397,N_1754);
and U3523 (N_3523,N_1724,N_2270);
nand U3524 (N_3524,N_1791,N_2316);
or U3525 (N_3525,N_1541,N_2120);
nand U3526 (N_3526,N_1479,N_1259);
nor U3527 (N_3527,N_2130,N_2226);
nand U3528 (N_3528,N_1676,N_1797);
nand U3529 (N_3529,N_2003,N_1658);
or U3530 (N_3530,N_2047,N_1414);
nand U3531 (N_3531,N_1251,N_2225);
nor U3532 (N_3532,N_2125,N_1738);
xor U3533 (N_3533,N_1392,N_2160);
xor U3534 (N_3534,N_2367,N_2214);
or U3535 (N_3535,N_2070,N_2189);
xnor U3536 (N_3536,N_1901,N_1347);
nor U3537 (N_3537,N_1490,N_2012);
and U3538 (N_3538,N_1408,N_1731);
or U3539 (N_3539,N_1762,N_1469);
or U3540 (N_3540,N_1437,N_1213);
xor U3541 (N_3541,N_1206,N_2068);
or U3542 (N_3542,N_1882,N_2315);
or U3543 (N_3543,N_2364,N_2243);
or U3544 (N_3544,N_2143,N_1833);
nand U3545 (N_3545,N_1896,N_2324);
xnor U3546 (N_3546,N_2146,N_2057);
and U3547 (N_3547,N_1258,N_1900);
nand U3548 (N_3548,N_1470,N_2055);
nor U3549 (N_3549,N_1886,N_1373);
or U3550 (N_3550,N_2318,N_1473);
xnor U3551 (N_3551,N_1750,N_1332);
nor U3552 (N_3552,N_1565,N_2352);
and U3553 (N_3553,N_1420,N_1674);
and U3554 (N_3554,N_1973,N_1454);
and U3555 (N_3555,N_1691,N_1965);
nor U3556 (N_3556,N_1228,N_1954);
nor U3557 (N_3557,N_1604,N_1253);
and U3558 (N_3558,N_1692,N_2346);
xor U3559 (N_3559,N_1620,N_1330);
nor U3560 (N_3560,N_2229,N_1752);
xor U3561 (N_3561,N_2395,N_2224);
nor U3562 (N_3562,N_1703,N_1527);
and U3563 (N_3563,N_1526,N_1738);
or U3564 (N_3564,N_2060,N_2157);
xor U3565 (N_3565,N_2101,N_1680);
and U3566 (N_3566,N_1900,N_1431);
xnor U3567 (N_3567,N_1932,N_1339);
and U3568 (N_3568,N_1569,N_1300);
nand U3569 (N_3569,N_1387,N_1342);
nor U3570 (N_3570,N_1307,N_1466);
and U3571 (N_3571,N_1536,N_2129);
and U3572 (N_3572,N_1969,N_1436);
and U3573 (N_3573,N_2126,N_2097);
nand U3574 (N_3574,N_2187,N_1411);
and U3575 (N_3575,N_1915,N_1612);
and U3576 (N_3576,N_1681,N_2029);
and U3577 (N_3577,N_2104,N_1532);
and U3578 (N_3578,N_1696,N_1548);
xor U3579 (N_3579,N_1674,N_2024);
nor U3580 (N_3580,N_1748,N_1781);
and U3581 (N_3581,N_1756,N_1405);
nand U3582 (N_3582,N_1414,N_2124);
nand U3583 (N_3583,N_1883,N_1254);
nor U3584 (N_3584,N_2069,N_1299);
or U3585 (N_3585,N_2356,N_1612);
xnor U3586 (N_3586,N_2396,N_2206);
nand U3587 (N_3587,N_1558,N_1801);
nand U3588 (N_3588,N_1302,N_2394);
or U3589 (N_3589,N_2379,N_1788);
nand U3590 (N_3590,N_1742,N_2177);
nor U3591 (N_3591,N_1535,N_2151);
xnor U3592 (N_3592,N_1939,N_2210);
or U3593 (N_3593,N_1319,N_1425);
or U3594 (N_3594,N_2297,N_2270);
or U3595 (N_3595,N_1498,N_2081);
nand U3596 (N_3596,N_2390,N_2327);
or U3597 (N_3597,N_1346,N_2078);
or U3598 (N_3598,N_2040,N_1449);
and U3599 (N_3599,N_1959,N_1883);
nand U3600 (N_3600,N_3480,N_2476);
nand U3601 (N_3601,N_3103,N_3573);
and U3602 (N_3602,N_2995,N_2924);
xnor U3603 (N_3603,N_2590,N_2471);
nand U3604 (N_3604,N_2403,N_3385);
or U3605 (N_3605,N_3083,N_3347);
nand U3606 (N_3606,N_2974,N_3412);
or U3607 (N_3607,N_2875,N_2427);
nand U3608 (N_3608,N_3210,N_3309);
and U3609 (N_3609,N_3066,N_3237);
xnor U3610 (N_3610,N_3097,N_2901);
or U3611 (N_3611,N_2543,N_3582);
nand U3612 (N_3612,N_3345,N_2931);
nor U3613 (N_3613,N_3213,N_3516);
and U3614 (N_3614,N_3088,N_2819);
nor U3615 (N_3615,N_2405,N_2447);
nor U3616 (N_3616,N_2404,N_2670);
or U3617 (N_3617,N_2797,N_3110);
and U3618 (N_3618,N_2867,N_2969);
or U3619 (N_3619,N_3553,N_2945);
nand U3620 (N_3620,N_3317,N_2870);
nand U3621 (N_3621,N_2676,N_3521);
xnor U3622 (N_3622,N_2673,N_2849);
nor U3623 (N_3623,N_2705,N_2840);
nand U3624 (N_3624,N_3489,N_2420);
nand U3625 (N_3625,N_2629,N_3334);
nor U3626 (N_3626,N_2448,N_3400);
and U3627 (N_3627,N_2845,N_2470);
and U3628 (N_3628,N_2806,N_2465);
and U3629 (N_3629,N_2780,N_3013);
and U3630 (N_3630,N_2973,N_2606);
nand U3631 (N_3631,N_3526,N_2909);
nand U3632 (N_3632,N_2879,N_3204);
and U3633 (N_3633,N_2712,N_2983);
nand U3634 (N_3634,N_3495,N_2768);
and U3635 (N_3635,N_3413,N_3207);
and U3636 (N_3636,N_2820,N_2791);
nand U3637 (N_3637,N_3322,N_2664);
and U3638 (N_3638,N_3409,N_3587);
or U3639 (N_3639,N_2921,N_2497);
and U3640 (N_3640,N_3435,N_3419);
and U3641 (N_3641,N_2766,N_2917);
nand U3642 (N_3642,N_3378,N_2511);
or U3643 (N_3643,N_3191,N_2654);
xor U3644 (N_3644,N_2898,N_3249);
and U3645 (N_3645,N_3168,N_2503);
xor U3646 (N_3646,N_3482,N_2523);
and U3647 (N_3647,N_2897,N_2796);
nand U3648 (N_3648,N_3186,N_2657);
xor U3649 (N_3649,N_3499,N_2770);
nand U3650 (N_3650,N_3515,N_3053);
or U3651 (N_3651,N_2699,N_2522);
nand U3652 (N_3652,N_3462,N_3355);
or U3653 (N_3653,N_2784,N_2740);
nand U3654 (N_3654,N_2978,N_2982);
and U3655 (N_3655,N_3371,N_3434);
nor U3656 (N_3656,N_3197,N_3483);
nor U3657 (N_3657,N_2490,N_3098);
or U3658 (N_3658,N_3260,N_3465);
or U3659 (N_3659,N_2759,N_3180);
or U3660 (N_3660,N_2442,N_3147);
nor U3661 (N_3661,N_2422,N_3161);
or U3662 (N_3662,N_2414,N_3145);
nand U3663 (N_3663,N_2941,N_3002);
or U3664 (N_3664,N_2496,N_2985);
or U3665 (N_3665,N_3230,N_3095);
xor U3666 (N_3666,N_3310,N_3177);
and U3667 (N_3667,N_2587,N_3092);
or U3668 (N_3668,N_3384,N_2762);
and U3669 (N_3669,N_2635,N_2871);
or U3670 (N_3670,N_2416,N_2900);
or U3671 (N_3671,N_2781,N_2491);
nor U3672 (N_3672,N_3386,N_3134);
nor U3673 (N_3673,N_3152,N_2609);
or U3674 (N_3674,N_2541,N_3308);
and U3675 (N_3675,N_3398,N_2869);
xnor U3676 (N_3676,N_3235,N_3358);
and U3677 (N_3677,N_2914,N_2918);
nand U3678 (N_3678,N_2536,N_2854);
and U3679 (N_3679,N_2807,N_2643);
nand U3680 (N_3680,N_3001,N_2610);
nor U3681 (N_3681,N_2611,N_3121);
and U3682 (N_3682,N_3157,N_3130);
nand U3683 (N_3683,N_3243,N_2883);
nor U3684 (N_3684,N_3262,N_3397);
or U3685 (N_3685,N_3323,N_3074);
or U3686 (N_3686,N_2481,N_3052);
or U3687 (N_3687,N_3045,N_3108);
and U3688 (N_3688,N_3138,N_2627);
or U3689 (N_3689,N_3264,N_3458);
and U3690 (N_3690,N_3354,N_3569);
nor U3691 (N_3691,N_3151,N_2679);
xnor U3692 (N_3692,N_3490,N_3129);
and U3693 (N_3693,N_2744,N_2719);
xnor U3694 (N_3694,N_3122,N_3202);
nand U3695 (N_3695,N_2561,N_3278);
and U3696 (N_3696,N_3477,N_2437);
nor U3697 (N_3697,N_2860,N_2691);
xor U3698 (N_3698,N_2721,N_3060);
xnor U3699 (N_3699,N_2817,N_2865);
or U3700 (N_3700,N_3443,N_2552);
nor U3701 (N_3701,N_3366,N_2655);
nor U3702 (N_3702,N_3252,N_2452);
and U3703 (N_3703,N_2802,N_3271);
and U3704 (N_3704,N_3194,N_2954);
xor U3705 (N_3705,N_2583,N_3519);
and U3706 (N_3706,N_2575,N_3256);
and U3707 (N_3707,N_3274,N_2778);
or U3708 (N_3708,N_3543,N_2932);
nand U3709 (N_3709,N_2929,N_2737);
or U3710 (N_3710,N_3268,N_2892);
nand U3711 (N_3711,N_3455,N_2736);
nor U3712 (N_3712,N_3055,N_2881);
or U3713 (N_3713,N_2410,N_3297);
nor U3714 (N_3714,N_2834,N_3033);
nor U3715 (N_3715,N_2632,N_2872);
and U3716 (N_3716,N_2605,N_3336);
xnor U3717 (N_3717,N_2813,N_2733);
nor U3718 (N_3718,N_2567,N_2707);
xor U3719 (N_3719,N_2928,N_2829);
or U3720 (N_3720,N_2585,N_2818);
and U3721 (N_3721,N_3373,N_3275);
nor U3722 (N_3722,N_2880,N_2863);
xor U3723 (N_3723,N_2446,N_3300);
nor U3724 (N_3724,N_3144,N_3041);
and U3725 (N_3725,N_3286,N_3281);
xor U3726 (N_3726,N_3380,N_2594);
or U3727 (N_3727,N_3290,N_2580);
xnor U3728 (N_3728,N_3171,N_3215);
or U3729 (N_3729,N_3481,N_2758);
and U3730 (N_3730,N_3212,N_3005);
and U3731 (N_3731,N_3029,N_2571);
xnor U3732 (N_3732,N_2935,N_2968);
nor U3733 (N_3733,N_3575,N_2714);
nor U3734 (N_3734,N_2506,N_2940);
nor U3735 (N_3735,N_2560,N_2559);
or U3736 (N_3736,N_3225,N_3228);
nand U3737 (N_3737,N_2663,N_2920);
and U3738 (N_3738,N_3198,N_2592);
nand U3739 (N_3739,N_2652,N_2556);
and U3740 (N_3740,N_3209,N_2462);
nor U3741 (N_3741,N_3285,N_2593);
nand U3742 (N_3742,N_3589,N_2577);
nor U3743 (N_3743,N_3367,N_3201);
xor U3744 (N_3744,N_3222,N_2785);
nand U3745 (N_3745,N_2772,N_2459);
and U3746 (N_3746,N_2513,N_2810);
nand U3747 (N_3747,N_2519,N_3474);
or U3748 (N_3748,N_2822,N_2775);
or U3749 (N_3749,N_2574,N_2599);
and U3750 (N_3750,N_3597,N_3174);
and U3751 (N_3751,N_3530,N_2678);
nor U3752 (N_3752,N_2458,N_2521);
nand U3753 (N_3753,N_2788,N_2615);
nor U3754 (N_3754,N_2938,N_3067);
nand U3755 (N_3755,N_2415,N_3303);
nor U3756 (N_3756,N_3100,N_2626);
or U3757 (N_3757,N_3580,N_2461);
nor U3758 (N_3758,N_2750,N_3036);
nor U3759 (N_3759,N_3541,N_3287);
and U3760 (N_3760,N_3472,N_2717);
nor U3761 (N_3761,N_2407,N_2455);
and U3762 (N_3762,N_2538,N_3189);
or U3763 (N_3763,N_2525,N_3135);
nor U3764 (N_3764,N_3500,N_3115);
or U3765 (N_3765,N_3184,N_3595);
nand U3766 (N_3766,N_3072,N_3313);
or U3767 (N_3767,N_2600,N_2760);
or U3768 (N_3768,N_3497,N_3105);
or U3769 (N_3769,N_3231,N_2518);
or U3770 (N_3770,N_3328,N_2682);
nor U3771 (N_3771,N_3248,N_2651);
and U3772 (N_3772,N_2753,N_2468);
and U3773 (N_3773,N_3208,N_2554);
or U3774 (N_3774,N_2527,N_3229);
nor U3775 (N_3775,N_3090,N_3009);
and U3776 (N_3776,N_3216,N_2984);
xor U3777 (N_3777,N_3169,N_2642);
or U3778 (N_3778,N_3450,N_2509);
and U3779 (N_3779,N_2769,N_2505);
nand U3780 (N_3780,N_2549,N_3059);
xor U3781 (N_3781,N_3533,N_3487);
nand U3782 (N_3782,N_2915,N_3578);
xor U3783 (N_3783,N_2662,N_3254);
xnor U3784 (N_3784,N_3096,N_3512);
or U3785 (N_3785,N_2586,N_2588);
xor U3786 (N_3786,N_3081,N_2836);
or U3787 (N_3787,N_3181,N_3289);
xnor U3788 (N_3788,N_3280,N_2680);
xor U3789 (N_3789,N_2478,N_2958);
and U3790 (N_3790,N_2835,N_2887);
and U3791 (N_3791,N_2540,N_3051);
nand U3792 (N_3792,N_2956,N_2765);
nor U3793 (N_3793,N_2489,N_3047);
and U3794 (N_3794,N_2756,N_2483);
or U3795 (N_3795,N_3405,N_3025);
nand U3796 (N_3796,N_2856,N_2884);
nand U3797 (N_3797,N_2450,N_2716);
or U3798 (N_3798,N_2440,N_3399);
xor U3799 (N_3799,N_3118,N_3247);
and U3800 (N_3800,N_3043,N_3391);
nand U3801 (N_3801,N_2454,N_3031);
or U3802 (N_3802,N_3457,N_3241);
or U3803 (N_3803,N_3104,N_2516);
nand U3804 (N_3804,N_2779,N_3596);
xor U3805 (N_3805,N_2946,N_3517);
nand U3806 (N_3806,N_3542,N_2754);
and U3807 (N_3807,N_3035,N_3227);
and U3808 (N_3808,N_2919,N_2911);
or U3809 (N_3809,N_2631,N_2908);
xor U3810 (N_3810,N_3292,N_3192);
and U3811 (N_3811,N_3319,N_2755);
or U3812 (N_3812,N_2853,N_3393);
xnor U3813 (N_3813,N_3574,N_3195);
xor U3814 (N_3814,N_3453,N_3236);
xor U3815 (N_3815,N_3266,N_2428);
xnor U3816 (N_3816,N_2443,N_2517);
xnor U3817 (N_3817,N_3350,N_2659);
and U3818 (N_3818,N_3305,N_2622);
or U3819 (N_3819,N_2463,N_3492);
nor U3820 (N_3820,N_3535,N_2423);
nand U3821 (N_3821,N_3217,N_2992);
and U3822 (N_3822,N_2930,N_2833);
xor U3823 (N_3823,N_3459,N_2972);
and U3824 (N_3824,N_3594,N_3353);
and U3825 (N_3825,N_3529,N_2949);
and U3826 (N_3826,N_3253,N_3321);
nor U3827 (N_3827,N_3514,N_3348);
nor U3828 (N_3828,N_2823,N_3479);
xor U3829 (N_3829,N_2479,N_3581);
xor U3830 (N_3830,N_2814,N_3437);
nand U3831 (N_3831,N_2832,N_3511);
xor U3832 (N_3832,N_2412,N_2805);
and U3833 (N_3833,N_3226,N_2665);
or U3834 (N_3834,N_2683,N_2494);
or U3835 (N_3835,N_3200,N_3117);
xnor U3836 (N_3836,N_3507,N_3579);
or U3837 (N_3837,N_3068,N_2725);
nand U3838 (N_3838,N_3344,N_3557);
xor U3839 (N_3839,N_3556,N_3263);
nand U3840 (N_3840,N_2706,N_2916);
or U3841 (N_3841,N_2885,N_2730);
nor U3842 (N_3842,N_2891,N_2617);
xnor U3843 (N_3843,N_2743,N_2537);
xnor U3844 (N_3844,N_2507,N_3383);
or U3845 (N_3845,N_2994,N_2927);
xnor U3846 (N_3846,N_2550,N_2539);
nand U3847 (N_3847,N_3346,N_3475);
xnor U3848 (N_3848,N_3456,N_3000);
xor U3849 (N_3849,N_3233,N_2787);
or U3850 (N_3850,N_2488,N_2542);
xor U3851 (N_3851,N_2961,N_2432);
nor U3852 (N_3852,N_3258,N_2722);
and U3853 (N_3853,N_3162,N_3561);
xor U3854 (N_3854,N_2894,N_2738);
nor U3855 (N_3855,N_3298,N_2852);
nor U3856 (N_3856,N_2444,N_3585);
nor U3857 (N_3857,N_3411,N_3078);
and U3858 (N_3858,N_3214,N_2576);
or U3859 (N_3859,N_3006,N_2597);
nand U3860 (N_3860,N_3357,N_3342);
or U3861 (N_3861,N_3082,N_2646);
xor U3862 (N_3862,N_2512,N_3014);
xnor U3863 (N_3863,N_3071,N_2612);
or U3864 (N_3864,N_2767,N_3113);
nand U3865 (N_3865,N_3562,N_3326);
xor U3866 (N_3866,N_2942,N_3167);
xor U3867 (N_3867,N_2798,N_3038);
nand U3868 (N_3868,N_2735,N_3304);
nor U3869 (N_3869,N_2809,N_2742);
nand U3870 (N_3870,N_3431,N_3565);
and U3871 (N_3871,N_3220,N_2906);
nor U3872 (N_3872,N_3364,N_3550);
nand U3873 (N_3873,N_3091,N_3560);
xor U3874 (N_3874,N_3592,N_3028);
or U3875 (N_3875,N_3424,N_2715);
nand U3876 (N_3876,N_3288,N_2837);
xor U3877 (N_3877,N_2970,N_2988);
and U3878 (N_3878,N_2649,N_2669);
and U3879 (N_3879,N_2851,N_2907);
nor U3880 (N_3880,N_3279,N_2528);
and U3881 (N_3881,N_3396,N_2508);
xor U3882 (N_3882,N_2966,N_3295);
and U3883 (N_3883,N_2710,N_3410);
and U3884 (N_3884,N_2456,N_3064);
and U3885 (N_3885,N_3566,N_3505);
xor U3886 (N_3886,N_2697,N_2620);
and U3887 (N_3887,N_2672,N_3020);
xnor U3888 (N_3888,N_3257,N_3586);
nand U3889 (N_3889,N_3250,N_3017);
and U3890 (N_3890,N_3427,N_2830);
xnor U3891 (N_3891,N_2411,N_3375);
and U3892 (N_3892,N_3244,N_3193);
nor U3893 (N_3893,N_3402,N_2677);
or U3894 (N_3894,N_2558,N_3065);
or U3895 (N_3895,N_2792,N_3125);
xor U3896 (N_3896,N_3486,N_3494);
xnor U3897 (N_3897,N_3080,N_2439);
nor U3898 (N_3898,N_3470,N_2573);
nor U3899 (N_3899,N_2431,N_2532);
nor U3900 (N_3900,N_3044,N_3547);
or U3901 (N_3901,N_3401,N_2993);
xor U3902 (N_3902,N_2990,N_2445);
nor U3903 (N_3903,N_2749,N_2406);
nand U3904 (N_3904,N_3154,N_2967);
xnor U3905 (N_3905,N_2704,N_3160);
and U3906 (N_3906,N_3361,N_3493);
or U3907 (N_3907,N_3141,N_2524);
nor U3908 (N_3908,N_2498,N_2531);
or U3909 (N_3909,N_3442,N_2645);
and U3910 (N_3910,N_3513,N_3032);
xnor U3911 (N_3911,N_2739,N_2696);
xnor U3912 (N_3912,N_3420,N_2713);
and U3913 (N_3913,N_3387,N_3270);
and U3914 (N_3914,N_2801,N_3294);
and U3915 (N_3915,N_3418,N_3504);
nand U3916 (N_3916,N_3498,N_2675);
nor U3917 (N_3917,N_2864,N_2838);
or U3918 (N_3918,N_2763,N_2861);
and U3919 (N_3919,N_2614,N_3407);
or U3920 (N_3920,N_3251,N_3452);
xor U3921 (N_3921,N_2402,N_2584);
nand U3922 (N_3922,N_3054,N_3449);
and U3923 (N_3923,N_3073,N_3164);
nor U3924 (N_3924,N_3107,N_2684);
and U3925 (N_3925,N_3272,N_2421);
xnor U3926 (N_3926,N_3485,N_3057);
or U3927 (N_3927,N_3027,N_2761);
and U3928 (N_3928,N_2500,N_3445);
nor U3929 (N_3929,N_2473,N_2628);
or U3930 (N_3930,N_2757,N_2482);
xor U3931 (N_3931,N_3299,N_3234);
xnor U3932 (N_3932,N_3008,N_3538);
xnor U3933 (N_3933,N_3165,N_2815);
xor U3934 (N_3934,N_2430,N_3050);
and U3935 (N_3935,N_2579,N_3218);
or U3936 (N_3936,N_2565,N_3245);
and U3937 (N_3937,N_3148,N_3219);
and U3938 (N_3938,N_3056,N_2874);
nor U3939 (N_3939,N_2734,N_2855);
or U3940 (N_3940,N_3018,N_2821);
and U3941 (N_3941,N_3163,N_2702);
and U3942 (N_3942,N_3085,N_3388);
and U3943 (N_3943,N_3558,N_3571);
xnor U3944 (N_3944,N_3362,N_2793);
or U3945 (N_3945,N_3451,N_3546);
nor U3946 (N_3946,N_2711,N_3079);
and U3947 (N_3947,N_2889,N_3316);
nor U3948 (N_3948,N_2487,N_3205);
and U3949 (N_3949,N_2979,N_3577);
and U3950 (N_3950,N_2841,N_3570);
nor U3951 (N_3951,N_2698,N_2466);
or U3952 (N_3952,N_2771,N_3438);
nor U3953 (N_3953,N_3484,N_3124);
xor U3954 (N_3954,N_3099,N_2746);
nor U3955 (N_3955,N_3101,N_2510);
nand U3956 (N_3956,N_3232,N_3211);
and U3957 (N_3957,N_2616,N_3150);
nand U3958 (N_3958,N_2533,N_3395);
nand U3959 (N_3959,N_2547,N_2526);
nand U3960 (N_3960,N_2441,N_3496);
nand U3961 (N_3961,N_2991,N_3433);
nor U3962 (N_3962,N_3554,N_3007);
xnor U3963 (N_3963,N_3394,N_2925);
and U3964 (N_3964,N_3267,N_2952);
nand U3965 (N_3965,N_2732,N_3448);
and U3966 (N_3966,N_2644,N_3491);
and U3967 (N_3967,N_2681,N_3341);
nor U3968 (N_3968,N_3352,N_2688);
xor U3969 (N_3969,N_2886,N_2986);
and U3970 (N_3970,N_2619,N_3070);
or U3971 (N_3971,N_3039,N_2882);
nand U3972 (N_3972,N_3440,N_2839);
nand U3973 (N_3973,N_2971,N_3374);
nor U3974 (N_3974,N_2557,N_3528);
xnor U3975 (N_3975,N_3119,N_2658);
nand U3976 (N_3976,N_3159,N_2453);
nor U3977 (N_3977,N_2640,N_3338);
or U3978 (N_3978,N_3414,N_3369);
or U3979 (N_3979,N_3133,N_3520);
nor U3980 (N_3980,N_2467,N_3042);
xor U3981 (N_3981,N_3093,N_3255);
nor U3982 (N_3982,N_2890,N_2727);
nor U3983 (N_3983,N_2703,N_3089);
or U3984 (N_3984,N_2495,N_2603);
or U3985 (N_3985,N_3203,N_2690);
nand U3986 (N_3986,N_3473,N_3333);
xnor U3987 (N_3987,N_3447,N_2996);
and U3988 (N_3988,N_2694,N_2634);
xor U3989 (N_3989,N_3502,N_3284);
or U3990 (N_3990,N_2569,N_3010);
nor U3991 (N_3991,N_2457,N_2903);
nor U3992 (N_3992,N_3325,N_2955);
nor U3993 (N_3993,N_3423,N_3015);
nand U3994 (N_3994,N_3016,N_3572);
nor U3995 (N_3995,N_3291,N_3559);
nand U3996 (N_3996,N_2435,N_3343);
nand U3997 (N_3997,N_2425,N_3408);
and U3998 (N_3998,N_2912,N_2553);
nor U3999 (N_3999,N_3406,N_3127);
nand U4000 (N_4000,N_2774,N_2484);
or U4001 (N_4001,N_3381,N_2502);
and U4002 (N_4002,N_3426,N_3172);
xor U4003 (N_4003,N_2695,N_2436);
or U4004 (N_4004,N_2623,N_3312);
nand U4005 (N_4005,N_3318,N_3175);
or U4006 (N_4006,N_2786,N_2893);
nor U4007 (N_4007,N_2876,N_2980);
xor U4008 (N_4008,N_2501,N_2486);
nor U4009 (N_4009,N_3432,N_2426);
or U4010 (N_4010,N_2723,N_3488);
nor U4011 (N_4011,N_2418,N_3086);
and U4012 (N_4012,N_2963,N_2551);
nor U4013 (N_4013,N_3185,N_2438);
nand U4014 (N_4014,N_3382,N_2962);
or U4015 (N_4015,N_2563,N_3436);
xor U4016 (N_4016,N_3311,N_2685);
nor U4017 (N_4017,N_3421,N_2578);
xor U4018 (N_4018,N_3293,N_3508);
or U4019 (N_4019,N_2514,N_3463);
or U4020 (N_4020,N_2824,N_3012);
nor U4021 (N_4021,N_2800,N_2811);
nor U4022 (N_4022,N_3324,N_2475);
and U4023 (N_4023,N_3004,N_3576);
or U4024 (N_4024,N_2731,N_3468);
and U4025 (N_4025,N_3040,N_2601);
nor U4026 (N_4026,N_3069,N_3536);
and U4027 (N_4027,N_3545,N_2472);
and U4028 (N_4028,N_3392,N_3276);
and U4029 (N_4029,N_2709,N_2844);
nand U4030 (N_4030,N_3188,N_2747);
nor U4031 (N_4031,N_2794,N_2764);
nand U4032 (N_4032,N_3331,N_2653);
nand U4033 (N_4033,N_3155,N_3469);
nor U4034 (N_4034,N_2751,N_2562);
or U4035 (N_4035,N_3471,N_2816);
nor U4036 (N_4036,N_2741,N_2773);
and U4037 (N_4037,N_2602,N_3501);
or U4038 (N_4038,N_2846,N_2724);
xor U4039 (N_4039,N_2943,N_2926);
xnor U4040 (N_4040,N_3525,N_3240);
and U4041 (N_4041,N_3094,N_3441);
nor U4042 (N_4042,N_2485,N_2803);
and U4043 (N_4043,N_3123,N_2999);
nor U4044 (N_4044,N_2812,N_2530);
or U4045 (N_4045,N_3555,N_2433);
and U4046 (N_4046,N_2981,N_3143);
xor U4047 (N_4047,N_3337,N_3548);
nand U4048 (N_4048,N_2904,N_2596);
or U4049 (N_4049,N_3061,N_3422);
nand U4050 (N_4050,N_2424,N_2647);
xor U4051 (N_4051,N_3510,N_2913);
and U4052 (N_4052,N_3339,N_2581);
nor U4053 (N_4053,N_2401,N_3179);
xnor U4054 (N_4054,N_3518,N_2888);
nor U4055 (N_4055,N_3126,N_3139);
and U4056 (N_4056,N_2671,N_2964);
and U4057 (N_4057,N_2923,N_2989);
nand U4058 (N_4058,N_2545,N_2804);
xnor U4059 (N_4059,N_3332,N_2933);
nand U4060 (N_4060,N_2667,N_2951);
xor U4061 (N_4061,N_2413,N_3593);
and U4062 (N_4062,N_2868,N_2409);
and U4063 (N_4063,N_3019,N_2570);
xor U4064 (N_4064,N_3532,N_3461);
or U4065 (N_4065,N_3446,N_2848);
nand U4066 (N_4066,N_2790,N_3349);
or U4067 (N_4067,N_3048,N_3142);
xor U4068 (N_4068,N_2776,N_2789);
and U4069 (N_4069,N_3590,N_2661);
or U4070 (N_4070,N_2902,N_3109);
and U4071 (N_4071,N_3178,N_2720);
or U4072 (N_4072,N_2826,N_3183);
xor U4073 (N_4073,N_3307,N_3182);
xor U4074 (N_4074,N_3460,N_2564);
or U4075 (N_4075,N_2451,N_3478);
and U4076 (N_4076,N_3390,N_2499);
or U4077 (N_4077,N_2858,N_3114);
nand U4078 (N_4078,N_2625,N_2666);
nand U4079 (N_4079,N_3330,N_3302);
xor U4080 (N_4080,N_2896,N_3136);
xnor U4081 (N_4081,N_3306,N_2534);
or U4082 (N_4082,N_2400,N_3140);
nand U4083 (N_4083,N_3282,N_3320);
xor U4084 (N_4084,N_3075,N_2828);
nor U4085 (N_4085,N_3037,N_3584);
nor U4086 (N_4086,N_2589,N_3046);
nand U4087 (N_4087,N_3261,N_2866);
nor U4088 (N_4088,N_3564,N_2937);
nand U4089 (N_4089,N_3102,N_3062);
or U4090 (N_4090,N_2639,N_3372);
and U4091 (N_4091,N_2660,N_3403);
or U4092 (N_4092,N_2492,N_3368);
nor U4093 (N_4093,N_3199,N_2608);
nor U4094 (N_4094,N_3552,N_2877);
and U4095 (N_4095,N_3503,N_3187);
nand U4096 (N_4096,N_3158,N_2604);
or U4097 (N_4097,N_2777,N_3301);
and U4098 (N_4098,N_3190,N_3076);
nor U4099 (N_4099,N_2975,N_2613);
nor U4100 (N_4100,N_3223,N_2630);
or U4101 (N_4101,N_2948,N_2520);
xor U4102 (N_4102,N_3022,N_2515);
nor U4103 (N_4103,N_3239,N_3176);
and U4104 (N_4104,N_2449,N_2429);
and U4105 (N_4105,N_2899,N_3077);
and U4106 (N_4106,N_3476,N_3429);
nand U4107 (N_4107,N_3549,N_3146);
nor U4108 (N_4108,N_2987,N_2504);
or U4109 (N_4109,N_3379,N_2529);
xnor U4110 (N_4110,N_2618,N_2795);
and U4111 (N_4111,N_3112,N_2718);
nand U4112 (N_4112,N_2477,N_2650);
xor U4113 (N_4113,N_3132,N_2638);
or U4114 (N_4114,N_3120,N_3021);
nand U4115 (N_4115,N_3340,N_2701);
nand U4116 (N_4116,N_2748,N_3522);
nand U4117 (N_4117,N_3359,N_3030);
and U4118 (N_4118,N_3296,N_3527);
nor U4119 (N_4119,N_2953,N_2700);
xnor U4120 (N_4120,N_3377,N_2959);
xor U4121 (N_4121,N_3356,N_2555);
nand U4122 (N_4122,N_2745,N_2808);
and U4123 (N_4123,N_3454,N_3540);
or U4124 (N_4124,N_2847,N_3087);
and U4125 (N_4125,N_3314,N_2729);
and U4126 (N_4126,N_3259,N_2910);
xor U4127 (N_4127,N_3523,N_3131);
nand U4128 (N_4128,N_2950,N_3265);
or U4129 (N_4129,N_2598,N_3531);
nand U4130 (N_4130,N_2572,N_3137);
nor U4131 (N_4131,N_2873,N_3238);
and U4132 (N_4132,N_2936,N_2656);
xnor U4133 (N_4133,N_3416,N_3524);
or U4134 (N_4134,N_2641,N_2434);
xor U4135 (N_4135,N_3327,N_3598);
xor U4136 (N_4136,N_3173,N_3011);
nand U4137 (N_4137,N_3221,N_3153);
or U4138 (N_4138,N_3149,N_2408);
or U4139 (N_4139,N_2977,N_3365);
nor U4140 (N_4140,N_3003,N_3277);
or U4141 (N_4141,N_2668,N_3425);
and U4142 (N_4142,N_2419,N_3206);
nand U4143 (N_4143,N_2493,N_3363);
or U4144 (N_4144,N_2637,N_2417);
nor U4145 (N_4145,N_3467,N_3023);
or U4146 (N_4146,N_3026,N_3315);
nor U4147 (N_4147,N_2905,N_3084);
and U4148 (N_4148,N_3024,N_2464);
nand U4149 (N_4149,N_3335,N_3273);
nor U4150 (N_4150,N_3583,N_3567);
nor U4151 (N_4151,N_2607,N_3539);
and U4152 (N_4152,N_3544,N_2957);
nor U4153 (N_4153,N_3329,N_2686);
nand U4154 (N_4154,N_3568,N_2997);
nand U4155 (N_4155,N_2591,N_3404);
nand U4156 (N_4156,N_2674,N_2922);
xnor U4157 (N_4157,N_2689,N_2831);
and U4158 (N_4158,N_2998,N_2783);
nor U4159 (N_4159,N_3417,N_2843);
xor U4160 (N_4160,N_2566,N_2752);
and U4161 (N_4161,N_3599,N_3360);
and U4162 (N_4162,N_2965,N_2708);
nand U4163 (N_4163,N_2480,N_3466);
nor U4164 (N_4164,N_2595,N_2693);
xor U4165 (N_4165,N_3063,N_3444);
or U4166 (N_4166,N_3464,N_3376);
and U4167 (N_4167,N_3034,N_2976);
nor U4168 (N_4168,N_2842,N_2934);
nor U4169 (N_4169,N_3534,N_2825);
and U4170 (N_4170,N_2895,N_3166);
nor U4171 (N_4171,N_3196,N_2827);
or U4172 (N_4172,N_2859,N_3428);
nor U4173 (N_4173,N_2939,N_2544);
xor U4174 (N_4174,N_2728,N_3283);
and U4175 (N_4175,N_3370,N_2862);
or U4176 (N_4176,N_3430,N_2636);
nand U4177 (N_4177,N_2726,N_2857);
and U4178 (N_4178,N_3588,N_2474);
and U4179 (N_4179,N_3591,N_3389);
xnor U4180 (N_4180,N_3111,N_2850);
and U4181 (N_4181,N_2878,N_2621);
xor U4182 (N_4182,N_3246,N_3049);
xor U4183 (N_4183,N_2947,N_3170);
nand U4184 (N_4184,N_2469,N_3224);
and U4185 (N_4185,N_3415,N_3506);
nor U4186 (N_4186,N_3242,N_3106);
xnor U4187 (N_4187,N_3439,N_2535);
and U4188 (N_4188,N_2799,N_2460);
or U4189 (N_4189,N_2692,N_3156);
and U4190 (N_4190,N_2944,N_2582);
nor U4191 (N_4191,N_3509,N_2568);
or U4192 (N_4192,N_3128,N_2687);
or U4193 (N_4193,N_2548,N_2648);
or U4194 (N_4194,N_2624,N_3351);
and U4195 (N_4195,N_3551,N_2960);
xor U4196 (N_4196,N_3269,N_3537);
and U4197 (N_4197,N_2782,N_2633);
nor U4198 (N_4198,N_3563,N_3058);
xnor U4199 (N_4199,N_2546,N_3116);
and U4200 (N_4200,N_2726,N_3576);
nand U4201 (N_4201,N_3404,N_2754);
and U4202 (N_4202,N_2679,N_2768);
and U4203 (N_4203,N_2902,N_3465);
or U4204 (N_4204,N_3437,N_3344);
and U4205 (N_4205,N_2480,N_3418);
and U4206 (N_4206,N_2990,N_3391);
nor U4207 (N_4207,N_2701,N_3530);
xnor U4208 (N_4208,N_3539,N_2426);
and U4209 (N_4209,N_2656,N_2911);
xnor U4210 (N_4210,N_3019,N_2611);
and U4211 (N_4211,N_2906,N_3474);
or U4212 (N_4212,N_3087,N_3199);
and U4213 (N_4213,N_2549,N_2759);
xnor U4214 (N_4214,N_3587,N_3316);
and U4215 (N_4215,N_3131,N_3293);
nor U4216 (N_4216,N_2796,N_2710);
xor U4217 (N_4217,N_3284,N_2512);
xnor U4218 (N_4218,N_2747,N_3126);
nor U4219 (N_4219,N_2444,N_3306);
nand U4220 (N_4220,N_2628,N_3350);
or U4221 (N_4221,N_2811,N_3376);
nand U4222 (N_4222,N_3026,N_2429);
nor U4223 (N_4223,N_2837,N_2792);
and U4224 (N_4224,N_3113,N_2495);
xnor U4225 (N_4225,N_2884,N_3520);
nor U4226 (N_4226,N_2639,N_3172);
nand U4227 (N_4227,N_3340,N_3548);
nand U4228 (N_4228,N_3395,N_3028);
xnor U4229 (N_4229,N_3584,N_2509);
nor U4230 (N_4230,N_2666,N_2605);
nand U4231 (N_4231,N_2918,N_2514);
nand U4232 (N_4232,N_2643,N_3560);
nor U4233 (N_4233,N_3457,N_2920);
nand U4234 (N_4234,N_2838,N_3098);
nand U4235 (N_4235,N_2570,N_2700);
or U4236 (N_4236,N_3233,N_3065);
or U4237 (N_4237,N_2601,N_2984);
nor U4238 (N_4238,N_3435,N_3362);
nor U4239 (N_4239,N_2698,N_2927);
nor U4240 (N_4240,N_3087,N_2591);
and U4241 (N_4241,N_3472,N_2522);
nand U4242 (N_4242,N_3056,N_2902);
nor U4243 (N_4243,N_3121,N_2612);
and U4244 (N_4244,N_3418,N_2550);
xnor U4245 (N_4245,N_2775,N_2584);
xor U4246 (N_4246,N_3457,N_2626);
or U4247 (N_4247,N_3087,N_3503);
nor U4248 (N_4248,N_2860,N_3228);
and U4249 (N_4249,N_3085,N_2831);
nor U4250 (N_4250,N_2863,N_3471);
or U4251 (N_4251,N_3483,N_3166);
nand U4252 (N_4252,N_3320,N_3081);
xor U4253 (N_4253,N_2538,N_3351);
nor U4254 (N_4254,N_2550,N_2548);
nand U4255 (N_4255,N_2958,N_3489);
and U4256 (N_4256,N_2656,N_2447);
nor U4257 (N_4257,N_3241,N_3587);
and U4258 (N_4258,N_3259,N_2450);
or U4259 (N_4259,N_2447,N_3441);
xnor U4260 (N_4260,N_2937,N_2532);
xnor U4261 (N_4261,N_3175,N_3325);
nand U4262 (N_4262,N_2781,N_2494);
and U4263 (N_4263,N_3356,N_3384);
or U4264 (N_4264,N_2890,N_2579);
xor U4265 (N_4265,N_2695,N_3053);
nand U4266 (N_4266,N_2469,N_3513);
nor U4267 (N_4267,N_3052,N_3483);
or U4268 (N_4268,N_3366,N_3241);
xor U4269 (N_4269,N_2882,N_3319);
and U4270 (N_4270,N_3374,N_3357);
xor U4271 (N_4271,N_3591,N_2432);
or U4272 (N_4272,N_3429,N_3125);
or U4273 (N_4273,N_3187,N_3571);
xnor U4274 (N_4274,N_3099,N_2731);
or U4275 (N_4275,N_2624,N_2946);
xor U4276 (N_4276,N_3525,N_3201);
nand U4277 (N_4277,N_2921,N_2772);
nand U4278 (N_4278,N_3515,N_3194);
nor U4279 (N_4279,N_3046,N_2497);
nor U4280 (N_4280,N_3213,N_2559);
nand U4281 (N_4281,N_3586,N_3438);
nand U4282 (N_4282,N_3234,N_3048);
xnor U4283 (N_4283,N_2881,N_2902);
nor U4284 (N_4284,N_2607,N_2405);
xor U4285 (N_4285,N_3129,N_2558);
and U4286 (N_4286,N_3136,N_3445);
nor U4287 (N_4287,N_3250,N_2818);
and U4288 (N_4288,N_2828,N_3524);
nor U4289 (N_4289,N_2911,N_2802);
and U4290 (N_4290,N_3094,N_2933);
nand U4291 (N_4291,N_2889,N_3116);
nor U4292 (N_4292,N_3577,N_3038);
or U4293 (N_4293,N_2451,N_2818);
and U4294 (N_4294,N_3476,N_3144);
nor U4295 (N_4295,N_3237,N_3567);
or U4296 (N_4296,N_2808,N_2967);
nand U4297 (N_4297,N_2609,N_2903);
xor U4298 (N_4298,N_2505,N_2706);
nand U4299 (N_4299,N_2709,N_3073);
and U4300 (N_4300,N_3322,N_2723);
or U4301 (N_4301,N_2730,N_2876);
and U4302 (N_4302,N_2532,N_2444);
or U4303 (N_4303,N_3331,N_2414);
or U4304 (N_4304,N_2469,N_3165);
nand U4305 (N_4305,N_3015,N_3065);
nand U4306 (N_4306,N_3283,N_3032);
and U4307 (N_4307,N_3124,N_2795);
or U4308 (N_4308,N_2724,N_3482);
or U4309 (N_4309,N_3429,N_3144);
and U4310 (N_4310,N_3069,N_3293);
or U4311 (N_4311,N_3222,N_3440);
nor U4312 (N_4312,N_3553,N_2457);
nor U4313 (N_4313,N_2600,N_3461);
nand U4314 (N_4314,N_2700,N_3212);
xor U4315 (N_4315,N_2687,N_2600);
or U4316 (N_4316,N_2673,N_3483);
or U4317 (N_4317,N_3016,N_2496);
xnor U4318 (N_4318,N_2639,N_3388);
nor U4319 (N_4319,N_2594,N_2482);
and U4320 (N_4320,N_3540,N_2528);
nor U4321 (N_4321,N_3111,N_3220);
xor U4322 (N_4322,N_2715,N_2889);
or U4323 (N_4323,N_3192,N_2955);
nor U4324 (N_4324,N_2510,N_2944);
or U4325 (N_4325,N_3569,N_2933);
nor U4326 (N_4326,N_2543,N_3142);
xnor U4327 (N_4327,N_3246,N_2680);
nand U4328 (N_4328,N_3008,N_2621);
nor U4329 (N_4329,N_2877,N_2482);
and U4330 (N_4330,N_2548,N_3226);
nor U4331 (N_4331,N_3102,N_2536);
or U4332 (N_4332,N_2928,N_3211);
nand U4333 (N_4333,N_3429,N_3087);
nor U4334 (N_4334,N_3465,N_3356);
or U4335 (N_4335,N_2901,N_3548);
and U4336 (N_4336,N_3043,N_3558);
and U4337 (N_4337,N_2958,N_3501);
xor U4338 (N_4338,N_2790,N_3580);
or U4339 (N_4339,N_2769,N_2608);
and U4340 (N_4340,N_2594,N_3537);
nand U4341 (N_4341,N_2900,N_3521);
xnor U4342 (N_4342,N_2497,N_2931);
or U4343 (N_4343,N_3063,N_3226);
and U4344 (N_4344,N_3064,N_2935);
or U4345 (N_4345,N_2704,N_3086);
nand U4346 (N_4346,N_3130,N_3321);
nand U4347 (N_4347,N_2501,N_2876);
and U4348 (N_4348,N_3251,N_2857);
and U4349 (N_4349,N_3510,N_2695);
nand U4350 (N_4350,N_2409,N_3598);
or U4351 (N_4351,N_3458,N_3188);
xor U4352 (N_4352,N_3580,N_2805);
and U4353 (N_4353,N_2821,N_2747);
or U4354 (N_4354,N_3489,N_3569);
nor U4355 (N_4355,N_3133,N_3266);
xor U4356 (N_4356,N_2429,N_3556);
or U4357 (N_4357,N_3185,N_3260);
or U4358 (N_4358,N_2499,N_3334);
or U4359 (N_4359,N_2625,N_2504);
xor U4360 (N_4360,N_2984,N_3420);
nor U4361 (N_4361,N_2912,N_3077);
nor U4362 (N_4362,N_3051,N_2447);
nor U4363 (N_4363,N_3427,N_2857);
nor U4364 (N_4364,N_3069,N_2744);
nor U4365 (N_4365,N_3380,N_3143);
nor U4366 (N_4366,N_3481,N_2680);
xnor U4367 (N_4367,N_2979,N_3363);
nor U4368 (N_4368,N_3022,N_3218);
and U4369 (N_4369,N_2496,N_3088);
nor U4370 (N_4370,N_2586,N_2536);
nand U4371 (N_4371,N_2467,N_2786);
or U4372 (N_4372,N_2686,N_2457);
or U4373 (N_4373,N_2973,N_2827);
nor U4374 (N_4374,N_2964,N_3451);
or U4375 (N_4375,N_2879,N_3463);
xor U4376 (N_4376,N_2855,N_3164);
or U4377 (N_4377,N_2810,N_2837);
or U4378 (N_4378,N_3221,N_3396);
nor U4379 (N_4379,N_3372,N_2666);
xor U4380 (N_4380,N_3115,N_3035);
xnor U4381 (N_4381,N_3485,N_2511);
and U4382 (N_4382,N_3430,N_3192);
nand U4383 (N_4383,N_2461,N_2420);
or U4384 (N_4384,N_2811,N_2738);
xnor U4385 (N_4385,N_3390,N_2946);
nand U4386 (N_4386,N_3062,N_2439);
nand U4387 (N_4387,N_2499,N_2697);
or U4388 (N_4388,N_2973,N_2680);
xnor U4389 (N_4389,N_3355,N_3134);
or U4390 (N_4390,N_2603,N_3490);
xor U4391 (N_4391,N_2578,N_2547);
nor U4392 (N_4392,N_3142,N_3417);
xnor U4393 (N_4393,N_3473,N_3061);
and U4394 (N_4394,N_2776,N_2926);
nand U4395 (N_4395,N_2980,N_3443);
and U4396 (N_4396,N_3202,N_2533);
xnor U4397 (N_4397,N_3167,N_3004);
and U4398 (N_4398,N_3268,N_2618);
nor U4399 (N_4399,N_3571,N_3347);
nand U4400 (N_4400,N_2816,N_3022);
or U4401 (N_4401,N_2577,N_2502);
nor U4402 (N_4402,N_3362,N_3132);
xor U4403 (N_4403,N_3271,N_2471);
nor U4404 (N_4404,N_3497,N_2405);
xor U4405 (N_4405,N_2428,N_3588);
and U4406 (N_4406,N_3409,N_3348);
xor U4407 (N_4407,N_3106,N_3158);
nand U4408 (N_4408,N_3057,N_3569);
and U4409 (N_4409,N_2584,N_2520);
or U4410 (N_4410,N_2768,N_2968);
nor U4411 (N_4411,N_3192,N_2557);
nor U4412 (N_4412,N_3013,N_2430);
nor U4413 (N_4413,N_3089,N_3042);
or U4414 (N_4414,N_3006,N_2416);
and U4415 (N_4415,N_2416,N_3218);
xor U4416 (N_4416,N_2672,N_2576);
nand U4417 (N_4417,N_2796,N_3333);
nor U4418 (N_4418,N_3205,N_2401);
xor U4419 (N_4419,N_2624,N_2676);
nor U4420 (N_4420,N_2671,N_2887);
or U4421 (N_4421,N_3157,N_3021);
and U4422 (N_4422,N_2989,N_3156);
or U4423 (N_4423,N_3002,N_3038);
xnor U4424 (N_4424,N_3367,N_3235);
nand U4425 (N_4425,N_2584,N_2544);
nand U4426 (N_4426,N_3248,N_2953);
nor U4427 (N_4427,N_3417,N_3130);
or U4428 (N_4428,N_2980,N_3341);
nand U4429 (N_4429,N_3216,N_3157);
xor U4430 (N_4430,N_3542,N_2412);
xnor U4431 (N_4431,N_3424,N_2831);
nor U4432 (N_4432,N_3002,N_3335);
nor U4433 (N_4433,N_2609,N_3310);
nor U4434 (N_4434,N_2887,N_3385);
nand U4435 (N_4435,N_3563,N_3312);
or U4436 (N_4436,N_3383,N_2907);
or U4437 (N_4437,N_2804,N_3376);
nand U4438 (N_4438,N_3539,N_3299);
or U4439 (N_4439,N_2879,N_2841);
and U4440 (N_4440,N_2562,N_2714);
or U4441 (N_4441,N_2461,N_3505);
nor U4442 (N_4442,N_3258,N_2968);
xor U4443 (N_4443,N_3474,N_3552);
nand U4444 (N_4444,N_2916,N_3572);
and U4445 (N_4445,N_3393,N_3490);
nor U4446 (N_4446,N_2778,N_3025);
xor U4447 (N_4447,N_2784,N_2752);
and U4448 (N_4448,N_2743,N_3583);
and U4449 (N_4449,N_2727,N_2692);
nor U4450 (N_4450,N_3353,N_2651);
and U4451 (N_4451,N_3416,N_3254);
nand U4452 (N_4452,N_3098,N_3278);
nor U4453 (N_4453,N_3327,N_3147);
and U4454 (N_4454,N_3576,N_3595);
nand U4455 (N_4455,N_3258,N_2469);
xnor U4456 (N_4456,N_3248,N_2987);
nor U4457 (N_4457,N_3200,N_3517);
and U4458 (N_4458,N_3569,N_3096);
or U4459 (N_4459,N_3549,N_3567);
nand U4460 (N_4460,N_2999,N_2686);
nand U4461 (N_4461,N_3028,N_2548);
xor U4462 (N_4462,N_3087,N_2805);
xnor U4463 (N_4463,N_3114,N_3145);
or U4464 (N_4464,N_2852,N_3477);
or U4465 (N_4465,N_2435,N_2590);
and U4466 (N_4466,N_2448,N_2753);
nand U4467 (N_4467,N_2967,N_3417);
nor U4468 (N_4468,N_2569,N_2952);
xor U4469 (N_4469,N_3290,N_2996);
nand U4470 (N_4470,N_3146,N_3286);
nand U4471 (N_4471,N_2850,N_2634);
xor U4472 (N_4472,N_3338,N_3420);
xor U4473 (N_4473,N_2646,N_2525);
nand U4474 (N_4474,N_3079,N_2665);
nand U4475 (N_4475,N_3098,N_2731);
nand U4476 (N_4476,N_2460,N_3057);
or U4477 (N_4477,N_2531,N_3397);
or U4478 (N_4478,N_2993,N_2628);
nand U4479 (N_4479,N_3049,N_3302);
nor U4480 (N_4480,N_2845,N_2938);
nand U4481 (N_4481,N_2415,N_2797);
nand U4482 (N_4482,N_2944,N_3186);
nand U4483 (N_4483,N_3367,N_3477);
or U4484 (N_4484,N_2458,N_3491);
and U4485 (N_4485,N_2853,N_3066);
and U4486 (N_4486,N_3075,N_3489);
nand U4487 (N_4487,N_2586,N_3011);
xnor U4488 (N_4488,N_2689,N_2443);
nor U4489 (N_4489,N_3069,N_2746);
xnor U4490 (N_4490,N_3064,N_3527);
and U4491 (N_4491,N_3150,N_2767);
and U4492 (N_4492,N_3468,N_3336);
or U4493 (N_4493,N_2612,N_3305);
nor U4494 (N_4494,N_2792,N_2415);
or U4495 (N_4495,N_3492,N_2710);
nand U4496 (N_4496,N_3015,N_3374);
xor U4497 (N_4497,N_3415,N_3054);
or U4498 (N_4498,N_3017,N_3292);
nand U4499 (N_4499,N_2840,N_3414);
nand U4500 (N_4500,N_2434,N_3031);
and U4501 (N_4501,N_3250,N_3151);
and U4502 (N_4502,N_2671,N_2569);
or U4503 (N_4503,N_3590,N_3128);
or U4504 (N_4504,N_2902,N_3237);
xor U4505 (N_4505,N_3107,N_3136);
xnor U4506 (N_4506,N_3555,N_3375);
xor U4507 (N_4507,N_2628,N_2757);
or U4508 (N_4508,N_3294,N_2545);
nand U4509 (N_4509,N_2814,N_2458);
and U4510 (N_4510,N_2935,N_3162);
nand U4511 (N_4511,N_3534,N_3498);
or U4512 (N_4512,N_3095,N_2589);
and U4513 (N_4513,N_2597,N_2485);
nor U4514 (N_4514,N_2979,N_2415);
and U4515 (N_4515,N_3312,N_2919);
and U4516 (N_4516,N_2640,N_3234);
xnor U4517 (N_4517,N_2467,N_3344);
xor U4518 (N_4518,N_2957,N_2984);
nand U4519 (N_4519,N_2651,N_2888);
xnor U4520 (N_4520,N_3383,N_3279);
nor U4521 (N_4521,N_2504,N_3419);
xnor U4522 (N_4522,N_2763,N_3436);
nand U4523 (N_4523,N_3598,N_2899);
nand U4524 (N_4524,N_3522,N_2653);
xor U4525 (N_4525,N_3163,N_2945);
xnor U4526 (N_4526,N_3274,N_2939);
xor U4527 (N_4527,N_2708,N_3152);
nor U4528 (N_4528,N_2998,N_3405);
nand U4529 (N_4529,N_3537,N_3270);
xor U4530 (N_4530,N_3521,N_2590);
and U4531 (N_4531,N_2822,N_3075);
nand U4532 (N_4532,N_3444,N_3453);
and U4533 (N_4533,N_2521,N_3496);
nor U4534 (N_4534,N_3561,N_3212);
and U4535 (N_4535,N_3495,N_2984);
xnor U4536 (N_4536,N_2690,N_3146);
or U4537 (N_4537,N_2629,N_2673);
nor U4538 (N_4538,N_2969,N_2462);
nand U4539 (N_4539,N_2896,N_3358);
and U4540 (N_4540,N_2504,N_3103);
nor U4541 (N_4541,N_3102,N_2791);
nand U4542 (N_4542,N_2875,N_2568);
xor U4543 (N_4543,N_3404,N_2750);
or U4544 (N_4544,N_3361,N_2857);
nand U4545 (N_4545,N_2994,N_2759);
and U4546 (N_4546,N_3350,N_3043);
nor U4547 (N_4547,N_2590,N_2799);
nand U4548 (N_4548,N_2598,N_2945);
nor U4549 (N_4549,N_2410,N_3301);
nand U4550 (N_4550,N_3126,N_2788);
xor U4551 (N_4551,N_3208,N_3365);
xor U4552 (N_4552,N_3425,N_3201);
nand U4553 (N_4553,N_3510,N_2582);
nor U4554 (N_4554,N_3578,N_3498);
xnor U4555 (N_4555,N_3003,N_3010);
nor U4556 (N_4556,N_3039,N_2773);
nand U4557 (N_4557,N_3429,N_3356);
nand U4558 (N_4558,N_2574,N_3345);
nand U4559 (N_4559,N_3530,N_3225);
xor U4560 (N_4560,N_2498,N_2916);
nor U4561 (N_4561,N_2654,N_2938);
nand U4562 (N_4562,N_3442,N_2418);
xor U4563 (N_4563,N_2793,N_3307);
xnor U4564 (N_4564,N_2615,N_3423);
nand U4565 (N_4565,N_2753,N_2972);
nor U4566 (N_4566,N_3449,N_3033);
nand U4567 (N_4567,N_2540,N_2402);
and U4568 (N_4568,N_2410,N_2503);
and U4569 (N_4569,N_2594,N_2891);
nor U4570 (N_4570,N_2827,N_3583);
or U4571 (N_4571,N_2976,N_2455);
nand U4572 (N_4572,N_2497,N_3352);
nand U4573 (N_4573,N_2493,N_3466);
nand U4574 (N_4574,N_3473,N_2946);
xor U4575 (N_4575,N_2578,N_3024);
xor U4576 (N_4576,N_3411,N_2711);
nor U4577 (N_4577,N_2954,N_2527);
and U4578 (N_4578,N_3398,N_3346);
nor U4579 (N_4579,N_2465,N_3504);
nand U4580 (N_4580,N_3322,N_3279);
nand U4581 (N_4581,N_3162,N_2597);
or U4582 (N_4582,N_3553,N_2423);
and U4583 (N_4583,N_2643,N_3179);
nand U4584 (N_4584,N_3558,N_3353);
nand U4585 (N_4585,N_3309,N_2908);
xor U4586 (N_4586,N_3012,N_2674);
xor U4587 (N_4587,N_3214,N_2640);
xor U4588 (N_4588,N_3104,N_3196);
or U4589 (N_4589,N_3421,N_2927);
or U4590 (N_4590,N_2436,N_2909);
xor U4591 (N_4591,N_2578,N_2425);
xor U4592 (N_4592,N_3556,N_2492);
and U4593 (N_4593,N_3367,N_3453);
nor U4594 (N_4594,N_3414,N_3335);
nand U4595 (N_4595,N_2534,N_2674);
and U4596 (N_4596,N_3451,N_3389);
and U4597 (N_4597,N_2743,N_3425);
nor U4598 (N_4598,N_3533,N_2593);
or U4599 (N_4599,N_3288,N_3392);
and U4600 (N_4600,N_2982,N_3013);
nor U4601 (N_4601,N_2430,N_2984);
nand U4602 (N_4602,N_2622,N_3395);
and U4603 (N_4603,N_2848,N_2746);
nand U4604 (N_4604,N_2680,N_3029);
nand U4605 (N_4605,N_3436,N_3463);
and U4606 (N_4606,N_2708,N_2719);
nand U4607 (N_4607,N_2464,N_2503);
nor U4608 (N_4608,N_3245,N_2889);
and U4609 (N_4609,N_2555,N_3056);
nand U4610 (N_4610,N_2447,N_3064);
xnor U4611 (N_4611,N_3182,N_3301);
nor U4612 (N_4612,N_2830,N_2587);
nand U4613 (N_4613,N_3469,N_2454);
xor U4614 (N_4614,N_3367,N_3220);
xnor U4615 (N_4615,N_2483,N_2976);
nor U4616 (N_4616,N_2494,N_2777);
nand U4617 (N_4617,N_3304,N_2943);
and U4618 (N_4618,N_2540,N_2623);
xor U4619 (N_4619,N_3577,N_2647);
and U4620 (N_4620,N_2874,N_3197);
xnor U4621 (N_4621,N_3029,N_3268);
nor U4622 (N_4622,N_2540,N_3130);
xnor U4623 (N_4623,N_3182,N_3534);
or U4624 (N_4624,N_2698,N_2539);
or U4625 (N_4625,N_2573,N_3017);
or U4626 (N_4626,N_3462,N_2765);
nand U4627 (N_4627,N_2526,N_2570);
or U4628 (N_4628,N_3140,N_3321);
xor U4629 (N_4629,N_3070,N_2609);
xor U4630 (N_4630,N_2603,N_3485);
xor U4631 (N_4631,N_3065,N_2729);
or U4632 (N_4632,N_2949,N_2538);
nor U4633 (N_4633,N_2676,N_2406);
or U4634 (N_4634,N_2513,N_2471);
nor U4635 (N_4635,N_2692,N_3193);
nand U4636 (N_4636,N_3431,N_2799);
nand U4637 (N_4637,N_2457,N_2533);
nor U4638 (N_4638,N_3188,N_3525);
and U4639 (N_4639,N_2829,N_3048);
nand U4640 (N_4640,N_3326,N_2486);
nand U4641 (N_4641,N_3119,N_3324);
xnor U4642 (N_4642,N_3388,N_2816);
and U4643 (N_4643,N_3400,N_2425);
and U4644 (N_4644,N_2696,N_3595);
or U4645 (N_4645,N_3452,N_2436);
and U4646 (N_4646,N_2550,N_3307);
xor U4647 (N_4647,N_2899,N_3112);
or U4648 (N_4648,N_2953,N_2913);
and U4649 (N_4649,N_3339,N_3400);
nand U4650 (N_4650,N_2840,N_3103);
nor U4651 (N_4651,N_2546,N_3201);
and U4652 (N_4652,N_3584,N_3436);
or U4653 (N_4653,N_3417,N_2517);
or U4654 (N_4654,N_3394,N_2787);
and U4655 (N_4655,N_3011,N_3165);
nor U4656 (N_4656,N_3022,N_3343);
or U4657 (N_4657,N_3525,N_2763);
or U4658 (N_4658,N_2636,N_2589);
nor U4659 (N_4659,N_3120,N_3332);
nor U4660 (N_4660,N_3315,N_2414);
xor U4661 (N_4661,N_2600,N_2491);
nand U4662 (N_4662,N_3525,N_2476);
nand U4663 (N_4663,N_3534,N_2901);
xnor U4664 (N_4664,N_2978,N_3136);
nand U4665 (N_4665,N_3493,N_2590);
nand U4666 (N_4666,N_3038,N_3556);
or U4667 (N_4667,N_3068,N_2783);
nand U4668 (N_4668,N_3151,N_3134);
nand U4669 (N_4669,N_3521,N_2423);
nand U4670 (N_4670,N_2897,N_2528);
nor U4671 (N_4671,N_3024,N_2687);
xor U4672 (N_4672,N_3004,N_2709);
nor U4673 (N_4673,N_3025,N_3270);
nand U4674 (N_4674,N_2625,N_3253);
and U4675 (N_4675,N_2494,N_2602);
xor U4676 (N_4676,N_3271,N_2668);
and U4677 (N_4677,N_2505,N_2563);
nor U4678 (N_4678,N_2515,N_3404);
or U4679 (N_4679,N_2580,N_2514);
or U4680 (N_4680,N_2712,N_3459);
nor U4681 (N_4681,N_2653,N_2904);
nand U4682 (N_4682,N_2598,N_3058);
nand U4683 (N_4683,N_3543,N_2678);
and U4684 (N_4684,N_3307,N_3396);
nor U4685 (N_4685,N_3478,N_2810);
nand U4686 (N_4686,N_3556,N_3310);
nand U4687 (N_4687,N_2911,N_2893);
xor U4688 (N_4688,N_2663,N_3016);
or U4689 (N_4689,N_2863,N_2641);
nor U4690 (N_4690,N_3254,N_2570);
or U4691 (N_4691,N_2993,N_2770);
nand U4692 (N_4692,N_3100,N_3437);
and U4693 (N_4693,N_2960,N_3581);
nand U4694 (N_4694,N_2502,N_2980);
nor U4695 (N_4695,N_3043,N_2857);
nor U4696 (N_4696,N_3501,N_2749);
or U4697 (N_4697,N_3051,N_2612);
nand U4698 (N_4698,N_3226,N_2485);
or U4699 (N_4699,N_2850,N_2983);
and U4700 (N_4700,N_2732,N_3004);
xor U4701 (N_4701,N_3563,N_3530);
xnor U4702 (N_4702,N_3475,N_2757);
nor U4703 (N_4703,N_3068,N_3318);
xnor U4704 (N_4704,N_2583,N_3264);
xor U4705 (N_4705,N_3426,N_3437);
nor U4706 (N_4706,N_2647,N_3488);
or U4707 (N_4707,N_2576,N_3007);
nand U4708 (N_4708,N_2759,N_2720);
xnor U4709 (N_4709,N_3450,N_3276);
nor U4710 (N_4710,N_2713,N_3234);
nor U4711 (N_4711,N_3050,N_2447);
and U4712 (N_4712,N_2798,N_3541);
nor U4713 (N_4713,N_3218,N_2647);
nor U4714 (N_4714,N_3577,N_3197);
and U4715 (N_4715,N_2606,N_2734);
and U4716 (N_4716,N_3395,N_2852);
and U4717 (N_4717,N_3364,N_2518);
or U4718 (N_4718,N_2879,N_3178);
and U4719 (N_4719,N_3117,N_3271);
or U4720 (N_4720,N_2548,N_2830);
or U4721 (N_4721,N_2719,N_3393);
nand U4722 (N_4722,N_3030,N_3487);
nand U4723 (N_4723,N_3256,N_2487);
nor U4724 (N_4724,N_2419,N_2887);
and U4725 (N_4725,N_2875,N_3196);
and U4726 (N_4726,N_2598,N_3553);
nand U4727 (N_4727,N_2679,N_3366);
or U4728 (N_4728,N_3023,N_2966);
nor U4729 (N_4729,N_2797,N_2614);
nand U4730 (N_4730,N_3492,N_2807);
xor U4731 (N_4731,N_3597,N_2727);
xnor U4732 (N_4732,N_3214,N_2414);
nor U4733 (N_4733,N_3126,N_3221);
xnor U4734 (N_4734,N_3529,N_3092);
and U4735 (N_4735,N_2907,N_3104);
nand U4736 (N_4736,N_3555,N_2730);
or U4737 (N_4737,N_2895,N_2695);
nor U4738 (N_4738,N_3001,N_2557);
or U4739 (N_4739,N_3519,N_2967);
nand U4740 (N_4740,N_3275,N_2617);
or U4741 (N_4741,N_3253,N_2554);
xor U4742 (N_4742,N_3031,N_3351);
nor U4743 (N_4743,N_2960,N_3057);
nor U4744 (N_4744,N_3135,N_2676);
xnor U4745 (N_4745,N_2854,N_2526);
xnor U4746 (N_4746,N_3407,N_3476);
nand U4747 (N_4747,N_2653,N_2578);
nor U4748 (N_4748,N_3241,N_3380);
nor U4749 (N_4749,N_3599,N_2936);
nand U4750 (N_4750,N_3449,N_2570);
xnor U4751 (N_4751,N_3120,N_2491);
xnor U4752 (N_4752,N_2574,N_2824);
xnor U4753 (N_4753,N_2502,N_3555);
nor U4754 (N_4754,N_3240,N_3156);
xnor U4755 (N_4755,N_2977,N_3104);
nand U4756 (N_4756,N_2915,N_3533);
nor U4757 (N_4757,N_3023,N_3002);
or U4758 (N_4758,N_2477,N_2701);
xor U4759 (N_4759,N_3297,N_3150);
xnor U4760 (N_4760,N_3477,N_3596);
xor U4761 (N_4761,N_2859,N_3356);
nand U4762 (N_4762,N_3164,N_3095);
nor U4763 (N_4763,N_3172,N_2507);
xor U4764 (N_4764,N_3082,N_3079);
xor U4765 (N_4765,N_2668,N_2550);
nor U4766 (N_4766,N_2424,N_2474);
nor U4767 (N_4767,N_2947,N_3504);
or U4768 (N_4768,N_2661,N_2437);
and U4769 (N_4769,N_2473,N_2915);
xnor U4770 (N_4770,N_2812,N_2705);
nand U4771 (N_4771,N_3159,N_3324);
nor U4772 (N_4772,N_2829,N_2534);
nor U4773 (N_4773,N_3080,N_3462);
or U4774 (N_4774,N_3210,N_2975);
and U4775 (N_4775,N_3067,N_3158);
nor U4776 (N_4776,N_2967,N_3438);
or U4777 (N_4777,N_2531,N_3435);
nor U4778 (N_4778,N_2961,N_2450);
nand U4779 (N_4779,N_2932,N_2586);
xor U4780 (N_4780,N_3260,N_2811);
xor U4781 (N_4781,N_3586,N_2907);
nand U4782 (N_4782,N_2986,N_3368);
and U4783 (N_4783,N_3588,N_3027);
nand U4784 (N_4784,N_3495,N_2504);
or U4785 (N_4785,N_2780,N_2990);
nand U4786 (N_4786,N_2801,N_2958);
nand U4787 (N_4787,N_3133,N_2490);
or U4788 (N_4788,N_2710,N_3036);
or U4789 (N_4789,N_3328,N_2601);
nand U4790 (N_4790,N_2644,N_3324);
nand U4791 (N_4791,N_3107,N_3193);
and U4792 (N_4792,N_2791,N_2872);
nand U4793 (N_4793,N_3484,N_3381);
or U4794 (N_4794,N_2830,N_2432);
xor U4795 (N_4795,N_3314,N_2993);
nor U4796 (N_4796,N_2825,N_3109);
nand U4797 (N_4797,N_2438,N_3332);
or U4798 (N_4798,N_3103,N_3229);
nor U4799 (N_4799,N_3111,N_3064);
and U4800 (N_4800,N_4442,N_4289);
and U4801 (N_4801,N_4444,N_3734);
xor U4802 (N_4802,N_4357,N_4416);
and U4803 (N_4803,N_4107,N_4235);
nand U4804 (N_4804,N_4712,N_3867);
or U4805 (N_4805,N_4630,N_4065);
or U4806 (N_4806,N_4632,N_4057);
xnor U4807 (N_4807,N_3646,N_4048);
and U4808 (N_4808,N_4350,N_3735);
or U4809 (N_4809,N_4422,N_4111);
xor U4810 (N_4810,N_4445,N_4251);
nand U4811 (N_4811,N_4672,N_4330);
nand U4812 (N_4812,N_4464,N_4655);
nand U4813 (N_4813,N_4227,N_4775);
xnor U4814 (N_4814,N_4402,N_3987);
xor U4815 (N_4815,N_4144,N_4301);
nand U4816 (N_4816,N_4625,N_4077);
or U4817 (N_4817,N_3747,N_3612);
nand U4818 (N_4818,N_3673,N_4224);
and U4819 (N_4819,N_4199,N_3997);
xor U4820 (N_4820,N_3977,N_4462);
xnor U4821 (N_4821,N_3767,N_4210);
nor U4822 (N_4822,N_3918,N_3848);
and U4823 (N_4823,N_4491,N_4501);
nor U4824 (N_4824,N_4098,N_4348);
and U4825 (N_4825,N_3793,N_3931);
and U4826 (N_4826,N_3781,N_4516);
or U4827 (N_4827,N_4038,N_4299);
xor U4828 (N_4828,N_4139,N_3661);
xnor U4829 (N_4829,N_3972,N_4087);
nor U4830 (N_4830,N_4668,N_3994);
nor U4831 (N_4831,N_4034,N_4053);
and U4832 (N_4832,N_4005,N_4008);
and U4833 (N_4833,N_3891,N_4537);
xor U4834 (N_4834,N_3785,N_4768);
or U4835 (N_4835,N_3899,N_3721);
nand U4836 (N_4836,N_4177,N_3946);
or U4837 (N_4837,N_3882,N_4322);
nand U4838 (N_4838,N_4435,N_4405);
nor U4839 (N_4839,N_4414,N_4636);
nor U4840 (N_4840,N_3700,N_4635);
and U4841 (N_4841,N_4453,N_3991);
and U4842 (N_4842,N_4595,N_4795);
or U4843 (N_4843,N_3880,N_4410);
and U4844 (N_4844,N_4764,N_4333);
nor U4845 (N_4845,N_4352,N_4508);
nand U4846 (N_4846,N_4606,N_4250);
xor U4847 (N_4847,N_3908,N_3716);
and U4848 (N_4848,N_4686,N_4489);
nand U4849 (N_4849,N_4398,N_3833);
xor U4850 (N_4850,N_4657,N_3690);
xnor U4851 (N_4851,N_3992,N_4495);
or U4852 (N_4852,N_4380,N_4736);
or U4853 (N_4853,N_4178,N_4497);
nand U4854 (N_4854,N_4066,N_4782);
xnor U4855 (N_4855,N_4571,N_4433);
xor U4856 (N_4856,N_4551,N_3702);
nand U4857 (N_4857,N_3657,N_4355);
and U4858 (N_4858,N_3851,N_4731);
nor U4859 (N_4859,N_3912,N_4513);
nor U4860 (N_4860,N_4628,N_3782);
and U4861 (N_4861,N_4786,N_4188);
xor U4862 (N_4862,N_4465,N_3671);
nor U4863 (N_4863,N_4600,N_4319);
or U4864 (N_4864,N_3663,N_3619);
and U4865 (N_4865,N_4158,N_4593);
nor U4866 (N_4866,N_3795,N_3729);
nand U4867 (N_4867,N_4719,N_4594);
nor U4868 (N_4868,N_4651,N_4585);
nor U4869 (N_4869,N_3834,N_3756);
and U4870 (N_4870,N_3944,N_4561);
nor U4871 (N_4871,N_3737,N_4086);
xor U4872 (N_4872,N_3950,N_4258);
xnor U4873 (N_4873,N_4016,N_4293);
nand U4874 (N_4874,N_4294,N_4223);
nand U4875 (N_4875,N_4679,N_3703);
nor U4876 (N_4876,N_3631,N_3772);
nor U4877 (N_4877,N_4316,N_4085);
and U4878 (N_4878,N_4794,N_3939);
and U4879 (N_4879,N_4225,N_4362);
or U4880 (N_4880,N_4543,N_4213);
nor U4881 (N_4881,N_4793,N_4326);
nand U4882 (N_4882,N_3965,N_4169);
xnor U4883 (N_4883,N_3879,N_3964);
or U4884 (N_4884,N_4419,N_4469);
nor U4885 (N_4885,N_4205,N_4649);
and U4886 (N_4886,N_4591,N_4529);
xor U4887 (N_4887,N_3788,N_4580);
nor U4888 (N_4888,N_3676,N_4041);
xnor U4889 (N_4889,N_4365,N_4612);
or U4890 (N_4890,N_4209,N_4351);
and U4891 (N_4891,N_4788,N_4339);
nand U4892 (N_4892,N_3632,N_3660);
and U4893 (N_4893,N_3794,N_3630);
nor U4894 (N_4894,N_3732,N_4661);
and U4895 (N_4895,N_3898,N_3618);
nand U4896 (N_4896,N_4285,N_4654);
xor U4897 (N_4897,N_4449,N_4153);
or U4898 (N_4898,N_3826,N_4597);
or U4899 (N_4899,N_4483,N_4259);
and U4900 (N_4900,N_4172,N_4438);
or U4901 (N_4901,N_3727,N_4255);
nand U4902 (N_4902,N_4109,N_4329);
nand U4903 (N_4903,N_4024,N_3780);
nor U4904 (N_4904,N_3865,N_4114);
xnor U4905 (N_4905,N_4072,N_4123);
nand U4906 (N_4906,N_3821,N_4187);
xor U4907 (N_4907,N_4681,N_4018);
or U4908 (N_4908,N_4396,N_4428);
nand U4909 (N_4909,N_4155,N_4650);
or U4910 (N_4910,N_3719,N_4602);
nor U4911 (N_4911,N_4700,N_4166);
or U4912 (N_4912,N_3850,N_3958);
or U4913 (N_4913,N_3973,N_4388);
xnor U4914 (N_4914,N_3776,N_4440);
nand U4915 (N_4915,N_4558,N_4590);
nor U4916 (N_4916,N_3611,N_4020);
xor U4917 (N_4917,N_4068,N_4218);
xnor U4918 (N_4918,N_4690,N_4372);
xor U4919 (N_4919,N_4532,N_3836);
nor U4920 (N_4920,N_4208,N_3853);
nand U4921 (N_4921,N_4554,N_4204);
nand U4922 (N_4922,N_3759,N_4479);
xor U4923 (N_4923,N_3903,N_3796);
xnor U4924 (N_4924,N_4017,N_4566);
or U4925 (N_4925,N_4658,N_4665);
nor U4926 (N_4926,N_4559,N_4673);
xor U4927 (N_4927,N_4079,N_4638);
and U4928 (N_4928,N_4785,N_4443);
and U4929 (N_4929,N_4182,N_4735);
or U4930 (N_4930,N_4070,N_3733);
nor U4931 (N_4931,N_3668,N_4173);
nor U4932 (N_4932,N_3600,N_4644);
nor U4933 (N_4933,N_4368,N_3815);
nand U4934 (N_4934,N_3686,N_4106);
xor U4935 (N_4935,N_3647,N_4674);
or U4936 (N_4936,N_3967,N_4721);
nor U4937 (N_4937,N_4221,N_4384);
or U4938 (N_4938,N_3816,N_4147);
nand U4939 (N_4939,N_4291,N_4090);
or U4940 (N_4940,N_4601,N_4050);
and U4941 (N_4941,N_3861,N_3937);
nand U4942 (N_4942,N_4001,N_4676);
xor U4943 (N_4943,N_4541,N_4014);
nor U4944 (N_4944,N_4143,N_3638);
nor U4945 (N_4945,N_3888,N_4149);
or U4946 (N_4946,N_4309,N_4547);
or U4947 (N_4947,N_4305,N_4332);
nor U4948 (N_4948,N_3860,N_3730);
nor U4949 (N_4949,N_4226,N_4728);
nor U4950 (N_4950,N_3909,N_4128);
and U4951 (N_4951,N_3707,N_4614);
xnor U4952 (N_4952,N_4525,N_4104);
xnor U4953 (N_4953,N_4279,N_3893);
and U4954 (N_4954,N_3910,N_4485);
nor U4955 (N_4955,N_4076,N_3832);
nand U4956 (N_4956,N_3731,N_4526);
nor U4957 (N_4957,N_4071,N_4015);
nor U4958 (N_4958,N_4287,N_4685);
nand U4959 (N_4959,N_3886,N_3960);
nor U4960 (N_4960,N_4539,N_3907);
or U4961 (N_4961,N_4011,N_4055);
xnor U4962 (N_4962,N_4564,N_4618);
or U4963 (N_4963,N_4583,N_3875);
or U4964 (N_4964,N_4371,N_3736);
nand U4965 (N_4965,N_3689,N_4069);
nand U4966 (N_4966,N_4607,N_4311);
xnor U4967 (N_4967,N_3890,N_4762);
and U4968 (N_4968,N_4779,N_4195);
nand U4969 (N_4969,N_3639,N_4113);
or U4970 (N_4970,N_3805,N_4254);
nand U4971 (N_4971,N_3922,N_3862);
and U4972 (N_4972,N_4486,N_3927);
xnor U4973 (N_4973,N_4133,N_4399);
and U4974 (N_4974,N_4103,N_4283);
nor U4975 (N_4975,N_3616,N_4563);
or U4976 (N_4976,N_4264,N_3644);
xor U4977 (N_4977,N_3741,N_4774);
xor U4978 (N_4978,N_3866,N_4385);
nand U4979 (N_4979,N_3985,N_3884);
nand U4980 (N_4980,N_4314,N_3629);
or U4981 (N_4981,N_4297,N_4022);
nand U4982 (N_4982,N_4688,N_4084);
nand U4983 (N_4983,N_3693,N_4027);
xor U4984 (N_4984,N_4080,N_3951);
nand U4985 (N_4985,N_4298,N_3758);
and U4986 (N_4986,N_4130,N_4303);
nand U4987 (N_4987,N_4490,N_3948);
nor U4988 (N_4988,N_4524,N_3718);
and U4989 (N_4989,N_3653,N_3670);
nand U4990 (N_4990,N_4536,N_4193);
xnor U4991 (N_4991,N_3803,N_4434);
nor U4992 (N_4992,N_4776,N_4167);
or U4993 (N_4993,N_3969,N_3777);
nor U4994 (N_4994,N_4129,N_3954);
or U4995 (N_4995,N_4122,N_4467);
or U4996 (N_4996,N_4540,N_4413);
nor U4997 (N_4997,N_3892,N_4457);
nand U4998 (N_4998,N_4589,N_4000);
xor U4999 (N_4999,N_3748,N_4089);
nand U5000 (N_5000,N_4535,N_3704);
and U5001 (N_5001,N_4270,N_3743);
nor U5002 (N_5002,N_4498,N_4707);
xnor U5003 (N_5003,N_4702,N_4450);
and U5004 (N_5004,N_4132,N_3986);
xnor U5005 (N_5005,N_4023,N_3620);
nor U5006 (N_5006,N_4184,N_4203);
nand U5007 (N_5007,N_4082,N_4722);
nor U5008 (N_5008,N_4765,N_4260);
nand U5009 (N_5009,N_4499,N_3911);
xnor U5010 (N_5010,N_3699,N_3941);
nor U5011 (N_5011,N_4755,N_4476);
nand U5012 (N_5012,N_4073,N_4494);
nor U5013 (N_5013,N_4481,N_4507);
and U5014 (N_5014,N_4401,N_4170);
xnor U5015 (N_5015,N_3768,N_4370);
nand U5016 (N_5016,N_4277,N_3666);
xor U5017 (N_5017,N_4427,N_3674);
nand U5018 (N_5018,N_4292,N_3936);
or U5019 (N_5019,N_4054,N_3827);
or U5020 (N_5020,N_4239,N_4318);
xnor U5021 (N_5021,N_4002,N_4036);
nor U5022 (N_5022,N_4281,N_3664);
xor U5023 (N_5023,N_4692,N_3685);
or U5024 (N_5024,N_4175,N_4390);
nor U5025 (N_5025,N_3728,N_4019);
and U5026 (N_5026,N_4096,N_4548);
or U5027 (N_5027,N_4446,N_3919);
xnor U5028 (N_5028,N_3824,N_4784);
nor U5029 (N_5029,N_3652,N_3672);
nor U5030 (N_5030,N_4186,N_4374);
and U5031 (N_5031,N_3812,N_3957);
and U5032 (N_5032,N_3831,N_4515);
and U5033 (N_5033,N_3687,N_4012);
and U5034 (N_5034,N_4615,N_4013);
xor U5035 (N_5035,N_3744,N_4771);
or U5036 (N_5036,N_4045,N_4337);
and U5037 (N_5037,N_3809,N_4117);
nor U5038 (N_5038,N_3988,N_4439);
nand U5039 (N_5039,N_4750,N_4431);
xnor U5040 (N_5040,N_3993,N_3874);
and U5041 (N_5041,N_4007,N_3738);
xor U5042 (N_5042,N_4200,N_4276);
xor U5043 (N_5043,N_3787,N_4032);
nand U5044 (N_5044,N_4101,N_3679);
nand U5045 (N_5045,N_4387,N_3749);
nand U5046 (N_5046,N_4544,N_4617);
nand U5047 (N_5047,N_4267,N_3692);
xnor U5048 (N_5048,N_4028,N_3771);
nand U5049 (N_5049,N_4509,N_4789);
or U5050 (N_5050,N_4487,N_3902);
nor U5051 (N_5051,N_3953,N_4646);
or U5052 (N_5052,N_3999,N_3746);
nand U5053 (N_5053,N_4713,N_4752);
xor U5054 (N_5054,N_3742,N_4461);
nor U5055 (N_5055,N_3799,N_3665);
xor U5056 (N_5056,N_4164,N_4408);
nand U5057 (N_5057,N_4426,N_3855);
xor U5058 (N_5058,N_4660,N_4029);
nand U5059 (N_5059,N_3921,N_4477);
nor U5060 (N_5060,N_4792,N_4386);
nand U5061 (N_5061,N_4502,N_4732);
nor U5062 (N_5062,N_4266,N_4631);
or U5063 (N_5063,N_3775,N_4466);
nand U5064 (N_5064,N_4772,N_4009);
nand U5065 (N_5065,N_3615,N_4474);
or U5066 (N_5066,N_4271,N_4748);
or U5067 (N_5067,N_3894,N_3872);
nor U5068 (N_5068,N_4582,N_4272);
or U5069 (N_5069,N_3932,N_3819);
xnor U5070 (N_5070,N_4245,N_4165);
nor U5071 (N_5071,N_3998,N_4237);
nor U5072 (N_5072,N_4240,N_3792);
nand U5073 (N_5073,N_4341,N_3636);
nand U5074 (N_5074,N_3797,N_4206);
nand U5075 (N_5075,N_4634,N_3650);
nor U5076 (N_5076,N_4244,N_4214);
xnor U5077 (N_5077,N_4436,N_4302);
and U5078 (N_5078,N_3962,N_4714);
xnor U5079 (N_5079,N_3895,N_4257);
and U5080 (N_5080,N_3837,N_3779);
and U5081 (N_5081,N_3971,N_4236);
and U5082 (N_5082,N_4609,N_4691);
and U5083 (N_5083,N_4137,N_4049);
xor U5084 (N_5084,N_4729,N_3938);
nor U5085 (N_5085,N_3889,N_3863);
nor U5086 (N_5086,N_4693,N_4003);
or U5087 (N_5087,N_4643,N_4740);
xor U5088 (N_5088,N_4246,N_3696);
xnor U5089 (N_5089,N_3930,N_4152);
or U5090 (N_5090,N_3983,N_4093);
and U5091 (N_5091,N_3876,N_4192);
and U5092 (N_5092,N_3975,N_4215);
and U5093 (N_5093,N_3801,N_3854);
nand U5094 (N_5094,N_3804,N_3655);
xor U5095 (N_5095,N_3818,N_4092);
xnor U5096 (N_5096,N_3712,N_4162);
xor U5097 (N_5097,N_4517,N_3789);
nand U5098 (N_5098,N_4799,N_4262);
or U5099 (N_5099,N_4503,N_3933);
nand U5100 (N_5100,N_4207,N_4656);
and U5101 (N_5101,N_4629,N_4340);
xnor U5102 (N_5102,N_4669,N_3949);
or U5103 (N_5103,N_3617,N_3849);
nor U5104 (N_5104,N_4230,N_4754);
nand U5105 (N_5105,N_4376,N_3887);
xnor U5106 (N_5106,N_4040,N_4542);
and U5107 (N_5107,N_4484,N_3607);
and U5108 (N_5108,N_4626,N_4611);
nor U5109 (N_5109,N_3806,N_3928);
xnor U5110 (N_5110,N_4640,N_4773);
and U5111 (N_5111,N_3979,N_4252);
xor U5112 (N_5112,N_4010,N_4409);
xor U5113 (N_5113,N_4778,N_4504);
or U5114 (N_5114,N_4592,N_4284);
nor U5115 (N_5115,N_4478,N_4201);
nand U5116 (N_5116,N_4286,N_3810);
and U5117 (N_5117,N_4342,N_4708);
nand U5118 (N_5118,N_3642,N_4531);
or U5119 (N_5119,N_3774,N_4421);
or U5120 (N_5120,N_3725,N_4154);
and U5121 (N_5121,N_3830,N_3978);
nand U5122 (N_5122,N_4480,N_4407);
xnor U5123 (N_5123,N_3996,N_4605);
xor U5124 (N_5124,N_4150,N_3681);
and U5125 (N_5125,N_4567,N_4705);
nor U5126 (N_5126,N_4671,N_4046);
nor U5127 (N_5127,N_4397,N_4569);
nor U5128 (N_5128,N_4088,N_3981);
or U5129 (N_5129,N_4021,N_3814);
or U5130 (N_5130,N_4608,N_3751);
xor U5131 (N_5131,N_3845,N_3745);
nand U5132 (N_5132,N_4345,N_4336);
nand U5133 (N_5133,N_3651,N_4288);
nand U5134 (N_5134,N_4623,N_3838);
xnor U5135 (N_5135,N_4570,N_4698);
and U5136 (N_5136,N_4232,N_4664);
and U5137 (N_5137,N_4482,N_3857);
and U5138 (N_5138,N_4417,N_4110);
xor U5139 (N_5139,N_4124,N_3995);
xor U5140 (N_5140,N_4620,N_4511);
xnor U5141 (N_5141,N_3858,N_4043);
nor U5142 (N_5142,N_3669,N_4538);
xor U5143 (N_5143,N_4358,N_4697);
or U5144 (N_5144,N_4361,N_4190);
nor U5145 (N_5145,N_3688,N_4727);
or U5146 (N_5146,N_4151,N_3705);
nand U5147 (N_5147,N_4521,N_4546);
nand U5148 (N_5148,N_4168,N_3641);
or U5149 (N_5149,N_4198,N_4556);
nand U5150 (N_5150,N_4471,N_4389);
and U5151 (N_5151,N_4052,N_3697);
or U5152 (N_5152,N_4217,N_3610);
nor U5153 (N_5153,N_4183,N_4115);
or U5154 (N_5154,N_4458,N_4378);
and U5155 (N_5155,N_3963,N_4747);
or U5156 (N_5156,N_4328,N_3701);
and U5157 (N_5157,N_4573,N_4031);
xor U5158 (N_5158,N_4300,N_4598);
nor U5159 (N_5159,N_4709,N_3913);
or U5160 (N_5160,N_3713,N_4621);
nor U5161 (N_5161,N_3762,N_3637);
or U5162 (N_5162,N_3813,N_3835);
and U5163 (N_5163,N_4488,N_4346);
nand U5164 (N_5164,N_4060,N_4758);
xnor U5165 (N_5165,N_4701,N_4759);
nand U5166 (N_5166,N_3869,N_3925);
or U5167 (N_5167,N_4159,N_3926);
nor U5168 (N_5168,N_4738,N_4290);
or U5169 (N_5169,N_3829,N_4095);
or U5170 (N_5170,N_3976,N_4734);
nor U5171 (N_5171,N_4145,N_4064);
nor U5172 (N_5172,N_4039,N_4797);
nand U5173 (N_5173,N_4062,N_4241);
and U5174 (N_5174,N_3843,N_3714);
xor U5175 (N_5175,N_3807,N_4506);
xnor U5176 (N_5176,N_4141,N_3739);
xor U5177 (N_5177,N_3773,N_4745);
nand U5178 (N_5178,N_4472,N_4131);
and U5179 (N_5179,N_3635,N_3622);
or U5180 (N_5180,N_4753,N_4717);
or U5181 (N_5181,N_4675,N_4560);
nand U5182 (N_5182,N_4798,N_3691);
xnor U5183 (N_5183,N_4059,N_4505);
and U5184 (N_5184,N_4704,N_4061);
nand U5185 (N_5185,N_4770,N_4706);
xor U5186 (N_5186,N_4033,N_4211);
and U5187 (N_5187,N_4557,N_4249);
nand U5188 (N_5188,N_3900,N_3760);
or U5189 (N_5189,N_3820,N_3839);
nand U5190 (N_5190,N_4194,N_3765);
or U5191 (N_5191,N_4716,N_4306);
nand U5192 (N_5192,N_4456,N_4603);
xnor U5193 (N_5193,N_4323,N_4581);
or U5194 (N_5194,N_3947,N_4148);
and U5195 (N_5195,N_4425,N_4500);
and U5196 (N_5196,N_4682,N_4663);
xnor U5197 (N_5197,N_3959,N_3915);
and U5198 (N_5198,N_4684,N_3723);
and U5199 (N_5199,N_3984,N_4613);
or U5200 (N_5200,N_4725,N_4596);
nor U5201 (N_5201,N_3766,N_4334);
xnor U5202 (N_5202,N_4231,N_4324);
xnor U5203 (N_5203,N_3614,N_3873);
xnor U5204 (N_5204,N_4174,N_4733);
nand U5205 (N_5205,N_4624,N_4238);
or U5206 (N_5206,N_4622,N_4633);
or U5207 (N_5207,N_4473,N_4599);
nand U5208 (N_5208,N_4379,N_4648);
nand U5209 (N_5209,N_4423,N_4761);
nand U5210 (N_5210,N_3790,N_3753);
nor U5211 (N_5211,N_3877,N_4575);
nor U5212 (N_5212,N_4261,N_4377);
and U5213 (N_5213,N_3924,N_4448);
nand U5214 (N_5214,N_4452,N_4138);
nand U5215 (N_5215,N_4746,N_3828);
or U5216 (N_5216,N_4578,N_4662);
nor U5217 (N_5217,N_3945,N_3694);
and U5218 (N_5218,N_4102,N_4185);
xnor U5219 (N_5219,N_4367,N_4268);
or U5220 (N_5220,N_4647,N_4263);
nor U5221 (N_5221,N_4530,N_4790);
and U5222 (N_5222,N_4097,N_4687);
xnor U5223 (N_5223,N_3761,N_4404);
nor U5224 (N_5224,N_4335,N_4562);
nor U5225 (N_5225,N_3608,N_3883);
nor U5226 (N_5226,N_3982,N_4741);
or U5227 (N_5227,N_3621,N_3906);
nand U5228 (N_5228,N_4363,N_4760);
or U5229 (N_5229,N_4455,N_4512);
xnor U5230 (N_5230,N_3659,N_4191);
xor U5231 (N_5231,N_4161,N_4459);
or U5232 (N_5232,N_3956,N_4395);
or U5233 (N_5233,N_3715,N_4220);
nor U5234 (N_5234,N_3808,N_4470);
xor U5235 (N_5235,N_3920,N_4550);
nor U5236 (N_5236,N_4689,N_3706);
and U5237 (N_5237,N_3648,N_3868);
and U5238 (N_5238,N_3800,N_4047);
nand U5239 (N_5239,N_4584,N_4075);
and U5240 (N_5240,N_4756,N_3859);
nor U5241 (N_5241,N_4763,N_4242);
or U5242 (N_5242,N_3825,N_3896);
nand U5243 (N_5243,N_4181,N_4534);
xor U5244 (N_5244,N_4694,N_4228);
or U5245 (N_5245,N_4121,N_4275);
or U5246 (N_5246,N_4766,N_4248);
nand U5247 (N_5247,N_4437,N_4383);
or U5248 (N_5248,N_3656,N_4780);
xnor U5249 (N_5249,N_4791,N_3940);
nor U5250 (N_5250,N_4025,N_3634);
and U5251 (N_5251,N_4222,N_4710);
xor U5252 (N_5252,N_4653,N_4321);
nand U5253 (N_5253,N_4418,N_4777);
nand U5254 (N_5254,N_4751,N_4545);
and U5255 (N_5255,N_4278,N_4394);
xor U5256 (N_5256,N_4347,N_4274);
nand U5257 (N_5257,N_4156,N_4296);
nand U5258 (N_5258,N_4269,N_4572);
xnor U5259 (N_5259,N_4447,N_4094);
and U5260 (N_5260,N_4724,N_3606);
nor U5261 (N_5261,N_4726,N_4680);
and U5262 (N_5262,N_4670,N_3904);
or U5263 (N_5263,N_3966,N_4247);
or U5264 (N_5264,N_4282,N_4796);
nand U5265 (N_5265,N_3840,N_4787);
or U5266 (N_5266,N_4140,N_3914);
or U5267 (N_5267,N_4699,N_4730);
nand U5268 (N_5268,N_4574,N_4233);
xor U5269 (N_5269,N_4677,N_4520);
xor U5270 (N_5270,N_4441,N_3717);
nor U5271 (N_5271,N_4415,N_3764);
nor U5272 (N_5272,N_4108,N_3624);
nor U5273 (N_5273,N_3989,N_3658);
nand U5274 (N_5274,N_4616,N_3802);
nand U5275 (N_5275,N_3625,N_4749);
and U5276 (N_5276,N_3602,N_4171);
and U5277 (N_5277,N_4100,N_4577);
nor U5278 (N_5278,N_3628,N_4586);
nand U5279 (N_5279,N_4392,N_3923);
or U5280 (N_5280,N_4134,N_3935);
nor U5281 (N_5281,N_4313,N_4783);
or U5282 (N_5282,N_4604,N_4619);
nor U5283 (N_5283,N_4645,N_3823);
and U5284 (N_5284,N_3881,N_4006);
nand U5285 (N_5285,N_4234,N_3757);
and U5286 (N_5286,N_4666,N_4667);
xor U5287 (N_5287,N_4696,N_4179);
and U5288 (N_5288,N_3968,N_4136);
nor U5289 (N_5289,N_3842,N_4781);
xor U5290 (N_5290,N_4579,N_4514);
nand U5291 (N_5291,N_3662,N_4492);
xor U5292 (N_5292,N_3677,N_3990);
nor U5293 (N_5293,N_3710,N_3955);
and U5294 (N_5294,N_4627,N_4081);
nand U5295 (N_5295,N_3609,N_4125);
nor U5296 (N_5296,N_3708,N_4051);
or U5297 (N_5297,N_4451,N_4099);
or U5298 (N_5298,N_3934,N_3871);
xor U5299 (N_5299,N_4127,N_3822);
nor U5300 (N_5300,N_4243,N_3916);
nor U5301 (N_5301,N_4202,N_4463);
nand U5302 (N_5302,N_4400,N_3878);
xor U5303 (N_5303,N_3952,N_3649);
and U5304 (N_5304,N_3841,N_4366);
nand U5305 (N_5305,N_4711,N_4430);
and U5306 (N_5306,N_4157,N_4118);
xor U5307 (N_5307,N_4338,N_4468);
nand U5308 (N_5308,N_4044,N_3791);
nand U5309 (N_5309,N_3846,N_4273);
and U5310 (N_5310,N_4256,N_4120);
nor U5311 (N_5311,N_4229,N_3740);
nor U5312 (N_5312,N_3942,N_3623);
xor U5313 (N_5313,N_4331,N_4349);
and U5314 (N_5314,N_4555,N_4105);
nor U5315 (N_5315,N_3605,N_4160);
nor U5316 (N_5316,N_4091,N_4119);
nor U5317 (N_5317,N_4610,N_4429);
and U5318 (N_5318,N_4343,N_3724);
or U5319 (N_5319,N_3682,N_3974);
or U5320 (N_5320,N_4126,N_4116);
or U5321 (N_5321,N_3769,N_4587);
and U5322 (N_5322,N_3763,N_4769);
and U5323 (N_5323,N_4354,N_3654);
nor U5324 (N_5324,N_4325,N_4359);
and U5325 (N_5325,N_4381,N_4063);
nor U5326 (N_5326,N_4637,N_4035);
xor U5327 (N_5327,N_4743,N_3667);
xor U5328 (N_5328,N_3885,N_3943);
xor U5329 (N_5329,N_3684,N_3601);
nor U5330 (N_5330,N_3778,N_4510);
or U5331 (N_5331,N_4420,N_4373);
or U5332 (N_5332,N_4533,N_4552);
and U5333 (N_5333,N_4742,N_3678);
xor U5334 (N_5334,N_4307,N_3929);
nor U5335 (N_5335,N_3711,N_3852);
or U5336 (N_5336,N_4360,N_3695);
xor U5337 (N_5337,N_4056,N_4432);
or U5338 (N_5338,N_3961,N_4553);
nor U5339 (N_5339,N_4744,N_3798);
or U5340 (N_5340,N_3698,N_3722);
nand U5341 (N_5341,N_3783,N_4315);
nand U5342 (N_5342,N_4652,N_4004);
nor U5343 (N_5343,N_3897,N_4767);
xor U5344 (N_5344,N_3754,N_4320);
xnor U5345 (N_5345,N_4026,N_3817);
nor U5346 (N_5346,N_3627,N_3752);
nand U5347 (N_5347,N_3640,N_4382);
or U5348 (N_5348,N_4083,N_4216);
or U5349 (N_5349,N_4720,N_3726);
and U5350 (N_5350,N_4424,N_4412);
or U5351 (N_5351,N_4037,N_4163);
nand U5352 (N_5352,N_4527,N_4518);
or U5353 (N_5353,N_3720,N_4523);
nor U5354 (N_5354,N_3755,N_4391);
or U5355 (N_5355,N_4723,N_4739);
nor U5356 (N_5356,N_3856,N_4310);
xnor U5357 (N_5357,N_3864,N_4030);
and U5358 (N_5358,N_4067,N_3980);
and U5359 (N_5359,N_3683,N_4393);
nand U5360 (N_5360,N_4568,N_4280);
xor U5361 (N_5361,N_4253,N_4454);
and U5362 (N_5362,N_4074,N_4212);
or U5363 (N_5363,N_4549,N_4308);
nand U5364 (N_5364,N_4496,N_4327);
nand U5365 (N_5365,N_4189,N_3770);
nor U5366 (N_5366,N_4683,N_4265);
and U5367 (N_5367,N_4715,N_3901);
nand U5368 (N_5368,N_4356,N_4353);
or U5369 (N_5369,N_4703,N_4522);
and U5370 (N_5370,N_4757,N_3970);
nor U5371 (N_5371,N_3613,N_4369);
and U5372 (N_5372,N_3643,N_3784);
and U5373 (N_5373,N_4058,N_4317);
nand U5374 (N_5374,N_4460,N_3633);
nor U5375 (N_5375,N_4219,N_4196);
or U5376 (N_5376,N_4406,N_3709);
nor U5377 (N_5377,N_3604,N_4659);
or U5378 (N_5378,N_3645,N_4176);
xnor U5379 (N_5379,N_4180,N_4364);
nand U5380 (N_5380,N_4588,N_3750);
nor U5381 (N_5381,N_3603,N_4146);
nor U5382 (N_5382,N_3626,N_3786);
or U5383 (N_5383,N_3844,N_4678);
and U5384 (N_5384,N_4639,N_3905);
xnor U5385 (N_5385,N_4493,N_4737);
nor U5386 (N_5386,N_4576,N_4312);
nor U5387 (N_5387,N_4375,N_3680);
and U5388 (N_5388,N_4642,N_3811);
nand U5389 (N_5389,N_4295,N_3870);
or U5390 (N_5390,N_4411,N_3675);
nor U5391 (N_5391,N_4344,N_4528);
nand U5392 (N_5392,N_3917,N_3847);
nand U5393 (N_5393,N_4641,N_4112);
xnor U5394 (N_5394,N_4695,N_4304);
nand U5395 (N_5395,N_4519,N_4042);
xor U5396 (N_5396,N_4197,N_4718);
nand U5397 (N_5397,N_4403,N_4142);
or U5398 (N_5398,N_4565,N_4078);
xnor U5399 (N_5399,N_4475,N_4135);
nor U5400 (N_5400,N_4090,N_4094);
nor U5401 (N_5401,N_3683,N_4191);
and U5402 (N_5402,N_4320,N_4038);
xnor U5403 (N_5403,N_3624,N_4650);
xor U5404 (N_5404,N_3913,N_3710);
and U5405 (N_5405,N_4034,N_3860);
xor U5406 (N_5406,N_3986,N_3785);
and U5407 (N_5407,N_4178,N_4714);
or U5408 (N_5408,N_4370,N_4742);
or U5409 (N_5409,N_3682,N_4512);
xor U5410 (N_5410,N_4093,N_4007);
xnor U5411 (N_5411,N_3920,N_3740);
nor U5412 (N_5412,N_3640,N_4087);
or U5413 (N_5413,N_4340,N_4283);
nand U5414 (N_5414,N_4435,N_3846);
or U5415 (N_5415,N_3608,N_3737);
and U5416 (N_5416,N_4032,N_4241);
nand U5417 (N_5417,N_3957,N_4592);
nand U5418 (N_5418,N_4475,N_4563);
nand U5419 (N_5419,N_3621,N_4667);
nor U5420 (N_5420,N_4281,N_3760);
or U5421 (N_5421,N_3783,N_4563);
or U5422 (N_5422,N_3948,N_4277);
or U5423 (N_5423,N_3993,N_4095);
and U5424 (N_5424,N_4019,N_4325);
nor U5425 (N_5425,N_4263,N_4255);
xnor U5426 (N_5426,N_3813,N_3742);
nor U5427 (N_5427,N_4416,N_3674);
nand U5428 (N_5428,N_3965,N_4707);
nand U5429 (N_5429,N_3793,N_4475);
nand U5430 (N_5430,N_4246,N_4492);
and U5431 (N_5431,N_3806,N_4601);
xor U5432 (N_5432,N_4307,N_4104);
xor U5433 (N_5433,N_3694,N_4009);
nor U5434 (N_5434,N_3738,N_4730);
and U5435 (N_5435,N_4030,N_3752);
and U5436 (N_5436,N_3927,N_4099);
nand U5437 (N_5437,N_4277,N_4011);
nor U5438 (N_5438,N_4466,N_4765);
nor U5439 (N_5439,N_4468,N_4513);
xor U5440 (N_5440,N_3659,N_3931);
nor U5441 (N_5441,N_4612,N_3867);
or U5442 (N_5442,N_3840,N_3617);
or U5443 (N_5443,N_4571,N_4247);
xnor U5444 (N_5444,N_4400,N_4752);
nor U5445 (N_5445,N_3739,N_4261);
xnor U5446 (N_5446,N_4744,N_4546);
nor U5447 (N_5447,N_4112,N_4619);
xor U5448 (N_5448,N_4113,N_4398);
xnor U5449 (N_5449,N_4435,N_3716);
xnor U5450 (N_5450,N_3718,N_3974);
nand U5451 (N_5451,N_3981,N_4097);
and U5452 (N_5452,N_4440,N_4615);
nand U5453 (N_5453,N_4411,N_4357);
nor U5454 (N_5454,N_4327,N_3780);
nand U5455 (N_5455,N_3983,N_4664);
xor U5456 (N_5456,N_4010,N_4568);
nor U5457 (N_5457,N_4435,N_4327);
nand U5458 (N_5458,N_4496,N_4547);
or U5459 (N_5459,N_3726,N_4286);
nand U5460 (N_5460,N_4279,N_4183);
nand U5461 (N_5461,N_4334,N_4436);
xor U5462 (N_5462,N_4782,N_3881);
and U5463 (N_5463,N_3713,N_4220);
nor U5464 (N_5464,N_4420,N_4018);
or U5465 (N_5465,N_4676,N_4537);
xnor U5466 (N_5466,N_4200,N_4664);
xor U5467 (N_5467,N_4248,N_3673);
or U5468 (N_5468,N_4279,N_4450);
and U5469 (N_5469,N_3728,N_3844);
or U5470 (N_5470,N_4308,N_3820);
nand U5471 (N_5471,N_4654,N_4160);
nand U5472 (N_5472,N_3612,N_3846);
nor U5473 (N_5473,N_3969,N_4213);
xnor U5474 (N_5474,N_4191,N_3602);
xor U5475 (N_5475,N_4714,N_4135);
nor U5476 (N_5476,N_4024,N_4183);
nand U5477 (N_5477,N_3816,N_3884);
and U5478 (N_5478,N_3753,N_3829);
or U5479 (N_5479,N_3829,N_3794);
xor U5480 (N_5480,N_4624,N_3767);
or U5481 (N_5481,N_4698,N_4497);
and U5482 (N_5482,N_3711,N_4633);
or U5483 (N_5483,N_3803,N_4008);
or U5484 (N_5484,N_3625,N_3697);
nor U5485 (N_5485,N_4271,N_3927);
and U5486 (N_5486,N_3999,N_3725);
xnor U5487 (N_5487,N_3948,N_3882);
nand U5488 (N_5488,N_4719,N_4622);
xnor U5489 (N_5489,N_4677,N_4739);
or U5490 (N_5490,N_3995,N_3892);
nor U5491 (N_5491,N_3677,N_3831);
and U5492 (N_5492,N_4064,N_4437);
or U5493 (N_5493,N_4418,N_4793);
nand U5494 (N_5494,N_4397,N_4541);
nor U5495 (N_5495,N_3789,N_4490);
nand U5496 (N_5496,N_4124,N_4651);
xnor U5497 (N_5497,N_4100,N_3768);
nand U5498 (N_5498,N_3839,N_4725);
nor U5499 (N_5499,N_4524,N_3943);
nand U5500 (N_5500,N_4353,N_4231);
xor U5501 (N_5501,N_4770,N_4003);
nor U5502 (N_5502,N_4040,N_4492);
or U5503 (N_5503,N_3773,N_4702);
and U5504 (N_5504,N_4238,N_4705);
nor U5505 (N_5505,N_4185,N_3738);
nor U5506 (N_5506,N_3756,N_4069);
nor U5507 (N_5507,N_4680,N_4723);
xnor U5508 (N_5508,N_3763,N_4059);
nor U5509 (N_5509,N_4789,N_3641);
xnor U5510 (N_5510,N_3609,N_3778);
and U5511 (N_5511,N_3904,N_3722);
nand U5512 (N_5512,N_3908,N_4610);
or U5513 (N_5513,N_4770,N_4238);
and U5514 (N_5514,N_3957,N_4367);
nand U5515 (N_5515,N_3789,N_4374);
and U5516 (N_5516,N_4176,N_4564);
and U5517 (N_5517,N_4010,N_4110);
nor U5518 (N_5518,N_4609,N_4413);
or U5519 (N_5519,N_4272,N_4610);
nand U5520 (N_5520,N_4376,N_4134);
or U5521 (N_5521,N_4498,N_4147);
nand U5522 (N_5522,N_3980,N_4553);
xnor U5523 (N_5523,N_4421,N_4096);
and U5524 (N_5524,N_4710,N_4120);
or U5525 (N_5525,N_4155,N_4597);
nand U5526 (N_5526,N_3933,N_3608);
nand U5527 (N_5527,N_3921,N_3923);
and U5528 (N_5528,N_4075,N_3672);
and U5529 (N_5529,N_4098,N_4674);
and U5530 (N_5530,N_4067,N_3609);
and U5531 (N_5531,N_3802,N_4169);
and U5532 (N_5532,N_4584,N_4307);
nand U5533 (N_5533,N_3606,N_3835);
nor U5534 (N_5534,N_4135,N_3617);
nor U5535 (N_5535,N_4280,N_4698);
nor U5536 (N_5536,N_4131,N_3730);
or U5537 (N_5537,N_3647,N_3793);
and U5538 (N_5538,N_3889,N_4092);
nand U5539 (N_5539,N_4104,N_4488);
xor U5540 (N_5540,N_4734,N_4501);
xor U5541 (N_5541,N_4066,N_3703);
nor U5542 (N_5542,N_4140,N_3832);
nor U5543 (N_5543,N_4414,N_4747);
or U5544 (N_5544,N_4654,N_4431);
and U5545 (N_5545,N_3712,N_4361);
and U5546 (N_5546,N_4727,N_3739);
nand U5547 (N_5547,N_4262,N_4213);
or U5548 (N_5548,N_3836,N_4186);
nor U5549 (N_5549,N_4739,N_3728);
xnor U5550 (N_5550,N_3699,N_4421);
nor U5551 (N_5551,N_3950,N_4588);
nand U5552 (N_5552,N_3974,N_4586);
xor U5553 (N_5553,N_4203,N_4577);
nor U5554 (N_5554,N_3706,N_4513);
nand U5555 (N_5555,N_4533,N_3832);
nor U5556 (N_5556,N_4773,N_4548);
nor U5557 (N_5557,N_3661,N_4001);
nor U5558 (N_5558,N_4071,N_4373);
xnor U5559 (N_5559,N_3608,N_4738);
or U5560 (N_5560,N_4330,N_4110);
xnor U5561 (N_5561,N_3717,N_3679);
nand U5562 (N_5562,N_3697,N_4618);
or U5563 (N_5563,N_3728,N_4303);
nor U5564 (N_5564,N_4051,N_3897);
and U5565 (N_5565,N_3696,N_3709);
or U5566 (N_5566,N_4385,N_3790);
nand U5567 (N_5567,N_3655,N_4096);
nand U5568 (N_5568,N_4361,N_3939);
nor U5569 (N_5569,N_4669,N_4798);
or U5570 (N_5570,N_4444,N_4652);
and U5571 (N_5571,N_4367,N_4255);
or U5572 (N_5572,N_4222,N_4023);
nand U5573 (N_5573,N_4105,N_3801);
nand U5574 (N_5574,N_3783,N_4673);
nor U5575 (N_5575,N_4478,N_4375);
nand U5576 (N_5576,N_3734,N_4679);
xnor U5577 (N_5577,N_3975,N_3969);
xor U5578 (N_5578,N_3760,N_4632);
nand U5579 (N_5579,N_4508,N_4662);
or U5580 (N_5580,N_4571,N_4070);
nor U5581 (N_5581,N_4235,N_3991);
nor U5582 (N_5582,N_4719,N_3664);
and U5583 (N_5583,N_4363,N_4527);
or U5584 (N_5584,N_4726,N_3856);
xor U5585 (N_5585,N_4293,N_3953);
or U5586 (N_5586,N_4234,N_4218);
nor U5587 (N_5587,N_4487,N_3692);
xor U5588 (N_5588,N_3782,N_3849);
and U5589 (N_5589,N_4078,N_4542);
or U5590 (N_5590,N_4741,N_4283);
or U5591 (N_5591,N_4615,N_3695);
nor U5592 (N_5592,N_4076,N_4132);
or U5593 (N_5593,N_3884,N_4610);
nor U5594 (N_5594,N_4142,N_4165);
and U5595 (N_5595,N_4193,N_4037);
nor U5596 (N_5596,N_3891,N_3945);
xnor U5597 (N_5597,N_4470,N_4559);
xor U5598 (N_5598,N_3801,N_4377);
or U5599 (N_5599,N_3908,N_4243);
nor U5600 (N_5600,N_4415,N_3938);
nand U5601 (N_5601,N_3741,N_3705);
or U5602 (N_5602,N_4684,N_3734);
or U5603 (N_5603,N_3789,N_4680);
and U5604 (N_5604,N_4568,N_4356);
and U5605 (N_5605,N_4717,N_4254);
xnor U5606 (N_5606,N_3808,N_3858);
and U5607 (N_5607,N_4657,N_3819);
or U5608 (N_5608,N_3658,N_3984);
nor U5609 (N_5609,N_3878,N_4200);
nand U5610 (N_5610,N_3747,N_3795);
or U5611 (N_5611,N_4264,N_4401);
xor U5612 (N_5612,N_4417,N_4633);
nand U5613 (N_5613,N_3668,N_4546);
or U5614 (N_5614,N_4705,N_4427);
or U5615 (N_5615,N_4121,N_4497);
and U5616 (N_5616,N_3793,N_3946);
xor U5617 (N_5617,N_3800,N_4796);
and U5618 (N_5618,N_4784,N_3944);
or U5619 (N_5619,N_4438,N_3980);
nor U5620 (N_5620,N_3894,N_3652);
nand U5621 (N_5621,N_4178,N_4669);
nand U5622 (N_5622,N_4553,N_4709);
and U5623 (N_5623,N_4405,N_4668);
nor U5624 (N_5624,N_4021,N_3834);
nand U5625 (N_5625,N_4201,N_4273);
xor U5626 (N_5626,N_4477,N_3818);
xor U5627 (N_5627,N_4141,N_4266);
nor U5628 (N_5628,N_3837,N_4060);
nand U5629 (N_5629,N_3971,N_4162);
nor U5630 (N_5630,N_4206,N_3665);
nor U5631 (N_5631,N_4448,N_4273);
nor U5632 (N_5632,N_4315,N_4494);
xor U5633 (N_5633,N_3695,N_4511);
nor U5634 (N_5634,N_3707,N_4474);
nand U5635 (N_5635,N_3730,N_4662);
or U5636 (N_5636,N_3693,N_3858);
and U5637 (N_5637,N_4196,N_4056);
xor U5638 (N_5638,N_4183,N_4708);
nor U5639 (N_5639,N_4726,N_4166);
nor U5640 (N_5640,N_4252,N_4386);
xor U5641 (N_5641,N_4626,N_4334);
or U5642 (N_5642,N_3828,N_3713);
nand U5643 (N_5643,N_4581,N_3725);
nor U5644 (N_5644,N_3725,N_4699);
xor U5645 (N_5645,N_3655,N_4551);
nor U5646 (N_5646,N_3614,N_4354);
or U5647 (N_5647,N_4575,N_3758);
xnor U5648 (N_5648,N_4174,N_4631);
nor U5649 (N_5649,N_4770,N_4515);
and U5650 (N_5650,N_4302,N_3685);
and U5651 (N_5651,N_4119,N_4306);
nand U5652 (N_5652,N_4722,N_3721);
xnor U5653 (N_5653,N_4605,N_4789);
nand U5654 (N_5654,N_3995,N_4070);
and U5655 (N_5655,N_4207,N_4103);
nand U5656 (N_5656,N_3900,N_4338);
nand U5657 (N_5657,N_3648,N_4799);
nand U5658 (N_5658,N_4755,N_3839);
or U5659 (N_5659,N_4445,N_4490);
xnor U5660 (N_5660,N_4764,N_3701);
and U5661 (N_5661,N_3957,N_3933);
or U5662 (N_5662,N_4120,N_4525);
nor U5663 (N_5663,N_3889,N_3739);
xnor U5664 (N_5664,N_3746,N_4215);
nor U5665 (N_5665,N_3767,N_4197);
or U5666 (N_5666,N_4016,N_4281);
xnor U5667 (N_5667,N_3833,N_4246);
nor U5668 (N_5668,N_3794,N_4154);
or U5669 (N_5669,N_4661,N_3621);
or U5670 (N_5670,N_4152,N_3636);
xnor U5671 (N_5671,N_4644,N_4453);
nand U5672 (N_5672,N_4278,N_4117);
nand U5673 (N_5673,N_3815,N_4332);
and U5674 (N_5674,N_4307,N_4306);
nor U5675 (N_5675,N_4568,N_4389);
and U5676 (N_5676,N_3790,N_3602);
nand U5677 (N_5677,N_3660,N_3859);
xnor U5678 (N_5678,N_3733,N_4083);
xor U5679 (N_5679,N_3931,N_4448);
nand U5680 (N_5680,N_4746,N_4771);
and U5681 (N_5681,N_4018,N_3677);
nand U5682 (N_5682,N_4672,N_3727);
nor U5683 (N_5683,N_4323,N_3770);
nor U5684 (N_5684,N_4332,N_4504);
nand U5685 (N_5685,N_4333,N_3604);
and U5686 (N_5686,N_4352,N_4733);
nor U5687 (N_5687,N_3993,N_4403);
and U5688 (N_5688,N_3604,N_3905);
and U5689 (N_5689,N_3673,N_4085);
xnor U5690 (N_5690,N_4269,N_4722);
nor U5691 (N_5691,N_3998,N_3985);
or U5692 (N_5692,N_4012,N_4650);
and U5693 (N_5693,N_3673,N_3747);
and U5694 (N_5694,N_4253,N_4386);
or U5695 (N_5695,N_4598,N_4436);
and U5696 (N_5696,N_4373,N_3947);
nor U5697 (N_5697,N_3624,N_3964);
xor U5698 (N_5698,N_4371,N_4667);
nor U5699 (N_5699,N_4662,N_3853);
nand U5700 (N_5700,N_4271,N_4375);
nand U5701 (N_5701,N_3674,N_4033);
nor U5702 (N_5702,N_4182,N_3724);
nand U5703 (N_5703,N_4401,N_4407);
xor U5704 (N_5704,N_3755,N_4785);
or U5705 (N_5705,N_4159,N_4278);
and U5706 (N_5706,N_4030,N_3756);
nor U5707 (N_5707,N_3649,N_4649);
or U5708 (N_5708,N_4049,N_4119);
or U5709 (N_5709,N_4412,N_4059);
and U5710 (N_5710,N_4541,N_3643);
nand U5711 (N_5711,N_4169,N_4157);
nand U5712 (N_5712,N_4394,N_4790);
or U5713 (N_5713,N_3630,N_4558);
nand U5714 (N_5714,N_3691,N_4632);
and U5715 (N_5715,N_3630,N_4422);
xor U5716 (N_5716,N_4799,N_4665);
and U5717 (N_5717,N_4701,N_4289);
nor U5718 (N_5718,N_4679,N_4412);
and U5719 (N_5719,N_4511,N_3872);
and U5720 (N_5720,N_4599,N_4472);
nor U5721 (N_5721,N_4731,N_4549);
xor U5722 (N_5722,N_4730,N_4024);
and U5723 (N_5723,N_4739,N_4656);
nor U5724 (N_5724,N_3735,N_4240);
and U5725 (N_5725,N_3730,N_3856);
or U5726 (N_5726,N_4123,N_4280);
and U5727 (N_5727,N_4080,N_4587);
xnor U5728 (N_5728,N_4152,N_3978);
nor U5729 (N_5729,N_4033,N_3851);
xor U5730 (N_5730,N_4693,N_4677);
nor U5731 (N_5731,N_4353,N_4759);
xor U5732 (N_5732,N_3618,N_3773);
nor U5733 (N_5733,N_4096,N_3972);
nor U5734 (N_5734,N_4335,N_4563);
xnor U5735 (N_5735,N_3827,N_4361);
or U5736 (N_5736,N_4247,N_3700);
xnor U5737 (N_5737,N_4364,N_3703);
or U5738 (N_5738,N_3743,N_4699);
xnor U5739 (N_5739,N_4781,N_4323);
nor U5740 (N_5740,N_4564,N_4706);
xnor U5741 (N_5741,N_4485,N_4461);
or U5742 (N_5742,N_4661,N_3772);
xor U5743 (N_5743,N_4442,N_3956);
or U5744 (N_5744,N_4265,N_4274);
nor U5745 (N_5745,N_3985,N_3622);
xnor U5746 (N_5746,N_4185,N_4182);
nor U5747 (N_5747,N_4659,N_4131);
xor U5748 (N_5748,N_4203,N_4050);
and U5749 (N_5749,N_4688,N_4542);
nor U5750 (N_5750,N_4233,N_4782);
nor U5751 (N_5751,N_4336,N_4608);
xnor U5752 (N_5752,N_3672,N_4488);
nor U5753 (N_5753,N_4107,N_4560);
nor U5754 (N_5754,N_4331,N_4485);
xor U5755 (N_5755,N_4428,N_3655);
nor U5756 (N_5756,N_4270,N_4558);
or U5757 (N_5757,N_4076,N_4089);
xnor U5758 (N_5758,N_4621,N_3736);
nand U5759 (N_5759,N_3702,N_3783);
nor U5760 (N_5760,N_4076,N_4600);
and U5761 (N_5761,N_4517,N_3960);
nor U5762 (N_5762,N_4242,N_3925);
and U5763 (N_5763,N_4477,N_4741);
or U5764 (N_5764,N_3666,N_3882);
or U5765 (N_5765,N_3694,N_4047);
and U5766 (N_5766,N_4292,N_3724);
nand U5767 (N_5767,N_3694,N_4464);
xor U5768 (N_5768,N_4676,N_4334);
nand U5769 (N_5769,N_3983,N_4660);
nand U5770 (N_5770,N_4152,N_3613);
or U5771 (N_5771,N_4198,N_4377);
and U5772 (N_5772,N_3664,N_4239);
and U5773 (N_5773,N_3941,N_4266);
xor U5774 (N_5774,N_4235,N_3684);
nand U5775 (N_5775,N_4066,N_4667);
nor U5776 (N_5776,N_4729,N_4698);
xnor U5777 (N_5777,N_4396,N_4671);
nand U5778 (N_5778,N_3601,N_4366);
and U5779 (N_5779,N_4166,N_4752);
nand U5780 (N_5780,N_4599,N_4188);
and U5781 (N_5781,N_4603,N_3784);
nor U5782 (N_5782,N_4067,N_4093);
or U5783 (N_5783,N_3812,N_3928);
or U5784 (N_5784,N_3810,N_4371);
or U5785 (N_5785,N_4607,N_4700);
nor U5786 (N_5786,N_4033,N_3607);
or U5787 (N_5787,N_3944,N_4646);
and U5788 (N_5788,N_3927,N_3769);
and U5789 (N_5789,N_4384,N_4603);
xnor U5790 (N_5790,N_4325,N_4010);
xor U5791 (N_5791,N_4160,N_4126);
xor U5792 (N_5792,N_3949,N_3641);
nor U5793 (N_5793,N_4037,N_3921);
nand U5794 (N_5794,N_4796,N_3887);
and U5795 (N_5795,N_4053,N_4507);
nand U5796 (N_5796,N_4287,N_3630);
xnor U5797 (N_5797,N_3762,N_4647);
or U5798 (N_5798,N_4613,N_3981);
xor U5799 (N_5799,N_4619,N_3906);
nand U5800 (N_5800,N_3901,N_4636);
or U5801 (N_5801,N_3715,N_3911);
nand U5802 (N_5802,N_4059,N_4002);
nand U5803 (N_5803,N_4598,N_4228);
nor U5804 (N_5804,N_4029,N_4517);
xor U5805 (N_5805,N_3609,N_4587);
and U5806 (N_5806,N_4122,N_4773);
nor U5807 (N_5807,N_4598,N_3832);
nand U5808 (N_5808,N_4298,N_3686);
xor U5809 (N_5809,N_4118,N_4408);
or U5810 (N_5810,N_4653,N_3878);
xnor U5811 (N_5811,N_4537,N_4351);
nand U5812 (N_5812,N_3792,N_4550);
or U5813 (N_5813,N_3696,N_4259);
and U5814 (N_5814,N_4053,N_4091);
xor U5815 (N_5815,N_3716,N_4139);
nand U5816 (N_5816,N_4573,N_4135);
nand U5817 (N_5817,N_4760,N_4212);
and U5818 (N_5818,N_4236,N_3822);
and U5819 (N_5819,N_4184,N_4070);
and U5820 (N_5820,N_4776,N_4674);
or U5821 (N_5821,N_4013,N_4726);
nand U5822 (N_5822,N_4650,N_3971);
nor U5823 (N_5823,N_4539,N_3981);
and U5824 (N_5824,N_4141,N_3609);
nor U5825 (N_5825,N_4726,N_4585);
and U5826 (N_5826,N_3619,N_4406);
or U5827 (N_5827,N_4339,N_4103);
nand U5828 (N_5828,N_4537,N_4112);
and U5829 (N_5829,N_4549,N_4280);
xor U5830 (N_5830,N_4217,N_3872);
and U5831 (N_5831,N_4357,N_4121);
or U5832 (N_5832,N_4592,N_4128);
and U5833 (N_5833,N_4249,N_3761);
and U5834 (N_5834,N_4321,N_3705);
nand U5835 (N_5835,N_4116,N_4505);
or U5836 (N_5836,N_3601,N_3937);
xnor U5837 (N_5837,N_3769,N_4116);
or U5838 (N_5838,N_4418,N_4302);
nand U5839 (N_5839,N_4400,N_4612);
and U5840 (N_5840,N_3632,N_4052);
or U5841 (N_5841,N_4294,N_3983);
nand U5842 (N_5842,N_4295,N_3855);
nand U5843 (N_5843,N_4185,N_4186);
and U5844 (N_5844,N_3840,N_4694);
or U5845 (N_5845,N_4723,N_4773);
xnor U5846 (N_5846,N_4412,N_4077);
nand U5847 (N_5847,N_4784,N_3600);
xor U5848 (N_5848,N_4594,N_4343);
and U5849 (N_5849,N_4434,N_4214);
nand U5850 (N_5850,N_4254,N_3807);
and U5851 (N_5851,N_4114,N_3725);
or U5852 (N_5852,N_4546,N_3856);
and U5853 (N_5853,N_4120,N_3874);
nand U5854 (N_5854,N_3627,N_4412);
and U5855 (N_5855,N_3632,N_4411);
xor U5856 (N_5856,N_4674,N_4668);
or U5857 (N_5857,N_3675,N_4265);
nor U5858 (N_5858,N_3672,N_4701);
xnor U5859 (N_5859,N_3962,N_4018);
and U5860 (N_5860,N_4060,N_3797);
nor U5861 (N_5861,N_4653,N_3792);
nand U5862 (N_5862,N_4110,N_4078);
xnor U5863 (N_5863,N_4640,N_3962);
and U5864 (N_5864,N_4597,N_4470);
or U5865 (N_5865,N_4629,N_3863);
nor U5866 (N_5866,N_4198,N_3895);
or U5867 (N_5867,N_3696,N_3659);
and U5868 (N_5868,N_4770,N_4136);
or U5869 (N_5869,N_4670,N_4783);
nand U5870 (N_5870,N_4110,N_4288);
nor U5871 (N_5871,N_4795,N_3940);
nand U5872 (N_5872,N_4660,N_3741);
nand U5873 (N_5873,N_4685,N_4185);
xnor U5874 (N_5874,N_4425,N_3679);
nand U5875 (N_5875,N_3681,N_4396);
and U5876 (N_5876,N_4571,N_3809);
or U5877 (N_5877,N_4612,N_4325);
nand U5878 (N_5878,N_4741,N_4029);
or U5879 (N_5879,N_3943,N_4705);
nand U5880 (N_5880,N_3944,N_3700);
and U5881 (N_5881,N_4758,N_4027);
nand U5882 (N_5882,N_3888,N_4349);
xor U5883 (N_5883,N_4373,N_4346);
nand U5884 (N_5884,N_4294,N_4078);
xnor U5885 (N_5885,N_4713,N_4162);
nor U5886 (N_5886,N_4136,N_4617);
nand U5887 (N_5887,N_3940,N_3694);
or U5888 (N_5888,N_4361,N_3949);
xor U5889 (N_5889,N_4686,N_4162);
or U5890 (N_5890,N_4056,N_3612);
nand U5891 (N_5891,N_4412,N_4780);
and U5892 (N_5892,N_4113,N_4144);
nand U5893 (N_5893,N_3857,N_4621);
nand U5894 (N_5894,N_4071,N_3922);
and U5895 (N_5895,N_4498,N_4367);
nor U5896 (N_5896,N_3853,N_3705);
xor U5897 (N_5897,N_3878,N_3735);
xor U5898 (N_5898,N_4236,N_4643);
nor U5899 (N_5899,N_3875,N_3920);
and U5900 (N_5900,N_4601,N_4434);
and U5901 (N_5901,N_4101,N_4173);
or U5902 (N_5902,N_4410,N_4225);
xor U5903 (N_5903,N_4666,N_3668);
or U5904 (N_5904,N_3784,N_4001);
nor U5905 (N_5905,N_4444,N_4023);
xor U5906 (N_5906,N_4791,N_4466);
nor U5907 (N_5907,N_4117,N_3954);
nand U5908 (N_5908,N_4624,N_4370);
xnor U5909 (N_5909,N_4578,N_4765);
nand U5910 (N_5910,N_4236,N_3847);
xnor U5911 (N_5911,N_4678,N_3639);
and U5912 (N_5912,N_4569,N_4249);
xor U5913 (N_5913,N_3991,N_4358);
or U5914 (N_5914,N_3961,N_4470);
or U5915 (N_5915,N_4476,N_4749);
nor U5916 (N_5916,N_3617,N_3972);
nand U5917 (N_5917,N_4580,N_4257);
nand U5918 (N_5918,N_4775,N_4252);
nand U5919 (N_5919,N_4286,N_4798);
nor U5920 (N_5920,N_4474,N_4112);
or U5921 (N_5921,N_4680,N_4023);
nor U5922 (N_5922,N_3623,N_4238);
and U5923 (N_5923,N_4088,N_3692);
xnor U5924 (N_5924,N_3826,N_4077);
and U5925 (N_5925,N_4279,N_4675);
and U5926 (N_5926,N_4410,N_4392);
nor U5927 (N_5927,N_3698,N_3855);
or U5928 (N_5928,N_3962,N_4328);
or U5929 (N_5929,N_3809,N_4648);
and U5930 (N_5930,N_3765,N_3728);
and U5931 (N_5931,N_3847,N_4592);
nor U5932 (N_5932,N_4347,N_4719);
or U5933 (N_5933,N_4228,N_4245);
or U5934 (N_5934,N_4351,N_4155);
or U5935 (N_5935,N_4765,N_4767);
or U5936 (N_5936,N_3654,N_4065);
and U5937 (N_5937,N_4727,N_3944);
or U5938 (N_5938,N_4755,N_4323);
nand U5939 (N_5939,N_4381,N_3934);
nand U5940 (N_5940,N_3624,N_4783);
and U5941 (N_5941,N_3949,N_4788);
nor U5942 (N_5942,N_3864,N_4238);
and U5943 (N_5943,N_4246,N_4504);
and U5944 (N_5944,N_4049,N_4339);
nand U5945 (N_5945,N_3650,N_3915);
nand U5946 (N_5946,N_3655,N_3989);
and U5947 (N_5947,N_4357,N_4370);
xor U5948 (N_5948,N_3733,N_4728);
and U5949 (N_5949,N_4587,N_4600);
nor U5950 (N_5950,N_4239,N_3947);
nor U5951 (N_5951,N_4517,N_3894);
nor U5952 (N_5952,N_4756,N_3706);
xnor U5953 (N_5953,N_4130,N_4558);
and U5954 (N_5954,N_3769,N_3741);
nand U5955 (N_5955,N_4791,N_3965);
and U5956 (N_5956,N_3942,N_4547);
and U5957 (N_5957,N_4273,N_4527);
or U5958 (N_5958,N_3776,N_4594);
nand U5959 (N_5959,N_4088,N_4068);
or U5960 (N_5960,N_4260,N_4529);
and U5961 (N_5961,N_3918,N_4390);
xor U5962 (N_5962,N_4558,N_3642);
xnor U5963 (N_5963,N_4237,N_4621);
xnor U5964 (N_5964,N_3729,N_4348);
nor U5965 (N_5965,N_3865,N_3911);
nand U5966 (N_5966,N_3822,N_4469);
and U5967 (N_5967,N_3974,N_3690);
or U5968 (N_5968,N_4650,N_4523);
nor U5969 (N_5969,N_4314,N_3667);
xor U5970 (N_5970,N_3935,N_3603);
and U5971 (N_5971,N_3631,N_4723);
xnor U5972 (N_5972,N_4773,N_4178);
and U5973 (N_5973,N_4581,N_4382);
xor U5974 (N_5974,N_4099,N_4756);
xor U5975 (N_5975,N_4008,N_4473);
and U5976 (N_5976,N_3734,N_4644);
nand U5977 (N_5977,N_4291,N_4704);
and U5978 (N_5978,N_4465,N_3908);
nand U5979 (N_5979,N_4140,N_4161);
or U5980 (N_5980,N_4587,N_4405);
xnor U5981 (N_5981,N_4722,N_4420);
nand U5982 (N_5982,N_4563,N_4579);
or U5983 (N_5983,N_4344,N_4607);
nand U5984 (N_5984,N_4363,N_4521);
and U5985 (N_5985,N_3711,N_4240);
nor U5986 (N_5986,N_4576,N_4400);
xnor U5987 (N_5987,N_3700,N_3992);
nand U5988 (N_5988,N_4289,N_4039);
xnor U5989 (N_5989,N_3935,N_3747);
or U5990 (N_5990,N_4537,N_4600);
or U5991 (N_5991,N_3904,N_4204);
and U5992 (N_5992,N_4142,N_4271);
xnor U5993 (N_5993,N_4000,N_3748);
nor U5994 (N_5994,N_4234,N_4265);
xnor U5995 (N_5995,N_4601,N_3855);
xnor U5996 (N_5996,N_4292,N_3800);
or U5997 (N_5997,N_4625,N_3929);
nand U5998 (N_5998,N_4630,N_4545);
nor U5999 (N_5999,N_3621,N_4476);
xnor U6000 (N_6000,N_4829,N_5457);
xnor U6001 (N_6001,N_5669,N_5445);
and U6002 (N_6002,N_5082,N_5160);
xnor U6003 (N_6003,N_5990,N_5043);
or U6004 (N_6004,N_5092,N_5866);
and U6005 (N_6005,N_5026,N_5788);
nor U6006 (N_6006,N_5109,N_5491);
and U6007 (N_6007,N_5860,N_5139);
nand U6008 (N_6008,N_5101,N_4849);
or U6009 (N_6009,N_5507,N_5071);
nand U6010 (N_6010,N_5471,N_5784);
or U6011 (N_6011,N_5137,N_5544);
xnor U6012 (N_6012,N_4900,N_5059);
xnor U6013 (N_6013,N_5234,N_5476);
nand U6014 (N_6014,N_5005,N_5487);
nor U6015 (N_6015,N_5126,N_5453);
nand U6016 (N_6016,N_5115,N_5244);
or U6017 (N_6017,N_5642,N_5470);
nor U6018 (N_6018,N_5818,N_5930);
nor U6019 (N_6019,N_5756,N_5655);
nor U6020 (N_6020,N_5151,N_5316);
nor U6021 (N_6021,N_5980,N_5436);
xnor U6022 (N_6022,N_5339,N_5834);
nand U6023 (N_6023,N_5743,N_5430);
or U6024 (N_6024,N_5185,N_5789);
xor U6025 (N_6025,N_5850,N_5737);
and U6026 (N_6026,N_5810,N_5439);
or U6027 (N_6027,N_5712,N_5839);
xnor U6028 (N_6028,N_5581,N_5978);
or U6029 (N_6029,N_5179,N_4891);
or U6030 (N_6030,N_5719,N_5191);
or U6031 (N_6031,N_5227,N_4979);
nor U6032 (N_6032,N_5266,N_5338);
nand U6033 (N_6033,N_5862,N_5557);
nor U6034 (N_6034,N_4922,N_5845);
or U6035 (N_6035,N_5093,N_5194);
nand U6036 (N_6036,N_5697,N_5699);
nand U6037 (N_6037,N_5490,N_5406);
and U6038 (N_6038,N_4805,N_5542);
nor U6039 (N_6039,N_5007,N_5364);
and U6040 (N_6040,N_5943,N_4882);
nand U6041 (N_6041,N_4934,N_5666);
or U6042 (N_6042,N_4892,N_5183);
nand U6043 (N_6043,N_4890,N_5523);
xnor U6044 (N_6044,N_5518,N_4959);
nor U6045 (N_6045,N_5963,N_4843);
nor U6046 (N_6046,N_5590,N_4901);
nor U6047 (N_6047,N_5512,N_5762);
xnor U6048 (N_6048,N_5887,N_5799);
or U6049 (N_6049,N_5173,N_5934);
or U6050 (N_6050,N_5131,N_5177);
or U6051 (N_6051,N_5468,N_5334);
and U6052 (N_6052,N_4984,N_5552);
nand U6053 (N_6053,N_5260,N_5998);
nor U6054 (N_6054,N_5226,N_5246);
nand U6055 (N_6055,N_5418,N_4937);
and U6056 (N_6056,N_5972,N_5107);
nor U6057 (N_6057,N_5665,N_5002);
nand U6058 (N_6058,N_5813,N_5910);
nand U6059 (N_6059,N_5938,N_5739);
nor U6060 (N_6060,N_5052,N_5335);
nand U6061 (N_6061,N_5601,N_5920);
nand U6062 (N_6062,N_5715,N_5859);
and U6063 (N_6063,N_4884,N_5248);
xor U6064 (N_6064,N_5794,N_5089);
and U6065 (N_6065,N_5599,N_5357);
nor U6066 (N_6066,N_5394,N_5024);
xor U6067 (N_6067,N_5270,N_5027);
and U6068 (N_6068,N_4951,N_5767);
or U6069 (N_6069,N_4991,N_4939);
xnor U6070 (N_6070,N_4813,N_4879);
nor U6071 (N_6071,N_5911,N_5856);
xor U6072 (N_6072,N_5158,N_5279);
and U6073 (N_6073,N_5233,N_5661);
nand U6074 (N_6074,N_5130,N_5128);
or U6075 (N_6075,N_5019,N_5050);
xnor U6076 (N_6076,N_4822,N_4970);
or U6077 (N_6077,N_5505,N_4842);
xnor U6078 (N_6078,N_5514,N_5317);
or U6079 (N_6079,N_5210,N_5770);
or U6080 (N_6080,N_5628,N_5957);
and U6081 (N_6081,N_5959,N_5632);
nand U6082 (N_6082,N_4883,N_5048);
xor U6083 (N_6083,N_5129,N_5981);
nand U6084 (N_6084,N_4885,N_5302);
or U6085 (N_6085,N_5055,N_4982);
xnor U6086 (N_6086,N_5051,N_5180);
or U6087 (N_6087,N_5517,N_4854);
nand U6088 (N_6088,N_4973,N_5836);
nor U6089 (N_6089,N_5045,N_5888);
nor U6090 (N_6090,N_4875,N_5230);
or U6091 (N_6091,N_4841,N_5873);
nand U6092 (N_6092,N_5408,N_4916);
and U6093 (N_6093,N_5782,N_5295);
nand U6094 (N_6094,N_5752,N_4861);
and U6095 (N_6095,N_5977,N_5448);
nand U6096 (N_6096,N_5387,N_4920);
and U6097 (N_6097,N_5150,N_4932);
xnor U6098 (N_6098,N_4802,N_5650);
xnor U6099 (N_6099,N_5738,N_5554);
xnor U6100 (N_6100,N_5876,N_5474);
or U6101 (N_6101,N_5263,N_5001);
nor U6102 (N_6102,N_5704,N_5508);
and U6103 (N_6103,N_5111,N_5361);
or U6104 (N_6104,N_5616,N_5730);
nor U6105 (N_6105,N_5192,N_4889);
and U6106 (N_6106,N_4943,N_5626);
and U6107 (N_6107,N_5708,N_5344);
xor U6108 (N_6108,N_5087,N_5374);
or U6109 (N_6109,N_5440,N_5740);
or U6110 (N_6110,N_5631,N_5922);
and U6111 (N_6111,N_5187,N_5985);
xnor U6112 (N_6112,N_5056,N_5321);
nand U6113 (N_6113,N_5376,N_5011);
or U6114 (N_6114,N_4872,N_5127);
or U6115 (N_6115,N_5821,N_5975);
xnor U6116 (N_6116,N_5256,N_5225);
xnor U6117 (N_6117,N_4828,N_5264);
or U6118 (N_6118,N_5433,N_5996);
nand U6119 (N_6119,N_5566,N_5675);
xnor U6120 (N_6120,N_5221,N_5349);
xor U6121 (N_6121,N_4995,N_4993);
nand U6122 (N_6122,N_5777,N_5638);
nor U6123 (N_6123,N_5067,N_4927);
and U6124 (N_6124,N_4856,N_5379);
nand U6125 (N_6125,N_4940,N_5322);
nand U6126 (N_6126,N_4800,N_5199);
nand U6127 (N_6127,N_5574,N_5742);
xor U6128 (N_6128,N_5319,N_5858);
and U6129 (N_6129,N_5423,N_5345);
or U6130 (N_6130,N_5694,N_5117);
nor U6131 (N_6131,N_5133,N_5359);
nand U6132 (N_6132,N_5294,N_5905);
and U6133 (N_6133,N_5034,N_5835);
and U6134 (N_6134,N_5659,N_5299);
or U6135 (N_6135,N_5409,N_5968);
nand U6136 (N_6136,N_5872,N_5202);
xnor U6137 (N_6137,N_5157,N_5152);
and U6138 (N_6138,N_4899,N_5410);
and U6139 (N_6139,N_5711,N_5598);
nand U6140 (N_6140,N_5278,N_5275);
xor U6141 (N_6141,N_5184,N_5933);
and U6142 (N_6142,N_5114,N_5413);
and U6143 (N_6143,N_5731,N_5994);
and U6144 (N_6144,N_5912,N_5219);
and U6145 (N_6145,N_4838,N_5309);
nand U6146 (N_6146,N_5627,N_5962);
xnor U6147 (N_6147,N_5506,N_5870);
nor U6148 (N_6148,N_5106,N_5944);
xnor U6149 (N_6149,N_5605,N_5691);
xnor U6150 (N_6150,N_5645,N_5393);
xnor U6151 (N_6151,N_5923,N_4873);
and U6152 (N_6152,N_5511,N_5563);
nand U6153 (N_6153,N_5161,N_4862);
and U6154 (N_6154,N_5012,N_5608);
or U6155 (N_6155,N_5330,N_5559);
and U6156 (N_6156,N_5496,N_4834);
nand U6157 (N_6157,N_5090,N_5113);
xor U6158 (N_6158,N_5656,N_5485);
nor U6159 (N_6159,N_5315,N_5431);
xnor U6160 (N_6160,N_5956,N_5172);
or U6161 (N_6161,N_5076,N_5372);
xor U6162 (N_6162,N_5000,N_5255);
nand U6163 (N_6163,N_5355,N_5806);
nand U6164 (N_6164,N_5567,N_5824);
or U6165 (N_6165,N_4987,N_5197);
nor U6166 (N_6166,N_4887,N_5607);
nand U6167 (N_6167,N_5816,N_5419);
nand U6168 (N_6168,N_4961,N_5366);
nand U6169 (N_6169,N_5036,N_5736);
nor U6170 (N_6170,N_5991,N_5018);
or U6171 (N_6171,N_5216,N_5884);
xnor U6172 (N_6172,N_4923,N_5369);
or U6173 (N_6173,N_5936,N_4860);
nand U6174 (N_6174,N_5982,N_5683);
and U6175 (N_6175,N_5979,N_5630);
or U6176 (N_6176,N_5099,N_5283);
nand U6177 (N_6177,N_5206,N_4953);
and U6178 (N_6178,N_5946,N_5636);
and U6179 (N_6179,N_5288,N_5973);
or U6180 (N_6180,N_5437,N_5205);
and U6181 (N_6181,N_5717,N_5597);
nand U6182 (N_6182,N_5997,N_5083);
and U6183 (N_6183,N_5392,N_5553);
and U6184 (N_6184,N_5571,N_5162);
and U6185 (N_6185,N_5837,N_5175);
or U6186 (N_6186,N_5240,N_5261);
or U6187 (N_6187,N_5336,N_5809);
nor U6188 (N_6188,N_5065,N_5267);
and U6189 (N_6189,N_5579,N_5624);
nor U6190 (N_6190,N_5776,N_5017);
or U6191 (N_6191,N_5706,N_5931);
or U6192 (N_6192,N_5612,N_5618);
nor U6193 (N_6193,N_5639,N_5588);
and U6194 (N_6194,N_5760,N_5124);
and U6195 (N_6195,N_5108,N_4977);
or U6196 (N_6196,N_5353,N_5976);
or U6197 (N_6197,N_5098,N_5967);
and U6198 (N_6198,N_5966,N_5477);
nor U6199 (N_6199,N_5575,N_4853);
nand U6200 (N_6200,N_5852,N_5144);
or U6201 (N_6201,N_5003,N_5692);
or U6202 (N_6202,N_4929,N_5503);
or U6203 (N_6203,N_5684,N_5781);
nor U6204 (N_6204,N_4878,N_5495);
xnor U6205 (N_6205,N_5759,N_5053);
nor U6206 (N_6206,N_5054,N_5497);
or U6207 (N_6207,N_5291,N_5218);
nand U6208 (N_6208,N_5698,N_5057);
xor U6209 (N_6209,N_4810,N_5695);
or U6210 (N_6210,N_5132,N_5796);
and U6211 (N_6211,N_5220,N_5049);
and U6212 (N_6212,N_5569,N_5595);
and U6213 (N_6213,N_5902,N_4972);
nand U6214 (N_6214,N_4909,N_5347);
nand U6215 (N_6215,N_5259,N_4832);
nor U6216 (N_6216,N_4988,N_5727);
xor U6217 (N_6217,N_5363,N_5449);
xnor U6218 (N_6218,N_5306,N_5536);
nor U6219 (N_6219,N_5416,N_5594);
or U6220 (N_6220,N_5383,N_5207);
xor U6221 (N_6221,N_5360,N_5892);
or U6222 (N_6222,N_5296,N_5060);
or U6223 (N_6223,N_5398,N_5530);
xnor U6224 (N_6224,N_5793,N_5549);
or U6225 (N_6225,N_5326,N_5375);
xnor U6226 (N_6226,N_4921,N_4888);
or U6227 (N_6227,N_5480,N_5258);
and U6228 (N_6228,N_5718,N_5949);
and U6229 (N_6229,N_5961,N_4985);
nor U6230 (N_6230,N_4954,N_5100);
xnor U6231 (N_6231,N_5720,N_5587);
xnor U6232 (N_6232,N_5894,N_5085);
nor U6233 (N_6233,N_5928,N_5526);
and U6234 (N_6234,N_5352,N_5800);
nor U6235 (N_6235,N_5122,N_5310);
or U6236 (N_6236,N_5772,N_4946);
or U6237 (N_6237,N_5041,N_5547);
xor U6238 (N_6238,N_5728,N_5138);
and U6239 (N_6239,N_5560,N_4836);
nor U6240 (N_6240,N_5438,N_5676);
xnor U6241 (N_6241,N_5614,N_5522);
xor U6242 (N_6242,N_5329,N_4983);
or U6243 (N_6243,N_5754,N_5913);
nor U6244 (N_6244,N_5572,N_4812);
nand U6245 (N_6245,N_5271,N_5539);
or U6246 (N_6246,N_5851,N_5297);
and U6247 (N_6247,N_5368,N_4804);
nor U6248 (N_6248,N_5120,N_5582);
nor U6249 (N_6249,N_5942,N_5779);
or U6250 (N_6250,N_5400,N_4801);
or U6251 (N_6251,N_4969,N_5390);
xor U6252 (N_6252,N_5145,N_5103);
nand U6253 (N_6253,N_5509,N_5686);
nand U6254 (N_6254,N_5236,N_5479);
and U6255 (N_6255,N_5212,N_5386);
or U6256 (N_6256,N_5875,N_5945);
or U6257 (N_6257,N_4928,N_5646);
nand U6258 (N_6258,N_4844,N_5868);
nor U6259 (N_6259,N_5484,N_4980);
or U6260 (N_6260,N_5110,N_4994);
nand U6261 (N_6261,N_5716,N_5825);
nand U6262 (N_6262,N_5679,N_4935);
and U6263 (N_6263,N_5622,N_5010);
nand U6264 (N_6264,N_5774,N_5685);
xnor U6265 (N_6265,N_5841,N_5343);
or U6266 (N_6266,N_4847,N_4868);
nand U6267 (N_6267,N_5424,N_5381);
nor U6268 (N_6268,N_5252,N_5970);
nand U6269 (N_6269,N_4926,N_5351);
nor U6270 (N_6270,N_5472,N_5066);
or U6271 (N_6271,N_5008,N_4914);
nor U6272 (N_6272,N_5042,N_5091);
or U6273 (N_6273,N_5488,N_5080);
and U6274 (N_6274,N_5570,N_4948);
xnor U6275 (N_6275,N_5033,N_5916);
and U6276 (N_6276,N_5254,N_5667);
nor U6277 (N_6277,N_5611,N_5354);
xor U6278 (N_6278,N_5148,N_5021);
and U6279 (N_6279,N_5181,N_4908);
and U6280 (N_6280,N_5358,N_5853);
or U6281 (N_6281,N_5702,N_5443);
xnor U6282 (N_6282,N_5886,N_5890);
nand U6283 (N_6283,N_5044,N_5201);
and U6284 (N_6284,N_5251,N_5528);
or U6285 (N_6285,N_5953,N_5584);
and U6286 (N_6286,N_5540,N_5425);
nor U6287 (N_6287,N_5014,N_5846);
and U6288 (N_6288,N_5874,N_5703);
nand U6289 (N_6289,N_5901,N_5281);
or U6290 (N_6290,N_5169,N_4852);
nor U6291 (N_6291,N_5290,N_5174);
or U6292 (N_6292,N_5932,N_5140);
or U6293 (N_6293,N_4894,N_5899);
xnor U6294 (N_6294,N_5245,N_4941);
or U6295 (N_6295,N_5812,N_4896);
nand U6296 (N_6296,N_5974,N_5591);
nand U6297 (N_6297,N_5242,N_5228);
nor U6298 (N_6298,N_5341,N_5696);
or U6299 (N_6299,N_5214,N_5926);
and U6300 (N_6300,N_4997,N_4819);
nor U6301 (N_6301,N_5434,N_5647);
xnor U6302 (N_6302,N_5829,N_5069);
nor U6303 (N_6303,N_5941,N_5746);
nor U6304 (N_6304,N_5558,N_4867);
xnor U6305 (N_6305,N_5342,N_4895);
nor U6306 (N_6306,N_5785,N_5195);
and U6307 (N_6307,N_5532,N_5960);
nand U6308 (N_6308,N_5613,N_5664);
or U6309 (N_6309,N_5826,N_5143);
nand U6310 (N_6310,N_5898,N_4814);
nand U6311 (N_6311,N_5965,N_5486);
nand U6312 (N_6312,N_5401,N_5726);
and U6313 (N_6313,N_5079,N_5925);
and U6314 (N_6314,N_5156,N_5885);
or U6315 (N_6315,N_5802,N_4958);
and U6316 (N_6316,N_5896,N_4947);
nor U6317 (N_6317,N_5586,N_5602);
xnor U6318 (N_6318,N_5748,N_5914);
or U6319 (N_6319,N_4839,N_5993);
nand U6320 (N_6320,N_5257,N_5768);
or U6321 (N_6321,N_5819,N_4996);
xnor U6322 (N_6322,N_4857,N_4963);
xnor U6323 (N_6323,N_5682,N_4866);
xor U6324 (N_6324,N_5805,N_5546);
nor U6325 (N_6325,N_5543,N_5389);
or U6326 (N_6326,N_5047,N_5678);
and U6327 (N_6327,N_5955,N_5037);
or U6328 (N_6328,N_5680,N_5016);
xnor U6329 (N_6329,N_5272,N_5116);
nor U6330 (N_6330,N_5830,N_5331);
and U6331 (N_6331,N_4924,N_5814);
and U6332 (N_6332,N_4952,N_5168);
nor U6333 (N_6333,N_5243,N_5154);
and U6334 (N_6334,N_4803,N_5637);
nor U6335 (N_6335,N_5435,N_5633);
nor U6336 (N_6336,N_5446,N_5280);
or U6337 (N_6337,N_5833,N_5723);
and U6338 (N_6338,N_5455,N_5915);
or U6339 (N_6339,N_5753,N_5939);
and U6340 (N_6340,N_5112,N_4905);
xor U6341 (N_6341,N_4848,N_5421);
nor U6342 (N_6342,N_4807,N_5502);
or U6343 (N_6343,N_5384,N_4874);
or U6344 (N_6344,N_5373,N_5534);
or U6345 (N_6345,N_5820,N_5783);
and U6346 (N_6346,N_5786,N_5780);
nand U6347 (N_6347,N_4975,N_4815);
xor U6348 (N_6348,N_5015,N_5889);
nand U6349 (N_6349,N_5849,N_5881);
or U6350 (N_6350,N_5769,N_5170);
nor U6351 (N_6351,N_5578,N_4998);
or U6352 (N_6352,N_5635,N_5167);
and U6353 (N_6353,N_4817,N_4960);
nand U6354 (N_6354,N_5013,N_5987);
nand U6355 (N_6355,N_5958,N_5396);
xnor U6356 (N_6356,N_5346,N_5188);
and U6357 (N_6357,N_5119,N_5104);
and U6358 (N_6358,N_4816,N_5348);
xor U6359 (N_6359,N_5077,N_5573);
xnor U6360 (N_6360,N_5735,N_5734);
nor U6361 (N_6361,N_5466,N_5451);
nor U6362 (N_6362,N_5478,N_5074);
xor U6363 (N_6363,N_4913,N_4911);
or U6364 (N_6364,N_5758,N_5600);
xor U6365 (N_6365,N_4904,N_5771);
or U6366 (N_6366,N_4859,N_5062);
nand U6367 (N_6367,N_4881,N_4818);
nand U6368 (N_6368,N_5551,N_5473);
or U6369 (N_6369,N_5422,N_4965);
and U6370 (N_6370,N_5285,N_4806);
xnor U6371 (N_6371,N_5235,N_5414);
or U6372 (N_6372,N_5857,N_5654);
and U6373 (N_6373,N_5411,N_5328);
and U6374 (N_6374,N_5653,N_5415);
and U6375 (N_6375,N_5378,N_5273);
nand U6376 (N_6376,N_4902,N_5159);
or U6377 (N_6377,N_5847,N_5840);
nor U6378 (N_6378,N_5969,N_5995);
and U6379 (N_6379,N_5456,N_5677);
nor U6380 (N_6380,N_4863,N_5237);
nand U6381 (N_6381,N_5795,N_4825);
and U6382 (N_6382,N_5039,N_5662);
xor U6383 (N_6383,N_5284,N_5950);
nand U6384 (N_6384,N_5729,N_5524);
nand U6385 (N_6385,N_5332,N_4925);
nor U6386 (N_6386,N_5229,N_5417);
or U6387 (N_6387,N_5450,N_4876);
and U6388 (N_6388,N_5651,N_5311);
xor U6389 (N_6389,N_5407,N_4976);
nand U6390 (N_6390,N_5196,N_5954);
or U6391 (N_6391,N_5861,N_5725);
nand U6392 (N_6392,N_5030,N_5623);
and U6393 (N_6393,N_5462,N_5211);
and U6394 (N_6394,N_5467,N_5118);
nand U6395 (N_6395,N_5094,N_4831);
xor U6396 (N_6396,N_4912,N_5215);
nor U6397 (N_6397,N_5828,N_5903);
and U6398 (N_6398,N_5864,N_5458);
and U6399 (N_6399,N_5701,N_5672);
or U6400 (N_6400,N_5525,N_4981);
or U6401 (N_6401,N_4989,N_5070);
nand U6402 (N_6402,N_5464,N_5232);
xnor U6403 (N_6403,N_5848,N_5146);
or U6404 (N_6404,N_4962,N_5031);
or U6405 (N_6405,N_5634,N_4938);
and U6406 (N_6406,N_5312,N_5541);
xor U6407 (N_6407,N_4910,N_5420);
xnor U6408 (N_6408,N_5935,N_5135);
and U6409 (N_6409,N_5564,N_5444);
nor U6410 (N_6410,N_5673,N_5465);
or U6411 (N_6411,N_5804,N_4871);
nand U6412 (N_6412,N_5163,N_5081);
or U6413 (N_6413,N_5555,N_5585);
or U6414 (N_6414,N_4903,N_5308);
or U6415 (N_6415,N_5609,N_5548);
and U6416 (N_6416,N_4830,N_4897);
nor U6417 (N_6417,N_5035,N_5519);
nor U6418 (N_6418,N_5871,N_5298);
nand U6419 (N_6419,N_5492,N_5324);
and U6420 (N_6420,N_5088,N_5660);
xnor U6421 (N_6421,N_5391,N_5463);
xnor U6422 (N_6422,N_5893,N_4811);
and U6423 (N_6423,N_5538,N_5741);
or U6424 (N_6424,N_5900,N_5693);
and U6425 (N_6425,N_5262,N_5992);
nand U6426 (N_6426,N_5937,N_5501);
or U6427 (N_6427,N_5644,N_5277);
or U6428 (N_6428,N_5520,N_5527);
nor U6429 (N_6429,N_5763,N_5086);
and U6430 (N_6430,N_5589,N_4950);
and U6431 (N_6431,N_5649,N_5687);
or U6432 (N_6432,N_5178,N_5757);
and U6433 (N_6433,N_5878,N_5801);
nor U6434 (N_6434,N_5493,N_5986);
xor U6435 (N_6435,N_5287,N_5200);
and U6436 (N_6436,N_5454,N_4850);
or U6437 (N_6437,N_5412,N_5854);
and U6438 (N_6438,N_5040,N_5038);
or U6439 (N_6439,N_4949,N_5617);
xor U6440 (N_6440,N_5136,N_5190);
xnor U6441 (N_6441,N_5948,N_5580);
xnor U6442 (N_6442,N_5253,N_4846);
nand U6443 (N_6443,N_5141,N_5545);
nand U6444 (N_6444,N_5790,N_5556);
and U6445 (N_6445,N_4840,N_5095);
xnor U6446 (N_6446,N_5583,N_4865);
xor U6447 (N_6447,N_4855,N_4893);
or U6448 (N_6448,N_5604,N_5025);
nor U6449 (N_6449,N_5984,N_5531);
nor U6450 (N_6450,N_5658,N_5313);
or U6451 (N_6451,N_5907,N_5293);
nand U6452 (N_6452,N_5286,N_4942);
nand U6453 (N_6453,N_5380,N_5149);
nor U6454 (N_6454,N_5766,N_5964);
nand U6455 (N_6455,N_5489,N_5515);
or U6456 (N_6456,N_5791,N_5231);
nand U6457 (N_6457,N_5362,N_5831);
nand U6458 (N_6458,N_5305,N_4864);
nand U6459 (N_6459,N_5189,N_5606);
nor U6460 (N_6460,N_5365,N_5072);
nor U6461 (N_6461,N_5822,N_5869);
xor U6462 (N_6462,N_5787,N_5193);
nor U6463 (N_6463,N_4826,N_5504);
xnor U6464 (N_6464,N_5843,N_5006);
nor U6465 (N_6465,N_5009,N_5500);
nand U6466 (N_6466,N_5426,N_5301);
xor U6467 (N_6467,N_5577,N_5842);
nor U6468 (N_6468,N_5880,N_5867);
and U6469 (N_6469,N_5482,N_4821);
or U6470 (N_6470,N_5182,N_5102);
nor U6471 (N_6471,N_5674,N_5610);
or U6472 (N_6472,N_5705,N_4971);
xor U6473 (N_6473,N_5565,N_5904);
nor U6474 (N_6474,N_4820,N_5710);
nand U6475 (N_6475,N_5276,N_5882);
nand U6476 (N_6476,N_5153,N_5300);
nand U6477 (N_6477,N_5778,N_5370);
or U6478 (N_6478,N_5971,N_5798);
and U6479 (N_6479,N_5883,N_5803);
and U6480 (N_6480,N_5908,N_5224);
and U6481 (N_6481,N_5459,N_5303);
xnor U6482 (N_6482,N_5832,N_5596);
nor U6483 (N_6483,N_5247,N_5707);
or U6484 (N_6484,N_5811,N_5382);
and U6485 (N_6485,N_5924,N_5371);
or U6486 (N_6486,N_5629,N_4886);
or U6487 (N_6487,N_5744,N_5921);
and U6488 (N_6488,N_5562,N_5125);
nand U6489 (N_6489,N_5340,N_5063);
xor U6490 (N_6490,N_4833,N_5621);
nand U6491 (N_6491,N_4992,N_5643);
xnor U6492 (N_6492,N_5709,N_5250);
nand U6493 (N_6493,N_5732,N_4931);
nand U6494 (N_6494,N_5947,N_5134);
and U6495 (N_6495,N_5314,N_4880);
xor U6496 (N_6496,N_4870,N_4898);
nor U6497 (N_6497,N_5249,N_4845);
xor U6498 (N_6498,N_4907,N_5681);
nor U6499 (N_6499,N_5377,N_5004);
nand U6500 (N_6500,N_5198,N_4955);
and U6501 (N_6501,N_5405,N_4957);
or U6502 (N_6502,N_5499,N_4930);
nand U6503 (N_6503,N_4936,N_5879);
and U6504 (N_6504,N_5469,N_5483);
nand U6505 (N_6505,N_5356,N_5652);
and U6506 (N_6506,N_5282,N_5640);
nand U6507 (N_6507,N_5663,N_5657);
and U6508 (N_6508,N_4915,N_5747);
xnor U6509 (N_6509,N_4823,N_5176);
xor U6510 (N_6510,N_4986,N_5203);
nor U6511 (N_6511,N_5751,N_4917);
or U6512 (N_6512,N_5529,N_5029);
nand U6513 (N_6513,N_5268,N_5121);
xor U6514 (N_6514,N_5615,N_5952);
xnor U6515 (N_6515,N_5807,N_5078);
or U6516 (N_6516,N_5917,N_4824);
and U6517 (N_6517,N_5940,N_5020);
nand U6518 (N_6518,N_4809,N_4906);
and U6519 (N_6519,N_5427,N_5327);
nor U6520 (N_6520,N_5442,N_5533);
and U6521 (N_6521,N_5603,N_5481);
and U6522 (N_6522,N_5028,N_5714);
xor U6523 (N_6523,N_5724,N_5690);
nand U6524 (N_6524,N_5620,N_5929);
nand U6525 (N_6525,N_5775,N_5441);
and U6526 (N_6526,N_5988,N_5337);
xor U6527 (N_6527,N_5641,N_4945);
xnor U6528 (N_6528,N_5265,N_4851);
nor U6529 (N_6529,N_5274,N_5918);
nor U6530 (N_6530,N_4858,N_5648);
or U6531 (N_6531,N_5863,N_5576);
nor U6532 (N_6532,N_5307,N_5333);
nor U6533 (N_6533,N_5289,N_4956);
and U6534 (N_6534,N_5494,N_5999);
nand U6535 (N_6535,N_5909,N_5164);
or U6536 (N_6536,N_5452,N_5619);
xnor U6537 (N_6537,N_5395,N_5550);
nand U6538 (N_6538,N_5064,N_4974);
xor U6539 (N_6539,N_5510,N_5765);
nand U6540 (N_6540,N_5292,N_5032);
or U6541 (N_6541,N_4918,N_5171);
xor U6542 (N_6542,N_5325,N_5222);
nor U6543 (N_6543,N_4967,N_5213);
xor U6544 (N_6544,N_5022,N_5061);
nor U6545 (N_6545,N_5068,N_5058);
or U6546 (N_6546,N_4990,N_5891);
or U6547 (N_6547,N_4877,N_5204);
or U6548 (N_6548,N_4999,N_5537);
nand U6549 (N_6549,N_5568,N_5593);
nor U6550 (N_6550,N_5142,N_4944);
xnor U6551 (N_6551,N_5865,N_4919);
and U6552 (N_6552,N_4968,N_5105);
nand U6553 (N_6553,N_4964,N_5223);
nand U6554 (N_6554,N_5761,N_4835);
nand U6555 (N_6555,N_5084,N_5241);
or U6556 (N_6556,N_5817,N_5764);
nand U6557 (N_6557,N_5208,N_5983);
nand U6558 (N_6558,N_5855,N_4837);
nand U6559 (N_6559,N_4808,N_5075);
and U6560 (N_6560,N_5096,N_5919);
xor U6561 (N_6561,N_5733,N_5388);
nand U6562 (N_6562,N_5447,N_5792);
and U6563 (N_6563,N_5320,N_5023);
nor U6564 (N_6564,N_5429,N_5186);
nor U6565 (N_6565,N_5670,N_5808);
nand U6566 (N_6566,N_5165,N_5521);
nand U6567 (N_6567,N_5385,N_5046);
or U6568 (N_6568,N_5797,N_5155);
xnor U6569 (N_6569,N_5749,N_5906);
nor U6570 (N_6570,N_5097,N_4827);
xnor U6571 (N_6571,N_5498,N_4869);
nor U6572 (N_6572,N_5689,N_5951);
and U6573 (N_6573,N_5460,N_5461);
or U6574 (N_6574,N_5668,N_4966);
nor U6575 (N_6575,N_5123,N_5318);
nand U6576 (N_6576,N_5403,N_5989);
or U6577 (N_6577,N_5671,N_5721);
nand U6578 (N_6578,N_5073,N_5688);
xor U6579 (N_6579,N_5844,N_5823);
or U6580 (N_6580,N_5239,N_5209);
and U6581 (N_6581,N_5269,N_5238);
xnor U6582 (N_6582,N_4978,N_5404);
nor U6583 (N_6583,N_5535,N_5304);
xor U6584 (N_6584,N_5399,N_5750);
or U6585 (N_6585,N_5217,N_5722);
nand U6586 (N_6586,N_5516,N_5428);
or U6587 (N_6587,N_5350,N_5745);
nor U6588 (N_6588,N_5561,N_5895);
or U6589 (N_6589,N_5713,N_5397);
nor U6590 (N_6590,N_5838,N_5367);
nand U6591 (N_6591,N_5475,N_5773);
and U6592 (N_6592,N_5147,N_5927);
xnor U6593 (N_6593,N_5513,N_5432);
nand U6594 (N_6594,N_5625,N_5815);
and U6595 (N_6595,N_5700,N_5592);
nor U6596 (N_6596,N_5897,N_5402);
or U6597 (N_6597,N_5755,N_4933);
and U6598 (N_6598,N_5166,N_5877);
and U6599 (N_6599,N_5827,N_5323);
nand U6600 (N_6600,N_5285,N_5274);
nand U6601 (N_6601,N_5415,N_5381);
or U6602 (N_6602,N_5262,N_5134);
or U6603 (N_6603,N_5952,N_5796);
nand U6604 (N_6604,N_5412,N_5677);
nor U6605 (N_6605,N_4833,N_5702);
xnor U6606 (N_6606,N_5440,N_5983);
nor U6607 (N_6607,N_4836,N_4802);
nand U6608 (N_6608,N_5908,N_5197);
or U6609 (N_6609,N_5680,N_5134);
nand U6610 (N_6610,N_5972,N_5461);
xor U6611 (N_6611,N_5244,N_5973);
and U6612 (N_6612,N_5178,N_5287);
or U6613 (N_6613,N_5754,N_4948);
nand U6614 (N_6614,N_5022,N_5003);
or U6615 (N_6615,N_4821,N_5656);
and U6616 (N_6616,N_5883,N_5270);
or U6617 (N_6617,N_5908,N_5201);
nand U6618 (N_6618,N_5607,N_5774);
nand U6619 (N_6619,N_5591,N_4890);
xor U6620 (N_6620,N_4987,N_4866);
nor U6621 (N_6621,N_5113,N_5495);
or U6622 (N_6622,N_4902,N_5001);
xor U6623 (N_6623,N_5731,N_5063);
nor U6624 (N_6624,N_5509,N_5514);
or U6625 (N_6625,N_5080,N_5182);
or U6626 (N_6626,N_5119,N_5780);
xor U6627 (N_6627,N_5700,N_5492);
nor U6628 (N_6628,N_4995,N_5310);
and U6629 (N_6629,N_4872,N_5079);
xor U6630 (N_6630,N_5570,N_5924);
nand U6631 (N_6631,N_5312,N_5788);
nand U6632 (N_6632,N_5028,N_4824);
nor U6633 (N_6633,N_5135,N_5871);
xor U6634 (N_6634,N_5948,N_5358);
and U6635 (N_6635,N_5338,N_5095);
xnor U6636 (N_6636,N_5197,N_5883);
nand U6637 (N_6637,N_5190,N_4805);
nor U6638 (N_6638,N_5995,N_5377);
nor U6639 (N_6639,N_5884,N_5589);
nand U6640 (N_6640,N_5457,N_5739);
nor U6641 (N_6641,N_5253,N_5870);
xor U6642 (N_6642,N_4960,N_4931);
nand U6643 (N_6643,N_5324,N_5788);
xor U6644 (N_6644,N_5767,N_5824);
nand U6645 (N_6645,N_5976,N_5318);
xor U6646 (N_6646,N_5807,N_5748);
xor U6647 (N_6647,N_5441,N_5383);
nand U6648 (N_6648,N_5558,N_5271);
or U6649 (N_6649,N_5419,N_5989);
nor U6650 (N_6650,N_5516,N_5017);
nand U6651 (N_6651,N_5518,N_5724);
and U6652 (N_6652,N_5969,N_5313);
nand U6653 (N_6653,N_5105,N_4823);
and U6654 (N_6654,N_4859,N_5074);
xor U6655 (N_6655,N_5953,N_5876);
and U6656 (N_6656,N_5126,N_5842);
nor U6657 (N_6657,N_5555,N_4906);
xor U6658 (N_6658,N_5306,N_5521);
nand U6659 (N_6659,N_5310,N_5697);
xnor U6660 (N_6660,N_5444,N_5298);
or U6661 (N_6661,N_5853,N_5967);
or U6662 (N_6662,N_5762,N_5197);
nor U6663 (N_6663,N_4951,N_5998);
xnor U6664 (N_6664,N_5351,N_5719);
nor U6665 (N_6665,N_5295,N_4831);
or U6666 (N_6666,N_5970,N_4949);
nor U6667 (N_6667,N_5066,N_5412);
and U6668 (N_6668,N_5760,N_5925);
nand U6669 (N_6669,N_5842,N_5926);
nand U6670 (N_6670,N_5659,N_5962);
nand U6671 (N_6671,N_5768,N_5560);
xor U6672 (N_6672,N_5028,N_5416);
xnor U6673 (N_6673,N_5677,N_5929);
or U6674 (N_6674,N_5415,N_5034);
xnor U6675 (N_6675,N_5378,N_5453);
nor U6676 (N_6676,N_5215,N_4937);
xor U6677 (N_6677,N_5525,N_5286);
nor U6678 (N_6678,N_5122,N_4907);
or U6679 (N_6679,N_5895,N_4907);
nand U6680 (N_6680,N_5131,N_5965);
and U6681 (N_6681,N_5440,N_5624);
or U6682 (N_6682,N_5722,N_5699);
nand U6683 (N_6683,N_4994,N_5483);
xor U6684 (N_6684,N_5264,N_5693);
xor U6685 (N_6685,N_5223,N_5653);
or U6686 (N_6686,N_4970,N_5663);
nand U6687 (N_6687,N_4934,N_5535);
nand U6688 (N_6688,N_5566,N_5437);
or U6689 (N_6689,N_5826,N_5723);
and U6690 (N_6690,N_5909,N_5076);
nand U6691 (N_6691,N_4999,N_5317);
nand U6692 (N_6692,N_4855,N_5626);
and U6693 (N_6693,N_5912,N_5082);
xor U6694 (N_6694,N_4961,N_4823);
nor U6695 (N_6695,N_4988,N_5734);
nor U6696 (N_6696,N_5306,N_5934);
nand U6697 (N_6697,N_5319,N_4990);
nor U6698 (N_6698,N_4988,N_5694);
nand U6699 (N_6699,N_5673,N_5726);
nand U6700 (N_6700,N_5300,N_5410);
nor U6701 (N_6701,N_5037,N_5433);
nand U6702 (N_6702,N_5778,N_5281);
xnor U6703 (N_6703,N_5684,N_5528);
xor U6704 (N_6704,N_5154,N_4977);
or U6705 (N_6705,N_5247,N_4884);
xor U6706 (N_6706,N_5860,N_4937);
or U6707 (N_6707,N_5081,N_5259);
xor U6708 (N_6708,N_5914,N_4882);
xor U6709 (N_6709,N_5414,N_5107);
xor U6710 (N_6710,N_5640,N_5468);
xnor U6711 (N_6711,N_5454,N_5593);
or U6712 (N_6712,N_5458,N_5381);
nand U6713 (N_6713,N_5266,N_4847);
or U6714 (N_6714,N_5167,N_5676);
nor U6715 (N_6715,N_5360,N_5891);
nand U6716 (N_6716,N_5983,N_4944);
xnor U6717 (N_6717,N_5529,N_5957);
xor U6718 (N_6718,N_5211,N_4975);
nor U6719 (N_6719,N_4866,N_5799);
and U6720 (N_6720,N_5826,N_5850);
nand U6721 (N_6721,N_5966,N_5097);
or U6722 (N_6722,N_5841,N_5247);
and U6723 (N_6723,N_5291,N_5233);
nor U6724 (N_6724,N_5615,N_4854);
xnor U6725 (N_6725,N_5905,N_5906);
and U6726 (N_6726,N_5188,N_4850);
and U6727 (N_6727,N_5791,N_5186);
nand U6728 (N_6728,N_4959,N_5825);
and U6729 (N_6729,N_5709,N_5880);
xnor U6730 (N_6730,N_5417,N_5135);
and U6731 (N_6731,N_5644,N_5508);
or U6732 (N_6732,N_5080,N_5739);
xnor U6733 (N_6733,N_5066,N_5913);
xnor U6734 (N_6734,N_5488,N_5858);
xnor U6735 (N_6735,N_5950,N_5742);
nand U6736 (N_6736,N_4943,N_5473);
or U6737 (N_6737,N_5338,N_5517);
xnor U6738 (N_6738,N_4955,N_5953);
and U6739 (N_6739,N_5892,N_5006);
or U6740 (N_6740,N_4901,N_5016);
and U6741 (N_6741,N_5089,N_5388);
nor U6742 (N_6742,N_5630,N_5025);
and U6743 (N_6743,N_5912,N_5834);
nand U6744 (N_6744,N_4910,N_5018);
xnor U6745 (N_6745,N_5028,N_5457);
nand U6746 (N_6746,N_5896,N_5434);
xnor U6747 (N_6747,N_5006,N_5709);
nand U6748 (N_6748,N_4898,N_5680);
and U6749 (N_6749,N_5046,N_5230);
or U6750 (N_6750,N_5307,N_5741);
nor U6751 (N_6751,N_5404,N_5443);
and U6752 (N_6752,N_5101,N_5255);
nand U6753 (N_6753,N_5838,N_4987);
or U6754 (N_6754,N_5331,N_5996);
nor U6755 (N_6755,N_4923,N_4993);
nand U6756 (N_6756,N_5670,N_5634);
nand U6757 (N_6757,N_5689,N_5187);
nand U6758 (N_6758,N_5126,N_5556);
or U6759 (N_6759,N_5074,N_5657);
nor U6760 (N_6760,N_5423,N_5451);
or U6761 (N_6761,N_5163,N_5856);
nor U6762 (N_6762,N_5758,N_5513);
nand U6763 (N_6763,N_5855,N_5392);
xnor U6764 (N_6764,N_5825,N_5531);
nand U6765 (N_6765,N_5135,N_5043);
nand U6766 (N_6766,N_5751,N_5831);
nand U6767 (N_6767,N_5273,N_5887);
and U6768 (N_6768,N_5900,N_5157);
and U6769 (N_6769,N_5240,N_5035);
xnor U6770 (N_6770,N_5018,N_5645);
nor U6771 (N_6771,N_4988,N_5948);
nor U6772 (N_6772,N_5352,N_4853);
nor U6773 (N_6773,N_4800,N_5416);
or U6774 (N_6774,N_4899,N_5459);
xor U6775 (N_6775,N_5346,N_5431);
xnor U6776 (N_6776,N_5227,N_5379);
nor U6777 (N_6777,N_5541,N_5167);
or U6778 (N_6778,N_5638,N_5717);
or U6779 (N_6779,N_5921,N_5814);
or U6780 (N_6780,N_5391,N_5826);
nor U6781 (N_6781,N_5676,N_5454);
nand U6782 (N_6782,N_5875,N_5784);
and U6783 (N_6783,N_5053,N_5597);
nor U6784 (N_6784,N_5160,N_5128);
or U6785 (N_6785,N_5763,N_5573);
or U6786 (N_6786,N_5150,N_5138);
nor U6787 (N_6787,N_5418,N_4913);
nor U6788 (N_6788,N_5211,N_5612);
or U6789 (N_6789,N_5781,N_5793);
nor U6790 (N_6790,N_5231,N_5358);
nand U6791 (N_6791,N_5921,N_5331);
xor U6792 (N_6792,N_5688,N_5792);
or U6793 (N_6793,N_5531,N_4863);
or U6794 (N_6794,N_5820,N_5835);
and U6795 (N_6795,N_5916,N_5702);
xor U6796 (N_6796,N_4834,N_5925);
and U6797 (N_6797,N_5901,N_5726);
xor U6798 (N_6798,N_5799,N_4952);
or U6799 (N_6799,N_5197,N_4933);
nor U6800 (N_6800,N_5321,N_5234);
xnor U6801 (N_6801,N_4908,N_5278);
or U6802 (N_6802,N_5431,N_4975);
nor U6803 (N_6803,N_5674,N_4985);
and U6804 (N_6804,N_4865,N_5708);
or U6805 (N_6805,N_5034,N_5504);
nor U6806 (N_6806,N_5571,N_5886);
nand U6807 (N_6807,N_5556,N_4883);
xnor U6808 (N_6808,N_5561,N_5900);
xor U6809 (N_6809,N_5685,N_4838);
xor U6810 (N_6810,N_5693,N_4869);
nor U6811 (N_6811,N_5224,N_5311);
or U6812 (N_6812,N_5636,N_5792);
and U6813 (N_6813,N_4996,N_4823);
nand U6814 (N_6814,N_5679,N_5444);
or U6815 (N_6815,N_5558,N_5984);
nor U6816 (N_6816,N_5959,N_5848);
nand U6817 (N_6817,N_5710,N_5619);
nor U6818 (N_6818,N_5022,N_5344);
nor U6819 (N_6819,N_5267,N_5278);
xor U6820 (N_6820,N_4965,N_5413);
nand U6821 (N_6821,N_5979,N_4842);
nor U6822 (N_6822,N_5740,N_5165);
nor U6823 (N_6823,N_5065,N_5614);
xnor U6824 (N_6824,N_5141,N_5930);
or U6825 (N_6825,N_5809,N_5460);
nor U6826 (N_6826,N_5265,N_5108);
xor U6827 (N_6827,N_5300,N_5102);
nand U6828 (N_6828,N_5907,N_5395);
xnor U6829 (N_6829,N_4852,N_5734);
or U6830 (N_6830,N_5138,N_5891);
and U6831 (N_6831,N_4907,N_5543);
or U6832 (N_6832,N_4968,N_5448);
or U6833 (N_6833,N_5855,N_5107);
nand U6834 (N_6834,N_5098,N_5659);
nand U6835 (N_6835,N_5283,N_5530);
xnor U6836 (N_6836,N_4919,N_5436);
nand U6837 (N_6837,N_4827,N_5757);
or U6838 (N_6838,N_5199,N_5640);
nor U6839 (N_6839,N_4967,N_5463);
nor U6840 (N_6840,N_5029,N_5116);
nand U6841 (N_6841,N_5597,N_5439);
or U6842 (N_6842,N_5264,N_5353);
or U6843 (N_6843,N_5814,N_5184);
xor U6844 (N_6844,N_4959,N_5881);
nor U6845 (N_6845,N_5683,N_5363);
xor U6846 (N_6846,N_5726,N_4888);
and U6847 (N_6847,N_5216,N_5830);
or U6848 (N_6848,N_5952,N_5503);
xnor U6849 (N_6849,N_5577,N_4916);
or U6850 (N_6850,N_5336,N_5703);
nand U6851 (N_6851,N_5144,N_5422);
nand U6852 (N_6852,N_5987,N_4990);
or U6853 (N_6853,N_5524,N_5487);
xor U6854 (N_6854,N_5076,N_5765);
nor U6855 (N_6855,N_4888,N_5432);
or U6856 (N_6856,N_5371,N_5769);
nand U6857 (N_6857,N_4931,N_5376);
and U6858 (N_6858,N_5064,N_4897);
and U6859 (N_6859,N_5647,N_5116);
or U6860 (N_6860,N_5593,N_5850);
or U6861 (N_6861,N_5335,N_5823);
and U6862 (N_6862,N_5801,N_5883);
xor U6863 (N_6863,N_5381,N_5219);
and U6864 (N_6864,N_5689,N_5011);
and U6865 (N_6865,N_5103,N_5009);
or U6866 (N_6866,N_4987,N_5994);
or U6867 (N_6867,N_4900,N_5169);
or U6868 (N_6868,N_5251,N_4937);
nand U6869 (N_6869,N_5411,N_5199);
nand U6870 (N_6870,N_5316,N_5780);
or U6871 (N_6871,N_5104,N_5309);
nor U6872 (N_6872,N_5886,N_5955);
or U6873 (N_6873,N_5266,N_5777);
and U6874 (N_6874,N_5090,N_5049);
and U6875 (N_6875,N_5088,N_5723);
nand U6876 (N_6876,N_5344,N_5005);
or U6877 (N_6877,N_5723,N_5408);
or U6878 (N_6878,N_5247,N_5160);
and U6879 (N_6879,N_5946,N_5191);
xnor U6880 (N_6880,N_4976,N_5343);
and U6881 (N_6881,N_5368,N_5486);
nor U6882 (N_6882,N_4964,N_5467);
or U6883 (N_6883,N_5382,N_5571);
or U6884 (N_6884,N_5234,N_5216);
or U6885 (N_6885,N_5622,N_5257);
nand U6886 (N_6886,N_5559,N_5667);
and U6887 (N_6887,N_5273,N_5865);
xor U6888 (N_6888,N_5936,N_5590);
xor U6889 (N_6889,N_5300,N_5924);
nand U6890 (N_6890,N_5406,N_5909);
xor U6891 (N_6891,N_5716,N_5458);
xnor U6892 (N_6892,N_5538,N_5144);
nand U6893 (N_6893,N_5864,N_5816);
nand U6894 (N_6894,N_5987,N_4952);
and U6895 (N_6895,N_5758,N_4922);
and U6896 (N_6896,N_5993,N_5756);
and U6897 (N_6897,N_5793,N_5858);
nand U6898 (N_6898,N_5225,N_5279);
xor U6899 (N_6899,N_5442,N_5036);
and U6900 (N_6900,N_5392,N_5017);
nor U6901 (N_6901,N_5171,N_5037);
xor U6902 (N_6902,N_4901,N_5561);
nor U6903 (N_6903,N_5541,N_5230);
and U6904 (N_6904,N_5166,N_5486);
or U6905 (N_6905,N_4842,N_5407);
and U6906 (N_6906,N_5549,N_5876);
nand U6907 (N_6907,N_5905,N_5262);
and U6908 (N_6908,N_5090,N_5686);
nand U6909 (N_6909,N_4939,N_5637);
nor U6910 (N_6910,N_4916,N_5492);
and U6911 (N_6911,N_5330,N_5189);
nor U6912 (N_6912,N_5317,N_5611);
xnor U6913 (N_6913,N_5205,N_5405);
nand U6914 (N_6914,N_5439,N_5351);
xnor U6915 (N_6915,N_4852,N_5008);
nor U6916 (N_6916,N_5853,N_4926);
nand U6917 (N_6917,N_5115,N_5420);
nor U6918 (N_6918,N_5315,N_5702);
and U6919 (N_6919,N_5212,N_5470);
nor U6920 (N_6920,N_4842,N_5332);
or U6921 (N_6921,N_5330,N_5253);
and U6922 (N_6922,N_5085,N_4908);
xnor U6923 (N_6923,N_5899,N_5493);
and U6924 (N_6924,N_5367,N_5926);
or U6925 (N_6925,N_5280,N_5659);
nand U6926 (N_6926,N_5335,N_5858);
nand U6927 (N_6927,N_5944,N_5839);
nor U6928 (N_6928,N_5232,N_4841);
and U6929 (N_6929,N_4801,N_4846);
xor U6930 (N_6930,N_5724,N_5948);
nor U6931 (N_6931,N_5337,N_5714);
xor U6932 (N_6932,N_4967,N_4805);
or U6933 (N_6933,N_5045,N_5410);
xnor U6934 (N_6934,N_5998,N_5537);
and U6935 (N_6935,N_5379,N_5561);
and U6936 (N_6936,N_4981,N_5481);
nand U6937 (N_6937,N_5382,N_5646);
nand U6938 (N_6938,N_5505,N_5877);
or U6939 (N_6939,N_5698,N_5810);
nor U6940 (N_6940,N_4928,N_5328);
nand U6941 (N_6941,N_5026,N_5006);
nor U6942 (N_6942,N_5101,N_4960);
and U6943 (N_6943,N_5220,N_5612);
nor U6944 (N_6944,N_5204,N_5793);
xnor U6945 (N_6945,N_5997,N_5784);
nand U6946 (N_6946,N_5399,N_5818);
and U6947 (N_6947,N_4857,N_5173);
and U6948 (N_6948,N_5944,N_5533);
nor U6949 (N_6949,N_5005,N_4849);
nand U6950 (N_6950,N_4903,N_5802);
and U6951 (N_6951,N_5982,N_5450);
xnor U6952 (N_6952,N_5049,N_5114);
xor U6953 (N_6953,N_5696,N_5733);
xnor U6954 (N_6954,N_5812,N_5963);
nor U6955 (N_6955,N_4895,N_5852);
nor U6956 (N_6956,N_5650,N_5384);
or U6957 (N_6957,N_5873,N_5423);
nor U6958 (N_6958,N_5848,N_5910);
nor U6959 (N_6959,N_5163,N_5102);
xnor U6960 (N_6960,N_5057,N_4856);
or U6961 (N_6961,N_5262,N_5141);
xor U6962 (N_6962,N_4980,N_4854);
and U6963 (N_6963,N_5730,N_5970);
or U6964 (N_6964,N_5239,N_5593);
nand U6965 (N_6965,N_5871,N_4853);
xor U6966 (N_6966,N_4954,N_5012);
or U6967 (N_6967,N_5494,N_5966);
and U6968 (N_6968,N_5838,N_5595);
and U6969 (N_6969,N_5170,N_5723);
or U6970 (N_6970,N_5056,N_5900);
nor U6971 (N_6971,N_5214,N_5198);
and U6972 (N_6972,N_5583,N_5783);
or U6973 (N_6973,N_5846,N_5739);
and U6974 (N_6974,N_5943,N_5244);
nand U6975 (N_6975,N_5365,N_4865);
nor U6976 (N_6976,N_5917,N_5506);
nor U6977 (N_6977,N_5979,N_5019);
or U6978 (N_6978,N_5433,N_5324);
and U6979 (N_6979,N_5080,N_5895);
and U6980 (N_6980,N_5908,N_5426);
nor U6981 (N_6981,N_5738,N_5802);
xnor U6982 (N_6982,N_5790,N_5813);
xor U6983 (N_6983,N_5944,N_5020);
nand U6984 (N_6984,N_5149,N_5105);
or U6985 (N_6985,N_4852,N_5840);
xnor U6986 (N_6986,N_5284,N_5400);
or U6987 (N_6987,N_5820,N_5330);
or U6988 (N_6988,N_5690,N_5190);
xnor U6989 (N_6989,N_5108,N_4961);
nor U6990 (N_6990,N_5232,N_5297);
and U6991 (N_6991,N_5098,N_5927);
xnor U6992 (N_6992,N_5801,N_5114);
nand U6993 (N_6993,N_5042,N_5312);
and U6994 (N_6994,N_5418,N_5960);
nand U6995 (N_6995,N_5064,N_5599);
nor U6996 (N_6996,N_5210,N_5790);
or U6997 (N_6997,N_5023,N_5720);
nand U6998 (N_6998,N_5187,N_5114);
and U6999 (N_6999,N_5295,N_5635);
and U7000 (N_7000,N_5864,N_5512);
xor U7001 (N_7001,N_5341,N_5981);
or U7002 (N_7002,N_4820,N_5271);
or U7003 (N_7003,N_5797,N_4939);
and U7004 (N_7004,N_5451,N_5359);
nor U7005 (N_7005,N_5048,N_5639);
and U7006 (N_7006,N_5365,N_5594);
nand U7007 (N_7007,N_5314,N_5377);
nand U7008 (N_7008,N_5988,N_5695);
or U7009 (N_7009,N_5059,N_4932);
or U7010 (N_7010,N_5465,N_5443);
and U7011 (N_7011,N_5155,N_5396);
nor U7012 (N_7012,N_5903,N_5130);
and U7013 (N_7013,N_5958,N_5911);
nor U7014 (N_7014,N_5452,N_4812);
nor U7015 (N_7015,N_5520,N_4972);
nor U7016 (N_7016,N_5915,N_4810);
xnor U7017 (N_7017,N_5913,N_5836);
xnor U7018 (N_7018,N_4964,N_5295);
and U7019 (N_7019,N_5358,N_5610);
xnor U7020 (N_7020,N_5423,N_5718);
nor U7021 (N_7021,N_5471,N_5674);
xor U7022 (N_7022,N_5670,N_5032);
or U7023 (N_7023,N_5002,N_5997);
nand U7024 (N_7024,N_5534,N_4955);
or U7025 (N_7025,N_5941,N_5813);
nand U7026 (N_7026,N_5551,N_4812);
and U7027 (N_7027,N_5535,N_5491);
nor U7028 (N_7028,N_4840,N_5797);
nor U7029 (N_7029,N_5902,N_5249);
and U7030 (N_7030,N_5638,N_5690);
nand U7031 (N_7031,N_5082,N_5799);
nand U7032 (N_7032,N_5845,N_5010);
xnor U7033 (N_7033,N_5971,N_4862);
nor U7034 (N_7034,N_4882,N_5134);
nor U7035 (N_7035,N_5296,N_5168);
nor U7036 (N_7036,N_4894,N_5653);
or U7037 (N_7037,N_5303,N_5164);
or U7038 (N_7038,N_5882,N_5446);
and U7039 (N_7039,N_5626,N_5397);
xor U7040 (N_7040,N_5733,N_5491);
xnor U7041 (N_7041,N_5612,N_5012);
nand U7042 (N_7042,N_5059,N_5430);
nor U7043 (N_7043,N_5095,N_5060);
xnor U7044 (N_7044,N_5174,N_5738);
and U7045 (N_7045,N_5778,N_5116);
or U7046 (N_7046,N_5494,N_5944);
nor U7047 (N_7047,N_5823,N_5895);
or U7048 (N_7048,N_5767,N_5953);
nand U7049 (N_7049,N_5182,N_5950);
nand U7050 (N_7050,N_5938,N_5258);
nand U7051 (N_7051,N_4898,N_4822);
nor U7052 (N_7052,N_5815,N_4929);
nand U7053 (N_7053,N_5671,N_4824);
or U7054 (N_7054,N_5667,N_5313);
nor U7055 (N_7055,N_5555,N_5303);
or U7056 (N_7056,N_5273,N_5138);
and U7057 (N_7057,N_5084,N_5633);
and U7058 (N_7058,N_5344,N_5687);
nor U7059 (N_7059,N_4878,N_5188);
and U7060 (N_7060,N_4868,N_5798);
or U7061 (N_7061,N_5001,N_5399);
nand U7062 (N_7062,N_5109,N_5562);
nor U7063 (N_7063,N_5342,N_5295);
xnor U7064 (N_7064,N_5763,N_5041);
or U7065 (N_7065,N_4824,N_5605);
or U7066 (N_7066,N_5767,N_5105);
or U7067 (N_7067,N_5263,N_5752);
or U7068 (N_7068,N_4906,N_5027);
nor U7069 (N_7069,N_5775,N_5360);
and U7070 (N_7070,N_5007,N_5049);
or U7071 (N_7071,N_5918,N_5456);
or U7072 (N_7072,N_4961,N_5627);
and U7073 (N_7073,N_5726,N_4982);
xor U7074 (N_7074,N_5244,N_5499);
nor U7075 (N_7075,N_5191,N_5797);
xor U7076 (N_7076,N_5378,N_5244);
and U7077 (N_7077,N_4889,N_5306);
or U7078 (N_7078,N_5094,N_5642);
and U7079 (N_7079,N_5129,N_5651);
and U7080 (N_7080,N_4891,N_4811);
xnor U7081 (N_7081,N_5633,N_5854);
and U7082 (N_7082,N_5670,N_5519);
and U7083 (N_7083,N_5048,N_5501);
nand U7084 (N_7084,N_5097,N_5509);
nand U7085 (N_7085,N_5539,N_5597);
or U7086 (N_7086,N_5669,N_5242);
nand U7087 (N_7087,N_5084,N_5527);
and U7088 (N_7088,N_5588,N_5704);
nand U7089 (N_7089,N_4979,N_5069);
or U7090 (N_7090,N_5284,N_5600);
or U7091 (N_7091,N_5087,N_5771);
nand U7092 (N_7092,N_5644,N_5662);
and U7093 (N_7093,N_4823,N_5671);
xor U7094 (N_7094,N_5877,N_5601);
nand U7095 (N_7095,N_5585,N_5949);
or U7096 (N_7096,N_5806,N_4873);
and U7097 (N_7097,N_5900,N_5200);
nor U7098 (N_7098,N_5240,N_5963);
nor U7099 (N_7099,N_5011,N_5481);
or U7100 (N_7100,N_5593,N_5502);
nor U7101 (N_7101,N_5652,N_5851);
nor U7102 (N_7102,N_4960,N_5618);
nor U7103 (N_7103,N_5669,N_5381);
or U7104 (N_7104,N_5556,N_5588);
and U7105 (N_7105,N_5806,N_5109);
xnor U7106 (N_7106,N_5083,N_5816);
nand U7107 (N_7107,N_5102,N_5266);
nor U7108 (N_7108,N_5902,N_5861);
xnor U7109 (N_7109,N_5531,N_4987);
nor U7110 (N_7110,N_5554,N_5388);
or U7111 (N_7111,N_4848,N_5487);
nor U7112 (N_7112,N_5569,N_4831);
xnor U7113 (N_7113,N_5591,N_5590);
and U7114 (N_7114,N_5454,N_5892);
xor U7115 (N_7115,N_5763,N_5376);
and U7116 (N_7116,N_5979,N_5514);
nand U7117 (N_7117,N_5505,N_5262);
or U7118 (N_7118,N_5340,N_5467);
nor U7119 (N_7119,N_5543,N_4938);
nor U7120 (N_7120,N_5623,N_5141);
or U7121 (N_7121,N_5791,N_5315);
nor U7122 (N_7122,N_5965,N_5634);
nor U7123 (N_7123,N_5902,N_4967);
xnor U7124 (N_7124,N_5366,N_5971);
and U7125 (N_7125,N_5274,N_5565);
xnor U7126 (N_7126,N_5762,N_5173);
or U7127 (N_7127,N_5665,N_5096);
or U7128 (N_7128,N_5452,N_5422);
nor U7129 (N_7129,N_5103,N_4883);
xor U7130 (N_7130,N_5102,N_4810);
or U7131 (N_7131,N_5080,N_5294);
nor U7132 (N_7132,N_5369,N_5528);
and U7133 (N_7133,N_5148,N_5681);
nor U7134 (N_7134,N_4859,N_5162);
xor U7135 (N_7135,N_5079,N_5365);
nand U7136 (N_7136,N_5315,N_5234);
or U7137 (N_7137,N_5108,N_5240);
nand U7138 (N_7138,N_5603,N_4866);
xnor U7139 (N_7139,N_4963,N_5886);
or U7140 (N_7140,N_5848,N_5631);
nor U7141 (N_7141,N_5344,N_5244);
or U7142 (N_7142,N_5323,N_5710);
and U7143 (N_7143,N_5782,N_5243);
nor U7144 (N_7144,N_4906,N_5625);
and U7145 (N_7145,N_5828,N_4899);
and U7146 (N_7146,N_5407,N_4854);
or U7147 (N_7147,N_5245,N_5027);
or U7148 (N_7148,N_5708,N_5951);
xor U7149 (N_7149,N_5119,N_5750);
xor U7150 (N_7150,N_5895,N_5465);
and U7151 (N_7151,N_5291,N_5510);
or U7152 (N_7152,N_5201,N_5239);
nor U7153 (N_7153,N_5779,N_5088);
or U7154 (N_7154,N_5351,N_5983);
nand U7155 (N_7155,N_5633,N_5211);
and U7156 (N_7156,N_5882,N_5523);
or U7157 (N_7157,N_4887,N_5665);
xor U7158 (N_7158,N_5888,N_5805);
nand U7159 (N_7159,N_5532,N_5051);
and U7160 (N_7160,N_5449,N_4818);
nor U7161 (N_7161,N_5877,N_5247);
and U7162 (N_7162,N_5794,N_4890);
and U7163 (N_7163,N_5019,N_4911);
and U7164 (N_7164,N_5099,N_5669);
nand U7165 (N_7165,N_5476,N_5450);
nor U7166 (N_7166,N_5419,N_5478);
or U7167 (N_7167,N_5386,N_5414);
and U7168 (N_7168,N_5228,N_5838);
nand U7169 (N_7169,N_5921,N_5276);
and U7170 (N_7170,N_4972,N_5929);
nor U7171 (N_7171,N_5953,N_5289);
nand U7172 (N_7172,N_5247,N_5126);
nand U7173 (N_7173,N_5322,N_5528);
or U7174 (N_7174,N_5587,N_5954);
and U7175 (N_7175,N_5619,N_4834);
nor U7176 (N_7176,N_5174,N_5075);
nor U7177 (N_7177,N_5019,N_5308);
or U7178 (N_7178,N_5858,N_4885);
and U7179 (N_7179,N_4987,N_5136);
and U7180 (N_7180,N_5004,N_5852);
nand U7181 (N_7181,N_5369,N_5552);
nand U7182 (N_7182,N_5005,N_5789);
or U7183 (N_7183,N_5909,N_5294);
nor U7184 (N_7184,N_5520,N_5513);
xnor U7185 (N_7185,N_5454,N_4990);
nand U7186 (N_7186,N_5485,N_4828);
xnor U7187 (N_7187,N_5203,N_5960);
xor U7188 (N_7188,N_5950,N_4869);
or U7189 (N_7189,N_5108,N_4998);
nand U7190 (N_7190,N_5870,N_5210);
nor U7191 (N_7191,N_5502,N_5257);
nor U7192 (N_7192,N_5955,N_5495);
nor U7193 (N_7193,N_5040,N_5683);
nor U7194 (N_7194,N_4875,N_5702);
or U7195 (N_7195,N_5972,N_5867);
xnor U7196 (N_7196,N_5390,N_4997);
nand U7197 (N_7197,N_5709,N_4866);
nor U7198 (N_7198,N_5047,N_5370);
and U7199 (N_7199,N_5890,N_5137);
or U7200 (N_7200,N_6535,N_6523);
and U7201 (N_7201,N_6021,N_6094);
nor U7202 (N_7202,N_6589,N_6949);
xnor U7203 (N_7203,N_6050,N_7036);
and U7204 (N_7204,N_7130,N_6294);
or U7205 (N_7205,N_6482,N_7051);
nor U7206 (N_7206,N_6798,N_6669);
nand U7207 (N_7207,N_7135,N_6499);
xnor U7208 (N_7208,N_6932,N_6440);
and U7209 (N_7209,N_6147,N_7001);
nor U7210 (N_7210,N_6348,N_7000);
nand U7211 (N_7211,N_6370,N_6944);
nor U7212 (N_7212,N_6681,N_6833);
or U7213 (N_7213,N_6113,N_7005);
and U7214 (N_7214,N_6001,N_6302);
xor U7215 (N_7215,N_6404,N_6301);
nor U7216 (N_7216,N_6808,N_6586);
and U7217 (N_7217,N_7089,N_6948);
or U7218 (N_7218,N_6189,N_6090);
xor U7219 (N_7219,N_6450,N_6079);
and U7220 (N_7220,N_7020,N_6522);
and U7221 (N_7221,N_6423,N_6082);
nor U7222 (N_7222,N_7068,N_6383);
xor U7223 (N_7223,N_7158,N_7050);
xnor U7224 (N_7224,N_7132,N_6595);
nor U7225 (N_7225,N_6594,N_6496);
nor U7226 (N_7226,N_6946,N_6143);
xor U7227 (N_7227,N_6843,N_7007);
or U7228 (N_7228,N_6489,N_6792);
xor U7229 (N_7229,N_6682,N_6157);
nor U7230 (N_7230,N_6823,N_6919);
xor U7231 (N_7231,N_6203,N_6719);
and U7232 (N_7232,N_6536,N_6610);
xor U7233 (N_7233,N_6498,N_6297);
nor U7234 (N_7234,N_6325,N_7029);
or U7235 (N_7235,N_6767,N_7094);
nand U7236 (N_7236,N_6227,N_6744);
xor U7237 (N_7237,N_6637,N_6564);
xnor U7238 (N_7238,N_6083,N_6593);
or U7239 (N_7239,N_6427,N_7017);
nor U7240 (N_7240,N_6525,N_6414);
xnor U7241 (N_7241,N_6013,N_6552);
xor U7242 (N_7242,N_6092,N_6000);
nand U7243 (N_7243,N_7079,N_6753);
and U7244 (N_7244,N_6696,N_6464);
or U7245 (N_7245,N_6969,N_6903);
nand U7246 (N_7246,N_6133,N_6983);
nor U7247 (N_7247,N_6774,N_6661);
xor U7248 (N_7248,N_6517,N_6668);
xnor U7249 (N_7249,N_6511,N_6803);
or U7250 (N_7250,N_6288,N_6353);
nor U7251 (N_7251,N_6282,N_6345);
xnor U7252 (N_7252,N_6878,N_6225);
and U7253 (N_7253,N_6501,N_7103);
xnor U7254 (N_7254,N_7146,N_6573);
or U7255 (N_7255,N_6715,N_7031);
xnor U7256 (N_7256,N_6816,N_6475);
nand U7257 (N_7257,N_6289,N_6628);
xor U7258 (N_7258,N_6705,N_6989);
nor U7259 (N_7259,N_7128,N_6468);
and U7260 (N_7260,N_6200,N_6743);
or U7261 (N_7261,N_6048,N_6388);
xor U7262 (N_7262,N_6670,N_6640);
xor U7263 (N_7263,N_6745,N_7117);
nand U7264 (N_7264,N_6747,N_6939);
xor U7265 (N_7265,N_6036,N_6198);
xor U7266 (N_7266,N_6003,N_6487);
nor U7267 (N_7267,N_6779,N_6902);
nand U7268 (N_7268,N_6035,N_6725);
or U7269 (N_7269,N_6754,N_6987);
and U7270 (N_7270,N_6925,N_6758);
nand U7271 (N_7271,N_7041,N_6002);
or U7272 (N_7272,N_6988,N_6343);
and U7273 (N_7273,N_6570,N_6030);
xnor U7274 (N_7274,N_6472,N_6274);
xor U7275 (N_7275,N_6955,N_6558);
and U7276 (N_7276,N_7012,N_6992);
or U7277 (N_7277,N_7184,N_6587);
or U7278 (N_7278,N_6395,N_6749);
nand U7279 (N_7279,N_6675,N_7198);
and U7280 (N_7280,N_7084,N_7160);
or U7281 (N_7281,N_7099,N_6645);
and U7282 (N_7282,N_6430,N_6951);
and U7283 (N_7283,N_7067,N_6249);
or U7284 (N_7284,N_6125,N_7043);
or U7285 (N_7285,N_7060,N_6034);
and U7286 (N_7286,N_6875,N_6060);
nor U7287 (N_7287,N_6124,N_6463);
xnor U7288 (N_7288,N_6602,N_6935);
or U7289 (N_7289,N_6802,N_7171);
nor U7290 (N_7290,N_6380,N_6695);
nor U7291 (N_7291,N_6757,N_6128);
and U7292 (N_7292,N_7155,N_6904);
and U7293 (N_7293,N_6748,N_6055);
and U7294 (N_7294,N_6694,N_6782);
nand U7295 (N_7295,N_6372,N_6152);
xnor U7296 (N_7296,N_7145,N_6677);
nor U7297 (N_7297,N_6484,N_6993);
nand U7298 (N_7298,N_6712,N_7070);
nand U7299 (N_7299,N_6374,N_7078);
and U7300 (N_7300,N_6963,N_7091);
or U7301 (N_7301,N_6797,N_6265);
nand U7302 (N_7302,N_6201,N_7149);
nand U7303 (N_7303,N_6834,N_6238);
nor U7304 (N_7304,N_6307,N_6512);
nand U7305 (N_7305,N_6876,N_6258);
xnor U7306 (N_7306,N_6391,N_6037);
or U7307 (N_7307,N_6477,N_6598);
nor U7308 (N_7308,N_6722,N_6017);
xnor U7309 (N_7309,N_6480,N_6112);
nand U7310 (N_7310,N_6340,N_6977);
or U7311 (N_7311,N_7055,N_6850);
xnor U7312 (N_7312,N_7147,N_6052);
nor U7313 (N_7313,N_6896,N_6106);
xnor U7314 (N_7314,N_6259,N_6316);
and U7315 (N_7315,N_6245,N_7129);
nand U7316 (N_7316,N_6364,N_6400);
xnor U7317 (N_7317,N_6365,N_6454);
nor U7318 (N_7318,N_6785,N_6350);
xnor U7319 (N_7319,N_6953,N_6699);
or U7320 (N_7320,N_6444,N_6691);
or U7321 (N_7321,N_6672,N_6917);
and U7322 (N_7322,N_6393,N_6402);
nor U7323 (N_7323,N_6369,N_6293);
and U7324 (N_7324,N_6028,N_6905);
nand U7325 (N_7325,N_6131,N_6280);
xnor U7326 (N_7326,N_6039,N_6019);
or U7327 (N_7327,N_6537,N_6229);
and U7328 (N_7328,N_6202,N_7112);
or U7329 (N_7329,N_6631,N_6979);
nor U7330 (N_7330,N_6271,N_6144);
nor U7331 (N_7331,N_6199,N_6132);
nand U7332 (N_7332,N_6267,N_7018);
nor U7333 (N_7333,N_6460,N_7056);
and U7334 (N_7334,N_6074,N_7090);
nand U7335 (N_7335,N_6295,N_6109);
nor U7336 (N_7336,N_6241,N_6807);
or U7337 (N_7337,N_7166,N_7006);
and U7338 (N_7338,N_6726,N_7151);
nand U7339 (N_7339,N_6663,N_6142);
nor U7340 (N_7340,N_6441,N_6111);
or U7341 (N_7341,N_6491,N_7190);
nand U7342 (N_7342,N_6016,N_6257);
and U7343 (N_7343,N_6762,N_6746);
xnor U7344 (N_7344,N_6795,N_6879);
xnor U7345 (N_7345,N_7064,N_6261);
xor U7346 (N_7346,N_7186,N_6967);
xor U7347 (N_7347,N_7052,N_6592);
or U7348 (N_7348,N_6553,N_7048);
nand U7349 (N_7349,N_6099,N_6260);
or U7350 (N_7350,N_6309,N_6248);
xnor U7351 (N_7351,N_6390,N_6780);
and U7352 (N_7352,N_6394,N_6997);
and U7353 (N_7353,N_6510,N_6930);
nand U7354 (N_7354,N_6545,N_6880);
and U7355 (N_7355,N_6086,N_7107);
nand U7356 (N_7356,N_6852,N_6772);
or U7357 (N_7357,N_6867,N_6004);
xor U7358 (N_7358,N_7077,N_6126);
nand U7359 (N_7359,N_6204,N_7042);
or U7360 (N_7360,N_7022,N_7110);
and U7361 (N_7361,N_6161,N_6130);
xnor U7362 (N_7362,N_6116,N_6541);
nor U7363 (N_7363,N_6217,N_6188);
nor U7364 (N_7364,N_7183,N_6599);
xor U7365 (N_7365,N_6135,N_6614);
nor U7366 (N_7366,N_6662,N_6693);
nor U7367 (N_7367,N_6974,N_7141);
nor U7368 (N_7368,N_6584,N_6874);
nand U7369 (N_7369,N_6296,N_6127);
nand U7370 (N_7370,N_6162,N_6713);
or U7371 (N_7371,N_7137,N_7027);
nor U7372 (N_7372,N_6462,N_6458);
nor U7373 (N_7373,N_6829,N_6508);
nor U7374 (N_7374,N_6585,N_7182);
or U7375 (N_7375,N_6165,N_6548);
or U7376 (N_7376,N_6976,N_6826);
nor U7377 (N_7377,N_6755,N_6539);
xnor U7378 (N_7378,N_6627,N_6591);
and U7379 (N_7379,N_7087,N_6886);
and U7380 (N_7380,N_6597,N_6686);
and U7381 (N_7381,N_6961,N_6980);
and U7382 (N_7382,N_6262,N_6190);
and U7383 (N_7383,N_6211,N_6895);
nand U7384 (N_7384,N_7081,N_6731);
and U7385 (N_7385,N_6366,N_6275);
or U7386 (N_7386,N_6168,N_7121);
or U7387 (N_7387,N_6428,N_6520);
nor U7388 (N_7388,N_6576,N_6840);
or U7389 (N_7389,N_6445,N_6054);
and U7390 (N_7390,N_6381,N_6407);
and U7391 (N_7391,N_6105,N_6721);
and U7392 (N_7392,N_6760,N_6174);
xnor U7393 (N_7393,N_6865,N_6115);
nor U7394 (N_7394,N_6065,N_6253);
nor U7395 (N_7395,N_7049,N_6818);
nor U7396 (N_7396,N_6853,N_6416);
or U7397 (N_7397,N_6192,N_7069);
nor U7398 (N_7398,N_6479,N_7045);
nor U7399 (N_7399,N_6089,N_7169);
nand U7400 (N_7400,N_6326,N_6418);
and U7401 (N_7401,N_6958,N_6351);
and U7402 (N_7402,N_6665,N_6146);
and U7403 (N_7403,N_6411,N_7122);
nand U7404 (N_7404,N_7100,N_6329);
and U7405 (N_7405,N_6333,N_7059);
nand U7406 (N_7406,N_6531,N_6352);
or U7407 (N_7407,N_6358,N_6473);
nor U7408 (N_7408,N_6942,N_6470);
xnor U7409 (N_7409,N_6179,N_6196);
nand U7410 (N_7410,N_6193,N_7024);
nand U7411 (N_7411,N_6616,N_6800);
xor U7412 (N_7412,N_6397,N_6172);
or U7413 (N_7413,N_6141,N_6442);
or U7414 (N_7414,N_6024,N_7011);
nand U7415 (N_7415,N_6098,N_6737);
and U7416 (N_7416,N_6457,N_6998);
and U7417 (N_7417,N_6776,N_6076);
and U7418 (N_7418,N_6509,N_6062);
or U7419 (N_7419,N_6007,N_6443);
nor U7420 (N_7420,N_6031,N_6424);
xnor U7421 (N_7421,N_6419,N_6488);
nand U7422 (N_7422,N_7126,N_7008);
or U7423 (N_7423,N_6654,N_6102);
nand U7424 (N_7424,N_6729,N_6505);
nand U7425 (N_7425,N_7080,N_6711);
or U7426 (N_7426,N_6866,N_6342);
nor U7427 (N_7427,N_6435,N_6909);
nand U7428 (N_7428,N_6331,N_6378);
nor U7429 (N_7429,N_6040,N_6611);
nand U7430 (N_7430,N_6367,N_6292);
nor U7431 (N_7431,N_6354,N_6735);
nor U7432 (N_7432,N_7074,N_6891);
xnor U7433 (N_7433,N_7014,N_6108);
and U7434 (N_7434,N_6384,N_6888);
or U7435 (N_7435,N_6844,N_6213);
xor U7436 (N_7436,N_6952,N_6945);
or U7437 (N_7437,N_6680,N_6566);
and U7438 (N_7438,N_6169,N_6527);
nor U7439 (N_7439,N_6349,N_7199);
nor U7440 (N_7440,N_6873,N_6330);
xnor U7441 (N_7441,N_6718,N_7082);
or U7442 (N_7442,N_6363,N_7072);
nand U7443 (N_7443,N_7021,N_6978);
or U7444 (N_7444,N_7123,N_7062);
xnor U7445 (N_7445,N_6129,N_6625);
nand U7446 (N_7446,N_6273,N_6756);
nor U7447 (N_7447,N_6839,N_6913);
or U7448 (N_7448,N_6250,N_6077);
and U7449 (N_7449,N_6042,N_6813);
nand U7450 (N_7450,N_6436,N_6860);
nand U7451 (N_7451,N_6892,N_6674);
nand U7452 (N_7452,N_6068,N_6810);
or U7453 (N_7453,N_6707,N_6927);
xnor U7454 (N_7454,N_6264,N_6559);
nand U7455 (N_7455,N_6177,N_7150);
or U7456 (N_7456,N_6449,N_6371);
and U7457 (N_7457,N_7019,N_7101);
nand U7458 (N_7458,N_6434,N_6461);
nor U7459 (N_7459,N_6377,N_6912);
or U7460 (N_7460,N_6555,N_6986);
and U7461 (N_7461,N_6059,N_6032);
nor U7462 (N_7462,N_7176,N_6359);
and U7463 (N_7463,N_6882,N_6690);
and U7464 (N_7464,N_6075,N_6619);
xor U7465 (N_7465,N_6409,N_7061);
or U7466 (N_7466,N_7088,N_6362);
or U7467 (N_7467,N_7044,N_6119);
or U7468 (N_7468,N_7115,N_6284);
or U7469 (N_7469,N_6734,N_6242);
xnor U7470 (N_7470,N_6455,N_6815);
or U7471 (N_7471,N_6982,N_6256);
xnor U7472 (N_7472,N_6981,N_6070);
or U7473 (N_7473,N_6306,N_7127);
xor U7474 (N_7474,N_6970,N_6583);
xnor U7475 (N_7475,N_6549,N_6012);
xor U7476 (N_7476,N_6581,N_7172);
or U7477 (N_7477,N_6825,N_6518);
nand U7478 (N_7478,N_6399,N_6123);
nand U7479 (N_7479,N_6830,N_6313);
and U7480 (N_7480,N_6376,N_6636);
nand U7481 (N_7481,N_6222,N_6255);
and U7482 (N_7482,N_6120,N_6417);
xnor U7483 (N_7483,N_6219,N_6730);
or U7484 (N_7484,N_6957,N_6228);
or U7485 (N_7485,N_6846,N_6994);
nand U7486 (N_7486,N_6101,N_6901);
or U7487 (N_7487,N_6182,N_7023);
and U7488 (N_7488,N_6678,N_7111);
or U7489 (N_7489,N_7065,N_6114);
nor U7490 (N_7490,N_6215,N_6740);
nor U7491 (N_7491,N_6160,N_6497);
nor U7492 (N_7492,N_6533,N_6838);
nor U7493 (N_7493,N_6732,N_6578);
and U7494 (N_7494,N_6990,N_6528);
nor U7495 (N_7495,N_6784,N_6622);
nor U7496 (N_7496,N_7047,N_6425);
and U7497 (N_7497,N_6053,N_6924);
or U7498 (N_7498,N_6574,N_6700);
nor U7499 (N_7499,N_6648,N_6907);
and U7500 (N_7500,N_6327,N_6438);
nor U7501 (N_7501,N_6685,N_7038);
nor U7502 (N_7502,N_6318,N_6618);
or U7503 (N_7503,N_6954,N_6596);
and U7504 (N_7504,N_6247,N_6831);
nor U7505 (N_7505,N_6185,N_6492);
nor U7506 (N_7506,N_6226,N_6991);
xor U7507 (N_7507,N_6170,N_7154);
or U7508 (N_7508,N_6601,N_6389);
and U7509 (N_7509,N_6656,N_6171);
or U7510 (N_7510,N_7098,N_6563);
nand U7511 (N_7511,N_6186,N_6936);
or U7512 (N_7512,N_6701,N_6051);
or U7513 (N_7513,N_6894,N_6044);
nand U7514 (N_7514,N_6794,N_7192);
or U7515 (N_7515,N_6557,N_6960);
nor U7516 (N_7516,N_6346,N_6720);
and U7517 (N_7517,N_7142,N_6565);
nand U7518 (N_7518,N_6214,N_6403);
nand U7519 (N_7519,N_6163,N_6504);
and U7520 (N_7520,N_6148,N_6612);
or U7521 (N_7521,N_6861,N_6777);
nand U7522 (N_7522,N_6739,N_6368);
and U7523 (N_7523,N_6856,N_6871);
nand U7524 (N_7524,N_6361,N_7073);
or U7525 (N_7525,N_7058,N_6975);
nor U7526 (N_7526,N_6862,N_6827);
xnor U7527 (N_7527,N_6630,N_6790);
and U7528 (N_7528,N_6918,N_6855);
nor U7529 (N_7529,N_6236,N_6684);
nor U7530 (N_7530,N_6095,N_7138);
nand U7531 (N_7531,N_6928,N_6658);
and U7532 (N_7532,N_6620,N_6526);
xnor U7533 (N_7533,N_6481,N_6530);
nor U7534 (N_7534,N_6929,N_6703);
or U7535 (N_7535,N_6937,N_7173);
nor U7536 (N_7536,N_6956,N_6893);
or U7537 (N_7537,N_6765,N_7136);
nand U7538 (N_7538,N_6439,N_6801);
or U7539 (N_7539,N_7095,N_6647);
or U7540 (N_7540,N_6623,N_6849);
xor U7541 (N_7541,N_6252,N_6920);
and U7542 (N_7542,N_6286,N_6884);
xnor U7543 (N_7543,N_6926,N_6809);
and U7544 (N_7544,N_6698,N_6736);
xor U7545 (N_7545,N_6448,N_6207);
xnor U7546 (N_7546,N_6011,N_6883);
xor U7547 (N_7547,N_7076,N_6379);
xnor U7548 (N_7548,N_6806,N_6476);
xor U7549 (N_7549,N_6206,N_6067);
or U7550 (N_7550,N_6406,N_6269);
xnor U7551 (N_7551,N_6870,N_6140);
xnor U7552 (N_7552,N_6465,N_6821);
or U7553 (N_7553,N_6889,N_6312);
or U7554 (N_7554,N_6154,N_6966);
nor U7555 (N_7555,N_7119,N_6532);
xnor U7556 (N_7556,N_6155,N_6164);
xor U7557 (N_7557,N_6266,N_6305);
xnor U7558 (N_7558,N_6910,N_6386);
or U7559 (N_7559,N_6317,N_6298);
xnor U7560 (N_7560,N_6344,N_6634);
nor U7561 (N_7561,N_6029,N_6704);
xor U7562 (N_7562,N_7162,N_6864);
nand U7563 (N_7563,N_6769,N_6308);
nor U7564 (N_7564,N_6290,N_7102);
and U7565 (N_7565,N_6940,N_7010);
xnor U7566 (N_7566,N_6791,N_6608);
xnor U7567 (N_7567,N_6793,N_7157);
and U7568 (N_7568,N_6649,N_6337);
nor U7569 (N_7569,N_6710,N_6321);
nand U7570 (N_7570,N_6943,N_7037);
nor U7571 (N_7571,N_6965,N_7174);
nor U7572 (N_7572,N_7164,N_6025);
nand U7573 (N_7573,N_6231,N_6385);
or U7574 (N_7574,N_6071,N_6651);
and U7575 (N_7575,N_6456,N_6159);
xor U7576 (N_7576,N_6716,N_6237);
and U7577 (N_7577,N_7168,N_6851);
or U7578 (N_7578,N_6804,N_6276);
and U7579 (N_7579,N_6666,N_6180);
or U7580 (N_7580,N_7034,N_7003);
and U7581 (N_7581,N_6121,N_6080);
nand U7582 (N_7582,N_6683,N_6322);
nor U7583 (N_7583,N_6431,N_6251);
nor U7584 (N_7584,N_6650,N_6629);
xor U7585 (N_7585,N_6515,N_6392);
or U7586 (N_7586,N_7152,N_6847);
and U7587 (N_7587,N_6224,N_7170);
nor U7588 (N_7588,N_6221,N_6659);
nand U7589 (N_7589,N_6572,N_6899);
xnor U7590 (N_7590,N_6513,N_7161);
nand U7591 (N_7591,N_6291,N_6773);
or U7592 (N_7592,N_7175,N_6263);
and U7593 (N_7593,N_6046,N_6150);
nand U7594 (N_7594,N_6551,N_7057);
xnor U7595 (N_7595,N_6660,N_6216);
or U7596 (N_7596,N_6941,N_7086);
or U7597 (N_7597,N_6569,N_6104);
nor U7598 (N_7598,N_6580,N_7032);
nor U7599 (N_7599,N_6209,N_6006);
nand U7600 (N_7600,N_6832,N_6923);
nand U7601 (N_7601,N_6087,N_6246);
or U7602 (N_7602,N_7116,N_6218);
xor U7603 (N_7603,N_6336,N_6194);
nand U7604 (N_7604,N_6724,N_6008);
xor U7605 (N_7605,N_6771,N_6277);
and U7606 (N_7606,N_6922,N_6931);
nand U7607 (N_7607,N_6934,N_6778);
or U7608 (N_7608,N_6822,N_6421);
or U7609 (N_7609,N_6401,N_6750);
xor U7610 (N_7610,N_6950,N_6692);
and U7611 (N_7611,N_6521,N_6781);
nand U7612 (N_7612,N_6287,N_6145);
or U7613 (N_7613,N_6588,N_6644);
or U7614 (N_7614,N_7028,N_6191);
and U7615 (N_7615,N_6835,N_6606);
xnor U7616 (N_7616,N_6562,N_7194);
xor U7617 (N_7617,N_7009,N_6972);
nor U7618 (N_7618,N_6540,N_6398);
nand U7619 (N_7619,N_6085,N_6023);
or U7620 (N_7620,N_6045,N_6600);
xnor U7621 (N_7621,N_6652,N_6962);
and U7622 (N_7622,N_6232,N_7026);
xnor U7623 (N_7623,N_6604,N_6347);
and U7624 (N_7624,N_7075,N_7013);
nand U7625 (N_7625,N_6728,N_6723);
nor U7626 (N_7626,N_6687,N_7131);
xnor U7627 (N_7627,N_7188,N_6529);
nor U7628 (N_7628,N_6010,N_6764);
xor U7629 (N_7629,N_6357,N_6096);
or U7630 (N_7630,N_6775,N_7093);
xor U7631 (N_7631,N_6234,N_6183);
or U7632 (N_7632,N_6617,N_6311);
xnor U7633 (N_7633,N_7156,N_6107);
nor U7634 (N_7634,N_6788,N_6877);
xor U7635 (N_7635,N_6020,N_6061);
xnor U7636 (N_7636,N_6524,N_6702);
nor U7637 (N_7637,N_6412,N_6181);
xnor U7638 (N_7638,N_6805,N_6653);
and U7639 (N_7639,N_6315,N_6947);
nor U7640 (N_7640,N_6063,N_6751);
and U7641 (N_7641,N_6270,N_6138);
or U7642 (N_7642,N_6579,N_7187);
nand U7643 (N_7643,N_7114,N_6088);
nand U7644 (N_7644,N_6733,N_6469);
or U7645 (N_7645,N_6985,N_6900);
xor U7646 (N_7646,N_6239,N_6210);
and U7647 (N_7647,N_6355,N_6100);
or U7648 (N_7648,N_6642,N_6848);
or U7649 (N_7649,N_6184,N_6243);
nor U7650 (N_7650,N_6546,N_7030);
nor U7651 (N_7651,N_7004,N_6208);
nand U7652 (N_7652,N_6117,N_6254);
or U7653 (N_7653,N_7120,N_6890);
nor U7654 (N_7654,N_7039,N_6033);
or U7655 (N_7655,N_6066,N_6568);
nand U7656 (N_7656,N_6519,N_6857);
nor U7657 (N_7657,N_6796,N_6220);
or U7658 (N_7658,N_6706,N_6471);
nand U7659 (N_7659,N_6466,N_6885);
and U7660 (N_7660,N_7179,N_6022);
and U7661 (N_7661,N_6657,N_7167);
nor U7662 (N_7662,N_6110,N_6233);
nor U7663 (N_7663,N_7163,N_7139);
and U7664 (N_7664,N_6996,N_6500);
xor U7665 (N_7665,N_6841,N_6688);
or U7666 (N_7666,N_7035,N_6405);
and U7667 (N_7667,N_6556,N_6429);
nor U7668 (N_7668,N_6836,N_6766);
and U7669 (N_7669,N_6485,N_7181);
xor U7670 (N_7670,N_6300,N_6741);
xnor U7671 (N_7671,N_6122,N_6633);
nor U7672 (N_7672,N_6026,N_6240);
and U7673 (N_7673,N_6828,N_6872);
nand U7674 (N_7674,N_6153,N_6453);
or U7675 (N_7675,N_6898,N_7191);
xnor U7676 (N_7676,N_6304,N_6671);
xnor U7677 (N_7677,N_6763,N_6420);
nand U7678 (N_7678,N_6887,N_6205);
nand U7679 (N_7679,N_7002,N_6136);
or U7680 (N_7680,N_6783,N_6058);
or U7681 (N_7681,N_6056,N_6230);
nor U7682 (N_7682,N_7106,N_6323);
and U7683 (N_7683,N_6303,N_7071);
and U7684 (N_7684,N_6655,N_6223);
and U7685 (N_7685,N_6915,N_6494);
and U7686 (N_7686,N_6921,N_6697);
xnor U7687 (N_7687,N_7189,N_6605);
and U7688 (N_7688,N_6310,N_6396);
nor U7689 (N_7689,N_6995,N_7085);
xor U7690 (N_7690,N_6167,N_7153);
nand U7691 (N_7691,N_6069,N_6507);
nor U7692 (N_7692,N_7025,N_6432);
and U7693 (N_7693,N_7133,N_6413);
and U7694 (N_7694,N_6968,N_6338);
and U7695 (N_7695,N_6502,N_6493);
nor U7696 (N_7696,N_6911,N_7054);
xor U7697 (N_7697,N_6863,N_7118);
nor U7698 (N_7698,N_6643,N_6752);
or U7699 (N_7699,N_6761,N_6073);
xor U7700 (N_7700,N_6149,N_6324);
nor U7701 (N_7701,N_6664,N_7185);
or U7702 (N_7702,N_6118,N_6639);
xnor U7703 (N_7703,N_6708,N_7177);
or U7704 (N_7704,N_6459,N_6582);
xnor U7705 (N_7705,N_6334,N_6770);
nand U7706 (N_7706,N_6447,N_6244);
and U7707 (N_7707,N_6285,N_6738);
or U7708 (N_7708,N_6868,N_7124);
nand U7709 (N_7709,N_6538,N_6005);
nand U7710 (N_7710,N_6156,N_6437);
nor U7711 (N_7711,N_7125,N_6158);
xor U7712 (N_7712,N_6103,N_6858);
and U7713 (N_7713,N_6603,N_6332);
nand U7714 (N_7714,N_6727,N_6609);
nor U7715 (N_7715,N_6786,N_6577);
nand U7716 (N_7716,N_7197,N_6817);
nor U7717 (N_7717,N_6938,N_6382);
nand U7718 (N_7718,N_6281,N_6799);
and U7719 (N_7719,N_6047,N_7159);
nand U7720 (N_7720,N_6408,N_7108);
and U7721 (N_7721,N_7033,N_6356);
or U7722 (N_7722,N_7053,N_6027);
or U7723 (N_7723,N_6544,N_6820);
and U7724 (N_7724,N_6081,N_6320);
xnor U7725 (N_7725,N_7063,N_6410);
or U7726 (N_7726,N_7015,N_6091);
nor U7727 (N_7727,N_6908,N_6195);
xor U7728 (N_7728,N_6514,N_7096);
nand U7729 (N_7729,N_7196,N_6709);
nor U7730 (N_7730,N_6933,N_6139);
nand U7731 (N_7731,N_6387,N_6984);
xnor U7732 (N_7732,N_6547,N_7016);
xor U7733 (N_7733,N_7092,N_6299);
and U7734 (N_7734,N_6789,N_6375);
nand U7735 (N_7735,N_6959,N_6768);
or U7736 (N_7736,N_6422,N_6014);
or U7737 (N_7737,N_6543,N_6667);
and U7738 (N_7738,N_7180,N_7134);
and U7739 (N_7739,N_6916,N_6516);
nor U7740 (N_7740,N_6134,N_6842);
nand U7741 (N_7741,N_6015,N_6339);
xor U7742 (N_7742,N_6814,N_6689);
xnor U7743 (N_7743,N_6971,N_6452);
or U7744 (N_7744,N_6635,N_6137);
nand U7745 (N_7745,N_6319,N_7097);
and U7746 (N_7746,N_6554,N_6426);
or U7747 (N_7747,N_6072,N_6151);
xnor U7748 (N_7748,N_6567,N_6049);
nand U7749 (N_7749,N_6845,N_6881);
nor U7750 (N_7750,N_7109,N_6607);
xor U7751 (N_7751,N_7178,N_7195);
and U7752 (N_7752,N_7193,N_6859);
and U7753 (N_7753,N_6503,N_7148);
or U7754 (N_7754,N_6575,N_6451);
nand U7755 (N_7755,N_6506,N_6854);
or U7756 (N_7756,N_6467,N_6084);
and U7757 (N_7757,N_6561,N_6283);
and U7758 (N_7758,N_6787,N_6314);
and U7759 (N_7759,N_6812,N_6235);
nand U7760 (N_7760,N_6964,N_6641);
nor U7761 (N_7761,N_6279,N_6341);
and U7762 (N_7762,N_6212,N_6613);
xor U7763 (N_7763,N_6197,N_6272);
or U7764 (N_7764,N_6433,N_6166);
and U7765 (N_7765,N_6759,N_6717);
xnor U7766 (N_7766,N_6043,N_6621);
or U7767 (N_7767,N_6869,N_6897);
nor U7768 (N_7768,N_6486,N_6446);
or U7769 (N_7769,N_6175,N_6078);
and U7770 (N_7770,N_6679,N_7144);
xnor U7771 (N_7771,N_6009,N_6590);
nand U7772 (N_7772,N_7165,N_6176);
xor U7773 (N_7773,N_7143,N_6646);
xnor U7774 (N_7774,N_7066,N_6542);
and U7775 (N_7775,N_6173,N_6676);
nand U7776 (N_7776,N_6093,N_6474);
xor U7777 (N_7777,N_6673,N_6638);
xnor U7778 (N_7778,N_6278,N_6268);
and U7779 (N_7779,N_6064,N_6819);
or U7780 (N_7780,N_6615,N_6824);
and U7781 (N_7781,N_6534,N_6742);
nand U7782 (N_7782,N_7046,N_6187);
or U7783 (N_7783,N_7040,N_6837);
and U7784 (N_7784,N_7113,N_6999);
and U7785 (N_7785,N_6038,N_6478);
xnor U7786 (N_7786,N_6415,N_6632);
nor U7787 (N_7787,N_6973,N_6714);
and U7788 (N_7788,N_7105,N_6490);
and U7789 (N_7789,N_6626,N_7104);
and U7790 (N_7790,N_6057,N_6483);
and U7791 (N_7791,N_6328,N_6373);
nand U7792 (N_7792,N_6906,N_6550);
and U7793 (N_7793,N_6018,N_7140);
nand U7794 (N_7794,N_6624,N_6811);
nor U7795 (N_7795,N_6571,N_6097);
xor U7796 (N_7796,N_6360,N_7083);
nand U7797 (N_7797,N_6178,N_6560);
nand U7798 (N_7798,N_6335,N_6041);
or U7799 (N_7799,N_6495,N_6914);
xnor U7800 (N_7800,N_6714,N_7017);
xor U7801 (N_7801,N_6155,N_6677);
xor U7802 (N_7802,N_6339,N_7009);
nand U7803 (N_7803,N_7049,N_6253);
or U7804 (N_7804,N_6842,N_6564);
and U7805 (N_7805,N_6702,N_6351);
xnor U7806 (N_7806,N_7001,N_6269);
xnor U7807 (N_7807,N_6666,N_6594);
nor U7808 (N_7808,N_6927,N_6114);
nand U7809 (N_7809,N_6579,N_7136);
nor U7810 (N_7810,N_6528,N_6443);
and U7811 (N_7811,N_7170,N_6913);
and U7812 (N_7812,N_6746,N_7043);
nor U7813 (N_7813,N_6961,N_6289);
nand U7814 (N_7814,N_6396,N_6869);
nor U7815 (N_7815,N_6591,N_6856);
nand U7816 (N_7816,N_6567,N_6469);
nand U7817 (N_7817,N_6869,N_6272);
or U7818 (N_7818,N_6713,N_6923);
and U7819 (N_7819,N_6179,N_6375);
nand U7820 (N_7820,N_6961,N_6473);
nor U7821 (N_7821,N_6470,N_6429);
xnor U7822 (N_7822,N_6777,N_6438);
nor U7823 (N_7823,N_6659,N_7140);
nand U7824 (N_7824,N_6651,N_6501);
nor U7825 (N_7825,N_6447,N_6453);
nand U7826 (N_7826,N_7104,N_6666);
nand U7827 (N_7827,N_6256,N_6616);
nor U7828 (N_7828,N_6961,N_6243);
or U7829 (N_7829,N_6823,N_6090);
and U7830 (N_7830,N_6745,N_6255);
xnor U7831 (N_7831,N_6426,N_6517);
and U7832 (N_7832,N_7017,N_6784);
nand U7833 (N_7833,N_6725,N_6098);
and U7834 (N_7834,N_6571,N_6487);
or U7835 (N_7835,N_7161,N_6278);
or U7836 (N_7836,N_6810,N_7129);
and U7837 (N_7837,N_6773,N_6957);
nor U7838 (N_7838,N_6925,N_7062);
and U7839 (N_7839,N_6471,N_6056);
nor U7840 (N_7840,N_6867,N_6497);
nand U7841 (N_7841,N_6598,N_7041);
or U7842 (N_7842,N_6342,N_7057);
or U7843 (N_7843,N_6379,N_6662);
or U7844 (N_7844,N_6144,N_7141);
or U7845 (N_7845,N_6881,N_7172);
nor U7846 (N_7846,N_7045,N_6902);
nor U7847 (N_7847,N_6092,N_6339);
nand U7848 (N_7848,N_7152,N_6396);
nand U7849 (N_7849,N_6867,N_7053);
nand U7850 (N_7850,N_7195,N_6858);
nand U7851 (N_7851,N_6496,N_6804);
or U7852 (N_7852,N_7099,N_6161);
nand U7853 (N_7853,N_6525,N_6566);
xor U7854 (N_7854,N_6216,N_7049);
or U7855 (N_7855,N_6927,N_6369);
and U7856 (N_7856,N_7018,N_7067);
nand U7857 (N_7857,N_6012,N_6347);
nand U7858 (N_7858,N_6937,N_6833);
or U7859 (N_7859,N_6684,N_6790);
xor U7860 (N_7860,N_7072,N_6238);
and U7861 (N_7861,N_6872,N_7058);
nand U7862 (N_7862,N_6878,N_6983);
or U7863 (N_7863,N_6286,N_6069);
or U7864 (N_7864,N_7060,N_6394);
or U7865 (N_7865,N_6971,N_6402);
or U7866 (N_7866,N_6796,N_6057);
nor U7867 (N_7867,N_6219,N_6095);
nand U7868 (N_7868,N_6539,N_6489);
or U7869 (N_7869,N_6822,N_6406);
and U7870 (N_7870,N_6160,N_6025);
and U7871 (N_7871,N_6180,N_7039);
or U7872 (N_7872,N_6531,N_7138);
or U7873 (N_7873,N_6507,N_6383);
or U7874 (N_7874,N_6626,N_7065);
nor U7875 (N_7875,N_7191,N_6558);
and U7876 (N_7876,N_6112,N_6310);
nand U7877 (N_7877,N_7020,N_6139);
and U7878 (N_7878,N_6664,N_6887);
nor U7879 (N_7879,N_6684,N_6674);
nand U7880 (N_7880,N_6766,N_6576);
nor U7881 (N_7881,N_6208,N_6798);
nor U7882 (N_7882,N_6259,N_6142);
nand U7883 (N_7883,N_6691,N_6696);
and U7884 (N_7884,N_6419,N_7112);
and U7885 (N_7885,N_6906,N_6057);
xor U7886 (N_7886,N_6435,N_7179);
or U7887 (N_7887,N_6154,N_6818);
nand U7888 (N_7888,N_6465,N_6010);
nand U7889 (N_7889,N_6612,N_7166);
xnor U7890 (N_7890,N_6451,N_6480);
or U7891 (N_7891,N_6258,N_6717);
nand U7892 (N_7892,N_6900,N_6481);
and U7893 (N_7893,N_6836,N_6190);
nor U7894 (N_7894,N_6708,N_6285);
nand U7895 (N_7895,N_6541,N_6717);
xor U7896 (N_7896,N_7025,N_6289);
or U7897 (N_7897,N_6983,N_6174);
or U7898 (N_7898,N_6994,N_6821);
or U7899 (N_7899,N_6500,N_6497);
nor U7900 (N_7900,N_6623,N_6541);
nand U7901 (N_7901,N_6593,N_6386);
nor U7902 (N_7902,N_6077,N_7018);
nand U7903 (N_7903,N_6877,N_6435);
and U7904 (N_7904,N_6800,N_6750);
or U7905 (N_7905,N_7016,N_7178);
and U7906 (N_7906,N_6040,N_6405);
nand U7907 (N_7907,N_6852,N_6047);
or U7908 (N_7908,N_6547,N_6829);
and U7909 (N_7909,N_6363,N_7160);
nor U7910 (N_7910,N_6869,N_6646);
nor U7911 (N_7911,N_7101,N_6015);
or U7912 (N_7912,N_6774,N_6628);
and U7913 (N_7913,N_6034,N_6380);
nor U7914 (N_7914,N_6781,N_6695);
nand U7915 (N_7915,N_6859,N_6921);
xor U7916 (N_7916,N_6136,N_6403);
or U7917 (N_7917,N_6976,N_7017);
nand U7918 (N_7918,N_6164,N_6361);
nand U7919 (N_7919,N_6925,N_6289);
xnor U7920 (N_7920,N_7057,N_6879);
nor U7921 (N_7921,N_6728,N_6067);
nor U7922 (N_7922,N_6518,N_6217);
nor U7923 (N_7923,N_7004,N_6771);
xor U7924 (N_7924,N_6061,N_6865);
or U7925 (N_7925,N_6052,N_6680);
nor U7926 (N_7926,N_6882,N_6503);
or U7927 (N_7927,N_6738,N_6144);
nor U7928 (N_7928,N_6293,N_6320);
and U7929 (N_7929,N_6928,N_6671);
or U7930 (N_7930,N_6141,N_6516);
nor U7931 (N_7931,N_7171,N_6110);
and U7932 (N_7932,N_6369,N_6047);
nand U7933 (N_7933,N_6960,N_6873);
nor U7934 (N_7934,N_7092,N_6633);
or U7935 (N_7935,N_7055,N_6786);
nor U7936 (N_7936,N_6460,N_7123);
or U7937 (N_7937,N_6730,N_6464);
nand U7938 (N_7938,N_6078,N_6900);
nor U7939 (N_7939,N_6350,N_6435);
nand U7940 (N_7940,N_6907,N_6523);
xor U7941 (N_7941,N_6967,N_6382);
or U7942 (N_7942,N_7187,N_6477);
nand U7943 (N_7943,N_6469,N_6453);
nand U7944 (N_7944,N_6583,N_6660);
xor U7945 (N_7945,N_6920,N_6308);
nand U7946 (N_7946,N_6264,N_7130);
xor U7947 (N_7947,N_6796,N_6886);
nor U7948 (N_7948,N_6401,N_6887);
nand U7949 (N_7949,N_6970,N_6395);
nor U7950 (N_7950,N_7082,N_6306);
xor U7951 (N_7951,N_6610,N_6119);
or U7952 (N_7952,N_6751,N_6221);
xnor U7953 (N_7953,N_6630,N_6769);
nor U7954 (N_7954,N_6339,N_6678);
nor U7955 (N_7955,N_6150,N_7189);
and U7956 (N_7956,N_7091,N_6004);
nand U7957 (N_7957,N_6303,N_7174);
xor U7958 (N_7958,N_7032,N_7130);
and U7959 (N_7959,N_6611,N_6325);
or U7960 (N_7960,N_6486,N_6686);
nor U7961 (N_7961,N_6068,N_6538);
or U7962 (N_7962,N_6636,N_6450);
or U7963 (N_7963,N_6318,N_6276);
or U7964 (N_7964,N_6874,N_6705);
xnor U7965 (N_7965,N_6880,N_6813);
or U7966 (N_7966,N_6726,N_6529);
xnor U7967 (N_7967,N_6600,N_6607);
or U7968 (N_7968,N_6763,N_6917);
or U7969 (N_7969,N_6162,N_6597);
and U7970 (N_7970,N_7144,N_7143);
nor U7971 (N_7971,N_6345,N_6829);
and U7972 (N_7972,N_7095,N_6473);
or U7973 (N_7973,N_6112,N_6868);
or U7974 (N_7974,N_6720,N_6388);
xor U7975 (N_7975,N_6222,N_6254);
xor U7976 (N_7976,N_6918,N_6039);
nor U7977 (N_7977,N_6672,N_7060);
xor U7978 (N_7978,N_6169,N_7017);
or U7979 (N_7979,N_6017,N_6811);
xnor U7980 (N_7980,N_6067,N_6994);
nand U7981 (N_7981,N_7074,N_6349);
xor U7982 (N_7982,N_6717,N_6607);
xor U7983 (N_7983,N_7184,N_6843);
and U7984 (N_7984,N_6677,N_7030);
nor U7985 (N_7985,N_6659,N_6516);
nand U7986 (N_7986,N_6188,N_6464);
nand U7987 (N_7987,N_6719,N_7113);
xor U7988 (N_7988,N_6704,N_6305);
nor U7989 (N_7989,N_6999,N_6658);
xor U7990 (N_7990,N_6278,N_6702);
or U7991 (N_7991,N_6073,N_6240);
xnor U7992 (N_7992,N_6079,N_6473);
xor U7993 (N_7993,N_6396,N_6947);
nor U7994 (N_7994,N_6984,N_6295);
or U7995 (N_7995,N_6434,N_6843);
xor U7996 (N_7996,N_7167,N_6402);
xnor U7997 (N_7997,N_6465,N_6748);
xnor U7998 (N_7998,N_6379,N_6166);
xor U7999 (N_7999,N_6387,N_6622);
xor U8000 (N_8000,N_6682,N_7019);
and U8001 (N_8001,N_7038,N_6697);
nand U8002 (N_8002,N_6565,N_6686);
nor U8003 (N_8003,N_6521,N_6499);
nor U8004 (N_8004,N_6306,N_6792);
xnor U8005 (N_8005,N_6900,N_6427);
nand U8006 (N_8006,N_6213,N_6168);
nand U8007 (N_8007,N_6763,N_6830);
nand U8008 (N_8008,N_6615,N_6280);
nor U8009 (N_8009,N_6801,N_6072);
nor U8010 (N_8010,N_6057,N_6273);
nand U8011 (N_8011,N_6118,N_7144);
nand U8012 (N_8012,N_6712,N_6940);
nor U8013 (N_8013,N_7157,N_6820);
xor U8014 (N_8014,N_6646,N_6526);
nor U8015 (N_8015,N_6340,N_7145);
nand U8016 (N_8016,N_6124,N_6606);
or U8017 (N_8017,N_6988,N_7054);
and U8018 (N_8018,N_6612,N_6758);
and U8019 (N_8019,N_6863,N_6173);
nand U8020 (N_8020,N_6487,N_6457);
xnor U8021 (N_8021,N_6154,N_7016);
xor U8022 (N_8022,N_6456,N_6681);
or U8023 (N_8023,N_6477,N_6489);
and U8024 (N_8024,N_6313,N_6493);
or U8025 (N_8025,N_6931,N_6187);
nand U8026 (N_8026,N_6534,N_7022);
or U8027 (N_8027,N_6225,N_6063);
xnor U8028 (N_8028,N_6937,N_6027);
nor U8029 (N_8029,N_6062,N_6559);
or U8030 (N_8030,N_6556,N_7158);
or U8031 (N_8031,N_6174,N_6283);
or U8032 (N_8032,N_7077,N_6962);
nor U8033 (N_8033,N_6068,N_6446);
nand U8034 (N_8034,N_6483,N_6697);
nand U8035 (N_8035,N_6747,N_6831);
nand U8036 (N_8036,N_6343,N_7046);
nor U8037 (N_8037,N_6152,N_6805);
xnor U8038 (N_8038,N_6183,N_6690);
xnor U8039 (N_8039,N_6385,N_6747);
nor U8040 (N_8040,N_6765,N_6443);
nor U8041 (N_8041,N_6408,N_6780);
nand U8042 (N_8042,N_6938,N_6557);
nand U8043 (N_8043,N_7037,N_6116);
xor U8044 (N_8044,N_7045,N_7024);
nor U8045 (N_8045,N_6715,N_6465);
nor U8046 (N_8046,N_6458,N_6584);
xor U8047 (N_8047,N_6889,N_6472);
xnor U8048 (N_8048,N_6705,N_6858);
nor U8049 (N_8049,N_6937,N_6910);
and U8050 (N_8050,N_6788,N_6398);
or U8051 (N_8051,N_6636,N_7097);
nand U8052 (N_8052,N_6371,N_7046);
and U8053 (N_8053,N_6361,N_6485);
and U8054 (N_8054,N_6914,N_6524);
nor U8055 (N_8055,N_7112,N_7139);
nand U8056 (N_8056,N_6944,N_7076);
nor U8057 (N_8057,N_7132,N_6990);
nor U8058 (N_8058,N_7197,N_6161);
nand U8059 (N_8059,N_6454,N_6240);
or U8060 (N_8060,N_6337,N_6925);
nand U8061 (N_8061,N_6902,N_6244);
nand U8062 (N_8062,N_6140,N_6811);
nor U8063 (N_8063,N_6041,N_6441);
xor U8064 (N_8064,N_6764,N_6415);
or U8065 (N_8065,N_6835,N_6492);
nor U8066 (N_8066,N_7018,N_7063);
xor U8067 (N_8067,N_6980,N_6047);
nand U8068 (N_8068,N_6598,N_6520);
and U8069 (N_8069,N_6762,N_6080);
or U8070 (N_8070,N_6357,N_6568);
or U8071 (N_8071,N_6050,N_6078);
or U8072 (N_8072,N_6374,N_6166);
xnor U8073 (N_8073,N_7046,N_7082);
nor U8074 (N_8074,N_6235,N_6312);
or U8075 (N_8075,N_6003,N_6859);
or U8076 (N_8076,N_6885,N_6510);
or U8077 (N_8077,N_6215,N_6847);
or U8078 (N_8078,N_7151,N_6360);
nor U8079 (N_8079,N_7170,N_6211);
nor U8080 (N_8080,N_6169,N_6988);
and U8081 (N_8081,N_6739,N_6745);
or U8082 (N_8082,N_6824,N_6633);
nand U8083 (N_8083,N_6301,N_6735);
or U8084 (N_8084,N_6502,N_6323);
nor U8085 (N_8085,N_6185,N_6971);
and U8086 (N_8086,N_6151,N_7092);
or U8087 (N_8087,N_6698,N_6024);
nand U8088 (N_8088,N_6292,N_6945);
nor U8089 (N_8089,N_6552,N_6958);
xnor U8090 (N_8090,N_6520,N_6089);
nand U8091 (N_8091,N_6842,N_6311);
nor U8092 (N_8092,N_7090,N_6573);
and U8093 (N_8093,N_6916,N_6321);
nor U8094 (N_8094,N_6303,N_7188);
nand U8095 (N_8095,N_6996,N_6549);
xor U8096 (N_8096,N_6968,N_6301);
nor U8097 (N_8097,N_6156,N_6693);
nand U8098 (N_8098,N_6632,N_6275);
or U8099 (N_8099,N_6452,N_7188);
nand U8100 (N_8100,N_7192,N_6800);
xor U8101 (N_8101,N_6131,N_6851);
nor U8102 (N_8102,N_6421,N_6003);
xor U8103 (N_8103,N_7002,N_6438);
and U8104 (N_8104,N_6971,N_6371);
or U8105 (N_8105,N_6047,N_6082);
or U8106 (N_8106,N_6759,N_6177);
and U8107 (N_8107,N_7037,N_6698);
nand U8108 (N_8108,N_6075,N_6479);
xnor U8109 (N_8109,N_6020,N_6754);
xnor U8110 (N_8110,N_6844,N_6471);
and U8111 (N_8111,N_6253,N_6797);
nand U8112 (N_8112,N_6038,N_6274);
xnor U8113 (N_8113,N_6202,N_6221);
xor U8114 (N_8114,N_6285,N_6386);
nor U8115 (N_8115,N_6841,N_6967);
or U8116 (N_8116,N_6048,N_6827);
nand U8117 (N_8117,N_7105,N_6952);
nand U8118 (N_8118,N_6745,N_6200);
xor U8119 (N_8119,N_6796,N_6688);
nor U8120 (N_8120,N_6001,N_6730);
xor U8121 (N_8121,N_6895,N_6027);
nor U8122 (N_8122,N_6514,N_7097);
nor U8123 (N_8123,N_6747,N_7159);
nand U8124 (N_8124,N_6244,N_6748);
nor U8125 (N_8125,N_6995,N_6118);
xor U8126 (N_8126,N_6936,N_6816);
or U8127 (N_8127,N_7017,N_6614);
or U8128 (N_8128,N_6291,N_6220);
nor U8129 (N_8129,N_6785,N_6181);
nand U8130 (N_8130,N_6312,N_6193);
and U8131 (N_8131,N_6612,N_6035);
xnor U8132 (N_8132,N_6813,N_7047);
nor U8133 (N_8133,N_6761,N_6780);
nor U8134 (N_8134,N_6195,N_6172);
nand U8135 (N_8135,N_6773,N_6481);
and U8136 (N_8136,N_6190,N_6769);
nor U8137 (N_8137,N_7113,N_7063);
xnor U8138 (N_8138,N_6137,N_6931);
nand U8139 (N_8139,N_6993,N_6248);
xnor U8140 (N_8140,N_6896,N_7095);
or U8141 (N_8141,N_6546,N_6319);
nand U8142 (N_8142,N_6862,N_6859);
and U8143 (N_8143,N_6832,N_6214);
nor U8144 (N_8144,N_6727,N_6166);
xnor U8145 (N_8145,N_7106,N_6358);
or U8146 (N_8146,N_6721,N_6928);
and U8147 (N_8147,N_7126,N_7059);
or U8148 (N_8148,N_6144,N_6598);
nand U8149 (N_8149,N_6940,N_6377);
xnor U8150 (N_8150,N_6121,N_6757);
nor U8151 (N_8151,N_6145,N_6916);
nor U8152 (N_8152,N_6906,N_6142);
or U8153 (N_8153,N_6888,N_6547);
and U8154 (N_8154,N_6350,N_7187);
nand U8155 (N_8155,N_6400,N_6751);
nor U8156 (N_8156,N_6983,N_6429);
and U8157 (N_8157,N_6407,N_7024);
or U8158 (N_8158,N_6873,N_6458);
and U8159 (N_8159,N_6718,N_6177);
nand U8160 (N_8160,N_6839,N_6008);
nor U8161 (N_8161,N_6157,N_7004);
nand U8162 (N_8162,N_6988,N_6175);
or U8163 (N_8163,N_6720,N_6894);
nand U8164 (N_8164,N_6693,N_7093);
or U8165 (N_8165,N_6372,N_7178);
nand U8166 (N_8166,N_7185,N_6713);
and U8167 (N_8167,N_6300,N_6711);
nand U8168 (N_8168,N_6164,N_6465);
nor U8169 (N_8169,N_6575,N_6632);
or U8170 (N_8170,N_6042,N_6786);
nand U8171 (N_8171,N_6271,N_6664);
xnor U8172 (N_8172,N_6158,N_6483);
nor U8173 (N_8173,N_6499,N_6964);
nor U8174 (N_8174,N_6879,N_6470);
nor U8175 (N_8175,N_6667,N_6789);
xor U8176 (N_8176,N_6678,N_6693);
and U8177 (N_8177,N_6080,N_7083);
nor U8178 (N_8178,N_7038,N_6015);
xor U8179 (N_8179,N_6494,N_7113);
xnor U8180 (N_8180,N_6417,N_6873);
nor U8181 (N_8181,N_6760,N_6179);
nor U8182 (N_8182,N_6921,N_6691);
nor U8183 (N_8183,N_6709,N_6371);
nand U8184 (N_8184,N_6106,N_6398);
and U8185 (N_8185,N_6116,N_6420);
and U8186 (N_8186,N_6606,N_6963);
and U8187 (N_8187,N_6638,N_6344);
xor U8188 (N_8188,N_6685,N_6650);
xnor U8189 (N_8189,N_7106,N_6295);
and U8190 (N_8190,N_6734,N_6482);
xor U8191 (N_8191,N_6686,N_6280);
nor U8192 (N_8192,N_6628,N_6532);
nor U8193 (N_8193,N_6254,N_6263);
nand U8194 (N_8194,N_6217,N_6120);
and U8195 (N_8195,N_7104,N_6040);
xnor U8196 (N_8196,N_6982,N_7096);
xor U8197 (N_8197,N_6533,N_6798);
or U8198 (N_8198,N_6821,N_6106);
nor U8199 (N_8199,N_7165,N_6032);
xnor U8200 (N_8200,N_6093,N_6841);
nor U8201 (N_8201,N_6040,N_6094);
nand U8202 (N_8202,N_7012,N_6969);
xnor U8203 (N_8203,N_6833,N_6547);
nor U8204 (N_8204,N_6094,N_6260);
and U8205 (N_8205,N_7180,N_6545);
nor U8206 (N_8206,N_6311,N_7157);
nor U8207 (N_8207,N_7025,N_6683);
or U8208 (N_8208,N_6605,N_6732);
nand U8209 (N_8209,N_6595,N_6755);
nor U8210 (N_8210,N_6649,N_6820);
nand U8211 (N_8211,N_6760,N_6966);
xor U8212 (N_8212,N_6108,N_6057);
xor U8213 (N_8213,N_6434,N_6480);
and U8214 (N_8214,N_6101,N_6027);
nand U8215 (N_8215,N_6932,N_6012);
nor U8216 (N_8216,N_6979,N_6168);
nand U8217 (N_8217,N_6148,N_7054);
xnor U8218 (N_8218,N_6412,N_6873);
and U8219 (N_8219,N_6669,N_7040);
nor U8220 (N_8220,N_6301,N_6063);
xnor U8221 (N_8221,N_6689,N_6336);
and U8222 (N_8222,N_6327,N_6618);
xnor U8223 (N_8223,N_6107,N_6764);
nand U8224 (N_8224,N_6327,N_6845);
and U8225 (N_8225,N_6034,N_6262);
nor U8226 (N_8226,N_6197,N_6440);
and U8227 (N_8227,N_6498,N_6670);
nor U8228 (N_8228,N_6264,N_6457);
xnor U8229 (N_8229,N_6307,N_6108);
or U8230 (N_8230,N_6979,N_6077);
nor U8231 (N_8231,N_6230,N_7191);
and U8232 (N_8232,N_6590,N_6839);
nor U8233 (N_8233,N_7121,N_6835);
and U8234 (N_8234,N_6433,N_6376);
nand U8235 (N_8235,N_7086,N_6927);
xnor U8236 (N_8236,N_7150,N_6353);
xnor U8237 (N_8237,N_6554,N_6088);
xor U8238 (N_8238,N_6424,N_6462);
or U8239 (N_8239,N_6878,N_6495);
or U8240 (N_8240,N_6384,N_6775);
xor U8241 (N_8241,N_6500,N_7012);
nand U8242 (N_8242,N_7080,N_6314);
or U8243 (N_8243,N_6977,N_6736);
xnor U8244 (N_8244,N_7182,N_6063);
and U8245 (N_8245,N_6835,N_6292);
nor U8246 (N_8246,N_6388,N_6351);
nand U8247 (N_8247,N_6500,N_6579);
and U8248 (N_8248,N_6506,N_6884);
nand U8249 (N_8249,N_6741,N_6037);
nor U8250 (N_8250,N_7182,N_6276);
xor U8251 (N_8251,N_6516,N_6661);
and U8252 (N_8252,N_6261,N_7038);
or U8253 (N_8253,N_7024,N_7117);
xnor U8254 (N_8254,N_6149,N_6731);
and U8255 (N_8255,N_6174,N_6032);
nand U8256 (N_8256,N_6208,N_6948);
xnor U8257 (N_8257,N_6429,N_6052);
or U8258 (N_8258,N_6008,N_6818);
or U8259 (N_8259,N_6922,N_6805);
or U8260 (N_8260,N_6149,N_7146);
or U8261 (N_8261,N_6983,N_6557);
nand U8262 (N_8262,N_6142,N_6984);
nand U8263 (N_8263,N_6968,N_6658);
or U8264 (N_8264,N_6598,N_6676);
nor U8265 (N_8265,N_7116,N_6471);
nor U8266 (N_8266,N_6748,N_6436);
nand U8267 (N_8267,N_7089,N_6709);
nand U8268 (N_8268,N_6066,N_6491);
nor U8269 (N_8269,N_6624,N_7103);
nor U8270 (N_8270,N_6346,N_6078);
and U8271 (N_8271,N_6794,N_6505);
xor U8272 (N_8272,N_6758,N_7075);
xnor U8273 (N_8273,N_7135,N_6144);
nor U8274 (N_8274,N_7164,N_6405);
nand U8275 (N_8275,N_6917,N_6541);
or U8276 (N_8276,N_6561,N_7092);
nand U8277 (N_8277,N_6642,N_6149);
and U8278 (N_8278,N_6398,N_6470);
and U8279 (N_8279,N_6689,N_7096);
and U8280 (N_8280,N_6710,N_6869);
nor U8281 (N_8281,N_6390,N_6061);
xnor U8282 (N_8282,N_7084,N_7015);
or U8283 (N_8283,N_6876,N_6133);
and U8284 (N_8284,N_6151,N_6915);
or U8285 (N_8285,N_6932,N_6196);
and U8286 (N_8286,N_6857,N_7044);
nor U8287 (N_8287,N_6342,N_6371);
nor U8288 (N_8288,N_6037,N_7016);
nand U8289 (N_8289,N_6713,N_6538);
xor U8290 (N_8290,N_6326,N_6661);
and U8291 (N_8291,N_6935,N_6845);
nor U8292 (N_8292,N_6405,N_6887);
nor U8293 (N_8293,N_6571,N_6414);
or U8294 (N_8294,N_6951,N_6985);
xor U8295 (N_8295,N_6823,N_6694);
nor U8296 (N_8296,N_7102,N_7082);
and U8297 (N_8297,N_6540,N_7016);
nand U8298 (N_8298,N_6863,N_6836);
or U8299 (N_8299,N_6031,N_6304);
and U8300 (N_8300,N_6650,N_6526);
xnor U8301 (N_8301,N_6540,N_6571);
or U8302 (N_8302,N_6317,N_6377);
nor U8303 (N_8303,N_6348,N_7112);
xor U8304 (N_8304,N_6953,N_6189);
xor U8305 (N_8305,N_6462,N_6819);
or U8306 (N_8306,N_6965,N_6005);
nor U8307 (N_8307,N_6414,N_7138);
nor U8308 (N_8308,N_6273,N_6963);
nor U8309 (N_8309,N_6994,N_6074);
or U8310 (N_8310,N_6382,N_6857);
and U8311 (N_8311,N_6140,N_7166);
xor U8312 (N_8312,N_6417,N_6624);
nand U8313 (N_8313,N_6762,N_6499);
nor U8314 (N_8314,N_6861,N_7180);
and U8315 (N_8315,N_7062,N_6298);
nor U8316 (N_8316,N_6008,N_7177);
or U8317 (N_8317,N_7019,N_6479);
or U8318 (N_8318,N_6404,N_6490);
nor U8319 (N_8319,N_6247,N_6745);
or U8320 (N_8320,N_6254,N_7033);
xor U8321 (N_8321,N_6314,N_6218);
nand U8322 (N_8322,N_7010,N_6634);
nand U8323 (N_8323,N_6304,N_6702);
nand U8324 (N_8324,N_7123,N_6617);
nor U8325 (N_8325,N_7168,N_6278);
nor U8326 (N_8326,N_6612,N_6570);
nand U8327 (N_8327,N_6417,N_6768);
nand U8328 (N_8328,N_6200,N_6207);
and U8329 (N_8329,N_7097,N_6574);
and U8330 (N_8330,N_6845,N_6285);
and U8331 (N_8331,N_6878,N_6579);
nor U8332 (N_8332,N_6675,N_6255);
nor U8333 (N_8333,N_6383,N_6825);
nor U8334 (N_8334,N_6851,N_6426);
nand U8335 (N_8335,N_6323,N_6186);
xnor U8336 (N_8336,N_6471,N_6494);
nand U8337 (N_8337,N_6412,N_6953);
nand U8338 (N_8338,N_6870,N_6675);
or U8339 (N_8339,N_7038,N_6240);
nor U8340 (N_8340,N_7011,N_6011);
nor U8341 (N_8341,N_6484,N_6771);
nor U8342 (N_8342,N_6546,N_6564);
nand U8343 (N_8343,N_6190,N_6097);
nand U8344 (N_8344,N_6587,N_6650);
and U8345 (N_8345,N_6159,N_6782);
nor U8346 (N_8346,N_6515,N_7035);
and U8347 (N_8347,N_6662,N_6774);
nor U8348 (N_8348,N_6921,N_6897);
nor U8349 (N_8349,N_6130,N_6876);
xor U8350 (N_8350,N_6913,N_6879);
xor U8351 (N_8351,N_6030,N_6117);
nand U8352 (N_8352,N_6168,N_7030);
nand U8353 (N_8353,N_6879,N_6729);
xor U8354 (N_8354,N_6602,N_6603);
nor U8355 (N_8355,N_6159,N_6337);
and U8356 (N_8356,N_6302,N_6352);
nor U8357 (N_8357,N_6314,N_6340);
or U8358 (N_8358,N_6998,N_6023);
nor U8359 (N_8359,N_6399,N_6291);
nand U8360 (N_8360,N_6611,N_6870);
and U8361 (N_8361,N_6870,N_7121);
nand U8362 (N_8362,N_7061,N_6630);
or U8363 (N_8363,N_6418,N_6976);
nand U8364 (N_8364,N_6699,N_6137);
and U8365 (N_8365,N_6935,N_6349);
or U8366 (N_8366,N_6868,N_6915);
nor U8367 (N_8367,N_7140,N_7080);
nor U8368 (N_8368,N_6351,N_6532);
nand U8369 (N_8369,N_6542,N_6571);
and U8370 (N_8370,N_6423,N_6697);
xor U8371 (N_8371,N_7157,N_6462);
or U8372 (N_8372,N_6830,N_6636);
or U8373 (N_8373,N_6736,N_6768);
and U8374 (N_8374,N_6732,N_6209);
nand U8375 (N_8375,N_6546,N_7045);
or U8376 (N_8376,N_6646,N_6764);
and U8377 (N_8377,N_6539,N_6939);
or U8378 (N_8378,N_6272,N_6698);
nand U8379 (N_8379,N_6151,N_6491);
or U8380 (N_8380,N_6668,N_6580);
or U8381 (N_8381,N_6133,N_6697);
or U8382 (N_8382,N_7141,N_6849);
xnor U8383 (N_8383,N_6646,N_6737);
xor U8384 (N_8384,N_7053,N_6763);
nand U8385 (N_8385,N_6926,N_7172);
nor U8386 (N_8386,N_6452,N_6018);
and U8387 (N_8387,N_6172,N_6184);
nor U8388 (N_8388,N_6016,N_7044);
or U8389 (N_8389,N_7194,N_6595);
nand U8390 (N_8390,N_7021,N_6834);
xnor U8391 (N_8391,N_6890,N_7177);
or U8392 (N_8392,N_6816,N_6085);
or U8393 (N_8393,N_6749,N_6507);
or U8394 (N_8394,N_6739,N_6135);
or U8395 (N_8395,N_6562,N_6871);
xor U8396 (N_8396,N_6339,N_6267);
or U8397 (N_8397,N_6451,N_7079);
nand U8398 (N_8398,N_7134,N_6411);
nor U8399 (N_8399,N_6021,N_6077);
and U8400 (N_8400,N_8157,N_7882);
nor U8401 (N_8401,N_7300,N_7989);
nand U8402 (N_8402,N_8240,N_8279);
xor U8403 (N_8403,N_7668,N_7879);
nor U8404 (N_8404,N_7485,N_8128);
and U8405 (N_8405,N_7975,N_7517);
xor U8406 (N_8406,N_7673,N_7527);
nor U8407 (N_8407,N_7672,N_8310);
and U8408 (N_8408,N_7738,N_7963);
or U8409 (N_8409,N_8189,N_8258);
nand U8410 (N_8410,N_7413,N_8174);
nor U8411 (N_8411,N_7640,N_8382);
nor U8412 (N_8412,N_7727,N_7752);
nor U8413 (N_8413,N_7506,N_7716);
nor U8414 (N_8414,N_7741,N_7750);
and U8415 (N_8415,N_8156,N_8251);
nand U8416 (N_8416,N_8350,N_7979);
or U8417 (N_8417,N_8160,N_8322);
or U8418 (N_8418,N_7575,N_8390);
or U8419 (N_8419,N_7595,N_7617);
nand U8420 (N_8420,N_7410,N_7837);
nand U8421 (N_8421,N_8264,N_7941);
xnor U8422 (N_8422,N_7256,N_7731);
and U8423 (N_8423,N_8301,N_7491);
and U8424 (N_8424,N_7743,N_7625);
nand U8425 (N_8425,N_7960,N_7890);
and U8426 (N_8426,N_7684,N_7859);
nand U8427 (N_8427,N_7510,N_7739);
and U8428 (N_8428,N_8152,N_7224);
xnor U8429 (N_8429,N_8176,N_8125);
nand U8430 (N_8430,N_8141,N_7481);
and U8431 (N_8431,N_8126,N_7223);
and U8432 (N_8432,N_7862,N_7714);
and U8433 (N_8433,N_7677,N_7993);
or U8434 (N_8434,N_7982,N_8150);
xor U8435 (N_8435,N_8120,N_8203);
nor U8436 (N_8436,N_7277,N_7965);
nand U8437 (N_8437,N_7285,N_7393);
nand U8438 (N_8438,N_7480,N_7292);
xor U8439 (N_8439,N_7220,N_7729);
or U8440 (N_8440,N_7608,N_8079);
xor U8441 (N_8441,N_7639,N_8099);
or U8442 (N_8442,N_8042,N_8341);
or U8443 (N_8443,N_7458,N_7453);
xnor U8444 (N_8444,N_8393,N_7650);
or U8445 (N_8445,N_7351,N_8065);
nor U8446 (N_8446,N_7665,N_7459);
nor U8447 (N_8447,N_7851,N_7400);
nand U8448 (N_8448,N_8223,N_7935);
nor U8449 (N_8449,N_7922,N_7991);
xor U8450 (N_8450,N_7662,N_8167);
nand U8451 (N_8451,N_7253,N_7611);
or U8452 (N_8452,N_7572,N_8312);
or U8453 (N_8453,N_7386,N_7726);
xnor U8454 (N_8454,N_7217,N_7498);
or U8455 (N_8455,N_7787,N_7892);
or U8456 (N_8456,N_8387,N_7471);
and U8457 (N_8457,N_8324,N_8013);
or U8458 (N_8458,N_8211,N_7556);
nand U8459 (N_8459,N_8031,N_7915);
nor U8460 (N_8460,N_7544,N_7775);
nand U8461 (N_8461,N_7380,N_7298);
or U8462 (N_8462,N_8355,N_8235);
and U8463 (N_8463,N_7293,N_7371);
nand U8464 (N_8464,N_7767,N_8139);
or U8465 (N_8465,N_8329,N_8164);
nor U8466 (N_8466,N_7692,N_7748);
and U8467 (N_8467,N_8015,N_8082);
nand U8468 (N_8468,N_8038,N_7440);
nand U8469 (N_8469,N_7985,N_8366);
and U8470 (N_8470,N_7387,N_8093);
or U8471 (N_8471,N_7609,N_7992);
xor U8472 (N_8472,N_7463,N_7315);
nand U8473 (N_8473,N_7833,N_8045);
xor U8474 (N_8474,N_7768,N_8311);
xnor U8475 (N_8475,N_7389,N_7344);
nand U8476 (N_8476,N_7549,N_7377);
nand U8477 (N_8477,N_7824,N_7274);
xor U8478 (N_8478,N_8179,N_8004);
nand U8479 (N_8479,N_7822,N_7327);
nand U8480 (N_8480,N_7412,N_8121);
xor U8481 (N_8481,N_8106,N_8232);
or U8482 (N_8482,N_7596,N_7206);
or U8483 (N_8483,N_7853,N_7318);
xor U8484 (N_8484,N_8025,N_8231);
or U8485 (N_8485,N_7845,N_7808);
or U8486 (N_8486,N_7202,N_8057);
xnor U8487 (N_8487,N_8305,N_8105);
nand U8488 (N_8488,N_8165,N_7350);
nand U8489 (N_8489,N_7500,N_7209);
nor U8490 (N_8490,N_8347,N_8196);
nor U8491 (N_8491,N_7604,N_7426);
nor U8492 (N_8492,N_7267,N_7854);
or U8493 (N_8493,N_8263,N_7411);
and U8494 (N_8494,N_7999,N_7683);
xnor U8495 (N_8495,N_7632,N_8010);
nor U8496 (N_8496,N_7693,N_7492);
or U8497 (N_8497,N_7995,N_7434);
and U8498 (N_8498,N_7273,N_7319);
xnor U8499 (N_8499,N_8171,N_7580);
and U8500 (N_8500,N_7359,N_7964);
xnor U8501 (N_8501,N_7573,N_7669);
nor U8502 (N_8502,N_8351,N_7836);
and U8503 (N_8503,N_7521,N_7357);
and U8504 (N_8504,N_8396,N_7353);
and U8505 (N_8505,N_7981,N_7241);
and U8506 (N_8506,N_7718,N_7687);
and U8507 (N_8507,N_8313,N_7366);
nor U8508 (N_8508,N_7451,N_7231);
nand U8509 (N_8509,N_7844,N_7303);
nor U8510 (N_8510,N_7652,N_8172);
nor U8511 (N_8511,N_7997,N_7712);
or U8512 (N_8512,N_7637,N_8256);
or U8513 (N_8513,N_8084,N_7244);
nor U8514 (N_8514,N_8288,N_7372);
or U8515 (N_8515,N_7381,N_7467);
xnor U8516 (N_8516,N_7832,N_7947);
nand U8517 (N_8517,N_7487,N_8083);
nor U8518 (N_8518,N_8208,N_7801);
xnor U8519 (N_8519,N_7899,N_7616);
and U8520 (N_8520,N_7555,N_8257);
xnor U8521 (N_8521,N_8289,N_8384);
or U8522 (N_8522,N_7259,N_7666);
and U8523 (N_8523,N_7651,N_7419);
and U8524 (N_8524,N_7403,N_8186);
xnor U8525 (N_8525,N_8369,N_8249);
and U8526 (N_8526,N_8006,N_7405);
or U8527 (N_8527,N_7522,N_8202);
and U8528 (N_8528,N_7382,N_7682);
nor U8529 (N_8529,N_7933,N_7793);
nand U8530 (N_8530,N_7321,N_7430);
and U8531 (N_8531,N_7856,N_7855);
nor U8532 (N_8532,N_7499,N_8229);
or U8533 (N_8533,N_7258,N_7326);
nand U8534 (N_8534,N_7635,N_7399);
or U8535 (N_8535,N_7356,N_8124);
nor U8536 (N_8536,N_8051,N_7501);
nand U8537 (N_8537,N_8030,N_7628);
or U8538 (N_8538,N_7479,N_8261);
nand U8539 (N_8539,N_7802,N_8236);
nand U8540 (N_8540,N_8303,N_7333);
or U8541 (N_8541,N_8153,N_8033);
nand U8542 (N_8542,N_7653,N_8335);
and U8543 (N_8543,N_8380,N_7641);
and U8544 (N_8544,N_7566,N_7810);
or U8545 (N_8545,N_7656,N_7654);
and U8546 (N_8546,N_7972,N_7532);
or U8547 (N_8547,N_7804,N_7423);
and U8548 (N_8548,N_8209,N_7661);
or U8549 (N_8549,N_7309,N_7286);
xor U8550 (N_8550,N_7539,N_7762);
xor U8551 (N_8551,N_7618,N_7870);
and U8552 (N_8552,N_7817,N_7944);
or U8553 (N_8553,N_7374,N_7331);
and U8554 (N_8554,N_7983,N_7547);
or U8555 (N_8555,N_7397,N_8195);
nor U8556 (N_8556,N_8358,N_8021);
nand U8557 (N_8557,N_7663,N_8316);
nor U8558 (N_8558,N_8060,N_8286);
nor U8559 (N_8559,N_7961,N_8277);
and U8560 (N_8560,N_8241,N_7959);
and U8561 (N_8561,N_8163,N_7408);
xor U8562 (N_8562,N_8048,N_7452);
nand U8563 (N_8563,N_8177,N_7424);
xnor U8564 (N_8564,N_7676,N_7446);
nor U8565 (N_8565,N_7365,N_7866);
and U8566 (N_8566,N_8294,N_8337);
or U8567 (N_8567,N_8326,N_7358);
nand U8568 (N_8568,N_7534,N_7520);
and U8569 (N_8569,N_7841,N_8087);
xnor U8570 (N_8570,N_7790,N_8035);
or U8571 (N_8571,N_8242,N_7347);
and U8572 (N_8572,N_8295,N_7585);
and U8573 (N_8573,N_7928,N_7966);
xor U8574 (N_8574,N_7305,N_8199);
nor U8575 (N_8575,N_7805,N_8067);
and U8576 (N_8576,N_7232,N_8017);
nand U8577 (N_8577,N_8331,N_8377);
nand U8578 (N_8578,N_8091,N_8169);
and U8579 (N_8579,N_7690,N_7378);
nand U8580 (N_8580,N_8161,N_7494);
nand U8581 (N_8581,N_7913,N_7807);
and U8582 (N_8582,N_8207,N_7296);
and U8583 (N_8583,N_7230,N_7987);
xor U8584 (N_8584,N_8246,N_8282);
nor U8585 (N_8585,N_7766,N_7794);
nand U8586 (N_8586,N_7770,N_8044);
or U8587 (N_8587,N_7717,N_7934);
nand U8588 (N_8588,N_8395,N_7797);
nand U8589 (N_8589,N_7986,N_7897);
or U8590 (N_8590,N_8287,N_8039);
nand U8591 (N_8591,N_7428,N_7936);
xnor U8592 (N_8592,N_7763,N_7704);
nor U8593 (N_8593,N_7222,N_7850);
xnor U8594 (N_8594,N_7212,N_7774);
nand U8595 (N_8595,N_7307,N_8354);
nor U8596 (N_8596,N_7869,N_7324);
or U8597 (N_8597,N_8088,N_7427);
xor U8598 (N_8598,N_7421,N_7251);
nor U8599 (N_8599,N_7877,N_7953);
xnor U8600 (N_8600,N_7476,N_7660);
xor U8601 (N_8601,N_7962,N_8255);
nand U8602 (N_8602,N_7917,N_8389);
xnor U8603 (N_8603,N_7278,N_7671);
nor U8604 (N_8604,N_7881,N_7831);
or U8605 (N_8605,N_7984,N_8233);
or U8606 (N_8606,N_7215,N_7271);
nand U8607 (N_8607,N_7415,N_8108);
nand U8608 (N_8608,N_7391,N_7893);
or U8609 (N_8609,N_8193,N_8367);
nor U8610 (N_8610,N_7889,N_7239);
nand U8611 (N_8611,N_7394,N_7624);
xor U8612 (N_8612,N_8080,N_8103);
or U8613 (N_8613,N_7909,N_7312);
xor U8614 (N_8614,N_8302,N_7569);
or U8615 (N_8615,N_8224,N_8388);
xnor U8616 (N_8616,N_7896,N_8012);
nand U8617 (N_8617,N_7644,N_8143);
or U8618 (N_8618,N_8119,N_7310);
nor U8619 (N_8619,N_8370,N_7468);
xnor U8620 (N_8620,N_8053,N_8063);
nand U8621 (N_8621,N_7756,N_8359);
or U8622 (N_8622,N_7858,N_7228);
or U8623 (N_8623,N_7249,N_7875);
and U8624 (N_8624,N_8398,N_7830);
nand U8625 (N_8625,N_7254,N_7543);
or U8626 (N_8626,N_8373,N_7425);
nand U8627 (N_8627,N_8011,N_7723);
nand U8628 (N_8628,N_7606,N_7670);
nand U8629 (N_8629,N_7871,N_8348);
or U8630 (N_8630,N_7819,N_7342);
and U8631 (N_8631,N_8149,N_7279);
and U8632 (N_8632,N_7289,N_7433);
nand U8633 (N_8633,N_7779,N_7436);
and U8634 (N_8634,N_7681,N_7200);
or U8635 (N_8635,N_8187,N_7548);
or U8636 (N_8636,N_7355,N_8096);
and U8637 (N_8637,N_7218,N_7269);
nand U8638 (N_8638,N_7942,N_7316);
and U8639 (N_8639,N_8345,N_8397);
or U8640 (N_8640,N_7950,N_7708);
or U8641 (N_8641,N_7806,N_8325);
and U8642 (N_8642,N_7559,N_7753);
nand U8643 (N_8643,N_8361,N_8375);
or U8644 (N_8644,N_7786,N_7929);
and U8645 (N_8645,N_7773,N_8314);
and U8646 (N_8646,N_7634,N_7973);
nand U8647 (N_8647,N_7646,N_7335);
or U8648 (N_8648,N_7345,N_8221);
or U8649 (N_8649,N_7435,N_8151);
and U8650 (N_8650,N_8001,N_7449);
or U8651 (N_8651,N_8297,N_7484);
nand U8652 (N_8652,N_7329,N_7633);
nand U8653 (N_8653,N_7605,N_8266);
or U8654 (N_8654,N_8107,N_7238);
nor U8655 (N_8655,N_8175,N_7516);
and U8656 (N_8656,N_7225,N_7341);
nand U8657 (N_8657,N_8173,N_8116);
or U8658 (N_8658,N_7582,N_8320);
or U8659 (N_8659,N_7838,N_7313);
or U8660 (N_8660,N_7593,N_8131);
nor U8661 (N_8661,N_8058,N_8034);
xnor U8662 (N_8662,N_8123,N_7242);
and U8663 (N_8663,N_7620,N_7343);
or U8664 (N_8664,N_7323,N_8159);
xor U8665 (N_8665,N_7328,N_7322);
xnor U8666 (N_8666,N_7957,N_8009);
or U8667 (N_8667,N_7252,N_7867);
nand U8668 (N_8668,N_8356,N_7615);
or U8669 (N_8669,N_7907,N_7648);
or U8670 (N_8670,N_8378,N_8029);
and U8671 (N_8671,N_8027,N_8285);
xor U8672 (N_8672,N_8309,N_7769);
nand U8673 (N_8673,N_7416,N_7940);
or U8674 (N_8674,N_8270,N_7619);
and U8675 (N_8675,N_7562,N_7336);
and U8676 (N_8676,N_7664,N_7900);
or U8677 (N_8677,N_7812,N_8075);
and U8678 (N_8678,N_7974,N_7234);
and U8679 (N_8679,N_7519,N_7542);
nor U8680 (N_8680,N_7864,N_8391);
or U8681 (N_8681,N_7280,N_7706);
and U8682 (N_8682,N_8142,N_8210);
or U8683 (N_8683,N_8333,N_7658);
nor U8684 (N_8684,N_7747,N_8147);
xnor U8685 (N_8685,N_8098,N_7332);
nand U8686 (N_8686,N_7969,N_8214);
xor U8687 (N_8687,N_8008,N_8228);
nand U8688 (N_8688,N_7771,N_7496);
and U8689 (N_8689,N_7590,N_8267);
and U8690 (N_8690,N_7887,N_7948);
xnor U8691 (N_8691,N_7270,N_8360);
or U8692 (N_8692,N_7919,N_7998);
nor U8693 (N_8693,N_7667,N_7297);
nor U8694 (N_8694,N_8217,N_7594);
xor U8695 (N_8695,N_7592,N_7514);
and U8696 (N_8696,N_8336,N_7375);
nand U8697 (N_8697,N_7438,N_7368);
and U8698 (N_8698,N_8061,N_7884);
or U8699 (N_8699,N_7733,N_7803);
or U8700 (N_8700,N_8100,N_7735);
xor U8701 (N_8701,N_7441,N_8050);
nand U8702 (N_8702,N_8024,N_8275);
xnor U8703 (N_8703,N_8086,N_7840);
nor U8704 (N_8704,N_8113,N_7390);
nor U8705 (N_8705,N_8074,N_8197);
or U8706 (N_8706,N_8014,N_7287);
and U8707 (N_8707,N_7246,N_7587);
and U8708 (N_8708,N_7724,N_7795);
nand U8709 (N_8709,N_7465,N_7788);
nor U8710 (N_8710,N_7570,N_8299);
or U8711 (N_8711,N_8317,N_8111);
nor U8712 (N_8712,N_8104,N_8268);
and U8713 (N_8713,N_8291,N_8192);
xor U8714 (N_8714,N_8332,N_8026);
and U8715 (N_8715,N_7630,N_7623);
and U8716 (N_8716,N_8115,N_8056);
nor U8717 (N_8717,N_7291,N_8290);
nor U8718 (N_8718,N_7227,N_8122);
or U8719 (N_8719,N_7385,N_8168);
nor U8720 (N_8720,N_7709,N_7931);
xor U8721 (N_8721,N_7749,N_7588);
xnor U8722 (N_8722,N_8078,N_7814);
xnor U8723 (N_8723,N_8304,N_8368);
nor U8724 (N_8724,N_8158,N_7951);
and U8725 (N_8725,N_7742,N_8054);
nand U8726 (N_8726,N_7925,N_7809);
nor U8727 (N_8727,N_7707,N_7406);
nand U8728 (N_8728,N_7655,N_7571);
or U8729 (N_8729,N_8040,N_7848);
nand U8730 (N_8730,N_7533,N_8260);
xnor U8731 (N_8731,N_7317,N_7949);
nand U8732 (N_8732,N_8308,N_7906);
nor U8733 (N_8733,N_7388,N_7872);
xor U8734 (N_8734,N_7777,N_8298);
and U8735 (N_8735,N_7462,N_7885);
nor U8736 (N_8736,N_7376,N_7861);
xnor U8737 (N_8737,N_7778,N_8385);
nand U8738 (N_8738,N_8095,N_7579);
nand U8739 (N_8739,N_8130,N_7761);
nand U8740 (N_8740,N_7923,N_8182);
nor U8741 (N_8741,N_7976,N_8253);
or U8742 (N_8742,N_8138,N_7488);
and U8743 (N_8743,N_7700,N_8049);
nor U8744 (N_8744,N_7364,N_7203);
or U8745 (N_8745,N_7395,N_8399);
or U8746 (N_8746,N_7612,N_7629);
nand U8747 (N_8747,N_8059,N_7214);
nor U8748 (N_8748,N_7338,N_8016);
nor U8749 (N_8749,N_7715,N_7711);
nor U8750 (N_8750,N_8372,N_7880);
or U8751 (N_8751,N_7988,N_7938);
xor U8752 (N_8752,N_7243,N_8181);
or U8753 (N_8753,N_7847,N_8386);
nand U8754 (N_8754,N_8023,N_8133);
xor U8755 (N_8755,N_7455,N_7247);
nand U8756 (N_8756,N_7791,N_8135);
nand U8757 (N_8757,N_8318,N_7493);
and U8758 (N_8758,N_7509,N_8218);
xor U8759 (N_8759,N_8072,N_8041);
and U8760 (N_8760,N_8248,N_8283);
or U8761 (N_8761,N_7578,N_7829);
xor U8762 (N_8762,N_7583,N_7396);
and U8763 (N_8763,N_7545,N_7523);
xnor U8764 (N_8764,N_7815,N_7828);
xnor U8765 (N_8765,N_7221,N_7260);
nand U8766 (N_8766,N_8306,N_8005);
nand U8767 (N_8767,N_8137,N_8145);
nor U8768 (N_8768,N_8328,N_8191);
xnor U8769 (N_8769,N_8018,N_7736);
nand U8770 (N_8770,N_8259,N_7529);
nor U8771 (N_8771,N_7448,N_7603);
nand U8772 (N_8772,N_7910,N_7264);
nand U8773 (N_8773,N_7302,N_7237);
nand U8774 (N_8774,N_7407,N_8076);
xnor U8775 (N_8775,N_7402,N_7505);
nand U8776 (N_8776,N_7235,N_7820);
nor U8777 (N_8777,N_7903,N_7626);
or U8778 (N_8778,N_7538,N_8206);
and U8779 (N_8779,N_7621,N_7703);
nand U8780 (N_8780,N_7956,N_8178);
or U8781 (N_8781,N_7930,N_8109);
or U8782 (N_8782,N_7272,N_8374);
or U8783 (N_8783,N_7213,N_7306);
or U8784 (N_8784,N_8247,N_8227);
or U8785 (N_8785,N_7461,N_8300);
or U8786 (N_8786,N_7314,N_7834);
or U8787 (N_8787,N_8272,N_7207);
xnor U8788 (N_8788,N_7883,N_7721);
and U8789 (N_8789,N_8352,N_7508);
or U8790 (N_8790,N_7912,N_7567);
and U8791 (N_8791,N_7240,N_7905);
and U8792 (N_8792,N_8327,N_8239);
nor U8793 (N_8793,N_7373,N_7362);
nor U8794 (N_8794,N_7211,N_8047);
or U8795 (N_8795,N_7486,N_8225);
nor U8796 (N_8796,N_8117,N_7927);
and U8797 (N_8797,N_7755,N_7210);
xnor U8798 (N_8798,N_7489,N_8296);
or U8799 (N_8799,N_7383,N_8069);
nor U8800 (N_8800,N_8180,N_7865);
nand U8801 (N_8801,N_7937,N_7918);
or U8802 (N_8802,N_8201,N_8371);
and U8803 (N_8803,N_8343,N_7996);
xnor U8804 (N_8804,N_8140,N_7340);
nor U8805 (N_8805,N_7698,N_7443);
and U8806 (N_8806,N_7414,N_7524);
or U8807 (N_8807,N_7781,N_7800);
or U8808 (N_8808,N_8043,N_8129);
and U8809 (N_8809,N_7601,N_7908);
nand U8810 (N_8810,N_7638,N_7361);
and U8811 (N_8811,N_7914,N_8362);
and U8812 (N_8812,N_7873,N_7924);
nor U8813 (N_8813,N_8066,N_7561);
xnor U8814 (N_8814,N_7901,N_7622);
nand U8815 (N_8815,N_8319,N_7921);
nand U8816 (N_8816,N_7835,N_7857);
or U8817 (N_8817,N_7442,N_7557);
nor U8818 (N_8818,N_7584,N_7248);
nand U8819 (N_8819,N_7275,N_8219);
or U8820 (N_8820,N_7888,N_8307);
and U8821 (N_8821,N_8346,N_8344);
and U8822 (N_8822,N_7728,N_8323);
or U8823 (N_8823,N_7348,N_7849);
nand U8824 (N_8824,N_8220,N_7600);
or U8825 (N_8825,N_7472,N_8090);
nor U8826 (N_8826,N_8365,N_7229);
nand U8827 (N_8827,N_8278,N_7284);
and U8828 (N_8828,N_8020,N_7450);
nor U8829 (N_8829,N_8073,N_7591);
xor U8830 (N_8830,N_7299,N_8185);
nand U8831 (N_8831,N_8146,N_8349);
nand U8832 (N_8832,N_7325,N_7874);
or U8833 (N_8833,N_7311,N_7552);
nor U8834 (N_8834,N_8215,N_7418);
nor U8835 (N_8835,N_7818,N_7261);
nor U8836 (N_8836,N_8068,N_7422);
nand U8837 (N_8837,N_8132,N_8244);
or U8838 (N_8838,N_8281,N_7971);
nor U8839 (N_8839,N_7478,N_7432);
or U8840 (N_8840,N_8166,N_8071);
xor U8841 (N_8841,N_7643,N_7863);
or U8842 (N_8842,N_8237,N_7751);
xnor U8843 (N_8843,N_7504,N_7429);
xnor U8844 (N_8844,N_7515,N_8170);
or U8845 (N_8845,N_8102,N_8245);
nand U8846 (N_8846,N_7689,N_8230);
or U8847 (N_8847,N_7645,N_7868);
nor U8848 (N_8848,N_8226,N_7958);
nor U8849 (N_8849,N_7282,N_7551);
nand U8850 (N_8850,N_8064,N_7233);
nor U8851 (N_8851,N_7464,N_7695);
xnor U8852 (N_8852,N_8338,N_7379);
or U8853 (N_8853,N_7691,N_7782);
xnor U8854 (N_8854,N_7688,N_7477);
and U8855 (N_8855,N_7852,N_7546);
xnor U8856 (N_8856,N_7226,N_7553);
nor U8857 (N_8857,N_7334,N_7697);
and U8858 (N_8858,N_7466,N_7554);
nor U8859 (N_8859,N_8110,N_7565);
and U8860 (N_8860,N_8002,N_7740);
nand U8861 (N_8861,N_8155,N_8037);
nor U8862 (N_8862,N_7642,N_7758);
or U8863 (N_8863,N_7990,N_7401);
or U8864 (N_8864,N_7843,N_7970);
and U8865 (N_8865,N_7507,N_7276);
xor U8866 (N_8866,N_7649,N_7470);
nand U8867 (N_8867,N_7685,N_7456);
nor U8868 (N_8868,N_7431,N_8055);
or U8869 (N_8869,N_7916,N_8212);
xor U8870 (N_8870,N_7977,N_7876);
or U8871 (N_8871,N_7980,N_7512);
xnor U8872 (N_8872,N_7513,N_8250);
and U8873 (N_8873,N_8077,N_7370);
and U8874 (N_8874,N_7911,N_8340);
xnor U8875 (N_8875,N_7878,N_7445);
and U8876 (N_8876,N_7827,N_7636);
nor U8877 (N_8877,N_7201,N_8046);
nand U8878 (N_8878,N_7541,N_7262);
nand U8879 (N_8879,N_8234,N_7659);
nor U8880 (N_8880,N_7776,N_7497);
and U8881 (N_8881,N_7994,N_7398);
xor U8882 (N_8882,N_7564,N_7540);
nand U8883 (N_8883,N_8273,N_8154);
xor U8884 (N_8884,N_7745,N_7764);
nand U8885 (N_8885,N_7360,N_8383);
and U8886 (N_8886,N_7265,N_8032);
nand U8887 (N_8887,N_8238,N_7257);
or U8888 (N_8888,N_7586,N_7288);
nand U8889 (N_8889,N_7531,N_7528);
nor U8890 (N_8890,N_7895,N_7263);
xnor U8891 (N_8891,N_8028,N_7503);
xnor U8892 (N_8892,N_7967,N_7204);
and U8893 (N_8893,N_7589,N_7679);
and U8894 (N_8894,N_7789,N_8184);
nor U8895 (N_8895,N_7576,N_7730);
nand U8896 (N_8896,N_8134,N_7320);
xnor U8897 (N_8897,N_7337,N_8144);
nor U8898 (N_8898,N_7657,N_8022);
xnor U8899 (N_8899,N_7473,N_8162);
xnor U8900 (N_8900,N_8292,N_8003);
xnor U8901 (N_8901,N_7613,N_7417);
nor U8902 (N_8902,N_8204,N_7354);
or U8903 (N_8903,N_7784,N_8097);
xnor U8904 (N_8904,N_7290,N_7563);
or U8905 (N_8905,N_7346,N_7255);
nand U8906 (N_8906,N_7475,N_7208);
and U8907 (N_8907,N_7369,N_7250);
xnor U8908 (N_8908,N_7886,N_7439);
xor U8909 (N_8909,N_8254,N_7483);
nand U8910 (N_8910,N_7686,N_8200);
or U8911 (N_8911,N_7558,N_7602);
xnor U8912 (N_8912,N_7469,N_7511);
or U8913 (N_8913,N_8284,N_8315);
nor U8914 (N_8914,N_7607,N_7631);
xor U8915 (N_8915,N_7839,N_7610);
nand U8916 (N_8916,N_7339,N_7367);
nand U8917 (N_8917,N_7783,N_8276);
or U8918 (N_8918,N_7447,N_8293);
or U8919 (N_8919,N_7955,N_8357);
nor U8920 (N_8920,N_7785,N_8007);
nand U8921 (N_8921,N_7550,N_7295);
xnor U8922 (N_8922,N_7943,N_8000);
and U8923 (N_8923,N_7826,N_7813);
nor U8924 (N_8924,N_7811,N_8280);
nand U8925 (N_8925,N_8089,N_7978);
nand U8926 (N_8926,N_7760,N_7454);
nand U8927 (N_8927,N_8274,N_7474);
nand U8928 (N_8928,N_8222,N_7725);
nor U8929 (N_8929,N_7678,N_7349);
xnor U8930 (N_8930,N_7409,N_7308);
nand U8931 (N_8931,N_7574,N_7392);
xor U8932 (N_8932,N_8243,N_7710);
and U8933 (N_8933,N_8085,N_8190);
nor U8934 (N_8934,N_7902,N_8376);
nor U8935 (N_8935,N_8183,N_7535);
nand U8936 (N_8936,N_8052,N_8334);
or U8937 (N_8937,N_7823,N_7599);
or U8938 (N_8938,N_8019,N_8364);
nand U8939 (N_8939,N_8271,N_7537);
nand U8940 (N_8940,N_8036,N_7894);
and U8941 (N_8941,N_7536,N_7495);
and U8942 (N_8942,N_8394,N_7699);
nand U8943 (N_8943,N_7568,N_7860);
xnor U8944 (N_8944,N_7744,N_7798);
nand U8945 (N_8945,N_7437,N_7420);
xnor U8946 (N_8946,N_7920,N_7680);
or U8947 (N_8947,N_7846,N_8114);
xnor U8948 (N_8948,N_7737,N_8198);
nand U8949 (N_8949,N_8213,N_7330);
xor U8950 (N_8950,N_8262,N_8188);
and U8951 (N_8951,N_7713,N_7352);
nand U8952 (N_8952,N_7842,N_7939);
and U8953 (N_8953,N_7825,N_7754);
or U8954 (N_8954,N_7266,N_7746);
or U8955 (N_8955,N_7301,N_7560);
and U8956 (N_8956,N_7722,N_8148);
nor U8957 (N_8957,N_7674,N_7799);
or U8958 (N_8958,N_7926,N_8205);
or U8959 (N_8959,N_7792,N_7968);
or U8960 (N_8960,N_7719,N_7702);
or U8961 (N_8961,N_7780,N_8342);
and U8962 (N_8962,N_7821,N_7757);
and U8963 (N_8963,N_8339,N_7205);
nor U8964 (N_8964,N_8321,N_7216);
nor U8965 (N_8965,N_8094,N_8216);
nor U8966 (N_8966,N_7363,N_8062);
nor U8967 (N_8967,N_8265,N_8194);
and U8968 (N_8968,N_7732,N_8252);
nand U8969 (N_8969,N_8118,N_7696);
nor U8970 (N_8970,N_7675,N_7236);
and U8971 (N_8971,N_7772,N_7759);
and U8972 (N_8972,N_8127,N_7898);
nor U8973 (N_8973,N_8136,N_7518);
and U8974 (N_8974,N_7701,N_7281);
and U8975 (N_8975,N_8269,N_7904);
xor U8976 (N_8976,N_7304,N_7457);
or U8977 (N_8977,N_7384,N_8392);
nand U8978 (N_8978,N_8081,N_7720);
nand U8979 (N_8979,N_8092,N_7765);
or U8980 (N_8980,N_7816,N_7891);
and U8981 (N_8981,N_7526,N_7490);
nor U8982 (N_8982,N_7245,N_7952);
xor U8983 (N_8983,N_8112,N_7268);
and U8984 (N_8984,N_7647,N_7734);
xnor U8985 (N_8985,N_8381,N_7614);
and U8986 (N_8986,N_7460,N_7482);
nor U8987 (N_8987,N_7444,N_7694);
nor U8988 (N_8988,N_8363,N_7577);
and U8989 (N_8989,N_7525,N_8070);
or U8990 (N_8990,N_8101,N_7294);
and U8991 (N_8991,N_7796,N_7283);
xor U8992 (N_8992,N_7502,N_7219);
nand U8993 (N_8993,N_7598,N_7581);
or U8994 (N_8994,N_7945,N_7932);
xnor U8995 (N_8995,N_7954,N_7946);
nor U8996 (N_8996,N_7705,N_8330);
or U8997 (N_8997,N_7404,N_8379);
or U8998 (N_8998,N_7530,N_8353);
xor U8999 (N_8999,N_7627,N_7597);
nor U9000 (N_9000,N_7765,N_7221);
xor U9001 (N_9001,N_7446,N_7904);
nor U9002 (N_9002,N_7403,N_7957);
and U9003 (N_9003,N_7212,N_8256);
and U9004 (N_9004,N_8289,N_7943);
and U9005 (N_9005,N_7531,N_8094);
and U9006 (N_9006,N_8273,N_7554);
and U9007 (N_9007,N_7678,N_8123);
or U9008 (N_9008,N_7536,N_8326);
and U9009 (N_9009,N_8217,N_8095);
xor U9010 (N_9010,N_8336,N_8397);
or U9011 (N_9011,N_8371,N_7589);
nor U9012 (N_9012,N_7700,N_7872);
xnor U9013 (N_9013,N_7871,N_7645);
xnor U9014 (N_9014,N_7991,N_7930);
nor U9015 (N_9015,N_8242,N_7384);
nor U9016 (N_9016,N_8145,N_7450);
nor U9017 (N_9017,N_7298,N_8069);
or U9018 (N_9018,N_8031,N_7556);
nor U9019 (N_9019,N_7828,N_7526);
and U9020 (N_9020,N_7963,N_7245);
nor U9021 (N_9021,N_8356,N_7248);
nor U9022 (N_9022,N_7283,N_7215);
nor U9023 (N_9023,N_7807,N_7805);
xor U9024 (N_9024,N_8109,N_7672);
nand U9025 (N_9025,N_7511,N_7339);
nor U9026 (N_9026,N_7718,N_7342);
nor U9027 (N_9027,N_8196,N_7502);
nand U9028 (N_9028,N_8074,N_7698);
or U9029 (N_9029,N_8332,N_7832);
nor U9030 (N_9030,N_7340,N_7626);
or U9031 (N_9031,N_7568,N_7322);
nor U9032 (N_9032,N_7484,N_7376);
and U9033 (N_9033,N_8285,N_7886);
xnor U9034 (N_9034,N_7222,N_8220);
xor U9035 (N_9035,N_7371,N_7417);
or U9036 (N_9036,N_7646,N_7350);
nand U9037 (N_9037,N_7758,N_7726);
xor U9038 (N_9038,N_8049,N_7468);
nand U9039 (N_9039,N_7553,N_7694);
nor U9040 (N_9040,N_7417,N_8183);
and U9041 (N_9041,N_7354,N_7505);
or U9042 (N_9042,N_7602,N_8132);
and U9043 (N_9043,N_7594,N_7887);
or U9044 (N_9044,N_7393,N_8212);
nor U9045 (N_9045,N_7582,N_7934);
or U9046 (N_9046,N_7910,N_8326);
or U9047 (N_9047,N_8389,N_7441);
xnor U9048 (N_9048,N_8183,N_7614);
nor U9049 (N_9049,N_7574,N_7374);
or U9050 (N_9050,N_8284,N_8050);
and U9051 (N_9051,N_8175,N_8016);
nand U9052 (N_9052,N_7261,N_7822);
and U9053 (N_9053,N_7759,N_7689);
and U9054 (N_9054,N_7277,N_7994);
or U9055 (N_9055,N_7904,N_7756);
or U9056 (N_9056,N_7812,N_7546);
nor U9057 (N_9057,N_7631,N_7249);
nand U9058 (N_9058,N_7782,N_7978);
nand U9059 (N_9059,N_7610,N_8005);
nor U9060 (N_9060,N_7355,N_7477);
xnor U9061 (N_9061,N_8104,N_7738);
nand U9062 (N_9062,N_8390,N_7430);
xnor U9063 (N_9063,N_7285,N_7514);
or U9064 (N_9064,N_7627,N_8365);
nand U9065 (N_9065,N_7813,N_8071);
nor U9066 (N_9066,N_7981,N_7536);
nand U9067 (N_9067,N_8041,N_7549);
xor U9068 (N_9068,N_7351,N_7903);
nor U9069 (N_9069,N_8050,N_7277);
or U9070 (N_9070,N_7879,N_7990);
and U9071 (N_9071,N_8152,N_7898);
or U9072 (N_9072,N_7254,N_8038);
xor U9073 (N_9073,N_8187,N_7635);
or U9074 (N_9074,N_7338,N_7473);
and U9075 (N_9075,N_8195,N_7598);
and U9076 (N_9076,N_8100,N_7813);
or U9077 (N_9077,N_8149,N_7892);
or U9078 (N_9078,N_7245,N_7516);
xor U9079 (N_9079,N_7341,N_7889);
nand U9080 (N_9080,N_7935,N_8238);
and U9081 (N_9081,N_8202,N_8224);
xnor U9082 (N_9082,N_7477,N_7980);
nand U9083 (N_9083,N_7758,N_7850);
xnor U9084 (N_9084,N_8096,N_8246);
nor U9085 (N_9085,N_7378,N_7924);
and U9086 (N_9086,N_7357,N_7622);
nand U9087 (N_9087,N_7895,N_7981);
nand U9088 (N_9088,N_7424,N_8267);
nor U9089 (N_9089,N_8074,N_7820);
xnor U9090 (N_9090,N_7503,N_7288);
xnor U9091 (N_9091,N_7961,N_7883);
and U9092 (N_9092,N_7770,N_7951);
nand U9093 (N_9093,N_7980,N_7203);
nand U9094 (N_9094,N_8036,N_7532);
or U9095 (N_9095,N_7680,N_7407);
xnor U9096 (N_9096,N_8323,N_7451);
xnor U9097 (N_9097,N_7263,N_8340);
xnor U9098 (N_9098,N_8188,N_7257);
nor U9099 (N_9099,N_7984,N_7452);
nor U9100 (N_9100,N_7970,N_7742);
and U9101 (N_9101,N_7345,N_7503);
and U9102 (N_9102,N_7387,N_8233);
xnor U9103 (N_9103,N_8358,N_7798);
nand U9104 (N_9104,N_7408,N_7882);
nand U9105 (N_9105,N_7968,N_7391);
nand U9106 (N_9106,N_7773,N_8042);
xnor U9107 (N_9107,N_7776,N_8180);
and U9108 (N_9108,N_7430,N_7882);
nor U9109 (N_9109,N_7412,N_7738);
xnor U9110 (N_9110,N_7972,N_7598);
xnor U9111 (N_9111,N_7399,N_8195);
xor U9112 (N_9112,N_7596,N_7655);
xor U9113 (N_9113,N_8238,N_7325);
nor U9114 (N_9114,N_8333,N_8262);
xor U9115 (N_9115,N_7596,N_7809);
nor U9116 (N_9116,N_8173,N_8076);
nor U9117 (N_9117,N_8168,N_7971);
or U9118 (N_9118,N_8125,N_7291);
nor U9119 (N_9119,N_8237,N_7921);
and U9120 (N_9120,N_7734,N_8280);
or U9121 (N_9121,N_7250,N_7580);
or U9122 (N_9122,N_8284,N_7552);
nand U9123 (N_9123,N_7340,N_8206);
xnor U9124 (N_9124,N_7264,N_7532);
and U9125 (N_9125,N_8056,N_8337);
nor U9126 (N_9126,N_7563,N_7415);
nand U9127 (N_9127,N_8161,N_8329);
xor U9128 (N_9128,N_8267,N_8255);
nor U9129 (N_9129,N_7882,N_8111);
nand U9130 (N_9130,N_7808,N_7254);
and U9131 (N_9131,N_7677,N_7549);
xnor U9132 (N_9132,N_8080,N_7835);
and U9133 (N_9133,N_7698,N_7716);
xor U9134 (N_9134,N_7913,N_7540);
nor U9135 (N_9135,N_8130,N_7493);
nand U9136 (N_9136,N_7876,N_8223);
xor U9137 (N_9137,N_7752,N_7739);
nor U9138 (N_9138,N_7805,N_7862);
nor U9139 (N_9139,N_7865,N_7438);
xnor U9140 (N_9140,N_7955,N_7552);
or U9141 (N_9141,N_8114,N_8270);
or U9142 (N_9142,N_7244,N_8218);
nand U9143 (N_9143,N_7899,N_7837);
xnor U9144 (N_9144,N_7257,N_7261);
nor U9145 (N_9145,N_7613,N_7316);
nor U9146 (N_9146,N_7489,N_8335);
nand U9147 (N_9147,N_8393,N_8311);
or U9148 (N_9148,N_7853,N_8166);
nand U9149 (N_9149,N_7422,N_8319);
nand U9150 (N_9150,N_7787,N_7257);
and U9151 (N_9151,N_7490,N_8311);
or U9152 (N_9152,N_8032,N_7740);
xor U9153 (N_9153,N_7406,N_8292);
and U9154 (N_9154,N_8347,N_7803);
and U9155 (N_9155,N_7986,N_7941);
and U9156 (N_9156,N_7243,N_7683);
nor U9157 (N_9157,N_8389,N_7770);
nand U9158 (N_9158,N_7589,N_8119);
nor U9159 (N_9159,N_7266,N_7781);
nor U9160 (N_9160,N_7871,N_7430);
xnor U9161 (N_9161,N_7570,N_8083);
and U9162 (N_9162,N_7805,N_7338);
nand U9163 (N_9163,N_7546,N_7831);
nand U9164 (N_9164,N_7873,N_8205);
nand U9165 (N_9165,N_7479,N_7381);
and U9166 (N_9166,N_7782,N_8344);
nand U9167 (N_9167,N_7945,N_7215);
nand U9168 (N_9168,N_7860,N_7687);
and U9169 (N_9169,N_8149,N_7248);
nand U9170 (N_9170,N_7948,N_8333);
nand U9171 (N_9171,N_8273,N_7231);
and U9172 (N_9172,N_7737,N_8066);
nand U9173 (N_9173,N_7543,N_7415);
nand U9174 (N_9174,N_8051,N_8246);
nand U9175 (N_9175,N_8335,N_7277);
and U9176 (N_9176,N_7282,N_7278);
nand U9177 (N_9177,N_7934,N_7835);
and U9178 (N_9178,N_7482,N_7801);
xor U9179 (N_9179,N_8320,N_7212);
and U9180 (N_9180,N_8250,N_7588);
nand U9181 (N_9181,N_7564,N_7834);
and U9182 (N_9182,N_8384,N_7592);
or U9183 (N_9183,N_8165,N_7803);
and U9184 (N_9184,N_7571,N_7792);
and U9185 (N_9185,N_8128,N_8142);
xor U9186 (N_9186,N_7792,N_7737);
xnor U9187 (N_9187,N_7522,N_8369);
or U9188 (N_9188,N_7317,N_7454);
or U9189 (N_9189,N_7342,N_7411);
or U9190 (N_9190,N_7871,N_7789);
or U9191 (N_9191,N_7416,N_8234);
xnor U9192 (N_9192,N_7978,N_7766);
and U9193 (N_9193,N_8290,N_7788);
nor U9194 (N_9194,N_7459,N_8210);
nand U9195 (N_9195,N_7612,N_7445);
xnor U9196 (N_9196,N_8245,N_8100);
nand U9197 (N_9197,N_8240,N_7352);
nand U9198 (N_9198,N_8214,N_8217);
xnor U9199 (N_9199,N_7518,N_7302);
or U9200 (N_9200,N_8397,N_7687);
or U9201 (N_9201,N_7339,N_7285);
nand U9202 (N_9202,N_7204,N_7767);
and U9203 (N_9203,N_7224,N_7393);
or U9204 (N_9204,N_8244,N_7933);
and U9205 (N_9205,N_7516,N_7263);
nand U9206 (N_9206,N_7759,N_7412);
and U9207 (N_9207,N_7962,N_7548);
and U9208 (N_9208,N_7498,N_7634);
nor U9209 (N_9209,N_7759,N_8072);
nor U9210 (N_9210,N_7596,N_8067);
nor U9211 (N_9211,N_7932,N_7767);
nor U9212 (N_9212,N_7856,N_8076);
and U9213 (N_9213,N_7637,N_7295);
and U9214 (N_9214,N_7334,N_7820);
and U9215 (N_9215,N_7612,N_7640);
or U9216 (N_9216,N_7250,N_8050);
and U9217 (N_9217,N_8101,N_8014);
xnor U9218 (N_9218,N_7672,N_8130);
nor U9219 (N_9219,N_8282,N_7544);
nor U9220 (N_9220,N_8012,N_8368);
and U9221 (N_9221,N_7371,N_7272);
and U9222 (N_9222,N_7853,N_7786);
xor U9223 (N_9223,N_8116,N_8112);
nor U9224 (N_9224,N_7875,N_7441);
nand U9225 (N_9225,N_7536,N_8199);
or U9226 (N_9226,N_8259,N_7866);
and U9227 (N_9227,N_8051,N_7240);
xnor U9228 (N_9228,N_7759,N_7332);
nand U9229 (N_9229,N_8385,N_7258);
and U9230 (N_9230,N_7975,N_7519);
nand U9231 (N_9231,N_7357,N_7566);
nand U9232 (N_9232,N_7336,N_8147);
nor U9233 (N_9233,N_7996,N_7556);
and U9234 (N_9234,N_8239,N_8030);
and U9235 (N_9235,N_8228,N_7283);
xnor U9236 (N_9236,N_7657,N_8179);
nor U9237 (N_9237,N_7991,N_7679);
nor U9238 (N_9238,N_7673,N_8124);
or U9239 (N_9239,N_7973,N_8114);
nand U9240 (N_9240,N_7916,N_7809);
or U9241 (N_9241,N_8270,N_7573);
and U9242 (N_9242,N_8142,N_7223);
xor U9243 (N_9243,N_7731,N_7774);
xnor U9244 (N_9244,N_7416,N_7874);
xor U9245 (N_9245,N_8200,N_7641);
nor U9246 (N_9246,N_7659,N_7884);
nor U9247 (N_9247,N_8354,N_7801);
nor U9248 (N_9248,N_7240,N_7672);
or U9249 (N_9249,N_7915,N_8256);
xnor U9250 (N_9250,N_7653,N_8209);
nor U9251 (N_9251,N_7805,N_8225);
nor U9252 (N_9252,N_7507,N_7613);
and U9253 (N_9253,N_7979,N_7776);
xnor U9254 (N_9254,N_7395,N_7569);
xnor U9255 (N_9255,N_7991,N_7758);
and U9256 (N_9256,N_8198,N_8154);
or U9257 (N_9257,N_8166,N_7632);
nor U9258 (N_9258,N_7331,N_7903);
xnor U9259 (N_9259,N_7867,N_7973);
or U9260 (N_9260,N_7307,N_7543);
and U9261 (N_9261,N_7849,N_8273);
and U9262 (N_9262,N_7627,N_7725);
or U9263 (N_9263,N_7520,N_8038);
nand U9264 (N_9264,N_7590,N_7945);
or U9265 (N_9265,N_7220,N_7589);
nor U9266 (N_9266,N_7485,N_8144);
and U9267 (N_9267,N_8247,N_7264);
or U9268 (N_9268,N_7478,N_7947);
or U9269 (N_9269,N_8062,N_8280);
nand U9270 (N_9270,N_7233,N_7333);
nand U9271 (N_9271,N_8192,N_8124);
nand U9272 (N_9272,N_7575,N_8204);
and U9273 (N_9273,N_8150,N_7959);
nand U9274 (N_9274,N_7657,N_7761);
nor U9275 (N_9275,N_7465,N_7727);
and U9276 (N_9276,N_8363,N_7907);
nand U9277 (N_9277,N_7617,N_7449);
nor U9278 (N_9278,N_7273,N_7900);
or U9279 (N_9279,N_7640,N_8381);
xor U9280 (N_9280,N_8337,N_7665);
nor U9281 (N_9281,N_7365,N_8149);
or U9282 (N_9282,N_7475,N_7830);
nor U9283 (N_9283,N_7358,N_7590);
xnor U9284 (N_9284,N_8239,N_7297);
nor U9285 (N_9285,N_8188,N_7280);
and U9286 (N_9286,N_8261,N_8253);
and U9287 (N_9287,N_7695,N_7443);
and U9288 (N_9288,N_7849,N_8393);
and U9289 (N_9289,N_7743,N_7965);
and U9290 (N_9290,N_7408,N_8337);
and U9291 (N_9291,N_7717,N_7315);
xnor U9292 (N_9292,N_7262,N_8056);
nor U9293 (N_9293,N_7895,N_8276);
or U9294 (N_9294,N_8112,N_7576);
nand U9295 (N_9295,N_7777,N_8012);
and U9296 (N_9296,N_7340,N_8053);
nand U9297 (N_9297,N_7514,N_7200);
xor U9298 (N_9298,N_7534,N_8387);
or U9299 (N_9299,N_7470,N_8237);
xnor U9300 (N_9300,N_7300,N_7343);
nor U9301 (N_9301,N_7585,N_8332);
xor U9302 (N_9302,N_8214,N_7832);
xor U9303 (N_9303,N_7524,N_7631);
xor U9304 (N_9304,N_7907,N_8231);
nand U9305 (N_9305,N_7387,N_7247);
or U9306 (N_9306,N_7278,N_7747);
nand U9307 (N_9307,N_7304,N_8009);
and U9308 (N_9308,N_8344,N_7656);
nor U9309 (N_9309,N_8335,N_7968);
xnor U9310 (N_9310,N_8187,N_7781);
or U9311 (N_9311,N_7648,N_8017);
nand U9312 (N_9312,N_7378,N_7645);
or U9313 (N_9313,N_7651,N_7740);
or U9314 (N_9314,N_7285,N_7933);
nor U9315 (N_9315,N_7712,N_7571);
nand U9316 (N_9316,N_7453,N_7791);
nand U9317 (N_9317,N_7954,N_7268);
or U9318 (N_9318,N_7324,N_7679);
nor U9319 (N_9319,N_8297,N_7648);
nor U9320 (N_9320,N_8321,N_7698);
or U9321 (N_9321,N_7717,N_7735);
nand U9322 (N_9322,N_8289,N_8097);
xnor U9323 (N_9323,N_7750,N_8221);
and U9324 (N_9324,N_7953,N_8059);
and U9325 (N_9325,N_7532,N_7629);
or U9326 (N_9326,N_7802,N_8076);
or U9327 (N_9327,N_7252,N_8384);
nand U9328 (N_9328,N_7899,N_8177);
nand U9329 (N_9329,N_8163,N_7538);
nand U9330 (N_9330,N_7334,N_7778);
nand U9331 (N_9331,N_8332,N_7631);
xor U9332 (N_9332,N_8321,N_7590);
or U9333 (N_9333,N_7215,N_7691);
nand U9334 (N_9334,N_7294,N_7534);
nand U9335 (N_9335,N_7911,N_7892);
and U9336 (N_9336,N_8368,N_8105);
nand U9337 (N_9337,N_7370,N_7287);
nor U9338 (N_9338,N_7280,N_7802);
nand U9339 (N_9339,N_8149,N_7326);
xnor U9340 (N_9340,N_7799,N_7870);
and U9341 (N_9341,N_7413,N_8242);
nor U9342 (N_9342,N_7973,N_7327);
or U9343 (N_9343,N_8078,N_8382);
xnor U9344 (N_9344,N_8237,N_7736);
or U9345 (N_9345,N_7656,N_7803);
nor U9346 (N_9346,N_8031,N_7673);
and U9347 (N_9347,N_7816,N_8111);
or U9348 (N_9348,N_7453,N_8046);
nor U9349 (N_9349,N_7226,N_7934);
or U9350 (N_9350,N_7849,N_8378);
and U9351 (N_9351,N_8294,N_8272);
nand U9352 (N_9352,N_8046,N_8108);
nor U9353 (N_9353,N_7275,N_7522);
nand U9354 (N_9354,N_8186,N_7627);
or U9355 (N_9355,N_7853,N_7674);
nor U9356 (N_9356,N_7906,N_7765);
nor U9357 (N_9357,N_7952,N_7319);
xor U9358 (N_9358,N_7227,N_7292);
xnor U9359 (N_9359,N_7868,N_8016);
xor U9360 (N_9360,N_8284,N_8061);
nor U9361 (N_9361,N_8170,N_7741);
and U9362 (N_9362,N_7320,N_7790);
or U9363 (N_9363,N_7728,N_7983);
nor U9364 (N_9364,N_8066,N_7378);
nand U9365 (N_9365,N_7612,N_7636);
nor U9366 (N_9366,N_7731,N_8013);
xor U9367 (N_9367,N_7285,N_8272);
nor U9368 (N_9368,N_7834,N_7635);
nand U9369 (N_9369,N_8013,N_7889);
xor U9370 (N_9370,N_7281,N_8243);
nand U9371 (N_9371,N_7998,N_7934);
nor U9372 (N_9372,N_7889,N_8158);
or U9373 (N_9373,N_7423,N_7997);
nor U9374 (N_9374,N_7967,N_8085);
and U9375 (N_9375,N_7994,N_7542);
or U9376 (N_9376,N_7387,N_7360);
or U9377 (N_9377,N_7916,N_7552);
xor U9378 (N_9378,N_8399,N_7457);
and U9379 (N_9379,N_8321,N_7675);
xnor U9380 (N_9380,N_7238,N_7252);
and U9381 (N_9381,N_7859,N_7552);
nand U9382 (N_9382,N_7317,N_8189);
or U9383 (N_9383,N_7398,N_7243);
nor U9384 (N_9384,N_8023,N_8025);
xnor U9385 (N_9385,N_7566,N_8068);
nor U9386 (N_9386,N_7544,N_7445);
and U9387 (N_9387,N_7262,N_7550);
or U9388 (N_9388,N_7224,N_7381);
and U9389 (N_9389,N_8137,N_8195);
xor U9390 (N_9390,N_8239,N_7572);
nand U9391 (N_9391,N_7544,N_7403);
nand U9392 (N_9392,N_7905,N_7740);
nand U9393 (N_9393,N_8162,N_7386);
xor U9394 (N_9394,N_8069,N_8248);
nand U9395 (N_9395,N_7999,N_7944);
or U9396 (N_9396,N_7804,N_7893);
nand U9397 (N_9397,N_8337,N_8076);
xnor U9398 (N_9398,N_8248,N_8240);
or U9399 (N_9399,N_8310,N_7542);
and U9400 (N_9400,N_7590,N_7614);
or U9401 (N_9401,N_7804,N_7699);
xnor U9402 (N_9402,N_7932,N_7578);
xnor U9403 (N_9403,N_7789,N_7860);
and U9404 (N_9404,N_8329,N_7222);
nand U9405 (N_9405,N_7810,N_7623);
and U9406 (N_9406,N_8349,N_7491);
or U9407 (N_9407,N_7421,N_8177);
and U9408 (N_9408,N_8161,N_7653);
xnor U9409 (N_9409,N_7641,N_7882);
xor U9410 (N_9410,N_8341,N_7710);
and U9411 (N_9411,N_8132,N_7747);
and U9412 (N_9412,N_8076,N_7615);
xor U9413 (N_9413,N_8088,N_8148);
or U9414 (N_9414,N_8139,N_8133);
nor U9415 (N_9415,N_7412,N_8104);
nand U9416 (N_9416,N_7821,N_7747);
and U9417 (N_9417,N_7897,N_7285);
and U9418 (N_9418,N_7327,N_7701);
nand U9419 (N_9419,N_7906,N_7937);
xnor U9420 (N_9420,N_7562,N_8017);
or U9421 (N_9421,N_8032,N_8104);
nor U9422 (N_9422,N_8248,N_8196);
xnor U9423 (N_9423,N_8219,N_7680);
nor U9424 (N_9424,N_8234,N_7290);
nor U9425 (N_9425,N_8243,N_8112);
or U9426 (N_9426,N_7469,N_8067);
and U9427 (N_9427,N_7838,N_8061);
or U9428 (N_9428,N_8240,N_7318);
nand U9429 (N_9429,N_7519,N_8129);
or U9430 (N_9430,N_7735,N_7659);
xor U9431 (N_9431,N_7374,N_8171);
or U9432 (N_9432,N_7627,N_8125);
nor U9433 (N_9433,N_7937,N_7688);
nand U9434 (N_9434,N_8392,N_7480);
or U9435 (N_9435,N_7280,N_7458);
nand U9436 (N_9436,N_8218,N_8391);
or U9437 (N_9437,N_8087,N_7393);
and U9438 (N_9438,N_8034,N_8339);
nand U9439 (N_9439,N_7313,N_7723);
or U9440 (N_9440,N_8334,N_7504);
nor U9441 (N_9441,N_7953,N_7475);
or U9442 (N_9442,N_8336,N_7615);
or U9443 (N_9443,N_7597,N_7874);
xnor U9444 (N_9444,N_7202,N_8051);
nor U9445 (N_9445,N_7531,N_7575);
nand U9446 (N_9446,N_8062,N_7763);
or U9447 (N_9447,N_7300,N_7327);
and U9448 (N_9448,N_7583,N_8360);
nand U9449 (N_9449,N_7588,N_7353);
nand U9450 (N_9450,N_7841,N_8375);
or U9451 (N_9451,N_8365,N_7521);
or U9452 (N_9452,N_8194,N_7977);
xor U9453 (N_9453,N_7671,N_7393);
xor U9454 (N_9454,N_8209,N_7647);
nand U9455 (N_9455,N_7500,N_7993);
xnor U9456 (N_9456,N_8340,N_7995);
or U9457 (N_9457,N_7966,N_7659);
xnor U9458 (N_9458,N_7377,N_8356);
xor U9459 (N_9459,N_7653,N_7445);
or U9460 (N_9460,N_7541,N_7695);
xnor U9461 (N_9461,N_7550,N_8194);
nand U9462 (N_9462,N_8229,N_7435);
and U9463 (N_9463,N_7308,N_7494);
nand U9464 (N_9464,N_8328,N_8103);
nand U9465 (N_9465,N_7637,N_7898);
nand U9466 (N_9466,N_8149,N_7758);
xnor U9467 (N_9467,N_8062,N_7516);
nor U9468 (N_9468,N_7316,N_7224);
and U9469 (N_9469,N_7366,N_7821);
xor U9470 (N_9470,N_7230,N_8195);
and U9471 (N_9471,N_8240,N_8165);
xnor U9472 (N_9472,N_8233,N_8259);
nor U9473 (N_9473,N_7414,N_7694);
nand U9474 (N_9474,N_7844,N_7228);
xor U9475 (N_9475,N_7411,N_7693);
xor U9476 (N_9476,N_8356,N_7563);
nor U9477 (N_9477,N_7827,N_7469);
and U9478 (N_9478,N_7528,N_8125);
xor U9479 (N_9479,N_8099,N_7935);
nor U9480 (N_9480,N_7299,N_8229);
and U9481 (N_9481,N_7890,N_7422);
nor U9482 (N_9482,N_8291,N_8391);
nand U9483 (N_9483,N_8139,N_8296);
and U9484 (N_9484,N_7378,N_8315);
xor U9485 (N_9485,N_8309,N_7978);
xnor U9486 (N_9486,N_7946,N_7895);
or U9487 (N_9487,N_7500,N_8085);
and U9488 (N_9488,N_7308,N_7746);
nand U9489 (N_9489,N_7956,N_7782);
nor U9490 (N_9490,N_7328,N_8271);
nand U9491 (N_9491,N_8036,N_8299);
nor U9492 (N_9492,N_7254,N_7417);
or U9493 (N_9493,N_7852,N_7482);
nand U9494 (N_9494,N_7692,N_7929);
nand U9495 (N_9495,N_8170,N_8177);
and U9496 (N_9496,N_7747,N_7459);
and U9497 (N_9497,N_7608,N_7850);
or U9498 (N_9498,N_7771,N_7588);
xor U9499 (N_9499,N_8239,N_7526);
or U9500 (N_9500,N_7357,N_7409);
nor U9501 (N_9501,N_7729,N_7864);
nor U9502 (N_9502,N_7679,N_7247);
nor U9503 (N_9503,N_7582,N_7345);
nand U9504 (N_9504,N_8237,N_8303);
xnor U9505 (N_9505,N_7712,N_7500);
or U9506 (N_9506,N_7700,N_7835);
and U9507 (N_9507,N_8175,N_7568);
or U9508 (N_9508,N_7682,N_8116);
nor U9509 (N_9509,N_8196,N_8256);
and U9510 (N_9510,N_7368,N_7593);
nand U9511 (N_9511,N_8349,N_7837);
or U9512 (N_9512,N_8184,N_7377);
and U9513 (N_9513,N_7966,N_7677);
and U9514 (N_9514,N_7201,N_7406);
or U9515 (N_9515,N_7944,N_7792);
or U9516 (N_9516,N_8345,N_8368);
and U9517 (N_9517,N_8118,N_7661);
nor U9518 (N_9518,N_7295,N_7766);
nand U9519 (N_9519,N_7951,N_7855);
or U9520 (N_9520,N_8239,N_7622);
xor U9521 (N_9521,N_8223,N_7717);
xor U9522 (N_9522,N_7771,N_7259);
or U9523 (N_9523,N_7327,N_8353);
nand U9524 (N_9524,N_8116,N_8249);
and U9525 (N_9525,N_7529,N_7915);
and U9526 (N_9526,N_7630,N_7213);
or U9527 (N_9527,N_8055,N_7421);
or U9528 (N_9528,N_8106,N_7223);
or U9529 (N_9529,N_7902,N_8399);
nand U9530 (N_9530,N_7802,N_7405);
nor U9531 (N_9531,N_7884,N_8121);
nand U9532 (N_9532,N_7299,N_7698);
nor U9533 (N_9533,N_7909,N_7228);
nor U9534 (N_9534,N_7226,N_8023);
nand U9535 (N_9535,N_7286,N_8320);
nand U9536 (N_9536,N_7655,N_7282);
nor U9537 (N_9537,N_7393,N_7455);
and U9538 (N_9538,N_7363,N_8067);
nor U9539 (N_9539,N_7439,N_8028);
and U9540 (N_9540,N_7737,N_7469);
nand U9541 (N_9541,N_7266,N_7369);
nor U9542 (N_9542,N_8393,N_7385);
and U9543 (N_9543,N_8031,N_7409);
xnor U9544 (N_9544,N_8005,N_8084);
nand U9545 (N_9545,N_7386,N_8071);
xnor U9546 (N_9546,N_8045,N_7660);
or U9547 (N_9547,N_7615,N_7993);
xnor U9548 (N_9548,N_8117,N_8052);
nor U9549 (N_9549,N_7422,N_7572);
nor U9550 (N_9550,N_7433,N_8051);
xor U9551 (N_9551,N_7377,N_7749);
nand U9552 (N_9552,N_8134,N_7475);
xnor U9553 (N_9553,N_8354,N_7680);
xor U9554 (N_9554,N_7382,N_8193);
nand U9555 (N_9555,N_7820,N_7233);
nand U9556 (N_9556,N_7827,N_8215);
or U9557 (N_9557,N_7369,N_8326);
xor U9558 (N_9558,N_7721,N_7233);
or U9559 (N_9559,N_7298,N_7601);
and U9560 (N_9560,N_8023,N_8195);
nor U9561 (N_9561,N_8343,N_7896);
or U9562 (N_9562,N_8178,N_7335);
nor U9563 (N_9563,N_7322,N_7495);
and U9564 (N_9564,N_8055,N_7393);
nand U9565 (N_9565,N_8154,N_8101);
and U9566 (N_9566,N_7242,N_7359);
nor U9567 (N_9567,N_7380,N_8127);
nor U9568 (N_9568,N_7752,N_8331);
nor U9569 (N_9569,N_8048,N_7651);
nor U9570 (N_9570,N_8207,N_7363);
nand U9571 (N_9571,N_7717,N_7513);
nand U9572 (N_9572,N_7950,N_8176);
nor U9573 (N_9573,N_7716,N_7829);
nand U9574 (N_9574,N_7264,N_8091);
nor U9575 (N_9575,N_7568,N_7536);
nor U9576 (N_9576,N_7552,N_7434);
nor U9577 (N_9577,N_8178,N_8103);
or U9578 (N_9578,N_7642,N_7725);
or U9579 (N_9579,N_8203,N_7221);
or U9580 (N_9580,N_7319,N_7971);
and U9581 (N_9581,N_7688,N_7521);
or U9582 (N_9582,N_8205,N_7896);
and U9583 (N_9583,N_7422,N_7394);
and U9584 (N_9584,N_7327,N_7204);
xnor U9585 (N_9585,N_7341,N_7340);
and U9586 (N_9586,N_7722,N_7551);
xnor U9587 (N_9587,N_8022,N_7956);
nand U9588 (N_9588,N_7955,N_7827);
or U9589 (N_9589,N_7515,N_7375);
nor U9590 (N_9590,N_8332,N_7532);
or U9591 (N_9591,N_7739,N_7722);
and U9592 (N_9592,N_7209,N_7409);
nor U9593 (N_9593,N_7433,N_7467);
or U9594 (N_9594,N_7405,N_7464);
nand U9595 (N_9595,N_7967,N_8273);
nand U9596 (N_9596,N_7406,N_8238);
or U9597 (N_9597,N_7402,N_7771);
xor U9598 (N_9598,N_7563,N_7327);
nand U9599 (N_9599,N_7269,N_7958);
xnor U9600 (N_9600,N_9197,N_9238);
nand U9601 (N_9601,N_9571,N_8901);
nand U9602 (N_9602,N_9275,N_9558);
and U9603 (N_9603,N_9024,N_8858);
nor U9604 (N_9604,N_8913,N_9041);
xnor U9605 (N_9605,N_8446,N_8874);
or U9606 (N_9606,N_9505,N_8632);
or U9607 (N_9607,N_8753,N_9004);
nand U9608 (N_9608,N_9577,N_8806);
nor U9609 (N_9609,N_9599,N_8769);
nor U9610 (N_9610,N_8415,N_9475);
nand U9611 (N_9611,N_9279,N_9454);
or U9612 (N_9612,N_9455,N_9163);
or U9613 (N_9613,N_8786,N_8688);
nor U9614 (N_9614,N_8687,N_8977);
xnor U9615 (N_9615,N_8684,N_9368);
nor U9616 (N_9616,N_9225,N_9261);
xor U9617 (N_9617,N_8610,N_9093);
or U9618 (N_9618,N_8867,N_9022);
or U9619 (N_9619,N_9509,N_8422);
and U9620 (N_9620,N_8706,N_8521);
and U9621 (N_9621,N_8408,N_8464);
and U9622 (N_9622,N_9292,N_8844);
or U9623 (N_9623,N_9109,N_8971);
and U9624 (N_9624,N_8961,N_9299);
nor U9625 (N_9625,N_8908,N_9144);
nor U9626 (N_9626,N_9335,N_9307);
or U9627 (N_9627,N_8525,N_9003);
xor U9628 (N_9628,N_9158,N_9512);
and U9629 (N_9629,N_9028,N_9593);
and U9630 (N_9630,N_8540,N_9546);
xor U9631 (N_9631,N_9116,N_9328);
nand U9632 (N_9632,N_9588,N_8893);
xnor U9633 (N_9633,N_8991,N_8578);
nor U9634 (N_9634,N_9502,N_8660);
nand U9635 (N_9635,N_8418,N_8878);
nor U9636 (N_9636,N_9528,N_8556);
nor U9637 (N_9637,N_8990,N_8775);
and U9638 (N_9638,N_9564,N_8881);
nand U9639 (N_9639,N_9085,N_8470);
and U9640 (N_9640,N_8850,N_8467);
xor U9641 (N_9641,N_8742,N_8537);
nor U9642 (N_9642,N_9229,N_9337);
or U9643 (N_9643,N_9316,N_8546);
or U9644 (N_9644,N_9412,N_9443);
nor U9645 (N_9645,N_8827,N_8960);
xnor U9646 (N_9646,N_9057,N_8992);
or U9647 (N_9647,N_9138,N_8608);
nor U9648 (N_9648,N_8488,N_8612);
or U9649 (N_9649,N_8561,N_9190);
or U9650 (N_9650,N_9483,N_9370);
and U9651 (N_9651,N_8939,N_8439);
nand U9652 (N_9652,N_8438,N_8749);
and U9653 (N_9653,N_9461,N_9516);
or U9654 (N_9654,N_9389,N_8657);
or U9655 (N_9655,N_8427,N_9569);
or U9656 (N_9656,N_8790,N_9269);
nand U9657 (N_9657,N_9213,N_8855);
and U9658 (N_9658,N_8633,N_9311);
nor U9659 (N_9659,N_9557,N_9131);
nor U9660 (N_9660,N_9205,N_9452);
and U9661 (N_9661,N_9011,N_8491);
xnor U9662 (N_9662,N_8982,N_8699);
or U9663 (N_9663,N_8412,N_8626);
or U9664 (N_9664,N_9545,N_9122);
nand U9665 (N_9665,N_9034,N_9556);
nand U9666 (N_9666,N_8936,N_9295);
xor U9667 (N_9667,N_8804,N_8948);
and U9668 (N_9668,N_8704,N_9203);
or U9669 (N_9669,N_8429,N_8555);
or U9670 (N_9670,N_8435,N_9302);
or U9671 (N_9671,N_9117,N_9110);
xor U9672 (N_9672,N_9182,N_9582);
or U9673 (N_9673,N_9542,N_8744);
and U9674 (N_9674,N_8778,N_8698);
or U9675 (N_9675,N_9460,N_8882);
and U9676 (N_9676,N_8647,N_8656);
and U9677 (N_9677,N_8835,N_9031);
xor U9678 (N_9678,N_8443,N_9027);
nor U9679 (N_9679,N_8695,N_8501);
nor U9680 (N_9680,N_8801,N_8539);
nor U9681 (N_9681,N_8950,N_9112);
or U9682 (N_9682,N_8883,N_9107);
or U9683 (N_9683,N_8962,N_8493);
or U9684 (N_9684,N_8425,N_8642);
nand U9685 (N_9685,N_8641,N_8606);
or U9686 (N_9686,N_9422,N_9060);
and U9687 (N_9687,N_9409,N_9527);
and U9688 (N_9688,N_9391,N_9322);
nand U9689 (N_9689,N_9142,N_9192);
and U9690 (N_9690,N_9375,N_9305);
xnor U9691 (N_9691,N_9589,N_9490);
nor U9692 (N_9692,N_9084,N_9145);
or U9693 (N_9693,N_8870,N_9477);
and U9694 (N_9694,N_8964,N_8536);
nor U9695 (N_9695,N_9345,N_9222);
nor U9696 (N_9696,N_9567,N_9478);
xnor U9697 (N_9697,N_9369,N_8617);
and U9698 (N_9698,N_9541,N_9399);
and U9699 (N_9699,N_9088,N_8869);
xnor U9700 (N_9700,N_8965,N_9223);
nand U9701 (N_9701,N_9153,N_8789);
nor U9702 (N_9702,N_9232,N_9230);
xnor U9703 (N_9703,N_9036,N_9427);
nor U9704 (N_9704,N_8995,N_9099);
nand U9705 (N_9705,N_8889,N_8559);
xnor U9706 (N_9706,N_9137,N_9277);
xor U9707 (N_9707,N_8853,N_8413);
and U9708 (N_9708,N_9414,N_9150);
or U9709 (N_9709,N_9543,N_8837);
nand U9710 (N_9710,N_9095,N_9470);
nand U9711 (N_9711,N_8922,N_9172);
nor U9712 (N_9712,N_8979,N_9576);
and U9713 (N_9713,N_8598,N_9198);
and U9714 (N_9714,N_9151,N_9220);
or U9715 (N_9715,N_9450,N_9518);
and U9716 (N_9716,N_9039,N_8891);
nand U9717 (N_9717,N_9333,N_9342);
or U9718 (N_9718,N_9212,N_9407);
xnor U9719 (N_9719,N_8524,N_9380);
nand U9720 (N_9720,N_9260,N_9425);
xor U9721 (N_9721,N_8416,N_9390);
xor U9722 (N_9722,N_9421,N_9585);
or U9723 (N_9723,N_9550,N_8862);
nor U9724 (N_9724,N_9224,N_8511);
nand U9725 (N_9725,N_8678,N_9308);
nor U9726 (N_9726,N_8831,N_8860);
nand U9727 (N_9727,N_8787,N_9489);
nor U9728 (N_9728,N_8940,N_9132);
and U9729 (N_9729,N_9064,N_8822);
or U9730 (N_9730,N_9276,N_9206);
and U9731 (N_9731,N_8692,N_8655);
or U9732 (N_9732,N_9395,N_9570);
or U9733 (N_9733,N_8444,N_8918);
nand U9734 (N_9734,N_9533,N_8662);
xnor U9735 (N_9735,N_9456,N_9320);
nand U9736 (N_9736,N_8782,N_9274);
and U9737 (N_9737,N_8934,N_9030);
and U9738 (N_9738,N_8711,N_8465);
and U9739 (N_9739,N_9310,N_9167);
nor U9740 (N_9740,N_8760,N_8989);
nand U9741 (N_9741,N_9418,N_9429);
or U9742 (N_9742,N_9524,N_9382);
and U9743 (N_9743,N_9139,N_8586);
nand U9744 (N_9744,N_8988,N_8800);
nand U9745 (N_9745,N_9549,N_9365);
nand U9746 (N_9746,N_8739,N_9514);
nor U9747 (N_9747,N_9068,N_9289);
or U9748 (N_9748,N_9248,N_8798);
or U9749 (N_9749,N_9372,N_9411);
or U9750 (N_9750,N_9048,N_9510);
and U9751 (N_9751,N_9339,N_8797);
nand U9752 (N_9752,N_8892,N_8522);
or U9753 (N_9753,N_9234,N_9101);
nand U9754 (N_9754,N_9530,N_9468);
and U9755 (N_9755,N_9330,N_9325);
and U9756 (N_9756,N_9464,N_8620);
nand U9757 (N_9757,N_8880,N_8592);
nand U9758 (N_9758,N_9251,N_8474);
nor U9759 (N_9759,N_9501,N_9447);
and U9760 (N_9760,N_9202,N_8597);
nor U9761 (N_9761,N_9007,N_8628);
xnor U9762 (N_9762,N_8589,N_9294);
nor U9763 (N_9763,N_9207,N_8843);
xor U9764 (N_9764,N_9059,N_9191);
and U9765 (N_9765,N_8799,N_8667);
nand U9766 (N_9766,N_9226,N_8693);
and U9767 (N_9767,N_9584,N_9002);
xor U9768 (N_9768,N_8538,N_9026);
nand U9769 (N_9769,N_9023,N_9423);
nor U9770 (N_9770,N_9033,N_9194);
and U9771 (N_9771,N_9351,N_9332);
nor U9772 (N_9772,N_8861,N_9381);
nand U9773 (N_9773,N_9241,N_8879);
nand U9774 (N_9774,N_9119,N_9526);
nor U9775 (N_9775,N_8468,N_9492);
nand U9776 (N_9776,N_9596,N_8857);
xnor U9777 (N_9777,N_9383,N_8809);
nand U9778 (N_9778,N_9480,N_8567);
and U9779 (N_9779,N_9597,N_8496);
or U9780 (N_9780,N_9309,N_9331);
xor U9781 (N_9781,N_8920,N_8820);
nand U9782 (N_9782,N_9396,N_9096);
and U9783 (N_9783,N_9338,N_8544);
and U9784 (N_9784,N_9349,N_9431);
or U9785 (N_9785,N_9487,N_9108);
xnor U9786 (N_9786,N_8752,N_8925);
or U9787 (N_9787,N_9075,N_9211);
xor U9788 (N_9788,N_9240,N_8735);
nand U9789 (N_9789,N_9352,N_9079);
xnor U9790 (N_9790,N_9195,N_8941);
and U9791 (N_9791,N_8651,N_9056);
xor U9792 (N_9792,N_9547,N_8436);
or U9793 (N_9793,N_8504,N_8566);
and U9794 (N_9794,N_8954,N_9231);
or U9795 (N_9795,N_8421,N_8840);
nor U9796 (N_9796,N_8519,N_8645);
nor U9797 (N_9797,N_9405,N_8803);
nand U9798 (N_9798,N_9436,N_8508);
or U9799 (N_9799,N_8485,N_9453);
and U9800 (N_9800,N_9484,N_8814);
nor U9801 (N_9801,N_8963,N_9280);
nand U9802 (N_9802,N_8685,N_8723);
nor U9803 (N_9803,N_9018,N_8607);
and U9804 (N_9804,N_8914,N_8587);
xor U9805 (N_9805,N_8463,N_8825);
nor U9806 (N_9806,N_9287,N_8477);
nor U9807 (N_9807,N_9265,N_9449);
nand U9808 (N_9808,N_9035,N_9268);
xnor U9809 (N_9809,N_8709,N_8957);
nor U9810 (N_9810,N_8535,N_8781);
xnor U9811 (N_9811,N_8864,N_9221);
xnor U9812 (N_9812,N_8875,N_9176);
nand U9813 (N_9813,N_9156,N_9152);
nand U9814 (N_9814,N_8935,N_9540);
or U9815 (N_9815,N_9482,N_8531);
or U9816 (N_9816,N_8621,N_9020);
or U9817 (N_9817,N_8527,N_8661);
and U9818 (N_9818,N_9008,N_9091);
nor U9819 (N_9819,N_9233,N_8552);
xnor U9820 (N_9820,N_9300,N_9485);
or U9821 (N_9821,N_8898,N_9081);
nor U9822 (N_9822,N_9270,N_8724);
nand U9823 (N_9823,N_8532,N_8772);
nand U9824 (N_9824,N_8952,N_8605);
xnor U9825 (N_9825,N_9105,N_8615);
and U9826 (N_9826,N_8955,N_8842);
nor U9827 (N_9827,N_9263,N_8663);
and U9828 (N_9828,N_8627,N_9419);
xnor U9829 (N_9829,N_8765,N_8691);
and U9830 (N_9830,N_8639,N_9147);
nand U9831 (N_9831,N_8849,N_9594);
xor U9832 (N_9832,N_8430,N_9155);
xnor U9833 (N_9833,N_8450,N_9317);
nand U9834 (N_9834,N_8750,N_8719);
xor U9835 (N_9835,N_8528,N_8747);
and U9836 (N_9836,N_8570,N_9189);
xor U9837 (N_9837,N_9272,N_9353);
and U9838 (N_9838,N_8829,N_9523);
or U9839 (N_9839,N_8927,N_8573);
or U9840 (N_9840,N_8953,N_9374);
xor U9841 (N_9841,N_8736,N_9417);
or U9842 (N_9842,N_9486,N_8833);
nand U9843 (N_9843,N_8679,N_8807);
or U9844 (N_9844,N_9394,N_9216);
nand U9845 (N_9845,N_9273,N_9130);
nand U9846 (N_9846,N_9135,N_9073);
nand U9847 (N_9847,N_9406,N_9078);
and U9848 (N_9848,N_8978,N_9578);
xnor U9849 (N_9849,N_9290,N_8818);
nand U9850 (N_9850,N_9362,N_8774);
and U9851 (N_9851,N_8912,N_9098);
or U9852 (N_9852,N_8677,N_9595);
xnor U9853 (N_9853,N_8784,N_9166);
nor U9854 (N_9854,N_8887,N_9162);
xnor U9855 (N_9855,N_8548,N_9520);
nor U9856 (N_9856,N_9178,N_8487);
nor U9857 (N_9857,N_8414,N_9356);
nand U9858 (N_9858,N_9448,N_8619);
xor U9859 (N_9859,N_8458,N_9364);
xnor U9860 (N_9860,N_9373,N_9267);
and U9861 (N_9861,N_9013,N_9367);
xnor U9862 (N_9862,N_8419,N_8495);
nand U9863 (N_9863,N_9296,N_9301);
xnor U9864 (N_9864,N_8646,N_9392);
nor U9865 (N_9865,N_9506,N_8808);
nor U9866 (N_9866,N_8529,N_8453);
or U9867 (N_9867,N_9559,N_9357);
nor U9868 (N_9868,N_9009,N_9143);
nor U9869 (N_9869,N_8622,N_9250);
and U9870 (N_9870,N_8530,N_9324);
nand U9871 (N_9871,N_8734,N_9044);
or U9872 (N_9872,N_9083,N_8517);
xnor U9873 (N_9873,N_8895,N_8406);
nor U9874 (N_9874,N_8515,N_8553);
and U9875 (N_9875,N_8956,N_9508);
or U9876 (N_9876,N_9283,N_9442);
nor U9877 (N_9877,N_9082,N_9074);
and U9878 (N_9878,N_9154,N_8967);
xnor U9879 (N_9879,N_8568,N_8958);
or U9880 (N_9880,N_9531,N_9433);
or U9881 (N_9881,N_8526,N_9115);
xor U9882 (N_9882,N_9111,N_8623);
or U9883 (N_9883,N_8763,N_8484);
xor U9884 (N_9884,N_9100,N_9149);
nand U9885 (N_9885,N_8788,N_8449);
nor U9886 (N_9886,N_8476,N_9055);
nand U9887 (N_9887,N_8503,N_9462);
or U9888 (N_9888,N_8473,N_8432);
or U9889 (N_9889,N_9552,N_8423);
or U9890 (N_9890,N_9386,N_9495);
nand U9891 (N_9891,N_8510,N_8923);
nor U9892 (N_9892,N_9070,N_9245);
nand U9893 (N_9893,N_9592,N_8745);
xnor U9894 (N_9894,N_8970,N_8582);
nand U9895 (N_9895,N_8697,N_9388);
xor U9896 (N_9896,N_9014,N_8830);
nand U9897 (N_9897,N_9566,N_9346);
nor U9898 (N_9898,N_9534,N_9517);
xnor U9899 (N_9899,N_9415,N_9262);
nor U9900 (N_9900,N_8947,N_9106);
nor U9901 (N_9901,N_9403,N_9385);
nand U9902 (N_9902,N_9579,N_9264);
and U9903 (N_9903,N_8928,N_9472);
nand U9904 (N_9904,N_9515,N_8766);
xor U9905 (N_9905,N_8634,N_9432);
or U9906 (N_9906,N_9244,N_9102);
nand U9907 (N_9907,N_8428,N_9255);
nand U9908 (N_9908,N_8732,N_8417);
and U9909 (N_9909,N_9430,N_8888);
nor U9910 (N_9910,N_8937,N_8871);
nor U9911 (N_9911,N_8671,N_9393);
or U9912 (N_9912,N_8509,N_8931);
and U9913 (N_9913,N_9053,N_9170);
or U9914 (N_9914,N_9537,N_9184);
or U9915 (N_9915,N_9377,N_8727);
nor U9916 (N_9916,N_9434,N_9323);
or U9917 (N_9917,N_8938,N_8672);
nor U9918 (N_9918,N_8886,N_9511);
or U9919 (N_9919,N_8588,N_8680);
nand U9920 (N_9920,N_9038,N_8554);
nand U9921 (N_9921,N_8638,N_9140);
xor U9922 (N_9922,N_8498,N_9355);
or U9923 (N_9923,N_9306,N_8845);
and U9924 (N_9924,N_9124,N_9249);
and U9925 (N_9925,N_8929,N_9384);
xor U9926 (N_9926,N_9575,N_8650);
nor U9927 (N_9927,N_9243,N_9525);
or U9928 (N_9928,N_9298,N_8653);
nor U9929 (N_9929,N_8783,N_9497);
nor U9930 (N_9930,N_8980,N_8591);
nand U9931 (N_9931,N_9319,N_8564);
or U9932 (N_9932,N_9437,N_8729);
nor U9933 (N_9933,N_8993,N_8601);
nand U9934 (N_9934,N_8461,N_8466);
nor U9935 (N_9935,N_8497,N_8557);
xor U9936 (N_9936,N_9371,N_8859);
nor U9937 (N_9937,N_9054,N_9253);
and U9938 (N_9938,N_9553,N_8437);
or U9939 (N_9939,N_9209,N_8409);
and U9940 (N_9940,N_9052,N_8549);
or U9941 (N_9941,N_8725,N_8580);
nand U9942 (N_9942,N_8821,N_9092);
and U9943 (N_9943,N_9348,N_8702);
and U9944 (N_9944,N_9463,N_9252);
nand U9945 (N_9945,N_8758,N_8696);
and U9946 (N_9946,N_9591,N_9025);
nor U9947 (N_9947,N_8599,N_8604);
nand U9948 (N_9948,N_8469,N_9363);
xnor U9949 (N_9949,N_8648,N_8730);
xor U9950 (N_9950,N_9161,N_8585);
and U9951 (N_9951,N_9257,N_8984);
or U9952 (N_9952,N_9513,N_8733);
nor U9953 (N_9953,N_9413,N_8951);
nand U9954 (N_9954,N_8603,N_9366);
nor U9955 (N_9955,N_8637,N_9313);
or U9956 (N_9956,N_8802,N_8490);
xor U9957 (N_9957,N_9076,N_9046);
or U9958 (N_9958,N_8854,N_9479);
nand U9959 (N_9959,N_9282,N_9572);
and U9960 (N_9960,N_8805,N_8722);
nor U9961 (N_9961,N_9476,N_8714);
and U9962 (N_9962,N_8847,N_9458);
or U9963 (N_9963,N_8791,N_8631);
nand U9964 (N_9964,N_8785,N_8533);
and U9965 (N_9965,N_8770,N_9129);
and U9966 (N_9966,N_9037,N_8579);
nor U9967 (N_9967,N_9104,N_9164);
xor U9968 (N_9968,N_8670,N_9573);
xor U9969 (N_9969,N_9016,N_8577);
and U9970 (N_9970,N_9017,N_9361);
nand U9971 (N_9971,N_9327,N_8593);
nand U9972 (N_9972,N_8410,N_8905);
and U9973 (N_9973,N_8676,N_9312);
xnor U9974 (N_9974,N_9493,N_8584);
xnor U9975 (N_9975,N_9005,N_8906);
nor U9976 (N_9976,N_9321,N_9186);
or U9977 (N_9977,N_8431,N_8900);
or U9978 (N_9978,N_8514,N_9303);
nor U9979 (N_9979,N_8877,N_9284);
and U9980 (N_9980,N_9185,N_9401);
nand U9981 (N_9981,N_8569,N_8518);
and U9982 (N_9982,N_8640,N_9521);
or U9983 (N_9983,N_9400,N_8897);
xor U9984 (N_9984,N_9239,N_9387);
nor U9985 (N_9985,N_8472,N_8401);
nand U9986 (N_9986,N_9583,N_8616);
nand U9987 (N_9987,N_9187,N_8594);
and U9988 (N_9988,N_8768,N_8944);
nand U9989 (N_9989,N_9160,N_9507);
nand U9990 (N_9990,N_8447,N_9503);
nor U9991 (N_9991,N_9113,N_9065);
nand U9992 (N_9992,N_9341,N_8924);
nor U9993 (N_9993,N_8903,N_9136);
nand U9994 (N_9994,N_9359,N_8492);
xor U9995 (N_9995,N_8618,N_8694);
nand U9996 (N_9996,N_8926,N_9378);
or U9997 (N_9997,N_9032,N_9043);
xor U9998 (N_9998,N_9175,N_8658);
nor U9999 (N_9999,N_9133,N_9285);
nor U10000 (N_10000,N_8771,N_9271);
xnor U10001 (N_10001,N_8455,N_8987);
nor U10002 (N_10002,N_8602,N_8635);
nand U10003 (N_10003,N_9590,N_9188);
or U10004 (N_10004,N_8707,N_9121);
and U10005 (N_10005,N_9288,N_9217);
xor U10006 (N_10006,N_9488,N_8451);
nand U10007 (N_10007,N_8715,N_9126);
or U10008 (N_10008,N_8916,N_9094);
or U10009 (N_10009,N_8575,N_9444);
nand U10010 (N_10010,N_8424,N_9291);
and U10011 (N_10011,N_8494,N_8630);
or U10012 (N_10012,N_8683,N_9159);
xnor U10013 (N_10013,N_8915,N_8946);
nand U10014 (N_10014,N_8550,N_9360);
nor U10015 (N_10015,N_8481,N_9058);
nand U10016 (N_10016,N_9146,N_9469);
nor U10017 (N_10017,N_9529,N_8480);
nor U10018 (N_10018,N_8996,N_8507);
nor U10019 (N_10019,N_8426,N_9334);
or U10020 (N_10020,N_8542,N_8483);
or U10021 (N_10021,N_9201,N_8502);
and U10022 (N_10022,N_9196,N_9087);
nor U10023 (N_10023,N_8674,N_8644);
nor U10024 (N_10024,N_9555,N_8565);
nand U10025 (N_10025,N_8754,N_8705);
and U10026 (N_10026,N_9500,N_9340);
and U10027 (N_10027,N_8523,N_8983);
nor U10028 (N_10028,N_8456,N_8999);
or U10029 (N_10029,N_8420,N_9473);
xnor U10030 (N_10030,N_8434,N_9286);
xnor U10031 (N_10031,N_9086,N_9535);
nand U10032 (N_10032,N_8479,N_8718);
xor U10033 (N_10033,N_8613,N_9029);
nor U10034 (N_10034,N_9544,N_8899);
nand U10035 (N_10035,N_8445,N_9097);
nand U10036 (N_10036,N_8966,N_9438);
nand U10037 (N_10037,N_9089,N_9179);
and U10038 (N_10038,N_8841,N_9183);
or U10039 (N_10039,N_8834,N_8741);
and U10040 (N_10040,N_8738,N_9047);
or U10041 (N_10041,N_8686,N_8907);
or U10042 (N_10042,N_9416,N_8933);
and U10043 (N_10043,N_9402,N_9010);
nand U10044 (N_10044,N_9071,N_8839);
xnor U10045 (N_10045,N_8649,N_9227);
nor U10046 (N_10046,N_8486,N_9439);
nand U10047 (N_10047,N_9554,N_9467);
xor U10048 (N_10048,N_8776,N_9471);
nor U10049 (N_10049,N_9397,N_9532);
xor U10050 (N_10050,N_9428,N_8780);
nand U10051 (N_10051,N_9315,N_9494);
or U10052 (N_10052,N_8812,N_8433);
xnor U10053 (N_10053,N_8932,N_9424);
xnor U10054 (N_10054,N_8690,N_8748);
or U10055 (N_10055,N_8942,N_8832);
xnor U10056 (N_10056,N_9568,N_8976);
nand U10057 (N_10057,N_9173,N_8411);
and U10058 (N_10058,N_8654,N_9562);
xnor U10059 (N_10059,N_9358,N_9019);
nand U10060 (N_10060,N_9134,N_9072);
nand U10061 (N_10061,N_9040,N_9148);
and U10062 (N_10062,N_9181,N_8836);
and U10063 (N_10063,N_8828,N_8624);
nor U10064 (N_10064,N_8563,N_8659);
and U10065 (N_10065,N_8972,N_9000);
and U10066 (N_10066,N_9062,N_9015);
or U10067 (N_10067,N_8817,N_8868);
or U10068 (N_10068,N_8767,N_9441);
xnor U10069 (N_10069,N_8757,N_9001);
xor U10070 (N_10070,N_8794,N_9171);
nor U10071 (N_10071,N_9214,N_9141);
and U10072 (N_10072,N_9247,N_9536);
and U10073 (N_10073,N_8460,N_9538);
nor U10074 (N_10074,N_9061,N_8998);
xnor U10075 (N_10075,N_8534,N_8746);
xor U10076 (N_10076,N_9077,N_9560);
nand U10077 (N_10077,N_8402,N_9281);
or U10078 (N_10078,N_9561,N_9347);
or U10079 (N_10079,N_8720,N_8462);
nand U10080 (N_10080,N_8700,N_8994);
and U10081 (N_10081,N_9127,N_8731);
xnor U10082 (N_10082,N_9219,N_9304);
nor U10083 (N_10083,N_8764,N_8823);
and U10084 (N_10084,N_9050,N_8974);
xor U10085 (N_10085,N_9499,N_8600);
xnor U10086 (N_10086,N_8609,N_8543);
or U10087 (N_10087,N_8673,N_9168);
nand U10088 (N_10088,N_9193,N_8930);
nand U10089 (N_10089,N_9398,N_8751);
nor U10090 (N_10090,N_8796,N_9258);
xnor U10091 (N_10091,N_9580,N_8943);
and U10092 (N_10092,N_9256,N_9006);
nand U10093 (N_10093,N_8755,N_8779);
nand U10094 (N_10094,N_8665,N_8777);
nand U10095 (N_10095,N_8675,N_8596);
and U10096 (N_10096,N_8716,N_9587);
xor U10097 (N_10097,N_8909,N_9177);
xnor U10098 (N_10098,N_9465,N_8894);
or U10099 (N_10099,N_9581,N_8664);
or U10100 (N_10100,N_8551,N_9466);
nor U10101 (N_10101,N_8848,N_9063);
and U10102 (N_10102,N_8838,N_9445);
xnor U10103 (N_10103,N_9551,N_9199);
nand U10104 (N_10104,N_9266,N_8701);
nor U10105 (N_10105,N_9174,N_9228);
nor U10106 (N_10106,N_8919,N_9069);
nor U10107 (N_10107,N_9067,N_9548);
nand U10108 (N_10108,N_9574,N_8959);
or U10109 (N_10109,N_8500,N_8708);
nand U10110 (N_10110,N_9123,N_8520);
or U10111 (N_10111,N_8973,N_8403);
xor U10112 (N_10112,N_9254,N_8873);
nor U10113 (N_10113,N_9326,N_8890);
or U10114 (N_10114,N_8583,N_9343);
nor U10115 (N_10115,N_9504,N_8921);
nor U10116 (N_10116,N_9459,N_8792);
xnor U10117 (N_10117,N_8852,N_8489);
nor U10118 (N_10118,N_8816,N_8541);
xor U10119 (N_10119,N_8571,N_9204);
and U10120 (N_10120,N_8762,N_9329);
and U10121 (N_10121,N_8558,N_9246);
xnor U10122 (N_10122,N_9491,N_9278);
nor U10123 (N_10123,N_8710,N_8773);
xnor U10124 (N_10124,N_8682,N_8866);
nor U10125 (N_10125,N_8547,N_8945);
and U10126 (N_10126,N_9586,N_8795);
xnor U10127 (N_10127,N_8872,N_9236);
nand U10128 (N_10128,N_9565,N_8400);
or U10129 (N_10129,N_8819,N_8949);
nand U10130 (N_10130,N_8902,N_8452);
or U10131 (N_10131,N_8448,N_8636);
or U10132 (N_10132,N_8793,N_9496);
and U10133 (N_10133,N_9165,N_8885);
and U10134 (N_10134,N_9090,N_8407);
or U10135 (N_10135,N_8590,N_9297);
and U10136 (N_10136,N_9379,N_9404);
xor U10137 (N_10137,N_8572,N_9235);
and U10138 (N_10138,N_9446,N_9426);
and U10139 (N_10139,N_9563,N_8454);
nor U10140 (N_10140,N_9350,N_9336);
and U10141 (N_10141,N_8728,N_9180);
xor U10142 (N_10142,N_8666,N_8482);
and U10143 (N_10143,N_9120,N_8712);
and U10144 (N_10144,N_8703,N_8499);
or U10145 (N_10145,N_8562,N_8478);
nand U10146 (N_10146,N_9410,N_9344);
nand U10147 (N_10147,N_8576,N_8986);
nand U10148 (N_10148,N_9118,N_9157);
xnor U10149 (N_10149,N_8824,N_8815);
and U10150 (N_10150,N_9049,N_9215);
nand U10151 (N_10151,N_8442,N_9293);
nor U10152 (N_10152,N_9200,N_8876);
and U10153 (N_10153,N_8652,N_9408);
nand U10154 (N_10154,N_9376,N_8985);
nand U10155 (N_10155,N_8440,N_8761);
xnor U10156 (N_10156,N_8595,N_8896);
and U10157 (N_10157,N_8516,N_8404);
xor U10158 (N_10158,N_9066,N_9208);
and U10159 (N_10159,N_9481,N_9042);
or U10160 (N_10160,N_9420,N_8726);
nor U10161 (N_10161,N_9237,N_8981);
nor U10162 (N_10162,N_8611,N_8721);
nand U10163 (N_10163,N_8911,N_8581);
nand U10164 (N_10164,N_8681,N_8737);
and U10165 (N_10165,N_9259,N_8457);
nand U10166 (N_10166,N_9218,N_9539);
nor U10167 (N_10167,N_8614,N_9519);
xnor U10168 (N_10168,N_9210,N_8668);
xnor U10169 (N_10169,N_9440,N_8743);
nand U10170 (N_10170,N_8405,N_8975);
nand U10171 (N_10171,N_8997,N_8689);
nand U10172 (N_10172,N_9021,N_9242);
or U10173 (N_10173,N_8826,N_8811);
nand U10174 (N_10174,N_9451,N_8560);
xor U10175 (N_10175,N_8969,N_8471);
xnor U10176 (N_10176,N_8459,N_8512);
and U10177 (N_10177,N_8713,N_9522);
xnor U10178 (N_10178,N_8441,N_9318);
xor U10179 (N_10179,N_8756,N_8506);
nand U10180 (N_10180,N_8545,N_8851);
xnor U10181 (N_10181,N_8740,N_8917);
or U10182 (N_10182,N_9435,N_8625);
and U10183 (N_10183,N_9457,N_9169);
nor U10184 (N_10184,N_9080,N_8856);
nor U10185 (N_10185,N_9114,N_8513);
xnor U10186 (N_10186,N_8629,N_8574);
xor U10187 (N_10187,N_9045,N_9474);
or U10188 (N_10188,N_8865,N_9051);
and U10189 (N_10189,N_8904,N_9125);
and U10190 (N_10190,N_8669,N_8884);
xor U10191 (N_10191,N_8643,N_8505);
and U10192 (N_10192,N_8475,N_8910);
xor U10193 (N_10193,N_8759,N_8968);
and U10194 (N_10194,N_8846,N_8717);
nand U10195 (N_10195,N_9012,N_9498);
nand U10196 (N_10196,N_8813,N_9128);
nand U10197 (N_10197,N_8863,N_8810);
or U10198 (N_10198,N_9103,N_9314);
and U10199 (N_10199,N_9354,N_9598);
or U10200 (N_10200,N_9497,N_8980);
or U10201 (N_10201,N_8485,N_8653);
or U10202 (N_10202,N_9417,N_9560);
xor U10203 (N_10203,N_8951,N_9221);
nand U10204 (N_10204,N_9305,N_8908);
nand U10205 (N_10205,N_9474,N_8657);
nor U10206 (N_10206,N_9451,N_8718);
nand U10207 (N_10207,N_9000,N_8894);
xor U10208 (N_10208,N_8835,N_8544);
xnor U10209 (N_10209,N_8819,N_8571);
nand U10210 (N_10210,N_9058,N_8764);
xnor U10211 (N_10211,N_8982,N_9058);
or U10212 (N_10212,N_8942,N_8548);
nand U10213 (N_10213,N_8464,N_8981);
nand U10214 (N_10214,N_8886,N_8932);
and U10215 (N_10215,N_8882,N_8542);
nor U10216 (N_10216,N_8853,N_9386);
or U10217 (N_10217,N_9549,N_9459);
and U10218 (N_10218,N_8569,N_9433);
xor U10219 (N_10219,N_8401,N_9363);
and U10220 (N_10220,N_9347,N_8661);
nand U10221 (N_10221,N_9466,N_8667);
xnor U10222 (N_10222,N_8538,N_9400);
or U10223 (N_10223,N_8465,N_9520);
xor U10224 (N_10224,N_9057,N_8608);
nand U10225 (N_10225,N_9437,N_9418);
nand U10226 (N_10226,N_9522,N_8854);
or U10227 (N_10227,N_9219,N_9203);
nand U10228 (N_10228,N_9215,N_8965);
xnor U10229 (N_10229,N_8656,N_8512);
or U10230 (N_10230,N_8949,N_8725);
or U10231 (N_10231,N_8429,N_8543);
or U10232 (N_10232,N_9519,N_9526);
nor U10233 (N_10233,N_9468,N_9058);
or U10234 (N_10234,N_9286,N_8675);
xnor U10235 (N_10235,N_8868,N_9028);
or U10236 (N_10236,N_9055,N_9368);
or U10237 (N_10237,N_8743,N_9413);
and U10238 (N_10238,N_9145,N_9560);
xnor U10239 (N_10239,N_8958,N_8466);
and U10240 (N_10240,N_8536,N_8700);
and U10241 (N_10241,N_8753,N_9348);
and U10242 (N_10242,N_9104,N_8400);
and U10243 (N_10243,N_9274,N_9154);
xnor U10244 (N_10244,N_9345,N_8554);
nand U10245 (N_10245,N_9576,N_8453);
or U10246 (N_10246,N_8891,N_8835);
xnor U10247 (N_10247,N_8860,N_9378);
or U10248 (N_10248,N_8830,N_9030);
or U10249 (N_10249,N_9067,N_8515);
nor U10250 (N_10250,N_9193,N_9034);
or U10251 (N_10251,N_9334,N_9085);
nor U10252 (N_10252,N_9438,N_9209);
nand U10253 (N_10253,N_9103,N_9443);
xnor U10254 (N_10254,N_9081,N_8852);
nand U10255 (N_10255,N_8585,N_8768);
and U10256 (N_10256,N_8574,N_9553);
or U10257 (N_10257,N_9520,N_8662);
nand U10258 (N_10258,N_9288,N_9475);
nor U10259 (N_10259,N_9457,N_8528);
or U10260 (N_10260,N_8644,N_8817);
nand U10261 (N_10261,N_8521,N_8941);
xor U10262 (N_10262,N_8805,N_9373);
or U10263 (N_10263,N_9431,N_8924);
and U10264 (N_10264,N_9354,N_8930);
or U10265 (N_10265,N_8816,N_9546);
and U10266 (N_10266,N_9354,N_9448);
or U10267 (N_10267,N_9130,N_9054);
and U10268 (N_10268,N_9299,N_9529);
nor U10269 (N_10269,N_9493,N_9205);
or U10270 (N_10270,N_8477,N_9092);
and U10271 (N_10271,N_9080,N_8985);
nor U10272 (N_10272,N_9251,N_9485);
xor U10273 (N_10273,N_8647,N_9072);
xor U10274 (N_10274,N_8939,N_9578);
nor U10275 (N_10275,N_8829,N_9562);
xor U10276 (N_10276,N_8791,N_9025);
xor U10277 (N_10277,N_8532,N_8739);
or U10278 (N_10278,N_9126,N_8695);
nand U10279 (N_10279,N_8641,N_8918);
and U10280 (N_10280,N_8758,N_9558);
and U10281 (N_10281,N_8422,N_8581);
nand U10282 (N_10282,N_8841,N_8741);
and U10283 (N_10283,N_9393,N_8590);
or U10284 (N_10284,N_8988,N_8426);
xor U10285 (N_10285,N_9306,N_9023);
nor U10286 (N_10286,N_9377,N_9064);
xor U10287 (N_10287,N_8436,N_8411);
and U10288 (N_10288,N_8546,N_9242);
and U10289 (N_10289,N_9204,N_8892);
nor U10290 (N_10290,N_9502,N_8429);
xor U10291 (N_10291,N_8898,N_8405);
and U10292 (N_10292,N_8897,N_8711);
nor U10293 (N_10293,N_9242,N_8468);
and U10294 (N_10294,N_8426,N_9599);
and U10295 (N_10295,N_8854,N_8838);
nor U10296 (N_10296,N_9115,N_9347);
and U10297 (N_10297,N_9162,N_8646);
nand U10298 (N_10298,N_8817,N_9367);
or U10299 (N_10299,N_8728,N_9129);
xnor U10300 (N_10300,N_8758,N_8545);
or U10301 (N_10301,N_8433,N_9239);
or U10302 (N_10302,N_8846,N_8715);
xnor U10303 (N_10303,N_9366,N_9136);
nand U10304 (N_10304,N_8988,N_9269);
or U10305 (N_10305,N_9145,N_8719);
xnor U10306 (N_10306,N_9147,N_8787);
nand U10307 (N_10307,N_8938,N_8516);
nand U10308 (N_10308,N_9401,N_9464);
nor U10309 (N_10309,N_8579,N_8514);
xnor U10310 (N_10310,N_8497,N_8646);
xor U10311 (N_10311,N_9423,N_8722);
nand U10312 (N_10312,N_8587,N_9296);
nand U10313 (N_10313,N_9069,N_9071);
xnor U10314 (N_10314,N_9448,N_9072);
or U10315 (N_10315,N_8460,N_9515);
nor U10316 (N_10316,N_8942,N_9113);
nand U10317 (N_10317,N_8590,N_8626);
or U10318 (N_10318,N_9107,N_9077);
or U10319 (N_10319,N_9476,N_9439);
or U10320 (N_10320,N_9559,N_8957);
and U10321 (N_10321,N_8870,N_9226);
nor U10322 (N_10322,N_9401,N_9142);
or U10323 (N_10323,N_9291,N_9553);
or U10324 (N_10324,N_8412,N_8504);
and U10325 (N_10325,N_9427,N_8738);
nand U10326 (N_10326,N_8932,N_9191);
xor U10327 (N_10327,N_9552,N_9187);
nand U10328 (N_10328,N_8775,N_9250);
nor U10329 (N_10329,N_8885,N_8741);
and U10330 (N_10330,N_8792,N_8788);
nand U10331 (N_10331,N_9581,N_8449);
nor U10332 (N_10332,N_9026,N_8706);
nand U10333 (N_10333,N_8407,N_8520);
or U10334 (N_10334,N_8532,N_8914);
nand U10335 (N_10335,N_8931,N_9354);
nand U10336 (N_10336,N_9234,N_9496);
nand U10337 (N_10337,N_8791,N_9110);
xnor U10338 (N_10338,N_8929,N_8876);
nor U10339 (N_10339,N_8764,N_8958);
and U10340 (N_10340,N_8688,N_8737);
nor U10341 (N_10341,N_8813,N_9278);
nor U10342 (N_10342,N_8454,N_8788);
xor U10343 (N_10343,N_9396,N_9411);
xnor U10344 (N_10344,N_9473,N_9131);
xor U10345 (N_10345,N_9123,N_9498);
nand U10346 (N_10346,N_9285,N_8686);
and U10347 (N_10347,N_9364,N_8803);
nor U10348 (N_10348,N_9222,N_8637);
nand U10349 (N_10349,N_9474,N_8614);
and U10350 (N_10350,N_8934,N_9533);
nor U10351 (N_10351,N_9385,N_9053);
xor U10352 (N_10352,N_9480,N_8737);
xor U10353 (N_10353,N_8577,N_8472);
nor U10354 (N_10354,N_8834,N_8484);
nand U10355 (N_10355,N_8670,N_8623);
nor U10356 (N_10356,N_8854,N_9049);
and U10357 (N_10357,N_9280,N_8913);
nor U10358 (N_10358,N_8532,N_9224);
nor U10359 (N_10359,N_9492,N_9457);
nor U10360 (N_10360,N_9467,N_9063);
nor U10361 (N_10361,N_9255,N_9268);
xor U10362 (N_10362,N_9535,N_9571);
xnor U10363 (N_10363,N_8668,N_8921);
xor U10364 (N_10364,N_8824,N_8844);
and U10365 (N_10365,N_8857,N_9466);
nor U10366 (N_10366,N_9199,N_9268);
and U10367 (N_10367,N_9534,N_9335);
nand U10368 (N_10368,N_8433,N_8743);
and U10369 (N_10369,N_8404,N_9382);
or U10370 (N_10370,N_9579,N_9524);
nand U10371 (N_10371,N_9239,N_8897);
nand U10372 (N_10372,N_8746,N_8937);
xor U10373 (N_10373,N_8443,N_9038);
and U10374 (N_10374,N_9511,N_9284);
and U10375 (N_10375,N_8469,N_9474);
nand U10376 (N_10376,N_8860,N_8720);
or U10377 (N_10377,N_8730,N_8908);
nand U10378 (N_10378,N_9423,N_9115);
nand U10379 (N_10379,N_9477,N_8775);
or U10380 (N_10380,N_9144,N_8664);
nand U10381 (N_10381,N_8811,N_9240);
or U10382 (N_10382,N_9217,N_8401);
xnor U10383 (N_10383,N_9274,N_8884);
xnor U10384 (N_10384,N_8825,N_8828);
or U10385 (N_10385,N_8837,N_8671);
or U10386 (N_10386,N_9051,N_9366);
or U10387 (N_10387,N_9046,N_8638);
xor U10388 (N_10388,N_8640,N_8833);
and U10389 (N_10389,N_8860,N_9515);
or U10390 (N_10390,N_8662,N_8633);
nor U10391 (N_10391,N_8788,N_9091);
nand U10392 (N_10392,N_9259,N_9426);
nand U10393 (N_10393,N_8472,N_9311);
or U10394 (N_10394,N_9241,N_9117);
xor U10395 (N_10395,N_9173,N_9201);
nor U10396 (N_10396,N_8615,N_9131);
nor U10397 (N_10397,N_8523,N_9429);
nor U10398 (N_10398,N_8691,N_8797);
nand U10399 (N_10399,N_8508,N_9257);
nand U10400 (N_10400,N_8922,N_8598);
nor U10401 (N_10401,N_8452,N_8561);
nand U10402 (N_10402,N_8423,N_9316);
or U10403 (N_10403,N_9075,N_9574);
nand U10404 (N_10404,N_8807,N_9479);
or U10405 (N_10405,N_8844,N_9385);
nor U10406 (N_10406,N_9472,N_9032);
xnor U10407 (N_10407,N_9018,N_9560);
or U10408 (N_10408,N_8404,N_9236);
nor U10409 (N_10409,N_8794,N_9192);
and U10410 (N_10410,N_9330,N_8622);
and U10411 (N_10411,N_8569,N_8478);
nand U10412 (N_10412,N_8654,N_8553);
or U10413 (N_10413,N_8711,N_8994);
nand U10414 (N_10414,N_9153,N_9186);
or U10415 (N_10415,N_9482,N_9472);
or U10416 (N_10416,N_8552,N_9130);
and U10417 (N_10417,N_8489,N_9154);
and U10418 (N_10418,N_8647,N_8525);
nand U10419 (N_10419,N_9145,N_9400);
and U10420 (N_10420,N_9155,N_8816);
and U10421 (N_10421,N_9074,N_9127);
and U10422 (N_10422,N_9524,N_9081);
or U10423 (N_10423,N_8996,N_9089);
or U10424 (N_10424,N_8799,N_9517);
or U10425 (N_10425,N_9082,N_9286);
nor U10426 (N_10426,N_9130,N_9381);
xor U10427 (N_10427,N_9330,N_9213);
and U10428 (N_10428,N_9137,N_9207);
and U10429 (N_10429,N_9357,N_9519);
nor U10430 (N_10430,N_8976,N_8486);
or U10431 (N_10431,N_8414,N_8659);
nand U10432 (N_10432,N_8677,N_9330);
nor U10433 (N_10433,N_8656,N_9415);
nand U10434 (N_10434,N_8880,N_8593);
xor U10435 (N_10435,N_8859,N_8704);
nor U10436 (N_10436,N_8912,N_9334);
nand U10437 (N_10437,N_9047,N_8469);
nand U10438 (N_10438,N_8996,N_9195);
xnor U10439 (N_10439,N_9518,N_8989);
nand U10440 (N_10440,N_8976,N_9428);
nor U10441 (N_10441,N_9573,N_9019);
nand U10442 (N_10442,N_9307,N_9558);
xor U10443 (N_10443,N_8861,N_9542);
xor U10444 (N_10444,N_9462,N_8697);
and U10445 (N_10445,N_9273,N_8916);
nand U10446 (N_10446,N_8701,N_8781);
and U10447 (N_10447,N_8853,N_9042);
xor U10448 (N_10448,N_8850,N_9349);
nand U10449 (N_10449,N_8416,N_8975);
nor U10450 (N_10450,N_8942,N_9224);
nor U10451 (N_10451,N_9532,N_9159);
xor U10452 (N_10452,N_8824,N_8883);
nor U10453 (N_10453,N_9256,N_9498);
nand U10454 (N_10454,N_8440,N_8682);
xnor U10455 (N_10455,N_9408,N_8807);
and U10456 (N_10456,N_9589,N_8430);
and U10457 (N_10457,N_9247,N_8843);
and U10458 (N_10458,N_9236,N_8864);
xor U10459 (N_10459,N_9131,N_9010);
and U10460 (N_10460,N_9369,N_9465);
or U10461 (N_10461,N_8632,N_8865);
or U10462 (N_10462,N_8893,N_8544);
nand U10463 (N_10463,N_8890,N_8920);
or U10464 (N_10464,N_8446,N_8574);
or U10465 (N_10465,N_8487,N_8929);
xnor U10466 (N_10466,N_8571,N_9557);
and U10467 (N_10467,N_9076,N_8848);
or U10468 (N_10468,N_8602,N_9068);
or U10469 (N_10469,N_8516,N_9204);
xnor U10470 (N_10470,N_8674,N_8889);
nor U10471 (N_10471,N_8598,N_8880);
nor U10472 (N_10472,N_8891,N_9073);
nand U10473 (N_10473,N_8999,N_8738);
and U10474 (N_10474,N_8488,N_8792);
nor U10475 (N_10475,N_8716,N_9459);
or U10476 (N_10476,N_9380,N_9442);
and U10477 (N_10477,N_9412,N_9371);
and U10478 (N_10478,N_9283,N_9333);
or U10479 (N_10479,N_9361,N_9102);
and U10480 (N_10480,N_9159,N_8777);
nor U10481 (N_10481,N_9397,N_8888);
or U10482 (N_10482,N_8702,N_9171);
nand U10483 (N_10483,N_9372,N_9282);
and U10484 (N_10484,N_8555,N_8606);
nor U10485 (N_10485,N_9466,N_8961);
xor U10486 (N_10486,N_8614,N_9372);
xor U10487 (N_10487,N_8885,N_8793);
and U10488 (N_10488,N_8690,N_8749);
nand U10489 (N_10489,N_8737,N_9030);
nand U10490 (N_10490,N_8423,N_8570);
or U10491 (N_10491,N_9532,N_8750);
or U10492 (N_10492,N_9141,N_8831);
and U10493 (N_10493,N_9283,N_8839);
nor U10494 (N_10494,N_9362,N_8729);
or U10495 (N_10495,N_9319,N_8754);
nor U10496 (N_10496,N_8453,N_9400);
nand U10497 (N_10497,N_9597,N_9060);
and U10498 (N_10498,N_8536,N_8611);
and U10499 (N_10499,N_9395,N_9036);
and U10500 (N_10500,N_9220,N_9519);
or U10501 (N_10501,N_8896,N_8519);
or U10502 (N_10502,N_8818,N_8646);
nand U10503 (N_10503,N_8676,N_9243);
nor U10504 (N_10504,N_9167,N_8400);
nor U10505 (N_10505,N_8688,N_8791);
nand U10506 (N_10506,N_9062,N_9006);
and U10507 (N_10507,N_9557,N_8947);
or U10508 (N_10508,N_9036,N_8860);
nor U10509 (N_10509,N_9366,N_9277);
nor U10510 (N_10510,N_9195,N_9504);
and U10511 (N_10511,N_8533,N_9176);
or U10512 (N_10512,N_9479,N_9161);
nand U10513 (N_10513,N_9261,N_9528);
nand U10514 (N_10514,N_8895,N_9032);
nor U10515 (N_10515,N_9413,N_9078);
or U10516 (N_10516,N_8601,N_9319);
nor U10517 (N_10517,N_9046,N_8596);
and U10518 (N_10518,N_9019,N_9434);
nor U10519 (N_10519,N_8403,N_8522);
nand U10520 (N_10520,N_9046,N_8521);
and U10521 (N_10521,N_9553,N_9098);
xor U10522 (N_10522,N_8684,N_8521);
nand U10523 (N_10523,N_9419,N_8979);
nor U10524 (N_10524,N_8699,N_8731);
and U10525 (N_10525,N_8411,N_9362);
and U10526 (N_10526,N_9087,N_9450);
nor U10527 (N_10527,N_8669,N_9484);
and U10528 (N_10528,N_9060,N_9325);
or U10529 (N_10529,N_9549,N_8952);
or U10530 (N_10530,N_8450,N_8526);
nand U10531 (N_10531,N_9257,N_9577);
xor U10532 (N_10532,N_9348,N_9560);
xor U10533 (N_10533,N_8766,N_9361);
nor U10534 (N_10534,N_9426,N_9072);
or U10535 (N_10535,N_9594,N_8706);
and U10536 (N_10536,N_9504,N_8903);
xor U10537 (N_10537,N_8502,N_9285);
xor U10538 (N_10538,N_8898,N_9493);
nor U10539 (N_10539,N_9168,N_8737);
nand U10540 (N_10540,N_8428,N_8704);
xnor U10541 (N_10541,N_8589,N_8708);
xor U10542 (N_10542,N_8914,N_8625);
nor U10543 (N_10543,N_9225,N_9426);
or U10544 (N_10544,N_9106,N_8547);
nor U10545 (N_10545,N_9440,N_8500);
nor U10546 (N_10546,N_8711,N_8676);
nor U10547 (N_10547,N_8485,N_9230);
nand U10548 (N_10548,N_8621,N_9519);
nand U10549 (N_10549,N_8972,N_9385);
nand U10550 (N_10550,N_9198,N_8778);
or U10551 (N_10551,N_9389,N_8507);
nor U10552 (N_10552,N_9189,N_9223);
nor U10553 (N_10553,N_8690,N_9396);
xor U10554 (N_10554,N_9342,N_8874);
and U10555 (N_10555,N_8999,N_8654);
nand U10556 (N_10556,N_8790,N_8668);
xnor U10557 (N_10557,N_8569,N_8870);
nand U10558 (N_10558,N_8436,N_9138);
xor U10559 (N_10559,N_9584,N_8666);
xnor U10560 (N_10560,N_9102,N_8643);
and U10561 (N_10561,N_9499,N_8816);
xor U10562 (N_10562,N_9314,N_9485);
xor U10563 (N_10563,N_9408,N_9159);
nand U10564 (N_10564,N_8956,N_9337);
xnor U10565 (N_10565,N_9030,N_8817);
xnor U10566 (N_10566,N_8438,N_8637);
and U10567 (N_10567,N_8652,N_8762);
nor U10568 (N_10568,N_9572,N_8445);
or U10569 (N_10569,N_9270,N_8592);
nand U10570 (N_10570,N_8793,N_8747);
xnor U10571 (N_10571,N_9287,N_9204);
nor U10572 (N_10572,N_8954,N_8719);
nor U10573 (N_10573,N_8929,N_9317);
nand U10574 (N_10574,N_8987,N_8930);
xor U10575 (N_10575,N_9175,N_8789);
nand U10576 (N_10576,N_9088,N_8504);
or U10577 (N_10577,N_9054,N_8614);
xor U10578 (N_10578,N_8880,N_8983);
and U10579 (N_10579,N_9218,N_8440);
xnor U10580 (N_10580,N_9058,N_8765);
and U10581 (N_10581,N_9109,N_9323);
nand U10582 (N_10582,N_9335,N_8566);
xnor U10583 (N_10583,N_9191,N_8683);
nor U10584 (N_10584,N_9258,N_8832);
and U10585 (N_10585,N_8880,N_9092);
or U10586 (N_10586,N_8408,N_8618);
xnor U10587 (N_10587,N_8751,N_8890);
nor U10588 (N_10588,N_9028,N_9116);
nor U10589 (N_10589,N_8694,N_9220);
and U10590 (N_10590,N_8917,N_8923);
xor U10591 (N_10591,N_9309,N_9496);
or U10592 (N_10592,N_9522,N_9432);
xnor U10593 (N_10593,N_8820,N_9177);
or U10594 (N_10594,N_9426,N_9358);
and U10595 (N_10595,N_9365,N_9448);
and U10596 (N_10596,N_8420,N_8783);
and U10597 (N_10597,N_8571,N_9359);
or U10598 (N_10598,N_9525,N_8507);
and U10599 (N_10599,N_8958,N_9126);
nand U10600 (N_10600,N_9324,N_8944);
and U10601 (N_10601,N_8699,N_9164);
nand U10602 (N_10602,N_9176,N_9374);
xor U10603 (N_10603,N_9124,N_9240);
or U10604 (N_10604,N_8439,N_9019);
and U10605 (N_10605,N_8751,N_8746);
and U10606 (N_10606,N_8456,N_8667);
nand U10607 (N_10607,N_8936,N_9127);
nand U10608 (N_10608,N_9441,N_8931);
or U10609 (N_10609,N_8846,N_9406);
and U10610 (N_10610,N_8812,N_9494);
xor U10611 (N_10611,N_8701,N_9217);
nor U10612 (N_10612,N_8835,N_9409);
and U10613 (N_10613,N_9257,N_9272);
nor U10614 (N_10614,N_9150,N_8875);
or U10615 (N_10615,N_8505,N_9050);
or U10616 (N_10616,N_8973,N_9029);
or U10617 (N_10617,N_8524,N_9416);
nand U10618 (N_10618,N_9283,N_8877);
xor U10619 (N_10619,N_9364,N_9305);
nand U10620 (N_10620,N_9241,N_8905);
nand U10621 (N_10621,N_8878,N_9074);
and U10622 (N_10622,N_9121,N_9302);
or U10623 (N_10623,N_8722,N_8687);
nor U10624 (N_10624,N_8806,N_9247);
xor U10625 (N_10625,N_8567,N_8498);
or U10626 (N_10626,N_8645,N_9064);
nor U10627 (N_10627,N_9190,N_8901);
nand U10628 (N_10628,N_9272,N_8676);
or U10629 (N_10629,N_8835,N_9197);
or U10630 (N_10630,N_8984,N_9350);
and U10631 (N_10631,N_9069,N_8618);
or U10632 (N_10632,N_9388,N_9151);
nor U10633 (N_10633,N_8680,N_8440);
and U10634 (N_10634,N_8743,N_9098);
and U10635 (N_10635,N_8782,N_8557);
and U10636 (N_10636,N_8849,N_9203);
and U10637 (N_10637,N_8861,N_9138);
and U10638 (N_10638,N_8832,N_8619);
nand U10639 (N_10639,N_9505,N_8741);
nor U10640 (N_10640,N_9357,N_9270);
and U10641 (N_10641,N_8843,N_8731);
or U10642 (N_10642,N_9553,N_9049);
nor U10643 (N_10643,N_8997,N_8478);
nand U10644 (N_10644,N_9094,N_8430);
and U10645 (N_10645,N_9480,N_8608);
xnor U10646 (N_10646,N_9312,N_8449);
nand U10647 (N_10647,N_8974,N_8503);
and U10648 (N_10648,N_8839,N_9169);
xnor U10649 (N_10649,N_9295,N_9120);
and U10650 (N_10650,N_9368,N_8722);
nand U10651 (N_10651,N_8688,N_8730);
nor U10652 (N_10652,N_8439,N_8722);
xor U10653 (N_10653,N_8958,N_8477);
nand U10654 (N_10654,N_9188,N_8670);
and U10655 (N_10655,N_9197,N_8805);
nand U10656 (N_10656,N_8659,N_9218);
xnor U10657 (N_10657,N_8804,N_9205);
and U10658 (N_10658,N_8687,N_8850);
and U10659 (N_10659,N_9048,N_8820);
nor U10660 (N_10660,N_8623,N_9178);
or U10661 (N_10661,N_8439,N_8655);
nand U10662 (N_10662,N_9038,N_9148);
nand U10663 (N_10663,N_9536,N_8991);
nor U10664 (N_10664,N_9119,N_8405);
and U10665 (N_10665,N_9407,N_9179);
nand U10666 (N_10666,N_9549,N_8648);
xnor U10667 (N_10667,N_8718,N_8605);
or U10668 (N_10668,N_8493,N_8574);
xnor U10669 (N_10669,N_9475,N_9363);
and U10670 (N_10670,N_8833,N_8630);
and U10671 (N_10671,N_8942,N_8803);
or U10672 (N_10672,N_9291,N_8661);
xnor U10673 (N_10673,N_9390,N_9280);
xnor U10674 (N_10674,N_9518,N_9452);
nand U10675 (N_10675,N_8634,N_8804);
and U10676 (N_10676,N_9149,N_8551);
or U10677 (N_10677,N_8726,N_8872);
nand U10678 (N_10678,N_9012,N_9305);
and U10679 (N_10679,N_8565,N_9570);
nand U10680 (N_10680,N_8615,N_8469);
nand U10681 (N_10681,N_8467,N_8662);
nand U10682 (N_10682,N_9399,N_8440);
or U10683 (N_10683,N_9209,N_9192);
or U10684 (N_10684,N_8550,N_8427);
or U10685 (N_10685,N_9210,N_8844);
xor U10686 (N_10686,N_8845,N_9187);
nand U10687 (N_10687,N_8639,N_9034);
or U10688 (N_10688,N_9543,N_9060);
and U10689 (N_10689,N_9385,N_9286);
nand U10690 (N_10690,N_9062,N_8874);
nor U10691 (N_10691,N_9406,N_9536);
nor U10692 (N_10692,N_8520,N_9538);
xnor U10693 (N_10693,N_8642,N_8685);
and U10694 (N_10694,N_8671,N_9114);
nand U10695 (N_10695,N_8839,N_8414);
nor U10696 (N_10696,N_8899,N_8776);
and U10697 (N_10697,N_9126,N_8700);
or U10698 (N_10698,N_8685,N_9317);
xor U10699 (N_10699,N_8423,N_9260);
and U10700 (N_10700,N_8520,N_8793);
and U10701 (N_10701,N_8531,N_8964);
or U10702 (N_10702,N_9159,N_8718);
xor U10703 (N_10703,N_8591,N_9316);
nor U10704 (N_10704,N_9591,N_8760);
or U10705 (N_10705,N_9290,N_8889);
xor U10706 (N_10706,N_8428,N_8534);
xor U10707 (N_10707,N_8523,N_8645);
xnor U10708 (N_10708,N_9465,N_9195);
and U10709 (N_10709,N_8747,N_9049);
nand U10710 (N_10710,N_9387,N_9222);
nand U10711 (N_10711,N_8993,N_9191);
and U10712 (N_10712,N_9401,N_8441);
nor U10713 (N_10713,N_8830,N_9208);
or U10714 (N_10714,N_8799,N_9107);
xnor U10715 (N_10715,N_9287,N_9564);
xnor U10716 (N_10716,N_8887,N_8992);
or U10717 (N_10717,N_9479,N_8988);
and U10718 (N_10718,N_8994,N_9279);
nand U10719 (N_10719,N_9242,N_9305);
and U10720 (N_10720,N_8786,N_9376);
and U10721 (N_10721,N_8488,N_8943);
or U10722 (N_10722,N_8892,N_8992);
nor U10723 (N_10723,N_9239,N_8580);
or U10724 (N_10724,N_9284,N_9309);
or U10725 (N_10725,N_9089,N_8756);
xnor U10726 (N_10726,N_9143,N_9047);
and U10727 (N_10727,N_8693,N_8460);
or U10728 (N_10728,N_9401,N_8611);
nor U10729 (N_10729,N_8919,N_9136);
or U10730 (N_10730,N_9488,N_8598);
xor U10731 (N_10731,N_9525,N_9331);
and U10732 (N_10732,N_9102,N_8863);
nand U10733 (N_10733,N_9553,N_9378);
nor U10734 (N_10734,N_8791,N_9149);
and U10735 (N_10735,N_9449,N_9086);
and U10736 (N_10736,N_9003,N_9592);
nand U10737 (N_10737,N_9402,N_9023);
nor U10738 (N_10738,N_9290,N_9201);
xnor U10739 (N_10739,N_8921,N_9307);
xor U10740 (N_10740,N_8598,N_9410);
or U10741 (N_10741,N_8789,N_9149);
nor U10742 (N_10742,N_9050,N_8402);
and U10743 (N_10743,N_9383,N_8870);
nand U10744 (N_10744,N_9070,N_9446);
nand U10745 (N_10745,N_9420,N_9035);
xor U10746 (N_10746,N_9457,N_8448);
nor U10747 (N_10747,N_8650,N_9293);
nor U10748 (N_10748,N_8831,N_8654);
nor U10749 (N_10749,N_8835,N_9098);
nand U10750 (N_10750,N_8952,N_8855);
and U10751 (N_10751,N_9011,N_8922);
nor U10752 (N_10752,N_8810,N_8864);
nand U10753 (N_10753,N_8521,N_9105);
xor U10754 (N_10754,N_9387,N_8836);
nand U10755 (N_10755,N_8564,N_9036);
nand U10756 (N_10756,N_8818,N_8637);
and U10757 (N_10757,N_8860,N_8689);
or U10758 (N_10758,N_8649,N_8978);
xnor U10759 (N_10759,N_9199,N_8914);
or U10760 (N_10760,N_9420,N_9235);
and U10761 (N_10761,N_9089,N_8855);
nand U10762 (N_10762,N_8449,N_8738);
and U10763 (N_10763,N_9144,N_9459);
or U10764 (N_10764,N_8772,N_8416);
or U10765 (N_10765,N_9329,N_9387);
and U10766 (N_10766,N_8728,N_9503);
nor U10767 (N_10767,N_9125,N_9195);
xor U10768 (N_10768,N_8716,N_8656);
nand U10769 (N_10769,N_8662,N_9096);
xnor U10770 (N_10770,N_8476,N_9053);
nand U10771 (N_10771,N_9172,N_9333);
and U10772 (N_10772,N_9316,N_9156);
or U10773 (N_10773,N_8705,N_8585);
and U10774 (N_10774,N_9456,N_9036);
or U10775 (N_10775,N_9182,N_8637);
and U10776 (N_10776,N_8405,N_9104);
or U10777 (N_10777,N_8786,N_8848);
or U10778 (N_10778,N_8902,N_9177);
nand U10779 (N_10779,N_9305,N_8433);
and U10780 (N_10780,N_8409,N_8448);
nor U10781 (N_10781,N_9028,N_8439);
and U10782 (N_10782,N_9521,N_8585);
or U10783 (N_10783,N_8942,N_9350);
xor U10784 (N_10784,N_8931,N_9480);
nor U10785 (N_10785,N_9323,N_9317);
or U10786 (N_10786,N_8921,N_9491);
nand U10787 (N_10787,N_8480,N_8845);
nand U10788 (N_10788,N_8654,N_9044);
nor U10789 (N_10789,N_8899,N_9518);
or U10790 (N_10790,N_9537,N_8561);
or U10791 (N_10791,N_9383,N_9465);
nand U10792 (N_10792,N_9419,N_8676);
or U10793 (N_10793,N_9140,N_9151);
nand U10794 (N_10794,N_9402,N_9369);
or U10795 (N_10795,N_9541,N_9248);
xnor U10796 (N_10796,N_9041,N_8417);
and U10797 (N_10797,N_8927,N_9165);
nor U10798 (N_10798,N_8501,N_8649);
or U10799 (N_10799,N_8909,N_8497);
and U10800 (N_10800,N_10451,N_10400);
xnor U10801 (N_10801,N_10606,N_10043);
nand U10802 (N_10802,N_10156,N_10212);
and U10803 (N_10803,N_9979,N_10372);
or U10804 (N_10804,N_10786,N_9742);
xor U10805 (N_10805,N_10251,N_10349);
xnor U10806 (N_10806,N_10151,N_9711);
xnor U10807 (N_10807,N_10505,N_10022);
nand U10808 (N_10808,N_10376,N_10727);
or U10809 (N_10809,N_10129,N_10631);
nand U10810 (N_10810,N_10615,N_9898);
nor U10811 (N_10811,N_10770,N_9886);
and U10812 (N_10812,N_10145,N_9967);
nor U10813 (N_10813,N_10160,N_10423);
xnor U10814 (N_10814,N_9725,N_9668);
xnor U10815 (N_10815,N_9770,N_10166);
nor U10816 (N_10816,N_10038,N_10000);
nand U10817 (N_10817,N_10256,N_10176);
nor U10818 (N_10818,N_10456,N_10626);
and U10819 (N_10819,N_10379,N_9970);
nor U10820 (N_10820,N_10206,N_10028);
or U10821 (N_10821,N_9690,N_9747);
or U10822 (N_10822,N_10403,N_10506);
or U10823 (N_10823,N_10331,N_10027);
and U10824 (N_10824,N_9663,N_10470);
and U10825 (N_10825,N_10224,N_10088);
or U10826 (N_10826,N_10309,N_10348);
and U10827 (N_10827,N_10278,N_9655);
and U10828 (N_10828,N_10593,N_9769);
and U10829 (N_10829,N_10313,N_10202);
nand U10830 (N_10830,N_10414,N_10655);
and U10831 (N_10831,N_10083,N_10014);
or U10832 (N_10832,N_10792,N_9635);
and U10833 (N_10833,N_10575,N_9790);
nor U10834 (N_10834,N_10262,N_10019);
nand U10835 (N_10835,N_10772,N_10102);
xnor U10836 (N_10836,N_9767,N_10387);
nor U10837 (N_10837,N_10696,N_9691);
or U10838 (N_10838,N_10679,N_10527);
nand U10839 (N_10839,N_10104,N_10069);
nor U10840 (N_10840,N_9906,N_10780);
nor U10841 (N_10841,N_9741,N_9986);
and U10842 (N_10842,N_9860,N_9638);
nand U10843 (N_10843,N_9706,N_10075);
and U10844 (N_10844,N_10633,N_10619);
xnor U10845 (N_10845,N_9908,N_10116);
or U10846 (N_10846,N_10107,N_9919);
or U10847 (N_10847,N_10471,N_9793);
nor U10848 (N_10848,N_10449,N_10360);
or U10849 (N_10849,N_10045,N_9708);
and U10850 (N_10850,N_10775,N_10308);
or U10851 (N_10851,N_9912,N_10258);
nor U10852 (N_10852,N_10316,N_9832);
or U10853 (N_10853,N_10194,N_9882);
nand U10854 (N_10854,N_10502,N_10443);
nor U10855 (N_10855,N_10171,N_10494);
or U10856 (N_10856,N_9870,N_10611);
xnor U10857 (N_10857,N_9651,N_9994);
and U10858 (N_10858,N_10179,N_9842);
and U10859 (N_10859,N_9649,N_9798);
xnor U10860 (N_10860,N_9892,N_10790);
and U10861 (N_10861,N_10073,N_10574);
and U10862 (N_10862,N_9686,N_9784);
xnor U10863 (N_10863,N_9625,N_9704);
or U10864 (N_10864,N_10568,N_10358);
or U10865 (N_10865,N_10534,N_10623);
or U10866 (N_10866,N_10667,N_9807);
and U10867 (N_10867,N_10498,N_9610);
xnor U10868 (N_10868,N_9838,N_10690);
xor U10869 (N_10869,N_9836,N_10023);
or U10870 (N_10870,N_10677,N_10473);
nor U10871 (N_10871,N_10647,N_9774);
xnor U10872 (N_10872,N_10742,N_9921);
nand U10873 (N_10873,N_10565,N_9978);
nor U10874 (N_10874,N_9626,N_10060);
nor U10875 (N_10875,N_10082,N_10612);
nand U10876 (N_10876,N_10672,N_10620);
nand U10877 (N_10877,N_9679,N_9710);
nor U10878 (N_10878,N_10148,N_10569);
nand U10879 (N_10879,N_10636,N_9909);
nand U10880 (N_10880,N_10207,N_9930);
nor U10881 (N_10881,N_9619,N_10217);
xnor U10882 (N_10882,N_9865,N_9781);
and U10883 (N_10883,N_10726,N_10366);
nor U10884 (N_10884,N_10136,N_10249);
or U10885 (N_10885,N_9731,N_10468);
or U10886 (N_10886,N_9857,N_10461);
or U10887 (N_10887,N_10455,N_10197);
or U10888 (N_10888,N_10791,N_9802);
nand U10889 (N_10889,N_10409,N_9702);
or U10890 (N_10890,N_10356,N_10120);
nand U10891 (N_10891,N_10297,N_10117);
xor U10892 (N_10892,N_9602,N_10531);
xnor U10893 (N_10893,N_9695,N_10472);
and U10894 (N_10894,N_9825,N_10537);
xor U10895 (N_10895,N_9714,N_10111);
xnor U10896 (N_10896,N_10335,N_10322);
or U10897 (N_10897,N_9947,N_9751);
nor U10898 (N_10898,N_10553,N_10225);
nand U10899 (N_10899,N_10610,N_10517);
or U10900 (N_10900,N_10720,N_9612);
and U10901 (N_10901,N_9843,N_10106);
nand U10902 (N_10902,N_9678,N_10552);
nand U10903 (N_10903,N_9687,N_10776);
xor U10904 (N_10904,N_9667,N_10657);
xor U10905 (N_10905,N_10706,N_9716);
xor U10906 (N_10906,N_9883,N_10412);
or U10907 (N_10907,N_10152,N_10269);
nand U10908 (N_10908,N_10535,N_10204);
or U10909 (N_10909,N_10296,N_10398);
nor U10910 (N_10910,N_10345,N_10496);
xor U10911 (N_10911,N_9778,N_9913);
nor U10912 (N_10912,N_10645,N_10718);
and U10913 (N_10913,N_10291,N_10497);
xnor U10914 (N_10914,N_10523,N_9922);
and U10915 (N_10915,N_10510,N_9964);
or U10916 (N_10916,N_10613,N_10085);
xor U10917 (N_10917,N_10637,N_10728);
or U10918 (N_10918,N_10103,N_10514);
nand U10919 (N_10919,N_10715,N_10500);
or U10920 (N_10920,N_10268,N_10259);
or U10921 (N_10921,N_10192,N_9760);
nor U10922 (N_10922,N_10036,N_10374);
and U10923 (N_10923,N_10722,N_9962);
and U10924 (N_10924,N_9879,N_9833);
or U10925 (N_10925,N_10702,N_10422);
nand U10926 (N_10926,N_9673,N_9664);
xnor U10927 (N_10927,N_10522,N_10601);
nor U10928 (N_10928,N_10438,N_9939);
or U10929 (N_10929,N_10035,N_10650);
or U10930 (N_10930,N_9739,N_10385);
xor U10931 (N_10931,N_9713,N_10177);
xor U10932 (N_10932,N_9800,N_10064);
or U10933 (N_10933,N_10245,N_9980);
nor U10934 (N_10934,N_10501,N_10688);
or U10935 (N_10935,N_10420,N_10150);
or U10936 (N_10936,N_9701,N_10214);
and U10937 (N_10937,N_10630,N_10652);
and U10938 (N_10938,N_10664,N_9779);
nor U10939 (N_10939,N_10643,N_10757);
nor U10940 (N_10940,N_10089,N_9944);
or U10941 (N_10941,N_9855,N_10208);
or U10942 (N_10942,N_10573,N_10238);
or U10943 (N_10943,N_10131,N_10754);
nor U10944 (N_10944,N_9943,N_10286);
and U10945 (N_10945,N_10598,N_10274);
or U10946 (N_10946,N_10109,N_9840);
or U10947 (N_10947,N_9814,N_10597);
nor U10948 (N_10948,N_10012,N_10283);
nor U10949 (N_10949,N_10067,N_10220);
or U10950 (N_10950,N_10056,N_10428);
and U10951 (N_10951,N_10063,N_9995);
and U10952 (N_10952,N_9854,N_10042);
nand U10953 (N_10953,N_10602,N_10175);
or U10954 (N_10954,N_9904,N_10448);
nand U10955 (N_10955,N_10065,N_10796);
nand U10956 (N_10956,N_9791,N_9754);
and U10957 (N_10957,N_9940,N_10680);
nand U10958 (N_10958,N_10763,N_10210);
xor U10959 (N_10959,N_9957,N_10549);
xnor U10960 (N_10960,N_10756,N_10797);
nand U10961 (N_10961,N_10137,N_10660);
xnor U10962 (N_10962,N_9866,N_9808);
xor U10963 (N_10963,N_10343,N_9736);
nand U10964 (N_10964,N_10550,N_10266);
or U10965 (N_10965,N_10339,N_10072);
or U10966 (N_10966,N_10653,N_10371);
nor U10967 (N_10967,N_10777,N_10429);
xnor U10968 (N_10968,N_10578,N_10458);
nand U10969 (N_10969,N_9672,N_10714);
or U10970 (N_10970,N_10669,N_9993);
or U10971 (N_10971,N_10144,N_10512);
or U10972 (N_10972,N_10017,N_10189);
and U10973 (N_10973,N_9888,N_10235);
nand U10974 (N_10974,N_10748,N_10388);
and U10975 (N_10975,N_9786,N_10282);
nand U10976 (N_10976,N_10676,N_10566);
nor U10977 (N_10977,N_9956,N_9758);
or U10978 (N_10978,N_10233,N_9862);
xor U10979 (N_10979,N_10557,N_10033);
nand U10980 (N_10980,N_10561,N_10218);
nor U10981 (N_10981,N_10052,N_10609);
nand U10982 (N_10982,N_10798,N_10094);
nand U10983 (N_10983,N_9744,N_10627);
or U10984 (N_10984,N_10591,N_10029);
nand U10985 (N_10985,N_10105,N_10751);
xnor U10986 (N_10986,N_10415,N_10289);
or U10987 (N_10987,N_10319,N_10689);
nor U10988 (N_10988,N_10250,N_10034);
nand U10989 (N_10989,N_10684,N_10205);
nor U10990 (N_10990,N_10671,N_10717);
nor U10991 (N_10991,N_10521,N_9705);
nor U10992 (N_10992,N_10070,N_10305);
nand U10993 (N_10993,N_9991,N_10273);
and U10994 (N_10994,N_10767,N_10768);
or U10995 (N_10995,N_10323,N_9941);
and U10996 (N_10996,N_10548,N_10723);
nand U10997 (N_10997,N_9960,N_9897);
nand U10998 (N_10998,N_10749,N_9927);
and U10999 (N_10999,N_9765,N_9834);
and U11000 (N_11000,N_10162,N_10541);
nand U11001 (N_11001,N_9934,N_9617);
and U11002 (N_11002,N_9887,N_10277);
and U11003 (N_11003,N_10232,N_10426);
nor U11004 (N_11004,N_9762,N_10304);
and U11005 (N_11005,N_10559,N_9606);
nor U11006 (N_11006,N_9863,N_10115);
nand U11007 (N_11007,N_10168,N_10730);
nand U11008 (N_11008,N_10050,N_10504);
nor U11009 (N_11009,N_10338,N_10607);
xor U11010 (N_11010,N_10396,N_10747);
and U11011 (N_11011,N_9605,N_10419);
nor U11012 (N_11012,N_9864,N_10011);
xor U11013 (N_11013,N_9818,N_10312);
or U11014 (N_11014,N_10554,N_9675);
nand U11015 (N_11015,N_10465,N_10632);
nor U11016 (N_11016,N_9928,N_9645);
nand U11017 (N_11017,N_10352,N_9682);
nor U11018 (N_11018,N_9620,N_9963);
xor U11019 (N_11019,N_10668,N_10333);
or U11020 (N_11020,N_10433,N_10087);
nor U11021 (N_11021,N_10294,N_10183);
or U11022 (N_11022,N_10203,N_9837);
nor U11023 (N_11023,N_10153,N_10579);
and U11024 (N_11024,N_10674,N_10533);
nor U11025 (N_11025,N_9873,N_9746);
xnor U11026 (N_11026,N_10406,N_10707);
xnor U11027 (N_11027,N_10519,N_10434);
xnor U11028 (N_11028,N_9847,N_10694);
or U11029 (N_11029,N_10764,N_9763);
xnor U11030 (N_11030,N_10622,N_10252);
and U11031 (N_11031,N_9910,N_10539);
or U11032 (N_11032,N_9955,N_9796);
xnor U11033 (N_11033,N_10771,N_10367);
nor U11034 (N_11034,N_9801,N_10698);
nor U11035 (N_11035,N_10134,N_9607);
nand U11036 (N_11036,N_10380,N_9875);
nor U11037 (N_11037,N_10234,N_9604);
xor U11038 (N_11038,N_10062,N_9665);
and U11039 (N_11039,N_10731,N_10783);
and U11040 (N_11040,N_10595,N_10544);
and U11041 (N_11041,N_10507,N_10200);
and U11042 (N_11042,N_10560,N_10529);
or U11043 (N_11043,N_9728,N_10229);
nor U11044 (N_11044,N_9715,N_10743);
xnor U11045 (N_11045,N_10354,N_10340);
and U11046 (N_11046,N_10157,N_10253);
and U11047 (N_11047,N_10442,N_9819);
xnor U11048 (N_11048,N_10002,N_9700);
xnor U11049 (N_11049,N_9601,N_10353);
and U11050 (N_11050,N_9637,N_10037);
and U11051 (N_11051,N_9899,N_10311);
or U11052 (N_11052,N_9968,N_10586);
nand U11053 (N_11053,N_10191,N_10344);
nand U11054 (N_11054,N_9724,N_9789);
and U11055 (N_11055,N_10605,N_10450);
and U11056 (N_11056,N_10737,N_10181);
or U11057 (N_11057,N_10418,N_10518);
or U11058 (N_11058,N_10264,N_10556);
or U11059 (N_11059,N_9684,N_10068);
nor U11060 (N_11060,N_10765,N_9926);
or U11061 (N_11061,N_10121,N_10469);
and U11062 (N_11062,N_10310,N_10365);
nand U11063 (N_11063,N_10161,N_10086);
xor U11064 (N_11064,N_10174,N_10048);
and U11065 (N_11065,N_10108,N_9821);
xnor U11066 (N_11066,N_10729,N_10397);
and U11067 (N_11067,N_9987,N_10099);
xor U11068 (N_11068,N_9976,N_10020);
nand U11069 (N_11069,N_9656,N_9661);
and U11070 (N_11070,N_10543,N_10716);
xnor U11071 (N_11071,N_9644,N_10713);
nand U11072 (N_11072,N_10604,N_10454);
xnor U11073 (N_11073,N_9810,N_10394);
and U11074 (N_11074,N_9831,N_10299);
xor U11075 (N_11075,N_9636,N_10039);
and U11076 (N_11076,N_10703,N_9916);
and U11077 (N_11077,N_10211,N_9952);
or U11078 (N_11078,N_10389,N_10571);
nor U11079 (N_11079,N_10375,N_10293);
and U11080 (N_11080,N_9654,N_10280);
or U11081 (N_11081,N_10329,N_10452);
and U11082 (N_11082,N_10378,N_9776);
or U11083 (N_11083,N_10377,N_9756);
or U11084 (N_11084,N_9698,N_10199);
xnor U11085 (N_11085,N_10363,N_9990);
nand U11086 (N_11086,N_10683,N_10746);
and U11087 (N_11087,N_10614,N_9680);
or U11088 (N_11088,N_9951,N_10782);
nor U11089 (N_11089,N_9642,N_9925);
or U11090 (N_11090,N_10328,N_10051);
and U11091 (N_11091,N_9975,N_10180);
or U11092 (N_11092,N_9827,N_9823);
and U11093 (N_11093,N_9653,N_9745);
nor U11094 (N_11094,N_10055,N_9845);
xor U11095 (N_11095,N_9856,N_9685);
or U11096 (N_11096,N_10444,N_10733);
nor U11097 (N_11097,N_10413,N_9905);
or U11098 (N_11098,N_9917,N_10324);
and U11099 (N_11099,N_10457,N_10386);
xnor U11100 (N_11100,N_10315,N_10432);
and U11101 (N_11101,N_10001,N_10074);
nor U11102 (N_11102,N_9616,N_9804);
or U11103 (N_11103,N_10477,N_9851);
or U11104 (N_11104,N_10638,N_9693);
nor U11105 (N_11105,N_10401,N_10018);
and U11106 (N_11106,N_10641,N_10480);
and U11107 (N_11107,N_10734,N_10079);
and U11108 (N_11108,N_10562,N_10185);
nand U11109 (N_11109,N_10583,N_10712);
or U11110 (N_11110,N_9813,N_10135);
xnor U11111 (N_11111,N_10320,N_10326);
nor U11112 (N_11112,N_10110,N_9861);
nand U11113 (N_11113,N_10678,N_9901);
xnor U11114 (N_11114,N_10705,N_10143);
nand U11115 (N_11115,N_10178,N_9902);
nand U11116 (N_11116,N_10755,N_10182);
or U11117 (N_11117,N_9624,N_9809);
nand U11118 (N_11118,N_9803,N_9752);
xor U11119 (N_11119,N_9877,N_9799);
nand U11120 (N_11120,N_9707,N_9871);
nand U11121 (N_11121,N_9671,N_10172);
or U11122 (N_11122,N_10327,N_10481);
and U11123 (N_11123,N_10475,N_10248);
xnor U11124 (N_11124,N_10084,N_10635);
nand U11125 (N_11125,N_9729,N_9629);
nor U11126 (N_11126,N_10355,N_10709);
and U11127 (N_11127,N_9923,N_10793);
or U11128 (N_11128,N_10681,N_9815);
and U11129 (N_11129,N_9611,N_9839);
or U11130 (N_11130,N_9829,N_9627);
nor U11131 (N_11131,N_10026,N_10100);
nor U11132 (N_11132,N_10260,N_9753);
nand U11133 (N_11133,N_9817,N_10546);
or U11134 (N_11134,N_10119,N_9938);
nand U11135 (N_11135,N_9792,N_9844);
or U11136 (N_11136,N_10302,N_10558);
or U11137 (N_11137,N_10138,N_10466);
or U11138 (N_11138,N_10009,N_10155);
nand U11139 (N_11139,N_10411,N_9785);
xor U11140 (N_11140,N_9722,N_10484);
xor U11141 (N_11141,N_10025,N_10330);
nor U11142 (N_11142,N_9949,N_10799);
nand U11143 (N_11143,N_10708,N_10659);
nand U11144 (N_11144,N_10752,N_9621);
nand U11145 (N_11145,N_10209,N_10113);
nor U11146 (N_11146,N_9717,N_10383);
xnor U11147 (N_11147,N_9757,N_10446);
xnor U11148 (N_11148,N_9982,N_10492);
nand U11149 (N_11149,N_10325,N_10795);
nand U11150 (N_11150,N_10342,N_9835);
nand U11151 (N_11151,N_10306,N_9755);
nand U11152 (N_11152,N_10096,N_10215);
or U11153 (N_11153,N_10053,N_10436);
nand U11154 (N_11154,N_10321,N_10163);
nand U11155 (N_11155,N_10361,N_9641);
nor U11156 (N_11156,N_10576,N_9683);
xnor U11157 (N_11157,N_9646,N_9894);
nor U11158 (N_11158,N_10254,N_10061);
nor U11159 (N_11159,N_10271,N_10402);
nand U11160 (N_11160,N_10687,N_9852);
and U11161 (N_11161,N_9609,N_9931);
nand U11162 (N_11162,N_10058,N_10230);
nor U11163 (N_11163,N_9999,N_10525);
nor U11164 (N_11164,N_9615,N_9853);
nand U11165 (N_11165,N_10059,N_9858);
and U11166 (N_11166,N_9735,N_9850);
nand U11167 (N_11167,N_9652,N_10692);
nand U11168 (N_11168,N_10164,N_10123);
and U11169 (N_11169,N_9761,N_10140);
xnor U11170 (N_11170,N_9948,N_10010);
xor U11171 (N_11171,N_10616,N_10785);
or U11172 (N_11172,N_10077,N_10098);
nor U11173 (N_11173,N_10464,N_10307);
nand U11174 (N_11174,N_10594,N_9658);
nor U11175 (N_11175,N_10758,N_10488);
or U11176 (N_11176,N_9650,N_9737);
or U11177 (N_11177,N_10127,N_10447);
nand U11178 (N_11178,N_10257,N_9872);
nor U11179 (N_11179,N_9712,N_10124);
and U11180 (N_11180,N_10314,N_10629);
or U11181 (N_11181,N_10691,N_9937);
xor U11182 (N_11182,N_10139,N_10459);
xor U11183 (N_11183,N_10003,N_10617);
xnor U11184 (N_11184,N_9777,N_10625);
nor U11185 (N_11185,N_10540,N_10370);
xnor U11186 (N_11186,N_10132,N_9694);
and U11187 (N_11187,N_10445,N_10287);
nor U11188 (N_11188,N_10133,N_9846);
nand U11189 (N_11189,N_9660,N_9797);
nor U11190 (N_11190,N_9895,N_10031);
or U11191 (N_11191,N_9726,N_10112);
or U11192 (N_11192,N_10649,N_10046);
nand U11193 (N_11193,N_9748,N_9878);
nand U11194 (N_11194,N_9911,N_10193);
or U11195 (N_11195,N_10318,N_10440);
nand U11196 (N_11196,N_10357,N_10169);
nor U11197 (N_11197,N_10198,N_9891);
and U11198 (N_11198,N_10350,N_10285);
nor U11199 (N_11199,N_9824,N_10013);
xor U11200 (N_11200,N_10049,N_10362);
nor U11201 (N_11201,N_9738,N_9775);
and U11202 (N_11202,N_9942,N_9953);
and U11203 (N_11203,N_9689,N_10592);
xor U11204 (N_11204,N_10281,N_10373);
nor U11205 (N_11205,N_10463,N_10016);
and U11206 (N_11206,N_10508,N_10582);
and U11207 (N_11207,N_10580,N_10644);
nor U11208 (N_11208,N_9772,N_10196);
and U11209 (N_11209,N_10509,N_10779);
xor U11210 (N_11210,N_10485,N_10794);
xnor U11211 (N_11211,N_9945,N_10317);
or U11212 (N_11212,N_10769,N_9732);
or U11213 (N_11213,N_10435,N_10301);
or U11214 (N_11214,N_10491,N_10292);
xnor U11215 (N_11215,N_10704,N_10670);
or U11216 (N_11216,N_9918,N_9730);
nor U11217 (N_11217,N_10228,N_9740);
xor U11218 (N_11218,N_10515,N_10697);
nor U11219 (N_11219,N_9764,N_10146);
xor U11220 (N_11220,N_10599,N_10516);
nor U11221 (N_11221,N_10261,N_9958);
nand U11222 (N_11222,N_10246,N_10467);
xor U11223 (N_11223,N_10588,N_9816);
and U11224 (N_11224,N_10745,N_9889);
nand U11225 (N_11225,N_9885,N_9634);
and U11226 (N_11226,N_10405,N_10195);
or U11227 (N_11227,N_10721,N_9628);
nand U11228 (N_11228,N_10167,N_9692);
nor U11229 (N_11229,N_10624,N_10490);
nand U11230 (N_11230,N_10787,N_10369);
xor U11231 (N_11231,N_9669,N_10476);
xnor U11232 (N_11232,N_9972,N_10462);
nand U11233 (N_11233,N_9743,N_9600);
nand U11234 (N_11234,N_9670,N_10532);
and U11235 (N_11235,N_9639,N_10524);
and U11236 (N_11236,N_10015,N_10760);
and U11237 (N_11237,N_9924,N_10404);
nand U11238 (N_11238,N_9721,N_10122);
xnor U11239 (N_11239,N_9632,N_9795);
or U11240 (N_11240,N_10416,N_10091);
and U11241 (N_11241,N_9859,N_10701);
and U11242 (N_11242,N_10024,N_9826);
xnor U11243 (N_11243,N_10732,N_10487);
nor U11244 (N_11244,N_10040,N_10242);
or U11245 (N_11245,N_10154,N_10646);
or U11246 (N_11246,N_9618,N_10538);
nor U11247 (N_11247,N_10572,N_10589);
nand U11248 (N_11248,N_10341,N_10226);
and U11249 (N_11249,N_10675,N_10288);
or U11250 (N_11250,N_9984,N_10431);
and U11251 (N_11251,N_10766,N_10608);
nor U11252 (N_11252,N_9734,N_10421);
nor U11253 (N_11253,N_10482,N_10596);
nand U11254 (N_11254,N_10545,N_9720);
and U11255 (N_11255,N_10577,N_10621);
and U11256 (N_11256,N_10030,N_9966);
nor U11257 (N_11257,N_10382,N_10738);
nor U11258 (N_11258,N_10739,N_10336);
xnor U11259 (N_11259,N_10044,N_9983);
nor U11260 (N_11260,N_10513,N_9974);
xor U11261 (N_11261,N_10662,N_10407);
nand U11262 (N_11262,N_10563,N_10231);
and U11263 (N_11263,N_10551,N_10744);
or U11264 (N_11264,N_10054,N_10227);
and U11265 (N_11265,N_10300,N_10095);
and U11266 (N_11266,N_9985,N_10710);
or U11267 (N_11267,N_10784,N_9959);
xnor U11268 (N_11268,N_10555,N_10618);
or U11269 (N_11269,N_10392,N_10359);
xnor U11270 (N_11270,N_9718,N_10590);
nand U11271 (N_11271,N_10526,N_10585);
nor U11272 (N_11272,N_9805,N_10699);
nand U11273 (N_11273,N_9914,N_9603);
nor U11274 (N_11274,N_9699,N_10789);
or U11275 (N_11275,N_10346,N_10390);
and U11276 (N_11276,N_10460,N_9780);
nand U11277 (N_11277,N_10520,N_10237);
nor U11278 (N_11278,N_9933,N_10188);
nand U11279 (N_11279,N_9662,N_9971);
nand U11280 (N_11280,N_10158,N_9841);
and U11281 (N_11281,N_10778,N_10528);
nand U11282 (N_11282,N_10685,N_10337);
and U11283 (N_11283,N_10651,N_10236);
nor U11284 (N_11284,N_9647,N_9659);
nor U11285 (N_11285,N_9688,N_10640);
or U11286 (N_11286,N_10725,N_10489);
xor U11287 (N_11287,N_9768,N_10190);
nand U11288 (N_11288,N_10682,N_10673);
xnor U11289 (N_11289,N_10334,N_10788);
nor U11290 (N_11290,N_10265,N_10474);
nand U11291 (N_11291,N_9881,N_9900);
nor U11292 (N_11292,N_10666,N_10695);
nor U11293 (N_11293,N_10781,N_10187);
and U11294 (N_11294,N_10542,N_9954);
or U11295 (N_11295,N_9766,N_9727);
xnor U11296 (N_11296,N_10093,N_10092);
nor U11297 (N_11297,N_10628,N_9812);
nand U11298 (N_11298,N_10005,N_9946);
and U11299 (N_11299,N_10128,N_9703);
and U11300 (N_11300,N_10658,N_9915);
nor U11301 (N_11301,N_10686,N_10564);
and U11302 (N_11302,N_10700,N_10536);
or U11303 (N_11303,N_10483,N_9903);
nor U11304 (N_11304,N_10284,N_9643);
nand U11305 (N_11305,N_10453,N_10439);
nor U11306 (N_11306,N_10759,N_9640);
nor U11307 (N_11307,N_10665,N_9630);
xnor U11308 (N_11308,N_10584,N_10735);
nand U11309 (N_11309,N_10384,N_10008);
nor U11310 (N_11310,N_9896,N_10057);
and U11311 (N_11311,N_10239,N_10241);
xor U11312 (N_11312,N_9992,N_10639);
and U11313 (N_11313,N_10170,N_9830);
and U11314 (N_11314,N_9920,N_9709);
and U11315 (N_11315,N_10441,N_10078);
and U11316 (N_11316,N_10654,N_9935);
xnor U11317 (N_11317,N_10149,N_10219);
and U11318 (N_11318,N_9783,N_9677);
xnor U11319 (N_11319,N_10486,N_9648);
nor U11320 (N_11320,N_10276,N_10351);
nand U11321 (N_11321,N_9907,N_9773);
or U11322 (N_11322,N_10750,N_9788);
or U11323 (N_11323,N_10774,N_10711);
xor U11324 (N_11324,N_10007,N_9977);
and U11325 (N_11325,N_9750,N_9965);
xor U11326 (N_11326,N_10101,N_9880);
and U11327 (N_11327,N_10503,N_10216);
or U11328 (N_11328,N_10080,N_9719);
nand U11329 (N_11329,N_10368,N_10047);
and U11330 (N_11330,N_10567,N_9828);
nand U11331 (N_11331,N_10761,N_10221);
nand U11332 (N_11332,N_9973,N_10303);
nand U11333 (N_11333,N_10587,N_9890);
and U11334 (N_11334,N_9771,N_10222);
xor U11335 (N_11335,N_9876,N_10570);
nor U11336 (N_11336,N_10332,N_9988);
and U11337 (N_11337,N_10391,N_10656);
xnor U11338 (N_11338,N_10648,N_9998);
nand U11339 (N_11339,N_10243,N_10399);
and U11340 (N_11340,N_10499,N_9961);
nor U11341 (N_11341,N_10661,N_10066);
and U11342 (N_11342,N_9848,N_9723);
nand U11343 (N_11343,N_10244,N_10634);
xnor U11344 (N_11344,N_9623,N_9806);
nor U11345 (N_11345,N_10410,N_10142);
or U11346 (N_11346,N_9614,N_10395);
nor U11347 (N_11347,N_10381,N_9884);
nor U11348 (N_11348,N_10240,N_10408);
or U11349 (N_11349,N_10663,N_9697);
xnor U11350 (N_11350,N_9666,N_10511);
nand U11351 (N_11351,N_10126,N_10493);
or U11352 (N_11352,N_9929,N_10118);
and U11353 (N_11353,N_9674,N_9782);
nor U11354 (N_11354,N_10530,N_10773);
or U11355 (N_11355,N_9932,N_10279);
and U11356 (N_11356,N_10427,N_10425);
xor U11357 (N_11357,N_10247,N_10417);
or U11358 (N_11358,N_10724,N_9811);
and U11359 (N_11359,N_10741,N_9997);
nor U11360 (N_11360,N_10295,N_10437);
xnor U11361 (N_11361,N_9794,N_10213);
and U11362 (N_11362,N_10021,N_9893);
or U11363 (N_11363,N_10125,N_9874);
xor U11364 (N_11364,N_10642,N_9759);
xnor U11365 (N_11365,N_10081,N_9696);
nand U11366 (N_11366,N_10159,N_10600);
and U11367 (N_11367,N_10130,N_9869);
or U11368 (N_11368,N_9613,N_10097);
nand U11369 (N_11369,N_10547,N_10275);
nor U11370 (N_11370,N_10201,N_9681);
or U11371 (N_11371,N_10165,N_9633);
nor U11372 (N_11372,N_9820,N_10478);
or U11373 (N_11373,N_10581,N_10290);
and U11374 (N_11374,N_10267,N_10347);
and U11375 (N_11375,N_9989,N_9936);
xor U11376 (N_11376,N_10298,N_10147);
nand U11377 (N_11377,N_10364,N_9822);
xor U11378 (N_11378,N_10186,N_10603);
nand U11379 (N_11379,N_10263,N_10424);
nor U11380 (N_11380,N_10430,N_10762);
xor U11381 (N_11381,N_9622,N_10495);
nand U11382 (N_11382,N_10740,N_10032);
nor U11383 (N_11383,N_10255,N_10090);
xor U11384 (N_11384,N_10004,N_9631);
xor U11385 (N_11385,N_10719,N_10076);
nor U11386 (N_11386,N_10114,N_10006);
xnor U11387 (N_11387,N_10223,N_10736);
xor U11388 (N_11388,N_10272,N_10393);
or U11389 (N_11389,N_10270,N_10479);
or U11390 (N_11390,N_10184,N_9981);
and U11391 (N_11391,N_9787,N_10141);
nand U11392 (N_11392,N_9950,N_10071);
or U11393 (N_11393,N_9749,N_10041);
or U11394 (N_11394,N_9868,N_9867);
nand U11395 (N_11395,N_9849,N_10753);
nor U11396 (N_11396,N_10173,N_9676);
and U11397 (N_11397,N_9996,N_9733);
xor U11398 (N_11398,N_9608,N_10693);
nand U11399 (N_11399,N_9969,N_9657);
xor U11400 (N_11400,N_9837,N_10784);
xnor U11401 (N_11401,N_10316,N_10663);
xor U11402 (N_11402,N_10490,N_10391);
or U11403 (N_11403,N_9707,N_9814);
or U11404 (N_11404,N_9616,N_10776);
and U11405 (N_11405,N_10558,N_10472);
nor U11406 (N_11406,N_10364,N_10200);
and U11407 (N_11407,N_10211,N_10575);
and U11408 (N_11408,N_9672,N_10189);
and U11409 (N_11409,N_10067,N_9917);
and U11410 (N_11410,N_9761,N_10221);
and U11411 (N_11411,N_9729,N_9656);
or U11412 (N_11412,N_10559,N_10570);
xor U11413 (N_11413,N_10755,N_9997);
and U11414 (N_11414,N_9996,N_10623);
nand U11415 (N_11415,N_10052,N_10056);
nor U11416 (N_11416,N_9940,N_10682);
nor U11417 (N_11417,N_9788,N_9853);
nand U11418 (N_11418,N_10370,N_9675);
and U11419 (N_11419,N_10134,N_9928);
nand U11420 (N_11420,N_10709,N_10505);
or U11421 (N_11421,N_10179,N_9945);
nor U11422 (N_11422,N_10361,N_10391);
nor U11423 (N_11423,N_9936,N_9877);
nor U11424 (N_11424,N_10174,N_10008);
nor U11425 (N_11425,N_10082,N_9689);
nor U11426 (N_11426,N_10122,N_9685);
and U11427 (N_11427,N_10040,N_9812);
nor U11428 (N_11428,N_10773,N_9637);
nor U11429 (N_11429,N_9727,N_9784);
and U11430 (N_11430,N_10238,N_9805);
or U11431 (N_11431,N_10766,N_10052);
xor U11432 (N_11432,N_9820,N_10400);
nor U11433 (N_11433,N_10551,N_9618);
xnor U11434 (N_11434,N_10128,N_10445);
xor U11435 (N_11435,N_10253,N_9775);
or U11436 (N_11436,N_9787,N_10213);
and U11437 (N_11437,N_10417,N_9690);
or U11438 (N_11438,N_10348,N_10287);
xor U11439 (N_11439,N_10243,N_10701);
nor U11440 (N_11440,N_10299,N_9902);
and U11441 (N_11441,N_9896,N_10445);
and U11442 (N_11442,N_10022,N_9773);
nor U11443 (N_11443,N_9636,N_10431);
xnor U11444 (N_11444,N_10474,N_10211);
xor U11445 (N_11445,N_10484,N_10302);
and U11446 (N_11446,N_10194,N_9912);
xnor U11447 (N_11447,N_10011,N_10128);
and U11448 (N_11448,N_10311,N_10643);
or U11449 (N_11449,N_9996,N_10048);
or U11450 (N_11450,N_10197,N_9990);
nand U11451 (N_11451,N_9691,N_10032);
or U11452 (N_11452,N_10793,N_10702);
nor U11453 (N_11453,N_10342,N_10492);
nand U11454 (N_11454,N_10061,N_10171);
nand U11455 (N_11455,N_9941,N_10222);
nor U11456 (N_11456,N_9671,N_9898);
and U11457 (N_11457,N_10262,N_10348);
and U11458 (N_11458,N_10662,N_10273);
or U11459 (N_11459,N_10483,N_9911);
or U11460 (N_11460,N_10058,N_10094);
nor U11461 (N_11461,N_9734,N_10416);
nor U11462 (N_11462,N_10793,N_10645);
and U11463 (N_11463,N_9622,N_10342);
nor U11464 (N_11464,N_10096,N_10075);
or U11465 (N_11465,N_10220,N_10477);
nor U11466 (N_11466,N_10317,N_10583);
nor U11467 (N_11467,N_9948,N_10385);
nand U11468 (N_11468,N_10100,N_10206);
or U11469 (N_11469,N_9793,N_10456);
nand U11470 (N_11470,N_10156,N_10052);
and U11471 (N_11471,N_10578,N_10412);
and U11472 (N_11472,N_10582,N_10403);
and U11473 (N_11473,N_10415,N_9726);
and U11474 (N_11474,N_9800,N_9653);
nand U11475 (N_11475,N_10627,N_9602);
nor U11476 (N_11476,N_10241,N_10729);
nor U11477 (N_11477,N_9937,N_10711);
xnor U11478 (N_11478,N_9955,N_10277);
xnor U11479 (N_11479,N_10247,N_10138);
xnor U11480 (N_11480,N_10410,N_9991);
xnor U11481 (N_11481,N_10686,N_10484);
xnor U11482 (N_11482,N_10269,N_10476);
or U11483 (N_11483,N_9802,N_10648);
and U11484 (N_11484,N_9677,N_10783);
nor U11485 (N_11485,N_10656,N_10367);
nand U11486 (N_11486,N_10311,N_10403);
nor U11487 (N_11487,N_10147,N_10296);
xor U11488 (N_11488,N_9617,N_9833);
xnor U11489 (N_11489,N_9994,N_10215);
nor U11490 (N_11490,N_10022,N_9748);
xor U11491 (N_11491,N_10600,N_9880);
and U11492 (N_11492,N_10692,N_10256);
and U11493 (N_11493,N_9913,N_10005);
xnor U11494 (N_11494,N_10159,N_10413);
nand U11495 (N_11495,N_10179,N_10104);
nor U11496 (N_11496,N_9679,N_10686);
nand U11497 (N_11497,N_10261,N_10134);
and U11498 (N_11498,N_10740,N_10679);
nor U11499 (N_11499,N_9726,N_10384);
nand U11500 (N_11500,N_9769,N_10514);
and U11501 (N_11501,N_10585,N_9635);
nor U11502 (N_11502,N_10767,N_10424);
xor U11503 (N_11503,N_10637,N_9672);
xnor U11504 (N_11504,N_10020,N_9948);
or U11505 (N_11505,N_9948,N_10634);
and U11506 (N_11506,N_9668,N_9731);
or U11507 (N_11507,N_9763,N_10276);
or U11508 (N_11508,N_9665,N_9776);
nand U11509 (N_11509,N_10292,N_10015);
nand U11510 (N_11510,N_10329,N_10543);
nor U11511 (N_11511,N_9707,N_9718);
or U11512 (N_11512,N_10265,N_10518);
xnor U11513 (N_11513,N_10246,N_9955);
and U11514 (N_11514,N_9754,N_10216);
nor U11515 (N_11515,N_10044,N_10255);
xor U11516 (N_11516,N_10421,N_10349);
or U11517 (N_11517,N_9782,N_9861);
nand U11518 (N_11518,N_9821,N_10299);
and U11519 (N_11519,N_10700,N_9667);
xnor U11520 (N_11520,N_10155,N_10287);
xor U11521 (N_11521,N_10032,N_10555);
or U11522 (N_11522,N_10687,N_9836);
xnor U11523 (N_11523,N_10278,N_10537);
xor U11524 (N_11524,N_10779,N_10277);
nor U11525 (N_11525,N_10793,N_9708);
xor U11526 (N_11526,N_9758,N_9975);
nand U11527 (N_11527,N_10418,N_10340);
xnor U11528 (N_11528,N_10262,N_9762);
or U11529 (N_11529,N_10781,N_9968);
and U11530 (N_11530,N_10216,N_10208);
xnor U11531 (N_11531,N_9610,N_9606);
nand U11532 (N_11532,N_9722,N_9788);
or U11533 (N_11533,N_10640,N_9898);
xnor U11534 (N_11534,N_9623,N_10331);
and U11535 (N_11535,N_9990,N_10547);
nand U11536 (N_11536,N_10363,N_9740);
nor U11537 (N_11537,N_10717,N_9699);
nor U11538 (N_11538,N_10580,N_10422);
or U11539 (N_11539,N_10344,N_9932);
nor U11540 (N_11540,N_10222,N_10105);
or U11541 (N_11541,N_10401,N_9673);
and U11542 (N_11542,N_10641,N_9922);
xor U11543 (N_11543,N_9824,N_10691);
or U11544 (N_11544,N_9616,N_9732);
and U11545 (N_11545,N_9898,N_10500);
nor U11546 (N_11546,N_9939,N_9983);
and U11547 (N_11547,N_10473,N_10398);
or U11548 (N_11548,N_10141,N_10626);
nor U11549 (N_11549,N_9944,N_10665);
nor U11550 (N_11550,N_10044,N_10637);
xnor U11551 (N_11551,N_10582,N_9944);
or U11552 (N_11552,N_10624,N_10349);
nor U11553 (N_11553,N_9627,N_10497);
nand U11554 (N_11554,N_10688,N_10145);
nand U11555 (N_11555,N_10019,N_9977);
nand U11556 (N_11556,N_10150,N_10709);
or U11557 (N_11557,N_10799,N_10617);
or U11558 (N_11558,N_10289,N_10738);
nand U11559 (N_11559,N_10561,N_10642);
nor U11560 (N_11560,N_9600,N_10391);
nand U11561 (N_11561,N_10088,N_10205);
or U11562 (N_11562,N_10150,N_9855);
nor U11563 (N_11563,N_9889,N_9615);
nor U11564 (N_11564,N_10651,N_10029);
or U11565 (N_11565,N_10225,N_10062);
nand U11566 (N_11566,N_10159,N_10429);
xnor U11567 (N_11567,N_10655,N_10118);
xnor U11568 (N_11568,N_9631,N_9908);
or U11569 (N_11569,N_10337,N_10015);
nor U11570 (N_11570,N_10110,N_9919);
nand U11571 (N_11571,N_10107,N_9988);
nand U11572 (N_11572,N_9821,N_10522);
nand U11573 (N_11573,N_10260,N_9765);
xnor U11574 (N_11574,N_10336,N_9824);
nor U11575 (N_11575,N_10084,N_10737);
nand U11576 (N_11576,N_10587,N_10172);
xor U11577 (N_11577,N_9604,N_10336);
nand U11578 (N_11578,N_10145,N_9718);
nor U11579 (N_11579,N_10493,N_9645);
or U11580 (N_11580,N_10656,N_10011);
and U11581 (N_11581,N_9637,N_9649);
or U11582 (N_11582,N_9686,N_10684);
and U11583 (N_11583,N_9870,N_10691);
nand U11584 (N_11584,N_10715,N_10304);
and U11585 (N_11585,N_9842,N_10214);
or U11586 (N_11586,N_10376,N_10509);
nor U11587 (N_11587,N_9624,N_9637);
and U11588 (N_11588,N_9610,N_9708);
xnor U11589 (N_11589,N_9972,N_10361);
and U11590 (N_11590,N_9658,N_10566);
xnor U11591 (N_11591,N_10315,N_10777);
or U11592 (N_11592,N_9871,N_9851);
nor U11593 (N_11593,N_10288,N_9683);
nor U11594 (N_11594,N_10445,N_10734);
nand U11595 (N_11595,N_10521,N_9754);
or U11596 (N_11596,N_9834,N_10358);
and U11597 (N_11597,N_10722,N_9913);
and U11598 (N_11598,N_10652,N_10027);
nand U11599 (N_11599,N_9722,N_10288);
xnor U11600 (N_11600,N_9604,N_9610);
or U11601 (N_11601,N_10184,N_9914);
nand U11602 (N_11602,N_9898,N_10034);
xor U11603 (N_11603,N_10581,N_9986);
nand U11604 (N_11604,N_10095,N_10528);
or U11605 (N_11605,N_9941,N_10430);
nor U11606 (N_11606,N_10276,N_9981);
or U11607 (N_11607,N_10325,N_10102);
nor U11608 (N_11608,N_9681,N_10390);
or U11609 (N_11609,N_9787,N_10627);
xnor U11610 (N_11610,N_9786,N_10444);
nand U11611 (N_11611,N_10566,N_9822);
nor U11612 (N_11612,N_10264,N_9845);
or U11613 (N_11613,N_10674,N_9796);
or U11614 (N_11614,N_10471,N_10078);
nand U11615 (N_11615,N_10571,N_10632);
nand U11616 (N_11616,N_10610,N_10394);
nor U11617 (N_11617,N_10694,N_10360);
or U11618 (N_11618,N_10616,N_9770);
and U11619 (N_11619,N_10016,N_10178);
nand U11620 (N_11620,N_10799,N_9885);
xnor U11621 (N_11621,N_10633,N_10548);
or U11622 (N_11622,N_9779,N_10573);
nand U11623 (N_11623,N_9687,N_9671);
and U11624 (N_11624,N_10468,N_9888);
xnor U11625 (N_11625,N_9608,N_9848);
nor U11626 (N_11626,N_10561,N_10338);
and U11627 (N_11627,N_9999,N_10129);
nor U11628 (N_11628,N_9681,N_9751);
xor U11629 (N_11629,N_10322,N_10268);
xor U11630 (N_11630,N_9789,N_10259);
nand U11631 (N_11631,N_10250,N_10472);
or U11632 (N_11632,N_10164,N_10731);
and U11633 (N_11633,N_9761,N_9864);
xnor U11634 (N_11634,N_10705,N_10423);
and U11635 (N_11635,N_10225,N_10183);
and U11636 (N_11636,N_10153,N_10411);
and U11637 (N_11637,N_9791,N_9973);
nor U11638 (N_11638,N_9667,N_9944);
nand U11639 (N_11639,N_10519,N_10498);
and U11640 (N_11640,N_10254,N_9859);
or U11641 (N_11641,N_10026,N_9789);
and U11642 (N_11642,N_9710,N_10203);
and U11643 (N_11643,N_9969,N_10692);
xor U11644 (N_11644,N_9659,N_9640);
and U11645 (N_11645,N_9829,N_10488);
or U11646 (N_11646,N_10205,N_10132);
or U11647 (N_11647,N_10480,N_9817);
xnor U11648 (N_11648,N_10326,N_10509);
or U11649 (N_11649,N_10799,N_10503);
nor U11650 (N_11650,N_9953,N_10343);
nor U11651 (N_11651,N_9853,N_9811);
nor U11652 (N_11652,N_10515,N_9706);
nand U11653 (N_11653,N_9699,N_9729);
and U11654 (N_11654,N_9989,N_9737);
nor U11655 (N_11655,N_10766,N_10219);
and U11656 (N_11656,N_9613,N_9607);
nor U11657 (N_11657,N_9962,N_10508);
xnor U11658 (N_11658,N_10349,N_9687);
and U11659 (N_11659,N_10686,N_10621);
nor U11660 (N_11660,N_10566,N_9947);
nor U11661 (N_11661,N_9636,N_10454);
nand U11662 (N_11662,N_9863,N_9716);
nor U11663 (N_11663,N_10558,N_10256);
nand U11664 (N_11664,N_9731,N_10283);
nand U11665 (N_11665,N_9800,N_9697);
nor U11666 (N_11666,N_10195,N_10706);
xnor U11667 (N_11667,N_10445,N_10631);
nand U11668 (N_11668,N_9869,N_10250);
and U11669 (N_11669,N_9667,N_10632);
nand U11670 (N_11670,N_9766,N_10099);
xor U11671 (N_11671,N_10306,N_9614);
xor U11672 (N_11672,N_10069,N_9612);
or U11673 (N_11673,N_10097,N_9674);
nor U11674 (N_11674,N_9729,N_10337);
or U11675 (N_11675,N_10455,N_10334);
xnor U11676 (N_11676,N_10650,N_10187);
nand U11677 (N_11677,N_10458,N_10376);
nor U11678 (N_11678,N_10780,N_9813);
or U11679 (N_11679,N_10555,N_10238);
xor U11680 (N_11680,N_10314,N_10298);
nand U11681 (N_11681,N_10635,N_10208);
nor U11682 (N_11682,N_10329,N_9619);
or U11683 (N_11683,N_10069,N_9626);
nor U11684 (N_11684,N_9672,N_10025);
and U11685 (N_11685,N_10294,N_10473);
xnor U11686 (N_11686,N_10278,N_10181);
or U11687 (N_11687,N_9945,N_9685);
or U11688 (N_11688,N_9875,N_10484);
xnor U11689 (N_11689,N_9792,N_10565);
or U11690 (N_11690,N_10293,N_10610);
nand U11691 (N_11691,N_9796,N_9689);
or U11692 (N_11692,N_10750,N_10788);
nand U11693 (N_11693,N_10745,N_10732);
and U11694 (N_11694,N_10225,N_10686);
xor U11695 (N_11695,N_10138,N_10372);
nor U11696 (N_11696,N_9749,N_10327);
nor U11697 (N_11697,N_10331,N_10180);
and U11698 (N_11698,N_9957,N_10394);
xor U11699 (N_11699,N_10695,N_9731);
nand U11700 (N_11700,N_10411,N_10679);
nand U11701 (N_11701,N_10715,N_10209);
nor U11702 (N_11702,N_10149,N_10174);
or U11703 (N_11703,N_9620,N_9623);
xor U11704 (N_11704,N_10503,N_10280);
nand U11705 (N_11705,N_10490,N_10758);
or U11706 (N_11706,N_10772,N_10224);
nor U11707 (N_11707,N_10798,N_10656);
nor U11708 (N_11708,N_10280,N_10356);
nand U11709 (N_11709,N_9816,N_9961);
xor U11710 (N_11710,N_10676,N_9864);
nor U11711 (N_11711,N_10166,N_10220);
nand U11712 (N_11712,N_10033,N_9849);
or U11713 (N_11713,N_10137,N_10648);
nor U11714 (N_11714,N_10699,N_10612);
or U11715 (N_11715,N_10339,N_10520);
or U11716 (N_11716,N_10104,N_10010);
and U11717 (N_11717,N_10602,N_10198);
or U11718 (N_11718,N_10447,N_9883);
nor U11719 (N_11719,N_10125,N_10040);
nand U11720 (N_11720,N_10029,N_10067);
and U11721 (N_11721,N_10623,N_10408);
and U11722 (N_11722,N_9947,N_9971);
and U11723 (N_11723,N_9990,N_10193);
and U11724 (N_11724,N_10376,N_9764);
xnor U11725 (N_11725,N_9726,N_10186);
nand U11726 (N_11726,N_10284,N_9938);
and U11727 (N_11727,N_9882,N_10707);
xor U11728 (N_11728,N_9749,N_10428);
and U11729 (N_11729,N_10300,N_10241);
nand U11730 (N_11730,N_10349,N_10333);
or U11731 (N_11731,N_10111,N_10766);
xor U11732 (N_11732,N_10253,N_10076);
or U11733 (N_11733,N_10143,N_10457);
or U11734 (N_11734,N_10609,N_9629);
nand U11735 (N_11735,N_10365,N_10545);
or U11736 (N_11736,N_10624,N_10688);
nor U11737 (N_11737,N_10752,N_10477);
xnor U11738 (N_11738,N_10578,N_10495);
or U11739 (N_11739,N_9803,N_10692);
or U11740 (N_11740,N_10081,N_10537);
or U11741 (N_11741,N_9746,N_10624);
or U11742 (N_11742,N_9886,N_10549);
nor U11743 (N_11743,N_9661,N_10789);
or U11744 (N_11744,N_10057,N_9730);
or U11745 (N_11745,N_10026,N_10536);
xor U11746 (N_11746,N_9626,N_10179);
nor U11747 (N_11747,N_9635,N_10101);
xnor U11748 (N_11748,N_10660,N_10705);
xnor U11749 (N_11749,N_10702,N_10788);
and U11750 (N_11750,N_10026,N_10373);
nand U11751 (N_11751,N_10020,N_10311);
or U11752 (N_11752,N_10219,N_10453);
nand U11753 (N_11753,N_10714,N_10513);
or U11754 (N_11754,N_10669,N_10277);
nand U11755 (N_11755,N_10119,N_10042);
nor U11756 (N_11756,N_9780,N_10041);
nor U11757 (N_11757,N_10712,N_9940);
and U11758 (N_11758,N_10775,N_10746);
nand U11759 (N_11759,N_10795,N_10775);
or U11760 (N_11760,N_9681,N_9625);
nand U11761 (N_11761,N_10385,N_10028);
nand U11762 (N_11762,N_10152,N_10287);
and U11763 (N_11763,N_9986,N_9735);
nor U11764 (N_11764,N_10625,N_10408);
nand U11765 (N_11765,N_10748,N_10527);
nand U11766 (N_11766,N_10560,N_10285);
or U11767 (N_11767,N_10772,N_10498);
xnor U11768 (N_11768,N_10575,N_9820);
xnor U11769 (N_11769,N_10599,N_10268);
or U11770 (N_11770,N_9827,N_9951);
nor U11771 (N_11771,N_9923,N_9750);
xnor U11772 (N_11772,N_10217,N_10681);
nor U11773 (N_11773,N_10719,N_10779);
nor U11774 (N_11774,N_10467,N_10699);
xnor U11775 (N_11775,N_10318,N_9711);
xor U11776 (N_11776,N_10406,N_10549);
nand U11777 (N_11777,N_10623,N_10658);
or U11778 (N_11778,N_9922,N_9865);
nor U11779 (N_11779,N_9651,N_10690);
nand U11780 (N_11780,N_9862,N_10424);
nor U11781 (N_11781,N_10150,N_10753);
xor U11782 (N_11782,N_10248,N_10703);
nand U11783 (N_11783,N_10690,N_10051);
and U11784 (N_11784,N_9908,N_10555);
nor U11785 (N_11785,N_10333,N_10119);
or U11786 (N_11786,N_10280,N_10553);
and U11787 (N_11787,N_10410,N_10684);
xnor U11788 (N_11788,N_10705,N_10639);
nand U11789 (N_11789,N_9806,N_10502);
and U11790 (N_11790,N_9693,N_9620);
xor U11791 (N_11791,N_9795,N_10203);
nand U11792 (N_11792,N_9802,N_9669);
xor U11793 (N_11793,N_10534,N_10575);
nor U11794 (N_11794,N_9628,N_9750);
and U11795 (N_11795,N_9805,N_9843);
nor U11796 (N_11796,N_9666,N_9600);
or U11797 (N_11797,N_10353,N_10680);
nor U11798 (N_11798,N_10134,N_10609);
or U11799 (N_11799,N_10323,N_10362);
or U11800 (N_11800,N_9766,N_10203);
and U11801 (N_11801,N_10133,N_10743);
nor U11802 (N_11802,N_10650,N_9647);
nor U11803 (N_11803,N_10256,N_10723);
xor U11804 (N_11804,N_10143,N_10034);
or U11805 (N_11805,N_10510,N_10492);
and U11806 (N_11806,N_9639,N_10709);
xnor U11807 (N_11807,N_10344,N_9636);
nand U11808 (N_11808,N_10150,N_9743);
nor U11809 (N_11809,N_10708,N_10036);
nor U11810 (N_11810,N_9668,N_10303);
nand U11811 (N_11811,N_9710,N_9985);
nor U11812 (N_11812,N_10255,N_10204);
nand U11813 (N_11813,N_10630,N_10014);
xor U11814 (N_11814,N_10604,N_10696);
xor U11815 (N_11815,N_9866,N_10632);
xor U11816 (N_11816,N_10670,N_10656);
nand U11817 (N_11817,N_10408,N_9895);
or U11818 (N_11818,N_10560,N_9918);
or U11819 (N_11819,N_9812,N_9934);
xor U11820 (N_11820,N_9853,N_10387);
and U11821 (N_11821,N_10125,N_10541);
xor U11822 (N_11822,N_9889,N_9755);
or U11823 (N_11823,N_10380,N_10027);
xnor U11824 (N_11824,N_9821,N_9758);
and U11825 (N_11825,N_9929,N_10433);
nand U11826 (N_11826,N_10168,N_10204);
nand U11827 (N_11827,N_10220,N_9962);
nand U11828 (N_11828,N_10583,N_9647);
nand U11829 (N_11829,N_10194,N_10690);
xnor U11830 (N_11830,N_9762,N_10447);
nand U11831 (N_11831,N_10255,N_9787);
xnor U11832 (N_11832,N_9903,N_9961);
xnor U11833 (N_11833,N_10097,N_10439);
xnor U11834 (N_11834,N_10712,N_9762);
nand U11835 (N_11835,N_9922,N_10355);
nand U11836 (N_11836,N_10759,N_10499);
nand U11837 (N_11837,N_10534,N_10598);
and U11838 (N_11838,N_9785,N_9970);
xor U11839 (N_11839,N_9793,N_10573);
nand U11840 (N_11840,N_10620,N_10422);
or U11841 (N_11841,N_10759,N_9839);
xor U11842 (N_11842,N_9818,N_9624);
nor U11843 (N_11843,N_9653,N_10727);
nand U11844 (N_11844,N_10016,N_10039);
nand U11845 (N_11845,N_9611,N_10484);
nor U11846 (N_11846,N_9917,N_10007);
nor U11847 (N_11847,N_9656,N_9986);
and U11848 (N_11848,N_10055,N_10232);
xor U11849 (N_11849,N_9978,N_9805);
nand U11850 (N_11850,N_10295,N_9936);
nand U11851 (N_11851,N_9677,N_10428);
and U11852 (N_11852,N_10156,N_10412);
and U11853 (N_11853,N_10291,N_10783);
or U11854 (N_11854,N_10262,N_10330);
nor U11855 (N_11855,N_10169,N_10747);
or U11856 (N_11856,N_9659,N_10468);
nor U11857 (N_11857,N_9879,N_10405);
nand U11858 (N_11858,N_9779,N_10420);
or U11859 (N_11859,N_9945,N_10717);
xor U11860 (N_11860,N_10521,N_10148);
nor U11861 (N_11861,N_10032,N_9749);
and U11862 (N_11862,N_10753,N_10124);
xnor U11863 (N_11863,N_9679,N_10675);
nand U11864 (N_11864,N_9788,N_10553);
xor U11865 (N_11865,N_9779,N_10584);
nor U11866 (N_11866,N_10260,N_10077);
nor U11867 (N_11867,N_10607,N_10081);
or U11868 (N_11868,N_9612,N_9771);
or U11869 (N_11869,N_10570,N_9983);
nor U11870 (N_11870,N_10271,N_9653);
xnor U11871 (N_11871,N_9876,N_9672);
nand U11872 (N_11872,N_10560,N_10144);
nor U11873 (N_11873,N_10408,N_9625);
xnor U11874 (N_11874,N_10258,N_9649);
xnor U11875 (N_11875,N_10135,N_9966);
or U11876 (N_11876,N_9657,N_10431);
nor U11877 (N_11877,N_10071,N_10653);
nand U11878 (N_11878,N_10450,N_10743);
and U11879 (N_11879,N_10714,N_10254);
nor U11880 (N_11880,N_9722,N_10179);
or U11881 (N_11881,N_9694,N_9897);
xnor U11882 (N_11882,N_9796,N_9612);
xnor U11883 (N_11883,N_10101,N_9636);
xnor U11884 (N_11884,N_10690,N_10313);
nor U11885 (N_11885,N_10305,N_10779);
and U11886 (N_11886,N_10683,N_10570);
nor U11887 (N_11887,N_9974,N_9744);
or U11888 (N_11888,N_10518,N_10545);
and U11889 (N_11889,N_10493,N_10204);
xnor U11890 (N_11890,N_10048,N_9861);
and U11891 (N_11891,N_10717,N_10252);
or U11892 (N_11892,N_10588,N_10694);
nor U11893 (N_11893,N_10450,N_9942);
nor U11894 (N_11894,N_9952,N_10539);
or U11895 (N_11895,N_10675,N_9939);
xnor U11896 (N_11896,N_10026,N_10464);
and U11897 (N_11897,N_9832,N_10115);
nand U11898 (N_11898,N_9956,N_10689);
xnor U11899 (N_11899,N_10688,N_9845);
and U11900 (N_11900,N_10492,N_10188);
and U11901 (N_11901,N_10762,N_9605);
or U11902 (N_11902,N_9621,N_10292);
nor U11903 (N_11903,N_10286,N_9657);
nand U11904 (N_11904,N_10160,N_10293);
xor U11905 (N_11905,N_9940,N_10355);
and U11906 (N_11906,N_9797,N_10074);
or U11907 (N_11907,N_10463,N_9699);
xnor U11908 (N_11908,N_10255,N_10607);
or U11909 (N_11909,N_10623,N_10336);
nand U11910 (N_11910,N_9639,N_10028);
nor U11911 (N_11911,N_9698,N_9970);
and U11912 (N_11912,N_10594,N_10431);
or U11913 (N_11913,N_10700,N_10466);
or U11914 (N_11914,N_10610,N_9650);
and U11915 (N_11915,N_9946,N_9942);
nand U11916 (N_11916,N_10762,N_10436);
nand U11917 (N_11917,N_9875,N_10035);
and U11918 (N_11918,N_10272,N_10190);
nand U11919 (N_11919,N_10742,N_9739);
and U11920 (N_11920,N_10752,N_10680);
nand U11921 (N_11921,N_9654,N_9667);
nand U11922 (N_11922,N_10026,N_10222);
and U11923 (N_11923,N_10102,N_10743);
or U11924 (N_11924,N_10248,N_10685);
and U11925 (N_11925,N_9862,N_10051);
and U11926 (N_11926,N_10402,N_10512);
nand U11927 (N_11927,N_9743,N_10250);
and U11928 (N_11928,N_10786,N_9829);
xnor U11929 (N_11929,N_10611,N_9750);
nor U11930 (N_11930,N_9694,N_10494);
or U11931 (N_11931,N_10604,N_10525);
and U11932 (N_11932,N_10297,N_10154);
xnor U11933 (N_11933,N_9887,N_9914);
and U11934 (N_11934,N_10437,N_10072);
nor U11935 (N_11935,N_9652,N_9672);
or U11936 (N_11936,N_9844,N_10712);
xor U11937 (N_11937,N_9754,N_10253);
xor U11938 (N_11938,N_9613,N_9639);
nand U11939 (N_11939,N_9866,N_10004);
and U11940 (N_11940,N_10260,N_9620);
or U11941 (N_11941,N_10440,N_10746);
nand U11942 (N_11942,N_10740,N_10680);
and U11943 (N_11943,N_9971,N_10018);
xor U11944 (N_11944,N_10122,N_9782);
and U11945 (N_11945,N_10293,N_10795);
nand U11946 (N_11946,N_10166,N_10736);
nor U11947 (N_11947,N_10484,N_10121);
nand U11948 (N_11948,N_10022,N_10537);
nand U11949 (N_11949,N_9954,N_9868);
and U11950 (N_11950,N_10454,N_10336);
and U11951 (N_11951,N_9648,N_10557);
nor U11952 (N_11952,N_10603,N_10086);
nand U11953 (N_11953,N_10400,N_10157);
and U11954 (N_11954,N_10576,N_10403);
nor U11955 (N_11955,N_10386,N_10642);
or U11956 (N_11956,N_10182,N_10640);
or U11957 (N_11957,N_9980,N_10288);
xor U11958 (N_11958,N_10697,N_9807);
nor U11959 (N_11959,N_10158,N_9773);
nor U11960 (N_11960,N_9741,N_9960);
or U11961 (N_11961,N_9821,N_10470);
nand U11962 (N_11962,N_10330,N_10782);
nor U11963 (N_11963,N_9675,N_9655);
xor U11964 (N_11964,N_10743,N_10608);
or U11965 (N_11965,N_10753,N_9951);
nor U11966 (N_11966,N_9722,N_10642);
or U11967 (N_11967,N_9912,N_10041);
or U11968 (N_11968,N_9760,N_10104);
nor U11969 (N_11969,N_10664,N_10266);
and U11970 (N_11970,N_9724,N_9908);
nor U11971 (N_11971,N_9909,N_10690);
nand U11972 (N_11972,N_10706,N_10583);
nor U11973 (N_11973,N_10343,N_9778);
or U11974 (N_11974,N_10395,N_10485);
and U11975 (N_11975,N_10100,N_9839);
and U11976 (N_11976,N_10389,N_10167);
nor U11977 (N_11977,N_10759,N_10658);
nand U11978 (N_11978,N_9948,N_9756);
xor U11979 (N_11979,N_10656,N_10143);
xor U11980 (N_11980,N_9739,N_10514);
nor U11981 (N_11981,N_10093,N_9932);
nor U11982 (N_11982,N_10765,N_10440);
xor U11983 (N_11983,N_9897,N_10023);
nand U11984 (N_11984,N_10405,N_10410);
or U11985 (N_11985,N_9900,N_10449);
nor U11986 (N_11986,N_9630,N_10581);
xnor U11987 (N_11987,N_10188,N_9619);
nand U11988 (N_11988,N_9774,N_9899);
or U11989 (N_11989,N_10429,N_9699);
nor U11990 (N_11990,N_9879,N_10724);
nor U11991 (N_11991,N_10000,N_10133);
and U11992 (N_11992,N_9841,N_10061);
xnor U11993 (N_11993,N_10562,N_10283);
nand U11994 (N_11994,N_10631,N_10037);
xnor U11995 (N_11995,N_9923,N_9911);
xnor U11996 (N_11996,N_9652,N_10357);
xor U11997 (N_11997,N_9865,N_10550);
and U11998 (N_11998,N_9898,N_9912);
or U11999 (N_11999,N_9641,N_9761);
nand U12000 (N_12000,N_11287,N_11554);
nor U12001 (N_12001,N_11926,N_11636);
or U12002 (N_12002,N_11604,N_11424);
nand U12003 (N_12003,N_11182,N_10969);
nor U12004 (N_12004,N_11267,N_10882);
nand U12005 (N_12005,N_11565,N_10970);
nor U12006 (N_12006,N_11129,N_11143);
or U12007 (N_12007,N_10808,N_11240);
or U12008 (N_12008,N_11208,N_11200);
xnor U12009 (N_12009,N_11079,N_10949);
and U12010 (N_12010,N_11893,N_11647);
nand U12011 (N_12011,N_11715,N_11545);
nor U12012 (N_12012,N_10896,N_11736);
nor U12013 (N_12013,N_11788,N_11070);
and U12014 (N_12014,N_11854,N_11247);
or U12015 (N_12015,N_11502,N_10888);
nor U12016 (N_12016,N_11995,N_11531);
nor U12017 (N_12017,N_11379,N_10804);
nor U12018 (N_12018,N_10943,N_11999);
nand U12019 (N_12019,N_11603,N_10884);
nor U12020 (N_12020,N_11054,N_11351);
nand U12021 (N_12021,N_11362,N_10957);
or U12022 (N_12022,N_11924,N_11477);
xor U12023 (N_12023,N_10862,N_10831);
xnor U12024 (N_12024,N_11506,N_11546);
or U12025 (N_12025,N_11642,N_11364);
or U12026 (N_12026,N_11931,N_11654);
nor U12027 (N_12027,N_10860,N_11163);
or U12028 (N_12028,N_11375,N_11831);
nor U12029 (N_12029,N_11946,N_10815);
xnor U12030 (N_12030,N_11433,N_11898);
nor U12031 (N_12031,N_11227,N_11073);
nor U12032 (N_12032,N_11314,N_11086);
nand U12033 (N_12033,N_11809,N_11431);
and U12034 (N_12034,N_11156,N_11657);
nor U12035 (N_12035,N_11274,N_11094);
nor U12036 (N_12036,N_11199,N_11869);
nor U12037 (N_12037,N_11519,N_11465);
and U12038 (N_12038,N_11386,N_10809);
and U12039 (N_12039,N_11009,N_11127);
nor U12040 (N_12040,N_11252,N_11515);
or U12041 (N_12041,N_11707,N_10936);
xnor U12042 (N_12042,N_11178,N_11296);
or U12043 (N_12043,N_10989,N_10976);
and U12044 (N_12044,N_10941,N_11663);
or U12045 (N_12045,N_11101,N_11555);
nor U12046 (N_12046,N_11705,N_11119);
or U12047 (N_12047,N_11138,N_11718);
or U12048 (N_12048,N_11695,N_11660);
nand U12049 (N_12049,N_11840,N_10820);
xnor U12050 (N_12050,N_11338,N_11332);
or U12051 (N_12051,N_11185,N_10986);
and U12052 (N_12052,N_10806,N_11441);
nand U12053 (N_12053,N_11579,N_11400);
nand U12054 (N_12054,N_11949,N_11453);
and U12055 (N_12055,N_11655,N_11624);
or U12056 (N_12056,N_11213,N_11838);
xnor U12057 (N_12057,N_11359,N_11861);
and U12058 (N_12058,N_11874,N_10801);
nor U12059 (N_12059,N_11971,N_11260);
xor U12060 (N_12060,N_11008,N_11571);
and U12061 (N_12061,N_11166,N_11035);
and U12062 (N_12062,N_11915,N_11281);
and U12063 (N_12063,N_11569,N_11610);
nand U12064 (N_12064,N_11959,N_11968);
nor U12065 (N_12065,N_11573,N_11850);
or U12066 (N_12066,N_11225,N_11394);
and U12067 (N_12067,N_11142,N_11455);
nand U12068 (N_12068,N_10994,N_10818);
xor U12069 (N_12069,N_11595,N_11914);
and U12070 (N_12070,N_11014,N_11120);
or U12071 (N_12071,N_11594,N_11757);
and U12072 (N_12072,N_11784,N_11262);
xor U12073 (N_12073,N_11940,N_11769);
and U12074 (N_12074,N_11964,N_11206);
nand U12075 (N_12075,N_11969,N_11589);
nor U12076 (N_12076,N_11732,N_11984);
nor U12077 (N_12077,N_11050,N_11948);
or U12078 (N_12078,N_11556,N_10861);
or U12079 (N_12079,N_11886,N_11268);
nor U12080 (N_12080,N_10915,N_11202);
and U12081 (N_12081,N_10865,N_11652);
xor U12082 (N_12082,N_11983,N_11640);
and U12083 (N_12083,N_11493,N_11828);
xor U12084 (N_12084,N_11765,N_11942);
or U12085 (N_12085,N_11567,N_11446);
nand U12086 (N_12086,N_11273,N_11108);
and U12087 (N_12087,N_11030,N_11685);
or U12088 (N_12088,N_11029,N_10902);
nor U12089 (N_12089,N_11986,N_11771);
nor U12090 (N_12090,N_11813,N_11904);
nand U12091 (N_12091,N_11929,N_10887);
nor U12092 (N_12092,N_11476,N_11945);
nand U12093 (N_12093,N_10958,N_11780);
nor U12094 (N_12094,N_11069,N_11532);
and U12095 (N_12095,N_11412,N_11102);
and U12096 (N_12096,N_11113,N_11656);
and U12097 (N_12097,N_11071,N_11128);
and U12098 (N_12098,N_11012,N_10833);
xnor U12099 (N_12099,N_10883,N_11851);
nand U12100 (N_12100,N_10853,N_11234);
and U12101 (N_12101,N_11615,N_10866);
xnor U12102 (N_12102,N_11888,N_11658);
and U12103 (N_12103,N_11155,N_10964);
nor U12104 (N_12104,N_11430,N_10810);
nand U12105 (N_12105,N_11885,N_10800);
nand U12106 (N_12106,N_11348,N_11489);
or U12107 (N_12107,N_11005,N_11833);
nand U12108 (N_12108,N_11614,N_10863);
nor U12109 (N_12109,N_11037,N_11717);
nand U12110 (N_12110,N_10946,N_11272);
and U12111 (N_12111,N_10814,N_11315);
xnor U12112 (N_12112,N_11100,N_11848);
xor U12113 (N_12113,N_11303,N_11318);
xor U12114 (N_12114,N_11048,N_11921);
nand U12115 (N_12115,N_11378,N_11807);
nor U12116 (N_12116,N_11798,N_11755);
and U12117 (N_12117,N_10891,N_11503);
xnor U12118 (N_12118,N_11853,N_11752);
nor U12119 (N_12119,N_11474,N_11162);
nor U12120 (N_12120,N_10857,N_10873);
xnor U12121 (N_12121,N_11242,N_10913);
xnor U12122 (N_12122,N_11870,N_11148);
nand U12123 (N_12123,N_10910,N_11421);
nor U12124 (N_12124,N_11814,N_11253);
and U12125 (N_12125,N_11751,N_11425);
or U12126 (N_12126,N_11360,N_10961);
and U12127 (N_12127,N_11961,N_11856);
and U12128 (N_12128,N_11323,N_11947);
or U12129 (N_12129,N_11533,N_11244);
or U12130 (N_12130,N_10911,N_11326);
nor U12131 (N_12131,N_11965,N_11080);
and U12132 (N_12132,N_11583,N_10907);
and U12133 (N_12133,N_11409,N_11927);
or U12134 (N_12134,N_11011,N_11665);
or U12135 (N_12135,N_11417,N_11028);
or U12136 (N_12136,N_11980,N_10988);
nand U12137 (N_12137,N_10802,N_11460);
and U12138 (N_12138,N_11026,N_11577);
xnor U12139 (N_12139,N_11301,N_10929);
nand U12140 (N_12140,N_11836,N_11509);
or U12141 (N_12141,N_10968,N_11955);
nor U12142 (N_12142,N_11538,N_10942);
or U12143 (N_12143,N_11782,N_11334);
or U12144 (N_12144,N_11313,N_11564);
nand U12145 (N_12145,N_11159,N_11495);
nor U12146 (N_12146,N_11612,N_11398);
nor U12147 (N_12147,N_10992,N_11889);
or U12148 (N_12148,N_11787,N_11250);
or U12149 (N_12149,N_11406,N_11371);
nor U12150 (N_12150,N_11237,N_10850);
xnor U12151 (N_12151,N_11543,N_11633);
or U12152 (N_12152,N_11077,N_11261);
and U12153 (N_12153,N_11778,N_11843);
or U12154 (N_12154,N_11471,N_10991);
nand U12155 (N_12155,N_11345,N_11270);
nand U12156 (N_12156,N_11684,N_11541);
nor U12157 (N_12157,N_11084,N_11115);
nand U12158 (N_12158,N_11203,N_11370);
nor U12159 (N_12159,N_11295,N_11672);
nor U12160 (N_12160,N_11741,N_11795);
nor U12161 (N_12161,N_11230,N_11057);
or U12162 (N_12162,N_11962,N_11910);
or U12163 (N_12163,N_11083,N_11329);
xor U12164 (N_12164,N_11561,N_11064);
xnor U12165 (N_12165,N_11095,N_10962);
or U12166 (N_12166,N_11863,N_11264);
xnor U12167 (N_12167,N_11469,N_11696);
nor U12168 (N_12168,N_11661,N_11047);
and U12169 (N_12169,N_11172,N_11111);
or U12170 (N_12170,N_11878,N_11606);
nor U12171 (N_12171,N_11664,N_10940);
or U12172 (N_12172,N_11330,N_11623);
xnor U12173 (N_12173,N_11808,N_10901);
or U12174 (N_12174,N_11093,N_11675);
xor U12175 (N_12175,N_11410,N_10864);
or U12176 (N_12176,N_11740,N_11586);
or U12177 (N_12177,N_10931,N_11671);
xnor U12178 (N_12178,N_11783,N_11207);
nand U12179 (N_12179,N_10978,N_11320);
nand U12180 (N_12180,N_11494,N_11620);
and U12181 (N_12181,N_10847,N_11444);
or U12182 (N_12182,N_10885,N_11676);
or U12183 (N_12183,N_11377,N_11149);
nor U12184 (N_12184,N_11716,N_11279);
or U12185 (N_12185,N_11639,N_11897);
nand U12186 (N_12186,N_11161,N_11144);
nand U12187 (N_12187,N_11286,N_11456);
nand U12188 (N_12188,N_11505,N_10995);
nand U12189 (N_12189,N_11951,N_11758);
nand U12190 (N_12190,N_11141,N_11151);
and U12191 (N_12191,N_11063,N_10980);
nand U12192 (N_12192,N_11974,N_11682);
nor U12193 (N_12193,N_10892,N_11060);
or U12194 (N_12194,N_10956,N_11068);
xor U12195 (N_12195,N_11059,N_11714);
nand U12196 (N_12196,N_11523,N_11087);
nand U12197 (N_12197,N_10816,N_11475);
nor U12198 (N_12198,N_11316,N_11906);
and U12199 (N_12199,N_10990,N_11801);
nor U12200 (N_12200,N_11125,N_11212);
xor U12201 (N_12201,N_11017,N_10881);
nand U12202 (N_12202,N_11490,N_11540);
and U12203 (N_12203,N_11634,N_11764);
nor U12204 (N_12204,N_11343,N_10997);
nand U12205 (N_12205,N_11447,N_10965);
xnor U12206 (N_12206,N_11641,N_11649);
or U12207 (N_12207,N_11601,N_11756);
xor U12208 (N_12208,N_11350,N_11452);
or U12209 (N_12209,N_10824,N_11294);
nand U12210 (N_12210,N_11407,N_11473);
nor U12211 (N_12211,N_11165,N_11582);
or U12212 (N_12212,N_11650,N_11750);
nor U12213 (N_12213,N_11592,N_11600);
nand U12214 (N_12214,N_11291,N_11401);
and U12215 (N_12215,N_11006,N_11157);
and U12216 (N_12216,N_11775,N_11283);
nand U12217 (N_12217,N_11428,N_11958);
xnor U12218 (N_12218,N_11399,N_11145);
nand U12219 (N_12219,N_11524,N_11786);
xnor U12220 (N_12220,N_11039,N_10813);
and U12221 (N_12221,N_11498,N_11858);
and U12222 (N_12222,N_11023,N_11591);
xor U12223 (N_12223,N_11632,N_11164);
and U12224 (N_12224,N_11271,N_11597);
xor U12225 (N_12225,N_11404,N_11966);
and U12226 (N_12226,N_11891,N_11817);
xnor U12227 (N_12227,N_11557,N_11305);
or U12228 (N_12228,N_11275,N_11464);
and U12229 (N_12229,N_11415,N_11923);
or U12230 (N_12230,N_11449,N_11133);
nor U12231 (N_12231,N_10846,N_10872);
xor U12232 (N_12232,N_11857,N_11669);
nand U12233 (N_12233,N_11859,N_10985);
and U12234 (N_12234,N_11539,N_10858);
nor U12235 (N_12235,N_11179,N_11900);
or U12236 (N_12236,N_11815,N_11566);
and U12237 (N_12237,N_11822,N_11180);
and U12238 (N_12238,N_10827,N_11304);
nor U12239 (N_12239,N_11729,N_11903);
or U12240 (N_12240,N_11440,N_11219);
and U12241 (N_12241,N_11251,N_11698);
or U12242 (N_12242,N_11562,N_11395);
xnor U12243 (N_12243,N_11584,N_11146);
nand U12244 (N_12244,N_11462,N_11062);
nand U12245 (N_12245,N_10944,N_10803);
nor U12246 (N_12246,N_11492,N_10889);
and U12247 (N_12247,N_11816,N_10947);
or U12248 (N_12248,N_10854,N_11486);
nor U12249 (N_12249,N_10939,N_11277);
and U12250 (N_12250,N_11307,N_11110);
nand U12251 (N_12251,N_11046,N_11920);
or U12252 (N_12252,N_11956,N_11733);
or U12253 (N_12253,N_11667,N_11290);
xor U12254 (N_12254,N_11434,N_11380);
and U12255 (N_12255,N_11558,N_11979);
and U12256 (N_12256,N_11336,N_11036);
nor U12257 (N_12257,N_11061,N_11837);
xor U12258 (N_12258,N_11723,N_10904);
nor U12259 (N_12259,N_11276,N_11402);
nand U12260 (N_12260,N_11154,N_11526);
nor U12261 (N_12261,N_11987,N_11683);
nor U12262 (N_12262,N_11293,N_11957);
or U12263 (N_12263,N_11645,N_11680);
or U12264 (N_12264,N_11628,N_11880);
nand U12265 (N_12265,N_11075,N_10925);
nor U12266 (N_12266,N_11703,N_11373);
or U12267 (N_12267,N_11528,N_10819);
nand U12268 (N_12268,N_11681,N_10906);
nor U12269 (N_12269,N_11529,N_11516);
nand U12270 (N_12270,N_11547,N_11468);
nand U12271 (N_12271,N_11311,N_11875);
and U12272 (N_12272,N_11845,N_11693);
or U12273 (N_12273,N_11692,N_10935);
or U12274 (N_12274,N_11231,N_11483);
and U12275 (N_12275,N_11298,N_11259);
nor U12276 (N_12276,N_10830,N_11883);
nand U12277 (N_12277,N_11881,N_11832);
xnor U12278 (N_12278,N_11712,N_11704);
or U12279 (N_12279,N_10973,N_11779);
nor U12280 (N_12280,N_11198,N_10953);
and U12281 (N_12281,N_11835,N_11147);
or U12282 (N_12282,N_11970,N_11701);
nor U12283 (N_12283,N_11744,N_11626);
and U12284 (N_12284,N_10945,N_11099);
nor U12285 (N_12285,N_10950,N_10982);
and U12286 (N_12286,N_10894,N_11024);
nand U12287 (N_12287,N_11013,N_11422);
nand U12288 (N_12288,N_10979,N_11461);
or U12289 (N_12289,N_10897,N_11092);
nand U12290 (N_12290,N_11170,N_11222);
and U12291 (N_12291,N_11353,N_11321);
nor U12292 (N_12292,N_11004,N_11580);
and U12293 (N_12293,N_11194,N_11297);
or U12294 (N_12294,N_10930,N_11943);
and U12295 (N_12295,N_11022,N_11001);
nand U12296 (N_12296,N_11896,N_11363);
nor U12297 (N_12297,N_11977,N_11003);
and U12298 (N_12298,N_11762,N_11629);
and U12299 (N_12299,N_11153,N_11892);
and U12300 (N_12300,N_11190,N_11387);
xor U12301 (N_12301,N_10981,N_11518);
xor U12302 (N_12302,N_11439,N_11674);
and U12303 (N_12303,N_11867,N_10952);
or U12304 (N_12304,N_11559,N_10852);
nand U12305 (N_12305,N_11085,N_11748);
nor U12306 (N_12306,N_11209,N_11432);
and U12307 (N_12307,N_11357,N_11568);
nor U12308 (N_12308,N_11221,N_11605);
xor U12309 (N_12309,N_11123,N_11916);
xnor U12310 (N_12310,N_11458,N_11791);
nor U12311 (N_12311,N_11443,N_10845);
nand U12312 (N_12312,N_11160,N_11934);
or U12313 (N_12313,N_11511,N_11072);
nand U12314 (N_12314,N_11188,N_11922);
nand U12315 (N_12315,N_11106,N_11513);
xor U12316 (N_12316,N_11590,N_10832);
nor U12317 (N_12317,N_11299,N_11542);
or U12318 (N_12318,N_11873,N_11834);
nor U12319 (N_12319,N_11719,N_10916);
and U12320 (N_12320,N_11382,N_10890);
or U12321 (N_12321,N_11917,N_10983);
nand U12322 (N_12322,N_10849,N_11708);
nand U12323 (N_12323,N_11510,N_11792);
xnor U12324 (N_12324,N_10807,N_11361);
nand U12325 (N_12325,N_11369,N_11255);
xnor U12326 (N_12326,N_11622,N_11997);
nand U12327 (N_12327,N_11021,N_11497);
xnor U12328 (N_12328,N_11333,N_11939);
nand U12329 (N_12329,N_11312,N_11451);
or U12330 (N_12330,N_11019,N_11191);
xnor U12331 (N_12331,N_11445,N_11668);
xor U12332 (N_12332,N_11913,N_11105);
xnor U12333 (N_12333,N_11824,N_10919);
xnor U12334 (N_12334,N_10895,N_10839);
or U12335 (N_12335,N_11694,N_11820);
nand U12336 (N_12336,N_11045,N_11197);
nand U12337 (N_12337,N_11285,N_11168);
xor U12338 (N_12338,N_11082,N_11027);
nor U12339 (N_12339,N_11195,N_11617);
nor U12340 (N_12340,N_11224,N_11936);
xor U12341 (N_12341,N_11536,N_11551);
nor U12342 (N_12342,N_11288,N_11482);
or U12343 (N_12343,N_11181,N_11572);
or U12344 (N_12344,N_11484,N_10874);
or U12345 (N_12345,N_11709,N_11284);
nor U12346 (N_12346,N_10921,N_11549);
nor U12347 (N_12347,N_11319,N_10927);
and U12348 (N_12348,N_11644,N_11521);
or U12349 (N_12349,N_11385,N_11501);
nand U12350 (N_12350,N_11204,N_10926);
nor U12351 (N_12351,N_11081,N_11653);
nand U12352 (N_12352,N_10868,N_11630);
and U12353 (N_12353,N_11871,N_11340);
and U12354 (N_12354,N_11390,N_11745);
nor U12355 (N_12355,N_11659,N_11799);
nor U12356 (N_12356,N_11183,N_11932);
nand U12357 (N_12357,N_11470,N_11265);
or U12358 (N_12358,N_11175,N_11699);
xor U12359 (N_12359,N_11941,N_11043);
nor U12360 (N_12360,N_10977,N_10867);
and U12361 (N_12361,N_11408,N_10836);
or U12362 (N_12362,N_10844,N_10840);
nand U12363 (N_12363,N_10893,N_11872);
xor U12364 (N_12364,N_10875,N_11908);
and U12365 (N_12365,N_11918,N_11103);
nor U12366 (N_12366,N_11339,N_10811);
xnor U12367 (N_12367,N_11308,N_11376);
and U12368 (N_12368,N_11058,N_11429);
xor U12369 (N_12369,N_11789,N_11418);
nor U12370 (N_12370,N_11651,N_10922);
xnor U12371 (N_12371,N_11673,N_11890);
xor U12372 (N_12372,N_11727,N_11548);
nor U12373 (N_12373,N_11877,N_11570);
xor U12374 (N_12374,N_11938,N_11776);
nand U12375 (N_12375,N_11720,N_11534);
nand U12376 (N_12376,N_11739,N_11608);
xor U12377 (N_12377,N_11352,N_11040);
and U12378 (N_12378,N_11420,N_11670);
xor U12379 (N_12379,N_11220,N_11090);
and U12380 (N_12380,N_11587,N_11767);
nand U12381 (N_12381,N_11342,N_11356);
xnor U12382 (N_12382,N_11067,N_11504);
xnor U12383 (N_12383,N_11618,N_11459);
xnor U12384 (N_12384,N_11937,N_10967);
xnor U12385 (N_12385,N_10954,N_11882);
nor U12386 (N_12386,N_11613,N_11576);
nand U12387 (N_12387,N_11619,N_11132);
and U12388 (N_12388,N_11855,N_11812);
or U12389 (N_12389,N_11097,N_11860);
or U12390 (N_12390,N_11876,N_11435);
or U12391 (N_12391,N_11347,N_11517);
or U12392 (N_12392,N_11602,N_10848);
xor U12393 (N_12393,N_11950,N_11137);
or U12394 (N_12394,N_10999,N_10878);
or U12395 (N_12395,N_11074,N_11124);
nor U12396 (N_12396,N_11849,N_11829);
or U12397 (N_12397,N_11588,N_11368);
and U12398 (N_12398,N_11463,N_11392);
and U12399 (N_12399,N_11734,N_11724);
nand U12400 (N_12400,N_11830,N_11514);
nand U12401 (N_12401,N_11550,N_11044);
nor U12402 (N_12402,N_11131,N_11053);
xnor U12403 (N_12403,N_11211,N_11864);
and U12404 (N_12404,N_11989,N_11768);
xnor U12405 (N_12405,N_11819,N_11902);
or U12406 (N_12406,N_10821,N_11803);
or U12407 (N_12407,N_11678,N_11215);
xor U12408 (N_12408,N_10898,N_11972);
nand U12409 (N_12409,N_11354,N_10928);
nand U12410 (N_12410,N_11089,N_11585);
xor U12411 (N_12411,N_11530,N_11763);
or U12412 (N_12412,N_11827,N_11616);
or U12413 (N_12413,N_11679,N_11388);
and U12414 (N_12414,N_11282,N_11793);
xnor U12415 (N_12415,N_11990,N_11800);
nand U12416 (N_12416,N_11335,N_11396);
nor U12417 (N_12417,N_11846,N_11328);
and U12418 (N_12418,N_11366,N_11662);
xor U12419 (N_12419,N_11121,N_11358);
nand U12420 (N_12420,N_10880,N_11527);
and U12421 (N_12421,N_10903,N_11467);
nor U12422 (N_12422,N_11437,N_11677);
nor U12423 (N_12423,N_11785,N_11991);
nor U12424 (N_12424,N_11811,N_11263);
nand U12425 (N_12425,N_11866,N_11055);
xnor U12426 (N_12426,N_11933,N_10870);
and U12427 (N_12427,N_11894,N_10886);
or U12428 (N_12428,N_11372,N_11735);
nand U12429 (N_12429,N_11091,N_10963);
nor U12430 (N_12430,N_11895,N_10823);
nor U12431 (N_12431,N_11772,N_11689);
or U12432 (N_12432,N_11416,N_11967);
and U12433 (N_12433,N_10920,N_10938);
and U12434 (N_12434,N_10899,N_11810);
nand U12435 (N_12435,N_11925,N_11512);
xor U12436 (N_12436,N_11574,N_11217);
or U12437 (N_12437,N_11448,N_11169);
or U12438 (N_12438,N_11427,N_10908);
nand U12439 (N_12439,N_11487,N_11839);
nand U12440 (N_12440,N_11245,N_11690);
nand U12441 (N_12441,N_11847,N_11563);
nor U12442 (N_12442,N_11051,N_11201);
nand U12443 (N_12443,N_10923,N_11706);
or U12444 (N_12444,N_10876,N_11246);
xor U12445 (N_12445,N_11508,N_11114);
nor U12446 (N_12446,N_11140,N_11173);
and U12447 (N_12447,N_11746,N_11257);
or U12448 (N_12448,N_10805,N_11552);
and U12449 (N_12449,N_11031,N_10812);
or U12450 (N_12450,N_11996,N_11993);
xnor U12451 (N_12451,N_10972,N_11507);
nor U12452 (N_12452,N_10842,N_11078);
and U12453 (N_12453,N_11553,N_11909);
and U12454 (N_12454,N_10837,N_11302);
xor U12455 (N_12455,N_11438,N_11258);
nor U12456 (N_12456,N_10822,N_11248);
xor U12457 (N_12457,N_11049,N_10828);
or U12458 (N_12458,N_11802,N_11522);
nor U12459 (N_12459,N_10914,N_11625);
nand U12460 (N_12460,N_11844,N_11702);
nand U12461 (N_12461,N_11988,N_11280);
nand U12462 (N_12462,N_11560,N_11825);
and U12463 (N_12463,N_11954,N_11158);
or U12464 (N_12464,N_11973,N_11722);
nor U12465 (N_12465,N_11749,N_11136);
xor U12466 (N_12466,N_11309,N_10835);
nor U12467 (N_12467,N_11032,N_11002);
nand U12468 (N_12468,N_11236,N_11112);
and U12469 (N_12469,N_11535,N_11887);
xor U12470 (N_12470,N_11804,N_11066);
nand U12471 (N_12471,N_11478,N_11713);
xor U12472 (N_12472,N_11365,N_11826);
nor U12473 (N_12473,N_11928,N_11341);
and U12474 (N_12474,N_11238,N_11994);
nor U12475 (N_12475,N_10843,N_11152);
or U12476 (N_12476,N_11963,N_11648);
and U12477 (N_12477,N_11426,N_11218);
or U12478 (N_12478,N_11052,N_11774);
nor U12479 (N_12479,N_11249,N_11982);
nand U12480 (N_12480,N_11331,N_11269);
nand U12481 (N_12481,N_11544,N_11731);
nand U12482 (N_12482,N_10909,N_11773);
xnor U12483 (N_12483,N_11174,N_11256);
and U12484 (N_12484,N_11189,N_11499);
nand U12485 (N_12485,N_11596,N_10984);
or U12486 (N_12486,N_11289,N_11737);
xnor U12487 (N_12487,N_11096,N_11985);
nor U12488 (N_12488,N_11056,N_11777);
nand U12489 (N_12489,N_10998,N_11761);
xor U12490 (N_12490,N_11635,N_11466);
and U12491 (N_12491,N_10932,N_11076);
or U12492 (N_12492,N_11135,N_10924);
nor U12493 (N_12493,N_11726,N_11821);
or U12494 (N_12494,N_11391,N_10851);
nand U12495 (N_12495,N_11038,N_11520);
or U12496 (N_12496,N_11930,N_11781);
or U12497 (N_12497,N_10912,N_11337);
nand U12498 (N_12498,N_11868,N_10951);
and U12499 (N_12499,N_10937,N_11759);
nand U12500 (N_12500,N_10971,N_11122);
nor U12501 (N_12501,N_11806,N_11754);
nor U12502 (N_12502,N_10905,N_11117);
nor U12503 (N_12503,N_10933,N_11907);
nand U12504 (N_12504,N_10877,N_11241);
xnor U12505 (N_12505,N_11646,N_10834);
and U12506 (N_12506,N_11397,N_11196);
and U12507 (N_12507,N_11638,N_10855);
and U12508 (N_12508,N_11593,N_11389);
nor U12509 (N_12509,N_11697,N_11126);
and U12510 (N_12510,N_11216,N_11953);
or U12511 (N_12511,N_11015,N_11794);
nor U12512 (N_12512,N_11381,N_11232);
nor U12513 (N_12513,N_11223,N_11393);
and U12514 (N_12514,N_11310,N_11065);
nor U12515 (N_12515,N_11384,N_11905);
xor U12516 (N_12516,N_11598,N_11728);
nor U12517 (N_12517,N_10948,N_11790);
nand U12518 (N_12518,N_11116,N_11346);
or U12519 (N_12519,N_10918,N_11007);
or U12520 (N_12520,N_11383,N_11919);
nand U12521 (N_12521,N_11355,N_11852);
nand U12522 (N_12522,N_11228,N_11643);
xnor U12523 (N_12523,N_11367,N_11186);
nand U12524 (N_12524,N_11177,N_11214);
nand U12525 (N_12525,N_10966,N_11118);
nor U12526 (N_12526,N_11975,N_11411);
nor U12527 (N_12527,N_11998,N_10829);
or U12528 (N_12528,N_11637,N_11952);
xor U12529 (N_12529,N_11730,N_10859);
nor U12530 (N_12530,N_11488,N_11344);
xnor U12531 (N_12531,N_11254,N_10960);
nand U12532 (N_12532,N_11317,N_11992);
nor U12533 (N_12533,N_11192,N_11235);
nor U12534 (N_12534,N_10959,N_10975);
or U12535 (N_12535,N_11578,N_11710);
and U12536 (N_12536,N_11300,N_11760);
xor U12537 (N_12537,N_11805,N_10825);
nand U12538 (N_12538,N_11187,N_11842);
or U12539 (N_12539,N_11450,N_11243);
xnor U12540 (N_12540,N_11020,N_11687);
or U12541 (N_12541,N_11481,N_11841);
xor U12542 (N_12542,N_10826,N_11327);
and U12543 (N_12543,N_10869,N_11098);
and U12544 (N_12544,N_11753,N_11325);
xor U12545 (N_12545,N_10917,N_11981);
xor U12546 (N_12546,N_11935,N_11107);
nand U12547 (N_12547,N_11322,N_11167);
and U12548 (N_12548,N_11688,N_10838);
and U12549 (N_12549,N_11374,N_11607);
nor U12550 (N_12550,N_11403,N_10856);
xor U12551 (N_12551,N_11631,N_11088);
nor U12552 (N_12552,N_11472,N_11413);
nand U12553 (N_12553,N_11205,N_10934);
and U12554 (N_12554,N_11442,N_11796);
nor U12555 (N_12555,N_11405,N_11738);
nand U12556 (N_12556,N_11770,N_11193);
and U12557 (N_12557,N_11109,N_11747);
nand U12558 (N_12558,N_11229,N_11278);
or U12559 (N_12559,N_10993,N_10974);
nand U12560 (N_12560,N_11130,N_11725);
or U12561 (N_12561,N_11865,N_11978);
nor U12562 (N_12562,N_11419,N_10900);
nor U12563 (N_12563,N_11899,N_11266);
xnor U12564 (N_12564,N_11944,N_11491);
nor U12565 (N_12565,N_11743,N_11233);
nor U12566 (N_12566,N_11797,N_11823);
nor U12567 (N_12567,N_11911,N_11912);
or U12568 (N_12568,N_11599,N_11818);
nand U12569 (N_12569,N_11150,N_11609);
nand U12570 (N_12570,N_11766,N_10987);
nor U12571 (N_12571,N_11666,N_11034);
nor U12572 (N_12572,N_11324,N_11349);
xor U12573 (N_12573,N_11306,N_11485);
nand U12574 (N_12574,N_11721,N_11479);
or U12575 (N_12575,N_11976,N_10879);
and U12576 (N_12576,N_11184,N_11879);
nand U12577 (N_12577,N_11104,N_11901);
nor U12578 (N_12578,N_11033,N_11691);
or U12579 (N_12579,N_11581,N_11010);
nor U12580 (N_12580,N_10871,N_11041);
nand U12581 (N_12581,N_11742,N_11000);
nand U12582 (N_12582,N_11018,N_11611);
nor U12583 (N_12583,N_11134,N_11627);
or U12584 (N_12584,N_11042,N_11960);
or U12585 (N_12585,N_11480,N_11292);
nand U12586 (N_12586,N_11537,N_11171);
nand U12587 (N_12587,N_11016,N_10996);
xnor U12588 (N_12588,N_11414,N_11621);
xnor U12589 (N_12589,N_11457,N_11239);
nand U12590 (N_12590,N_11496,N_10841);
and U12591 (N_12591,N_11700,N_11686);
nor U12592 (N_12592,N_11176,N_11436);
xor U12593 (N_12593,N_10955,N_11226);
xnor U12594 (N_12594,N_11454,N_10817);
or U12595 (N_12595,N_11884,N_11711);
nor U12596 (N_12596,N_11500,N_11025);
nand U12597 (N_12597,N_11139,N_11423);
nand U12598 (N_12598,N_11210,N_11525);
and U12599 (N_12599,N_11862,N_11575);
and U12600 (N_12600,N_11517,N_11437);
xnor U12601 (N_12601,N_11573,N_11877);
and U12602 (N_12602,N_11088,N_11047);
and U12603 (N_12603,N_11739,N_11272);
xor U12604 (N_12604,N_10923,N_11373);
nor U12605 (N_12605,N_11344,N_11064);
or U12606 (N_12606,N_11833,N_11337);
and U12607 (N_12607,N_10860,N_11585);
xor U12608 (N_12608,N_11811,N_11181);
xor U12609 (N_12609,N_11564,N_11521);
xnor U12610 (N_12610,N_11102,N_11482);
xor U12611 (N_12611,N_10931,N_11864);
nor U12612 (N_12612,N_11813,N_11261);
and U12613 (N_12613,N_11318,N_11704);
xor U12614 (N_12614,N_11937,N_10847);
or U12615 (N_12615,N_11984,N_11280);
xor U12616 (N_12616,N_10981,N_11303);
nand U12617 (N_12617,N_11051,N_11852);
nor U12618 (N_12618,N_11313,N_11290);
xor U12619 (N_12619,N_11282,N_11885);
and U12620 (N_12620,N_11345,N_11101);
or U12621 (N_12621,N_11139,N_11787);
xor U12622 (N_12622,N_11145,N_11308);
and U12623 (N_12623,N_11901,N_11841);
or U12624 (N_12624,N_11737,N_11718);
nor U12625 (N_12625,N_11405,N_11013);
and U12626 (N_12626,N_11845,N_10973);
or U12627 (N_12627,N_11338,N_11496);
nand U12628 (N_12628,N_11906,N_11522);
or U12629 (N_12629,N_10875,N_11253);
xor U12630 (N_12630,N_11783,N_11357);
nand U12631 (N_12631,N_10874,N_11291);
or U12632 (N_12632,N_10877,N_11048);
and U12633 (N_12633,N_11905,N_11816);
or U12634 (N_12634,N_10832,N_10965);
nor U12635 (N_12635,N_11394,N_11974);
nand U12636 (N_12636,N_11261,N_10896);
and U12637 (N_12637,N_10947,N_11042);
or U12638 (N_12638,N_11452,N_11208);
xor U12639 (N_12639,N_11535,N_11061);
or U12640 (N_12640,N_11338,N_11383);
xor U12641 (N_12641,N_10962,N_11385);
xor U12642 (N_12642,N_10870,N_11754);
xnor U12643 (N_12643,N_11053,N_10937);
or U12644 (N_12644,N_11452,N_11975);
nor U12645 (N_12645,N_11734,N_11404);
or U12646 (N_12646,N_10811,N_11225);
nand U12647 (N_12647,N_11435,N_11854);
nand U12648 (N_12648,N_11068,N_11151);
and U12649 (N_12649,N_11920,N_11533);
nor U12650 (N_12650,N_11679,N_11303);
nand U12651 (N_12651,N_11095,N_11013);
xnor U12652 (N_12652,N_11939,N_11459);
and U12653 (N_12653,N_11893,N_11616);
nor U12654 (N_12654,N_11325,N_11162);
or U12655 (N_12655,N_11233,N_10962);
or U12656 (N_12656,N_10853,N_11712);
or U12657 (N_12657,N_11720,N_11340);
and U12658 (N_12658,N_11124,N_11866);
nand U12659 (N_12659,N_11583,N_11490);
xnor U12660 (N_12660,N_11328,N_11473);
nand U12661 (N_12661,N_10946,N_11622);
and U12662 (N_12662,N_11281,N_11480);
xnor U12663 (N_12663,N_11384,N_11128);
and U12664 (N_12664,N_11091,N_11943);
nand U12665 (N_12665,N_11948,N_11602);
nor U12666 (N_12666,N_11669,N_10997);
nand U12667 (N_12667,N_11946,N_11003);
nand U12668 (N_12668,N_11154,N_11227);
or U12669 (N_12669,N_11917,N_11033);
nor U12670 (N_12670,N_11114,N_11236);
nor U12671 (N_12671,N_11347,N_11472);
or U12672 (N_12672,N_11396,N_11032);
nand U12673 (N_12673,N_10986,N_10821);
or U12674 (N_12674,N_11652,N_11631);
nand U12675 (N_12675,N_11390,N_11532);
or U12676 (N_12676,N_11501,N_11838);
nand U12677 (N_12677,N_11332,N_10814);
and U12678 (N_12678,N_11684,N_11523);
or U12679 (N_12679,N_10810,N_11721);
or U12680 (N_12680,N_11140,N_10936);
xor U12681 (N_12681,N_11392,N_11037);
nor U12682 (N_12682,N_11971,N_11753);
and U12683 (N_12683,N_10953,N_10993);
and U12684 (N_12684,N_11046,N_11935);
or U12685 (N_12685,N_11479,N_11104);
nor U12686 (N_12686,N_11398,N_11701);
nand U12687 (N_12687,N_11699,N_11666);
xnor U12688 (N_12688,N_11542,N_11573);
or U12689 (N_12689,N_11143,N_11763);
and U12690 (N_12690,N_10926,N_11910);
nor U12691 (N_12691,N_11136,N_11997);
and U12692 (N_12692,N_11978,N_11875);
and U12693 (N_12693,N_11005,N_11712);
nor U12694 (N_12694,N_11645,N_11412);
or U12695 (N_12695,N_11121,N_11596);
nor U12696 (N_12696,N_11007,N_11014);
nor U12697 (N_12697,N_11819,N_11168);
or U12698 (N_12698,N_11077,N_11369);
nand U12699 (N_12699,N_10960,N_11491);
and U12700 (N_12700,N_11380,N_11105);
nor U12701 (N_12701,N_11148,N_11541);
nor U12702 (N_12702,N_11568,N_10915);
or U12703 (N_12703,N_11965,N_10960);
nand U12704 (N_12704,N_11716,N_11258);
xor U12705 (N_12705,N_11643,N_11364);
and U12706 (N_12706,N_10956,N_10874);
nor U12707 (N_12707,N_11348,N_11506);
xnor U12708 (N_12708,N_11542,N_11109);
xor U12709 (N_12709,N_11048,N_11329);
nor U12710 (N_12710,N_11933,N_11878);
and U12711 (N_12711,N_11806,N_11677);
nor U12712 (N_12712,N_11550,N_11388);
xnor U12713 (N_12713,N_11446,N_11209);
and U12714 (N_12714,N_11956,N_11587);
nor U12715 (N_12715,N_11058,N_11611);
xnor U12716 (N_12716,N_11564,N_11188);
nor U12717 (N_12717,N_11919,N_11455);
nand U12718 (N_12718,N_10857,N_10865);
or U12719 (N_12719,N_11539,N_11721);
and U12720 (N_12720,N_11251,N_11846);
xnor U12721 (N_12721,N_11875,N_11680);
nand U12722 (N_12722,N_11359,N_11546);
or U12723 (N_12723,N_11322,N_11373);
nor U12724 (N_12724,N_11640,N_11183);
or U12725 (N_12725,N_11752,N_11171);
and U12726 (N_12726,N_11330,N_11724);
xor U12727 (N_12727,N_11415,N_11008);
or U12728 (N_12728,N_11281,N_11548);
and U12729 (N_12729,N_11726,N_11937);
or U12730 (N_12730,N_11065,N_10844);
nor U12731 (N_12731,N_11030,N_11065);
nor U12732 (N_12732,N_11099,N_11872);
nor U12733 (N_12733,N_10948,N_11600);
and U12734 (N_12734,N_10932,N_10810);
nand U12735 (N_12735,N_11637,N_11766);
and U12736 (N_12736,N_10853,N_11653);
and U12737 (N_12737,N_11199,N_11986);
nand U12738 (N_12738,N_11921,N_11078);
xnor U12739 (N_12739,N_10959,N_11160);
and U12740 (N_12740,N_11482,N_11030);
and U12741 (N_12741,N_11550,N_11403);
or U12742 (N_12742,N_11682,N_11259);
xor U12743 (N_12743,N_11955,N_11685);
and U12744 (N_12744,N_11656,N_11803);
nand U12745 (N_12745,N_11940,N_11999);
xnor U12746 (N_12746,N_11570,N_11783);
or U12747 (N_12747,N_11394,N_10975);
xnor U12748 (N_12748,N_11684,N_11937);
and U12749 (N_12749,N_11584,N_11525);
or U12750 (N_12750,N_11889,N_11420);
and U12751 (N_12751,N_11964,N_11735);
or U12752 (N_12752,N_11742,N_11309);
nor U12753 (N_12753,N_11911,N_11335);
or U12754 (N_12754,N_11952,N_11745);
and U12755 (N_12755,N_11095,N_11947);
xnor U12756 (N_12756,N_11448,N_11845);
and U12757 (N_12757,N_11012,N_11988);
nor U12758 (N_12758,N_11141,N_11937);
xor U12759 (N_12759,N_11880,N_11864);
nor U12760 (N_12760,N_11932,N_11207);
and U12761 (N_12761,N_11422,N_11792);
nand U12762 (N_12762,N_11837,N_11080);
and U12763 (N_12763,N_11828,N_11856);
xor U12764 (N_12764,N_11545,N_11112);
and U12765 (N_12765,N_11794,N_11121);
nor U12766 (N_12766,N_11544,N_11568);
nand U12767 (N_12767,N_10925,N_11872);
or U12768 (N_12768,N_11237,N_11322);
or U12769 (N_12769,N_11300,N_10879);
nand U12770 (N_12770,N_11108,N_11903);
and U12771 (N_12771,N_10947,N_11166);
or U12772 (N_12772,N_11426,N_10880);
and U12773 (N_12773,N_11162,N_11972);
and U12774 (N_12774,N_11946,N_11582);
nor U12775 (N_12775,N_11336,N_11437);
xor U12776 (N_12776,N_11434,N_11241);
nor U12777 (N_12777,N_11989,N_10946);
nand U12778 (N_12778,N_11154,N_10934);
and U12779 (N_12779,N_11078,N_11593);
nand U12780 (N_12780,N_11813,N_10837);
or U12781 (N_12781,N_11225,N_10886);
nand U12782 (N_12782,N_11912,N_11888);
and U12783 (N_12783,N_11862,N_11371);
nand U12784 (N_12784,N_11738,N_10875);
xnor U12785 (N_12785,N_11175,N_11650);
nor U12786 (N_12786,N_10883,N_11164);
nor U12787 (N_12787,N_11975,N_11266);
nand U12788 (N_12788,N_11440,N_11370);
or U12789 (N_12789,N_11019,N_11259);
xnor U12790 (N_12790,N_11253,N_11443);
or U12791 (N_12791,N_11245,N_11134);
or U12792 (N_12792,N_11627,N_11604);
or U12793 (N_12793,N_11837,N_11015);
or U12794 (N_12794,N_11884,N_11448);
nor U12795 (N_12795,N_11765,N_10893);
xor U12796 (N_12796,N_10916,N_11810);
nand U12797 (N_12797,N_11900,N_11434);
or U12798 (N_12798,N_11988,N_11859);
or U12799 (N_12799,N_11605,N_11773);
or U12800 (N_12800,N_11443,N_10808);
nand U12801 (N_12801,N_10800,N_11344);
and U12802 (N_12802,N_11282,N_11486);
and U12803 (N_12803,N_11254,N_11672);
nand U12804 (N_12804,N_11375,N_11499);
and U12805 (N_12805,N_10971,N_11170);
and U12806 (N_12806,N_10806,N_11121);
nor U12807 (N_12807,N_11754,N_11890);
or U12808 (N_12808,N_11724,N_11343);
nor U12809 (N_12809,N_11825,N_11657);
and U12810 (N_12810,N_11148,N_10820);
nor U12811 (N_12811,N_10896,N_11112);
or U12812 (N_12812,N_11712,N_11516);
nor U12813 (N_12813,N_11793,N_11431);
and U12814 (N_12814,N_10988,N_11257);
or U12815 (N_12815,N_11840,N_10894);
and U12816 (N_12816,N_10873,N_11950);
and U12817 (N_12817,N_11676,N_11754);
and U12818 (N_12818,N_11200,N_11841);
nand U12819 (N_12819,N_11767,N_11614);
nand U12820 (N_12820,N_11628,N_11386);
nor U12821 (N_12821,N_11326,N_11689);
xnor U12822 (N_12822,N_10919,N_11145);
xor U12823 (N_12823,N_11985,N_11841);
and U12824 (N_12824,N_11035,N_11162);
nand U12825 (N_12825,N_11697,N_11662);
or U12826 (N_12826,N_11513,N_11940);
nor U12827 (N_12827,N_11706,N_11950);
and U12828 (N_12828,N_11644,N_11059);
and U12829 (N_12829,N_11458,N_11270);
nor U12830 (N_12830,N_11597,N_11907);
nor U12831 (N_12831,N_11905,N_11365);
or U12832 (N_12832,N_11535,N_11039);
nor U12833 (N_12833,N_11766,N_11477);
and U12834 (N_12834,N_11915,N_11183);
xnor U12835 (N_12835,N_11733,N_10985);
nor U12836 (N_12836,N_11014,N_11013);
xor U12837 (N_12837,N_11889,N_10987);
or U12838 (N_12838,N_11616,N_11572);
xor U12839 (N_12839,N_11691,N_11305);
nand U12840 (N_12840,N_11126,N_11597);
nand U12841 (N_12841,N_11030,N_10861);
and U12842 (N_12842,N_10827,N_11660);
and U12843 (N_12843,N_11001,N_11947);
xnor U12844 (N_12844,N_11022,N_11285);
or U12845 (N_12845,N_11151,N_11519);
nor U12846 (N_12846,N_10996,N_11444);
and U12847 (N_12847,N_11444,N_11307);
nand U12848 (N_12848,N_10903,N_11204);
nor U12849 (N_12849,N_11928,N_11634);
or U12850 (N_12850,N_11265,N_11837);
and U12851 (N_12851,N_11781,N_11029);
or U12852 (N_12852,N_11581,N_11783);
or U12853 (N_12853,N_11647,N_11915);
nor U12854 (N_12854,N_11482,N_11076);
nand U12855 (N_12855,N_11600,N_11634);
xnor U12856 (N_12856,N_11325,N_11655);
xor U12857 (N_12857,N_11347,N_11238);
and U12858 (N_12858,N_11716,N_11489);
and U12859 (N_12859,N_11612,N_11787);
nand U12860 (N_12860,N_11324,N_11851);
or U12861 (N_12861,N_10889,N_10954);
nand U12862 (N_12862,N_11267,N_11498);
and U12863 (N_12863,N_11877,N_10803);
or U12864 (N_12864,N_11579,N_11227);
xnor U12865 (N_12865,N_11678,N_11719);
xnor U12866 (N_12866,N_11016,N_11193);
nand U12867 (N_12867,N_11077,N_11393);
nand U12868 (N_12868,N_10882,N_11750);
nor U12869 (N_12869,N_10842,N_11751);
nand U12870 (N_12870,N_11172,N_11762);
xor U12871 (N_12871,N_11587,N_11602);
or U12872 (N_12872,N_11213,N_11111);
or U12873 (N_12873,N_10985,N_11388);
xor U12874 (N_12874,N_11526,N_10809);
nor U12875 (N_12875,N_11150,N_11941);
and U12876 (N_12876,N_11066,N_11202);
and U12877 (N_12877,N_11855,N_11955);
nor U12878 (N_12878,N_11348,N_11027);
nor U12879 (N_12879,N_11330,N_11254);
xnor U12880 (N_12880,N_11171,N_11468);
xor U12881 (N_12881,N_11134,N_11620);
xnor U12882 (N_12882,N_11390,N_11295);
nand U12883 (N_12883,N_11365,N_11932);
and U12884 (N_12884,N_10994,N_11988);
xnor U12885 (N_12885,N_10811,N_11761);
and U12886 (N_12886,N_10931,N_11433);
and U12887 (N_12887,N_11332,N_10818);
xor U12888 (N_12888,N_11979,N_11642);
xnor U12889 (N_12889,N_11694,N_11222);
nor U12890 (N_12890,N_11405,N_10897);
xor U12891 (N_12891,N_11983,N_11711);
nand U12892 (N_12892,N_10838,N_10876);
and U12893 (N_12893,N_11110,N_11144);
xor U12894 (N_12894,N_11877,N_11860);
xor U12895 (N_12895,N_11175,N_11627);
and U12896 (N_12896,N_11827,N_11951);
and U12897 (N_12897,N_11464,N_11834);
nand U12898 (N_12898,N_11144,N_11872);
and U12899 (N_12899,N_11172,N_11099);
and U12900 (N_12900,N_10828,N_11630);
nand U12901 (N_12901,N_11490,N_11684);
and U12902 (N_12902,N_11952,N_10858);
nand U12903 (N_12903,N_10911,N_11663);
nor U12904 (N_12904,N_11759,N_10894);
xnor U12905 (N_12905,N_11196,N_11087);
or U12906 (N_12906,N_11496,N_11503);
nand U12907 (N_12907,N_11243,N_11182);
and U12908 (N_12908,N_11797,N_11776);
and U12909 (N_12909,N_11835,N_11336);
nor U12910 (N_12910,N_11906,N_11659);
nor U12911 (N_12911,N_11686,N_11750);
and U12912 (N_12912,N_10880,N_11620);
nand U12913 (N_12913,N_10901,N_11108);
or U12914 (N_12914,N_11262,N_11996);
nand U12915 (N_12915,N_11962,N_10825);
nor U12916 (N_12916,N_11849,N_11286);
xor U12917 (N_12917,N_11837,N_11670);
nor U12918 (N_12918,N_11682,N_11946);
or U12919 (N_12919,N_11519,N_11874);
nor U12920 (N_12920,N_11632,N_11222);
xor U12921 (N_12921,N_11694,N_11261);
nand U12922 (N_12922,N_10927,N_11662);
and U12923 (N_12923,N_11995,N_11562);
nor U12924 (N_12924,N_11377,N_11289);
and U12925 (N_12925,N_11389,N_11565);
nor U12926 (N_12926,N_11160,N_11155);
and U12927 (N_12927,N_10848,N_11362);
or U12928 (N_12928,N_11452,N_10826);
xnor U12929 (N_12929,N_11433,N_11325);
or U12930 (N_12930,N_11022,N_11305);
or U12931 (N_12931,N_10875,N_11518);
xnor U12932 (N_12932,N_11805,N_11539);
or U12933 (N_12933,N_11791,N_10812);
and U12934 (N_12934,N_11203,N_11653);
and U12935 (N_12935,N_11610,N_11257);
or U12936 (N_12936,N_11745,N_11291);
and U12937 (N_12937,N_11741,N_11677);
xnor U12938 (N_12938,N_11155,N_11607);
nand U12939 (N_12939,N_11736,N_11645);
xnor U12940 (N_12940,N_11703,N_10804);
xor U12941 (N_12941,N_11152,N_11162);
and U12942 (N_12942,N_11301,N_10864);
or U12943 (N_12943,N_11460,N_11158);
or U12944 (N_12944,N_11842,N_11092);
and U12945 (N_12945,N_10984,N_11247);
nand U12946 (N_12946,N_11839,N_11874);
nor U12947 (N_12947,N_11905,N_11098);
xnor U12948 (N_12948,N_10842,N_11604);
xor U12949 (N_12949,N_11564,N_11210);
or U12950 (N_12950,N_11411,N_11382);
nor U12951 (N_12951,N_11698,N_11762);
nand U12952 (N_12952,N_11808,N_11903);
or U12953 (N_12953,N_11109,N_11432);
nand U12954 (N_12954,N_10810,N_11489);
or U12955 (N_12955,N_10954,N_11958);
xor U12956 (N_12956,N_11647,N_11639);
nor U12957 (N_12957,N_10861,N_11478);
nand U12958 (N_12958,N_11125,N_11467);
xnor U12959 (N_12959,N_11633,N_10943);
and U12960 (N_12960,N_11676,N_11748);
nor U12961 (N_12961,N_11983,N_11933);
nor U12962 (N_12962,N_11754,N_11321);
or U12963 (N_12963,N_11354,N_11896);
xor U12964 (N_12964,N_11412,N_10952);
xor U12965 (N_12965,N_11661,N_11482);
nor U12966 (N_12966,N_11962,N_11629);
xnor U12967 (N_12967,N_11827,N_11351);
or U12968 (N_12968,N_11197,N_10900);
nand U12969 (N_12969,N_11594,N_11753);
or U12970 (N_12970,N_11543,N_11652);
and U12971 (N_12971,N_11846,N_11763);
and U12972 (N_12972,N_11748,N_10966);
nor U12973 (N_12973,N_10901,N_11089);
xnor U12974 (N_12974,N_11034,N_10873);
or U12975 (N_12975,N_11336,N_11163);
nand U12976 (N_12976,N_11819,N_11412);
or U12977 (N_12977,N_11341,N_11130);
and U12978 (N_12978,N_11755,N_11260);
or U12979 (N_12979,N_11909,N_11019);
and U12980 (N_12980,N_11285,N_11653);
nor U12981 (N_12981,N_11849,N_11791);
nand U12982 (N_12982,N_11152,N_11498);
nand U12983 (N_12983,N_11744,N_11538);
nand U12984 (N_12984,N_11388,N_11614);
xor U12985 (N_12985,N_11486,N_11544);
and U12986 (N_12986,N_10870,N_11152);
nand U12987 (N_12987,N_11578,N_11412);
nor U12988 (N_12988,N_11883,N_11701);
or U12989 (N_12989,N_11427,N_10807);
xnor U12990 (N_12990,N_11174,N_11638);
or U12991 (N_12991,N_11543,N_11535);
and U12992 (N_12992,N_11005,N_11502);
or U12993 (N_12993,N_11266,N_11888);
or U12994 (N_12994,N_11590,N_11113);
nor U12995 (N_12995,N_11870,N_11705);
nor U12996 (N_12996,N_11970,N_11429);
or U12997 (N_12997,N_11441,N_11621);
and U12998 (N_12998,N_11076,N_11040);
xor U12999 (N_12999,N_11637,N_11976);
nor U13000 (N_13000,N_11701,N_11575);
and U13001 (N_13001,N_11526,N_11234);
nand U13002 (N_13002,N_10961,N_11305);
nand U13003 (N_13003,N_11569,N_11032);
and U13004 (N_13004,N_11070,N_10960);
and U13005 (N_13005,N_11771,N_11039);
and U13006 (N_13006,N_10968,N_11917);
nor U13007 (N_13007,N_11040,N_11399);
nand U13008 (N_13008,N_10933,N_11256);
xor U13009 (N_13009,N_11083,N_11363);
nor U13010 (N_13010,N_11437,N_11971);
and U13011 (N_13011,N_11422,N_11288);
nand U13012 (N_13012,N_10871,N_11158);
nand U13013 (N_13013,N_11947,N_11117);
and U13014 (N_13014,N_11719,N_11177);
nor U13015 (N_13015,N_11514,N_11873);
or U13016 (N_13016,N_11175,N_11586);
or U13017 (N_13017,N_11618,N_10923);
and U13018 (N_13018,N_11293,N_11142);
nor U13019 (N_13019,N_11023,N_11219);
xnor U13020 (N_13020,N_11131,N_11269);
and U13021 (N_13021,N_11151,N_11196);
xnor U13022 (N_13022,N_11303,N_11142);
nor U13023 (N_13023,N_11902,N_11551);
xnor U13024 (N_13024,N_11574,N_11224);
nor U13025 (N_13025,N_10965,N_11094);
or U13026 (N_13026,N_11712,N_10857);
and U13027 (N_13027,N_11932,N_11215);
or U13028 (N_13028,N_11651,N_11481);
nand U13029 (N_13029,N_11403,N_11085);
nor U13030 (N_13030,N_11911,N_11608);
xnor U13031 (N_13031,N_11971,N_11539);
and U13032 (N_13032,N_11094,N_11453);
nand U13033 (N_13033,N_10958,N_11696);
and U13034 (N_13034,N_10822,N_11193);
nand U13035 (N_13035,N_11490,N_11247);
or U13036 (N_13036,N_11543,N_11128);
nor U13037 (N_13037,N_11024,N_11123);
xor U13038 (N_13038,N_10958,N_11100);
and U13039 (N_13039,N_11719,N_11663);
nand U13040 (N_13040,N_11861,N_11278);
and U13041 (N_13041,N_11827,N_11288);
nand U13042 (N_13042,N_11884,N_10845);
nand U13043 (N_13043,N_10878,N_11829);
or U13044 (N_13044,N_11398,N_10915);
or U13045 (N_13045,N_11617,N_11247);
nor U13046 (N_13046,N_11663,N_10948);
nor U13047 (N_13047,N_11399,N_10855);
nor U13048 (N_13048,N_11774,N_10831);
xnor U13049 (N_13049,N_11413,N_11797);
or U13050 (N_13050,N_11106,N_11476);
nand U13051 (N_13051,N_11722,N_11853);
xnor U13052 (N_13052,N_10882,N_11923);
and U13053 (N_13053,N_11393,N_11011);
xnor U13054 (N_13054,N_11413,N_10890);
and U13055 (N_13055,N_10947,N_11585);
nand U13056 (N_13056,N_11197,N_11188);
and U13057 (N_13057,N_11627,N_11978);
xnor U13058 (N_13058,N_11952,N_10931);
and U13059 (N_13059,N_11614,N_11592);
nor U13060 (N_13060,N_11548,N_11056);
and U13061 (N_13061,N_11713,N_11399);
or U13062 (N_13062,N_11132,N_11637);
or U13063 (N_13063,N_11036,N_11040);
xnor U13064 (N_13064,N_11188,N_11293);
nand U13065 (N_13065,N_11197,N_11788);
or U13066 (N_13066,N_10846,N_11212);
or U13067 (N_13067,N_11725,N_11145);
and U13068 (N_13068,N_11589,N_11156);
or U13069 (N_13069,N_11323,N_11679);
nand U13070 (N_13070,N_10978,N_11716);
nand U13071 (N_13071,N_11050,N_11527);
xor U13072 (N_13072,N_10872,N_11681);
nand U13073 (N_13073,N_11696,N_11502);
and U13074 (N_13074,N_11046,N_10834);
or U13075 (N_13075,N_11659,N_11898);
nor U13076 (N_13076,N_11363,N_10958);
or U13077 (N_13077,N_11061,N_11851);
xnor U13078 (N_13078,N_11071,N_11950);
or U13079 (N_13079,N_11180,N_11071);
nand U13080 (N_13080,N_10868,N_11230);
and U13081 (N_13081,N_11725,N_11074);
and U13082 (N_13082,N_10836,N_11656);
nand U13083 (N_13083,N_11976,N_11844);
nor U13084 (N_13084,N_10966,N_11867);
nor U13085 (N_13085,N_11422,N_10966);
nand U13086 (N_13086,N_11521,N_11379);
nor U13087 (N_13087,N_11755,N_10883);
xnor U13088 (N_13088,N_11684,N_11441);
xor U13089 (N_13089,N_11056,N_10977);
nor U13090 (N_13090,N_11272,N_11354);
and U13091 (N_13091,N_11308,N_11164);
and U13092 (N_13092,N_11419,N_10807);
nand U13093 (N_13093,N_10878,N_10909);
xor U13094 (N_13094,N_11389,N_11027);
or U13095 (N_13095,N_10800,N_11137);
or U13096 (N_13096,N_10827,N_11518);
xnor U13097 (N_13097,N_10913,N_11104);
or U13098 (N_13098,N_11877,N_11473);
or U13099 (N_13099,N_11910,N_11337);
and U13100 (N_13100,N_11770,N_11062);
nor U13101 (N_13101,N_10901,N_11684);
xnor U13102 (N_13102,N_11270,N_11273);
nor U13103 (N_13103,N_11057,N_11113);
nor U13104 (N_13104,N_11497,N_11363);
nor U13105 (N_13105,N_11670,N_11228);
nand U13106 (N_13106,N_11094,N_11762);
xor U13107 (N_13107,N_11824,N_11964);
xor U13108 (N_13108,N_11057,N_11788);
or U13109 (N_13109,N_11159,N_11978);
and U13110 (N_13110,N_11429,N_11608);
nor U13111 (N_13111,N_11259,N_11869);
nor U13112 (N_13112,N_11236,N_11467);
xnor U13113 (N_13113,N_11435,N_11587);
nor U13114 (N_13114,N_11842,N_11648);
xnor U13115 (N_13115,N_11799,N_10953);
xor U13116 (N_13116,N_11010,N_11224);
or U13117 (N_13117,N_11585,N_11756);
nor U13118 (N_13118,N_11864,N_11788);
nand U13119 (N_13119,N_11157,N_11401);
and U13120 (N_13120,N_10854,N_11817);
nand U13121 (N_13121,N_11722,N_11666);
nor U13122 (N_13122,N_11515,N_11033);
and U13123 (N_13123,N_11900,N_10893);
xor U13124 (N_13124,N_11809,N_11420);
xor U13125 (N_13125,N_11656,N_11581);
nand U13126 (N_13126,N_11334,N_11177);
nor U13127 (N_13127,N_11503,N_10800);
or U13128 (N_13128,N_11230,N_11597);
and U13129 (N_13129,N_11009,N_11261);
xor U13130 (N_13130,N_11633,N_11269);
xor U13131 (N_13131,N_10925,N_11166);
and U13132 (N_13132,N_11373,N_11220);
nand U13133 (N_13133,N_11776,N_11963);
nand U13134 (N_13134,N_11853,N_11154);
nand U13135 (N_13135,N_11671,N_11898);
xor U13136 (N_13136,N_11642,N_11889);
and U13137 (N_13137,N_11752,N_10916);
and U13138 (N_13138,N_11472,N_11246);
xnor U13139 (N_13139,N_11573,N_11360);
and U13140 (N_13140,N_11968,N_11055);
or U13141 (N_13141,N_11339,N_11447);
or U13142 (N_13142,N_11596,N_11400);
nor U13143 (N_13143,N_10916,N_11575);
or U13144 (N_13144,N_10905,N_11708);
nand U13145 (N_13145,N_10827,N_10981);
nand U13146 (N_13146,N_11955,N_11337);
xor U13147 (N_13147,N_10926,N_11754);
and U13148 (N_13148,N_10872,N_11137);
xnor U13149 (N_13149,N_11105,N_11412);
xnor U13150 (N_13150,N_11621,N_11077);
and U13151 (N_13151,N_11256,N_11294);
nand U13152 (N_13152,N_11861,N_11085);
nor U13153 (N_13153,N_11105,N_11094);
and U13154 (N_13154,N_10833,N_11554);
nor U13155 (N_13155,N_11924,N_11263);
nand U13156 (N_13156,N_10907,N_11411);
or U13157 (N_13157,N_11119,N_11173);
nor U13158 (N_13158,N_11130,N_11044);
and U13159 (N_13159,N_11542,N_11190);
xnor U13160 (N_13160,N_11299,N_11235);
nor U13161 (N_13161,N_11571,N_11640);
nand U13162 (N_13162,N_10977,N_11466);
nand U13163 (N_13163,N_11120,N_10829);
and U13164 (N_13164,N_11915,N_11637);
xnor U13165 (N_13165,N_11816,N_11144);
nand U13166 (N_13166,N_11804,N_11289);
or U13167 (N_13167,N_10983,N_11480);
nand U13168 (N_13168,N_11923,N_11015);
and U13169 (N_13169,N_11752,N_11570);
and U13170 (N_13170,N_11012,N_10857);
nor U13171 (N_13171,N_10862,N_11831);
and U13172 (N_13172,N_11297,N_11626);
and U13173 (N_13173,N_11955,N_11320);
nor U13174 (N_13174,N_11181,N_11788);
nand U13175 (N_13175,N_10985,N_10999);
nand U13176 (N_13176,N_11876,N_11341);
or U13177 (N_13177,N_11264,N_11705);
nor U13178 (N_13178,N_11053,N_11604);
or U13179 (N_13179,N_11153,N_11384);
or U13180 (N_13180,N_11212,N_10935);
xnor U13181 (N_13181,N_11725,N_11688);
nand U13182 (N_13182,N_11165,N_11894);
and U13183 (N_13183,N_11103,N_11514);
xor U13184 (N_13184,N_11276,N_11777);
nor U13185 (N_13185,N_10831,N_11829);
nor U13186 (N_13186,N_11559,N_11245);
xnor U13187 (N_13187,N_11498,N_11854);
nand U13188 (N_13188,N_11145,N_10975);
nor U13189 (N_13189,N_11632,N_11162);
and U13190 (N_13190,N_11245,N_11545);
nor U13191 (N_13191,N_11733,N_11009);
xnor U13192 (N_13192,N_11400,N_11587);
nand U13193 (N_13193,N_11731,N_11043);
xor U13194 (N_13194,N_10845,N_10842);
and U13195 (N_13195,N_11725,N_10849);
and U13196 (N_13196,N_11999,N_11569);
or U13197 (N_13197,N_11305,N_11236);
nor U13198 (N_13198,N_10819,N_11063);
and U13199 (N_13199,N_11055,N_10904);
or U13200 (N_13200,N_12768,N_13095);
nor U13201 (N_13201,N_12437,N_12970);
nand U13202 (N_13202,N_12564,N_12965);
nand U13203 (N_13203,N_12741,N_13128);
xor U13204 (N_13204,N_12602,N_12210);
or U13205 (N_13205,N_12953,N_12081);
and U13206 (N_13206,N_12509,N_12826);
nand U13207 (N_13207,N_12146,N_12102);
nor U13208 (N_13208,N_12460,N_12021);
and U13209 (N_13209,N_12462,N_12205);
nor U13210 (N_13210,N_12083,N_12891);
and U13211 (N_13211,N_12774,N_12998);
and U13212 (N_13212,N_12890,N_12230);
nand U13213 (N_13213,N_12655,N_12139);
nor U13214 (N_13214,N_12914,N_12666);
and U13215 (N_13215,N_12504,N_12757);
nand U13216 (N_13216,N_12783,N_12024);
xnor U13217 (N_13217,N_12821,N_12915);
nand U13218 (N_13218,N_12060,N_12232);
nor U13219 (N_13219,N_12517,N_12313);
and U13220 (N_13220,N_12004,N_12173);
nor U13221 (N_13221,N_12677,N_12749);
and U13222 (N_13222,N_12419,N_12416);
or U13223 (N_13223,N_12179,N_13132);
nand U13224 (N_13224,N_13153,N_12928);
nand U13225 (N_13225,N_12219,N_13069);
and U13226 (N_13226,N_13135,N_12761);
nand U13227 (N_13227,N_12856,N_12239);
xnor U13228 (N_13228,N_12265,N_12901);
or U13229 (N_13229,N_12252,N_12626);
nor U13230 (N_13230,N_12364,N_12939);
nand U13231 (N_13231,N_12849,N_12759);
nor U13232 (N_13232,N_12196,N_12334);
and U13233 (N_13233,N_12022,N_12777);
or U13234 (N_13234,N_12264,N_12199);
nand U13235 (N_13235,N_12319,N_12431);
xor U13236 (N_13236,N_12474,N_12440);
nand U13237 (N_13237,N_13166,N_12430);
xor U13238 (N_13238,N_13092,N_12015);
xor U13239 (N_13239,N_12845,N_13102);
xnor U13240 (N_13240,N_12244,N_13001);
nor U13241 (N_13241,N_12417,N_12320);
nor U13242 (N_13242,N_13124,N_12099);
nor U13243 (N_13243,N_12858,N_12609);
nand U13244 (N_13244,N_13007,N_12508);
nand U13245 (N_13245,N_13081,N_12895);
nand U13246 (N_13246,N_12436,N_12046);
nand U13247 (N_13247,N_12753,N_12715);
or U13248 (N_13248,N_12710,N_12218);
xnor U13249 (N_13249,N_12043,N_12036);
xnor U13250 (N_13250,N_12461,N_12476);
nand U13251 (N_13251,N_12876,N_12916);
nand U13252 (N_13252,N_13099,N_12041);
nand U13253 (N_13253,N_12190,N_12289);
xor U13254 (N_13254,N_12296,N_12925);
xor U13255 (N_13255,N_12276,N_13074);
or U13256 (N_13256,N_13080,N_13048);
nand U13257 (N_13257,N_12087,N_13054);
nor U13258 (N_13258,N_12639,N_12279);
nand U13259 (N_13259,N_12799,N_12378);
and U13260 (N_13260,N_13148,N_12852);
xnor U13261 (N_13261,N_12026,N_12412);
or U13262 (N_13262,N_12310,N_12348);
nand U13263 (N_13263,N_12453,N_12217);
nand U13264 (N_13264,N_12178,N_13088);
or U13265 (N_13265,N_12381,N_12337);
nand U13266 (N_13266,N_12134,N_12595);
xnor U13267 (N_13267,N_12784,N_12750);
and U13268 (N_13268,N_12803,N_13006);
or U13269 (N_13269,N_12933,N_12158);
nor U13270 (N_13270,N_12851,N_13056);
nor U13271 (N_13271,N_12306,N_12778);
nand U13272 (N_13272,N_12137,N_13175);
and U13273 (N_13273,N_12760,N_12231);
nand U13274 (N_13274,N_12128,N_12580);
nor U13275 (N_13275,N_13022,N_12883);
xnor U13276 (N_13276,N_12367,N_12910);
or U13277 (N_13277,N_12305,N_12186);
nand U13278 (N_13278,N_12303,N_12284);
nand U13279 (N_13279,N_12815,N_12391);
xor U13280 (N_13280,N_12725,N_12513);
nor U13281 (N_13281,N_12469,N_12325);
xor U13282 (N_13282,N_12298,N_12059);
and U13283 (N_13283,N_12604,N_12383);
or U13284 (N_13284,N_12827,N_12828);
and U13285 (N_13285,N_12432,N_12308);
nor U13286 (N_13286,N_12726,N_12954);
xnor U13287 (N_13287,N_12703,N_12272);
nor U13288 (N_13288,N_12119,N_12352);
or U13289 (N_13289,N_13151,N_13199);
nor U13290 (N_13290,N_12615,N_13017);
nand U13291 (N_13291,N_12896,N_12999);
nor U13292 (N_13292,N_12012,N_12680);
xnor U13293 (N_13293,N_13012,N_12285);
nor U13294 (N_13294,N_13093,N_12660);
and U13295 (N_13295,N_12009,N_12067);
xnor U13296 (N_13296,N_12362,N_12687);
nand U13297 (N_13297,N_12528,N_12645);
nor U13298 (N_13298,N_12003,N_12405);
xor U13299 (N_13299,N_13169,N_12862);
or U13300 (N_13300,N_12736,N_12958);
nor U13301 (N_13301,N_12150,N_12502);
or U13302 (N_13302,N_13068,N_12397);
nor U13303 (N_13303,N_13086,N_12399);
nor U13304 (N_13304,N_12247,N_12038);
and U13305 (N_13305,N_12125,N_12002);
and U13306 (N_13306,N_12425,N_12568);
nand U13307 (N_13307,N_12787,N_12743);
nor U13308 (N_13308,N_13129,N_12452);
nor U13309 (N_13309,N_12200,N_13127);
xnor U13310 (N_13310,N_13005,N_12396);
and U13311 (N_13311,N_12734,N_12174);
and U13312 (N_13312,N_12940,N_13105);
xnor U13313 (N_13313,N_12457,N_12818);
nand U13314 (N_13314,N_12701,N_12160);
and U13315 (N_13315,N_12882,N_12535);
nor U13316 (N_13316,N_12945,N_12149);
nand U13317 (N_13317,N_12288,N_12658);
or U13318 (N_13318,N_12921,N_12860);
and U13319 (N_13319,N_12554,N_13042);
nor U13320 (N_13320,N_13167,N_13123);
and U13321 (N_13321,N_12808,N_13192);
nand U13322 (N_13322,N_13020,N_12147);
nor U13323 (N_13323,N_12506,N_12542);
nor U13324 (N_13324,N_12010,N_12114);
nand U13325 (N_13325,N_13030,N_12642);
nand U13326 (N_13326,N_12249,N_12817);
nor U13327 (N_13327,N_12105,N_12256);
or U13328 (N_13328,N_12985,N_12867);
and U13329 (N_13329,N_13155,N_12112);
xnor U13330 (N_13330,N_12014,N_12665);
xor U13331 (N_13331,N_12782,N_12234);
and U13332 (N_13332,N_13008,N_12855);
nor U13333 (N_13333,N_12592,N_12032);
xor U13334 (N_13334,N_12492,N_12468);
nor U13335 (N_13335,N_12488,N_12690);
or U13336 (N_13336,N_12140,N_12875);
or U13337 (N_13337,N_12421,N_12957);
nor U13338 (N_13338,N_12005,N_12829);
nand U13339 (N_13339,N_13004,N_12769);
nand U13340 (N_13340,N_13113,N_12669);
and U13341 (N_13341,N_13137,N_12300);
xor U13342 (N_13342,N_12129,N_12066);
or U13343 (N_13343,N_12152,N_12923);
nand U13344 (N_13344,N_12132,N_12772);
xor U13345 (N_13345,N_12964,N_13104);
and U13346 (N_13346,N_12547,N_13089);
nor U13347 (N_13347,N_12280,N_13110);
nor U13348 (N_13348,N_12667,N_12278);
or U13349 (N_13349,N_13173,N_12536);
or U13350 (N_13350,N_12927,N_13183);
nor U13351 (N_13351,N_12235,N_12368);
nand U13352 (N_13352,N_12865,N_12507);
xor U13353 (N_13353,N_12410,N_12512);
or U13354 (N_13354,N_12834,N_12044);
or U13355 (N_13355,N_12662,N_12541);
xnor U13356 (N_13356,N_13144,N_12900);
and U13357 (N_13357,N_12588,N_13186);
and U13358 (N_13358,N_12344,N_12972);
or U13359 (N_13359,N_12028,N_12409);
nand U13360 (N_13360,N_13114,N_13165);
or U13361 (N_13361,N_12880,N_12946);
and U13362 (N_13362,N_12806,N_13176);
xor U13363 (N_13363,N_13094,N_12370);
nor U13364 (N_13364,N_12093,N_12587);
xor U13365 (N_13365,N_12889,N_12637);
or U13366 (N_13366,N_12086,N_12020);
or U13367 (N_13367,N_12668,N_12395);
or U13368 (N_13368,N_13109,N_13061);
and U13369 (N_13369,N_12581,N_12401);
nand U13370 (N_13370,N_13096,N_12501);
or U13371 (N_13371,N_12908,N_12579);
or U13372 (N_13372,N_12560,N_12794);
xor U13373 (N_13373,N_12758,N_12649);
or U13374 (N_13374,N_12857,N_12089);
nand U13375 (N_13375,N_12268,N_12471);
nor U13376 (N_13376,N_13016,N_12798);
xor U13377 (N_13377,N_12770,N_12326);
or U13378 (N_13378,N_13120,N_12350);
nand U13379 (N_13379,N_12981,N_12311);
nor U13380 (N_13380,N_12566,N_13161);
and U13381 (N_13381,N_13041,N_12165);
and U13382 (N_13382,N_12553,N_12571);
xnor U13383 (N_13383,N_12648,N_12001);
xnor U13384 (N_13384,N_12072,N_12853);
or U13385 (N_13385,N_12459,N_12611);
or U13386 (N_13386,N_12766,N_12521);
or U13387 (N_13387,N_12586,N_12295);
nand U13388 (N_13388,N_12122,N_12810);
nor U13389 (N_13389,N_13097,N_12537);
nand U13390 (N_13390,N_12572,N_12847);
or U13391 (N_13391,N_12624,N_12569);
xor U13392 (N_13392,N_12540,N_13077);
and U13393 (N_13393,N_12355,N_12243);
nand U13394 (N_13394,N_12062,N_12627);
nand U13395 (N_13395,N_12106,N_12282);
xnor U13396 (N_13396,N_12893,N_13112);
nor U13397 (N_13397,N_12490,N_12640);
and U13398 (N_13398,N_12215,N_12483);
or U13399 (N_13399,N_12975,N_13023);
nor U13400 (N_13400,N_12987,N_12739);
and U13401 (N_13401,N_12878,N_12008);
xnor U13402 (N_13402,N_12992,N_12269);
nand U13403 (N_13403,N_13002,N_12248);
or U13404 (N_13404,N_13066,N_13131);
and U13405 (N_13405,N_13111,N_12470);
or U13406 (N_13406,N_12995,N_12450);
nor U13407 (N_13407,N_12404,N_13100);
nor U13408 (N_13408,N_13179,N_12061);
nor U13409 (N_13409,N_12562,N_12780);
and U13410 (N_13410,N_12740,N_12563);
xor U13411 (N_13411,N_12299,N_12717);
and U13412 (N_13412,N_13140,N_12793);
xor U13413 (N_13413,N_12451,N_12389);
or U13414 (N_13414,N_12127,N_13190);
xor U13415 (N_13415,N_13053,N_12801);
and U13416 (N_13416,N_12610,N_12063);
or U13417 (N_13417,N_12962,N_12156);
or U13418 (N_13418,N_12433,N_12455);
nand U13419 (N_13419,N_12124,N_12868);
nor U13420 (N_13420,N_12844,N_12598);
nand U13421 (N_13421,N_12790,N_12283);
nand U13422 (N_13422,N_12172,N_12816);
or U13423 (N_13423,N_12727,N_12123);
or U13424 (N_13424,N_12497,N_12966);
xnor U13425 (N_13425,N_12903,N_12529);
or U13426 (N_13426,N_12013,N_12924);
nand U13427 (N_13427,N_12719,N_12621);
and U13428 (N_13428,N_12053,N_13143);
xnor U13429 (N_13429,N_13130,N_12809);
nor U13430 (N_13430,N_13025,N_12700);
and U13431 (N_13431,N_12194,N_13082);
and U13432 (N_13432,N_12304,N_12275);
xor U13433 (N_13433,N_12494,N_13011);
and U13434 (N_13434,N_12804,N_12722);
xnor U13435 (N_13435,N_12735,N_12623);
xor U13436 (N_13436,N_12549,N_13058);
and U13437 (N_13437,N_12077,N_13116);
nand U13438 (N_13438,N_13121,N_12387);
xor U13439 (N_13439,N_12057,N_12162);
and U13440 (N_13440,N_12000,N_12756);
nand U13441 (N_13441,N_12336,N_12380);
nor U13442 (N_13442,N_12351,N_12438);
or U13443 (N_13443,N_12518,N_12088);
or U13444 (N_13444,N_13154,N_13098);
nand U13445 (N_13445,N_13091,N_12824);
xnor U13446 (N_13446,N_12820,N_12406);
xor U13447 (N_13447,N_12225,N_12271);
nor U13448 (N_13448,N_12187,N_12084);
xnor U13449 (N_13449,N_12616,N_13162);
and U13450 (N_13450,N_12175,N_13052);
nor U13451 (N_13451,N_12767,N_12257);
nor U13452 (N_13452,N_12585,N_13073);
and U13453 (N_13453,N_12797,N_12045);
xor U13454 (N_13454,N_12449,N_12565);
nand U13455 (N_13455,N_12170,N_12789);
and U13456 (N_13456,N_12415,N_12944);
and U13457 (N_13457,N_12143,N_12974);
and U13458 (N_13458,N_12653,N_12467);
xor U13459 (N_13459,N_12906,N_12591);
nand U13460 (N_13460,N_12188,N_12839);
or U13461 (N_13461,N_12751,N_13015);
xnor U13462 (N_13462,N_12407,N_13046);
xor U13463 (N_13463,N_12493,N_12811);
or U13464 (N_13464,N_12447,N_12967);
nand U13465 (N_13465,N_12241,N_12495);
nand U13466 (N_13466,N_12643,N_12500);
and U13467 (N_13467,N_13037,N_12076);
or U13468 (N_13468,N_12301,N_12154);
or U13469 (N_13469,N_13139,N_12221);
xor U13470 (N_13470,N_12683,N_12078);
and U13471 (N_13471,N_12646,N_12894);
and U13472 (N_13472,N_12525,N_12385);
nand U13473 (N_13473,N_12211,N_12245);
and U13474 (N_13474,N_12531,N_12636);
nand U13475 (N_13475,N_12222,N_12532);
nand U13476 (N_13476,N_12443,N_12873);
nor U13477 (N_13477,N_12049,N_12273);
nand U13478 (N_13478,N_12403,N_12213);
nor U13479 (N_13479,N_12161,N_12812);
or U13480 (N_13480,N_13071,N_12842);
nand U13481 (N_13481,N_12699,N_12167);
and U13482 (N_13482,N_12929,N_13163);
and U13483 (N_13483,N_12075,N_12181);
nor U13484 (N_13484,N_12590,N_12074);
or U13485 (N_13485,N_12177,N_12208);
nand U13486 (N_13486,N_12679,N_12613);
nor U13487 (N_13487,N_12333,N_12055);
and U13488 (N_13488,N_12664,N_12192);
nand U13489 (N_13489,N_12557,N_12422);
nand U13490 (N_13490,N_12442,N_12328);
nor U13491 (N_13491,N_12386,N_12491);
and U13492 (N_13492,N_12229,N_12551);
nor U13493 (N_13493,N_12212,N_12850);
xor U13494 (N_13494,N_12109,N_13152);
xor U13495 (N_13495,N_13141,N_12704);
or U13496 (N_13496,N_12477,N_12654);
or U13497 (N_13497,N_12582,N_12548);
or U13498 (N_13498,N_12047,N_12169);
nor U13499 (N_13499,N_12733,N_12151);
or U13500 (N_13500,N_12358,N_12366);
xnor U13501 (N_13501,N_12323,N_12515);
and U13502 (N_13502,N_13159,N_12672);
nand U13503 (N_13503,N_12103,N_12365);
xnor U13504 (N_13504,N_12176,N_12498);
nand U13505 (N_13505,N_12496,N_12201);
xor U13506 (N_13506,N_12423,N_12136);
and U13507 (N_13507,N_12071,N_12971);
or U13508 (N_13508,N_12155,N_12746);
nand U13509 (N_13509,N_12877,N_12872);
nor U13510 (N_13510,N_12342,N_12792);
or U13511 (N_13511,N_12262,N_12372);
or U13512 (N_13512,N_12373,N_12718);
or U13513 (N_13513,N_12731,N_12835);
nor U13514 (N_13514,N_12538,N_12561);
xnor U13515 (N_13515,N_12870,N_12110);
nand U13516 (N_13516,N_12938,N_12258);
xor U13517 (N_13517,N_12831,N_12897);
nor U13518 (N_13518,N_13138,N_12133);
xnor U13519 (N_13519,N_12085,N_12730);
or U13520 (N_13520,N_12315,N_12499);
xor U13521 (N_13521,N_12121,N_12709);
and U13522 (N_13522,N_12577,N_12879);
nor U13523 (N_13523,N_12448,N_12327);
xnor U13524 (N_13524,N_12206,N_13064);
nand U13525 (N_13525,N_12312,N_12054);
xnor U13526 (N_13526,N_12426,N_12707);
nand U13527 (N_13527,N_12597,N_13039);
and U13528 (N_13528,N_12874,N_13031);
xnor U13529 (N_13529,N_12101,N_12356);
nor U13530 (N_13530,N_12374,N_12822);
or U13531 (N_13531,N_13196,N_12267);
nor U13532 (N_13532,N_12104,N_12632);
nor U13533 (N_13533,N_12745,N_12318);
or U13534 (N_13534,N_12260,N_13055);
or U13535 (N_13535,N_12228,N_12107);
and U13536 (N_13536,N_13085,N_13119);
xnor U13537 (N_13537,N_12435,N_12684);
nor U13538 (N_13538,N_13146,N_12473);
xor U13539 (N_13539,N_12785,N_12918);
xnor U13540 (N_13540,N_12837,N_12293);
nor U13541 (N_13541,N_13014,N_12781);
or U13542 (N_13542,N_12520,N_13003);
xor U13543 (N_13543,N_12223,N_12691);
and U13544 (N_13544,N_12543,N_12661);
or U13545 (N_13545,N_12070,N_13084);
and U13546 (N_13546,N_13051,N_12016);
xnor U13547 (N_13547,N_12936,N_12130);
nor U13548 (N_13548,N_12911,N_12742);
nand U13549 (N_13549,N_13028,N_12487);
and U13550 (N_13550,N_12763,N_12384);
xor U13551 (N_13551,N_13072,N_12899);
nand U13552 (N_13552,N_12912,N_12671);
or U13553 (N_13553,N_12343,N_12287);
nor U13554 (N_13554,N_13009,N_13194);
nand U13555 (N_13555,N_12266,N_13065);
or U13556 (N_13556,N_12398,N_12802);
or U13557 (N_13557,N_12111,N_12614);
nand U13558 (N_13558,N_12065,N_12377);
xnor U13559 (N_13559,N_12148,N_13156);
nor U13560 (N_13560,N_12204,N_12079);
nor U13561 (N_13561,N_13024,N_12574);
and U13562 (N_13562,N_12338,N_12465);
nand U13563 (N_13563,N_13060,N_12920);
or U13564 (N_13564,N_12138,N_12961);
or U13565 (N_13565,N_12676,N_13126);
xnor U13566 (N_13566,N_12558,N_13150);
and U13567 (N_13567,N_12729,N_13164);
and U13568 (N_13568,N_12446,N_13021);
xnor U13569 (N_13569,N_12357,N_13171);
xor U13570 (N_13570,N_12902,N_12854);
nand U13571 (N_13571,N_12080,N_12686);
nand U13572 (N_13572,N_12779,N_12570);
and U13573 (N_13573,N_12556,N_12479);
nor U13574 (N_13574,N_13103,N_12048);
nor U13575 (N_13575,N_12108,N_12115);
nor U13576 (N_13576,N_12445,N_12776);
or U13577 (N_13577,N_12420,N_12051);
xnor U13578 (N_13578,N_12552,N_13087);
xnor U13579 (N_13579,N_12935,N_12913);
xor U13580 (N_13580,N_12317,N_12250);
nand U13581 (N_13581,N_12600,N_12444);
and U13582 (N_13582,N_12594,N_12884);
xnor U13583 (N_13583,N_12788,N_12530);
or U13584 (N_13584,N_13045,N_12991);
xor U13585 (N_13585,N_12764,N_12029);
nor U13586 (N_13586,N_13083,N_13117);
and U13587 (N_13587,N_13115,N_12682);
and U13588 (N_13588,N_12097,N_12830);
nand U13589 (N_13589,N_12263,N_13108);
nand U13590 (N_13590,N_12932,N_12617);
and U13591 (N_13591,N_12599,N_12237);
nor U13592 (N_13592,N_12486,N_13178);
nand U13593 (N_13593,N_12324,N_12618);
nand U13594 (N_13594,N_12361,N_12836);
and U13595 (N_13595,N_12354,N_13147);
xnor U13596 (N_13596,N_12706,N_12456);
nor U13597 (N_13597,N_12322,N_12724);
nand U13598 (N_13598,N_13181,N_12567);
or U13599 (N_13599,N_12534,N_12064);
xor U13600 (N_13600,N_12331,N_12674);
nand U13601 (N_13601,N_12702,N_12441);
nor U13602 (N_13602,N_12650,N_12379);
nand U13603 (N_13603,N_12226,N_12904);
and U13604 (N_13604,N_12197,N_12031);
nor U13605 (N_13605,N_12400,N_12994);
nand U13606 (N_13606,N_12346,N_12207);
nor U13607 (N_13607,N_12771,N_13174);
or U13608 (N_13608,N_12345,N_12330);
and U13609 (N_13609,N_12959,N_12622);
or U13610 (N_13610,N_12692,N_13191);
and U13611 (N_13611,N_12120,N_12737);
nor U13612 (N_13612,N_12340,N_12795);
nor U13613 (N_13613,N_13172,N_12678);
or U13614 (N_13614,N_12011,N_12369);
and U13615 (N_13615,N_12034,N_12117);
nand U13616 (N_13616,N_12628,N_13142);
xnor U13617 (N_13617,N_12869,N_12100);
xor U13618 (N_13618,N_12814,N_12428);
and U13619 (N_13619,N_12688,N_12274);
or U13620 (N_13620,N_12673,N_12171);
nand U13621 (N_13621,N_12307,N_12711);
nand U13622 (N_13622,N_12480,N_12620);
nand U13623 (N_13623,N_12976,N_12198);
nor U13624 (N_13624,N_13049,N_12286);
and U13625 (N_13625,N_13149,N_12805);
nor U13626 (N_13626,N_13198,N_12708);
or U13627 (N_13627,N_12630,N_12716);
nor U13628 (N_13628,N_12813,N_12555);
or U13629 (N_13629,N_12863,N_12848);
nand U13630 (N_13630,N_12596,N_12052);
or U13631 (N_13631,N_12224,N_13076);
and U13632 (N_13632,N_12712,N_12728);
xnor U13633 (N_13633,N_12159,N_12291);
nor U13634 (N_13634,N_12720,N_12098);
or U13635 (N_13635,N_12481,N_12589);
or U13636 (N_13636,N_12017,N_12157);
nand U13637 (N_13637,N_12281,N_12941);
nor U13638 (N_13638,N_12791,N_12978);
or U13639 (N_13639,N_12220,N_12754);
nor U13640 (N_13640,N_13013,N_12027);
nor U13641 (N_13641,N_13079,N_12183);
xor U13642 (N_13642,N_12090,N_13038);
nand U13643 (N_13643,N_12885,N_12464);
xnor U13644 (N_13644,N_12696,N_12619);
and U13645 (N_13645,N_12184,N_12638);
and U13646 (N_13646,N_12018,N_12539);
nor U13647 (N_13647,N_12576,N_13185);
or U13648 (N_13648,N_12656,N_12341);
nor U13649 (N_13649,N_12982,N_12533);
nor U13650 (N_13650,N_12056,N_13122);
nor U13651 (N_13651,N_12871,N_12675);
nor U13652 (N_13652,N_12261,N_12888);
xnor U13653 (N_13653,N_12775,N_12898);
xor U13654 (N_13654,N_12454,N_13044);
nor U13655 (N_13655,N_12050,N_12092);
nand U13656 (N_13656,N_12838,N_13043);
nand U13657 (N_13657,N_12182,N_12503);
or U13658 (N_13658,N_12514,N_12153);
and U13659 (N_13659,N_12697,N_12607);
xnor U13660 (N_13660,N_12713,N_12209);
nand U13661 (N_13661,N_12516,N_13189);
nor U13662 (N_13662,N_12359,N_13032);
nor U13663 (N_13663,N_12526,N_12037);
nor U13664 (N_13664,N_12141,N_12006);
xor U13665 (N_13665,N_12807,N_12524);
xnor U13666 (N_13666,N_12191,N_13134);
and U13667 (N_13667,N_13026,N_12253);
nand U13668 (N_13668,N_12892,N_13067);
and U13669 (N_13669,N_12723,N_12394);
xnor U13670 (N_13670,N_12511,N_13193);
and U13671 (N_13671,N_12773,N_12390);
xor U13672 (N_13672,N_13187,N_12068);
xor U13673 (N_13673,N_12113,N_12796);
and U13674 (N_13674,N_12952,N_12960);
nor U13675 (N_13675,N_13035,N_12866);
nand U13676 (N_13676,N_12189,N_12685);
and U13677 (N_13677,N_13063,N_13070);
or U13678 (N_13678,N_12040,N_12236);
nand U13679 (N_13679,N_12095,N_12408);
or U13680 (N_13680,N_12573,N_13078);
and U13681 (N_13681,N_12485,N_13195);
and U13682 (N_13682,N_12545,N_12996);
xnor U13683 (N_13683,N_12254,N_12919);
nor U13684 (N_13684,N_12193,N_12007);
nor U13685 (N_13685,N_12427,N_12909);
nor U13686 (N_13686,N_13027,N_12907);
and U13687 (N_13687,N_12145,N_12951);
nor U13688 (N_13688,N_12418,N_12732);
nand U13689 (N_13689,N_12681,N_13062);
nor U13690 (N_13690,N_12371,N_12644);
nor U13691 (N_13691,N_12332,N_12039);
nor U13692 (N_13692,N_13145,N_12575);
and U13693 (N_13693,N_12131,N_12942);
and U13694 (N_13694,N_12144,N_13157);
or U13695 (N_13695,N_13050,N_12466);
or U13696 (N_13696,N_12625,N_12376);
nor U13697 (N_13697,N_12360,N_12629);
and U13698 (N_13698,N_12527,N_12329);
and U13699 (N_13699,N_12631,N_12321);
xnor U13700 (N_13700,N_12986,N_12969);
or U13701 (N_13701,N_12864,N_12846);
nor U13702 (N_13702,N_12840,N_12096);
xnor U13703 (N_13703,N_12948,N_12375);
nand U13704 (N_13704,N_13184,N_12983);
xnor U13705 (N_13705,N_12135,N_12233);
nor U13706 (N_13706,N_13177,N_12990);
or U13707 (N_13707,N_12744,N_12434);
or U13708 (N_13708,N_13197,N_12475);
xnor U13709 (N_13709,N_13107,N_13000);
and U13710 (N_13710,N_12292,N_12314);
nand U13711 (N_13711,N_12823,N_13118);
xor U13712 (N_13712,N_13034,N_12216);
and U13713 (N_13713,N_12349,N_12227);
nand U13714 (N_13714,N_12424,N_12163);
nand U13715 (N_13715,N_12762,N_12116);
nor U13716 (N_13716,N_12290,N_12082);
nand U13717 (N_13717,N_12294,N_12142);
nor U13718 (N_13718,N_12550,N_12819);
nand U13719 (N_13719,N_12094,N_12950);
and U13720 (N_13720,N_12606,N_12489);
nor U13721 (N_13721,N_13033,N_12979);
nand U13722 (N_13722,N_12363,N_12603);
xnor U13723 (N_13723,N_13133,N_12747);
and U13724 (N_13724,N_12641,N_12670);
and U13725 (N_13725,N_13168,N_12259);
and U13726 (N_13726,N_13018,N_12353);
xor U13727 (N_13727,N_13101,N_12651);
or U13728 (N_13728,N_12214,N_12605);
xor U13729 (N_13729,N_12905,N_12393);
nand U13730 (N_13730,N_12593,N_13125);
or U13731 (N_13731,N_12633,N_12202);
and U13732 (N_13732,N_12881,N_12705);
xor U13733 (N_13733,N_12168,N_12195);
nand U13734 (N_13734,N_12984,N_12484);
or U13735 (N_13735,N_12023,N_12980);
nor U13736 (N_13736,N_12238,N_12663);
xnor U13737 (N_13737,N_12689,N_12859);
nand U13738 (N_13738,N_12392,N_12973);
or U13739 (N_13739,N_12989,N_12931);
nand U13740 (N_13740,N_12402,N_12522);
and U13741 (N_13741,N_13136,N_12861);
and U13742 (N_13742,N_12180,N_13090);
nor U13743 (N_13743,N_12714,N_12635);
nor U13744 (N_13744,N_12335,N_12414);
and U13745 (N_13745,N_12968,N_12956);
nand U13746 (N_13746,N_12612,N_12069);
nand U13747 (N_13747,N_12841,N_12752);
or U13748 (N_13748,N_12472,N_12523);
xor U13749 (N_13749,N_13182,N_12608);
xnor U13750 (N_13750,N_12164,N_13040);
and U13751 (N_13751,N_12652,N_12019);
nor U13752 (N_13752,N_12277,N_12185);
or U13753 (N_13753,N_12058,N_12073);
xnor U13754 (N_13754,N_12955,N_12930);
or U13755 (N_13755,N_12519,N_12997);
or U13756 (N_13756,N_12316,N_12246);
or U13757 (N_13757,N_12825,N_13158);
and U13758 (N_13758,N_12886,N_12843);
nand U13759 (N_13759,N_12949,N_12458);
xor U13760 (N_13760,N_12382,N_13106);
nand U13761 (N_13761,N_13170,N_13180);
and U13762 (N_13762,N_12347,N_12478);
nand U13763 (N_13763,N_12765,N_12339);
or U13764 (N_13764,N_13188,N_12832);
and U13765 (N_13765,N_12786,N_12695);
xnor U13766 (N_13766,N_12559,N_12917);
nand U13767 (N_13767,N_12297,N_13047);
xor U13768 (N_13768,N_12937,N_12634);
nor U13769 (N_13769,N_13010,N_12388);
or U13770 (N_13770,N_12738,N_12413);
and U13771 (N_13771,N_12887,N_12030);
nand U13772 (N_13772,N_12546,N_12583);
or U13773 (N_13773,N_12242,N_12800);
or U13774 (N_13774,N_13160,N_12578);
or U13775 (N_13775,N_12118,N_12721);
or U13776 (N_13776,N_12429,N_12544);
or U13777 (N_13777,N_13057,N_12042);
xnor U13778 (N_13778,N_12270,N_12833);
nor U13779 (N_13779,N_13019,N_12463);
nand U13780 (N_13780,N_12977,N_12943);
xnor U13781 (N_13781,N_12601,N_12922);
or U13782 (N_13782,N_12584,N_12025);
nand U13783 (N_13783,N_13029,N_12411);
or U13784 (N_13784,N_12698,N_12309);
nor U13785 (N_13785,N_12091,N_12251);
or U13786 (N_13786,N_12988,N_12302);
nand U13787 (N_13787,N_12255,N_12755);
and U13788 (N_13788,N_13059,N_12126);
nand U13789 (N_13789,N_12505,N_13075);
nor U13790 (N_13790,N_12659,N_12439);
or U13791 (N_13791,N_12657,N_12203);
xnor U13792 (N_13792,N_12926,N_12993);
or U13793 (N_13793,N_12694,N_12934);
nor U13794 (N_13794,N_12963,N_12693);
nor U13795 (N_13795,N_12647,N_12035);
nor U13796 (N_13796,N_12510,N_12748);
xor U13797 (N_13797,N_12033,N_13036);
nor U13798 (N_13798,N_12240,N_12166);
xor U13799 (N_13799,N_12947,N_12482);
xor U13800 (N_13800,N_12003,N_12038);
or U13801 (N_13801,N_12526,N_12924);
and U13802 (N_13802,N_13030,N_13021);
xnor U13803 (N_13803,N_12222,N_13167);
and U13804 (N_13804,N_12075,N_12190);
nand U13805 (N_13805,N_12721,N_13025);
and U13806 (N_13806,N_12865,N_12600);
xnor U13807 (N_13807,N_12226,N_12969);
nor U13808 (N_13808,N_12560,N_12300);
or U13809 (N_13809,N_12505,N_13099);
and U13810 (N_13810,N_12755,N_12524);
and U13811 (N_13811,N_12597,N_12889);
or U13812 (N_13812,N_12806,N_12327);
and U13813 (N_13813,N_12773,N_12529);
nor U13814 (N_13814,N_12680,N_12140);
nor U13815 (N_13815,N_12054,N_12395);
nor U13816 (N_13816,N_12769,N_12857);
or U13817 (N_13817,N_12172,N_12870);
xnor U13818 (N_13818,N_12126,N_12855);
and U13819 (N_13819,N_12146,N_12649);
nor U13820 (N_13820,N_12207,N_12786);
nand U13821 (N_13821,N_12688,N_12895);
and U13822 (N_13822,N_12257,N_12044);
or U13823 (N_13823,N_12807,N_12791);
and U13824 (N_13824,N_13191,N_12926);
nand U13825 (N_13825,N_12824,N_13060);
xnor U13826 (N_13826,N_13090,N_12609);
xor U13827 (N_13827,N_12395,N_12079);
xor U13828 (N_13828,N_13163,N_12275);
xor U13829 (N_13829,N_12534,N_12974);
and U13830 (N_13830,N_12980,N_12658);
and U13831 (N_13831,N_13090,N_12412);
nor U13832 (N_13832,N_12576,N_12254);
nor U13833 (N_13833,N_12652,N_12570);
xnor U13834 (N_13834,N_12659,N_13030);
nor U13835 (N_13835,N_12006,N_12089);
and U13836 (N_13836,N_12964,N_12266);
or U13837 (N_13837,N_12858,N_12996);
nand U13838 (N_13838,N_12325,N_12003);
or U13839 (N_13839,N_12452,N_12733);
and U13840 (N_13840,N_12469,N_12100);
xnor U13841 (N_13841,N_12648,N_12151);
or U13842 (N_13842,N_12847,N_12428);
or U13843 (N_13843,N_12633,N_12233);
xor U13844 (N_13844,N_12352,N_12632);
nor U13845 (N_13845,N_12679,N_13144);
nor U13846 (N_13846,N_12640,N_12391);
and U13847 (N_13847,N_12107,N_12495);
xor U13848 (N_13848,N_12104,N_12801);
nor U13849 (N_13849,N_12017,N_12874);
nand U13850 (N_13850,N_12586,N_12597);
xnor U13851 (N_13851,N_12709,N_12919);
nand U13852 (N_13852,N_12226,N_12837);
or U13853 (N_13853,N_12343,N_12735);
nand U13854 (N_13854,N_12110,N_13011);
or U13855 (N_13855,N_12042,N_12774);
and U13856 (N_13856,N_12930,N_12386);
and U13857 (N_13857,N_12074,N_12734);
or U13858 (N_13858,N_13151,N_12347);
and U13859 (N_13859,N_13127,N_12648);
nor U13860 (N_13860,N_12841,N_12693);
nand U13861 (N_13861,N_12442,N_12236);
and U13862 (N_13862,N_12515,N_12309);
and U13863 (N_13863,N_12986,N_12996);
xor U13864 (N_13864,N_12252,N_13021);
or U13865 (N_13865,N_12305,N_12807);
xnor U13866 (N_13866,N_13161,N_12764);
xor U13867 (N_13867,N_13043,N_12542);
and U13868 (N_13868,N_12197,N_13074);
and U13869 (N_13869,N_12894,N_12909);
nor U13870 (N_13870,N_12213,N_12811);
nand U13871 (N_13871,N_12445,N_12015);
and U13872 (N_13872,N_12406,N_13088);
xor U13873 (N_13873,N_13115,N_12994);
nor U13874 (N_13874,N_13183,N_13121);
xnor U13875 (N_13875,N_12017,N_12417);
nand U13876 (N_13876,N_12397,N_12572);
nor U13877 (N_13877,N_12677,N_13125);
nor U13878 (N_13878,N_12848,N_12677);
nand U13879 (N_13879,N_12736,N_12157);
or U13880 (N_13880,N_12605,N_12246);
and U13881 (N_13881,N_12444,N_12087);
nor U13882 (N_13882,N_12250,N_12154);
xnor U13883 (N_13883,N_12284,N_12850);
and U13884 (N_13884,N_13140,N_12922);
or U13885 (N_13885,N_12884,N_13036);
nand U13886 (N_13886,N_13087,N_12394);
nor U13887 (N_13887,N_13168,N_12171);
and U13888 (N_13888,N_12735,N_12412);
and U13889 (N_13889,N_12627,N_13115);
nor U13890 (N_13890,N_12828,N_12829);
and U13891 (N_13891,N_12205,N_12291);
nor U13892 (N_13892,N_12186,N_12525);
or U13893 (N_13893,N_12279,N_12320);
nand U13894 (N_13894,N_12011,N_12906);
and U13895 (N_13895,N_12673,N_12481);
and U13896 (N_13896,N_12617,N_12273);
or U13897 (N_13897,N_12442,N_12420);
nand U13898 (N_13898,N_12157,N_12236);
nand U13899 (N_13899,N_13023,N_12791);
and U13900 (N_13900,N_12168,N_12072);
nor U13901 (N_13901,N_12058,N_12872);
nand U13902 (N_13902,N_12425,N_13097);
nand U13903 (N_13903,N_12183,N_13055);
xnor U13904 (N_13904,N_13101,N_13111);
and U13905 (N_13905,N_12289,N_12097);
xnor U13906 (N_13906,N_12822,N_12364);
nor U13907 (N_13907,N_13035,N_12969);
and U13908 (N_13908,N_12296,N_13080);
nor U13909 (N_13909,N_12527,N_12554);
and U13910 (N_13910,N_12546,N_12140);
or U13911 (N_13911,N_12938,N_12824);
nand U13912 (N_13912,N_12819,N_12917);
or U13913 (N_13913,N_13054,N_12414);
nor U13914 (N_13914,N_12169,N_12374);
xnor U13915 (N_13915,N_12717,N_12291);
xor U13916 (N_13916,N_12974,N_12268);
or U13917 (N_13917,N_12079,N_12127);
or U13918 (N_13918,N_13104,N_12946);
or U13919 (N_13919,N_12401,N_12975);
xnor U13920 (N_13920,N_12698,N_12767);
nor U13921 (N_13921,N_13165,N_12738);
xnor U13922 (N_13922,N_12066,N_12997);
or U13923 (N_13923,N_12761,N_12619);
xnor U13924 (N_13924,N_12660,N_13167);
nand U13925 (N_13925,N_12563,N_12477);
nand U13926 (N_13926,N_12921,N_13068);
xnor U13927 (N_13927,N_12202,N_12589);
nor U13928 (N_13928,N_12154,N_12531);
xnor U13929 (N_13929,N_12202,N_12713);
xor U13930 (N_13930,N_12806,N_13105);
and U13931 (N_13931,N_13118,N_12277);
nor U13932 (N_13932,N_12424,N_13049);
nand U13933 (N_13933,N_12575,N_12023);
nor U13934 (N_13934,N_13169,N_12545);
xnor U13935 (N_13935,N_12791,N_13037);
xor U13936 (N_13936,N_12264,N_12273);
nor U13937 (N_13937,N_13052,N_12865);
and U13938 (N_13938,N_12068,N_12086);
xor U13939 (N_13939,N_12481,N_12463);
nand U13940 (N_13940,N_12644,N_12806);
nand U13941 (N_13941,N_12299,N_12747);
nand U13942 (N_13942,N_12341,N_13124);
nor U13943 (N_13943,N_12922,N_12554);
or U13944 (N_13944,N_12994,N_12915);
nand U13945 (N_13945,N_12061,N_12815);
and U13946 (N_13946,N_12812,N_12902);
nand U13947 (N_13947,N_13051,N_12023);
nand U13948 (N_13948,N_12929,N_13004);
nand U13949 (N_13949,N_12537,N_12363);
and U13950 (N_13950,N_12577,N_12591);
nor U13951 (N_13951,N_13120,N_12822);
nand U13952 (N_13952,N_13118,N_12111);
nand U13953 (N_13953,N_12374,N_12062);
or U13954 (N_13954,N_12666,N_13091);
nor U13955 (N_13955,N_12080,N_13175);
and U13956 (N_13956,N_12096,N_12776);
or U13957 (N_13957,N_12784,N_12009);
and U13958 (N_13958,N_12597,N_13087);
and U13959 (N_13959,N_12837,N_12745);
nand U13960 (N_13960,N_12830,N_12964);
nand U13961 (N_13961,N_12074,N_12763);
xnor U13962 (N_13962,N_12732,N_12079);
nor U13963 (N_13963,N_12076,N_12441);
nor U13964 (N_13964,N_12298,N_12587);
and U13965 (N_13965,N_12103,N_13012);
nand U13966 (N_13966,N_12396,N_12616);
or U13967 (N_13967,N_12509,N_12695);
or U13968 (N_13968,N_12968,N_13013);
nand U13969 (N_13969,N_13019,N_12716);
nor U13970 (N_13970,N_13170,N_12874);
xor U13971 (N_13971,N_12550,N_12731);
nor U13972 (N_13972,N_12320,N_12241);
and U13973 (N_13973,N_12773,N_12210);
and U13974 (N_13974,N_12836,N_12925);
nor U13975 (N_13975,N_12723,N_12339);
and U13976 (N_13976,N_12970,N_12760);
and U13977 (N_13977,N_12400,N_12800);
xnor U13978 (N_13978,N_12171,N_13075);
nor U13979 (N_13979,N_13018,N_12019);
and U13980 (N_13980,N_13004,N_12619);
nor U13981 (N_13981,N_12072,N_12613);
and U13982 (N_13982,N_13165,N_13109);
nor U13983 (N_13983,N_12474,N_12406);
nor U13984 (N_13984,N_12681,N_12508);
nand U13985 (N_13985,N_13155,N_12858);
nand U13986 (N_13986,N_12342,N_12898);
or U13987 (N_13987,N_12308,N_12549);
or U13988 (N_13988,N_12171,N_12060);
or U13989 (N_13989,N_12554,N_13197);
and U13990 (N_13990,N_12637,N_12819);
and U13991 (N_13991,N_12638,N_12138);
xor U13992 (N_13992,N_12792,N_12026);
and U13993 (N_13993,N_12979,N_12949);
xor U13994 (N_13994,N_12798,N_12473);
xnor U13995 (N_13995,N_12795,N_12250);
or U13996 (N_13996,N_12313,N_12976);
nor U13997 (N_13997,N_12681,N_12465);
nor U13998 (N_13998,N_12626,N_12544);
and U13999 (N_13999,N_12420,N_12035);
xnor U14000 (N_14000,N_12653,N_13032);
or U14001 (N_14001,N_12510,N_13173);
and U14002 (N_14002,N_12940,N_13010);
or U14003 (N_14003,N_12401,N_13135);
or U14004 (N_14004,N_12268,N_12914);
and U14005 (N_14005,N_13088,N_12848);
or U14006 (N_14006,N_12814,N_12972);
xnor U14007 (N_14007,N_12397,N_13135);
nand U14008 (N_14008,N_12589,N_12939);
nand U14009 (N_14009,N_12567,N_13007);
nor U14010 (N_14010,N_13081,N_12072);
or U14011 (N_14011,N_12416,N_12094);
and U14012 (N_14012,N_12706,N_12315);
xnor U14013 (N_14013,N_13091,N_12847);
and U14014 (N_14014,N_12774,N_13032);
nand U14015 (N_14015,N_12476,N_12347);
xor U14016 (N_14016,N_12577,N_12659);
and U14017 (N_14017,N_12012,N_12089);
nor U14018 (N_14018,N_13151,N_12724);
nor U14019 (N_14019,N_12257,N_12228);
and U14020 (N_14020,N_13158,N_12872);
nand U14021 (N_14021,N_12739,N_12698);
nand U14022 (N_14022,N_12946,N_12950);
and U14023 (N_14023,N_12466,N_12409);
nand U14024 (N_14024,N_12209,N_12960);
nand U14025 (N_14025,N_13155,N_12188);
and U14026 (N_14026,N_12313,N_13075);
nor U14027 (N_14027,N_13127,N_12673);
or U14028 (N_14028,N_12399,N_12557);
or U14029 (N_14029,N_13018,N_12862);
xnor U14030 (N_14030,N_12347,N_12607);
or U14031 (N_14031,N_13000,N_12943);
and U14032 (N_14032,N_13115,N_12744);
nor U14033 (N_14033,N_12535,N_12098);
xor U14034 (N_14034,N_12230,N_12032);
nor U14035 (N_14035,N_12237,N_12939);
xor U14036 (N_14036,N_12708,N_12054);
and U14037 (N_14037,N_12478,N_12333);
nor U14038 (N_14038,N_12740,N_12803);
nor U14039 (N_14039,N_12344,N_12368);
nor U14040 (N_14040,N_12207,N_12516);
nor U14041 (N_14041,N_12837,N_12427);
or U14042 (N_14042,N_13139,N_12505);
or U14043 (N_14043,N_12721,N_12400);
or U14044 (N_14044,N_12814,N_12675);
nor U14045 (N_14045,N_13043,N_12947);
and U14046 (N_14046,N_12575,N_12064);
nor U14047 (N_14047,N_12820,N_12056);
or U14048 (N_14048,N_12183,N_12101);
or U14049 (N_14049,N_12765,N_12451);
nand U14050 (N_14050,N_12699,N_12941);
and U14051 (N_14051,N_13116,N_12255);
nand U14052 (N_14052,N_12129,N_13121);
nand U14053 (N_14053,N_12323,N_12275);
nand U14054 (N_14054,N_12726,N_12143);
nor U14055 (N_14055,N_12082,N_12639);
nand U14056 (N_14056,N_12749,N_13131);
nand U14057 (N_14057,N_12742,N_12487);
nor U14058 (N_14058,N_12558,N_12493);
nor U14059 (N_14059,N_12229,N_12488);
nor U14060 (N_14060,N_12797,N_12937);
nand U14061 (N_14061,N_12948,N_12572);
nor U14062 (N_14062,N_12698,N_12237);
and U14063 (N_14063,N_12164,N_12786);
and U14064 (N_14064,N_12440,N_12554);
nor U14065 (N_14065,N_12949,N_12825);
or U14066 (N_14066,N_12740,N_12841);
nor U14067 (N_14067,N_12090,N_12969);
xor U14068 (N_14068,N_12704,N_12526);
and U14069 (N_14069,N_13123,N_13051);
nand U14070 (N_14070,N_13046,N_12376);
nand U14071 (N_14071,N_12259,N_13054);
nor U14072 (N_14072,N_12541,N_12273);
and U14073 (N_14073,N_12985,N_12647);
and U14074 (N_14074,N_13079,N_12563);
nor U14075 (N_14075,N_12638,N_12408);
nor U14076 (N_14076,N_12950,N_12716);
or U14077 (N_14077,N_12914,N_12789);
and U14078 (N_14078,N_12191,N_12985);
xnor U14079 (N_14079,N_12876,N_13128);
and U14080 (N_14080,N_12146,N_12686);
xnor U14081 (N_14081,N_12314,N_12470);
or U14082 (N_14082,N_12051,N_12418);
nand U14083 (N_14083,N_13138,N_13159);
or U14084 (N_14084,N_12786,N_13069);
or U14085 (N_14085,N_12698,N_12748);
xor U14086 (N_14086,N_12384,N_12888);
nor U14087 (N_14087,N_12829,N_12236);
and U14088 (N_14088,N_13089,N_12459);
and U14089 (N_14089,N_12100,N_12636);
and U14090 (N_14090,N_12827,N_12198);
nor U14091 (N_14091,N_12615,N_13003);
and U14092 (N_14092,N_12255,N_12832);
and U14093 (N_14093,N_12525,N_12757);
nand U14094 (N_14094,N_12747,N_12077);
or U14095 (N_14095,N_12864,N_12651);
nor U14096 (N_14096,N_12577,N_13110);
nor U14097 (N_14097,N_12652,N_12332);
nand U14098 (N_14098,N_12078,N_12613);
nand U14099 (N_14099,N_12972,N_12633);
nand U14100 (N_14100,N_13123,N_13034);
nor U14101 (N_14101,N_12936,N_12556);
nand U14102 (N_14102,N_13055,N_12793);
and U14103 (N_14103,N_13138,N_12866);
xor U14104 (N_14104,N_12177,N_12012);
and U14105 (N_14105,N_12288,N_12952);
xnor U14106 (N_14106,N_13085,N_12949);
xor U14107 (N_14107,N_13150,N_12520);
or U14108 (N_14108,N_12352,N_12273);
nor U14109 (N_14109,N_12737,N_12651);
nor U14110 (N_14110,N_12509,N_13152);
nand U14111 (N_14111,N_13116,N_12797);
or U14112 (N_14112,N_12945,N_12576);
and U14113 (N_14113,N_13103,N_13101);
or U14114 (N_14114,N_12007,N_12706);
nor U14115 (N_14115,N_12268,N_12023);
and U14116 (N_14116,N_12920,N_12413);
or U14117 (N_14117,N_12764,N_12404);
nor U14118 (N_14118,N_12290,N_12288);
and U14119 (N_14119,N_12200,N_12083);
or U14120 (N_14120,N_12421,N_13154);
xnor U14121 (N_14121,N_12060,N_12411);
and U14122 (N_14122,N_12638,N_12547);
xnor U14123 (N_14123,N_12079,N_12830);
and U14124 (N_14124,N_12544,N_12578);
and U14125 (N_14125,N_12962,N_12077);
xor U14126 (N_14126,N_12355,N_12201);
nand U14127 (N_14127,N_12110,N_13095);
or U14128 (N_14128,N_12445,N_12535);
nand U14129 (N_14129,N_13053,N_12698);
nand U14130 (N_14130,N_12097,N_12320);
and U14131 (N_14131,N_12220,N_13094);
or U14132 (N_14132,N_12471,N_12570);
or U14133 (N_14133,N_12132,N_12449);
and U14134 (N_14134,N_12975,N_12818);
nor U14135 (N_14135,N_12168,N_12356);
and U14136 (N_14136,N_12428,N_12028);
and U14137 (N_14137,N_13024,N_12239);
or U14138 (N_14138,N_13111,N_12515);
and U14139 (N_14139,N_13035,N_12241);
nor U14140 (N_14140,N_13045,N_12251);
or U14141 (N_14141,N_12047,N_12538);
nand U14142 (N_14142,N_12765,N_12264);
or U14143 (N_14143,N_12927,N_12042);
xor U14144 (N_14144,N_12698,N_12621);
nand U14145 (N_14145,N_12625,N_12338);
nand U14146 (N_14146,N_13170,N_13064);
or U14147 (N_14147,N_12620,N_12090);
xor U14148 (N_14148,N_12471,N_12430);
xor U14149 (N_14149,N_12403,N_12884);
or U14150 (N_14150,N_12793,N_12423);
or U14151 (N_14151,N_12802,N_13077);
nor U14152 (N_14152,N_13123,N_12763);
xor U14153 (N_14153,N_12836,N_12229);
nand U14154 (N_14154,N_12104,N_12726);
xnor U14155 (N_14155,N_13190,N_12475);
xor U14156 (N_14156,N_13182,N_12595);
xnor U14157 (N_14157,N_12339,N_12630);
xor U14158 (N_14158,N_12211,N_13041);
nand U14159 (N_14159,N_12091,N_12952);
xnor U14160 (N_14160,N_12987,N_12100);
and U14161 (N_14161,N_12909,N_12063);
or U14162 (N_14162,N_12376,N_12599);
nand U14163 (N_14163,N_12433,N_12208);
or U14164 (N_14164,N_12321,N_12850);
and U14165 (N_14165,N_13188,N_12029);
nand U14166 (N_14166,N_12691,N_12215);
nand U14167 (N_14167,N_13191,N_12389);
nor U14168 (N_14168,N_13085,N_12556);
nor U14169 (N_14169,N_12352,N_13154);
and U14170 (N_14170,N_12911,N_12368);
or U14171 (N_14171,N_13047,N_12663);
or U14172 (N_14172,N_12580,N_12859);
and U14173 (N_14173,N_12078,N_12634);
nand U14174 (N_14174,N_12996,N_12478);
or U14175 (N_14175,N_13198,N_12982);
or U14176 (N_14176,N_13139,N_12682);
or U14177 (N_14177,N_12705,N_12457);
and U14178 (N_14178,N_12548,N_12793);
or U14179 (N_14179,N_12412,N_12464);
nand U14180 (N_14180,N_12569,N_12628);
xor U14181 (N_14181,N_12601,N_12655);
or U14182 (N_14182,N_12072,N_12167);
and U14183 (N_14183,N_13170,N_12332);
and U14184 (N_14184,N_13100,N_12778);
or U14185 (N_14185,N_12189,N_12240);
nor U14186 (N_14186,N_13011,N_12851);
and U14187 (N_14187,N_12364,N_12249);
nor U14188 (N_14188,N_12926,N_13193);
or U14189 (N_14189,N_12975,N_13191);
or U14190 (N_14190,N_12201,N_13002);
or U14191 (N_14191,N_12502,N_12799);
nor U14192 (N_14192,N_13007,N_12438);
nor U14193 (N_14193,N_12879,N_12025);
nor U14194 (N_14194,N_12540,N_13068);
or U14195 (N_14195,N_12820,N_12851);
and U14196 (N_14196,N_12021,N_12315);
nor U14197 (N_14197,N_12786,N_12287);
nor U14198 (N_14198,N_13178,N_13030);
nor U14199 (N_14199,N_13169,N_12365);
and U14200 (N_14200,N_12940,N_12360);
xor U14201 (N_14201,N_12308,N_13180);
nor U14202 (N_14202,N_13102,N_12904);
nor U14203 (N_14203,N_12902,N_12954);
nor U14204 (N_14204,N_12604,N_12798);
or U14205 (N_14205,N_12469,N_12315);
xor U14206 (N_14206,N_12304,N_12586);
nand U14207 (N_14207,N_12608,N_12926);
and U14208 (N_14208,N_12018,N_12862);
nand U14209 (N_14209,N_12619,N_12319);
nor U14210 (N_14210,N_12644,N_13184);
or U14211 (N_14211,N_12196,N_12193);
or U14212 (N_14212,N_12721,N_12540);
or U14213 (N_14213,N_12119,N_12788);
nand U14214 (N_14214,N_12207,N_12998);
xor U14215 (N_14215,N_12864,N_13130);
or U14216 (N_14216,N_12731,N_12777);
nand U14217 (N_14217,N_12246,N_12503);
and U14218 (N_14218,N_12150,N_12328);
and U14219 (N_14219,N_12864,N_13137);
xnor U14220 (N_14220,N_12680,N_12221);
or U14221 (N_14221,N_13101,N_12683);
and U14222 (N_14222,N_12892,N_12305);
or U14223 (N_14223,N_12017,N_13064);
or U14224 (N_14224,N_12729,N_12159);
nor U14225 (N_14225,N_12576,N_12829);
xnor U14226 (N_14226,N_12269,N_12439);
or U14227 (N_14227,N_12454,N_12912);
or U14228 (N_14228,N_12000,N_12979);
and U14229 (N_14229,N_12757,N_12484);
and U14230 (N_14230,N_12699,N_12208);
and U14231 (N_14231,N_12255,N_12691);
xor U14232 (N_14232,N_12264,N_12229);
xor U14233 (N_14233,N_13113,N_12113);
xor U14234 (N_14234,N_12181,N_12548);
nand U14235 (N_14235,N_13131,N_12394);
or U14236 (N_14236,N_12170,N_12156);
and U14237 (N_14237,N_13057,N_12822);
and U14238 (N_14238,N_12921,N_12772);
xor U14239 (N_14239,N_13108,N_12461);
and U14240 (N_14240,N_12719,N_12374);
and U14241 (N_14241,N_12917,N_12384);
nand U14242 (N_14242,N_12284,N_13170);
nor U14243 (N_14243,N_12269,N_12349);
xor U14244 (N_14244,N_12192,N_12864);
nand U14245 (N_14245,N_12365,N_12204);
nand U14246 (N_14246,N_12666,N_12708);
nor U14247 (N_14247,N_12150,N_12392);
or U14248 (N_14248,N_12686,N_12331);
or U14249 (N_14249,N_12210,N_13066);
xnor U14250 (N_14250,N_12256,N_12043);
nand U14251 (N_14251,N_12225,N_13022);
xor U14252 (N_14252,N_12360,N_12992);
or U14253 (N_14253,N_12816,N_12624);
nor U14254 (N_14254,N_12887,N_12534);
nand U14255 (N_14255,N_13087,N_12791);
nor U14256 (N_14256,N_12132,N_12907);
and U14257 (N_14257,N_12954,N_12635);
nor U14258 (N_14258,N_12643,N_13050);
or U14259 (N_14259,N_12167,N_13049);
nor U14260 (N_14260,N_12311,N_12342);
xnor U14261 (N_14261,N_12958,N_12204);
xor U14262 (N_14262,N_12749,N_13118);
or U14263 (N_14263,N_13186,N_12392);
nand U14264 (N_14264,N_12572,N_12636);
nand U14265 (N_14265,N_12598,N_12943);
nor U14266 (N_14266,N_12162,N_13002);
xor U14267 (N_14267,N_12776,N_12729);
nor U14268 (N_14268,N_12512,N_12540);
or U14269 (N_14269,N_12317,N_12438);
xor U14270 (N_14270,N_12867,N_12864);
and U14271 (N_14271,N_12378,N_12929);
nand U14272 (N_14272,N_12156,N_12941);
or U14273 (N_14273,N_12540,N_12863);
xnor U14274 (N_14274,N_12547,N_12672);
xnor U14275 (N_14275,N_13078,N_13155);
and U14276 (N_14276,N_12092,N_12393);
xor U14277 (N_14277,N_12205,N_12081);
nand U14278 (N_14278,N_12269,N_12617);
xor U14279 (N_14279,N_12490,N_13035);
nor U14280 (N_14280,N_12400,N_12843);
nand U14281 (N_14281,N_12998,N_12769);
nor U14282 (N_14282,N_12346,N_12997);
nor U14283 (N_14283,N_12531,N_13198);
and U14284 (N_14284,N_12170,N_13122);
or U14285 (N_14285,N_12139,N_12681);
or U14286 (N_14286,N_12703,N_12646);
nand U14287 (N_14287,N_12204,N_12879);
nand U14288 (N_14288,N_12275,N_12208);
xor U14289 (N_14289,N_12414,N_12916);
or U14290 (N_14290,N_13100,N_12525);
nor U14291 (N_14291,N_12018,N_12040);
or U14292 (N_14292,N_12374,N_12644);
or U14293 (N_14293,N_12307,N_13028);
nor U14294 (N_14294,N_12234,N_13036);
and U14295 (N_14295,N_12729,N_12921);
or U14296 (N_14296,N_12464,N_12114);
nor U14297 (N_14297,N_12540,N_12501);
nand U14298 (N_14298,N_12239,N_12639);
nor U14299 (N_14299,N_12067,N_12383);
nand U14300 (N_14300,N_13150,N_12433);
xor U14301 (N_14301,N_12168,N_12769);
or U14302 (N_14302,N_12155,N_12348);
or U14303 (N_14303,N_12135,N_12838);
nor U14304 (N_14304,N_12192,N_12803);
and U14305 (N_14305,N_12333,N_12641);
xnor U14306 (N_14306,N_12184,N_12559);
xor U14307 (N_14307,N_12937,N_12359);
nand U14308 (N_14308,N_13004,N_12469);
xnor U14309 (N_14309,N_12600,N_13170);
xnor U14310 (N_14310,N_12864,N_13006);
xor U14311 (N_14311,N_13161,N_12279);
or U14312 (N_14312,N_12555,N_12626);
and U14313 (N_14313,N_12191,N_12717);
nor U14314 (N_14314,N_12881,N_12220);
nand U14315 (N_14315,N_12135,N_12417);
xor U14316 (N_14316,N_12275,N_12244);
nor U14317 (N_14317,N_12536,N_13102);
or U14318 (N_14318,N_12714,N_12254);
nor U14319 (N_14319,N_12961,N_12569);
or U14320 (N_14320,N_13007,N_12877);
xnor U14321 (N_14321,N_12110,N_13124);
and U14322 (N_14322,N_12193,N_12232);
nand U14323 (N_14323,N_12912,N_12594);
or U14324 (N_14324,N_12802,N_12644);
nor U14325 (N_14325,N_12786,N_12660);
and U14326 (N_14326,N_12411,N_12504);
and U14327 (N_14327,N_12562,N_13064);
nand U14328 (N_14328,N_12941,N_12275);
nor U14329 (N_14329,N_12789,N_12356);
nor U14330 (N_14330,N_12383,N_13087);
and U14331 (N_14331,N_12646,N_12325);
nor U14332 (N_14332,N_12777,N_12350);
and U14333 (N_14333,N_12037,N_12833);
nor U14334 (N_14334,N_12243,N_12965);
nand U14335 (N_14335,N_12185,N_12414);
or U14336 (N_14336,N_12865,N_12449);
nand U14337 (N_14337,N_12445,N_12243);
and U14338 (N_14338,N_13111,N_12003);
and U14339 (N_14339,N_12189,N_12361);
and U14340 (N_14340,N_12979,N_12619);
and U14341 (N_14341,N_13122,N_13119);
xnor U14342 (N_14342,N_12496,N_12977);
nor U14343 (N_14343,N_13064,N_12214);
and U14344 (N_14344,N_13058,N_12712);
and U14345 (N_14345,N_12771,N_12877);
and U14346 (N_14346,N_12245,N_12333);
xnor U14347 (N_14347,N_13044,N_12688);
nand U14348 (N_14348,N_12526,N_12511);
and U14349 (N_14349,N_12514,N_13197);
nor U14350 (N_14350,N_12829,N_12638);
xor U14351 (N_14351,N_12263,N_12742);
or U14352 (N_14352,N_12617,N_12531);
xor U14353 (N_14353,N_13195,N_12307);
or U14354 (N_14354,N_12122,N_12438);
nand U14355 (N_14355,N_12352,N_12969);
or U14356 (N_14356,N_13018,N_12892);
and U14357 (N_14357,N_13130,N_12562);
nor U14358 (N_14358,N_12846,N_12493);
nor U14359 (N_14359,N_12888,N_12228);
and U14360 (N_14360,N_12923,N_12199);
or U14361 (N_14361,N_12582,N_12141);
or U14362 (N_14362,N_12922,N_12515);
nor U14363 (N_14363,N_12943,N_12299);
or U14364 (N_14364,N_13067,N_13120);
or U14365 (N_14365,N_12947,N_13193);
and U14366 (N_14366,N_12064,N_12872);
or U14367 (N_14367,N_12474,N_12546);
or U14368 (N_14368,N_12153,N_12233);
or U14369 (N_14369,N_12337,N_12245);
xnor U14370 (N_14370,N_12472,N_12919);
nand U14371 (N_14371,N_12252,N_12216);
and U14372 (N_14372,N_12738,N_12895);
or U14373 (N_14373,N_12789,N_12975);
or U14374 (N_14374,N_13023,N_13085);
nor U14375 (N_14375,N_13167,N_12319);
or U14376 (N_14376,N_12661,N_12248);
xor U14377 (N_14377,N_13037,N_12196);
nand U14378 (N_14378,N_12951,N_12365);
nand U14379 (N_14379,N_12414,N_12886);
xnor U14380 (N_14380,N_12895,N_12505);
nor U14381 (N_14381,N_12486,N_13007);
nor U14382 (N_14382,N_13147,N_12470);
xor U14383 (N_14383,N_12054,N_12985);
and U14384 (N_14384,N_13168,N_12675);
and U14385 (N_14385,N_12919,N_12747);
and U14386 (N_14386,N_12752,N_12929);
or U14387 (N_14387,N_13151,N_12127);
nand U14388 (N_14388,N_12186,N_12201);
or U14389 (N_14389,N_12124,N_13156);
or U14390 (N_14390,N_13152,N_13134);
xor U14391 (N_14391,N_12953,N_12951);
xor U14392 (N_14392,N_12463,N_12920);
nor U14393 (N_14393,N_12203,N_13098);
xnor U14394 (N_14394,N_12797,N_12204);
and U14395 (N_14395,N_12454,N_12325);
xor U14396 (N_14396,N_12760,N_13069);
or U14397 (N_14397,N_12931,N_12147);
xnor U14398 (N_14398,N_12059,N_12390);
xor U14399 (N_14399,N_12089,N_13083);
nor U14400 (N_14400,N_13371,N_13458);
xnor U14401 (N_14401,N_13966,N_13226);
or U14402 (N_14402,N_13473,N_14283);
nor U14403 (N_14403,N_13322,N_14094);
or U14404 (N_14404,N_14046,N_14083);
nand U14405 (N_14405,N_13965,N_13265);
nand U14406 (N_14406,N_13994,N_13868);
nand U14407 (N_14407,N_13310,N_14114);
or U14408 (N_14408,N_13350,N_14330);
or U14409 (N_14409,N_13843,N_14150);
or U14410 (N_14410,N_14235,N_14021);
and U14411 (N_14411,N_13715,N_14204);
and U14412 (N_14412,N_13943,N_14014);
nor U14413 (N_14413,N_14143,N_14101);
nand U14414 (N_14414,N_13910,N_14389);
nor U14415 (N_14415,N_14091,N_13789);
or U14416 (N_14416,N_13945,N_13738);
and U14417 (N_14417,N_13316,N_14023);
and U14418 (N_14418,N_14369,N_13591);
or U14419 (N_14419,N_13555,N_13233);
or U14420 (N_14420,N_14220,N_13589);
nand U14421 (N_14421,N_13321,N_14076);
xor U14422 (N_14422,N_13225,N_14266);
xor U14423 (N_14423,N_13202,N_13342);
and U14424 (N_14424,N_14261,N_13506);
xnor U14425 (N_14425,N_13681,N_13696);
nand U14426 (N_14426,N_14335,N_13973);
nor U14427 (N_14427,N_13949,N_13934);
nand U14428 (N_14428,N_14270,N_14038);
or U14429 (N_14429,N_13730,N_13406);
nor U14430 (N_14430,N_14146,N_13753);
nor U14431 (N_14431,N_14297,N_13381);
and U14432 (N_14432,N_13499,N_13706);
or U14433 (N_14433,N_13273,N_13338);
nand U14434 (N_14434,N_14151,N_14368);
nand U14435 (N_14435,N_13243,N_13262);
or U14436 (N_14436,N_13391,N_14182);
xnor U14437 (N_14437,N_13411,N_14218);
xnor U14438 (N_14438,N_13514,N_14184);
or U14439 (N_14439,N_14349,N_13883);
or U14440 (N_14440,N_13685,N_14118);
xor U14441 (N_14441,N_13729,N_14319);
xnor U14442 (N_14442,N_14117,N_13800);
nor U14443 (N_14443,N_13324,N_13556);
or U14444 (N_14444,N_13305,N_14345);
nor U14445 (N_14445,N_13308,N_14234);
nor U14446 (N_14446,N_13891,N_14308);
nor U14447 (N_14447,N_14274,N_13732);
or U14448 (N_14448,N_13951,N_13505);
or U14449 (N_14449,N_13817,N_13278);
xor U14450 (N_14450,N_13645,N_14060);
nand U14451 (N_14451,N_13410,N_14269);
nand U14452 (N_14452,N_13213,N_14122);
nand U14453 (N_14453,N_13769,N_13529);
xor U14454 (N_14454,N_14065,N_14115);
xor U14455 (N_14455,N_13660,N_14129);
xor U14456 (N_14456,N_13489,N_14306);
nor U14457 (N_14457,N_13720,N_14179);
nor U14458 (N_14458,N_14396,N_13621);
and U14459 (N_14459,N_13286,N_13630);
or U14460 (N_14460,N_13852,N_13849);
xor U14461 (N_14461,N_13758,N_13520);
and U14462 (N_14462,N_14121,N_13954);
or U14463 (N_14463,N_13357,N_13527);
nand U14464 (N_14464,N_13221,N_14217);
and U14465 (N_14465,N_13483,N_13404);
and U14466 (N_14466,N_13393,N_14350);
and U14467 (N_14467,N_13407,N_13533);
or U14468 (N_14468,N_13811,N_13770);
or U14469 (N_14469,N_13318,N_14099);
nor U14470 (N_14470,N_14289,N_14207);
nor U14471 (N_14471,N_13797,N_13628);
and U14472 (N_14472,N_13613,N_13959);
nor U14473 (N_14473,N_13932,N_13263);
xnor U14474 (N_14474,N_14035,N_13384);
nand U14475 (N_14475,N_14252,N_14176);
nand U14476 (N_14476,N_13232,N_13260);
and U14477 (N_14477,N_14189,N_13633);
and U14478 (N_14478,N_13481,N_13281);
xnor U14479 (N_14479,N_14028,N_13616);
and U14480 (N_14480,N_14267,N_13986);
xnor U14481 (N_14481,N_14079,N_13500);
or U14482 (N_14482,N_14344,N_13756);
nor U14483 (N_14483,N_13869,N_13256);
xor U14484 (N_14484,N_13953,N_13284);
nand U14485 (N_14485,N_13831,N_13415);
and U14486 (N_14486,N_14359,N_13474);
nor U14487 (N_14487,N_14026,N_13223);
nor U14488 (N_14488,N_14001,N_13676);
nor U14489 (N_14489,N_13542,N_13351);
xor U14490 (N_14490,N_13475,N_13352);
or U14491 (N_14491,N_14087,N_13921);
xnor U14492 (N_14492,N_14363,N_13703);
or U14493 (N_14493,N_13752,N_14066);
and U14494 (N_14494,N_13331,N_14120);
or U14495 (N_14495,N_13295,N_13689);
or U14496 (N_14496,N_13925,N_13445);
nor U14497 (N_14497,N_13477,N_14342);
nand U14498 (N_14498,N_14320,N_13740);
nor U14499 (N_14499,N_14136,N_13508);
nand U14500 (N_14500,N_14047,N_13801);
and U14501 (N_14501,N_14242,N_13772);
nor U14502 (N_14502,N_14196,N_14382);
or U14503 (N_14503,N_13437,N_13942);
nand U14504 (N_14504,N_14109,N_13725);
or U14505 (N_14505,N_13240,N_13261);
or U14506 (N_14506,N_13999,N_14003);
xnor U14507 (N_14507,N_13599,N_14107);
and U14508 (N_14508,N_13258,N_13736);
nand U14509 (N_14509,N_13767,N_13625);
xor U14510 (N_14510,N_13960,N_14338);
nand U14511 (N_14511,N_13257,N_14103);
nor U14512 (N_14512,N_13662,N_13490);
xor U14513 (N_14513,N_13755,N_13201);
and U14514 (N_14514,N_13356,N_13691);
xor U14515 (N_14515,N_13878,N_13453);
xor U14516 (N_14516,N_13346,N_14215);
or U14517 (N_14517,N_13782,N_13493);
xor U14518 (N_14518,N_13530,N_13980);
nand U14519 (N_14519,N_13884,N_13567);
nand U14520 (N_14520,N_13640,N_14098);
nand U14521 (N_14521,N_13632,N_13979);
nand U14522 (N_14522,N_14321,N_13909);
and U14523 (N_14523,N_13803,N_14195);
nand U14524 (N_14524,N_13516,N_13347);
xnor U14525 (N_14525,N_14371,N_13480);
nand U14526 (N_14526,N_14004,N_13726);
nor U14527 (N_14527,N_13813,N_13398);
nor U14528 (N_14528,N_14208,N_14383);
and U14529 (N_14529,N_14116,N_14237);
xor U14530 (N_14530,N_14246,N_14209);
nand U14531 (N_14531,N_14203,N_14393);
and U14532 (N_14532,N_14154,N_13837);
xnor U14533 (N_14533,N_13307,N_13557);
nand U14534 (N_14534,N_13559,N_13325);
and U14535 (N_14535,N_14077,N_14163);
and U14536 (N_14536,N_13209,N_13866);
xor U14537 (N_14537,N_14041,N_13677);
or U14538 (N_14538,N_14288,N_13619);
and U14539 (N_14539,N_13903,N_14048);
and U14540 (N_14540,N_14212,N_14024);
or U14541 (N_14541,N_13807,N_14398);
and U14542 (N_14542,N_13264,N_14172);
or U14543 (N_14543,N_13930,N_14200);
nor U14544 (N_14544,N_13641,N_13648);
xnor U14545 (N_14545,N_13798,N_13902);
nand U14546 (N_14546,N_13655,N_14340);
nand U14547 (N_14547,N_14075,N_14223);
nor U14548 (N_14548,N_14126,N_14216);
or U14549 (N_14549,N_13386,N_14029);
xor U14550 (N_14550,N_14284,N_13778);
or U14551 (N_14551,N_13362,N_14167);
or U14552 (N_14552,N_13337,N_14175);
nand U14553 (N_14553,N_14222,N_14385);
xnor U14554 (N_14554,N_13997,N_14304);
nor U14555 (N_14555,N_13749,N_13606);
or U14556 (N_14556,N_14247,N_14331);
and U14557 (N_14557,N_14156,N_14232);
xnor U14558 (N_14558,N_13333,N_14248);
or U14559 (N_14559,N_14236,N_13546);
nand U14560 (N_14560,N_13880,N_13306);
xor U14561 (N_14561,N_13531,N_13908);
or U14562 (N_14562,N_13417,N_13698);
and U14563 (N_14563,N_14124,N_13564);
or U14564 (N_14564,N_13541,N_14293);
nand U14565 (N_14565,N_13224,N_13867);
and U14566 (N_14566,N_13560,N_13777);
and U14567 (N_14567,N_13502,N_13896);
or U14568 (N_14568,N_13563,N_14272);
nand U14569 (N_14569,N_13824,N_13566);
nand U14570 (N_14570,N_13455,N_14224);
and U14571 (N_14571,N_13579,N_13626);
xnor U14572 (N_14572,N_13554,N_13792);
xnor U14573 (N_14573,N_13297,N_14199);
xnor U14574 (N_14574,N_14260,N_13919);
or U14575 (N_14575,N_14108,N_13956);
and U14576 (N_14576,N_13609,N_14392);
xnor U14577 (N_14577,N_14142,N_13614);
xor U14578 (N_14578,N_13534,N_14059);
nand U14579 (N_14579,N_13612,N_13916);
nor U14580 (N_14580,N_13915,N_13585);
and U14581 (N_14581,N_14348,N_13728);
nor U14582 (N_14582,N_14226,N_14258);
nand U14583 (N_14583,N_13374,N_13938);
nor U14584 (N_14584,N_14053,N_13724);
nor U14585 (N_14585,N_13844,N_14372);
nand U14586 (N_14586,N_13372,N_13744);
or U14587 (N_14587,N_14399,N_13543);
and U14588 (N_14588,N_13886,N_14257);
and U14589 (N_14589,N_13832,N_13793);
and U14590 (N_14590,N_13504,N_13378);
nand U14591 (N_14591,N_13366,N_13978);
and U14592 (N_14592,N_14082,N_13252);
or U14593 (N_14593,N_14080,N_14262);
xor U14594 (N_14594,N_13227,N_13989);
nor U14595 (N_14595,N_13851,N_14290);
nor U14596 (N_14596,N_13710,N_13230);
and U14597 (N_14597,N_13812,N_14051);
xnor U14598 (N_14598,N_13219,N_14190);
and U14599 (N_14599,N_13383,N_14366);
xnor U14600 (N_14600,N_13668,N_14005);
or U14601 (N_14601,N_13678,N_13864);
xnor U14602 (N_14602,N_14378,N_13215);
xnor U14603 (N_14603,N_13570,N_13746);
or U14604 (N_14604,N_14279,N_14188);
xor U14605 (N_14605,N_14373,N_13451);
and U14606 (N_14606,N_14171,N_14058);
nand U14607 (N_14607,N_13211,N_13838);
and U14608 (N_14608,N_14202,N_13229);
or U14609 (N_14609,N_13716,N_14322);
nor U14610 (N_14610,N_13548,N_13401);
nor U14611 (N_14611,N_13962,N_13363);
and U14612 (N_14612,N_14213,N_13783);
or U14613 (N_14613,N_14084,N_14127);
nor U14614 (N_14614,N_13466,N_14379);
xor U14615 (N_14615,N_13637,N_14158);
nor U14616 (N_14616,N_13430,N_14181);
and U14617 (N_14617,N_14100,N_14111);
and U14618 (N_14618,N_13487,N_13242);
nand U14619 (N_14619,N_14249,N_13472);
nand U14620 (N_14620,N_13513,N_13898);
xnor U14621 (N_14621,N_14317,N_13507);
and U14622 (N_14622,N_13427,N_13561);
or U14623 (N_14623,N_14211,N_14197);
xnor U14624 (N_14624,N_13890,N_13329);
or U14625 (N_14625,N_13808,N_13247);
nor U14626 (N_14626,N_13418,N_14064);
or U14627 (N_14627,N_13822,N_14314);
and U14628 (N_14628,N_13551,N_13906);
xor U14629 (N_14629,N_13319,N_13488);
nor U14630 (N_14630,N_13775,N_14137);
or U14631 (N_14631,N_13235,N_14072);
xor U14632 (N_14632,N_13857,N_13988);
and U14633 (N_14633,N_14356,N_14134);
nand U14634 (N_14634,N_13425,N_13713);
and U14635 (N_14635,N_13920,N_13390);
and U14636 (N_14636,N_13791,N_13287);
nor U14637 (N_14637,N_13663,N_14300);
or U14638 (N_14638,N_13463,N_13309);
and U14639 (N_14639,N_13433,N_13471);
nand U14640 (N_14640,N_13478,N_13972);
xnor U14641 (N_14641,N_13279,N_13638);
or U14642 (N_14642,N_14110,N_13617);
nor U14643 (N_14643,N_13742,N_14093);
or U14644 (N_14644,N_14280,N_13210);
nand U14645 (N_14645,N_13537,N_14165);
nor U14646 (N_14646,N_14205,N_13829);
nand U14647 (N_14647,N_14239,N_13348);
or U14648 (N_14648,N_13259,N_13911);
nand U14649 (N_14649,N_13359,N_13344);
xnor U14650 (N_14650,N_14113,N_13739);
xor U14651 (N_14651,N_14169,N_13816);
nor U14652 (N_14652,N_14302,N_13611);
and U14653 (N_14653,N_13436,N_14380);
and U14654 (N_14654,N_13647,N_13465);
and U14655 (N_14655,N_13624,N_13873);
or U14656 (N_14656,N_14141,N_13553);
and U14657 (N_14657,N_13571,N_13802);
nor U14658 (N_14658,N_13737,N_13723);
nor U14659 (N_14659,N_14161,N_13833);
xnor U14660 (N_14660,N_13562,N_13690);
nor U14661 (N_14661,N_13301,N_13627);
nor U14662 (N_14662,N_14390,N_13448);
and U14663 (N_14663,N_13521,N_13821);
or U14664 (N_14664,N_13581,N_13538);
nand U14665 (N_14665,N_13620,N_13584);
or U14666 (N_14666,N_13693,N_14244);
and U14667 (N_14667,N_13766,N_14362);
xor U14668 (N_14668,N_13961,N_14063);
or U14669 (N_14669,N_14253,N_14255);
xnor U14670 (N_14670,N_14016,N_13858);
nor U14671 (N_14671,N_13540,N_13389);
or U14672 (N_14672,N_13940,N_13405);
xnor U14673 (N_14673,N_13275,N_13918);
nor U14674 (N_14674,N_14311,N_13313);
and U14675 (N_14675,N_13470,N_14240);
or U14676 (N_14676,N_14395,N_13320);
nand U14677 (N_14677,N_14015,N_14243);
nand U14678 (N_14678,N_14125,N_13426);
nor U14679 (N_14679,N_13601,N_14281);
and U14680 (N_14680,N_13532,N_13872);
or U14681 (N_14681,N_13987,N_13456);
nand U14682 (N_14682,N_13774,N_13524);
xor U14683 (N_14683,N_13283,N_13618);
xnor U14684 (N_14684,N_13670,N_13600);
nand U14685 (N_14685,N_13365,N_13269);
and U14686 (N_14686,N_13674,N_14153);
and U14687 (N_14687,N_13790,N_13879);
xor U14688 (N_14688,N_13340,N_14358);
or U14689 (N_14689,N_13776,N_13786);
xor U14690 (N_14690,N_14173,N_13654);
and U14691 (N_14691,N_14049,N_13497);
nor U14692 (N_14692,N_13395,N_13796);
nand U14693 (N_14693,N_14312,N_13323);
nand U14694 (N_14694,N_13651,N_13957);
or U14695 (N_14695,N_14259,N_13454);
nor U14696 (N_14696,N_13280,N_13828);
xor U14697 (N_14697,N_13496,N_14241);
or U14698 (N_14698,N_13985,N_13893);
and U14699 (N_14699,N_13661,N_14376);
xor U14700 (N_14700,N_13239,N_13892);
xor U14701 (N_14701,N_13709,N_14354);
or U14702 (N_14702,N_13452,N_13860);
and U14703 (N_14703,N_13300,N_14140);
xor U14704 (N_14704,N_13492,N_13969);
nor U14705 (N_14705,N_13349,N_14364);
nor U14706 (N_14706,N_13771,N_13667);
xnor U14707 (N_14707,N_13214,N_13971);
xnor U14708 (N_14708,N_13547,N_13721);
nor U14709 (N_14709,N_13745,N_14042);
xor U14710 (N_14710,N_13205,N_13923);
nand U14711 (N_14711,N_14271,N_13751);
nand U14712 (N_14712,N_14201,N_13231);
xor U14713 (N_14713,N_13788,N_14296);
xor U14714 (N_14714,N_13586,N_14011);
xnor U14715 (N_14715,N_14069,N_13901);
nand U14716 (N_14716,N_13941,N_13409);
and U14717 (N_14717,N_13964,N_14353);
nor U14718 (N_14718,N_13604,N_13784);
nor U14719 (N_14719,N_14263,N_13760);
and U14720 (N_14720,N_13912,N_14286);
or U14721 (N_14721,N_14268,N_13679);
and U14722 (N_14722,N_14013,N_13993);
or U14723 (N_14723,N_13944,N_14273);
nor U14724 (N_14724,N_13761,N_13871);
and U14725 (N_14725,N_13330,N_14198);
or U14726 (N_14726,N_13810,N_14078);
nand U14727 (N_14727,N_14214,N_13248);
or U14728 (N_14728,N_13929,N_13469);
nor U14729 (N_14729,N_13336,N_14020);
nand U14730 (N_14730,N_13615,N_13402);
or U14731 (N_14731,N_13491,N_14339);
or U14732 (N_14732,N_14132,N_14238);
or U14733 (N_14733,N_13268,N_13485);
and U14734 (N_14734,N_14360,N_13768);
and U14735 (N_14735,N_13501,N_13370);
or U14736 (N_14736,N_13569,N_13271);
xnor U14737 (N_14737,N_13535,N_13447);
xnor U14738 (N_14738,N_13577,N_13467);
and U14739 (N_14739,N_13757,N_13913);
nand U14740 (N_14740,N_13422,N_14256);
nand U14741 (N_14741,N_13583,N_14295);
or U14742 (N_14742,N_13644,N_14228);
nand U14743 (N_14743,N_13686,N_14164);
nand U14744 (N_14744,N_13597,N_13603);
nand U14745 (N_14745,N_14105,N_13605);
nand U14746 (N_14746,N_13368,N_13717);
xnor U14747 (N_14747,N_13266,N_13228);
and U14748 (N_14748,N_13594,N_13596);
xnor U14749 (N_14749,N_13805,N_13818);
nor U14750 (N_14750,N_13899,N_13827);
nor U14751 (N_14751,N_13894,N_13545);
xor U14752 (N_14752,N_13429,N_13876);
nor U14753 (N_14753,N_14394,N_13982);
or U14754 (N_14754,N_13396,N_14365);
or U14755 (N_14755,N_13787,N_13765);
xor U14756 (N_14756,N_13423,N_14387);
nor U14757 (N_14757,N_14250,N_14152);
or U14758 (N_14758,N_13332,N_14017);
nor U14759 (N_14759,N_13441,N_13664);
nor U14760 (N_14760,N_14018,N_14225);
xor U14761 (N_14761,N_13317,N_14149);
xnor U14762 (N_14762,N_13438,N_13509);
nand U14763 (N_14763,N_13649,N_13639);
nor U14764 (N_14764,N_13515,N_14370);
nor U14765 (N_14765,N_14159,N_14309);
nor U14766 (N_14766,N_13711,N_13650);
or U14767 (N_14767,N_13510,N_13743);
nor U14768 (N_14768,N_14278,N_14043);
nand U14769 (N_14769,N_13274,N_13935);
nor U14770 (N_14770,N_13326,N_13354);
and U14771 (N_14771,N_13220,N_14265);
or U14772 (N_14772,N_14007,N_13568);
nand U14773 (N_14773,N_13412,N_13573);
or U14774 (N_14774,N_14055,N_13853);
and U14775 (N_14775,N_13253,N_13636);
nand U14776 (N_14776,N_14194,N_14139);
xnor U14777 (N_14777,N_13652,N_13719);
nor U14778 (N_14778,N_13590,N_13841);
and U14779 (N_14779,N_13865,N_13981);
xor U14780 (N_14780,N_13970,N_13293);
or U14781 (N_14781,N_13684,N_14282);
xor U14782 (N_14782,N_13635,N_13276);
xnor U14783 (N_14783,N_13394,N_13482);
nand U14784 (N_14784,N_14233,N_13486);
and U14785 (N_14785,N_13905,N_13328);
nor U14786 (N_14786,N_13922,N_14030);
nand U14787 (N_14787,N_13291,N_14287);
nand U14788 (N_14788,N_13519,N_14131);
or U14789 (N_14789,N_13544,N_14334);
xnor U14790 (N_14790,N_14033,N_13705);
and U14791 (N_14791,N_13272,N_13387);
or U14792 (N_14792,N_14130,N_14298);
and U14793 (N_14793,N_14361,N_13267);
or U14794 (N_14794,N_13718,N_14148);
or U14795 (N_14795,N_13208,N_13446);
and U14796 (N_14796,N_13460,N_14135);
or U14797 (N_14797,N_13255,N_13897);
xor U14798 (N_14798,N_14081,N_14251);
nand U14799 (N_14799,N_13804,N_14231);
and U14800 (N_14800,N_13552,N_14050);
and U14801 (N_14801,N_13392,N_13439);
and U14802 (N_14802,N_13610,N_13825);
and U14803 (N_14803,N_13675,N_14031);
or U14804 (N_14804,N_13361,N_13550);
nand U14805 (N_14805,N_13939,N_13643);
and U14806 (N_14806,N_13733,N_14144);
and U14807 (N_14807,N_14210,N_13207);
nor U14808 (N_14808,N_13494,N_13882);
and U14809 (N_14809,N_13285,N_13495);
xor U14810 (N_14810,N_13399,N_13773);
nand U14811 (N_14811,N_14316,N_14157);
or U14812 (N_14812,N_13558,N_14355);
nand U14813 (N_14813,N_13450,N_13992);
nor U14814 (N_14814,N_14347,N_13397);
xor U14815 (N_14815,N_13216,N_14086);
nor U14816 (N_14816,N_13377,N_13536);
and U14817 (N_14817,N_13850,N_13355);
and U14818 (N_14818,N_14039,N_13794);
and U14819 (N_14819,N_13304,N_13692);
xor U14820 (N_14820,N_13296,N_14002);
nand U14821 (N_14821,N_13288,N_13484);
nand U14822 (N_14822,N_14323,N_13400);
nand U14823 (N_14823,N_14000,N_13646);
or U14824 (N_14824,N_14206,N_14088);
nor U14825 (N_14825,N_13292,N_13498);
nand U14826 (N_14826,N_14276,N_13565);
xnor U14827 (N_14827,N_13479,N_14229);
and U14828 (N_14828,N_14052,N_13442);
xnor U14829 (N_14829,N_13958,N_13870);
nor U14830 (N_14830,N_14332,N_13299);
nand U14831 (N_14831,N_13952,N_13428);
xnor U14832 (N_14832,N_13592,N_13251);
or U14833 (N_14833,N_13924,N_13420);
or U14834 (N_14834,N_14328,N_14102);
or U14835 (N_14835,N_13602,N_14377);
nand U14836 (N_14836,N_13700,N_13673);
and U14837 (N_14837,N_14329,N_13382);
xnor U14838 (N_14838,N_13735,N_13539);
nand U14839 (N_14839,N_14138,N_14009);
xor U14840 (N_14840,N_13200,N_13373);
nand U14841 (N_14841,N_13975,N_13385);
nand U14842 (N_14842,N_14112,N_13444);
nand U14843 (N_14843,N_13875,N_13701);
and U14844 (N_14844,N_13888,N_14391);
or U14845 (N_14845,N_13806,N_13819);
xor U14846 (N_14846,N_14006,N_13984);
and U14847 (N_14847,N_14337,N_14336);
or U14848 (N_14848,N_13522,N_13823);
or U14849 (N_14849,N_13926,N_14067);
nand U14850 (N_14850,N_14397,N_14174);
and U14851 (N_14851,N_13687,N_13623);
xor U14852 (N_14852,N_13526,N_13834);
and U14853 (N_14853,N_14034,N_13877);
nor U14854 (N_14854,N_13995,N_13968);
nor U14855 (N_14855,N_13863,N_14106);
or U14856 (N_14856,N_13244,N_14128);
nand U14857 (N_14857,N_14012,N_14357);
nor U14858 (N_14858,N_13830,N_13298);
or U14859 (N_14859,N_13353,N_13461);
or U14860 (N_14860,N_13889,N_14333);
or U14861 (N_14861,N_13795,N_13861);
nand U14862 (N_14862,N_13574,N_14221);
xnor U14863 (N_14863,N_13762,N_13593);
nor U14864 (N_14864,N_14032,N_13419);
or U14865 (N_14865,N_14254,N_14160);
or U14866 (N_14866,N_14073,N_13303);
nand U14867 (N_14867,N_14375,N_14325);
or U14868 (N_14868,N_14147,N_13518);
and U14869 (N_14869,N_14324,N_13669);
or U14870 (N_14870,N_14022,N_13234);
and U14871 (N_14871,N_14045,N_13250);
or U14872 (N_14872,N_13785,N_13874);
or U14873 (N_14873,N_13665,N_13582);
nor U14874 (N_14874,N_14186,N_13622);
or U14875 (N_14875,N_14245,N_13376);
xnor U14876 (N_14876,N_13511,N_14318);
nand U14877 (N_14877,N_14010,N_14019);
nor U14878 (N_14878,N_14096,N_14374);
xor U14879 (N_14879,N_13809,N_13311);
nand U14880 (N_14880,N_13727,N_13440);
and U14881 (N_14881,N_13826,N_13416);
or U14882 (N_14882,N_13588,N_14341);
nand U14883 (N_14883,N_13996,N_14054);
xor U14884 (N_14884,N_14070,N_13836);
and U14885 (N_14885,N_13580,N_14074);
and U14886 (N_14886,N_13549,N_13462);
xnor U14887 (N_14887,N_13763,N_13991);
xnor U14888 (N_14888,N_13388,N_13656);
and U14889 (N_14889,N_13702,N_13937);
nor U14890 (N_14890,N_14277,N_13671);
xnor U14891 (N_14891,N_13854,N_13697);
and U14892 (N_14892,N_14166,N_13236);
nor U14893 (N_14893,N_13708,N_13955);
and U14894 (N_14894,N_13927,N_13341);
or U14895 (N_14895,N_13855,N_13820);
xor U14896 (N_14896,N_13950,N_13443);
xor U14897 (N_14897,N_13948,N_13468);
nand U14898 (N_14898,N_14145,N_13249);
or U14899 (N_14899,N_14061,N_13699);
or U14900 (N_14900,N_13900,N_13327);
nand U14901 (N_14901,N_13666,N_13974);
or U14902 (N_14902,N_13294,N_14381);
nor U14903 (N_14903,N_14313,N_13435);
xor U14904 (N_14904,N_13928,N_13212);
nor U14905 (N_14905,N_13434,N_13845);
nand U14906 (N_14906,N_14343,N_13334);
or U14907 (N_14907,N_13895,N_14095);
nor U14908 (N_14908,N_13862,N_13459);
nand U14909 (N_14909,N_13414,N_13432);
nor U14910 (N_14910,N_14230,N_14275);
xor U14911 (N_14911,N_13314,N_13631);
and U14912 (N_14912,N_13931,N_13403);
nor U14913 (N_14913,N_13222,N_13642);
xor U14914 (N_14914,N_14346,N_13449);
and U14915 (N_14915,N_13967,N_13245);
xor U14916 (N_14916,N_14180,N_14036);
or U14917 (N_14917,N_14294,N_13847);
nand U14918 (N_14918,N_14170,N_13367);
and U14919 (N_14919,N_13204,N_13421);
and U14920 (N_14920,N_13815,N_13578);
nand U14921 (N_14921,N_13512,N_13315);
or U14922 (N_14922,N_14299,N_14327);
and U14923 (N_14923,N_14037,N_13848);
or U14924 (N_14924,N_13379,N_13653);
or U14925 (N_14925,N_13206,N_13607);
nand U14926 (N_14926,N_14104,N_13682);
xnor U14927 (N_14927,N_14183,N_13237);
or U14928 (N_14928,N_14307,N_13754);
xnor U14929 (N_14929,N_13704,N_14367);
xor U14930 (N_14930,N_13842,N_14352);
nor U14931 (N_14931,N_13722,N_13780);
nor U14932 (N_14932,N_13343,N_14162);
nor U14933 (N_14933,N_13523,N_13431);
and U14934 (N_14934,N_13907,N_13695);
nand U14935 (N_14935,N_13608,N_13595);
or U14936 (N_14936,N_14071,N_13312);
or U14937 (N_14937,N_13277,N_14193);
or U14938 (N_14938,N_14264,N_13933);
or U14939 (N_14939,N_14187,N_13270);
xor U14940 (N_14940,N_14025,N_13759);
or U14941 (N_14941,N_13413,N_13598);
nor U14942 (N_14942,N_13358,N_13936);
nand U14943 (N_14943,N_13380,N_14386);
or U14944 (N_14944,N_13998,N_13840);
nand U14945 (N_14945,N_13963,N_14068);
or U14946 (N_14946,N_13712,N_13707);
or U14947 (N_14947,N_13799,N_14310);
and U14948 (N_14948,N_13856,N_14168);
nand U14949 (N_14949,N_13904,N_13887);
xor U14950 (N_14950,N_13634,N_13503);
nand U14951 (N_14951,N_13881,N_14062);
and U14952 (N_14952,N_13241,N_13302);
xor U14953 (N_14953,N_14291,N_13714);
or U14954 (N_14954,N_13408,N_13683);
and U14955 (N_14955,N_14185,N_14326);
nand U14956 (N_14956,N_13688,N_13917);
and U14957 (N_14957,N_13339,N_13885);
xor U14958 (N_14958,N_13859,N_13835);
or U14959 (N_14959,N_13914,N_13983);
and U14960 (N_14960,N_13781,N_13375);
and U14961 (N_14961,N_13694,N_13576);
nand U14962 (N_14962,N_14133,N_13525);
and U14963 (N_14963,N_13764,N_14303);
and U14964 (N_14964,N_13238,N_13731);
nor U14965 (N_14965,N_13947,N_13587);
xor U14966 (N_14966,N_14384,N_14092);
or U14967 (N_14967,N_13517,N_13369);
or U14968 (N_14968,N_13246,N_13282);
and U14969 (N_14969,N_14123,N_14191);
nor U14970 (N_14970,N_13217,N_13464);
nand U14971 (N_14971,N_14155,N_14057);
xor U14972 (N_14972,N_14089,N_13424);
or U14973 (N_14973,N_13203,N_14192);
or U14974 (N_14974,N_14090,N_13476);
xor U14975 (N_14975,N_14388,N_14027);
and U14976 (N_14976,N_13360,N_14008);
or U14977 (N_14977,N_13289,N_13658);
and U14978 (N_14978,N_13254,N_14056);
xnor U14979 (N_14979,N_13575,N_13814);
nor U14980 (N_14980,N_13218,N_13976);
or U14981 (N_14981,N_14177,N_14040);
or U14982 (N_14982,N_13335,N_13528);
nor U14983 (N_14983,N_13734,N_13741);
xor U14984 (N_14984,N_13747,N_14292);
nor U14985 (N_14985,N_13364,N_14178);
or U14986 (N_14986,N_13977,N_13672);
or U14987 (N_14987,N_13750,N_13345);
and U14988 (N_14988,N_13846,N_13572);
xor U14989 (N_14989,N_14097,N_13657);
xor U14990 (N_14990,N_13946,N_14351);
nor U14991 (N_14991,N_14315,N_14285);
nor U14992 (N_14992,N_13457,N_13629);
or U14993 (N_14993,N_14085,N_14305);
nor U14994 (N_14994,N_14219,N_13839);
xnor U14995 (N_14995,N_13659,N_13680);
xnor U14996 (N_14996,N_14227,N_14119);
nand U14997 (N_14997,N_13748,N_13290);
nor U14998 (N_14998,N_13990,N_14301);
nor U14999 (N_14999,N_14044,N_13779);
nand U15000 (N_15000,N_13517,N_14001);
nor U15001 (N_15001,N_13751,N_13376);
xnor U15002 (N_15002,N_13881,N_13703);
nand U15003 (N_15003,N_14041,N_13859);
or U15004 (N_15004,N_14146,N_14274);
or U15005 (N_15005,N_13682,N_13811);
xor U15006 (N_15006,N_13397,N_14211);
nor U15007 (N_15007,N_14147,N_13336);
nor U15008 (N_15008,N_13347,N_14119);
nand U15009 (N_15009,N_13815,N_13465);
nor U15010 (N_15010,N_13868,N_13850);
or U15011 (N_15011,N_14363,N_13947);
and U15012 (N_15012,N_13613,N_13518);
and U15013 (N_15013,N_14331,N_13975);
xnor U15014 (N_15014,N_14232,N_14090);
nor U15015 (N_15015,N_13571,N_14256);
nor U15016 (N_15016,N_14074,N_14380);
xnor U15017 (N_15017,N_13554,N_13385);
and U15018 (N_15018,N_13663,N_14138);
nand U15019 (N_15019,N_13591,N_14076);
or U15020 (N_15020,N_13412,N_13650);
and U15021 (N_15021,N_13930,N_13675);
nand U15022 (N_15022,N_14128,N_14116);
nor U15023 (N_15023,N_13274,N_13538);
xnor U15024 (N_15024,N_13735,N_13254);
nor U15025 (N_15025,N_13792,N_13363);
xnor U15026 (N_15026,N_14231,N_13741);
nor U15027 (N_15027,N_14292,N_13797);
or U15028 (N_15028,N_14370,N_13753);
nand U15029 (N_15029,N_13304,N_13676);
nor U15030 (N_15030,N_14033,N_14236);
or U15031 (N_15031,N_13327,N_14310);
nand U15032 (N_15032,N_13702,N_14277);
nand U15033 (N_15033,N_14017,N_13959);
and U15034 (N_15034,N_14284,N_14243);
nand U15035 (N_15035,N_13826,N_13816);
and U15036 (N_15036,N_14341,N_13327);
or U15037 (N_15037,N_13246,N_13409);
and U15038 (N_15038,N_13800,N_13352);
and U15039 (N_15039,N_14097,N_14295);
or U15040 (N_15040,N_13855,N_14321);
and U15041 (N_15041,N_13253,N_13972);
and U15042 (N_15042,N_13565,N_13235);
and U15043 (N_15043,N_14393,N_14241);
and U15044 (N_15044,N_13947,N_13207);
nor U15045 (N_15045,N_14146,N_14262);
xor U15046 (N_15046,N_14149,N_13711);
or U15047 (N_15047,N_13281,N_14184);
nand U15048 (N_15048,N_13902,N_14244);
nand U15049 (N_15049,N_14166,N_13569);
nor U15050 (N_15050,N_14037,N_14297);
nor U15051 (N_15051,N_13519,N_14119);
or U15052 (N_15052,N_14369,N_13687);
or U15053 (N_15053,N_13827,N_13429);
xnor U15054 (N_15054,N_13661,N_13761);
nor U15055 (N_15055,N_14118,N_13653);
xor U15056 (N_15056,N_13204,N_13212);
xnor U15057 (N_15057,N_14382,N_13443);
nand U15058 (N_15058,N_13269,N_13425);
and U15059 (N_15059,N_13565,N_13415);
and U15060 (N_15060,N_13285,N_14370);
nand U15061 (N_15061,N_13429,N_13915);
and U15062 (N_15062,N_13957,N_14285);
or U15063 (N_15063,N_13519,N_13657);
nand U15064 (N_15064,N_13551,N_13200);
and U15065 (N_15065,N_13825,N_13920);
nor U15066 (N_15066,N_14076,N_13278);
xor U15067 (N_15067,N_13996,N_14302);
xnor U15068 (N_15068,N_14329,N_13209);
nor U15069 (N_15069,N_13615,N_14397);
and U15070 (N_15070,N_14242,N_14115);
or U15071 (N_15071,N_13339,N_14365);
or U15072 (N_15072,N_13621,N_13749);
or U15073 (N_15073,N_13991,N_14287);
nand U15074 (N_15074,N_13967,N_14097);
nor U15075 (N_15075,N_13273,N_13474);
nor U15076 (N_15076,N_14187,N_13997);
nor U15077 (N_15077,N_14052,N_13916);
and U15078 (N_15078,N_13813,N_14182);
or U15079 (N_15079,N_13564,N_13651);
nor U15080 (N_15080,N_14278,N_13339);
nand U15081 (N_15081,N_13210,N_13369);
nor U15082 (N_15082,N_13263,N_13862);
or U15083 (N_15083,N_14351,N_13565);
or U15084 (N_15084,N_14390,N_14362);
or U15085 (N_15085,N_14361,N_13654);
or U15086 (N_15086,N_13989,N_13622);
nor U15087 (N_15087,N_14342,N_13200);
nand U15088 (N_15088,N_13279,N_13999);
and U15089 (N_15089,N_13979,N_13528);
xnor U15090 (N_15090,N_13898,N_14372);
and U15091 (N_15091,N_14267,N_13334);
and U15092 (N_15092,N_13931,N_14324);
nand U15093 (N_15093,N_13704,N_14088);
xor U15094 (N_15094,N_13584,N_13335);
and U15095 (N_15095,N_13313,N_14362);
xor U15096 (N_15096,N_14356,N_13275);
nand U15097 (N_15097,N_13499,N_13977);
nor U15098 (N_15098,N_14125,N_13525);
and U15099 (N_15099,N_13711,N_13661);
xnor U15100 (N_15100,N_13797,N_13210);
and U15101 (N_15101,N_13445,N_14151);
or U15102 (N_15102,N_14023,N_13366);
nand U15103 (N_15103,N_13934,N_13860);
nand U15104 (N_15104,N_13835,N_13972);
nor U15105 (N_15105,N_13498,N_13945);
nor U15106 (N_15106,N_13597,N_13414);
nor U15107 (N_15107,N_14262,N_14325);
and U15108 (N_15108,N_14351,N_14112);
nand U15109 (N_15109,N_13966,N_13301);
and U15110 (N_15110,N_14391,N_13952);
and U15111 (N_15111,N_13516,N_13773);
xnor U15112 (N_15112,N_13514,N_14272);
nor U15113 (N_15113,N_13323,N_14015);
or U15114 (N_15114,N_14168,N_14170);
nand U15115 (N_15115,N_14204,N_13442);
nor U15116 (N_15116,N_14187,N_14153);
and U15117 (N_15117,N_13666,N_14024);
or U15118 (N_15118,N_13968,N_13202);
or U15119 (N_15119,N_14039,N_13958);
or U15120 (N_15120,N_14374,N_14104);
and U15121 (N_15121,N_13904,N_14039);
nor U15122 (N_15122,N_13967,N_13447);
nor U15123 (N_15123,N_13943,N_13208);
or U15124 (N_15124,N_13780,N_13936);
or U15125 (N_15125,N_13671,N_14318);
or U15126 (N_15126,N_13717,N_14004);
xor U15127 (N_15127,N_13457,N_14239);
nand U15128 (N_15128,N_13658,N_13351);
xnor U15129 (N_15129,N_14116,N_13467);
nand U15130 (N_15130,N_13861,N_14114);
nor U15131 (N_15131,N_13228,N_13757);
nand U15132 (N_15132,N_13398,N_14263);
and U15133 (N_15133,N_13653,N_13811);
and U15134 (N_15134,N_14228,N_13828);
or U15135 (N_15135,N_14067,N_14230);
or U15136 (N_15136,N_13330,N_13220);
or U15137 (N_15137,N_13708,N_13939);
and U15138 (N_15138,N_13857,N_13292);
nor U15139 (N_15139,N_13564,N_14368);
nand U15140 (N_15140,N_14019,N_13764);
xnor U15141 (N_15141,N_13772,N_13519);
and U15142 (N_15142,N_13825,N_14081);
or U15143 (N_15143,N_13391,N_13992);
xnor U15144 (N_15144,N_13837,N_14059);
and U15145 (N_15145,N_13826,N_14225);
nand U15146 (N_15146,N_14046,N_14069);
or U15147 (N_15147,N_14049,N_13926);
or U15148 (N_15148,N_13404,N_13746);
nand U15149 (N_15149,N_13200,N_13507);
or U15150 (N_15150,N_13965,N_13392);
or U15151 (N_15151,N_13803,N_13481);
nor U15152 (N_15152,N_13561,N_13538);
nand U15153 (N_15153,N_13505,N_13286);
nor U15154 (N_15154,N_13241,N_13723);
nor U15155 (N_15155,N_13918,N_13626);
xnor U15156 (N_15156,N_14029,N_14071);
xor U15157 (N_15157,N_13345,N_14306);
nand U15158 (N_15158,N_13705,N_13325);
nand U15159 (N_15159,N_14356,N_13857);
and U15160 (N_15160,N_13805,N_13726);
xor U15161 (N_15161,N_13539,N_14178);
and U15162 (N_15162,N_13794,N_13649);
nor U15163 (N_15163,N_13767,N_13849);
nor U15164 (N_15164,N_13496,N_14099);
nand U15165 (N_15165,N_14389,N_13300);
nor U15166 (N_15166,N_13316,N_14193);
and U15167 (N_15167,N_13214,N_13541);
xnor U15168 (N_15168,N_13494,N_13474);
nor U15169 (N_15169,N_14084,N_13339);
nor U15170 (N_15170,N_14227,N_13883);
nor U15171 (N_15171,N_13947,N_13683);
nand U15172 (N_15172,N_14087,N_13737);
xnor U15173 (N_15173,N_13281,N_13393);
nand U15174 (N_15174,N_14380,N_14389);
nand U15175 (N_15175,N_14315,N_13424);
xnor U15176 (N_15176,N_13477,N_13654);
nand U15177 (N_15177,N_14222,N_13583);
or U15178 (N_15178,N_13322,N_14136);
or U15179 (N_15179,N_13279,N_13475);
nor U15180 (N_15180,N_13976,N_13610);
and U15181 (N_15181,N_14002,N_14304);
or U15182 (N_15182,N_13367,N_13387);
and U15183 (N_15183,N_13456,N_14264);
nand U15184 (N_15184,N_13787,N_14372);
nor U15185 (N_15185,N_13779,N_14058);
nand U15186 (N_15186,N_14369,N_14362);
or U15187 (N_15187,N_13592,N_13219);
nand U15188 (N_15188,N_13491,N_13512);
nor U15189 (N_15189,N_14077,N_13938);
xor U15190 (N_15190,N_14281,N_13238);
nor U15191 (N_15191,N_14190,N_13909);
nand U15192 (N_15192,N_13360,N_14368);
or U15193 (N_15193,N_13994,N_14008);
nand U15194 (N_15194,N_14316,N_14330);
or U15195 (N_15195,N_14295,N_13750);
nor U15196 (N_15196,N_14239,N_13715);
xnor U15197 (N_15197,N_13976,N_14303);
nor U15198 (N_15198,N_13412,N_13950);
and U15199 (N_15199,N_13549,N_14266);
xnor U15200 (N_15200,N_13396,N_13316);
and U15201 (N_15201,N_14211,N_14076);
nand U15202 (N_15202,N_13900,N_14382);
and U15203 (N_15203,N_13753,N_13886);
or U15204 (N_15204,N_14364,N_13414);
nand U15205 (N_15205,N_13631,N_14113);
nor U15206 (N_15206,N_13906,N_13487);
or U15207 (N_15207,N_13313,N_13867);
nor U15208 (N_15208,N_13941,N_13895);
nand U15209 (N_15209,N_13467,N_13511);
nor U15210 (N_15210,N_13727,N_13582);
xor U15211 (N_15211,N_13523,N_14160);
nand U15212 (N_15212,N_13794,N_14097);
nand U15213 (N_15213,N_13456,N_13861);
xor U15214 (N_15214,N_13755,N_13723);
nand U15215 (N_15215,N_13780,N_13529);
nand U15216 (N_15216,N_13455,N_13758);
or U15217 (N_15217,N_13632,N_14234);
nor U15218 (N_15218,N_13513,N_14012);
xor U15219 (N_15219,N_13232,N_13890);
or U15220 (N_15220,N_13746,N_13474);
xor U15221 (N_15221,N_14220,N_14320);
nand U15222 (N_15222,N_13586,N_13925);
nand U15223 (N_15223,N_13533,N_13618);
or U15224 (N_15224,N_14240,N_14128);
nor U15225 (N_15225,N_13242,N_13700);
or U15226 (N_15226,N_13666,N_14226);
xor U15227 (N_15227,N_13596,N_13859);
xnor U15228 (N_15228,N_13651,N_14139);
nor U15229 (N_15229,N_13294,N_13535);
xnor U15230 (N_15230,N_13462,N_14001);
nor U15231 (N_15231,N_13762,N_14236);
or U15232 (N_15232,N_13895,N_14368);
or U15233 (N_15233,N_13416,N_13550);
nand U15234 (N_15234,N_13725,N_13251);
and U15235 (N_15235,N_13592,N_13252);
or U15236 (N_15236,N_13724,N_13579);
nand U15237 (N_15237,N_13280,N_14178);
or U15238 (N_15238,N_13625,N_13771);
or U15239 (N_15239,N_13346,N_13824);
or U15240 (N_15240,N_13667,N_13485);
xnor U15241 (N_15241,N_13594,N_13794);
and U15242 (N_15242,N_14188,N_14104);
and U15243 (N_15243,N_14085,N_14121);
or U15244 (N_15244,N_13533,N_13960);
nor U15245 (N_15245,N_14334,N_14280);
and U15246 (N_15246,N_13980,N_13840);
nor U15247 (N_15247,N_14262,N_13517);
nand U15248 (N_15248,N_14057,N_13486);
or U15249 (N_15249,N_13962,N_14398);
nor U15250 (N_15250,N_13284,N_13417);
nor U15251 (N_15251,N_14072,N_14211);
and U15252 (N_15252,N_13255,N_13283);
nand U15253 (N_15253,N_14036,N_14072);
or U15254 (N_15254,N_13860,N_13700);
and U15255 (N_15255,N_13927,N_13781);
xnor U15256 (N_15256,N_13977,N_13435);
and U15257 (N_15257,N_14203,N_13990);
and U15258 (N_15258,N_13897,N_14163);
or U15259 (N_15259,N_13811,N_14306);
and U15260 (N_15260,N_13463,N_13435);
or U15261 (N_15261,N_14257,N_13215);
or U15262 (N_15262,N_13300,N_13792);
and U15263 (N_15263,N_13249,N_13303);
xor U15264 (N_15264,N_13881,N_13826);
or U15265 (N_15265,N_13825,N_13303);
xor U15266 (N_15266,N_13519,N_13520);
xnor U15267 (N_15267,N_13816,N_13764);
xnor U15268 (N_15268,N_14119,N_13859);
xnor U15269 (N_15269,N_13531,N_13561);
or U15270 (N_15270,N_13477,N_14117);
or U15271 (N_15271,N_13230,N_14114);
nor U15272 (N_15272,N_13425,N_14278);
nand U15273 (N_15273,N_13647,N_13900);
and U15274 (N_15274,N_13678,N_14392);
nand U15275 (N_15275,N_13927,N_13257);
xor U15276 (N_15276,N_13877,N_13230);
nor U15277 (N_15277,N_13606,N_13965);
or U15278 (N_15278,N_13854,N_13834);
or U15279 (N_15279,N_13367,N_13851);
or U15280 (N_15280,N_14112,N_13829);
nand U15281 (N_15281,N_13432,N_13692);
nor U15282 (N_15282,N_13504,N_14368);
nand U15283 (N_15283,N_14325,N_14047);
nor U15284 (N_15284,N_13970,N_13296);
nand U15285 (N_15285,N_13989,N_13553);
or U15286 (N_15286,N_13631,N_13621);
nand U15287 (N_15287,N_13302,N_13545);
xor U15288 (N_15288,N_13626,N_13517);
or U15289 (N_15289,N_13822,N_13814);
and U15290 (N_15290,N_13673,N_13667);
xnor U15291 (N_15291,N_13746,N_13319);
and U15292 (N_15292,N_13678,N_13604);
xnor U15293 (N_15293,N_14186,N_13331);
nand U15294 (N_15294,N_13443,N_13663);
nand U15295 (N_15295,N_14248,N_13399);
xnor U15296 (N_15296,N_13337,N_13950);
nor U15297 (N_15297,N_13938,N_13920);
xor U15298 (N_15298,N_14320,N_14381);
xor U15299 (N_15299,N_14353,N_14183);
nand U15300 (N_15300,N_14057,N_13695);
xor U15301 (N_15301,N_13420,N_13683);
nor U15302 (N_15302,N_13696,N_13499);
nor U15303 (N_15303,N_13410,N_13377);
xnor U15304 (N_15304,N_14130,N_13290);
xor U15305 (N_15305,N_13502,N_13292);
xnor U15306 (N_15306,N_13902,N_13515);
nor U15307 (N_15307,N_13945,N_13555);
or U15308 (N_15308,N_14279,N_13758);
nand U15309 (N_15309,N_13456,N_14179);
or U15310 (N_15310,N_13781,N_13682);
xnor U15311 (N_15311,N_13335,N_13947);
xor U15312 (N_15312,N_13258,N_13855);
and U15313 (N_15313,N_14355,N_14369);
xnor U15314 (N_15314,N_13222,N_13472);
or U15315 (N_15315,N_13399,N_13727);
nand U15316 (N_15316,N_13269,N_14027);
xor U15317 (N_15317,N_13483,N_13554);
or U15318 (N_15318,N_13738,N_13204);
xnor U15319 (N_15319,N_14005,N_13758);
and U15320 (N_15320,N_13255,N_13790);
nand U15321 (N_15321,N_13718,N_14309);
nand U15322 (N_15322,N_13889,N_13792);
nor U15323 (N_15323,N_14042,N_13438);
nor U15324 (N_15324,N_13989,N_13446);
or U15325 (N_15325,N_13562,N_13441);
nand U15326 (N_15326,N_13935,N_14103);
nor U15327 (N_15327,N_13261,N_13908);
xnor U15328 (N_15328,N_14362,N_13364);
or U15329 (N_15329,N_14294,N_13313);
xnor U15330 (N_15330,N_14345,N_14292);
nor U15331 (N_15331,N_14270,N_13738);
xnor U15332 (N_15332,N_13204,N_13277);
and U15333 (N_15333,N_14348,N_13989);
nand U15334 (N_15334,N_14181,N_14101);
or U15335 (N_15335,N_14255,N_13603);
and U15336 (N_15336,N_13275,N_13820);
nor U15337 (N_15337,N_13474,N_14149);
nor U15338 (N_15338,N_13403,N_13218);
and U15339 (N_15339,N_14085,N_13429);
xnor U15340 (N_15340,N_13785,N_13271);
xor U15341 (N_15341,N_13892,N_13280);
or U15342 (N_15342,N_13819,N_14274);
xnor U15343 (N_15343,N_14376,N_14035);
or U15344 (N_15344,N_14017,N_14093);
and U15345 (N_15345,N_13755,N_14153);
nor U15346 (N_15346,N_14075,N_13763);
xor U15347 (N_15347,N_14057,N_13748);
nand U15348 (N_15348,N_14076,N_14141);
xnor U15349 (N_15349,N_13387,N_13441);
xor U15350 (N_15350,N_13751,N_13839);
nor U15351 (N_15351,N_13969,N_13498);
nand U15352 (N_15352,N_14166,N_13307);
or U15353 (N_15353,N_13405,N_13974);
nor U15354 (N_15354,N_13701,N_13655);
nand U15355 (N_15355,N_13264,N_13832);
nand U15356 (N_15356,N_13615,N_13270);
nand U15357 (N_15357,N_14066,N_13936);
nand U15358 (N_15358,N_13457,N_14219);
and U15359 (N_15359,N_13305,N_14330);
nor U15360 (N_15360,N_13718,N_13691);
or U15361 (N_15361,N_13674,N_14241);
nor U15362 (N_15362,N_14316,N_13723);
and U15363 (N_15363,N_14338,N_14393);
and U15364 (N_15364,N_14095,N_13940);
and U15365 (N_15365,N_13651,N_14090);
nor U15366 (N_15366,N_13898,N_13821);
nor U15367 (N_15367,N_13493,N_13299);
nor U15368 (N_15368,N_13710,N_13214);
nand U15369 (N_15369,N_14044,N_13963);
xor U15370 (N_15370,N_14374,N_14181);
or U15371 (N_15371,N_13738,N_14072);
and U15372 (N_15372,N_14297,N_13611);
or U15373 (N_15373,N_14194,N_14104);
nand U15374 (N_15374,N_13848,N_13293);
and U15375 (N_15375,N_14337,N_13864);
or U15376 (N_15376,N_13675,N_13206);
xor U15377 (N_15377,N_14186,N_13497);
nor U15378 (N_15378,N_13787,N_14075);
nor U15379 (N_15379,N_13735,N_14273);
and U15380 (N_15380,N_13630,N_14054);
nor U15381 (N_15381,N_13846,N_13254);
nor U15382 (N_15382,N_13704,N_13288);
and U15383 (N_15383,N_14198,N_13639);
or U15384 (N_15384,N_14150,N_13462);
or U15385 (N_15385,N_13790,N_13280);
nor U15386 (N_15386,N_13616,N_13239);
nand U15387 (N_15387,N_13654,N_13777);
nand U15388 (N_15388,N_13976,N_13840);
and U15389 (N_15389,N_13752,N_13635);
and U15390 (N_15390,N_13963,N_14236);
nand U15391 (N_15391,N_13479,N_13209);
nand U15392 (N_15392,N_13336,N_13335);
xor U15393 (N_15393,N_13451,N_13786);
or U15394 (N_15394,N_13542,N_13633);
nand U15395 (N_15395,N_14084,N_14344);
and U15396 (N_15396,N_14263,N_13887);
and U15397 (N_15397,N_13838,N_13654);
nand U15398 (N_15398,N_14060,N_13269);
and U15399 (N_15399,N_13295,N_13503);
and U15400 (N_15400,N_13256,N_14251);
xor U15401 (N_15401,N_13600,N_13514);
xor U15402 (N_15402,N_14048,N_14182);
or U15403 (N_15403,N_14333,N_14026);
nand U15404 (N_15404,N_14386,N_13719);
nor U15405 (N_15405,N_13618,N_13547);
nor U15406 (N_15406,N_14263,N_14032);
or U15407 (N_15407,N_13427,N_14208);
nor U15408 (N_15408,N_13437,N_13310);
or U15409 (N_15409,N_13432,N_13545);
and U15410 (N_15410,N_13567,N_14093);
nand U15411 (N_15411,N_14107,N_13319);
nor U15412 (N_15412,N_13681,N_14116);
or U15413 (N_15413,N_13240,N_13793);
or U15414 (N_15414,N_14209,N_13437);
nand U15415 (N_15415,N_13653,N_14166);
and U15416 (N_15416,N_14115,N_13713);
xor U15417 (N_15417,N_13842,N_13258);
or U15418 (N_15418,N_13562,N_13328);
xnor U15419 (N_15419,N_13551,N_14294);
nor U15420 (N_15420,N_13330,N_13302);
xor U15421 (N_15421,N_13371,N_13356);
or U15422 (N_15422,N_13283,N_13555);
nor U15423 (N_15423,N_14007,N_13332);
nand U15424 (N_15424,N_13484,N_14157);
and U15425 (N_15425,N_13336,N_13974);
xnor U15426 (N_15426,N_13464,N_13598);
nand U15427 (N_15427,N_13764,N_13701);
nand U15428 (N_15428,N_14307,N_14334);
nand U15429 (N_15429,N_13291,N_14169);
xor U15430 (N_15430,N_14152,N_13796);
or U15431 (N_15431,N_13972,N_14347);
nor U15432 (N_15432,N_13805,N_13420);
nor U15433 (N_15433,N_14041,N_14216);
xnor U15434 (N_15434,N_13691,N_13527);
or U15435 (N_15435,N_14399,N_14082);
nor U15436 (N_15436,N_13613,N_13255);
or U15437 (N_15437,N_13625,N_13200);
nand U15438 (N_15438,N_14123,N_13309);
nand U15439 (N_15439,N_14177,N_13677);
xor U15440 (N_15440,N_13864,N_14030);
xnor U15441 (N_15441,N_13544,N_14184);
nor U15442 (N_15442,N_13875,N_14170);
xor U15443 (N_15443,N_13520,N_13890);
or U15444 (N_15444,N_14365,N_13476);
or U15445 (N_15445,N_13320,N_13910);
nand U15446 (N_15446,N_13449,N_13922);
or U15447 (N_15447,N_13228,N_13509);
and U15448 (N_15448,N_13492,N_13573);
xnor U15449 (N_15449,N_13715,N_14294);
nor U15450 (N_15450,N_13678,N_13603);
and U15451 (N_15451,N_14044,N_14286);
or U15452 (N_15452,N_14142,N_14278);
and U15453 (N_15453,N_14392,N_13887);
nand U15454 (N_15454,N_13598,N_14300);
nand U15455 (N_15455,N_13248,N_13683);
nand U15456 (N_15456,N_13440,N_13847);
and U15457 (N_15457,N_13990,N_14145);
or U15458 (N_15458,N_13312,N_13281);
nor U15459 (N_15459,N_13614,N_14265);
xor U15460 (N_15460,N_14053,N_14085);
xnor U15461 (N_15461,N_13742,N_14216);
nor U15462 (N_15462,N_13313,N_13239);
nand U15463 (N_15463,N_14377,N_13709);
and U15464 (N_15464,N_13374,N_14293);
nor U15465 (N_15465,N_13378,N_14093);
and U15466 (N_15466,N_13920,N_13969);
nor U15467 (N_15467,N_14365,N_13268);
and U15468 (N_15468,N_14267,N_14192);
nand U15469 (N_15469,N_14279,N_13370);
nor U15470 (N_15470,N_13467,N_13855);
xnor U15471 (N_15471,N_13948,N_14101);
nand U15472 (N_15472,N_14351,N_13797);
nand U15473 (N_15473,N_14283,N_14233);
nor U15474 (N_15474,N_13213,N_14272);
nor U15475 (N_15475,N_13982,N_14185);
and U15476 (N_15476,N_13246,N_13937);
or U15477 (N_15477,N_13580,N_13238);
nor U15478 (N_15478,N_13357,N_14112);
or U15479 (N_15479,N_14174,N_14033);
and U15480 (N_15480,N_14375,N_13360);
and U15481 (N_15481,N_13550,N_13910);
xnor U15482 (N_15482,N_13975,N_13588);
nor U15483 (N_15483,N_13814,N_13877);
xnor U15484 (N_15484,N_13287,N_13310);
and U15485 (N_15485,N_13529,N_13569);
or U15486 (N_15486,N_13832,N_13548);
xor U15487 (N_15487,N_13775,N_13327);
and U15488 (N_15488,N_13659,N_13820);
and U15489 (N_15489,N_13399,N_13341);
and U15490 (N_15490,N_14213,N_13327);
nor U15491 (N_15491,N_14266,N_13756);
xor U15492 (N_15492,N_13398,N_13504);
or U15493 (N_15493,N_14386,N_13230);
nand U15494 (N_15494,N_13552,N_13617);
or U15495 (N_15495,N_13243,N_13672);
or U15496 (N_15496,N_13768,N_14358);
nor U15497 (N_15497,N_13762,N_13416);
or U15498 (N_15498,N_13341,N_13241);
or U15499 (N_15499,N_14073,N_13418);
nand U15500 (N_15500,N_13425,N_14043);
or U15501 (N_15501,N_13514,N_13889);
or U15502 (N_15502,N_13621,N_13654);
nand U15503 (N_15503,N_14225,N_13810);
nand U15504 (N_15504,N_14177,N_13564);
and U15505 (N_15505,N_13676,N_14156);
xor U15506 (N_15506,N_13602,N_13500);
nand U15507 (N_15507,N_13255,N_13896);
and U15508 (N_15508,N_14187,N_13648);
nand U15509 (N_15509,N_13469,N_13298);
nor U15510 (N_15510,N_13744,N_14162);
nand U15511 (N_15511,N_13316,N_14235);
or U15512 (N_15512,N_13688,N_13925);
nor U15513 (N_15513,N_13807,N_13488);
nand U15514 (N_15514,N_13987,N_14207);
nor U15515 (N_15515,N_13881,N_13403);
and U15516 (N_15516,N_13221,N_13302);
or U15517 (N_15517,N_14371,N_13671);
nor U15518 (N_15518,N_13440,N_14206);
and U15519 (N_15519,N_13593,N_13839);
nand U15520 (N_15520,N_13871,N_13501);
nor U15521 (N_15521,N_13820,N_14246);
nor U15522 (N_15522,N_13310,N_13911);
or U15523 (N_15523,N_14376,N_13534);
xor U15524 (N_15524,N_13780,N_14177);
or U15525 (N_15525,N_13701,N_13743);
or U15526 (N_15526,N_13933,N_14394);
and U15527 (N_15527,N_14197,N_13402);
or U15528 (N_15528,N_13388,N_13302);
xor U15529 (N_15529,N_13909,N_13983);
nor U15530 (N_15530,N_14199,N_13466);
and U15531 (N_15531,N_14137,N_14241);
or U15532 (N_15532,N_13697,N_13501);
and U15533 (N_15533,N_13549,N_13644);
xor U15534 (N_15534,N_13593,N_14210);
or U15535 (N_15535,N_13318,N_13275);
and U15536 (N_15536,N_13724,N_14224);
nor U15537 (N_15537,N_13950,N_13235);
and U15538 (N_15538,N_14270,N_14254);
and U15539 (N_15539,N_14254,N_13464);
nor U15540 (N_15540,N_14048,N_14371);
nor U15541 (N_15541,N_13806,N_13745);
nand U15542 (N_15542,N_13745,N_13546);
xnor U15543 (N_15543,N_13451,N_13794);
xnor U15544 (N_15544,N_14018,N_14082);
xor U15545 (N_15545,N_13360,N_13766);
xnor U15546 (N_15546,N_14299,N_13635);
and U15547 (N_15547,N_14025,N_13992);
and U15548 (N_15548,N_13602,N_14164);
or U15549 (N_15549,N_13836,N_13531);
or U15550 (N_15550,N_13901,N_13774);
nand U15551 (N_15551,N_13872,N_13699);
xor U15552 (N_15552,N_13372,N_14173);
and U15553 (N_15553,N_14283,N_13696);
nor U15554 (N_15554,N_13383,N_13703);
xnor U15555 (N_15555,N_13699,N_13364);
or U15556 (N_15556,N_14361,N_13934);
nor U15557 (N_15557,N_14254,N_13633);
or U15558 (N_15558,N_13791,N_13931);
nand U15559 (N_15559,N_13903,N_14129);
and U15560 (N_15560,N_13451,N_13430);
and U15561 (N_15561,N_13841,N_13441);
xor U15562 (N_15562,N_14131,N_13306);
xnor U15563 (N_15563,N_14180,N_13288);
xnor U15564 (N_15564,N_13251,N_13956);
nand U15565 (N_15565,N_14159,N_13248);
nand U15566 (N_15566,N_14070,N_13566);
or U15567 (N_15567,N_13949,N_13386);
or U15568 (N_15568,N_14050,N_13450);
or U15569 (N_15569,N_13920,N_13327);
nor U15570 (N_15570,N_13683,N_13805);
or U15571 (N_15571,N_13749,N_13320);
and U15572 (N_15572,N_14234,N_14271);
xor U15573 (N_15573,N_13547,N_14131);
and U15574 (N_15574,N_13835,N_14267);
nand U15575 (N_15575,N_14255,N_14153);
and U15576 (N_15576,N_13225,N_13630);
xor U15577 (N_15577,N_13624,N_14243);
and U15578 (N_15578,N_14151,N_13467);
or U15579 (N_15579,N_13932,N_13799);
xor U15580 (N_15580,N_14357,N_13783);
and U15581 (N_15581,N_13244,N_13278);
xnor U15582 (N_15582,N_13859,N_13287);
or U15583 (N_15583,N_14179,N_13890);
and U15584 (N_15584,N_14295,N_13804);
and U15585 (N_15585,N_13426,N_13412);
or U15586 (N_15586,N_13333,N_13925);
nor U15587 (N_15587,N_13846,N_13514);
and U15588 (N_15588,N_13828,N_13327);
nor U15589 (N_15589,N_13847,N_13764);
and U15590 (N_15590,N_14309,N_13808);
xnor U15591 (N_15591,N_13577,N_14039);
nor U15592 (N_15592,N_13639,N_14298);
and U15593 (N_15593,N_13922,N_13870);
xnor U15594 (N_15594,N_13454,N_13761);
and U15595 (N_15595,N_14282,N_13816);
nand U15596 (N_15596,N_14375,N_14352);
nand U15597 (N_15597,N_13243,N_13571);
nor U15598 (N_15598,N_13840,N_14076);
or U15599 (N_15599,N_13673,N_13228);
nor U15600 (N_15600,N_15127,N_14787);
nand U15601 (N_15601,N_14894,N_14730);
nand U15602 (N_15602,N_15391,N_15599);
or U15603 (N_15603,N_15445,N_15207);
nor U15604 (N_15604,N_15189,N_14904);
or U15605 (N_15605,N_14648,N_15296);
nand U15606 (N_15606,N_14589,N_14825);
xnor U15607 (N_15607,N_15508,N_15437);
or U15608 (N_15608,N_14429,N_15527);
xnor U15609 (N_15609,N_15455,N_15151);
or U15610 (N_15610,N_14609,N_14569);
nor U15611 (N_15611,N_15278,N_14536);
nand U15612 (N_15612,N_14942,N_15359);
nor U15613 (N_15613,N_15308,N_15261);
and U15614 (N_15614,N_14434,N_15317);
xor U15615 (N_15615,N_15130,N_14982);
xnor U15616 (N_15616,N_15526,N_14956);
xor U15617 (N_15617,N_14987,N_15371);
or U15618 (N_15618,N_14647,N_14808);
xnor U15619 (N_15619,N_15260,N_14509);
and U15620 (N_15620,N_15262,N_15223);
xnor U15621 (N_15621,N_15511,N_14916);
xnor U15622 (N_15622,N_14959,N_15501);
and U15623 (N_15623,N_15123,N_14439);
xor U15624 (N_15624,N_14506,N_15072);
and U15625 (N_15625,N_14793,N_15341);
nand U15626 (N_15626,N_14641,N_15494);
nand U15627 (N_15627,N_15576,N_14917);
nor U15628 (N_15628,N_14535,N_15280);
xor U15629 (N_15629,N_15333,N_14731);
and U15630 (N_15630,N_15517,N_15214);
and U15631 (N_15631,N_14546,N_15303);
xor U15632 (N_15632,N_15139,N_14813);
nand U15633 (N_15633,N_14636,N_15178);
nor U15634 (N_15634,N_14447,N_15361);
nor U15635 (N_15635,N_14412,N_14550);
xnor U15636 (N_15636,N_15101,N_14596);
and U15637 (N_15637,N_15003,N_15297);
or U15638 (N_15638,N_14737,N_14865);
nand U15639 (N_15639,N_15363,N_15227);
and U15640 (N_15640,N_14833,N_14419);
nor U15641 (N_15641,N_14459,N_14965);
xnor U15642 (N_15642,N_15555,N_14992);
xor U15643 (N_15643,N_14911,N_15345);
or U15644 (N_15644,N_14574,N_14836);
and U15645 (N_15645,N_15109,N_14415);
xor U15646 (N_15646,N_15427,N_14954);
xnor U15647 (N_15647,N_14462,N_14504);
nand U15648 (N_15648,N_15150,N_14537);
nand U15649 (N_15649,N_15183,N_15116);
nand U15650 (N_15650,N_14963,N_14642);
xnor U15651 (N_15651,N_14771,N_14719);
nor U15652 (N_15652,N_15406,N_14879);
or U15653 (N_15653,N_14762,N_14923);
xor U15654 (N_15654,N_14875,N_14856);
nand U15655 (N_15655,N_15336,N_15170);
or U15656 (N_15656,N_15018,N_14699);
or U15657 (N_15657,N_14926,N_15167);
or U15658 (N_15658,N_15131,N_14500);
xor U15659 (N_15659,N_15563,N_14665);
nand U15660 (N_15660,N_14756,N_15186);
nor U15661 (N_15661,N_15153,N_15006);
xor U15662 (N_15662,N_15162,N_14708);
or U15663 (N_15663,N_15039,N_15340);
or U15664 (N_15664,N_14616,N_14451);
or U15665 (N_15665,N_15114,N_15536);
or U15666 (N_15666,N_14639,N_14860);
xor U15667 (N_15667,N_15430,N_14886);
or U15668 (N_15668,N_15082,N_15379);
or U15669 (N_15669,N_14423,N_14652);
nor U15670 (N_15670,N_15537,N_15273);
nand U15671 (N_15671,N_15103,N_15370);
nor U15672 (N_15672,N_14581,N_14850);
nand U15673 (N_15673,N_14832,N_14874);
nor U15674 (N_15674,N_15196,N_14814);
nand U15675 (N_15675,N_15444,N_15432);
nand U15676 (N_15676,N_14921,N_14409);
and U15677 (N_15677,N_14725,N_15401);
nor U15678 (N_15678,N_14945,N_14547);
and U15679 (N_15679,N_14918,N_15257);
or U15680 (N_15680,N_15433,N_14576);
nor U15681 (N_15681,N_14656,N_14745);
nand U15682 (N_15682,N_15144,N_14818);
nand U15683 (N_15683,N_14599,N_15202);
xor U15684 (N_15684,N_14908,N_15120);
nand U15685 (N_15685,N_14826,N_15276);
xnor U15686 (N_15686,N_14678,N_15334);
xnor U15687 (N_15687,N_14852,N_15512);
and U15688 (N_15688,N_14655,N_14951);
and U15689 (N_15689,N_15031,N_15483);
or U15690 (N_15690,N_14407,N_15272);
and U15691 (N_15691,N_14883,N_15442);
nor U15692 (N_15692,N_14948,N_15480);
xnor U15693 (N_15693,N_15215,N_14566);
nor U15694 (N_15694,N_14915,N_15330);
nand U15695 (N_15695,N_14897,N_14796);
nand U15696 (N_15696,N_14455,N_15023);
and U15697 (N_15697,N_15395,N_14677);
nor U15698 (N_15698,N_14727,N_15008);
nand U15699 (N_15699,N_15165,N_15241);
and U15700 (N_15700,N_14501,N_14659);
nand U15701 (N_15701,N_15492,N_15212);
nor U15702 (N_15702,N_15115,N_15270);
xnor U15703 (N_15703,N_15233,N_15424);
or U15704 (N_15704,N_15594,N_15047);
and U15705 (N_15705,N_15365,N_15259);
or U15706 (N_15706,N_14533,N_15035);
and U15707 (N_15707,N_14595,N_15493);
and U15708 (N_15708,N_15052,N_14700);
and U15709 (N_15709,N_14687,N_15528);
and U15710 (N_15710,N_15096,N_14611);
or U15711 (N_15711,N_14681,N_14411);
nand U15712 (N_15712,N_14843,N_14543);
nor U15713 (N_15713,N_14950,N_14529);
or U15714 (N_15714,N_15568,N_15429);
nand U15715 (N_15715,N_14770,N_14910);
nor U15716 (N_15716,N_15454,N_14792);
nand U15717 (N_15717,N_15590,N_15347);
xor U15718 (N_15718,N_15304,N_14585);
or U15719 (N_15719,N_14811,N_14711);
or U15720 (N_15720,N_14736,N_15598);
and U15721 (N_15721,N_15258,N_15204);
or U15722 (N_15722,N_15463,N_15591);
or U15723 (N_15723,N_15218,N_14458);
xor U15724 (N_15724,N_14943,N_15025);
or U15725 (N_15725,N_15390,N_15095);
or U15726 (N_15726,N_15350,N_14572);
nand U15727 (N_15727,N_14588,N_14885);
or U15728 (N_15728,N_14619,N_15058);
nand U15729 (N_15729,N_14929,N_15172);
xnor U15730 (N_15730,N_15473,N_14754);
or U15731 (N_15731,N_15174,N_14804);
or U15732 (N_15732,N_14488,N_14735);
nand U15733 (N_15733,N_15410,N_14512);
nand U15734 (N_15734,N_14782,N_14510);
nor U15735 (N_15735,N_15292,N_15344);
or U15736 (N_15736,N_14601,N_15486);
xnor U15737 (N_15737,N_14823,N_15168);
nand U15738 (N_15738,N_15519,N_15074);
nand U15739 (N_15739,N_14666,N_14763);
nor U15740 (N_15740,N_15251,N_15237);
and U15741 (N_15741,N_15245,N_15065);
or U15742 (N_15742,N_15305,N_15017);
nand U15743 (N_15743,N_15135,N_14888);
xor U15744 (N_15744,N_15325,N_14542);
or U15745 (N_15745,N_15085,N_14706);
nand U15746 (N_15746,N_15431,N_14957);
nor U15747 (N_15747,N_15570,N_14769);
and U15748 (N_15748,N_15099,N_15573);
and U15749 (N_15749,N_14734,N_14723);
xnor U15750 (N_15750,N_14752,N_15489);
nor U15751 (N_15751,N_14819,N_14822);
nor U15752 (N_15752,N_14671,N_15435);
nor U15753 (N_15753,N_14967,N_14788);
xnor U15754 (N_15754,N_15213,N_14695);
or U15755 (N_15755,N_14739,N_15324);
xnor U15756 (N_15756,N_15319,N_14985);
and U15757 (N_15757,N_15554,N_14562);
nor U15758 (N_15758,N_14774,N_15546);
nor U15759 (N_15759,N_15574,N_15515);
xor U15760 (N_15760,N_14805,N_14777);
or U15761 (N_15761,N_14870,N_14976);
nand U15762 (N_15762,N_14548,N_15263);
nor U15763 (N_15763,N_14980,N_14496);
xor U15764 (N_15764,N_14552,N_14520);
and U15765 (N_15765,N_15053,N_14930);
nor U15766 (N_15766,N_14851,N_15453);
nand U15767 (N_15767,N_15077,N_15523);
nand U15768 (N_15768,N_15316,N_15136);
nand U15769 (N_15769,N_15412,N_14584);
and U15770 (N_15770,N_14797,N_14847);
and U15771 (N_15771,N_14807,N_14620);
nand U15772 (N_15772,N_15567,N_14604);
nand U15773 (N_15773,N_14768,N_14773);
and U15774 (N_15774,N_15503,N_15446);
nor U15775 (N_15775,N_14765,N_14485);
nor U15776 (N_15776,N_14997,N_15256);
nand U15777 (N_15777,N_14617,N_14709);
or U15778 (N_15778,N_15155,N_15373);
nand U15779 (N_15779,N_15119,N_14848);
and U15780 (N_15780,N_15143,N_15206);
and U15781 (N_15781,N_15028,N_15211);
nand U15782 (N_15782,N_14443,N_14523);
or U15783 (N_15783,N_14448,N_15240);
and U15784 (N_15784,N_14564,N_14891);
xor U15785 (N_15785,N_15219,N_15529);
nor U15786 (N_15786,N_14484,N_15128);
nor U15787 (N_15787,N_15425,N_15271);
xor U15788 (N_15788,N_14514,N_15556);
xor U15789 (N_15789,N_14909,N_14486);
or U15790 (N_15790,N_15073,N_14670);
nor U15791 (N_15791,N_15420,N_15071);
and U15792 (N_15792,N_14772,N_15352);
xor U15793 (N_15793,N_15593,N_15022);
and U15794 (N_15794,N_14863,N_14622);
xnor U15795 (N_15795,N_15383,N_14563);
or U15796 (N_15796,N_15548,N_15544);
nor U15797 (N_15797,N_15088,N_14638);
nand U15798 (N_15798,N_15339,N_14603);
xnor U15799 (N_15799,N_15138,N_15440);
and U15800 (N_15800,N_15147,N_15266);
nor U15801 (N_15801,N_15531,N_14473);
and U15802 (N_15802,N_15107,N_15002);
nor U15803 (N_15803,N_15291,N_14544);
or U15804 (N_15804,N_14612,N_14789);
and U15805 (N_15805,N_15315,N_15354);
and U15806 (N_15806,N_15397,N_15279);
nand U15807 (N_15807,N_15329,N_14714);
and U15808 (N_15808,N_15045,N_14966);
nand U15809 (N_15809,N_15498,N_14645);
or U15810 (N_15810,N_15566,N_15318);
nand U15811 (N_15811,N_15495,N_14471);
nor U15812 (N_15812,N_15274,N_14962);
xor U15813 (N_15813,N_15331,N_15530);
nor U15814 (N_15814,N_14990,N_15436);
nor U15815 (N_15815,N_15122,N_15580);
nand U15816 (N_15816,N_14508,N_14416);
nand U15817 (N_15817,N_14437,N_15166);
or U15818 (N_15818,N_14607,N_15385);
nand U15819 (N_15819,N_14880,N_14949);
nor U15820 (N_15820,N_14895,N_15220);
xnor U15821 (N_15821,N_15060,N_15389);
nand U15822 (N_15822,N_15061,N_14668);
or U15823 (N_15823,N_15479,N_14593);
nand U15824 (N_15824,N_14854,N_15076);
nand U15825 (N_15825,N_14890,N_14554);
nor U15826 (N_15826,N_15141,N_14482);
nor U15827 (N_15827,N_14912,N_14786);
xor U15828 (N_15828,N_15541,N_14442);
xor U15829 (N_15829,N_15532,N_15111);
nor U15830 (N_15830,N_15094,N_15137);
nor U15831 (N_15831,N_14503,N_14449);
and U15832 (N_15832,N_14869,N_14927);
or U15833 (N_15833,N_15295,N_14707);
nor U15834 (N_15834,N_15046,N_14806);
nand U15835 (N_15835,N_14624,N_14436);
nand U15836 (N_15836,N_14901,N_15221);
and U15837 (N_15837,N_15408,N_14696);
and U15838 (N_15838,N_15294,N_15374);
or U15839 (N_15839,N_15441,N_14534);
nor U15840 (N_15840,N_15507,N_14682);
nor U15841 (N_15841,N_15024,N_14791);
or U15842 (N_15842,N_15110,N_15396);
and U15843 (N_15843,N_15393,N_15496);
nor U15844 (N_15844,N_14937,N_15067);
and U15845 (N_15845,N_14802,N_14483);
xnor U15846 (N_15846,N_15521,N_15449);
nand U15847 (N_15847,N_15367,N_15327);
nor U15848 (N_15848,N_15014,N_15553);
or U15849 (N_15849,N_15264,N_14887);
or U15850 (N_15850,N_14685,N_15232);
nor U15851 (N_15851,N_14582,N_15514);
nand U15852 (N_15852,N_14560,N_14519);
xor U15853 (N_15853,N_15000,N_15392);
or U15854 (N_15854,N_15175,N_14644);
and U15855 (N_15855,N_15542,N_15267);
and U15856 (N_15856,N_15098,N_14672);
or U15857 (N_15857,N_14633,N_15252);
nor U15858 (N_15858,N_14575,N_15439);
and U15859 (N_15859,N_15062,N_15070);
or U15860 (N_15860,N_15015,N_15021);
nand U15861 (N_15861,N_15417,N_14984);
xor U15862 (N_15862,N_15364,N_14871);
nor U15863 (N_15863,N_14433,N_15118);
or U15864 (N_15864,N_14914,N_15129);
nor U15865 (N_15865,N_15581,N_14651);
or U15866 (N_15866,N_14868,N_15197);
nor U15867 (N_15867,N_15328,N_14898);
xor U15868 (N_15868,N_14830,N_15589);
or U15869 (N_15869,N_14615,N_15375);
or U15870 (N_15870,N_15321,N_15466);
xnor U15871 (N_15871,N_14474,N_14540);
nand U15872 (N_15872,N_14749,N_15100);
or U15873 (N_15873,N_14872,N_15491);
nor U15874 (N_15874,N_15461,N_14801);
and U15875 (N_15875,N_14996,N_14750);
xor U15876 (N_15876,N_15090,N_14663);
xor U15877 (N_15877,N_14691,N_14515);
or U15878 (N_15878,N_14861,N_14968);
nand U15879 (N_15879,N_15476,N_14628);
nand U15880 (N_15880,N_14470,N_15368);
nor U15881 (N_15881,N_14972,N_15048);
and U15882 (N_15882,N_15578,N_14521);
nor U15883 (N_15883,N_14590,N_15587);
nand U15884 (N_15884,N_14518,N_15465);
xnor U15885 (N_15885,N_15369,N_14946);
or U15886 (N_15886,N_14829,N_14559);
or U15887 (N_15887,N_14664,N_14775);
or U15888 (N_15888,N_15203,N_15434);
nand U15889 (N_15889,N_14551,N_14413);
and U15890 (N_15890,N_14827,N_15419);
nand U15891 (N_15891,N_14605,N_14790);
xor U15892 (N_15892,N_15038,N_15012);
nand U15893 (N_15893,N_15386,N_15343);
or U15894 (N_15894,N_15113,N_15055);
xor U15895 (N_15895,N_15475,N_14757);
nand U15896 (N_15896,N_15231,N_14837);
xor U15897 (N_15897,N_15459,N_14936);
nor U15898 (N_15898,N_14408,N_14922);
xor U15899 (N_15899,N_15510,N_15450);
nand U15900 (N_15900,N_14674,N_14755);
nor U15901 (N_15901,N_15299,N_15400);
or U15902 (N_15902,N_15372,N_14689);
xnor U15903 (N_15903,N_15524,N_14631);
xor U15904 (N_15904,N_15505,N_15106);
xor U15905 (N_15905,N_14993,N_15269);
nand U15906 (N_15906,N_14776,N_15583);
or U15907 (N_15907,N_14899,N_15195);
nor U15908 (N_15908,N_14643,N_14417);
nor U15909 (N_15909,N_15380,N_15290);
nand U15910 (N_15910,N_15353,N_15335);
nor U15911 (N_15911,N_14487,N_15288);
or U15912 (N_15912,N_14799,N_15187);
nor U15913 (N_15913,N_15588,N_15201);
and U15914 (N_15914,N_15585,N_15500);
xor U15915 (N_15915,N_14919,N_15457);
and U15916 (N_15916,N_15163,N_15081);
xor U15917 (N_15917,N_15481,N_15597);
nand U15918 (N_15918,N_14586,N_14613);
and U15919 (N_15919,N_14903,N_15447);
nand U15920 (N_15920,N_14466,N_14857);
xnor U15921 (N_15921,N_15152,N_15286);
xnor U15922 (N_15922,N_15504,N_14452);
nand U15923 (N_15923,N_15133,N_14953);
or U15924 (N_15924,N_15312,N_15477);
and U15925 (N_15925,N_15117,N_14958);
and U15926 (N_15926,N_14427,N_14673);
and U15927 (N_15927,N_15009,N_15171);
nand U15928 (N_15928,N_14640,N_14545);
nand U15929 (N_15929,N_14809,N_15007);
xor U15930 (N_15930,N_15044,N_15205);
nand U15931 (N_15931,N_14401,N_14421);
and U15932 (N_15932,N_14573,N_14658);
and U15933 (N_15933,N_14630,N_14472);
and U15934 (N_15934,N_15423,N_14810);
or U15935 (N_15935,N_15157,N_15194);
nor U15936 (N_15936,N_15236,N_15191);
xnor U15937 (N_15937,N_15019,N_15066);
nor U15938 (N_15938,N_14438,N_14753);
or U15939 (N_15939,N_15284,N_14705);
xnor U15940 (N_15940,N_15485,N_15049);
xnor U15941 (N_15941,N_15337,N_15356);
nor U15942 (N_15942,N_15443,N_15471);
nor U15943 (N_15943,N_15487,N_14492);
and U15944 (N_15944,N_14414,N_14974);
nor U15945 (N_15945,N_14717,N_14446);
nand U15946 (N_15946,N_14866,N_15360);
and U15947 (N_15947,N_15228,N_14410);
or U15948 (N_15948,N_14979,N_15474);
or U15949 (N_15949,N_14499,N_15407);
xor U15950 (N_15950,N_15346,N_15125);
nand U15951 (N_15951,N_14977,N_14692);
and U15952 (N_15952,N_14679,N_14680);
xnor U15953 (N_15953,N_15411,N_14568);
and U15954 (N_15954,N_15216,N_14481);
nand U15955 (N_15955,N_15399,N_14460);
or U15956 (N_15956,N_15582,N_15161);
nor U15957 (N_15957,N_15042,N_14742);
xnor U15958 (N_15958,N_15253,N_15464);
nand U15959 (N_15959,N_14565,N_15293);
nor U15960 (N_15960,N_14587,N_14635);
nand U15961 (N_15961,N_15016,N_14513);
or U15962 (N_15962,N_15230,N_15059);
nand U15963 (N_15963,N_15239,N_15323);
nand U15964 (N_15964,N_15063,N_14713);
nand U15965 (N_15965,N_14924,N_14457);
or U15966 (N_15966,N_15289,N_14718);
or U15967 (N_15967,N_15121,N_15032);
or U15968 (N_15968,N_14732,N_15033);
xnor U15969 (N_15969,N_15409,N_14539);
nand U15970 (N_15970,N_15394,N_15518);
xnor U15971 (N_15971,N_14567,N_14722);
nor U15972 (N_15972,N_15547,N_15357);
nand U15973 (N_15973,N_15254,N_14973);
nor U15974 (N_15974,N_15078,N_14669);
nor U15975 (N_15975,N_15285,N_14900);
xnor U15976 (N_15976,N_14441,N_14431);
or U15977 (N_15977,N_15093,N_15247);
xnor U15978 (N_15978,N_15404,N_14400);
nand U15979 (N_15979,N_14743,N_15322);
nand U15980 (N_15980,N_14600,N_14420);
xor U15981 (N_15981,N_15525,N_15132);
xor U15982 (N_15982,N_14527,N_15338);
or U15983 (N_15983,N_15562,N_15506);
nor U15984 (N_15984,N_14815,N_14906);
nor U15985 (N_15985,N_15248,N_15124);
or U15986 (N_15986,N_14698,N_15142);
xor U15987 (N_15987,N_15456,N_15079);
and U15988 (N_15988,N_14989,N_14444);
or U15989 (N_15989,N_15484,N_15190);
nor U15990 (N_15990,N_14784,N_15438);
xnor U15991 (N_15991,N_14970,N_14932);
nor U15992 (N_15992,N_14779,N_15467);
xor U15993 (N_15993,N_15382,N_15559);
or U15994 (N_15994,N_14940,N_14944);
xnor U15995 (N_15995,N_15413,N_14928);
nor U15996 (N_15996,N_14876,N_14969);
or U15997 (N_15997,N_15560,N_14741);
or U15998 (N_15998,N_14728,N_15134);
or U15999 (N_15999,N_15056,N_15243);
or U16000 (N_16000,N_15180,N_14740);
nand U16001 (N_16001,N_14627,N_15040);
xnor U16002 (N_16002,N_15080,N_15298);
and U16003 (N_16003,N_14526,N_14841);
xnor U16004 (N_16004,N_15185,N_15540);
and U16005 (N_16005,N_14798,N_14862);
or U16006 (N_16006,N_14964,N_15179);
xor U16007 (N_16007,N_14435,N_15550);
or U16008 (N_16008,N_14694,N_14817);
or U16009 (N_16009,N_14450,N_15358);
nor U16010 (N_16010,N_14858,N_15287);
or U16011 (N_16011,N_15545,N_14594);
nor U16012 (N_16012,N_14637,N_14701);
xnor U16013 (N_16013,N_15149,N_15020);
nor U16014 (N_16014,N_14491,N_14597);
nand U16015 (N_16015,N_15029,N_14878);
nor U16016 (N_16016,N_15310,N_14555);
and U16017 (N_16017,N_14816,N_14978);
xor U16018 (N_16018,N_14893,N_14842);
or U16019 (N_16019,N_14626,N_15307);
xor U16020 (N_16020,N_15558,N_15234);
or U16021 (N_16021,N_14729,N_15577);
and U16022 (N_16022,N_15277,N_15092);
and U16023 (N_16023,N_14661,N_14889);
xnor U16024 (N_16024,N_14426,N_14432);
nand U16025 (N_16025,N_15217,N_14835);
nand U16026 (N_16026,N_15126,N_14955);
or U16027 (N_16027,N_15198,N_14598);
or U16028 (N_16028,N_14580,N_15268);
nand U16029 (N_16029,N_15458,N_15229);
nor U16030 (N_16030,N_14583,N_15146);
nor U16031 (N_16031,N_14475,N_15366);
and U16032 (N_16032,N_14592,N_14676);
nand U16033 (N_16033,N_14538,N_14994);
nor U16034 (N_16034,N_14961,N_14995);
and U16035 (N_16035,N_15027,N_15104);
and U16036 (N_16036,N_15572,N_14505);
nand U16037 (N_16037,N_15381,N_14553);
xnor U16038 (N_16038,N_15516,N_14716);
xnor U16039 (N_16039,N_14941,N_15102);
nand U16040 (N_16040,N_15154,N_15314);
or U16041 (N_16041,N_14490,N_15472);
or U16042 (N_16042,N_15034,N_15300);
and U16043 (N_16043,N_15428,N_14532);
xor U16044 (N_16044,N_15342,N_14760);
xnor U16045 (N_16045,N_15502,N_14498);
nand U16046 (N_16046,N_14690,N_15188);
and U16047 (N_16047,N_15557,N_15509);
or U16048 (N_16048,N_14845,N_15398);
nor U16049 (N_16049,N_14812,N_14502);
or U16050 (N_16050,N_14577,N_14783);
xnor U16051 (N_16051,N_14465,N_15415);
nor U16052 (N_16052,N_14758,N_14884);
or U16053 (N_16053,N_14947,N_15037);
xnor U16054 (N_16054,N_15140,N_14516);
nand U16055 (N_16055,N_15148,N_14720);
and U16056 (N_16056,N_15470,N_15520);
and U16057 (N_16057,N_15311,N_14934);
and U16058 (N_16058,N_15199,N_14522);
and U16059 (N_16059,N_15565,N_15160);
nor U16060 (N_16060,N_14864,N_14618);
nor U16061 (N_16061,N_14430,N_14913);
and U16062 (N_16062,N_15208,N_14873);
nand U16063 (N_16063,N_14726,N_15426);
xnor U16064 (N_16064,N_14881,N_14902);
nand U16065 (N_16065,N_15387,N_14999);
nor U16066 (N_16066,N_15448,N_15586);
and U16067 (N_16067,N_15283,N_15050);
nor U16068 (N_16068,N_15086,N_14489);
or U16069 (N_16069,N_14952,N_14998);
nand U16070 (N_16070,N_14767,N_15482);
xor U16071 (N_16071,N_15173,N_15535);
xnor U16072 (N_16072,N_14625,N_14780);
or U16073 (N_16073,N_14761,N_14724);
and U16074 (N_16074,N_15156,N_14528);
xnor U16075 (N_16075,N_14803,N_14463);
or U16076 (N_16076,N_14759,N_14855);
or U16077 (N_16077,N_14404,N_14892);
nand U16078 (N_16078,N_14800,N_14834);
or U16079 (N_16079,N_15112,N_14991);
and U16080 (N_16080,N_14853,N_14424);
xor U16081 (N_16081,N_15376,N_14703);
xor U16082 (N_16082,N_14988,N_15348);
and U16083 (N_16083,N_14606,N_15549);
nor U16084 (N_16084,N_15224,N_14556);
or U16085 (N_16085,N_15301,N_14778);
nor U16086 (N_16086,N_14525,N_15384);
or U16087 (N_16087,N_15320,N_15054);
nor U16088 (N_16088,N_14684,N_15158);
nor U16089 (N_16089,N_14738,N_15418);
and U16090 (N_16090,N_15051,N_15192);
and U16091 (N_16091,N_14697,N_14610);
or U16092 (N_16092,N_14667,N_15083);
xor U16093 (N_16093,N_14907,N_15378);
xor U16094 (N_16094,N_15250,N_14517);
xnor U16095 (N_16095,N_15026,N_15226);
and U16096 (N_16096,N_15362,N_14428);
xor U16097 (N_16097,N_14785,N_14495);
and U16098 (N_16098,N_14712,N_14896);
nor U16099 (N_16099,N_14933,N_14831);
nor U16100 (N_16100,N_15057,N_14747);
and U16101 (N_16101,N_15488,N_14846);
and U16102 (N_16102,N_14493,N_14454);
or U16103 (N_16103,N_14981,N_14480);
and U16104 (N_16104,N_14425,N_15200);
and U16105 (N_16105,N_14925,N_14766);
or U16106 (N_16106,N_15451,N_14721);
nor U16107 (N_16107,N_15235,N_15182);
and U16108 (N_16108,N_14561,N_15468);
nand U16109 (N_16109,N_15043,N_15422);
xor U16110 (N_16110,N_14507,N_15238);
xor U16111 (N_16111,N_14675,N_14541);
xor U16112 (N_16112,N_15177,N_15209);
xnor U16113 (N_16113,N_15564,N_15571);
xor U16114 (N_16114,N_15497,N_14821);
or U16115 (N_16115,N_14828,N_15533);
xnor U16116 (N_16116,N_14477,N_14975);
nor U16117 (N_16117,N_14653,N_15579);
nand U16118 (N_16118,N_14905,N_15036);
or U16119 (N_16119,N_15569,N_14764);
or U16120 (N_16120,N_14478,N_14549);
or U16121 (N_16121,N_15105,N_15469);
and U16122 (N_16122,N_14558,N_14602);
xor U16123 (N_16123,N_14662,N_15064);
or U16124 (N_16124,N_15462,N_14467);
and U16125 (N_16125,N_15164,N_15551);
or U16126 (N_16126,N_14931,N_15265);
nand U16127 (N_16127,N_14971,N_15089);
nand U16128 (N_16128,N_14654,N_15539);
nor U16129 (N_16129,N_14571,N_14748);
nor U16130 (N_16130,N_14751,N_14795);
nor U16131 (N_16131,N_14578,N_15403);
and U16132 (N_16132,N_15041,N_15005);
nand U16133 (N_16133,N_15306,N_15210);
nand U16134 (N_16134,N_15242,N_14461);
or U16135 (N_16135,N_15452,N_15302);
nand U16136 (N_16136,N_15313,N_15499);
and U16137 (N_16137,N_14794,N_15004);
nor U16138 (N_16138,N_15181,N_14511);
and U16139 (N_16139,N_15249,N_15075);
and U16140 (N_16140,N_14524,N_15534);
nor U16141 (N_16141,N_15169,N_15222);
xnor U16142 (N_16142,N_14838,N_14986);
xnor U16143 (N_16143,N_14849,N_15108);
and U16144 (N_16144,N_14468,N_14479);
nand U16145 (N_16145,N_15478,N_15282);
and U16146 (N_16146,N_15377,N_14882);
and U16147 (N_16147,N_14744,N_15460);
nor U16148 (N_16148,N_14418,N_15584);
and U16149 (N_16149,N_14456,N_14646);
nor U16150 (N_16150,N_14440,N_15030);
nand U16151 (N_16151,N_14939,N_15159);
xnor U16152 (N_16152,N_15091,N_15275);
nor U16153 (N_16153,N_14938,N_14715);
nor U16154 (N_16154,N_14464,N_15355);
xor U16155 (N_16155,N_15176,N_15001);
xor U16156 (N_16156,N_14608,N_15575);
nor U16157 (N_16157,N_15087,N_14557);
nor U16158 (N_16158,N_14683,N_15013);
and U16159 (N_16159,N_14704,N_15010);
xnor U16160 (N_16160,N_15405,N_14445);
or U16161 (N_16161,N_15552,N_14820);
nand U16162 (N_16162,N_14710,N_14530);
nor U16163 (N_16163,N_15490,N_15193);
nand U16164 (N_16164,N_14453,N_14824);
or U16165 (N_16165,N_14403,N_14983);
nor U16166 (N_16166,N_14494,N_14629);
nor U16167 (N_16167,N_15351,N_15244);
or U16168 (N_16168,N_14591,N_15011);
xor U16169 (N_16169,N_14650,N_14632);
or U16170 (N_16170,N_14840,N_14702);
nor U16171 (N_16171,N_14688,N_14657);
xor U16172 (N_16172,N_15349,N_14476);
nor U16173 (N_16173,N_14402,N_14960);
xor U16174 (N_16174,N_14733,N_14649);
or U16175 (N_16175,N_14877,N_15402);
or U16176 (N_16176,N_15069,N_14935);
or U16177 (N_16177,N_15414,N_14920);
nand U16178 (N_16178,N_15097,N_15332);
nand U16179 (N_16179,N_15561,N_14469);
nor U16180 (N_16180,N_14839,N_14693);
nand U16181 (N_16181,N_15309,N_15543);
or U16182 (N_16182,N_14621,N_14570);
xnor U16183 (N_16183,N_15225,N_15592);
nand U16184 (N_16184,N_15388,N_14614);
nand U16185 (N_16185,N_15281,N_15596);
xor U16186 (N_16186,N_15246,N_15184);
nand U16187 (N_16187,N_15595,N_15421);
or U16188 (N_16188,N_14579,N_15538);
and U16189 (N_16189,N_14623,N_14660);
and U16190 (N_16190,N_14844,N_15084);
xnor U16191 (N_16191,N_14867,N_15326);
and U16192 (N_16192,N_15513,N_15068);
nor U16193 (N_16193,N_14686,N_14781);
or U16194 (N_16194,N_14422,N_14531);
nor U16195 (N_16195,N_15145,N_15255);
nor U16196 (N_16196,N_14634,N_14406);
xor U16197 (N_16197,N_15416,N_15522);
and U16198 (N_16198,N_14405,N_14746);
and U16199 (N_16199,N_14497,N_14859);
and U16200 (N_16200,N_15599,N_14569);
or U16201 (N_16201,N_15583,N_14954);
xor U16202 (N_16202,N_15397,N_14547);
and U16203 (N_16203,N_14973,N_15295);
and U16204 (N_16204,N_15457,N_14888);
or U16205 (N_16205,N_14923,N_15417);
xor U16206 (N_16206,N_15029,N_15277);
and U16207 (N_16207,N_14891,N_15104);
nor U16208 (N_16208,N_15262,N_15564);
nand U16209 (N_16209,N_15082,N_14685);
and U16210 (N_16210,N_15098,N_15507);
and U16211 (N_16211,N_15537,N_14946);
and U16212 (N_16212,N_14845,N_15183);
xnor U16213 (N_16213,N_15287,N_14564);
nor U16214 (N_16214,N_14711,N_14519);
xor U16215 (N_16215,N_14756,N_14893);
xnor U16216 (N_16216,N_14852,N_15131);
or U16217 (N_16217,N_14839,N_14939);
or U16218 (N_16218,N_14870,N_14604);
and U16219 (N_16219,N_14422,N_15163);
nand U16220 (N_16220,N_15367,N_14888);
and U16221 (N_16221,N_14932,N_14620);
and U16222 (N_16222,N_14915,N_15142);
nand U16223 (N_16223,N_14945,N_15484);
and U16224 (N_16224,N_15281,N_14828);
and U16225 (N_16225,N_14935,N_15053);
nor U16226 (N_16226,N_14897,N_14982);
nand U16227 (N_16227,N_15220,N_15514);
nor U16228 (N_16228,N_15366,N_14694);
or U16229 (N_16229,N_14603,N_14610);
nand U16230 (N_16230,N_15132,N_15428);
and U16231 (N_16231,N_14989,N_15029);
and U16232 (N_16232,N_15258,N_14489);
and U16233 (N_16233,N_15181,N_15000);
nor U16234 (N_16234,N_14587,N_15567);
or U16235 (N_16235,N_15152,N_15133);
nor U16236 (N_16236,N_15246,N_14821);
and U16237 (N_16237,N_14762,N_15528);
or U16238 (N_16238,N_14886,N_15405);
and U16239 (N_16239,N_15063,N_15208);
or U16240 (N_16240,N_15028,N_14552);
and U16241 (N_16241,N_15256,N_14523);
xnor U16242 (N_16242,N_14707,N_15139);
and U16243 (N_16243,N_15401,N_14580);
and U16244 (N_16244,N_15345,N_14853);
or U16245 (N_16245,N_15569,N_14545);
xor U16246 (N_16246,N_15584,N_14758);
and U16247 (N_16247,N_15444,N_15437);
or U16248 (N_16248,N_14916,N_14873);
nand U16249 (N_16249,N_14540,N_15513);
nor U16250 (N_16250,N_15270,N_15444);
or U16251 (N_16251,N_15039,N_14872);
and U16252 (N_16252,N_14591,N_14598);
and U16253 (N_16253,N_15506,N_14424);
nor U16254 (N_16254,N_14515,N_15289);
nand U16255 (N_16255,N_14659,N_15306);
nand U16256 (N_16256,N_14770,N_14998);
nand U16257 (N_16257,N_14505,N_14662);
nor U16258 (N_16258,N_15478,N_14885);
and U16259 (N_16259,N_14983,N_14894);
and U16260 (N_16260,N_14929,N_14410);
or U16261 (N_16261,N_14744,N_15016);
xor U16262 (N_16262,N_14838,N_15111);
and U16263 (N_16263,N_15259,N_14958);
or U16264 (N_16264,N_15364,N_15337);
xor U16265 (N_16265,N_14755,N_14831);
nor U16266 (N_16266,N_14507,N_14795);
xor U16267 (N_16267,N_14782,N_15574);
xnor U16268 (N_16268,N_15378,N_15065);
nand U16269 (N_16269,N_15458,N_14844);
and U16270 (N_16270,N_14541,N_15105);
and U16271 (N_16271,N_14920,N_15157);
nor U16272 (N_16272,N_15506,N_14890);
and U16273 (N_16273,N_15426,N_15420);
or U16274 (N_16274,N_14637,N_14443);
xnor U16275 (N_16275,N_14970,N_14580);
xnor U16276 (N_16276,N_14477,N_14529);
nand U16277 (N_16277,N_15488,N_14544);
and U16278 (N_16278,N_15123,N_15465);
and U16279 (N_16279,N_14541,N_14782);
and U16280 (N_16280,N_14956,N_15128);
nor U16281 (N_16281,N_15366,N_15322);
nand U16282 (N_16282,N_14425,N_15545);
and U16283 (N_16283,N_14737,N_14987);
xor U16284 (N_16284,N_15477,N_15537);
nor U16285 (N_16285,N_14722,N_15530);
and U16286 (N_16286,N_15017,N_15468);
nor U16287 (N_16287,N_14979,N_15540);
xnor U16288 (N_16288,N_15140,N_15239);
nand U16289 (N_16289,N_15594,N_14971);
xor U16290 (N_16290,N_14634,N_15027);
nor U16291 (N_16291,N_15445,N_15335);
xnor U16292 (N_16292,N_14907,N_14550);
xor U16293 (N_16293,N_15449,N_14748);
nand U16294 (N_16294,N_14504,N_14449);
or U16295 (N_16295,N_15254,N_14802);
xor U16296 (N_16296,N_15422,N_14558);
and U16297 (N_16297,N_14759,N_14427);
nand U16298 (N_16298,N_15180,N_15252);
nand U16299 (N_16299,N_15256,N_15207);
xor U16300 (N_16300,N_15530,N_15204);
xor U16301 (N_16301,N_15391,N_15163);
nor U16302 (N_16302,N_14812,N_15551);
nand U16303 (N_16303,N_14502,N_14912);
or U16304 (N_16304,N_14828,N_14775);
or U16305 (N_16305,N_14767,N_15255);
nor U16306 (N_16306,N_14641,N_14560);
nor U16307 (N_16307,N_15504,N_15471);
nand U16308 (N_16308,N_15474,N_15559);
nand U16309 (N_16309,N_14406,N_15126);
nand U16310 (N_16310,N_15148,N_14688);
and U16311 (N_16311,N_15062,N_15120);
nand U16312 (N_16312,N_15073,N_15394);
and U16313 (N_16313,N_15315,N_15203);
and U16314 (N_16314,N_15125,N_14937);
xnor U16315 (N_16315,N_14560,N_14898);
nand U16316 (N_16316,N_14733,N_15285);
nand U16317 (N_16317,N_15363,N_14866);
xnor U16318 (N_16318,N_15432,N_14875);
nor U16319 (N_16319,N_15316,N_15455);
xor U16320 (N_16320,N_14723,N_15167);
nand U16321 (N_16321,N_14609,N_14580);
nand U16322 (N_16322,N_14502,N_14547);
xnor U16323 (N_16323,N_14520,N_14739);
or U16324 (N_16324,N_14772,N_14843);
nand U16325 (N_16325,N_14659,N_15352);
or U16326 (N_16326,N_14403,N_14422);
nor U16327 (N_16327,N_14524,N_14427);
nor U16328 (N_16328,N_15568,N_14452);
and U16329 (N_16329,N_14607,N_14631);
nor U16330 (N_16330,N_14570,N_15441);
and U16331 (N_16331,N_14672,N_14702);
or U16332 (N_16332,N_15118,N_14813);
nor U16333 (N_16333,N_15333,N_15541);
or U16334 (N_16334,N_14946,N_14557);
or U16335 (N_16335,N_15438,N_15171);
or U16336 (N_16336,N_14525,N_14905);
or U16337 (N_16337,N_14955,N_15197);
nand U16338 (N_16338,N_14579,N_14588);
nor U16339 (N_16339,N_15271,N_14687);
and U16340 (N_16340,N_15563,N_14931);
and U16341 (N_16341,N_15109,N_14508);
xnor U16342 (N_16342,N_15546,N_15262);
nand U16343 (N_16343,N_15281,N_15085);
nor U16344 (N_16344,N_14824,N_14591);
and U16345 (N_16345,N_14712,N_14721);
xnor U16346 (N_16346,N_14721,N_15418);
nand U16347 (N_16347,N_14746,N_15104);
or U16348 (N_16348,N_14969,N_15595);
nor U16349 (N_16349,N_15094,N_15428);
or U16350 (N_16350,N_15415,N_15133);
xnor U16351 (N_16351,N_15150,N_14468);
and U16352 (N_16352,N_15498,N_14506);
or U16353 (N_16353,N_15580,N_15198);
and U16354 (N_16354,N_15251,N_15511);
xor U16355 (N_16355,N_15049,N_14404);
and U16356 (N_16356,N_14802,N_14607);
or U16357 (N_16357,N_15113,N_14928);
nor U16358 (N_16358,N_14855,N_14653);
xor U16359 (N_16359,N_15175,N_15183);
nor U16360 (N_16360,N_14771,N_14665);
nand U16361 (N_16361,N_15167,N_15560);
nand U16362 (N_16362,N_15504,N_14896);
nand U16363 (N_16363,N_14681,N_15051);
xor U16364 (N_16364,N_15239,N_15386);
or U16365 (N_16365,N_15397,N_15293);
nand U16366 (N_16366,N_14762,N_14726);
nand U16367 (N_16367,N_15597,N_15022);
or U16368 (N_16368,N_15479,N_15181);
xor U16369 (N_16369,N_14681,N_15145);
nand U16370 (N_16370,N_14541,N_15595);
and U16371 (N_16371,N_15497,N_14628);
or U16372 (N_16372,N_14709,N_14809);
and U16373 (N_16373,N_14945,N_15582);
or U16374 (N_16374,N_15469,N_14908);
xor U16375 (N_16375,N_15374,N_14855);
xor U16376 (N_16376,N_15468,N_14917);
xor U16377 (N_16377,N_15183,N_15075);
or U16378 (N_16378,N_15479,N_14509);
and U16379 (N_16379,N_15255,N_14860);
nand U16380 (N_16380,N_15099,N_14405);
nor U16381 (N_16381,N_15252,N_14884);
or U16382 (N_16382,N_14865,N_14516);
or U16383 (N_16383,N_14706,N_15195);
and U16384 (N_16384,N_14546,N_15462);
or U16385 (N_16385,N_14498,N_14949);
and U16386 (N_16386,N_14942,N_14823);
nand U16387 (N_16387,N_15391,N_14863);
nor U16388 (N_16388,N_15177,N_14586);
and U16389 (N_16389,N_15491,N_14848);
nor U16390 (N_16390,N_14584,N_14696);
or U16391 (N_16391,N_15326,N_14608);
nor U16392 (N_16392,N_14981,N_15264);
nor U16393 (N_16393,N_15587,N_14935);
or U16394 (N_16394,N_15336,N_15298);
nor U16395 (N_16395,N_14778,N_15207);
xnor U16396 (N_16396,N_14403,N_14527);
nor U16397 (N_16397,N_14467,N_14536);
xor U16398 (N_16398,N_15191,N_14954);
nand U16399 (N_16399,N_14552,N_15376);
xnor U16400 (N_16400,N_15297,N_14955);
nand U16401 (N_16401,N_15113,N_15075);
nand U16402 (N_16402,N_15511,N_14842);
xnor U16403 (N_16403,N_14976,N_15485);
nand U16404 (N_16404,N_14837,N_14442);
nor U16405 (N_16405,N_14800,N_14943);
and U16406 (N_16406,N_14996,N_14728);
and U16407 (N_16407,N_15140,N_15517);
nand U16408 (N_16408,N_15234,N_15277);
or U16409 (N_16409,N_14661,N_14975);
and U16410 (N_16410,N_14911,N_14740);
and U16411 (N_16411,N_15494,N_15124);
nand U16412 (N_16412,N_15368,N_14437);
xor U16413 (N_16413,N_14839,N_14596);
or U16414 (N_16414,N_15498,N_15025);
xor U16415 (N_16415,N_15016,N_14960);
or U16416 (N_16416,N_15346,N_14679);
nand U16417 (N_16417,N_14709,N_15027);
or U16418 (N_16418,N_15591,N_15426);
nand U16419 (N_16419,N_14506,N_15229);
nand U16420 (N_16420,N_15096,N_15046);
nor U16421 (N_16421,N_14619,N_15412);
and U16422 (N_16422,N_14938,N_15149);
xor U16423 (N_16423,N_14719,N_14968);
nor U16424 (N_16424,N_14500,N_15197);
xnor U16425 (N_16425,N_15419,N_14826);
nand U16426 (N_16426,N_15124,N_15137);
nand U16427 (N_16427,N_15466,N_14563);
and U16428 (N_16428,N_15141,N_15336);
nor U16429 (N_16429,N_15588,N_15220);
or U16430 (N_16430,N_14640,N_15418);
or U16431 (N_16431,N_14641,N_15495);
or U16432 (N_16432,N_14423,N_15028);
or U16433 (N_16433,N_14414,N_14870);
nor U16434 (N_16434,N_14458,N_14911);
and U16435 (N_16435,N_14718,N_15110);
xnor U16436 (N_16436,N_14521,N_14957);
xor U16437 (N_16437,N_14529,N_15325);
and U16438 (N_16438,N_14780,N_14861);
or U16439 (N_16439,N_14601,N_14655);
xor U16440 (N_16440,N_14938,N_14797);
and U16441 (N_16441,N_14962,N_15493);
and U16442 (N_16442,N_14725,N_15521);
or U16443 (N_16443,N_15060,N_15433);
and U16444 (N_16444,N_15265,N_15169);
xor U16445 (N_16445,N_15301,N_14516);
nor U16446 (N_16446,N_15120,N_14941);
xnor U16447 (N_16447,N_15408,N_14404);
and U16448 (N_16448,N_15151,N_15473);
and U16449 (N_16449,N_14999,N_14933);
and U16450 (N_16450,N_15512,N_15588);
nand U16451 (N_16451,N_15008,N_15271);
xor U16452 (N_16452,N_14555,N_14800);
nand U16453 (N_16453,N_14813,N_15472);
and U16454 (N_16454,N_15291,N_14750);
nand U16455 (N_16455,N_15179,N_15104);
or U16456 (N_16456,N_14605,N_15359);
xnor U16457 (N_16457,N_14446,N_15054);
nor U16458 (N_16458,N_14540,N_14488);
xor U16459 (N_16459,N_15271,N_14845);
xor U16460 (N_16460,N_14771,N_15510);
and U16461 (N_16461,N_14476,N_15414);
xnor U16462 (N_16462,N_15582,N_15341);
and U16463 (N_16463,N_15560,N_14833);
xor U16464 (N_16464,N_14617,N_15233);
nand U16465 (N_16465,N_14919,N_15343);
nor U16466 (N_16466,N_14619,N_15358);
and U16467 (N_16467,N_14491,N_14673);
nand U16468 (N_16468,N_15151,N_14416);
or U16469 (N_16469,N_15143,N_15469);
xor U16470 (N_16470,N_15556,N_14688);
and U16471 (N_16471,N_14900,N_15286);
or U16472 (N_16472,N_14411,N_14673);
nor U16473 (N_16473,N_15509,N_14640);
nor U16474 (N_16474,N_14691,N_15147);
nor U16475 (N_16475,N_14441,N_14935);
nor U16476 (N_16476,N_14815,N_14928);
and U16477 (N_16477,N_15511,N_14793);
xnor U16478 (N_16478,N_14772,N_14869);
nand U16479 (N_16479,N_15098,N_15170);
or U16480 (N_16480,N_15094,N_15198);
xnor U16481 (N_16481,N_14668,N_15187);
nand U16482 (N_16482,N_15598,N_15115);
xor U16483 (N_16483,N_14854,N_15334);
or U16484 (N_16484,N_15337,N_14918);
nor U16485 (N_16485,N_14935,N_14937);
nor U16486 (N_16486,N_15141,N_15245);
and U16487 (N_16487,N_15525,N_15596);
and U16488 (N_16488,N_14658,N_14590);
xor U16489 (N_16489,N_15503,N_15010);
or U16490 (N_16490,N_14635,N_15484);
nand U16491 (N_16491,N_15566,N_14913);
or U16492 (N_16492,N_14797,N_14450);
or U16493 (N_16493,N_15477,N_14881);
or U16494 (N_16494,N_14779,N_15428);
xor U16495 (N_16495,N_15476,N_15037);
nand U16496 (N_16496,N_15346,N_15049);
or U16497 (N_16497,N_14789,N_15406);
and U16498 (N_16498,N_15124,N_14687);
xor U16499 (N_16499,N_14968,N_15072);
and U16500 (N_16500,N_14785,N_14710);
nand U16501 (N_16501,N_15399,N_15439);
and U16502 (N_16502,N_14425,N_15398);
xnor U16503 (N_16503,N_15425,N_14526);
or U16504 (N_16504,N_15415,N_14961);
or U16505 (N_16505,N_14865,N_15306);
and U16506 (N_16506,N_15230,N_15094);
and U16507 (N_16507,N_14781,N_14990);
nor U16508 (N_16508,N_15270,N_15541);
xnor U16509 (N_16509,N_15179,N_14924);
and U16510 (N_16510,N_15535,N_14658);
and U16511 (N_16511,N_15252,N_15008);
xnor U16512 (N_16512,N_14935,N_14886);
and U16513 (N_16513,N_14432,N_14631);
and U16514 (N_16514,N_15247,N_14719);
or U16515 (N_16515,N_15129,N_15301);
or U16516 (N_16516,N_14772,N_14680);
or U16517 (N_16517,N_14748,N_15047);
nand U16518 (N_16518,N_15371,N_14753);
nor U16519 (N_16519,N_15248,N_14730);
or U16520 (N_16520,N_14944,N_14677);
nor U16521 (N_16521,N_15142,N_14801);
nor U16522 (N_16522,N_14420,N_14456);
and U16523 (N_16523,N_14665,N_14627);
nor U16524 (N_16524,N_15380,N_15278);
and U16525 (N_16525,N_14833,N_15518);
nor U16526 (N_16526,N_15049,N_15171);
or U16527 (N_16527,N_15326,N_15323);
nor U16528 (N_16528,N_14554,N_14711);
nor U16529 (N_16529,N_14591,N_15016);
nor U16530 (N_16530,N_14609,N_15232);
and U16531 (N_16531,N_14476,N_14502);
or U16532 (N_16532,N_14424,N_15503);
nand U16533 (N_16533,N_14778,N_14753);
and U16534 (N_16534,N_14734,N_15564);
xnor U16535 (N_16535,N_14472,N_15309);
nor U16536 (N_16536,N_14415,N_15065);
and U16537 (N_16537,N_15397,N_15210);
nand U16538 (N_16538,N_14401,N_15570);
or U16539 (N_16539,N_14873,N_14910);
and U16540 (N_16540,N_14546,N_14549);
nor U16541 (N_16541,N_15174,N_14596);
nor U16542 (N_16542,N_15004,N_14771);
xor U16543 (N_16543,N_15265,N_14443);
nor U16544 (N_16544,N_14447,N_15207);
or U16545 (N_16545,N_15547,N_14921);
or U16546 (N_16546,N_15037,N_14970);
xor U16547 (N_16547,N_15515,N_14663);
or U16548 (N_16548,N_14603,N_14683);
and U16549 (N_16549,N_14529,N_15238);
and U16550 (N_16550,N_14922,N_14884);
nor U16551 (N_16551,N_14428,N_15072);
xor U16552 (N_16552,N_14759,N_14869);
xor U16553 (N_16553,N_14940,N_15525);
nand U16554 (N_16554,N_15580,N_14672);
xor U16555 (N_16555,N_15356,N_15051);
and U16556 (N_16556,N_15061,N_15078);
and U16557 (N_16557,N_14780,N_15318);
nor U16558 (N_16558,N_14556,N_15213);
and U16559 (N_16559,N_15123,N_15328);
and U16560 (N_16560,N_14448,N_14563);
nor U16561 (N_16561,N_14765,N_14558);
nand U16562 (N_16562,N_14739,N_14430);
xnor U16563 (N_16563,N_14428,N_15224);
and U16564 (N_16564,N_15597,N_14973);
or U16565 (N_16565,N_15131,N_15490);
xnor U16566 (N_16566,N_15317,N_15460);
nor U16567 (N_16567,N_15301,N_15136);
or U16568 (N_16568,N_14755,N_14731);
nor U16569 (N_16569,N_15016,N_15247);
xor U16570 (N_16570,N_14792,N_15158);
xnor U16571 (N_16571,N_15114,N_14834);
nand U16572 (N_16572,N_15160,N_14687);
xnor U16573 (N_16573,N_14977,N_14633);
and U16574 (N_16574,N_14967,N_14976);
nand U16575 (N_16575,N_14794,N_14427);
nor U16576 (N_16576,N_15079,N_15341);
or U16577 (N_16577,N_15574,N_14881);
nand U16578 (N_16578,N_15435,N_15552);
or U16579 (N_16579,N_14707,N_14776);
or U16580 (N_16580,N_15323,N_15115);
or U16581 (N_16581,N_14523,N_14537);
and U16582 (N_16582,N_14419,N_14835);
and U16583 (N_16583,N_14587,N_14457);
and U16584 (N_16584,N_14855,N_15598);
and U16585 (N_16585,N_14495,N_14608);
nor U16586 (N_16586,N_14400,N_14998);
or U16587 (N_16587,N_14620,N_15094);
or U16588 (N_16588,N_14600,N_14977);
xor U16589 (N_16589,N_14724,N_15013);
or U16590 (N_16590,N_15539,N_15580);
nand U16591 (N_16591,N_14863,N_15205);
nor U16592 (N_16592,N_14683,N_14443);
xnor U16593 (N_16593,N_14740,N_15341);
or U16594 (N_16594,N_14850,N_15201);
or U16595 (N_16595,N_14591,N_15224);
or U16596 (N_16596,N_14922,N_14451);
nand U16597 (N_16597,N_15325,N_15255);
nand U16598 (N_16598,N_14444,N_15113);
nor U16599 (N_16599,N_14871,N_14842);
xnor U16600 (N_16600,N_15048,N_14743);
or U16601 (N_16601,N_15042,N_15315);
nor U16602 (N_16602,N_15531,N_15597);
nor U16603 (N_16603,N_14846,N_14498);
nand U16604 (N_16604,N_15086,N_15037);
xor U16605 (N_16605,N_15199,N_15142);
nand U16606 (N_16606,N_15397,N_14579);
and U16607 (N_16607,N_15212,N_14703);
or U16608 (N_16608,N_14452,N_14693);
nand U16609 (N_16609,N_14469,N_15586);
or U16610 (N_16610,N_14418,N_15417);
or U16611 (N_16611,N_15196,N_15252);
or U16612 (N_16612,N_14734,N_15417);
or U16613 (N_16613,N_14411,N_14543);
and U16614 (N_16614,N_14662,N_14897);
xnor U16615 (N_16615,N_14549,N_14941);
and U16616 (N_16616,N_15492,N_14553);
and U16617 (N_16617,N_14900,N_15225);
and U16618 (N_16618,N_15468,N_15201);
or U16619 (N_16619,N_14986,N_14790);
or U16620 (N_16620,N_14406,N_15066);
xor U16621 (N_16621,N_15002,N_15270);
and U16622 (N_16622,N_14998,N_14918);
or U16623 (N_16623,N_14648,N_14854);
xor U16624 (N_16624,N_15323,N_14609);
xnor U16625 (N_16625,N_15078,N_14631);
and U16626 (N_16626,N_15463,N_14658);
nor U16627 (N_16627,N_15204,N_15170);
nor U16628 (N_16628,N_15595,N_14884);
nand U16629 (N_16629,N_14525,N_14783);
and U16630 (N_16630,N_15561,N_15434);
nor U16631 (N_16631,N_15279,N_14823);
nand U16632 (N_16632,N_14460,N_15018);
nand U16633 (N_16633,N_14709,N_14550);
nand U16634 (N_16634,N_15419,N_14770);
and U16635 (N_16635,N_15586,N_15225);
nand U16636 (N_16636,N_15548,N_15382);
and U16637 (N_16637,N_15450,N_15084);
nor U16638 (N_16638,N_14530,N_14664);
xor U16639 (N_16639,N_15272,N_14855);
or U16640 (N_16640,N_14963,N_14540);
and U16641 (N_16641,N_15132,N_15124);
nand U16642 (N_16642,N_14720,N_14950);
or U16643 (N_16643,N_15579,N_14646);
xor U16644 (N_16644,N_14947,N_15229);
nand U16645 (N_16645,N_14774,N_14968);
and U16646 (N_16646,N_14931,N_15582);
nand U16647 (N_16647,N_15291,N_15505);
nor U16648 (N_16648,N_14636,N_14940);
or U16649 (N_16649,N_14627,N_14961);
or U16650 (N_16650,N_14604,N_15191);
xor U16651 (N_16651,N_15187,N_15275);
and U16652 (N_16652,N_15495,N_15585);
or U16653 (N_16653,N_15374,N_14868);
nor U16654 (N_16654,N_15380,N_15452);
or U16655 (N_16655,N_14956,N_15213);
or U16656 (N_16656,N_14970,N_15416);
nand U16657 (N_16657,N_15035,N_14723);
nor U16658 (N_16658,N_15535,N_15449);
nor U16659 (N_16659,N_14440,N_15598);
nor U16660 (N_16660,N_14814,N_14403);
or U16661 (N_16661,N_14651,N_14825);
xor U16662 (N_16662,N_14695,N_14572);
or U16663 (N_16663,N_14989,N_15299);
nand U16664 (N_16664,N_15589,N_14808);
nand U16665 (N_16665,N_14527,N_14578);
or U16666 (N_16666,N_15552,N_15467);
nand U16667 (N_16667,N_15514,N_14820);
xnor U16668 (N_16668,N_14633,N_14557);
xor U16669 (N_16669,N_14916,N_15049);
nand U16670 (N_16670,N_15372,N_14651);
nand U16671 (N_16671,N_14602,N_14575);
and U16672 (N_16672,N_14695,N_14504);
or U16673 (N_16673,N_14585,N_15509);
nor U16674 (N_16674,N_15545,N_14952);
or U16675 (N_16675,N_14535,N_15457);
and U16676 (N_16676,N_15107,N_14708);
or U16677 (N_16677,N_14875,N_14818);
and U16678 (N_16678,N_14708,N_14660);
nor U16679 (N_16679,N_15400,N_14783);
xor U16680 (N_16680,N_15203,N_15074);
or U16681 (N_16681,N_14998,N_14823);
xnor U16682 (N_16682,N_15119,N_15044);
or U16683 (N_16683,N_14822,N_15178);
nand U16684 (N_16684,N_14700,N_14691);
or U16685 (N_16685,N_14842,N_15260);
nand U16686 (N_16686,N_14529,N_15510);
or U16687 (N_16687,N_15251,N_14626);
xor U16688 (N_16688,N_15350,N_15174);
or U16689 (N_16689,N_14988,N_14842);
xnor U16690 (N_16690,N_15078,N_14588);
and U16691 (N_16691,N_14809,N_15463);
or U16692 (N_16692,N_14487,N_15440);
nor U16693 (N_16693,N_14583,N_14704);
nor U16694 (N_16694,N_15153,N_15437);
and U16695 (N_16695,N_14879,N_14562);
nand U16696 (N_16696,N_15412,N_14736);
or U16697 (N_16697,N_15305,N_14992);
nor U16698 (N_16698,N_14839,N_15529);
xnor U16699 (N_16699,N_15313,N_14959);
and U16700 (N_16700,N_14685,N_15216);
and U16701 (N_16701,N_15231,N_15435);
nor U16702 (N_16702,N_15107,N_15162);
nand U16703 (N_16703,N_15201,N_15394);
nand U16704 (N_16704,N_14565,N_15280);
xor U16705 (N_16705,N_15598,N_15285);
nand U16706 (N_16706,N_14595,N_15580);
nor U16707 (N_16707,N_14973,N_15216);
nor U16708 (N_16708,N_15075,N_15425);
nor U16709 (N_16709,N_14629,N_14656);
and U16710 (N_16710,N_15463,N_14518);
or U16711 (N_16711,N_14785,N_15095);
nor U16712 (N_16712,N_15072,N_14554);
xnor U16713 (N_16713,N_14707,N_14451);
or U16714 (N_16714,N_15162,N_15159);
nand U16715 (N_16715,N_14610,N_14695);
or U16716 (N_16716,N_14724,N_15547);
nand U16717 (N_16717,N_14690,N_15357);
nor U16718 (N_16718,N_14543,N_15211);
and U16719 (N_16719,N_15090,N_14657);
xor U16720 (N_16720,N_15560,N_15327);
and U16721 (N_16721,N_15199,N_15323);
nor U16722 (N_16722,N_15257,N_15060);
xor U16723 (N_16723,N_14656,N_15011);
xor U16724 (N_16724,N_14920,N_14719);
nand U16725 (N_16725,N_14629,N_14549);
or U16726 (N_16726,N_15139,N_14491);
nand U16727 (N_16727,N_15241,N_15124);
nor U16728 (N_16728,N_14719,N_15353);
nand U16729 (N_16729,N_14665,N_15488);
nor U16730 (N_16730,N_14911,N_15479);
nand U16731 (N_16731,N_15019,N_14644);
xor U16732 (N_16732,N_14435,N_15128);
or U16733 (N_16733,N_14481,N_14482);
nor U16734 (N_16734,N_14842,N_15470);
nor U16735 (N_16735,N_14888,N_14536);
nor U16736 (N_16736,N_14739,N_15491);
or U16737 (N_16737,N_14945,N_14851);
nor U16738 (N_16738,N_14929,N_15290);
xnor U16739 (N_16739,N_14939,N_14691);
xnor U16740 (N_16740,N_15107,N_15324);
xor U16741 (N_16741,N_15395,N_15472);
nor U16742 (N_16742,N_15500,N_14500);
and U16743 (N_16743,N_15216,N_15332);
xnor U16744 (N_16744,N_14524,N_15423);
xnor U16745 (N_16745,N_14870,N_14952);
or U16746 (N_16746,N_14425,N_14591);
nand U16747 (N_16747,N_15238,N_14599);
xor U16748 (N_16748,N_14907,N_14844);
nand U16749 (N_16749,N_14691,N_14401);
or U16750 (N_16750,N_15358,N_15469);
or U16751 (N_16751,N_14523,N_14778);
or U16752 (N_16752,N_14599,N_15223);
nand U16753 (N_16753,N_14873,N_15155);
and U16754 (N_16754,N_15391,N_15092);
and U16755 (N_16755,N_14605,N_15598);
or U16756 (N_16756,N_14482,N_15585);
and U16757 (N_16757,N_14422,N_15519);
or U16758 (N_16758,N_14581,N_15325);
xnor U16759 (N_16759,N_15562,N_15119);
nand U16760 (N_16760,N_15365,N_14528);
nand U16761 (N_16761,N_14814,N_15291);
nand U16762 (N_16762,N_14997,N_14856);
and U16763 (N_16763,N_14651,N_14962);
or U16764 (N_16764,N_14891,N_15084);
xor U16765 (N_16765,N_15521,N_14616);
nand U16766 (N_16766,N_14502,N_14513);
and U16767 (N_16767,N_15074,N_14713);
and U16768 (N_16768,N_15369,N_14811);
and U16769 (N_16769,N_14854,N_14469);
xnor U16770 (N_16770,N_14444,N_15215);
nand U16771 (N_16771,N_14454,N_14538);
or U16772 (N_16772,N_14824,N_15403);
xnor U16773 (N_16773,N_15009,N_15058);
or U16774 (N_16774,N_14803,N_14899);
and U16775 (N_16775,N_15589,N_14930);
and U16776 (N_16776,N_14507,N_15226);
nor U16777 (N_16777,N_15336,N_15197);
or U16778 (N_16778,N_15097,N_15591);
xnor U16779 (N_16779,N_14824,N_14757);
xor U16780 (N_16780,N_15010,N_14614);
nor U16781 (N_16781,N_15246,N_14700);
and U16782 (N_16782,N_15129,N_14749);
nand U16783 (N_16783,N_15248,N_15020);
nand U16784 (N_16784,N_15277,N_15152);
xnor U16785 (N_16785,N_15402,N_15152);
or U16786 (N_16786,N_14528,N_15370);
nor U16787 (N_16787,N_14779,N_14430);
nor U16788 (N_16788,N_14578,N_14654);
and U16789 (N_16789,N_14446,N_14492);
and U16790 (N_16790,N_14797,N_14859);
and U16791 (N_16791,N_15269,N_15570);
nor U16792 (N_16792,N_15053,N_14897);
nor U16793 (N_16793,N_14567,N_14492);
nor U16794 (N_16794,N_14519,N_14556);
and U16795 (N_16795,N_14579,N_14661);
nand U16796 (N_16796,N_15166,N_14642);
xnor U16797 (N_16797,N_15151,N_15397);
nor U16798 (N_16798,N_15584,N_15315);
or U16799 (N_16799,N_14641,N_15355);
or U16800 (N_16800,N_16293,N_16202);
nor U16801 (N_16801,N_16419,N_15707);
nor U16802 (N_16802,N_16731,N_15956);
or U16803 (N_16803,N_16283,N_16073);
or U16804 (N_16804,N_15808,N_16199);
nand U16805 (N_16805,N_16372,N_15861);
xor U16806 (N_16806,N_16373,N_16516);
or U16807 (N_16807,N_16680,N_15799);
xnor U16808 (N_16808,N_16125,N_15982);
or U16809 (N_16809,N_15983,N_16299);
or U16810 (N_16810,N_15782,N_16296);
and U16811 (N_16811,N_15710,N_16257);
xnor U16812 (N_16812,N_15683,N_15600);
nor U16813 (N_16813,N_16721,N_16263);
or U16814 (N_16814,N_16077,N_16677);
nor U16815 (N_16815,N_15976,N_16784);
or U16816 (N_16816,N_15796,N_15879);
and U16817 (N_16817,N_16595,N_16094);
or U16818 (N_16818,N_16301,N_16122);
nand U16819 (N_16819,N_16069,N_15787);
xnor U16820 (N_16820,N_16130,N_16398);
nor U16821 (N_16821,N_15711,N_16729);
xnor U16822 (N_16822,N_15862,N_16749);
nand U16823 (N_16823,N_15809,N_16639);
nand U16824 (N_16824,N_16783,N_16205);
or U16825 (N_16825,N_15853,N_15999);
nor U16826 (N_16826,N_15623,N_16110);
xor U16827 (N_16827,N_16324,N_16294);
and U16828 (N_16828,N_16087,N_16287);
nand U16829 (N_16829,N_15951,N_16507);
nor U16830 (N_16830,N_16367,N_16111);
or U16831 (N_16831,N_16173,N_16082);
nor U16832 (N_16832,N_16102,N_16103);
or U16833 (N_16833,N_16148,N_16559);
xnor U16834 (N_16834,N_16341,N_15829);
or U16835 (N_16835,N_16260,N_16186);
or U16836 (N_16836,N_16676,N_15653);
xnor U16837 (N_16837,N_16161,N_15668);
or U16838 (N_16838,N_16190,N_15677);
nor U16839 (N_16839,N_16621,N_16646);
xor U16840 (N_16840,N_16259,N_16175);
xor U16841 (N_16841,N_15775,N_16389);
xnor U16842 (N_16842,N_16782,N_16185);
or U16843 (N_16843,N_16264,N_16158);
nor U16844 (N_16844,N_16041,N_15715);
nand U16845 (N_16845,N_16157,N_15661);
nor U16846 (N_16846,N_16654,N_15871);
xor U16847 (N_16847,N_15902,N_15795);
and U16848 (N_16848,N_16514,N_16617);
nor U16849 (N_16849,N_15953,N_16121);
nand U16850 (N_16850,N_16156,N_16775);
xor U16851 (N_16851,N_16402,N_16705);
xnor U16852 (N_16852,N_15603,N_16285);
nor U16853 (N_16853,N_16028,N_16583);
nor U16854 (N_16854,N_16049,N_16127);
and U16855 (N_16855,N_16180,N_15842);
xor U16856 (N_16856,N_16115,N_16144);
nor U16857 (N_16857,N_16723,N_16416);
and U16858 (N_16858,N_15629,N_16358);
nand U16859 (N_16859,N_16756,N_15967);
and U16860 (N_16860,N_15865,N_15877);
or U16861 (N_16861,N_16136,N_15770);
xnor U16862 (N_16862,N_15634,N_16504);
nand U16863 (N_16863,N_15726,N_16669);
xnor U16864 (N_16864,N_16235,N_15759);
nor U16865 (N_16865,N_16265,N_16084);
and U16866 (N_16866,N_16500,N_15984);
xnor U16867 (N_16867,N_16492,N_16386);
nand U16868 (N_16868,N_16089,N_15636);
and U16869 (N_16869,N_16760,N_16607);
or U16870 (N_16870,N_16138,N_16380);
and U16871 (N_16871,N_15693,N_16425);
or U16872 (N_16872,N_15851,N_16441);
and U16873 (N_16873,N_16155,N_16550);
xnor U16874 (N_16874,N_16465,N_16240);
xnor U16875 (N_16875,N_15971,N_16593);
nand U16876 (N_16876,N_16390,N_16776);
xor U16877 (N_16877,N_16479,N_16740);
and U16878 (N_16878,N_16295,N_15901);
nor U16879 (N_16879,N_16651,N_16472);
nand U16880 (N_16880,N_16707,N_15631);
nor U16881 (N_16881,N_16636,N_16460);
and U16882 (N_16882,N_15699,N_16739);
or U16883 (N_16883,N_16236,N_16542);
xnor U16884 (N_16884,N_16489,N_15972);
nor U16885 (N_16885,N_15671,N_16284);
and U16886 (N_16886,N_16513,N_16759);
or U16887 (N_16887,N_16698,N_15942);
or U16888 (N_16888,N_16043,N_16768);
or U16889 (N_16889,N_16750,N_16498);
or U16890 (N_16890,N_15687,N_16228);
nand U16891 (N_16891,N_15977,N_16382);
and U16892 (N_16892,N_16015,N_15614);
and U16893 (N_16893,N_16563,N_16001);
xor U16894 (N_16894,N_16469,N_16422);
xor U16895 (N_16895,N_15692,N_16256);
nand U16896 (N_16896,N_16211,N_16374);
and U16897 (N_16897,N_15788,N_16747);
xor U16898 (N_16898,N_16695,N_16413);
xnor U16899 (N_16899,N_16455,N_16360);
nand U16900 (N_16900,N_15811,N_16400);
xor U16901 (N_16901,N_16742,N_16449);
and U16902 (N_16902,N_16376,N_15756);
xnor U16903 (N_16903,N_16451,N_16107);
xnor U16904 (N_16904,N_16735,N_15914);
xnor U16905 (N_16905,N_16765,N_15663);
nor U16906 (N_16906,N_16524,N_15718);
xor U16907 (N_16907,N_15749,N_16053);
or U16908 (N_16908,N_16799,N_15651);
and U16909 (N_16909,N_15695,N_16629);
or U16910 (N_16910,N_16409,N_16335);
or U16911 (N_16911,N_16456,N_16364);
nor U16912 (N_16912,N_16706,N_15689);
nand U16913 (N_16913,N_15819,N_15728);
nor U16914 (N_16914,N_16063,N_15860);
nand U16915 (N_16915,N_16201,N_16589);
nor U16916 (N_16916,N_16569,N_15913);
nand U16917 (N_16917,N_15934,N_16781);
xnor U16918 (N_16918,N_16744,N_15680);
or U16919 (N_16919,N_16601,N_15832);
nor U16920 (N_16920,N_16525,N_16603);
xnor U16921 (N_16921,N_16671,N_15607);
nand U16922 (N_16922,N_16548,N_16659);
nor U16923 (N_16923,N_15605,N_15817);
xor U16924 (N_16924,N_15713,N_15735);
nor U16925 (N_16925,N_16541,N_16309);
xor U16926 (N_16926,N_16033,N_15827);
xnor U16927 (N_16927,N_16143,N_16270);
nor U16928 (N_16928,N_16345,N_16027);
xor U16929 (N_16929,N_15880,N_15868);
xor U16930 (N_16930,N_15968,N_16463);
nor U16931 (N_16931,N_16062,N_16553);
xor U16932 (N_16932,N_16332,N_16697);
or U16933 (N_16933,N_16474,N_15667);
xnor U16934 (N_16934,N_16690,N_16442);
nor U16935 (N_16935,N_16058,N_16401);
and U16936 (N_16936,N_16040,N_15950);
nor U16937 (N_16937,N_15685,N_15890);
nor U16938 (N_16938,N_16701,N_16773);
nor U16939 (N_16939,N_15815,N_16610);
and U16940 (N_16940,N_15801,N_15924);
nor U16941 (N_16941,N_15980,N_16439);
or U16942 (N_16942,N_16579,N_16317);
nor U16943 (N_16943,N_16162,N_16286);
nand U16944 (N_16944,N_15821,N_15993);
or U16945 (N_16945,N_15618,N_16414);
and U16946 (N_16946,N_16710,N_16220);
xnor U16947 (N_16947,N_16101,N_16300);
nor U16948 (N_16948,N_16667,N_16291);
xor U16949 (N_16949,N_16734,N_16793);
nand U16950 (N_16950,N_15622,N_16711);
and U16951 (N_16951,N_15732,N_15873);
and U16952 (N_16952,N_15978,N_16511);
or U16953 (N_16953,N_16509,N_16704);
nor U16954 (N_16954,N_15790,N_16237);
xnor U16955 (N_16955,N_16097,N_16246);
or U16956 (N_16956,N_16369,N_16245);
or U16957 (N_16957,N_16243,N_15784);
nand U16958 (N_16958,N_15818,N_15656);
nor U16959 (N_16959,N_16433,N_15994);
and U16960 (N_16960,N_16571,N_15985);
nor U16961 (N_16961,N_15665,N_16017);
xor U16962 (N_16962,N_16078,N_16010);
and U16963 (N_16963,N_16716,N_15601);
nor U16964 (N_16964,N_16528,N_16356);
and U16965 (N_16965,N_15814,N_16444);
xnor U16966 (N_16966,N_15813,N_16774);
nand U16967 (N_16967,N_15965,N_15996);
nand U16968 (N_16968,N_16537,N_15910);
and U16969 (N_16969,N_16539,N_16391);
nand U16970 (N_16970,N_16653,N_16616);
nor U16971 (N_16971,N_16663,N_16351);
nand U16972 (N_16972,N_15893,N_16751);
or U16973 (N_16973,N_16503,N_16549);
or U16974 (N_16974,N_16334,N_15630);
xnor U16975 (N_16975,N_16435,N_16008);
nor U16976 (N_16976,N_16722,N_15625);
and U16977 (N_16977,N_15849,N_16383);
nor U16978 (N_16978,N_15803,N_16418);
nor U16979 (N_16979,N_15908,N_15744);
or U16980 (N_16980,N_16182,N_16066);
nand U16981 (N_16981,N_16683,N_15964);
or U16982 (N_16982,N_16798,N_15643);
nand U16983 (N_16983,N_15941,N_15812);
nand U16984 (N_16984,N_15963,N_16321);
nand U16985 (N_16985,N_16557,N_16044);
nand U16986 (N_16986,N_16530,N_16496);
nand U16987 (N_16987,N_16666,N_16737);
nor U16988 (N_16988,N_16709,N_16311);
or U16989 (N_16989,N_16458,N_16596);
or U16990 (N_16990,N_15785,N_15768);
nor U16991 (N_16991,N_16404,N_16067);
nand U16992 (N_16992,N_16393,N_15940);
nor U16993 (N_16993,N_16230,N_16794);
or U16994 (N_16994,N_16167,N_15872);
nor U16995 (N_16995,N_16766,N_15611);
or U16996 (N_16996,N_16743,N_15616);
and U16997 (N_16997,N_16209,N_16253);
or U16998 (N_16998,N_15904,N_15739);
nand U16999 (N_16999,N_16114,N_15640);
and U17000 (N_17000,N_16649,N_16502);
nand U17001 (N_17001,N_15991,N_15959);
nand U17002 (N_17002,N_16598,N_16092);
or U17003 (N_17003,N_15754,N_16397);
nand U17004 (N_17004,N_16289,N_16061);
and U17005 (N_17005,N_16518,N_16031);
nor U17006 (N_17006,N_15684,N_15751);
and U17007 (N_17007,N_16515,N_16764);
nand U17008 (N_17008,N_15706,N_16674);
xor U17009 (N_17009,N_16178,N_16552);
nand U17010 (N_17010,N_16785,N_16415);
nand U17011 (N_17011,N_16468,N_16079);
nand U17012 (N_17012,N_15780,N_16672);
nand U17013 (N_17013,N_16531,N_16277);
and U17014 (N_17014,N_16778,N_16080);
nand U17015 (N_17015,N_15610,N_15792);
and U17016 (N_17016,N_16223,N_16032);
nand U17017 (N_17017,N_15762,N_16357);
xor U17018 (N_17018,N_15774,N_16745);
nand U17019 (N_17019,N_15837,N_16151);
and U17020 (N_17020,N_16184,N_16189);
xor U17021 (N_17021,N_15866,N_15800);
xnor U17022 (N_17022,N_16484,N_16347);
xnor U17023 (N_17023,N_16577,N_16312);
xor U17024 (N_17024,N_16034,N_16030);
or U17025 (N_17025,N_16007,N_16466);
and U17026 (N_17026,N_16700,N_16478);
and U17027 (N_17027,N_16226,N_15719);
xor U17028 (N_17028,N_16141,N_15828);
nand U17029 (N_17029,N_15724,N_16005);
and U17030 (N_17030,N_16540,N_15670);
nand U17031 (N_17031,N_15928,N_15926);
and U17032 (N_17032,N_15835,N_16188);
nand U17033 (N_17033,N_16399,N_15781);
nand U17034 (N_17034,N_15620,N_16592);
and U17035 (N_17035,N_16385,N_15907);
nor U17036 (N_17036,N_16055,N_15944);
and U17037 (N_17037,N_15712,N_16483);
nand U17038 (N_17038,N_16568,N_15645);
xor U17039 (N_17039,N_16655,N_15777);
nand U17040 (N_17040,N_15672,N_15826);
nand U17041 (N_17041,N_16308,N_16318);
nand U17042 (N_17042,N_15697,N_16306);
and U17043 (N_17043,N_16430,N_16462);
nor U17044 (N_17044,N_16229,N_16591);
or U17045 (N_17045,N_15648,N_15845);
or U17046 (N_17046,N_15676,N_16543);
or U17047 (N_17047,N_15738,N_16322);
nand U17048 (N_17048,N_16355,N_16112);
xnor U17049 (N_17049,N_16426,N_16072);
xor U17050 (N_17050,N_16625,N_16247);
xnor U17051 (N_17051,N_16251,N_15617);
or U17052 (N_17052,N_16753,N_15825);
nor U17053 (N_17053,N_15824,N_15854);
nor U17054 (N_17054,N_15764,N_16123);
nand U17055 (N_17055,N_15624,N_16586);
or U17056 (N_17056,N_15874,N_16482);
nand U17057 (N_17057,N_16224,N_16023);
or U17058 (N_17058,N_15938,N_15917);
nor U17059 (N_17059,N_16686,N_16396);
or U17060 (N_17060,N_16748,N_16198);
xor U17061 (N_17061,N_16656,N_16488);
and U17062 (N_17062,N_16522,N_16298);
nand U17063 (N_17063,N_15752,N_16420);
or U17064 (N_17064,N_16417,N_16403);
and U17065 (N_17065,N_16575,N_16349);
or U17066 (N_17066,N_16445,N_16570);
or U17067 (N_17067,N_16556,N_15935);
nand U17068 (N_17068,N_16217,N_16523);
and U17069 (N_17069,N_16611,N_16780);
nor U17070 (N_17070,N_16025,N_15615);
nor U17071 (N_17071,N_16641,N_16786);
nor U17072 (N_17072,N_16368,N_16673);
nor U17073 (N_17073,N_16447,N_16431);
xnor U17074 (N_17074,N_16736,N_15887);
xor U17075 (N_17075,N_16637,N_16423);
or U17076 (N_17076,N_16521,N_15923);
nand U17077 (N_17077,N_16137,N_15740);
xor U17078 (N_17078,N_16567,N_15834);
xnor U17079 (N_17079,N_16056,N_15939);
nor U17080 (N_17080,N_16310,N_16682);
and U17081 (N_17081,N_16119,N_16154);
xor U17082 (N_17082,N_16446,N_16378);
and U17083 (N_17083,N_16631,N_16730);
and U17084 (N_17084,N_15981,N_16377);
nand U17085 (N_17085,N_16304,N_16754);
nor U17086 (N_17086,N_16566,N_16083);
or U17087 (N_17087,N_16485,N_15779);
nand U17088 (N_17088,N_16068,N_16075);
xnor U17089 (N_17089,N_16580,N_15836);
xnor U17090 (N_17090,N_16713,N_16267);
xnor U17091 (N_17091,N_16279,N_15875);
and U17092 (N_17092,N_15882,N_16536);
and U17093 (N_17093,N_15903,N_15638);
or U17094 (N_17094,N_16517,N_16273);
xnor U17095 (N_17095,N_15957,N_16292);
nand U17096 (N_17096,N_15716,N_16275);
or U17097 (N_17097,N_16266,N_15906);
nor U17098 (N_17098,N_16234,N_15899);
xor U17099 (N_17099,N_15883,N_16715);
nand U17100 (N_17100,N_15804,N_16694);
or U17101 (N_17101,N_16022,N_15946);
nand U17102 (N_17102,N_15772,N_16379);
or U17103 (N_17103,N_16519,N_15839);
and U17104 (N_17104,N_16219,N_16633);
nand U17105 (N_17105,N_16020,N_15723);
nor U17106 (N_17106,N_15992,N_16490);
nand U17107 (N_17107,N_15721,N_15840);
nor U17108 (N_17108,N_16330,N_15627);
xnor U17109 (N_17109,N_16626,N_16693);
xnor U17110 (N_17110,N_16620,N_16771);
or U17111 (N_17111,N_16555,N_16363);
and U17112 (N_17112,N_16535,N_15997);
nand U17113 (N_17113,N_16564,N_16011);
or U17114 (N_17114,N_16619,N_16448);
nand U17115 (N_17115,N_16120,N_15736);
or U17116 (N_17116,N_16315,N_16192);
nor U17117 (N_17117,N_16026,N_15626);
nand U17118 (N_17118,N_16065,N_15641);
nor U17119 (N_17119,N_16493,N_16642);
and U17120 (N_17120,N_15652,N_15681);
nand U17121 (N_17121,N_16795,N_16359);
nand U17122 (N_17122,N_15912,N_16091);
xor U17123 (N_17123,N_15743,N_16371);
nand U17124 (N_17124,N_16233,N_16106);
xor U17125 (N_17125,N_16685,N_16012);
and U17126 (N_17126,N_15786,N_16687);
and U17127 (N_17127,N_15889,N_16238);
xor U17128 (N_17128,N_16278,N_16004);
xor U17129 (N_17129,N_16168,N_16692);
nand U17130 (N_17130,N_16689,N_16717);
nand U17131 (N_17131,N_15783,N_16297);
nand U17132 (N_17132,N_16787,N_16074);
nor U17133 (N_17133,N_16558,N_16452);
and U17134 (N_17134,N_16486,N_16585);
or U17135 (N_17135,N_15613,N_15869);
or U17136 (N_17136,N_16221,N_16272);
or U17137 (N_17137,N_16738,N_16081);
nand U17138 (N_17138,N_16029,N_16720);
or U17139 (N_17139,N_16381,N_16169);
nor U17140 (N_17140,N_15969,N_16443);
xor U17141 (N_17141,N_16222,N_15714);
nand U17142 (N_17142,N_16623,N_16340);
xor U17143 (N_17143,N_16395,N_15816);
nand U17144 (N_17144,N_15919,N_16627);
nor U17145 (N_17145,N_16394,N_15698);
xor U17146 (N_17146,N_16551,N_16652);
and U17147 (N_17147,N_15741,N_16353);
xnor U17148 (N_17148,N_16648,N_16255);
xnor U17149 (N_17149,N_16196,N_16204);
xor U17150 (N_17150,N_15916,N_15897);
xor U17151 (N_17151,N_16437,N_16370);
and U17152 (N_17152,N_16471,N_15922);
or U17153 (N_17153,N_15961,N_16407);
and U17154 (N_17154,N_16792,N_16450);
nand U17155 (N_17155,N_16269,N_15898);
nand U17156 (N_17156,N_16139,N_15609);
nor U17157 (N_17157,N_15807,N_16319);
nor U17158 (N_17158,N_16421,N_15635);
xor U17159 (N_17159,N_15700,N_15664);
or U17160 (N_17160,N_16520,N_16467);
or U17161 (N_17161,N_16758,N_16581);
nor U17162 (N_17162,N_16573,N_16014);
or U17163 (N_17163,N_15888,N_15918);
nand U17164 (N_17164,N_16789,N_16241);
nor U17165 (N_17165,N_15843,N_16207);
and U17166 (N_17166,N_16142,N_15979);
and U17167 (N_17167,N_16658,N_15674);
xnor U17168 (N_17168,N_15765,N_15930);
xor U17169 (N_17169,N_16424,N_15844);
nand U17170 (N_17170,N_16615,N_16327);
and U17171 (N_17171,N_16038,N_16149);
or U17172 (N_17172,N_16208,N_16757);
and U17173 (N_17173,N_15850,N_15990);
nand U17174 (N_17174,N_16250,N_15647);
nor U17175 (N_17175,N_16153,N_15864);
nand U17176 (N_17176,N_16763,N_16526);
nand U17177 (N_17177,N_15760,N_16752);
xnor U17178 (N_17178,N_16665,N_16118);
xor U17179 (N_17179,N_16086,N_16194);
or U17180 (N_17180,N_16529,N_16675);
xor U17181 (N_17181,N_16045,N_15702);
xor U17182 (N_17182,N_16172,N_15686);
nor U17183 (N_17183,N_16645,N_15704);
nand U17184 (N_17184,N_15885,N_16762);
xnor U17185 (N_17185,N_16505,N_16387);
or U17186 (N_17186,N_16338,N_16042);
or U17187 (N_17187,N_16006,N_16303);
and U17188 (N_17188,N_16160,N_15633);
nand U17189 (N_17189,N_16606,N_16475);
nor U17190 (N_17190,N_16016,N_15920);
nand U17191 (N_17191,N_15895,N_16732);
and U17192 (N_17192,N_16634,N_15943);
xnor U17193 (N_17193,N_15688,N_16177);
nand U17194 (N_17194,N_16337,N_15646);
or U17195 (N_17195,N_16024,N_16129);
xnor U17196 (N_17196,N_16288,N_16733);
or U17197 (N_17197,N_16454,N_16314);
nand U17198 (N_17198,N_16225,N_15820);
nand U17199 (N_17199,N_16021,N_16608);
nor U17200 (N_17200,N_16133,N_16788);
nor U17201 (N_17201,N_16290,N_15856);
xnor U17202 (N_17202,N_16533,N_16746);
and U17203 (N_17203,N_15673,N_15847);
and U17204 (N_17204,N_15662,N_15733);
or U17205 (N_17205,N_16244,N_16644);
or U17206 (N_17206,N_15657,N_15761);
nor U17207 (N_17207,N_15608,N_16100);
xor U17208 (N_17208,N_16282,N_16688);
nor U17209 (N_17209,N_16152,N_16494);
nor U17210 (N_17210,N_16035,N_16206);
nand U17211 (N_17211,N_16609,N_15960);
xor U17212 (N_17212,N_15746,N_15937);
xor U17213 (N_17213,N_16109,N_16057);
or U17214 (N_17214,N_16544,N_16565);
or U17215 (N_17215,N_16366,N_16432);
and U17216 (N_17216,N_16510,N_16036);
nand U17217 (N_17217,N_15748,N_15810);
xnor U17218 (N_17218,N_16002,N_16473);
nor U17219 (N_17219,N_16305,N_16406);
and U17220 (N_17220,N_15691,N_16797);
nor U17221 (N_17221,N_16183,N_15892);
nand U17222 (N_17222,N_15722,N_16790);
or U17223 (N_17223,N_16668,N_16331);
xor U17224 (N_17224,N_16679,N_16547);
and U17225 (N_17225,N_16491,N_16163);
and U17226 (N_17226,N_16098,N_15658);
xor U17227 (N_17227,N_15823,N_16343);
or U17228 (N_17228,N_16325,N_15876);
xor U17229 (N_17229,N_15948,N_15773);
or U17230 (N_17230,N_15966,N_16104);
or U17231 (N_17231,N_16588,N_15998);
and U17232 (N_17232,N_15863,N_16203);
or U17233 (N_17233,N_15945,N_16274);
nand U17234 (N_17234,N_15701,N_15859);
nor U17235 (N_17235,N_15797,N_15886);
nand U17236 (N_17236,N_15932,N_16019);
xor U17237 (N_17237,N_16534,N_16117);
and U17238 (N_17238,N_15753,N_16336);
nor U17239 (N_17239,N_16594,N_15729);
or U17240 (N_17240,N_16147,N_15891);
xnor U17241 (N_17241,N_16661,N_16691);
or U17242 (N_17242,N_16048,N_16796);
and U17243 (N_17243,N_16070,N_15669);
and U17244 (N_17244,N_16268,N_16622);
and U17245 (N_17245,N_16436,N_15870);
nor U17246 (N_17246,N_16587,N_16718);
and U17247 (N_17247,N_16499,N_15745);
nor U17248 (N_17248,N_16280,N_16339);
nand U17249 (N_17249,N_15954,N_16597);
or U17250 (N_17250,N_16262,N_16476);
nor U17251 (N_17251,N_16193,N_15696);
and U17252 (N_17252,N_16232,N_16712);
xor U17253 (N_17253,N_15915,N_16361);
xnor U17254 (N_17254,N_15659,N_16670);
or U17255 (N_17255,N_15858,N_15717);
and U17256 (N_17256,N_16703,N_16171);
nand U17257 (N_17257,N_16313,N_16664);
xnor U17258 (N_17258,N_15975,N_16166);
nor U17259 (N_17259,N_16046,N_16384);
nor U17260 (N_17260,N_15802,N_15933);
xnor U17261 (N_17261,N_16231,N_15793);
xnor U17262 (N_17262,N_16093,N_16126);
nand U17263 (N_17263,N_16362,N_16635);
and U17264 (N_17264,N_16392,N_15986);
xor U17265 (N_17265,N_16135,N_16590);
nand U17266 (N_17266,N_15841,N_15642);
nor U17267 (N_17267,N_15952,N_15766);
xor U17268 (N_17268,N_16248,N_15690);
xnor U17269 (N_17269,N_16076,N_15838);
nor U17270 (N_17270,N_15988,N_15900);
nor U17271 (N_17271,N_15639,N_16578);
or U17272 (N_17272,N_16348,N_16560);
or U17273 (N_17273,N_16191,N_15955);
and U17274 (N_17274,N_16767,N_16727);
nor U17275 (N_17275,N_16791,N_16599);
xor U17276 (N_17276,N_15602,N_16561);
and U17277 (N_17277,N_15989,N_16640);
and U17278 (N_17278,N_15987,N_15805);
and U17279 (N_17279,N_16638,N_16538);
or U17280 (N_17280,N_15737,N_15973);
and U17281 (N_17281,N_16254,N_16329);
nor U17282 (N_17282,N_16113,N_16412);
nor U17283 (N_17283,N_16060,N_15848);
xor U17284 (N_17284,N_16572,N_16769);
nor U17285 (N_17285,N_15708,N_15878);
xnor U17286 (N_17286,N_16346,N_15758);
or U17287 (N_17287,N_15857,N_16054);
or U17288 (N_17288,N_15855,N_16187);
xor U17289 (N_17289,N_16051,N_16218);
and U17290 (N_17290,N_16242,N_16495);
nor U17291 (N_17291,N_16770,N_15612);
nor U17292 (N_17292,N_16064,N_15750);
xnor U17293 (N_17293,N_16003,N_15927);
or U17294 (N_17294,N_16481,N_16037);
or U17295 (N_17295,N_16613,N_16438);
and U17296 (N_17296,N_16328,N_16427);
or U17297 (N_17297,N_16410,N_16681);
xor U17298 (N_17298,N_16252,N_15852);
nand U17299 (N_17299,N_16216,N_15682);
or U17300 (N_17300,N_15936,N_15771);
nand U17301 (N_17301,N_15831,N_16772);
nor U17302 (N_17302,N_16643,N_16140);
and U17303 (N_17303,N_16071,N_16699);
or U17304 (N_17304,N_16375,N_16650);
nor U17305 (N_17305,N_16320,N_15884);
or U17306 (N_17306,N_16464,N_16047);
nand U17307 (N_17307,N_15731,N_15675);
nand U17308 (N_17308,N_15846,N_16741);
or U17309 (N_17309,N_15778,N_16724);
and U17310 (N_17310,N_16105,N_16000);
xor U17311 (N_17311,N_16453,N_16365);
or U17312 (N_17312,N_16227,N_16600);
nor U17313 (N_17313,N_16527,N_16728);
nand U17314 (N_17314,N_15727,N_16408);
or U17315 (N_17315,N_15947,N_16388);
nor U17316 (N_17316,N_15896,N_16013);
nor U17317 (N_17317,N_15709,N_15678);
xor U17318 (N_17318,N_15776,N_16461);
and U17319 (N_17319,N_16725,N_16059);
nand U17320 (N_17320,N_16261,N_16333);
nor U17321 (N_17321,N_15757,N_16326);
or U17322 (N_17322,N_15929,N_16009);
nand U17323 (N_17323,N_15734,N_16195);
nor U17324 (N_17324,N_16145,N_16428);
or U17325 (N_17325,N_16124,N_16210);
nor U17326 (N_17326,N_16116,N_16150);
or U17327 (N_17327,N_16562,N_16696);
nand U17328 (N_17328,N_16678,N_15763);
nor U17329 (N_17329,N_16302,N_15833);
or U17330 (N_17330,N_16576,N_16440);
nor U17331 (N_17331,N_16271,N_15894);
nand U17332 (N_17332,N_16307,N_16605);
or U17333 (N_17333,N_16352,N_15606);
nand U17334 (N_17334,N_16630,N_16429);
nand U17335 (N_17335,N_16487,N_15679);
xor U17336 (N_17336,N_16657,N_16532);
or U17337 (N_17337,N_16470,N_16405);
or U17338 (N_17338,N_15655,N_16276);
and U17339 (N_17339,N_16647,N_16618);
xor U17340 (N_17340,N_16602,N_16512);
xnor U17341 (N_17341,N_15654,N_16249);
nor U17342 (N_17342,N_15806,N_16239);
or U17343 (N_17343,N_15703,N_15867);
xor U17344 (N_17344,N_15909,N_16088);
xor U17345 (N_17345,N_16281,N_15769);
xor U17346 (N_17346,N_15798,N_16501);
nor U17347 (N_17347,N_16612,N_15931);
and U17348 (N_17348,N_16128,N_16108);
nand U17349 (N_17349,N_15974,N_16777);
nand U17350 (N_17350,N_15830,N_15911);
nand U17351 (N_17351,N_15905,N_15720);
xnor U17352 (N_17352,N_16755,N_15619);
xor U17353 (N_17353,N_16660,N_16179);
or U17354 (N_17354,N_16574,N_15925);
and U17355 (N_17355,N_16459,N_16354);
or U17356 (N_17356,N_16662,N_16096);
xnor U17357 (N_17357,N_16164,N_16506);
nor U17358 (N_17358,N_15628,N_15705);
or U17359 (N_17359,N_15881,N_16411);
nor U17360 (N_17360,N_16434,N_15742);
nand U17361 (N_17361,N_16614,N_16213);
or U17362 (N_17362,N_16545,N_16554);
nand U17363 (N_17363,N_16726,N_16132);
and U17364 (N_17364,N_15767,N_15949);
and U17365 (N_17365,N_16085,N_16632);
nor U17366 (N_17366,N_15747,N_16099);
xnor U17367 (N_17367,N_16624,N_16176);
nand U17368 (N_17368,N_16323,N_15921);
and U17369 (N_17369,N_16761,N_16497);
xnor U17370 (N_17370,N_16316,N_16457);
or U17371 (N_17371,N_15725,N_16708);
xnor U17372 (N_17372,N_16779,N_15621);
xnor U17373 (N_17373,N_16159,N_16200);
nand U17374 (N_17374,N_15822,N_16050);
and U17375 (N_17375,N_16477,N_16214);
nand U17376 (N_17376,N_16095,N_16546);
nor U17377 (N_17377,N_15604,N_16170);
and U17378 (N_17378,N_15970,N_16215);
nor U17379 (N_17379,N_16628,N_15666);
and U17380 (N_17380,N_15962,N_16131);
and U17381 (N_17381,N_16480,N_15958);
nor U17382 (N_17382,N_16165,N_15694);
xor U17383 (N_17383,N_16604,N_16702);
and U17384 (N_17384,N_15632,N_15995);
nand U17385 (N_17385,N_16197,N_16508);
nand U17386 (N_17386,N_15730,N_16342);
or U17387 (N_17387,N_16018,N_15789);
nor U17388 (N_17388,N_16584,N_16134);
or U17389 (N_17389,N_16719,N_15644);
or U17390 (N_17390,N_15650,N_16090);
nand U17391 (N_17391,N_15660,N_15755);
or U17392 (N_17392,N_15791,N_16052);
nand U17393 (N_17393,N_16181,N_16582);
and U17394 (N_17394,N_15637,N_16174);
nor U17395 (N_17395,N_16039,N_15649);
nor U17396 (N_17396,N_16146,N_15794);
nor U17397 (N_17397,N_16212,N_16258);
xnor U17398 (N_17398,N_16344,N_16350);
nand U17399 (N_17399,N_16714,N_16684);
xnor U17400 (N_17400,N_15897,N_16158);
xor U17401 (N_17401,N_15736,N_16632);
nor U17402 (N_17402,N_16329,N_16389);
xnor U17403 (N_17403,N_16440,N_16449);
xnor U17404 (N_17404,N_16132,N_16409);
nor U17405 (N_17405,N_15846,N_16075);
xor U17406 (N_17406,N_16130,N_16020);
nor U17407 (N_17407,N_16499,N_15782);
xor U17408 (N_17408,N_16769,N_16017);
nor U17409 (N_17409,N_15797,N_15726);
xnor U17410 (N_17410,N_16279,N_16021);
nor U17411 (N_17411,N_16131,N_15752);
nor U17412 (N_17412,N_15802,N_16759);
nand U17413 (N_17413,N_16206,N_15692);
or U17414 (N_17414,N_16666,N_15662);
nand U17415 (N_17415,N_16284,N_15837);
xnor U17416 (N_17416,N_16671,N_16122);
and U17417 (N_17417,N_16708,N_16196);
xor U17418 (N_17418,N_16752,N_15812);
nand U17419 (N_17419,N_16466,N_16572);
nand U17420 (N_17420,N_16637,N_15923);
or U17421 (N_17421,N_16374,N_16435);
or U17422 (N_17422,N_16024,N_16647);
xor U17423 (N_17423,N_16121,N_16387);
nor U17424 (N_17424,N_15765,N_15766);
and U17425 (N_17425,N_16464,N_16114);
nand U17426 (N_17426,N_15670,N_16238);
and U17427 (N_17427,N_16178,N_16373);
nand U17428 (N_17428,N_15697,N_15617);
nor U17429 (N_17429,N_16112,N_16480);
nor U17430 (N_17430,N_16296,N_16684);
and U17431 (N_17431,N_15961,N_16474);
nor U17432 (N_17432,N_16426,N_16789);
and U17433 (N_17433,N_16684,N_16506);
nand U17434 (N_17434,N_16074,N_16518);
or U17435 (N_17435,N_16053,N_15681);
and U17436 (N_17436,N_15752,N_15685);
xor U17437 (N_17437,N_15937,N_15871);
xor U17438 (N_17438,N_16437,N_16450);
xor U17439 (N_17439,N_15968,N_16388);
and U17440 (N_17440,N_15968,N_16489);
xor U17441 (N_17441,N_15934,N_15676);
nand U17442 (N_17442,N_16329,N_16175);
and U17443 (N_17443,N_15647,N_16078);
nor U17444 (N_17444,N_16738,N_16238);
and U17445 (N_17445,N_15957,N_16131);
and U17446 (N_17446,N_16726,N_16343);
xor U17447 (N_17447,N_16254,N_16424);
nor U17448 (N_17448,N_16343,N_16614);
nor U17449 (N_17449,N_16710,N_16111);
xnor U17450 (N_17450,N_16696,N_15943);
xor U17451 (N_17451,N_15892,N_16277);
nand U17452 (N_17452,N_16417,N_16657);
and U17453 (N_17453,N_15883,N_15945);
nor U17454 (N_17454,N_16631,N_16105);
and U17455 (N_17455,N_16563,N_16358);
or U17456 (N_17456,N_16338,N_15651);
and U17457 (N_17457,N_16577,N_16138);
and U17458 (N_17458,N_16156,N_15963);
xnor U17459 (N_17459,N_16736,N_16182);
or U17460 (N_17460,N_16770,N_16063);
nand U17461 (N_17461,N_16688,N_15673);
or U17462 (N_17462,N_15918,N_16207);
nand U17463 (N_17463,N_16577,N_15636);
and U17464 (N_17464,N_16773,N_16200);
nand U17465 (N_17465,N_16740,N_16100);
nand U17466 (N_17466,N_16505,N_16642);
nand U17467 (N_17467,N_15978,N_16076);
and U17468 (N_17468,N_15965,N_15653);
xor U17469 (N_17469,N_16605,N_16187);
or U17470 (N_17470,N_16017,N_16648);
and U17471 (N_17471,N_16384,N_16416);
or U17472 (N_17472,N_16334,N_15661);
and U17473 (N_17473,N_16395,N_16192);
xnor U17474 (N_17474,N_16234,N_16220);
and U17475 (N_17475,N_16360,N_16747);
nor U17476 (N_17476,N_16022,N_16091);
and U17477 (N_17477,N_15927,N_16244);
xnor U17478 (N_17478,N_16094,N_16530);
nor U17479 (N_17479,N_16123,N_16074);
nand U17480 (N_17480,N_16655,N_15951);
xor U17481 (N_17481,N_16511,N_16489);
and U17482 (N_17482,N_16365,N_16108);
and U17483 (N_17483,N_16263,N_16383);
nor U17484 (N_17484,N_16478,N_15930);
xnor U17485 (N_17485,N_15830,N_16355);
or U17486 (N_17486,N_16342,N_15911);
xor U17487 (N_17487,N_15867,N_16483);
or U17488 (N_17488,N_16397,N_16518);
xnor U17489 (N_17489,N_16756,N_16340);
nand U17490 (N_17490,N_16148,N_16162);
xnor U17491 (N_17491,N_16673,N_16786);
and U17492 (N_17492,N_16575,N_16448);
or U17493 (N_17493,N_15812,N_16095);
nor U17494 (N_17494,N_16049,N_16036);
nor U17495 (N_17495,N_15735,N_16390);
xor U17496 (N_17496,N_15856,N_15680);
nor U17497 (N_17497,N_15675,N_15912);
or U17498 (N_17498,N_16251,N_15700);
or U17499 (N_17499,N_16066,N_15930);
and U17500 (N_17500,N_16024,N_16109);
and U17501 (N_17501,N_15733,N_15812);
nand U17502 (N_17502,N_16287,N_16498);
or U17503 (N_17503,N_16607,N_16181);
and U17504 (N_17504,N_16273,N_15895);
nor U17505 (N_17505,N_16557,N_15839);
xnor U17506 (N_17506,N_16669,N_16069);
xor U17507 (N_17507,N_16753,N_15806);
nand U17508 (N_17508,N_15756,N_16450);
xnor U17509 (N_17509,N_15664,N_16751);
xor U17510 (N_17510,N_15651,N_16395);
and U17511 (N_17511,N_15854,N_15951);
and U17512 (N_17512,N_15973,N_16013);
nor U17513 (N_17513,N_16219,N_16569);
or U17514 (N_17514,N_16523,N_16553);
or U17515 (N_17515,N_16006,N_15831);
and U17516 (N_17516,N_16191,N_16048);
xor U17517 (N_17517,N_15869,N_16292);
xnor U17518 (N_17518,N_16342,N_16515);
nand U17519 (N_17519,N_16431,N_16008);
and U17520 (N_17520,N_15758,N_16002);
or U17521 (N_17521,N_15858,N_16469);
or U17522 (N_17522,N_15970,N_16564);
nand U17523 (N_17523,N_16295,N_15866);
nand U17524 (N_17524,N_15941,N_15774);
nor U17525 (N_17525,N_16653,N_16136);
xnor U17526 (N_17526,N_16581,N_16611);
nor U17527 (N_17527,N_16204,N_16496);
xor U17528 (N_17528,N_16491,N_15937);
nor U17529 (N_17529,N_16004,N_16730);
nand U17530 (N_17530,N_15903,N_16010);
or U17531 (N_17531,N_16526,N_16558);
nor U17532 (N_17532,N_16356,N_16135);
and U17533 (N_17533,N_15639,N_15953);
or U17534 (N_17534,N_16476,N_15867);
nor U17535 (N_17535,N_16633,N_15672);
xnor U17536 (N_17536,N_16221,N_15972);
nand U17537 (N_17537,N_15837,N_16197);
or U17538 (N_17538,N_16403,N_15755);
xnor U17539 (N_17539,N_16660,N_16352);
nor U17540 (N_17540,N_15910,N_16409);
nor U17541 (N_17541,N_15963,N_15739);
nand U17542 (N_17542,N_16729,N_16726);
or U17543 (N_17543,N_16376,N_16790);
or U17544 (N_17544,N_16426,N_16743);
nand U17545 (N_17545,N_15799,N_16644);
and U17546 (N_17546,N_15782,N_15830);
and U17547 (N_17547,N_16425,N_15850);
or U17548 (N_17548,N_15663,N_15664);
or U17549 (N_17549,N_16481,N_15816);
nand U17550 (N_17550,N_16710,N_16487);
nor U17551 (N_17551,N_16528,N_15955);
xnor U17552 (N_17552,N_16118,N_16610);
xnor U17553 (N_17553,N_15885,N_16243);
and U17554 (N_17554,N_16263,N_15835);
nand U17555 (N_17555,N_15655,N_15818);
nand U17556 (N_17556,N_15972,N_15897);
xnor U17557 (N_17557,N_15835,N_16515);
xnor U17558 (N_17558,N_16470,N_16423);
nand U17559 (N_17559,N_16148,N_16458);
nor U17560 (N_17560,N_16043,N_15776);
xor U17561 (N_17561,N_16314,N_15896);
nand U17562 (N_17562,N_16029,N_16743);
or U17563 (N_17563,N_15806,N_15890);
nand U17564 (N_17564,N_16327,N_16428);
xnor U17565 (N_17565,N_16166,N_15616);
or U17566 (N_17566,N_16463,N_16154);
nand U17567 (N_17567,N_15817,N_15746);
or U17568 (N_17568,N_15835,N_16478);
or U17569 (N_17569,N_15769,N_15753);
nor U17570 (N_17570,N_16140,N_16426);
and U17571 (N_17571,N_15782,N_15909);
and U17572 (N_17572,N_16797,N_16305);
nand U17573 (N_17573,N_15684,N_16241);
nor U17574 (N_17574,N_16360,N_15600);
nand U17575 (N_17575,N_15927,N_16147);
or U17576 (N_17576,N_16515,N_16560);
xnor U17577 (N_17577,N_16445,N_16365);
or U17578 (N_17578,N_15680,N_15830);
or U17579 (N_17579,N_16082,N_16551);
and U17580 (N_17580,N_16651,N_15758);
nor U17581 (N_17581,N_15872,N_16273);
nand U17582 (N_17582,N_16620,N_15716);
nor U17583 (N_17583,N_16748,N_15641);
xnor U17584 (N_17584,N_15739,N_15887);
and U17585 (N_17585,N_16623,N_16395);
nor U17586 (N_17586,N_15687,N_16251);
or U17587 (N_17587,N_16110,N_15981);
nand U17588 (N_17588,N_16069,N_16130);
and U17589 (N_17589,N_16529,N_15923);
nor U17590 (N_17590,N_15615,N_16087);
xnor U17591 (N_17591,N_16655,N_15768);
nand U17592 (N_17592,N_15993,N_16476);
xor U17593 (N_17593,N_16197,N_16531);
nor U17594 (N_17594,N_16331,N_16233);
nor U17595 (N_17595,N_16245,N_15821);
nor U17596 (N_17596,N_16581,N_15886);
or U17597 (N_17597,N_15975,N_16079);
xnor U17598 (N_17598,N_15971,N_16354);
xnor U17599 (N_17599,N_16137,N_16584);
xnor U17600 (N_17600,N_15899,N_15705);
xnor U17601 (N_17601,N_15706,N_16425);
xnor U17602 (N_17602,N_15850,N_16392);
nand U17603 (N_17603,N_15750,N_16735);
or U17604 (N_17604,N_15689,N_16379);
nand U17605 (N_17605,N_16725,N_16685);
nor U17606 (N_17606,N_16552,N_15855);
nand U17607 (N_17607,N_15974,N_15720);
nand U17608 (N_17608,N_16270,N_16686);
nor U17609 (N_17609,N_15651,N_15791);
nor U17610 (N_17610,N_16123,N_15812);
and U17611 (N_17611,N_15793,N_15765);
xor U17612 (N_17612,N_16527,N_16128);
nand U17613 (N_17613,N_16192,N_15921);
or U17614 (N_17614,N_15663,N_16539);
and U17615 (N_17615,N_16788,N_15619);
nand U17616 (N_17616,N_16237,N_16426);
and U17617 (N_17617,N_16622,N_16346);
and U17618 (N_17618,N_15858,N_16182);
or U17619 (N_17619,N_16268,N_16645);
nor U17620 (N_17620,N_15719,N_16144);
xnor U17621 (N_17621,N_16263,N_16555);
and U17622 (N_17622,N_16049,N_15863);
and U17623 (N_17623,N_15813,N_16106);
xnor U17624 (N_17624,N_16530,N_16248);
or U17625 (N_17625,N_16499,N_16760);
or U17626 (N_17626,N_15649,N_16074);
nand U17627 (N_17627,N_15712,N_16155);
or U17628 (N_17628,N_15674,N_16789);
nor U17629 (N_17629,N_16032,N_16727);
nor U17630 (N_17630,N_16235,N_16588);
and U17631 (N_17631,N_15956,N_15929);
xor U17632 (N_17632,N_15692,N_16332);
nor U17633 (N_17633,N_16405,N_16733);
or U17634 (N_17634,N_16734,N_16487);
or U17635 (N_17635,N_15810,N_15838);
and U17636 (N_17636,N_16629,N_15708);
nand U17637 (N_17637,N_16766,N_16463);
or U17638 (N_17638,N_16713,N_15927);
or U17639 (N_17639,N_16282,N_16109);
nand U17640 (N_17640,N_16373,N_16218);
xnor U17641 (N_17641,N_16590,N_16779);
nand U17642 (N_17642,N_15624,N_16699);
or U17643 (N_17643,N_16754,N_16009);
and U17644 (N_17644,N_15762,N_16719);
xnor U17645 (N_17645,N_15846,N_16069);
or U17646 (N_17646,N_15803,N_15787);
or U17647 (N_17647,N_16260,N_16449);
nor U17648 (N_17648,N_15931,N_16463);
nor U17649 (N_17649,N_15945,N_16323);
xnor U17650 (N_17650,N_16360,N_16059);
or U17651 (N_17651,N_15873,N_16461);
nor U17652 (N_17652,N_16033,N_16455);
nand U17653 (N_17653,N_16248,N_16376);
xor U17654 (N_17654,N_16663,N_16222);
or U17655 (N_17655,N_16450,N_15823);
nor U17656 (N_17656,N_15885,N_16349);
xor U17657 (N_17657,N_15909,N_16018);
nand U17658 (N_17658,N_16051,N_16048);
nand U17659 (N_17659,N_16111,N_15667);
nand U17660 (N_17660,N_16343,N_16321);
nand U17661 (N_17661,N_16646,N_16308);
nor U17662 (N_17662,N_16207,N_16108);
nor U17663 (N_17663,N_16442,N_16320);
xnor U17664 (N_17664,N_15715,N_16147);
nor U17665 (N_17665,N_16199,N_16435);
or U17666 (N_17666,N_16668,N_15899);
nor U17667 (N_17667,N_15675,N_16723);
nor U17668 (N_17668,N_16663,N_15835);
or U17669 (N_17669,N_16416,N_16207);
and U17670 (N_17670,N_16718,N_15810);
xor U17671 (N_17671,N_16495,N_16635);
or U17672 (N_17672,N_16297,N_16414);
nand U17673 (N_17673,N_16358,N_15775);
or U17674 (N_17674,N_16344,N_16031);
nor U17675 (N_17675,N_16725,N_15625);
or U17676 (N_17676,N_16095,N_16636);
nor U17677 (N_17677,N_16050,N_16342);
or U17678 (N_17678,N_16415,N_15667);
xor U17679 (N_17679,N_16735,N_15821);
and U17680 (N_17680,N_16216,N_15921);
nand U17681 (N_17681,N_16378,N_15607);
xnor U17682 (N_17682,N_15995,N_16236);
nand U17683 (N_17683,N_16201,N_16008);
nor U17684 (N_17684,N_16677,N_16126);
nor U17685 (N_17685,N_16482,N_16577);
nand U17686 (N_17686,N_15951,N_16680);
nor U17687 (N_17687,N_16499,N_16130);
xnor U17688 (N_17688,N_16660,N_16149);
and U17689 (N_17689,N_16032,N_16531);
and U17690 (N_17690,N_15749,N_16604);
nor U17691 (N_17691,N_16399,N_16473);
and U17692 (N_17692,N_16107,N_16122);
nand U17693 (N_17693,N_16452,N_16646);
nor U17694 (N_17694,N_16051,N_16519);
nor U17695 (N_17695,N_16406,N_15881);
or U17696 (N_17696,N_15979,N_16424);
xor U17697 (N_17697,N_15912,N_15902);
and U17698 (N_17698,N_16352,N_15781);
xor U17699 (N_17699,N_16194,N_15973);
nor U17700 (N_17700,N_16715,N_16174);
and U17701 (N_17701,N_16137,N_15628);
xor U17702 (N_17702,N_16681,N_16544);
nand U17703 (N_17703,N_15885,N_16109);
nor U17704 (N_17704,N_16369,N_15804);
or U17705 (N_17705,N_15750,N_16561);
nor U17706 (N_17706,N_16362,N_16014);
xnor U17707 (N_17707,N_16532,N_16055);
xnor U17708 (N_17708,N_15954,N_15738);
and U17709 (N_17709,N_16387,N_16319);
or U17710 (N_17710,N_16321,N_16791);
nand U17711 (N_17711,N_15935,N_15602);
xnor U17712 (N_17712,N_15803,N_15660);
or U17713 (N_17713,N_16046,N_16123);
or U17714 (N_17714,N_16682,N_15645);
or U17715 (N_17715,N_16215,N_15853);
nor U17716 (N_17716,N_15824,N_16597);
nor U17717 (N_17717,N_16277,N_15891);
nand U17718 (N_17718,N_16406,N_15741);
or U17719 (N_17719,N_16343,N_16431);
and U17720 (N_17720,N_15817,N_16038);
nand U17721 (N_17721,N_16793,N_16790);
xnor U17722 (N_17722,N_16465,N_16188);
or U17723 (N_17723,N_16589,N_16067);
xnor U17724 (N_17724,N_16409,N_16730);
or U17725 (N_17725,N_16237,N_16350);
or U17726 (N_17726,N_15796,N_16664);
nor U17727 (N_17727,N_16401,N_16690);
nand U17728 (N_17728,N_15955,N_15823);
nor U17729 (N_17729,N_16578,N_16642);
nand U17730 (N_17730,N_16150,N_15695);
or U17731 (N_17731,N_16321,N_15646);
nand U17732 (N_17732,N_16626,N_15922);
and U17733 (N_17733,N_16358,N_15942);
nand U17734 (N_17734,N_15837,N_16413);
or U17735 (N_17735,N_16558,N_16601);
and U17736 (N_17736,N_16616,N_16182);
nand U17737 (N_17737,N_15668,N_16317);
and U17738 (N_17738,N_15829,N_16034);
nor U17739 (N_17739,N_16104,N_16431);
xnor U17740 (N_17740,N_16382,N_16134);
nand U17741 (N_17741,N_16234,N_15858);
or U17742 (N_17742,N_16139,N_15698);
nor U17743 (N_17743,N_16422,N_16331);
nand U17744 (N_17744,N_16372,N_15695);
nand U17745 (N_17745,N_15815,N_15771);
and U17746 (N_17746,N_16099,N_16439);
nand U17747 (N_17747,N_16639,N_16027);
xor U17748 (N_17748,N_16652,N_16504);
nor U17749 (N_17749,N_15683,N_16721);
xor U17750 (N_17750,N_15839,N_15619);
xnor U17751 (N_17751,N_15929,N_16064);
nand U17752 (N_17752,N_16558,N_15720);
xnor U17753 (N_17753,N_15688,N_16051);
nand U17754 (N_17754,N_16677,N_16541);
or U17755 (N_17755,N_15872,N_16060);
nor U17756 (N_17756,N_16241,N_16143);
xor U17757 (N_17757,N_16177,N_15617);
and U17758 (N_17758,N_16283,N_16090);
and U17759 (N_17759,N_16413,N_16669);
xor U17760 (N_17760,N_16387,N_16214);
xor U17761 (N_17761,N_16427,N_15879);
nand U17762 (N_17762,N_15718,N_16532);
nand U17763 (N_17763,N_16585,N_16012);
or U17764 (N_17764,N_16628,N_15912);
nand U17765 (N_17765,N_15644,N_16360);
xor U17766 (N_17766,N_16536,N_16296);
and U17767 (N_17767,N_16775,N_15920);
xor U17768 (N_17768,N_16205,N_16469);
xor U17769 (N_17769,N_15749,N_16047);
and U17770 (N_17770,N_16797,N_16637);
xnor U17771 (N_17771,N_16517,N_16143);
nand U17772 (N_17772,N_15645,N_15736);
and U17773 (N_17773,N_15659,N_16329);
nor U17774 (N_17774,N_15750,N_15974);
nand U17775 (N_17775,N_16057,N_16630);
or U17776 (N_17776,N_15869,N_16526);
xnor U17777 (N_17777,N_16691,N_15695);
or U17778 (N_17778,N_15732,N_15760);
nand U17779 (N_17779,N_15908,N_15685);
xor U17780 (N_17780,N_16206,N_16692);
xnor U17781 (N_17781,N_16030,N_16131);
or U17782 (N_17782,N_16604,N_16442);
and U17783 (N_17783,N_15935,N_16380);
nor U17784 (N_17784,N_15653,N_16679);
and U17785 (N_17785,N_16237,N_16096);
nor U17786 (N_17786,N_15881,N_15992);
or U17787 (N_17787,N_16095,N_16084);
xor U17788 (N_17788,N_16376,N_15968);
nand U17789 (N_17789,N_15842,N_16722);
or U17790 (N_17790,N_15764,N_16631);
and U17791 (N_17791,N_16565,N_16360);
or U17792 (N_17792,N_15755,N_15993);
xnor U17793 (N_17793,N_15905,N_16074);
xnor U17794 (N_17794,N_16388,N_16162);
nand U17795 (N_17795,N_15894,N_16365);
and U17796 (N_17796,N_15985,N_16304);
or U17797 (N_17797,N_16413,N_15673);
xnor U17798 (N_17798,N_15700,N_15845);
nor U17799 (N_17799,N_16161,N_16458);
xnor U17800 (N_17800,N_15738,N_16047);
nor U17801 (N_17801,N_16096,N_16560);
xnor U17802 (N_17802,N_15956,N_16603);
xnor U17803 (N_17803,N_15845,N_16447);
and U17804 (N_17804,N_15992,N_15960);
nand U17805 (N_17805,N_15967,N_16082);
xnor U17806 (N_17806,N_15972,N_16747);
xnor U17807 (N_17807,N_16138,N_15688);
nand U17808 (N_17808,N_16394,N_16358);
and U17809 (N_17809,N_15972,N_16232);
and U17810 (N_17810,N_16778,N_15918);
or U17811 (N_17811,N_16674,N_16556);
nand U17812 (N_17812,N_16683,N_16291);
or U17813 (N_17813,N_16206,N_16236);
xor U17814 (N_17814,N_15740,N_16514);
nor U17815 (N_17815,N_15974,N_16277);
nor U17816 (N_17816,N_16122,N_16773);
and U17817 (N_17817,N_16773,N_16786);
nor U17818 (N_17818,N_16791,N_16764);
or U17819 (N_17819,N_16164,N_16290);
nand U17820 (N_17820,N_15837,N_16228);
xor U17821 (N_17821,N_16493,N_16558);
nor U17822 (N_17822,N_16209,N_15990);
and U17823 (N_17823,N_16544,N_16196);
nand U17824 (N_17824,N_16314,N_16538);
nand U17825 (N_17825,N_16571,N_16413);
or U17826 (N_17826,N_15825,N_16285);
and U17827 (N_17827,N_15787,N_16665);
and U17828 (N_17828,N_16125,N_16460);
xnor U17829 (N_17829,N_16758,N_16299);
nand U17830 (N_17830,N_16633,N_15652);
or U17831 (N_17831,N_15861,N_15690);
or U17832 (N_17832,N_15801,N_16263);
nor U17833 (N_17833,N_16080,N_16079);
xnor U17834 (N_17834,N_16772,N_16632);
xnor U17835 (N_17835,N_16293,N_16701);
nor U17836 (N_17836,N_16392,N_16475);
xor U17837 (N_17837,N_15876,N_16505);
and U17838 (N_17838,N_15786,N_16063);
and U17839 (N_17839,N_15716,N_16616);
or U17840 (N_17840,N_16001,N_16705);
or U17841 (N_17841,N_16271,N_15715);
nand U17842 (N_17842,N_16068,N_16430);
nand U17843 (N_17843,N_15872,N_15852);
or U17844 (N_17844,N_16671,N_16229);
or U17845 (N_17845,N_15895,N_15893);
or U17846 (N_17846,N_16160,N_16393);
or U17847 (N_17847,N_16311,N_16561);
xnor U17848 (N_17848,N_16408,N_16745);
nand U17849 (N_17849,N_16235,N_16063);
and U17850 (N_17850,N_16509,N_16414);
nand U17851 (N_17851,N_15640,N_15953);
nand U17852 (N_17852,N_16652,N_16701);
or U17853 (N_17853,N_16043,N_16619);
xor U17854 (N_17854,N_16100,N_16659);
and U17855 (N_17855,N_15778,N_15954);
nand U17856 (N_17856,N_16560,N_16010);
nand U17857 (N_17857,N_16473,N_15804);
or U17858 (N_17858,N_15816,N_16019);
nand U17859 (N_17859,N_16644,N_16625);
nand U17860 (N_17860,N_16682,N_15738);
and U17861 (N_17861,N_16053,N_16321);
or U17862 (N_17862,N_16277,N_16657);
xor U17863 (N_17863,N_15683,N_16758);
or U17864 (N_17864,N_16258,N_16552);
nand U17865 (N_17865,N_16073,N_16640);
nor U17866 (N_17866,N_16223,N_16176);
or U17867 (N_17867,N_16032,N_16239);
and U17868 (N_17868,N_16014,N_15701);
and U17869 (N_17869,N_16761,N_16284);
nor U17870 (N_17870,N_16492,N_15841);
xnor U17871 (N_17871,N_16533,N_16504);
xnor U17872 (N_17872,N_16366,N_16313);
nor U17873 (N_17873,N_15946,N_15944);
or U17874 (N_17874,N_16608,N_16373);
nand U17875 (N_17875,N_16076,N_15635);
and U17876 (N_17876,N_16200,N_16700);
or U17877 (N_17877,N_15610,N_16265);
and U17878 (N_17878,N_16365,N_16627);
nor U17879 (N_17879,N_15612,N_15800);
or U17880 (N_17880,N_16504,N_16142);
nand U17881 (N_17881,N_16519,N_16493);
nand U17882 (N_17882,N_16707,N_16454);
or U17883 (N_17883,N_15799,N_16635);
nand U17884 (N_17884,N_16466,N_15852);
xnor U17885 (N_17885,N_16095,N_15880);
and U17886 (N_17886,N_16075,N_16620);
and U17887 (N_17887,N_15633,N_15883);
and U17888 (N_17888,N_16683,N_16021);
or U17889 (N_17889,N_15641,N_16785);
or U17890 (N_17890,N_16615,N_16289);
nor U17891 (N_17891,N_16478,N_16262);
or U17892 (N_17892,N_15888,N_15853);
and U17893 (N_17893,N_16158,N_16083);
and U17894 (N_17894,N_16414,N_15696);
xnor U17895 (N_17895,N_15903,N_16160);
nand U17896 (N_17896,N_16668,N_15853);
or U17897 (N_17897,N_15834,N_15804);
xor U17898 (N_17898,N_16057,N_16562);
and U17899 (N_17899,N_16219,N_15863);
xnor U17900 (N_17900,N_15956,N_15817);
nor U17901 (N_17901,N_16645,N_16202);
xor U17902 (N_17902,N_16289,N_16547);
nand U17903 (N_17903,N_16493,N_15765);
nor U17904 (N_17904,N_15884,N_15908);
nor U17905 (N_17905,N_16324,N_16021);
nor U17906 (N_17906,N_15940,N_16059);
and U17907 (N_17907,N_16099,N_15905);
and U17908 (N_17908,N_15794,N_15878);
nor U17909 (N_17909,N_16360,N_16027);
and U17910 (N_17910,N_16700,N_15903);
or U17911 (N_17911,N_16292,N_16087);
nor U17912 (N_17912,N_16355,N_16085);
xor U17913 (N_17913,N_16103,N_16085);
nor U17914 (N_17914,N_15723,N_15676);
or U17915 (N_17915,N_15763,N_16673);
nor U17916 (N_17916,N_16493,N_16630);
xor U17917 (N_17917,N_15680,N_16213);
or U17918 (N_17918,N_16369,N_15772);
nor U17919 (N_17919,N_16443,N_16164);
and U17920 (N_17920,N_16211,N_16703);
xnor U17921 (N_17921,N_15621,N_16777);
and U17922 (N_17922,N_15746,N_15985);
or U17923 (N_17923,N_15852,N_16102);
xnor U17924 (N_17924,N_16680,N_16058);
xnor U17925 (N_17925,N_16103,N_15983);
and U17926 (N_17926,N_16581,N_16440);
xor U17927 (N_17927,N_16641,N_15832);
and U17928 (N_17928,N_16637,N_16359);
and U17929 (N_17929,N_15897,N_15955);
and U17930 (N_17930,N_16792,N_16138);
nor U17931 (N_17931,N_15733,N_16039);
and U17932 (N_17932,N_16242,N_16609);
or U17933 (N_17933,N_16314,N_15720);
xor U17934 (N_17934,N_15671,N_16753);
xnor U17935 (N_17935,N_16373,N_15934);
nor U17936 (N_17936,N_16042,N_15698);
and U17937 (N_17937,N_16623,N_15689);
nor U17938 (N_17938,N_15630,N_16625);
nand U17939 (N_17939,N_15761,N_16777);
xor U17940 (N_17940,N_16578,N_16483);
nand U17941 (N_17941,N_16345,N_15646);
or U17942 (N_17942,N_15637,N_15743);
or U17943 (N_17943,N_15672,N_15821);
and U17944 (N_17944,N_16195,N_16621);
and U17945 (N_17945,N_15706,N_16707);
xnor U17946 (N_17946,N_15631,N_16064);
nor U17947 (N_17947,N_15998,N_16384);
xnor U17948 (N_17948,N_16160,N_16326);
nor U17949 (N_17949,N_16751,N_15763);
nor U17950 (N_17950,N_15924,N_15647);
xnor U17951 (N_17951,N_16427,N_16219);
xnor U17952 (N_17952,N_16782,N_16292);
nand U17953 (N_17953,N_16373,N_16354);
nor U17954 (N_17954,N_16227,N_16528);
xor U17955 (N_17955,N_16165,N_16487);
nand U17956 (N_17956,N_16321,N_15760);
nor U17957 (N_17957,N_16259,N_16129);
or U17958 (N_17958,N_16153,N_15685);
nand U17959 (N_17959,N_16222,N_15731);
xnor U17960 (N_17960,N_16551,N_16051);
xnor U17961 (N_17961,N_15830,N_15669);
or U17962 (N_17962,N_16626,N_15754);
xnor U17963 (N_17963,N_15885,N_16755);
nor U17964 (N_17964,N_16678,N_16662);
nand U17965 (N_17965,N_16634,N_16435);
and U17966 (N_17966,N_15691,N_15995);
or U17967 (N_17967,N_16568,N_16665);
nor U17968 (N_17968,N_15927,N_15690);
nand U17969 (N_17969,N_16239,N_16586);
nand U17970 (N_17970,N_15678,N_16619);
nor U17971 (N_17971,N_16384,N_16058);
nor U17972 (N_17972,N_15748,N_16100);
nand U17973 (N_17973,N_16343,N_16417);
nand U17974 (N_17974,N_16669,N_16139);
nor U17975 (N_17975,N_16155,N_16371);
or U17976 (N_17976,N_16142,N_15957);
and U17977 (N_17977,N_16780,N_16638);
nand U17978 (N_17978,N_16444,N_16718);
or U17979 (N_17979,N_16644,N_16054);
nand U17980 (N_17980,N_15600,N_16707);
and U17981 (N_17981,N_16698,N_16540);
nand U17982 (N_17982,N_16314,N_16158);
nand U17983 (N_17983,N_16489,N_16180);
xor U17984 (N_17984,N_16069,N_16656);
nand U17985 (N_17985,N_16272,N_16688);
and U17986 (N_17986,N_15752,N_16293);
xnor U17987 (N_17987,N_16501,N_16171);
and U17988 (N_17988,N_15602,N_16343);
or U17989 (N_17989,N_16018,N_16275);
or U17990 (N_17990,N_16720,N_15604);
or U17991 (N_17991,N_15983,N_15632);
or U17992 (N_17992,N_16411,N_16741);
nand U17993 (N_17993,N_16194,N_16034);
or U17994 (N_17994,N_16367,N_16027);
nand U17995 (N_17995,N_16086,N_16709);
nand U17996 (N_17996,N_15952,N_16362);
and U17997 (N_17997,N_16657,N_16732);
or U17998 (N_17998,N_16140,N_16352);
nor U17999 (N_17999,N_15759,N_16620);
xor U18000 (N_18000,N_17815,N_17330);
nand U18001 (N_18001,N_17871,N_17604);
and U18002 (N_18002,N_17717,N_17046);
nand U18003 (N_18003,N_17148,N_17327);
and U18004 (N_18004,N_17881,N_17964);
and U18005 (N_18005,N_17137,N_16937);
nor U18006 (N_18006,N_17666,N_17443);
and U18007 (N_18007,N_16967,N_17105);
and U18008 (N_18008,N_17654,N_17566);
nand U18009 (N_18009,N_17447,N_17638);
or U18010 (N_18010,N_17298,N_17322);
nor U18011 (N_18011,N_17492,N_17957);
xor U18012 (N_18012,N_17488,N_17350);
and U18013 (N_18013,N_17089,N_16866);
and U18014 (N_18014,N_17071,N_17238);
and U18015 (N_18015,N_17361,N_17428);
nand U18016 (N_18016,N_17049,N_17683);
nor U18017 (N_18017,N_17213,N_17326);
and U18018 (N_18018,N_17214,N_17934);
or U18019 (N_18019,N_17992,N_17693);
nand U18020 (N_18020,N_17817,N_17570);
xor U18021 (N_18021,N_17739,N_17596);
nand U18022 (N_18022,N_17112,N_17824);
xor U18023 (N_18023,N_17880,N_16806);
and U18024 (N_18024,N_17907,N_17540);
or U18025 (N_18025,N_17651,N_17844);
nor U18026 (N_18026,N_17026,N_17846);
nand U18027 (N_18027,N_16865,N_16813);
and U18028 (N_18028,N_17133,N_16844);
and U18029 (N_18029,N_17920,N_17670);
nor U18030 (N_18030,N_16905,N_17261);
and U18031 (N_18031,N_16921,N_17543);
nor U18032 (N_18032,N_17953,N_17382);
or U18033 (N_18033,N_17775,N_17094);
and U18034 (N_18034,N_17370,N_17098);
and U18035 (N_18035,N_17658,N_17041);
and U18036 (N_18036,N_17211,N_17687);
nor U18037 (N_18037,N_17667,N_17411);
xor U18038 (N_18038,N_17042,N_17988);
xor U18039 (N_18039,N_16944,N_17664);
xor U18040 (N_18040,N_16912,N_17724);
or U18041 (N_18041,N_17710,N_17416);
and U18042 (N_18042,N_17955,N_16919);
and U18043 (N_18043,N_17099,N_17021);
and U18044 (N_18044,N_17414,N_17622);
or U18045 (N_18045,N_16805,N_17561);
nand U18046 (N_18046,N_17475,N_17500);
nor U18047 (N_18047,N_17378,N_17199);
nor U18048 (N_18048,N_17508,N_16933);
nand U18049 (N_18049,N_17158,N_16942);
nor U18050 (N_18050,N_16842,N_17061);
xnor U18051 (N_18051,N_17713,N_17234);
and U18052 (N_18052,N_16927,N_17737);
nor U18053 (N_18053,N_17147,N_17006);
nand U18054 (N_18054,N_17987,N_17360);
and U18055 (N_18055,N_17757,N_17966);
nand U18056 (N_18056,N_16854,N_17497);
and U18057 (N_18057,N_17504,N_16962);
or U18058 (N_18058,N_17828,N_17534);
xnor U18059 (N_18059,N_17085,N_16926);
nand U18060 (N_18060,N_17554,N_16969);
nor U18061 (N_18061,N_17841,N_17547);
nand U18062 (N_18062,N_17176,N_17262);
nand U18063 (N_18063,N_17827,N_17195);
nand U18064 (N_18064,N_17449,N_17362);
xor U18065 (N_18065,N_17458,N_17192);
xnor U18066 (N_18066,N_17559,N_17585);
and U18067 (N_18067,N_16949,N_17059);
nor U18068 (N_18068,N_17791,N_17588);
nor U18069 (N_18069,N_17338,N_16939);
and U18070 (N_18070,N_17927,N_17519);
nand U18071 (N_18071,N_17028,N_17947);
nand U18072 (N_18072,N_17406,N_17183);
nor U18073 (N_18073,N_17936,N_16879);
and U18074 (N_18074,N_17022,N_17044);
xnor U18075 (N_18075,N_17040,N_17560);
nand U18076 (N_18076,N_17229,N_17201);
xor U18077 (N_18077,N_17251,N_17943);
nor U18078 (N_18078,N_17033,N_17720);
nand U18079 (N_18079,N_17535,N_17931);
or U18080 (N_18080,N_17976,N_17851);
xnor U18081 (N_18081,N_17869,N_17445);
nand U18082 (N_18082,N_17744,N_17108);
nor U18083 (N_18083,N_17103,N_17623);
nor U18084 (N_18084,N_17865,N_17132);
and U18085 (N_18085,N_17695,N_17677);
nand U18086 (N_18086,N_17905,N_17563);
nand U18087 (N_18087,N_17075,N_17948);
or U18088 (N_18088,N_17355,N_17233);
nor U18089 (N_18089,N_17823,N_17109);
and U18090 (N_18090,N_17690,N_16841);
nor U18091 (N_18091,N_16907,N_17008);
or U18092 (N_18092,N_17082,N_16849);
and U18093 (N_18093,N_17138,N_17027);
and U18094 (N_18094,N_17276,N_17272);
nor U18095 (N_18095,N_17896,N_17180);
or U18096 (N_18096,N_16913,N_17373);
or U18097 (N_18097,N_17446,N_17968);
nand U18098 (N_18098,N_17128,N_17169);
nor U18099 (N_18099,N_17923,N_17848);
nand U18100 (N_18100,N_16824,N_17241);
xor U18101 (N_18101,N_17538,N_17104);
and U18102 (N_18102,N_17131,N_17727);
xor U18103 (N_18103,N_17043,N_16818);
or U18104 (N_18104,N_17785,N_17808);
nand U18105 (N_18105,N_17198,N_17753);
nor U18106 (N_18106,N_17424,N_17288);
and U18107 (N_18107,N_17281,N_16859);
and U18108 (N_18108,N_17691,N_17462);
nand U18109 (N_18109,N_16995,N_16993);
or U18110 (N_18110,N_17455,N_17155);
or U18111 (N_18111,N_17228,N_17476);
nand U18112 (N_18112,N_16823,N_17478);
xor U18113 (N_18113,N_17834,N_17096);
xor U18114 (N_18114,N_17883,N_17311);
nor U18115 (N_18115,N_17263,N_17888);
xnor U18116 (N_18116,N_17110,N_17982);
or U18117 (N_18117,N_17782,N_17810);
nor U18118 (N_18118,N_16924,N_17002);
and U18119 (N_18119,N_17627,N_17598);
nor U18120 (N_18120,N_17379,N_17423);
nor U18121 (N_18121,N_16888,N_16925);
nor U18122 (N_18122,N_16821,N_17429);
nand U18123 (N_18123,N_17859,N_17226);
and U18124 (N_18124,N_16943,N_17277);
nand U18125 (N_18125,N_17703,N_17221);
nor U18126 (N_18126,N_17750,N_17126);
nor U18127 (N_18127,N_17240,N_17307);
nor U18128 (N_18128,N_17501,N_17742);
nand U18129 (N_18129,N_17235,N_17767);
xor U18130 (N_18130,N_17921,N_17020);
and U18131 (N_18131,N_17090,N_17190);
xor U18132 (N_18132,N_17611,N_17925);
and U18133 (N_18133,N_16965,N_17755);
nand U18134 (N_18134,N_17116,N_17437);
nor U18135 (N_18135,N_17799,N_17393);
xnor U18136 (N_18136,N_17358,N_17084);
xnor U18137 (N_18137,N_17079,N_16994);
nor U18138 (N_18138,N_16941,N_17961);
nand U18139 (N_18139,N_16903,N_17356);
xor U18140 (N_18140,N_17840,N_17838);
or U18141 (N_18141,N_17701,N_17291);
nor U18142 (N_18142,N_17657,N_16974);
or U18143 (N_18143,N_17818,N_17230);
or U18144 (N_18144,N_16809,N_17731);
nor U18145 (N_18145,N_16828,N_17119);
and U18146 (N_18146,N_17625,N_17822);
or U18147 (N_18147,N_17532,N_17659);
xnor U18148 (N_18148,N_17673,N_16838);
xnor U18149 (N_18149,N_17210,N_17018);
or U18150 (N_18150,N_17232,N_17390);
nand U18151 (N_18151,N_17351,N_17702);
or U18152 (N_18152,N_16989,N_17541);
nand U18153 (N_18153,N_16910,N_17552);
and U18154 (N_18154,N_17086,N_16977);
or U18155 (N_18155,N_17980,N_17067);
nand U18156 (N_18156,N_17299,N_17969);
nand U18157 (N_18157,N_17495,N_16826);
and U18158 (N_18158,N_17487,N_17452);
nor U18159 (N_18159,N_17886,N_17152);
and U18160 (N_18160,N_17024,N_17707);
nand U18161 (N_18161,N_17223,N_17107);
and U18162 (N_18162,N_17819,N_17345);
or U18163 (N_18163,N_16884,N_17442);
and U18164 (N_18164,N_17302,N_17854);
nor U18165 (N_18165,N_17906,N_16922);
xor U18166 (N_18166,N_16901,N_17582);
xnor U18167 (N_18167,N_16930,N_17460);
xnor U18168 (N_18168,N_17903,N_17124);
and U18169 (N_18169,N_17680,N_16929);
and U18170 (N_18170,N_17542,N_17178);
and U18171 (N_18171,N_17830,N_17275);
nor U18172 (N_18172,N_17127,N_17990);
nand U18173 (N_18173,N_17050,N_17965);
and U18174 (N_18174,N_17450,N_17062);
and U18175 (N_18175,N_17154,N_17674);
or U18176 (N_18176,N_17315,N_16986);
xnor U18177 (N_18177,N_17397,N_16848);
xor U18178 (N_18178,N_17682,N_16964);
and U18179 (N_18179,N_17718,N_17575);
and U18180 (N_18180,N_17902,N_17811);
xor U18181 (N_18181,N_17522,N_17765);
or U18182 (N_18182,N_16851,N_17974);
nand U18183 (N_18183,N_17016,N_17796);
nor U18184 (N_18184,N_16820,N_16880);
nand U18185 (N_18185,N_16860,N_17072);
nor U18186 (N_18186,N_17877,N_16920);
nor U18187 (N_18187,N_17679,N_17282);
nor U18188 (N_18188,N_17081,N_17493);
and U18189 (N_18189,N_16804,N_17203);
nor U18190 (N_18190,N_16875,N_17245);
nand U18191 (N_18191,N_17309,N_17479);
xnor U18192 (N_18192,N_17465,N_16847);
or U18193 (N_18193,N_17781,N_16947);
or U18194 (N_18194,N_16963,N_17219);
nand U18195 (N_18195,N_17637,N_17312);
nor U18196 (N_18196,N_17448,N_17332);
xnor U18197 (N_18197,N_17646,N_17440);
nand U18198 (N_18198,N_17911,N_17951);
nand U18199 (N_18199,N_16834,N_17320);
xnor U18200 (N_18200,N_17856,N_16990);
nor U18201 (N_18201,N_17857,N_17359);
xnor U18202 (N_18202,N_17185,N_17608);
and U18203 (N_18203,N_17058,N_17209);
xnor U18204 (N_18204,N_17945,N_17369);
and U18205 (N_18205,N_17599,N_17520);
nand U18206 (N_18206,N_17285,N_16890);
xnor U18207 (N_18207,N_17662,N_17463);
or U18208 (N_18208,N_17615,N_16981);
or U18209 (N_18209,N_17162,N_17944);
xnor U18210 (N_18210,N_17655,N_17496);
nand U18211 (N_18211,N_17916,N_17438);
nand U18212 (N_18212,N_17997,N_17172);
and U18213 (N_18213,N_17453,N_17432);
nand U18214 (N_18214,N_17733,N_17716);
or U18215 (N_18215,N_17630,N_17528);
and U18216 (N_18216,N_17803,N_17427);
nor U18217 (N_18217,N_17353,N_17583);
nor U18218 (N_18218,N_17597,N_17308);
or U18219 (N_18219,N_17617,N_17741);
and U18220 (N_18220,N_17885,N_16971);
and U18221 (N_18221,N_17314,N_17486);
and U18222 (N_18222,N_17959,N_16846);
xor U18223 (N_18223,N_17456,N_17760);
xor U18224 (N_18224,N_17417,N_17653);
nor U18225 (N_18225,N_16812,N_17776);
and U18226 (N_18226,N_17053,N_17239);
or U18227 (N_18227,N_17933,N_17783);
nor U18228 (N_18228,N_17420,N_17650);
and U18229 (N_18229,N_17914,N_16999);
nor U18230 (N_18230,N_17052,N_16914);
and U18231 (N_18231,N_17624,N_17193);
nor U18232 (N_18232,N_17231,N_17407);
nor U18233 (N_18233,N_17287,N_17763);
nor U18234 (N_18234,N_17971,N_17200);
or U18235 (N_18235,N_17578,N_17381);
and U18236 (N_18236,N_17498,N_17732);
nand U18237 (N_18237,N_17752,N_17594);
xor U18238 (N_18238,N_16839,N_17484);
and U18239 (N_18239,N_17227,N_17550);
nor U18240 (N_18240,N_17433,N_17114);
nand U18241 (N_18241,N_17507,N_17410);
nor U18242 (N_18242,N_17619,N_16872);
or U18243 (N_18243,N_17122,N_17849);
nor U18244 (N_18244,N_17708,N_17212);
nor U18245 (N_18245,N_17013,N_17768);
and U18246 (N_18246,N_17389,N_17418);
or U18247 (N_18247,N_16951,N_17618);
or U18248 (N_18248,N_17736,N_16959);
xnor U18249 (N_18249,N_17303,N_16807);
nand U18250 (N_18250,N_17402,N_17592);
or U18251 (N_18251,N_16840,N_17893);
xnor U18252 (N_18252,N_17790,N_17884);
nand U18253 (N_18253,N_17807,N_17749);
nand U18254 (N_18254,N_17632,N_17586);
xor U18255 (N_18255,N_17215,N_17347);
and U18256 (N_18256,N_17401,N_17962);
xnor U18257 (N_18257,N_17405,N_17143);
and U18258 (N_18258,N_16992,N_16861);
xor U18259 (N_18259,N_17593,N_17784);
or U18260 (N_18260,N_17474,N_16803);
nand U18261 (N_18261,N_17932,N_17115);
nor U18262 (N_18262,N_17372,N_17343);
xor U18263 (N_18263,N_16952,N_17083);
nand U18264 (N_18264,N_17426,N_17055);
or U18265 (N_18265,N_17093,N_17661);
nor U18266 (N_18266,N_16985,N_17101);
xor U18267 (N_18267,N_17120,N_17340);
nor U18268 (N_18268,N_17709,N_16889);
nand U18269 (N_18269,N_17515,N_17034);
nor U18270 (N_18270,N_17204,N_17259);
or U18271 (N_18271,N_16960,N_16909);
and U18272 (N_18272,N_16957,N_17660);
and U18273 (N_18273,N_17714,N_17000);
xor U18274 (N_18274,N_17584,N_17721);
and U18275 (N_18275,N_17258,N_17635);
nor U18276 (N_18276,N_17477,N_17526);
and U18277 (N_18277,N_17826,N_17007);
nor U18278 (N_18278,N_17640,N_16816);
or U18279 (N_18279,N_17734,N_16893);
or U18280 (N_18280,N_17745,N_17743);
and U18281 (N_18281,N_16867,N_16877);
and U18282 (N_18282,N_17253,N_17140);
nand U18283 (N_18283,N_17786,N_17153);
nand U18284 (N_18284,N_17989,N_16948);
and U18285 (N_18285,N_17206,N_17631);
and U18286 (N_18286,N_16996,N_17789);
nand U18287 (N_18287,N_17573,N_17060);
nor U18288 (N_18288,N_17567,N_16945);
xor U18289 (N_18289,N_17422,N_17861);
xnor U18290 (N_18290,N_17644,N_17950);
or U18291 (N_18291,N_16800,N_17697);
xnor U18292 (N_18292,N_17415,N_17323);
xor U18293 (N_18293,N_16873,N_16853);
xor U18294 (N_18294,N_17265,N_16978);
nor U18295 (N_18295,N_17793,N_17257);
and U18296 (N_18296,N_17876,N_17014);
nand U18297 (N_18297,N_17960,N_17170);
nor U18298 (N_18298,N_17891,N_17915);
or U18299 (N_18299,N_17802,N_17439);
or U18300 (N_18300,N_17904,N_16832);
or U18301 (N_18301,N_17758,N_17409);
or U18302 (N_18302,N_16908,N_17847);
and U18303 (N_18303,N_16954,N_17300);
xnor U18304 (N_18304,N_17145,N_17078);
nand U18305 (N_18305,N_17080,N_16998);
and U18306 (N_18306,N_17357,N_17935);
and U18307 (N_18307,N_17237,N_17688);
nor U18308 (N_18308,N_17333,N_17771);
xor U18309 (N_18309,N_17468,N_17266);
xor U18310 (N_18310,N_16871,N_17978);
nand U18311 (N_18311,N_17529,N_16988);
nand U18312 (N_18312,N_17929,N_17537);
or U18313 (N_18313,N_17816,N_16918);
nor U18314 (N_18314,N_17339,N_17365);
xnor U18315 (N_18315,N_17770,N_17797);
nand U18316 (N_18316,N_17831,N_17324);
and U18317 (N_18317,N_17305,N_17247);
xnor U18318 (N_18318,N_17572,N_17037);
nand U18319 (N_18319,N_17202,N_17384);
or U18320 (N_18320,N_17764,N_17738);
and U18321 (N_18321,N_16883,N_17813);
and U18322 (N_18322,N_17244,N_17289);
xnor U18323 (N_18323,N_17521,N_17530);
nand U18324 (N_18324,N_17348,N_17364);
or U18325 (N_18325,N_17607,N_17250);
and U18326 (N_18326,N_17470,N_17694);
xnor U18327 (N_18327,N_17994,N_17336);
nor U18328 (N_18328,N_16991,N_17242);
nor U18329 (N_18329,N_17825,N_16886);
nor U18330 (N_18330,N_16982,N_17301);
xnor U18331 (N_18331,N_17161,N_17341);
or U18332 (N_18332,N_17391,N_17868);
or U18333 (N_18333,N_17236,N_17380);
or U18334 (N_18334,N_17867,N_17175);
nand U18335 (N_18335,N_17606,N_16936);
and U18336 (N_18336,N_17792,N_17678);
or U18337 (N_18337,N_17441,N_17246);
or U18338 (N_18338,N_17489,N_17171);
nor U18339 (N_18339,N_17207,N_16980);
xor U18340 (N_18340,N_16825,N_16900);
and U18341 (N_18341,N_17248,N_17769);
nand U18342 (N_18342,N_16902,N_17224);
xor U18343 (N_18343,N_17574,N_16881);
nor U18344 (N_18344,N_17118,N_17385);
nor U18345 (N_18345,N_17523,N_17981);
and U18346 (N_18346,N_17562,N_16808);
nand U18347 (N_18347,N_16894,N_17820);
nor U18348 (N_18348,N_17954,N_17001);
or U18349 (N_18349,N_17106,N_17938);
or U18350 (N_18350,N_17074,N_17472);
nand U18351 (N_18351,N_17064,N_17620);
or U18352 (N_18352,N_16968,N_17012);
xor U18353 (N_18353,N_17457,N_17100);
nand U18354 (N_18354,N_16931,N_17882);
nand U18355 (N_18355,N_17996,N_16869);
xnor U18356 (N_18356,N_17806,N_17063);
nand U18357 (N_18357,N_17481,N_17613);
or U18358 (N_18358,N_16946,N_17590);
or U18359 (N_18359,N_16895,N_17983);
nand U18360 (N_18360,N_17863,N_17387);
nor U18361 (N_18361,N_17647,N_17220);
and U18362 (N_18362,N_17832,N_16885);
and U18363 (N_18363,N_17068,N_17600);
or U18364 (N_18364,N_17003,N_16897);
and U18365 (N_18365,N_17912,N_17698);
xor U18366 (N_18366,N_17436,N_17511);
nor U18367 (N_18367,N_17696,N_17998);
nor U18368 (N_18368,N_17165,N_17243);
nand U18369 (N_18369,N_17366,N_17991);
nand U18370 (N_18370,N_17149,N_16802);
nand U18371 (N_18371,N_17761,N_16997);
nor U18372 (N_18372,N_17711,N_17225);
nand U18373 (N_18373,N_17910,N_17167);
and U18374 (N_18374,N_16857,N_17367);
and U18375 (N_18375,N_17480,N_17181);
or U18376 (N_18376,N_17917,N_17940);
and U18377 (N_18377,N_17264,N_17306);
nor U18378 (N_18378,N_17591,N_17310);
and U18379 (N_18379,N_17352,N_17568);
nor U18380 (N_18380,N_17870,N_16958);
nand U18381 (N_18381,N_17860,N_17643);
or U18382 (N_18382,N_17371,N_17787);
nand U18383 (N_18383,N_16836,N_17928);
nand U18384 (N_18384,N_17374,N_17451);
or U18385 (N_18385,N_16915,N_17151);
xnor U18386 (N_18386,N_17842,N_17286);
and U18387 (N_18387,N_17553,N_17772);
nor U18388 (N_18388,N_17942,N_16882);
nor U18389 (N_18389,N_17054,N_17853);
xor U18390 (N_18390,N_17166,N_17656);
and U18391 (N_18391,N_17836,N_17609);
nor U18392 (N_18392,N_16970,N_17156);
and U18393 (N_18393,N_17773,N_17524);
or U18394 (N_18394,N_17835,N_16856);
xor U18395 (N_18395,N_16917,N_17396);
or U18396 (N_18396,N_17270,N_17412);
and U18397 (N_18397,N_16837,N_17924);
xor U18398 (N_18398,N_17454,N_16850);
nand U18399 (N_18399,N_17077,N_17399);
xor U18400 (N_18400,N_17821,N_17862);
and U18401 (N_18401,N_17179,N_16911);
or U18402 (N_18402,N_17461,N_17756);
nor U18403 (N_18403,N_17469,N_17531);
nor U18404 (N_18404,N_17913,N_17939);
nor U18405 (N_18405,N_17892,N_17070);
xor U18406 (N_18406,N_17873,N_17605);
nand U18407 (N_18407,N_17164,N_17814);
nor U18408 (N_18408,N_17400,N_17864);
xor U18409 (N_18409,N_17648,N_17459);
or U18410 (N_18410,N_17740,N_16983);
nand U18411 (N_18411,N_17845,N_17073);
and U18412 (N_18412,N_17895,N_17325);
and U18413 (N_18413,N_17548,N_16972);
xnor U18414 (N_18414,N_17284,N_17377);
or U18415 (N_18415,N_17901,N_17509);
nand U18416 (N_18416,N_17502,N_17675);
and U18417 (N_18417,N_17774,N_16928);
nand U18418 (N_18418,N_17930,N_17900);
nor U18419 (N_18419,N_17681,N_17706);
nand U18420 (N_18420,N_17194,N_17386);
nor U18421 (N_18421,N_17395,N_17260);
nand U18422 (N_18422,N_16835,N_16938);
xor U18423 (N_18423,N_16863,N_17017);
nand U18424 (N_18424,N_17805,N_17545);
nor U18425 (N_18425,N_17273,N_16950);
or U18426 (N_18426,N_17977,N_16934);
or U18427 (N_18427,N_17595,N_17267);
and U18428 (N_18428,N_17919,N_17986);
xor U18429 (N_18429,N_17189,N_17722);
nor U18430 (N_18430,N_17795,N_17875);
nor U18431 (N_18431,N_17649,N_17283);
xnor U18432 (N_18432,N_17095,N_17196);
nor U18433 (N_18433,N_17011,N_17217);
xor U18434 (N_18434,N_17612,N_17676);
and U18435 (N_18435,N_17467,N_17536);
xor U18436 (N_18436,N_17546,N_17191);
nand U18437 (N_18437,N_16898,N_17091);
nand U18438 (N_18438,N_17464,N_17652);
nand U18439 (N_18439,N_17730,N_17759);
or U18440 (N_18440,N_17280,N_17829);
and U18441 (N_18441,N_16896,N_17269);
nor U18442 (N_18442,N_17689,N_17004);
xnor U18443 (N_18443,N_17316,N_17328);
nand U18444 (N_18444,N_16932,N_17946);
xnor U18445 (N_18445,N_17958,N_17576);
or U18446 (N_18446,N_17254,N_17321);
and U18447 (N_18447,N_17967,N_16973);
or U18448 (N_18448,N_17421,N_17146);
xor U18449 (N_18449,N_17368,N_17894);
nand U18450 (N_18450,N_17066,N_17641);
or U18451 (N_18451,N_17728,N_17130);
xnor U18452 (N_18452,N_17136,N_17296);
xnor U18453 (N_18453,N_16979,N_16801);
or U18454 (N_18454,N_17304,N_17705);
xor U18455 (N_18455,N_16976,N_17601);
and U18456 (N_18456,N_17956,N_16955);
or U18457 (N_18457,N_17473,N_17610);
xor U18458 (N_18458,N_17937,N_17047);
xor U18459 (N_18459,N_17111,N_17471);
or U18460 (N_18460,N_17636,N_16868);
xnor U18461 (N_18461,N_17375,N_17342);
nor U18462 (N_18462,N_17491,N_17890);
nor U18463 (N_18463,N_17581,N_17252);
and U18464 (N_18464,N_17317,N_17051);
or U18465 (N_18465,N_17163,N_16940);
nand U18466 (N_18466,N_17329,N_16858);
nand U18467 (N_18467,N_17123,N_17056);
nor U18468 (N_18468,N_17569,N_17483);
xnor U18469 (N_18469,N_17088,N_17278);
nor U18470 (N_18470,N_17952,N_17376);
nand U18471 (N_18471,N_16887,N_16819);
nand U18472 (N_18472,N_17218,N_17125);
xnor U18473 (N_18473,N_17866,N_17404);
nand U18474 (N_18474,N_17941,N_16984);
or U18475 (N_18475,N_17999,N_17392);
nor U18476 (N_18476,N_17850,N_17626);
nor U18477 (N_18477,N_17922,N_17413);
or U18478 (N_18478,N_17889,N_17346);
nand U18479 (N_18479,N_17801,N_17113);
and U18480 (N_18480,N_16811,N_17160);
nor U18481 (N_18481,N_17057,N_17879);
nand U18482 (N_18482,N_17249,N_16833);
xnor U18483 (N_18483,N_17735,N_17293);
or U18484 (N_18484,N_17949,N_17794);
nor U18485 (N_18485,N_16899,N_17579);
nand U18486 (N_18486,N_17510,N_17926);
nor U18487 (N_18487,N_17274,N_17533);
nor U18488 (N_18488,N_16874,N_16961);
and U18489 (N_18489,N_17777,N_17494);
nand U18490 (N_18490,N_17580,N_17645);
nand U18491 (N_18491,N_16814,N_17255);
xnor U18492 (N_18492,N_17430,N_17015);
nor U18493 (N_18493,N_17045,N_17036);
nor U18494 (N_18494,N_17517,N_17556);
xnor U18495 (N_18495,N_16870,N_17855);
and U18496 (N_18496,N_17294,N_17642);
or U18497 (N_18497,N_17684,N_17295);
xnor U18498 (N_18498,N_16852,N_16953);
xor U18499 (N_18499,N_17503,N_17010);
or U18500 (N_18500,N_16829,N_17506);
nand U18501 (N_18501,N_17256,N_16935);
or U18502 (N_18502,N_17798,N_17577);
nand U18503 (N_18503,N_17672,N_17751);
xnor U18504 (N_18504,N_17686,N_17539);
xnor U18505 (N_18505,N_17628,N_17704);
nand U18506 (N_18506,N_17555,N_17023);
nor U18507 (N_18507,N_17973,N_17979);
or U18508 (N_18508,N_17425,N_17669);
nor U18509 (N_18509,N_17897,N_17383);
and U18510 (N_18510,N_16966,N_16916);
xor U18511 (N_18511,N_17766,N_17319);
xnor U18512 (N_18512,N_17208,N_16822);
nor U18513 (N_18513,N_17268,N_17725);
and U18514 (N_18514,N_17908,N_17833);
and U18515 (N_18515,N_17513,N_17134);
nand U18516 (N_18516,N_16864,N_17009);
xor U18517 (N_18517,N_17839,N_17184);
and U18518 (N_18518,N_17565,N_17621);
nand U18519 (N_18519,N_17715,N_17729);
nor U18520 (N_18520,N_17723,N_17334);
and U18521 (N_18521,N_17544,N_17097);
and U18522 (N_18522,N_17514,N_17159);
or U18523 (N_18523,N_17019,N_17102);
nor U18524 (N_18524,N_17435,N_17800);
nor U18525 (N_18525,N_17963,N_17144);
nand U18526 (N_18526,N_17038,N_17685);
and U18527 (N_18527,N_17878,N_17852);
or U18528 (N_18528,N_16862,N_17292);
nand U18529 (N_18529,N_17177,N_17671);
nor U18530 (N_18530,N_17571,N_16810);
nor U18531 (N_18531,N_17335,N_17076);
xnor U18532 (N_18532,N_17918,N_17505);
and U18533 (N_18533,N_16831,N_17564);
and U18534 (N_18534,N_17388,N_17394);
nand U18535 (N_18535,N_17985,N_17482);
nand U18536 (N_18536,N_17187,N_17129);
nor U18537 (N_18537,N_17290,N_17031);
and U18538 (N_18538,N_17762,N_17135);
or U18539 (N_18539,N_17874,N_16904);
nand U18540 (N_18540,N_17812,N_17150);
nor U18541 (N_18541,N_17837,N_17168);
xnor U18542 (N_18542,N_17972,N_17712);
nor U18543 (N_18543,N_17551,N_17216);
xnor U18544 (N_18544,N_16830,N_17444);
and U18545 (N_18545,N_16878,N_17271);
xnor U18546 (N_18546,N_17747,N_17898);
xnor U18547 (N_18547,N_17634,N_17331);
or U18548 (N_18548,N_17726,N_17403);
xnor U18549 (N_18549,N_16855,N_17665);
nor U18550 (N_18550,N_16817,N_17512);
and U18551 (N_18551,N_16843,N_17039);
xor U18552 (N_18552,N_16923,N_17297);
nand U18553 (N_18553,N_17408,N_17318);
xor U18554 (N_18554,N_17668,N_17746);
xnor U18555 (N_18555,N_17490,N_16906);
nand U18556 (N_18556,N_17975,N_16891);
xor U18557 (N_18557,N_17065,N_17970);
xnor U18558 (N_18558,N_17466,N_17349);
and U18559 (N_18559,N_17629,N_17363);
nor U18560 (N_18560,N_16892,N_17780);
or U18561 (N_18561,N_17700,N_17692);
nor U18562 (N_18562,N_17434,N_17899);
nand U18563 (N_18563,N_17779,N_17035);
or U18564 (N_18564,N_17663,N_17558);
nor U18565 (N_18565,N_17398,N_17344);
nand U18566 (N_18566,N_17633,N_17337);
nand U18567 (N_18567,N_17748,N_17516);
nand U18568 (N_18568,N_17030,N_17499);
and U18569 (N_18569,N_17182,N_17843);
and U18570 (N_18570,N_17222,N_17174);
and U18571 (N_18571,N_17205,N_16827);
or U18572 (N_18572,N_17887,N_17186);
and U18573 (N_18573,N_17788,N_17616);
and U18574 (N_18574,N_17197,N_17029);
nand U18575 (N_18575,N_17141,N_17142);
xor U18576 (N_18576,N_17005,N_17639);
xor U18577 (N_18577,N_17354,N_17092);
or U18578 (N_18578,N_17872,N_17557);
or U18579 (N_18579,N_17419,N_17139);
xnor U18580 (N_18580,N_17527,N_17909);
xnor U18581 (N_18581,N_17069,N_16987);
nor U18582 (N_18582,N_17485,N_16956);
nor U18583 (N_18583,N_16876,N_17313);
or U18584 (N_18584,N_17525,N_17032);
and U18585 (N_18585,N_16975,N_17699);
or U18586 (N_18586,N_17431,N_17602);
or U18587 (N_18587,N_17173,N_16845);
nor U18588 (N_18588,N_17809,N_17188);
or U18589 (N_18589,N_17993,N_17719);
and U18590 (N_18590,N_17754,N_17279);
nand U18591 (N_18591,N_17121,N_17858);
or U18592 (N_18592,N_17157,N_17804);
nand U18593 (N_18593,N_17995,N_17117);
nand U18594 (N_18594,N_17778,N_16815);
and U18595 (N_18595,N_17614,N_17518);
xor U18596 (N_18596,N_17587,N_17984);
or U18597 (N_18597,N_17048,N_17025);
xor U18598 (N_18598,N_17549,N_17589);
and U18599 (N_18599,N_17603,N_17087);
or U18600 (N_18600,N_16982,N_17260);
nand U18601 (N_18601,N_17410,N_17906);
and U18602 (N_18602,N_17938,N_16846);
or U18603 (N_18603,N_17063,N_17389);
nand U18604 (N_18604,N_17323,N_16969);
or U18605 (N_18605,N_17049,N_17822);
or U18606 (N_18606,N_17995,N_17008);
nand U18607 (N_18607,N_17526,N_17695);
nor U18608 (N_18608,N_17059,N_17702);
and U18609 (N_18609,N_17629,N_17112);
nand U18610 (N_18610,N_17771,N_17302);
nand U18611 (N_18611,N_17584,N_16941);
nor U18612 (N_18612,N_17425,N_17127);
and U18613 (N_18613,N_17384,N_17367);
nand U18614 (N_18614,N_17519,N_17507);
or U18615 (N_18615,N_17789,N_17670);
and U18616 (N_18616,N_17980,N_17042);
nor U18617 (N_18617,N_17390,N_17342);
or U18618 (N_18618,N_17789,N_17401);
nand U18619 (N_18619,N_17296,N_17168);
nor U18620 (N_18620,N_17939,N_17972);
or U18621 (N_18621,N_17725,N_16853);
nand U18622 (N_18622,N_17026,N_17593);
nand U18623 (N_18623,N_17862,N_17647);
nand U18624 (N_18624,N_17038,N_17673);
xor U18625 (N_18625,N_17666,N_16825);
or U18626 (N_18626,N_17500,N_17311);
xnor U18627 (N_18627,N_17217,N_17224);
or U18628 (N_18628,N_17859,N_17800);
nand U18629 (N_18629,N_17817,N_17632);
xor U18630 (N_18630,N_17955,N_17373);
or U18631 (N_18631,N_16961,N_17272);
and U18632 (N_18632,N_17016,N_17094);
nor U18633 (N_18633,N_16908,N_17744);
or U18634 (N_18634,N_17997,N_16908);
nand U18635 (N_18635,N_17923,N_17484);
xnor U18636 (N_18636,N_17070,N_17019);
nand U18637 (N_18637,N_17151,N_17203);
or U18638 (N_18638,N_17292,N_17919);
and U18639 (N_18639,N_17620,N_17165);
or U18640 (N_18640,N_17140,N_17921);
nand U18641 (N_18641,N_17251,N_17989);
nor U18642 (N_18642,N_17645,N_17848);
xnor U18643 (N_18643,N_17659,N_17357);
and U18644 (N_18644,N_17031,N_17830);
or U18645 (N_18645,N_17384,N_17571);
or U18646 (N_18646,N_17267,N_16870);
and U18647 (N_18647,N_17661,N_17331);
or U18648 (N_18648,N_17363,N_17679);
nor U18649 (N_18649,N_17038,N_17483);
xnor U18650 (N_18650,N_17129,N_17584);
or U18651 (N_18651,N_16812,N_17752);
xor U18652 (N_18652,N_16956,N_17469);
nor U18653 (N_18653,N_17085,N_17580);
nand U18654 (N_18654,N_17390,N_17393);
xnor U18655 (N_18655,N_16886,N_16983);
nor U18656 (N_18656,N_16916,N_17303);
nand U18657 (N_18657,N_17926,N_17102);
xnor U18658 (N_18658,N_17660,N_17316);
xor U18659 (N_18659,N_17825,N_17239);
or U18660 (N_18660,N_17506,N_16903);
and U18661 (N_18661,N_17288,N_17192);
nor U18662 (N_18662,N_17869,N_16923);
nor U18663 (N_18663,N_17014,N_16859);
and U18664 (N_18664,N_17675,N_17109);
nor U18665 (N_18665,N_17612,N_17137);
or U18666 (N_18666,N_17227,N_16837);
and U18667 (N_18667,N_17606,N_17743);
or U18668 (N_18668,N_17287,N_17284);
or U18669 (N_18669,N_16875,N_17319);
or U18670 (N_18670,N_17042,N_17690);
or U18671 (N_18671,N_17723,N_17252);
nand U18672 (N_18672,N_17034,N_17198);
nand U18673 (N_18673,N_17033,N_17706);
or U18674 (N_18674,N_17464,N_17968);
and U18675 (N_18675,N_17651,N_16987);
or U18676 (N_18676,N_17121,N_17156);
and U18677 (N_18677,N_17979,N_17116);
xnor U18678 (N_18678,N_17425,N_16936);
nor U18679 (N_18679,N_17956,N_17799);
and U18680 (N_18680,N_17967,N_17136);
nor U18681 (N_18681,N_17496,N_16865);
xor U18682 (N_18682,N_17950,N_17084);
nand U18683 (N_18683,N_17072,N_17553);
or U18684 (N_18684,N_17695,N_17799);
and U18685 (N_18685,N_17309,N_17313);
or U18686 (N_18686,N_17489,N_17004);
nor U18687 (N_18687,N_17392,N_17099);
nand U18688 (N_18688,N_17629,N_17119);
nor U18689 (N_18689,N_17888,N_17476);
or U18690 (N_18690,N_17140,N_17245);
nand U18691 (N_18691,N_17795,N_17580);
xnor U18692 (N_18692,N_17156,N_17095);
and U18693 (N_18693,N_16856,N_17884);
and U18694 (N_18694,N_17686,N_17568);
or U18695 (N_18695,N_17947,N_17380);
or U18696 (N_18696,N_17576,N_17361);
xor U18697 (N_18697,N_17390,N_17150);
nor U18698 (N_18698,N_16965,N_17934);
and U18699 (N_18699,N_17203,N_17638);
and U18700 (N_18700,N_17040,N_17666);
and U18701 (N_18701,N_17619,N_16861);
xnor U18702 (N_18702,N_17907,N_17567);
or U18703 (N_18703,N_16834,N_17625);
xor U18704 (N_18704,N_17324,N_17077);
nand U18705 (N_18705,N_17746,N_17497);
or U18706 (N_18706,N_17322,N_17853);
nor U18707 (N_18707,N_16863,N_17115);
xor U18708 (N_18708,N_17280,N_17432);
and U18709 (N_18709,N_17870,N_17496);
xor U18710 (N_18710,N_17857,N_17221);
or U18711 (N_18711,N_16948,N_17649);
and U18712 (N_18712,N_17823,N_17148);
or U18713 (N_18713,N_16861,N_17691);
xor U18714 (N_18714,N_17135,N_17168);
nor U18715 (N_18715,N_17475,N_17828);
or U18716 (N_18716,N_17405,N_17428);
nor U18717 (N_18717,N_17005,N_17089);
nor U18718 (N_18718,N_17884,N_17379);
xor U18719 (N_18719,N_17181,N_17749);
and U18720 (N_18720,N_17189,N_17107);
and U18721 (N_18721,N_17383,N_17733);
and U18722 (N_18722,N_16893,N_17394);
and U18723 (N_18723,N_16996,N_17919);
xor U18724 (N_18724,N_17845,N_17436);
xor U18725 (N_18725,N_16810,N_17489);
or U18726 (N_18726,N_17688,N_17755);
nor U18727 (N_18727,N_17582,N_17576);
or U18728 (N_18728,N_17683,N_17094);
nor U18729 (N_18729,N_16952,N_17002);
nand U18730 (N_18730,N_17320,N_17616);
nor U18731 (N_18731,N_17530,N_16821);
or U18732 (N_18732,N_17248,N_17505);
nand U18733 (N_18733,N_16827,N_17218);
and U18734 (N_18734,N_17136,N_17215);
nand U18735 (N_18735,N_17508,N_16827);
nor U18736 (N_18736,N_16926,N_17885);
and U18737 (N_18737,N_17951,N_17807);
or U18738 (N_18738,N_16872,N_17926);
nand U18739 (N_18739,N_17451,N_17643);
or U18740 (N_18740,N_17124,N_17934);
or U18741 (N_18741,N_16820,N_17237);
nor U18742 (N_18742,N_17882,N_17879);
or U18743 (N_18743,N_16882,N_17626);
nand U18744 (N_18744,N_17387,N_17858);
xnor U18745 (N_18745,N_17332,N_16837);
nor U18746 (N_18746,N_17601,N_17196);
and U18747 (N_18747,N_17237,N_17010);
or U18748 (N_18748,N_17342,N_17045);
and U18749 (N_18749,N_17207,N_17877);
nor U18750 (N_18750,N_17165,N_17994);
nor U18751 (N_18751,N_17404,N_17723);
and U18752 (N_18752,N_17416,N_17716);
or U18753 (N_18753,N_17126,N_17738);
nor U18754 (N_18754,N_16971,N_16840);
nor U18755 (N_18755,N_17891,N_16820);
nand U18756 (N_18756,N_17042,N_17864);
nor U18757 (N_18757,N_17670,N_16902);
and U18758 (N_18758,N_17728,N_17436);
and U18759 (N_18759,N_17823,N_17665);
nor U18760 (N_18760,N_17565,N_17461);
and U18761 (N_18761,N_16868,N_16930);
and U18762 (N_18762,N_17338,N_16865);
or U18763 (N_18763,N_16886,N_17998);
or U18764 (N_18764,N_17290,N_17333);
nand U18765 (N_18765,N_17917,N_17137);
xnor U18766 (N_18766,N_17863,N_17413);
and U18767 (N_18767,N_17387,N_16856);
nand U18768 (N_18768,N_17874,N_17043);
nand U18769 (N_18769,N_16870,N_17345);
nand U18770 (N_18770,N_17178,N_17158);
and U18771 (N_18771,N_17945,N_17327);
nor U18772 (N_18772,N_17480,N_17464);
nand U18773 (N_18773,N_17101,N_16854);
nor U18774 (N_18774,N_16915,N_16930);
and U18775 (N_18775,N_17090,N_17136);
nand U18776 (N_18776,N_17489,N_17583);
xnor U18777 (N_18777,N_17717,N_17517);
nor U18778 (N_18778,N_17181,N_17192);
or U18779 (N_18779,N_16967,N_16913);
and U18780 (N_18780,N_17461,N_17274);
nand U18781 (N_18781,N_17609,N_17201);
nand U18782 (N_18782,N_17714,N_17583);
nor U18783 (N_18783,N_17732,N_17537);
nand U18784 (N_18784,N_17910,N_17925);
and U18785 (N_18785,N_17491,N_17000);
or U18786 (N_18786,N_17532,N_17649);
nor U18787 (N_18787,N_17148,N_17149);
nor U18788 (N_18788,N_17392,N_17762);
nor U18789 (N_18789,N_17901,N_17218);
or U18790 (N_18790,N_17629,N_17517);
and U18791 (N_18791,N_17941,N_17651);
nor U18792 (N_18792,N_16867,N_17283);
and U18793 (N_18793,N_17645,N_16872);
and U18794 (N_18794,N_16951,N_17729);
nand U18795 (N_18795,N_17641,N_17859);
nor U18796 (N_18796,N_17631,N_16954);
and U18797 (N_18797,N_17260,N_17815);
and U18798 (N_18798,N_16898,N_17054);
nand U18799 (N_18799,N_17726,N_17173);
xnor U18800 (N_18800,N_17924,N_17820);
or U18801 (N_18801,N_16988,N_16918);
nand U18802 (N_18802,N_17789,N_17057);
or U18803 (N_18803,N_16925,N_17473);
nor U18804 (N_18804,N_17220,N_17087);
nand U18805 (N_18805,N_17905,N_17191);
nand U18806 (N_18806,N_17626,N_17058);
and U18807 (N_18807,N_16993,N_17227);
and U18808 (N_18808,N_17776,N_17573);
xnor U18809 (N_18809,N_17851,N_17932);
nor U18810 (N_18810,N_17877,N_17121);
or U18811 (N_18811,N_16964,N_16973);
nand U18812 (N_18812,N_17250,N_17372);
nand U18813 (N_18813,N_16900,N_17858);
and U18814 (N_18814,N_17893,N_17822);
or U18815 (N_18815,N_17641,N_17579);
nor U18816 (N_18816,N_17135,N_17177);
or U18817 (N_18817,N_17173,N_17425);
xnor U18818 (N_18818,N_16895,N_17939);
xor U18819 (N_18819,N_17248,N_17951);
and U18820 (N_18820,N_17315,N_17092);
or U18821 (N_18821,N_17651,N_17174);
or U18822 (N_18822,N_17187,N_17625);
xor U18823 (N_18823,N_17292,N_17869);
xor U18824 (N_18824,N_17771,N_17915);
and U18825 (N_18825,N_17824,N_17267);
nand U18826 (N_18826,N_16871,N_17475);
xor U18827 (N_18827,N_17175,N_17733);
and U18828 (N_18828,N_17902,N_17340);
xor U18829 (N_18829,N_17861,N_17588);
nand U18830 (N_18830,N_17335,N_17260);
and U18831 (N_18831,N_17196,N_17703);
and U18832 (N_18832,N_17721,N_17670);
nor U18833 (N_18833,N_16889,N_17348);
and U18834 (N_18834,N_17956,N_17252);
xor U18835 (N_18835,N_17866,N_17757);
xnor U18836 (N_18836,N_17973,N_17123);
xor U18837 (N_18837,N_17285,N_17274);
nand U18838 (N_18838,N_17716,N_17661);
nand U18839 (N_18839,N_17699,N_16970);
xnor U18840 (N_18840,N_17507,N_17822);
nor U18841 (N_18841,N_17693,N_17501);
or U18842 (N_18842,N_17409,N_17248);
or U18843 (N_18843,N_17277,N_17156);
xnor U18844 (N_18844,N_17936,N_16957);
and U18845 (N_18845,N_17305,N_17384);
nand U18846 (N_18846,N_17993,N_16951);
nor U18847 (N_18847,N_16904,N_16943);
nand U18848 (N_18848,N_16830,N_17333);
nor U18849 (N_18849,N_17111,N_17604);
xnor U18850 (N_18850,N_17343,N_17921);
nor U18851 (N_18851,N_16899,N_17298);
nor U18852 (N_18852,N_17874,N_17362);
nand U18853 (N_18853,N_17591,N_16859);
nand U18854 (N_18854,N_16992,N_17092);
or U18855 (N_18855,N_17188,N_17488);
xnor U18856 (N_18856,N_17565,N_17762);
xnor U18857 (N_18857,N_17648,N_17546);
nand U18858 (N_18858,N_17449,N_17813);
nand U18859 (N_18859,N_17977,N_17346);
and U18860 (N_18860,N_17788,N_17921);
nand U18861 (N_18861,N_17545,N_17218);
or U18862 (N_18862,N_17896,N_16924);
nand U18863 (N_18863,N_16841,N_17393);
xor U18864 (N_18864,N_17041,N_17722);
xor U18865 (N_18865,N_17253,N_17748);
nand U18866 (N_18866,N_17360,N_17124);
and U18867 (N_18867,N_17135,N_17914);
or U18868 (N_18868,N_17040,N_17527);
nand U18869 (N_18869,N_17819,N_17513);
or U18870 (N_18870,N_17549,N_17136);
nor U18871 (N_18871,N_17411,N_17809);
or U18872 (N_18872,N_17707,N_17339);
xnor U18873 (N_18873,N_17244,N_17834);
xnor U18874 (N_18874,N_17888,N_17241);
or U18875 (N_18875,N_16841,N_17252);
and U18876 (N_18876,N_17967,N_17720);
nand U18877 (N_18877,N_17464,N_17179);
xnor U18878 (N_18878,N_17046,N_17199);
xnor U18879 (N_18879,N_17978,N_17804);
xor U18880 (N_18880,N_17704,N_17436);
nand U18881 (N_18881,N_17497,N_17823);
and U18882 (N_18882,N_17907,N_17372);
xor U18883 (N_18883,N_17380,N_17848);
and U18884 (N_18884,N_17983,N_16880);
and U18885 (N_18885,N_16922,N_17650);
or U18886 (N_18886,N_17867,N_17797);
nor U18887 (N_18887,N_17433,N_17421);
and U18888 (N_18888,N_17317,N_17895);
or U18889 (N_18889,N_17489,N_17518);
nand U18890 (N_18890,N_17840,N_16952);
nor U18891 (N_18891,N_16907,N_17659);
nand U18892 (N_18892,N_16986,N_17248);
nand U18893 (N_18893,N_17487,N_17195);
nor U18894 (N_18894,N_16908,N_16831);
or U18895 (N_18895,N_17299,N_17882);
or U18896 (N_18896,N_17708,N_17654);
and U18897 (N_18897,N_17050,N_17163);
nor U18898 (N_18898,N_16971,N_17474);
nor U18899 (N_18899,N_17819,N_17024);
or U18900 (N_18900,N_17319,N_17208);
nor U18901 (N_18901,N_17003,N_17125);
and U18902 (N_18902,N_16921,N_17391);
nor U18903 (N_18903,N_17662,N_17159);
nand U18904 (N_18904,N_17686,N_17336);
or U18905 (N_18905,N_17028,N_17737);
nor U18906 (N_18906,N_17438,N_17346);
xor U18907 (N_18907,N_17445,N_17811);
or U18908 (N_18908,N_17391,N_17770);
nand U18909 (N_18909,N_17592,N_17971);
or U18910 (N_18910,N_17281,N_17259);
or U18911 (N_18911,N_17906,N_17338);
nor U18912 (N_18912,N_17899,N_17223);
nor U18913 (N_18913,N_17481,N_16870);
nand U18914 (N_18914,N_17564,N_17283);
xnor U18915 (N_18915,N_17795,N_16880);
nor U18916 (N_18916,N_17274,N_17453);
or U18917 (N_18917,N_17463,N_16882);
xor U18918 (N_18918,N_17447,N_16830);
xnor U18919 (N_18919,N_17142,N_17602);
nor U18920 (N_18920,N_16886,N_17669);
nor U18921 (N_18921,N_17248,N_17184);
nor U18922 (N_18922,N_16948,N_17534);
or U18923 (N_18923,N_17846,N_17449);
and U18924 (N_18924,N_17012,N_17912);
nor U18925 (N_18925,N_17377,N_17174);
or U18926 (N_18926,N_17865,N_17102);
or U18927 (N_18927,N_16847,N_17439);
xor U18928 (N_18928,N_17312,N_17624);
or U18929 (N_18929,N_17580,N_16938);
and U18930 (N_18930,N_17462,N_17851);
or U18931 (N_18931,N_16911,N_17209);
nor U18932 (N_18932,N_17290,N_17292);
nand U18933 (N_18933,N_17350,N_17352);
nor U18934 (N_18934,N_17527,N_17315);
and U18935 (N_18935,N_17083,N_16865);
xor U18936 (N_18936,N_17297,N_17967);
xor U18937 (N_18937,N_16954,N_16861);
xnor U18938 (N_18938,N_17091,N_16977);
xor U18939 (N_18939,N_17410,N_17002);
xor U18940 (N_18940,N_17211,N_17239);
and U18941 (N_18941,N_17069,N_17202);
xnor U18942 (N_18942,N_17361,N_17022);
or U18943 (N_18943,N_17434,N_17797);
nand U18944 (N_18944,N_17623,N_17209);
or U18945 (N_18945,N_16983,N_16961);
and U18946 (N_18946,N_17790,N_17308);
nor U18947 (N_18947,N_17655,N_17632);
or U18948 (N_18948,N_17583,N_17628);
xnor U18949 (N_18949,N_17139,N_17072);
and U18950 (N_18950,N_17935,N_17277);
nor U18951 (N_18951,N_17813,N_16872);
xor U18952 (N_18952,N_17282,N_17673);
nand U18953 (N_18953,N_17790,N_17727);
nand U18954 (N_18954,N_17889,N_17922);
and U18955 (N_18955,N_17098,N_17182);
and U18956 (N_18956,N_16884,N_17553);
nand U18957 (N_18957,N_16895,N_17514);
nor U18958 (N_18958,N_17283,N_17478);
nand U18959 (N_18959,N_17462,N_17701);
nand U18960 (N_18960,N_17898,N_17529);
and U18961 (N_18961,N_17359,N_16819);
or U18962 (N_18962,N_17490,N_16910);
xor U18963 (N_18963,N_17288,N_17246);
nor U18964 (N_18964,N_16992,N_16909);
nor U18965 (N_18965,N_17175,N_17240);
xnor U18966 (N_18966,N_17356,N_17404);
and U18967 (N_18967,N_17987,N_17283);
xor U18968 (N_18968,N_17480,N_17023);
nor U18969 (N_18969,N_17933,N_17761);
nor U18970 (N_18970,N_17182,N_17109);
or U18971 (N_18971,N_17257,N_17445);
or U18972 (N_18972,N_17196,N_17110);
nand U18973 (N_18973,N_17336,N_17912);
or U18974 (N_18974,N_17599,N_16808);
nor U18975 (N_18975,N_17292,N_17539);
and U18976 (N_18976,N_17940,N_16933);
xor U18977 (N_18977,N_17369,N_16937);
xor U18978 (N_18978,N_17621,N_17460);
or U18979 (N_18979,N_17414,N_17278);
nand U18980 (N_18980,N_17369,N_17315);
nand U18981 (N_18981,N_17653,N_17309);
nand U18982 (N_18982,N_16993,N_17528);
nor U18983 (N_18983,N_17273,N_17185);
and U18984 (N_18984,N_16999,N_17727);
and U18985 (N_18985,N_17345,N_16932);
nand U18986 (N_18986,N_17767,N_17474);
xor U18987 (N_18987,N_17269,N_16982);
nor U18988 (N_18988,N_16832,N_16919);
and U18989 (N_18989,N_17944,N_17197);
xnor U18990 (N_18990,N_17186,N_17745);
or U18991 (N_18991,N_17833,N_17625);
nor U18992 (N_18992,N_17309,N_17285);
nor U18993 (N_18993,N_17124,N_17277);
nand U18994 (N_18994,N_17053,N_17404);
and U18995 (N_18995,N_16827,N_17929);
or U18996 (N_18996,N_17264,N_17017);
nand U18997 (N_18997,N_17901,N_17997);
or U18998 (N_18998,N_17797,N_16956);
xor U18999 (N_18999,N_17708,N_17747);
or U19000 (N_19000,N_16971,N_17512);
nand U19001 (N_19001,N_17769,N_17671);
and U19002 (N_19002,N_17144,N_17431);
or U19003 (N_19003,N_17645,N_17051);
and U19004 (N_19004,N_17114,N_17498);
nand U19005 (N_19005,N_17128,N_16868);
and U19006 (N_19006,N_17255,N_17670);
or U19007 (N_19007,N_17389,N_17303);
xor U19008 (N_19008,N_17604,N_17496);
xor U19009 (N_19009,N_17143,N_17780);
xnor U19010 (N_19010,N_17906,N_17136);
xor U19011 (N_19011,N_17627,N_17591);
and U19012 (N_19012,N_16818,N_17476);
nor U19013 (N_19013,N_17265,N_17362);
xnor U19014 (N_19014,N_17277,N_17221);
or U19015 (N_19015,N_17207,N_17847);
nor U19016 (N_19016,N_16890,N_17116);
nor U19017 (N_19017,N_17417,N_17466);
nand U19018 (N_19018,N_17589,N_17522);
and U19019 (N_19019,N_17049,N_16904);
and U19020 (N_19020,N_17598,N_16930);
and U19021 (N_19021,N_16817,N_17299);
xor U19022 (N_19022,N_17587,N_17627);
xor U19023 (N_19023,N_17844,N_17343);
xor U19024 (N_19024,N_17259,N_17410);
or U19025 (N_19025,N_17403,N_17720);
xor U19026 (N_19026,N_17403,N_17144);
nor U19027 (N_19027,N_17103,N_17215);
nor U19028 (N_19028,N_17149,N_17885);
xor U19029 (N_19029,N_17054,N_17006);
and U19030 (N_19030,N_16849,N_17228);
nand U19031 (N_19031,N_17790,N_16810);
nand U19032 (N_19032,N_17599,N_17991);
and U19033 (N_19033,N_17300,N_17670);
nor U19034 (N_19034,N_17916,N_17757);
and U19035 (N_19035,N_17627,N_17772);
xor U19036 (N_19036,N_17856,N_17642);
nor U19037 (N_19037,N_17940,N_17668);
nor U19038 (N_19038,N_16825,N_16952);
and U19039 (N_19039,N_17546,N_17733);
or U19040 (N_19040,N_17897,N_17738);
xnor U19041 (N_19041,N_17505,N_16858);
nand U19042 (N_19042,N_17672,N_17973);
nand U19043 (N_19043,N_17940,N_17667);
nand U19044 (N_19044,N_17140,N_16982);
xor U19045 (N_19045,N_17076,N_17972);
or U19046 (N_19046,N_17260,N_17072);
or U19047 (N_19047,N_17924,N_17992);
nand U19048 (N_19048,N_17737,N_17026);
xnor U19049 (N_19049,N_16927,N_16844);
nand U19050 (N_19050,N_17448,N_17017);
xor U19051 (N_19051,N_17665,N_17857);
and U19052 (N_19052,N_17185,N_17239);
nor U19053 (N_19053,N_17239,N_17090);
or U19054 (N_19054,N_17010,N_17975);
or U19055 (N_19055,N_17344,N_17526);
xnor U19056 (N_19056,N_16885,N_17617);
nor U19057 (N_19057,N_17341,N_17573);
and U19058 (N_19058,N_17531,N_17484);
xnor U19059 (N_19059,N_17655,N_17458);
nor U19060 (N_19060,N_17538,N_17816);
xnor U19061 (N_19061,N_17229,N_17267);
and U19062 (N_19062,N_17182,N_17987);
nand U19063 (N_19063,N_17517,N_17330);
xnor U19064 (N_19064,N_17423,N_17119);
xor U19065 (N_19065,N_17778,N_17768);
or U19066 (N_19066,N_17999,N_17628);
and U19067 (N_19067,N_16965,N_17100);
nand U19068 (N_19068,N_17773,N_17110);
nand U19069 (N_19069,N_17542,N_17169);
nand U19070 (N_19070,N_17305,N_16957);
and U19071 (N_19071,N_16844,N_17421);
and U19072 (N_19072,N_17704,N_17077);
xor U19073 (N_19073,N_17907,N_17475);
nor U19074 (N_19074,N_17314,N_17341);
nand U19075 (N_19075,N_16906,N_17020);
xnor U19076 (N_19076,N_16860,N_17897);
nand U19077 (N_19077,N_17040,N_17211);
nor U19078 (N_19078,N_17451,N_17677);
or U19079 (N_19079,N_17632,N_17723);
and U19080 (N_19080,N_17859,N_17912);
xor U19081 (N_19081,N_17135,N_17473);
xor U19082 (N_19082,N_17003,N_17557);
or U19083 (N_19083,N_17485,N_17488);
nand U19084 (N_19084,N_17619,N_17123);
or U19085 (N_19085,N_17588,N_17280);
nand U19086 (N_19086,N_17291,N_16846);
xor U19087 (N_19087,N_17853,N_17911);
and U19088 (N_19088,N_17498,N_17620);
nand U19089 (N_19089,N_17578,N_17897);
and U19090 (N_19090,N_17271,N_17732);
xor U19091 (N_19091,N_17355,N_16895);
nand U19092 (N_19092,N_16806,N_16868);
xor U19093 (N_19093,N_16915,N_17048);
nand U19094 (N_19094,N_17928,N_17568);
nand U19095 (N_19095,N_17267,N_16959);
nor U19096 (N_19096,N_17993,N_17264);
nor U19097 (N_19097,N_17233,N_17929);
nor U19098 (N_19098,N_17990,N_17187);
xor U19099 (N_19099,N_16930,N_16987);
nand U19100 (N_19100,N_17095,N_17451);
nand U19101 (N_19101,N_17501,N_17594);
nor U19102 (N_19102,N_17064,N_17601);
or U19103 (N_19103,N_17541,N_17120);
nor U19104 (N_19104,N_17484,N_17838);
xor U19105 (N_19105,N_17295,N_17964);
or U19106 (N_19106,N_16907,N_17501);
nor U19107 (N_19107,N_17429,N_16984);
xnor U19108 (N_19108,N_17293,N_17058);
nand U19109 (N_19109,N_17882,N_17434);
nor U19110 (N_19110,N_17770,N_17311);
nor U19111 (N_19111,N_17667,N_17632);
nor U19112 (N_19112,N_17738,N_16994);
or U19113 (N_19113,N_17103,N_17422);
nand U19114 (N_19114,N_17101,N_17828);
and U19115 (N_19115,N_16989,N_17184);
nor U19116 (N_19116,N_17855,N_17858);
or U19117 (N_19117,N_17791,N_17678);
or U19118 (N_19118,N_17050,N_17910);
and U19119 (N_19119,N_17270,N_17493);
nand U19120 (N_19120,N_17797,N_17392);
nor U19121 (N_19121,N_17696,N_17667);
and U19122 (N_19122,N_17915,N_17674);
nand U19123 (N_19123,N_17652,N_17552);
xor U19124 (N_19124,N_17586,N_17212);
xor U19125 (N_19125,N_16980,N_17758);
nor U19126 (N_19126,N_17586,N_17566);
and U19127 (N_19127,N_17254,N_17640);
nor U19128 (N_19128,N_17389,N_17606);
nand U19129 (N_19129,N_17247,N_16801);
xnor U19130 (N_19130,N_17223,N_17359);
xor U19131 (N_19131,N_16911,N_16831);
nor U19132 (N_19132,N_17436,N_17492);
and U19133 (N_19133,N_17343,N_16814);
and U19134 (N_19134,N_17267,N_17834);
nand U19135 (N_19135,N_17535,N_17168);
xor U19136 (N_19136,N_17110,N_17615);
nand U19137 (N_19137,N_16815,N_17476);
nor U19138 (N_19138,N_16803,N_17137);
nand U19139 (N_19139,N_17395,N_17006);
xor U19140 (N_19140,N_17724,N_17684);
xor U19141 (N_19141,N_17644,N_17393);
xor U19142 (N_19142,N_16982,N_17054);
xnor U19143 (N_19143,N_16801,N_16994);
and U19144 (N_19144,N_17255,N_17598);
or U19145 (N_19145,N_16966,N_17151);
or U19146 (N_19146,N_17451,N_17397);
nor U19147 (N_19147,N_17789,N_16979);
xor U19148 (N_19148,N_17308,N_17442);
and U19149 (N_19149,N_17400,N_17658);
or U19150 (N_19150,N_17428,N_16903);
nand U19151 (N_19151,N_17538,N_17690);
nor U19152 (N_19152,N_17164,N_17604);
nor U19153 (N_19153,N_16977,N_17528);
or U19154 (N_19154,N_16953,N_17697);
xor U19155 (N_19155,N_17331,N_17215);
xor U19156 (N_19156,N_17894,N_17832);
xor U19157 (N_19157,N_17377,N_17563);
or U19158 (N_19158,N_16821,N_16838);
nor U19159 (N_19159,N_17398,N_17636);
nand U19160 (N_19160,N_17937,N_17516);
and U19161 (N_19161,N_17190,N_17312);
nor U19162 (N_19162,N_17215,N_17164);
or U19163 (N_19163,N_17877,N_16986);
xnor U19164 (N_19164,N_16871,N_16999);
or U19165 (N_19165,N_17707,N_17288);
nand U19166 (N_19166,N_17012,N_17229);
xor U19167 (N_19167,N_17494,N_17162);
xnor U19168 (N_19168,N_17194,N_17690);
nor U19169 (N_19169,N_17957,N_16970);
nor U19170 (N_19170,N_17481,N_17452);
nand U19171 (N_19171,N_16886,N_17253);
xor U19172 (N_19172,N_17096,N_17431);
and U19173 (N_19173,N_17513,N_17237);
or U19174 (N_19174,N_17150,N_17249);
xnor U19175 (N_19175,N_16946,N_16814);
and U19176 (N_19176,N_16900,N_17645);
and U19177 (N_19177,N_17762,N_17339);
and U19178 (N_19178,N_17197,N_17902);
nor U19179 (N_19179,N_17396,N_17286);
and U19180 (N_19180,N_17829,N_17091);
nor U19181 (N_19181,N_17566,N_16883);
xnor U19182 (N_19182,N_17089,N_17986);
and U19183 (N_19183,N_17710,N_17627);
xnor U19184 (N_19184,N_16968,N_16872);
nor U19185 (N_19185,N_16971,N_17879);
xor U19186 (N_19186,N_17503,N_17216);
xor U19187 (N_19187,N_17939,N_17636);
or U19188 (N_19188,N_17635,N_17267);
xnor U19189 (N_19189,N_17808,N_16836);
xor U19190 (N_19190,N_17777,N_17209);
or U19191 (N_19191,N_17135,N_17529);
or U19192 (N_19192,N_17614,N_17506);
nor U19193 (N_19193,N_17692,N_17846);
nand U19194 (N_19194,N_17993,N_17060);
or U19195 (N_19195,N_17188,N_17693);
xor U19196 (N_19196,N_17942,N_17905);
xor U19197 (N_19197,N_17729,N_17273);
xnor U19198 (N_19198,N_16834,N_17951);
nor U19199 (N_19199,N_17369,N_17557);
and U19200 (N_19200,N_18592,N_19149);
or U19201 (N_19201,N_18033,N_18569);
nor U19202 (N_19202,N_18908,N_18965);
nand U19203 (N_19203,N_18882,N_18359);
nor U19204 (N_19204,N_18385,N_19167);
nand U19205 (N_19205,N_19101,N_18835);
and U19206 (N_19206,N_18585,N_18500);
nand U19207 (N_19207,N_18910,N_18373);
and U19208 (N_19208,N_18217,N_18461);
and U19209 (N_19209,N_19145,N_18184);
and U19210 (N_19210,N_18686,N_18090);
nand U19211 (N_19211,N_18327,N_18788);
or U19212 (N_19212,N_18924,N_18824);
nand U19213 (N_19213,N_18257,N_18319);
or U19214 (N_19214,N_18392,N_18915);
and U19215 (N_19215,N_18346,N_18450);
and U19216 (N_19216,N_19059,N_18503);
xnor U19217 (N_19217,N_18622,N_18008);
or U19218 (N_19218,N_18940,N_18984);
or U19219 (N_19219,N_19098,N_18037);
nand U19220 (N_19220,N_18260,N_18493);
xor U19221 (N_19221,N_19150,N_19161);
or U19222 (N_19222,N_19136,N_18634);
or U19223 (N_19223,N_18961,N_18483);
and U19224 (N_19224,N_18253,N_18064);
xnor U19225 (N_19225,N_18818,N_18449);
nand U19226 (N_19226,N_18360,N_19164);
or U19227 (N_19227,N_18967,N_18110);
nand U19228 (N_19228,N_19188,N_19192);
nand U19229 (N_19229,N_19093,N_18609);
or U19230 (N_19230,N_18689,N_18921);
and U19231 (N_19231,N_18925,N_18696);
nand U19232 (N_19232,N_18939,N_18790);
and U19233 (N_19233,N_18948,N_18866);
nor U19234 (N_19234,N_18863,N_18955);
xor U19235 (N_19235,N_18928,N_18776);
or U19236 (N_19236,N_19115,N_18869);
and U19237 (N_19237,N_18054,N_18862);
xor U19238 (N_19238,N_19199,N_18071);
xnor U19239 (N_19239,N_18840,N_19133);
nor U19240 (N_19240,N_19050,N_19006);
or U19241 (N_19241,N_18045,N_18743);
or U19242 (N_19242,N_18182,N_18584);
or U19243 (N_19243,N_18263,N_19086);
nor U19244 (N_19244,N_18521,N_19121);
xnor U19245 (N_19245,N_19124,N_18886);
nor U19246 (N_19246,N_18390,N_18951);
xor U19247 (N_19247,N_18301,N_18713);
nand U19248 (N_19248,N_18844,N_18799);
and U19249 (N_19249,N_18411,N_19159);
xor U19250 (N_19250,N_19062,N_18953);
xor U19251 (N_19251,N_18593,N_18982);
xnor U19252 (N_19252,N_18185,N_18504);
and U19253 (N_19253,N_18399,N_18073);
nand U19254 (N_19254,N_18701,N_18752);
nor U19255 (N_19255,N_18100,N_18662);
and U19256 (N_19256,N_18415,N_18465);
and U19257 (N_19257,N_19032,N_18375);
and U19258 (N_19258,N_18349,N_18439);
and U19259 (N_19259,N_18499,N_18561);
and U19260 (N_19260,N_18291,N_18116);
nand U19261 (N_19261,N_18995,N_18758);
nand U19262 (N_19262,N_18270,N_18739);
and U19263 (N_19263,N_18698,N_18983);
nor U19264 (N_19264,N_18423,N_18909);
nand U19265 (N_19265,N_18446,N_18672);
nor U19266 (N_19266,N_18014,N_18784);
nor U19267 (N_19267,N_18136,N_18543);
or U19268 (N_19268,N_19076,N_18538);
nand U19269 (N_19269,N_18141,N_19047);
nor U19270 (N_19270,N_18825,N_18205);
nor U19271 (N_19271,N_18254,N_18345);
xnor U19272 (N_19272,N_18552,N_18297);
nand U19273 (N_19273,N_18239,N_18936);
or U19274 (N_19274,N_18053,N_18657);
xnor U19275 (N_19275,N_18566,N_18229);
nand U19276 (N_19276,N_18860,N_18979);
nand U19277 (N_19277,N_18645,N_18002);
xor U19278 (N_19278,N_18626,N_18681);
nor U19279 (N_19279,N_18087,N_18625);
nand U19280 (N_19280,N_18410,N_18639);
or U19281 (N_19281,N_19118,N_18877);
or U19282 (N_19282,N_18188,N_18803);
or U19283 (N_19283,N_18588,N_18150);
nand U19284 (N_19284,N_18582,N_18800);
and U19285 (N_19285,N_19169,N_18200);
nand U19286 (N_19286,N_18772,N_18997);
and U19287 (N_19287,N_19095,N_18697);
nand U19288 (N_19288,N_18378,N_18206);
or U19289 (N_19289,N_18601,N_18541);
xor U19290 (N_19290,N_18989,N_19168);
or U19291 (N_19291,N_18782,N_18711);
nor U19292 (N_19292,N_19067,N_18880);
xnor U19293 (N_19293,N_19162,N_18660);
and U19294 (N_19294,N_18666,N_18655);
xnor U19295 (N_19295,N_18082,N_18377);
or U19296 (N_19296,N_18421,N_18658);
nor U19297 (N_19297,N_18092,N_18751);
xor U19298 (N_19298,N_18337,N_18514);
xor U19299 (N_19299,N_18821,N_18613);
nor U19300 (N_19300,N_18780,N_18210);
nand U19301 (N_19301,N_18748,N_18023);
nor U19302 (N_19302,N_18395,N_18475);
or U19303 (N_19303,N_19141,N_18786);
nand U19304 (N_19304,N_18534,N_19019);
nor U19305 (N_19305,N_19097,N_18550);
nand U19306 (N_19306,N_19185,N_18633);
and U19307 (N_19307,N_18520,N_19198);
nor U19308 (N_19308,N_19001,N_18652);
and U19309 (N_19309,N_19166,N_18610);
xor U19310 (N_19310,N_19132,N_18098);
and U19311 (N_19311,N_18874,N_18604);
xnor U19312 (N_19312,N_19057,N_18460);
nor U19313 (N_19313,N_19137,N_19108);
xor U19314 (N_19314,N_19143,N_18306);
xor U19315 (N_19315,N_18553,N_18564);
and U19316 (N_19316,N_18669,N_18467);
nor U19317 (N_19317,N_18224,N_18762);
or U19318 (N_19318,N_18730,N_18489);
and U19319 (N_19319,N_18030,N_19060);
nand U19320 (N_19320,N_18854,N_18196);
nand U19321 (N_19321,N_18436,N_18498);
and U19322 (N_19322,N_18783,N_18557);
or U19323 (N_19323,N_19134,N_18817);
and U19324 (N_19324,N_18080,N_18403);
or U19325 (N_19325,N_19154,N_18878);
nor U19326 (N_19326,N_18061,N_18548);
xor U19327 (N_19327,N_18187,N_18820);
nor U19328 (N_19328,N_18382,N_19068);
nor U19329 (N_19329,N_18275,N_18024);
or U19330 (N_19330,N_18941,N_19195);
or U19331 (N_19331,N_18488,N_18281);
nor U19332 (N_19332,N_19158,N_18268);
nand U19333 (N_19333,N_18340,N_18511);
or U19334 (N_19334,N_18323,N_18114);
xnor U19335 (N_19335,N_18213,N_18770);
xnor U19336 (N_19336,N_18810,N_18348);
nor U19337 (N_19337,N_19025,N_18962);
or U19338 (N_19338,N_19085,N_19171);
or U19339 (N_19339,N_18353,N_18219);
xnor U19340 (N_19340,N_18177,N_18842);
nor U19341 (N_19341,N_18393,N_18523);
nand U19342 (N_19342,N_18019,N_18547);
or U19343 (N_19343,N_19042,N_18966);
nor U19344 (N_19344,N_18321,N_18903);
xnor U19345 (N_19345,N_18599,N_18331);
nand U19346 (N_19346,N_18906,N_18675);
nor U19347 (N_19347,N_18285,N_18777);
nand U19348 (N_19348,N_18357,N_18001);
or U19349 (N_19349,N_18478,N_18401);
and U19350 (N_19350,N_18320,N_18720);
nor U19351 (N_19351,N_18883,N_18247);
nor U19352 (N_19352,N_18424,N_18282);
and U19353 (N_19353,N_18137,N_18428);
nor U19354 (N_19354,N_18513,N_18994);
and U19355 (N_19355,N_18248,N_18108);
and U19356 (N_19356,N_18245,N_18085);
nor U19357 (N_19357,N_18069,N_18572);
nand U19358 (N_19358,N_18383,N_18335);
nor U19359 (N_19359,N_18620,N_19036);
and U19360 (N_19360,N_18964,N_18204);
or U19361 (N_19361,N_18916,N_18041);
and U19362 (N_19362,N_18885,N_18149);
xnor U19363 (N_19363,N_18771,N_18744);
xnor U19364 (N_19364,N_19135,N_18822);
or U19365 (N_19365,N_18304,N_18084);
nor U19366 (N_19366,N_18811,N_18929);
or U19367 (N_19367,N_19090,N_18011);
nor U19368 (N_19368,N_18841,N_18067);
and U19369 (N_19369,N_18186,N_18351);
nor U19370 (N_19370,N_18389,N_18221);
and U19371 (N_19371,N_18457,N_18753);
nor U19372 (N_19372,N_18443,N_18191);
nand U19373 (N_19373,N_18950,N_19183);
nor U19374 (N_19374,N_18009,N_19012);
nand U19375 (N_19375,N_18872,N_18207);
and U19376 (N_19376,N_18105,N_18693);
nor U19377 (N_19377,N_18524,N_18763);
or U19378 (N_19378,N_19088,N_18554);
nand U19379 (N_19379,N_18025,N_18040);
xor U19380 (N_19380,N_19079,N_18352);
nor U19381 (N_19381,N_18220,N_18235);
and U19382 (N_19382,N_18325,N_19146);
nor U19383 (N_19383,N_18830,N_18691);
nor U19384 (N_19384,N_19151,N_18234);
and U19385 (N_19385,N_18904,N_18459);
nand U19386 (N_19386,N_18451,N_18202);
nand U19387 (N_19387,N_18945,N_18138);
nor U19388 (N_19388,N_18227,N_18287);
xor U19389 (N_19389,N_18126,N_19038);
xor U19390 (N_19390,N_18688,N_18463);
and U19391 (N_19391,N_18232,N_18153);
and U19392 (N_19392,N_18250,N_19152);
or U19393 (N_19393,N_18692,N_18759);
xnor U19394 (N_19394,N_18198,N_18725);
or U19395 (N_19395,N_19089,N_18454);
and U19396 (N_19396,N_18448,N_18761);
and U19397 (N_19397,N_19070,N_18833);
and U19398 (N_19398,N_18708,N_19071);
nand U19399 (N_19399,N_18308,N_18881);
xor U19400 (N_19400,N_19084,N_18670);
or U19401 (N_19401,N_18211,N_18288);
and U19402 (N_19402,N_18259,N_18152);
or U19403 (N_19403,N_18839,N_18852);
nor U19404 (N_19404,N_18704,N_18322);
nor U19405 (N_19405,N_18571,N_18021);
xor U19406 (N_19406,N_19147,N_18875);
and U19407 (N_19407,N_18684,N_18103);
and U19408 (N_19408,N_18059,N_18712);
nand U19409 (N_19409,N_18189,N_18855);
xor U19410 (N_19410,N_18314,N_18627);
nand U19411 (N_19411,N_18266,N_18765);
nand U19412 (N_19412,N_18076,N_18891);
xnor U19413 (N_19413,N_18931,N_18476);
or U19414 (N_19414,N_18764,N_18212);
nand U19415 (N_19415,N_18974,N_18918);
xor U19416 (N_19416,N_18118,N_18174);
nand U19417 (N_19417,N_18749,N_18055);
or U19418 (N_19418,N_19160,N_18365);
nand U19419 (N_19419,N_18612,N_18618);
xnor U19420 (N_19420,N_18063,N_19120);
nor U19421 (N_19421,N_18699,N_18674);
or U19422 (N_19422,N_18829,N_19096);
nand U19423 (N_19423,N_18649,N_18381);
xnor U19424 (N_19424,N_18496,N_18721);
nand U19425 (N_19425,N_18058,N_18180);
xnor U19426 (N_19426,N_18156,N_18723);
nand U19427 (N_19427,N_19181,N_19055);
or U19428 (N_19428,N_18330,N_18968);
nand U19429 (N_19429,N_18583,N_18066);
nand U19430 (N_19430,N_18237,N_18350);
xor U19431 (N_19431,N_19191,N_18119);
nand U19432 (N_19432,N_18298,N_18522);
and U19433 (N_19433,N_18176,N_18648);
nand U19434 (N_19434,N_18201,N_18473);
and U19435 (N_19435,N_18106,N_18386);
and U19436 (N_19436,N_18034,N_18826);
nand U19437 (N_19437,N_18536,N_18683);
and U19438 (N_19438,N_18754,N_18431);
or U19439 (N_19439,N_18068,N_18981);
nor U19440 (N_19440,N_18740,N_18396);
or U19441 (N_19441,N_18163,N_19029);
or U19442 (N_19442,N_18151,N_18732);
xnor U19443 (N_19443,N_18570,N_18900);
and U19444 (N_19444,N_18603,N_19107);
nand U19445 (N_19445,N_18927,N_18052);
nand U19446 (N_19446,N_18539,N_18663);
and U19447 (N_19447,N_19010,N_18495);
or U19448 (N_19448,N_19129,N_18518);
or U19449 (N_19449,N_18121,N_18678);
or U19450 (N_19450,N_18728,N_18047);
or U19451 (N_19451,N_19005,N_18228);
or U19452 (N_19452,N_18175,N_18781);
and U19453 (N_19453,N_18142,N_18930);
or U19454 (N_19454,N_18072,N_18404);
or U19455 (N_19455,N_18208,N_19112);
and U19456 (N_19456,N_18233,N_18241);
and U19457 (N_19457,N_18792,N_18089);
nor U19458 (N_19458,N_18414,N_18707);
nand U19459 (N_19459,N_18850,N_18644);
xnor U19460 (N_19460,N_18356,N_19189);
and U19461 (N_19461,N_19065,N_18664);
nor U19462 (N_19462,N_18214,N_18022);
xor U19463 (N_19463,N_18734,N_18292);
or U19464 (N_19464,N_18480,N_19073);
nor U19465 (N_19465,N_19049,N_19123);
nand U19466 (N_19466,N_18647,N_18530);
nor U19467 (N_19467,N_18278,N_19190);
or U19468 (N_19468,N_18370,N_18120);
or U19469 (N_19469,N_18636,N_18243);
or U19470 (N_19470,N_18244,N_18231);
xnor U19471 (N_19471,N_18051,N_18296);
or U19472 (N_19472,N_18172,N_18785);
and U19473 (N_19473,N_18102,N_19187);
xor U19474 (N_19474,N_18261,N_18629);
nand U19475 (N_19475,N_18432,N_18474);
xor U19476 (N_19476,N_18774,N_18124);
nand U19477 (N_19477,N_18486,N_18887);
xnor U19478 (N_19478,N_18796,N_18471);
nor U19479 (N_19479,N_19034,N_18549);
nor U19480 (N_19480,N_19082,N_18902);
nor U19481 (N_19481,N_19061,N_18843);
or U19482 (N_19482,N_18715,N_18256);
xor U19483 (N_19483,N_18746,N_18814);
and U19484 (N_19484,N_19083,N_19178);
nor U19485 (N_19485,N_18895,N_18420);
and U19486 (N_19486,N_18433,N_18870);
nand U19487 (N_19487,N_18363,N_18508);
and U19488 (N_19488,N_18238,N_18767);
nor U19489 (N_19489,N_19156,N_18075);
nand U19490 (N_19490,N_18628,N_18230);
or U19491 (N_19491,N_18417,N_18005);
and U19492 (N_19492,N_19155,N_18606);
and U19493 (N_19493,N_18650,N_19116);
or U19494 (N_19494,N_18766,N_18893);
xnor U19495 (N_19495,N_19018,N_19144);
xnor U19496 (N_19496,N_18544,N_18668);
xor U19497 (N_19497,N_18440,N_18032);
and U19498 (N_19498,N_18405,N_18990);
or U19499 (N_19499,N_18409,N_19008);
nor U19500 (N_19500,N_18289,N_18805);
xnor U19501 (N_19501,N_19002,N_18344);
and U19502 (N_19502,N_18309,N_18249);
and U19503 (N_19503,N_19125,N_18959);
or U19504 (N_19504,N_18577,N_18343);
nand U19505 (N_19505,N_18970,N_18737);
and U19506 (N_19506,N_18507,N_18223);
and U19507 (N_19507,N_18050,N_19028);
or U19508 (N_19508,N_18795,N_18651);
or U19509 (N_19509,N_18797,N_18605);
or U19510 (N_19510,N_18576,N_18438);
nor U19511 (N_19511,N_19026,N_18608);
xor U19512 (N_19512,N_19023,N_18515);
or U19513 (N_19513,N_18097,N_18416);
nor U19514 (N_19514,N_19109,N_18303);
nor U19515 (N_19515,N_18659,N_18775);
and U19516 (N_19516,N_19100,N_18726);
or U19517 (N_19517,N_18857,N_18132);
nand U19518 (N_19518,N_18876,N_18333);
nand U19519 (N_19519,N_18954,N_18901);
xor U19520 (N_19520,N_18773,N_18859);
and U19521 (N_19521,N_18718,N_18717);
or U19522 (N_19522,N_18445,N_18646);
xor U19523 (N_19523,N_18526,N_18996);
and U19524 (N_19524,N_19148,N_18255);
nor U19525 (N_19525,N_18004,N_18258);
xnor U19526 (N_19526,N_18505,N_19051);
nand U19527 (N_19527,N_18745,N_19003);
or U19528 (N_19528,N_19126,N_18640);
or U19529 (N_19529,N_18510,N_18943);
xor U19530 (N_19530,N_18398,N_18162);
nor U19531 (N_19531,N_18133,N_19091);
xor U19532 (N_19532,N_18435,N_18529);
nand U19533 (N_19533,N_18044,N_18595);
xnor U19534 (N_19534,N_18519,N_18560);
nor U19535 (N_19535,N_18685,N_18006);
or U19536 (N_19536,N_19110,N_18594);
and U19537 (N_19537,N_18779,N_18299);
or U19538 (N_19538,N_18896,N_18284);
or U19539 (N_19539,N_18159,N_18179);
nand U19540 (N_19540,N_18706,N_18123);
nor U19541 (N_19541,N_18768,N_18099);
or U19542 (N_19542,N_18919,N_18867);
nand U19543 (N_19543,N_19046,N_18656);
nand U19544 (N_19544,N_18987,N_18332);
and U19545 (N_19545,N_19017,N_18171);
xnor U19546 (N_19546,N_18049,N_18935);
nand U19547 (N_19547,N_18086,N_18980);
xnor U19548 (N_19548,N_18828,N_18148);
nand U19549 (N_19549,N_18374,N_18665);
xor U19550 (N_19550,N_19111,N_18978);
or U19551 (N_19551,N_18532,N_18568);
nor U19552 (N_19552,N_18048,N_18949);
nor U19553 (N_19553,N_19072,N_18369);
nand U19554 (N_19554,N_18671,N_19015);
nand U19555 (N_19555,N_18551,N_18621);
or U19556 (N_19556,N_19022,N_18018);
xor U19557 (N_19557,N_18139,N_18376);
and U19558 (N_19558,N_18484,N_18798);
and U19559 (N_19559,N_18899,N_19194);
and U19560 (N_19560,N_19014,N_19000);
or U19561 (N_19561,N_18203,N_18026);
and U19562 (N_19562,N_18305,N_18236);
nand U19563 (N_19563,N_18641,N_18992);
and U19564 (N_19564,N_19064,N_18556);
xor U19565 (N_19565,N_18264,N_18165);
xor U19566 (N_19566,N_18479,N_18611);
xnor U19567 (N_19567,N_18324,N_18093);
nand U19568 (N_19568,N_18000,N_18988);
xor U19569 (N_19569,N_18755,N_18400);
nor U19570 (N_19570,N_18199,N_18317);
or U19571 (N_19571,N_19182,N_18274);
nor U19572 (N_19572,N_18487,N_18341);
or U19573 (N_19573,N_19139,N_18328);
or U19574 (N_19574,N_18590,N_18143);
and U19575 (N_19575,N_18555,N_19104);
nand U19576 (N_19576,N_18157,N_19165);
xor U19577 (N_19577,N_18756,N_18338);
or U19578 (N_19578,N_18193,N_19021);
nor U19579 (N_19579,N_18430,N_18028);
xnor U19580 (N_19580,N_19011,N_18716);
and U19581 (N_19581,N_18631,N_18591);
xor U19582 (N_19582,N_18074,N_18969);
nand U19583 (N_19583,N_18013,N_18834);
xnor U19584 (N_19584,N_18267,N_18702);
nand U19585 (N_19585,N_18942,N_18868);
and U19586 (N_19586,N_18455,N_18907);
or U19587 (N_19587,N_18687,N_18750);
and U19588 (N_19588,N_18837,N_18793);
nor U19589 (N_19589,N_18293,N_18643);
nor U19590 (N_19590,N_18190,N_18789);
or U19591 (N_19591,N_18889,N_18388);
xnor U19592 (N_19592,N_19024,N_18963);
nand U19593 (N_19593,N_18589,N_18131);
nor U19594 (N_19594,N_18676,N_19138);
and U19595 (N_19595,N_18957,N_18482);
xnor U19596 (N_19596,N_18537,N_18397);
nand U19597 (N_19597,N_18690,N_18160);
xor U19598 (N_19598,N_18312,N_18525);
and U19599 (N_19599,N_18823,N_18240);
nand U19600 (N_19600,N_18361,N_18279);
nand U19601 (N_19601,N_18661,N_18181);
xnor U19602 (N_19602,N_18413,N_18700);
nor U19603 (N_19603,N_18884,N_18911);
or U19604 (N_19604,N_18845,N_18677);
nand U19605 (N_19605,N_18574,N_18973);
and U19606 (N_19606,N_18029,N_19007);
and U19607 (N_19607,N_19106,N_18587);
nor U19608 (N_19608,N_18441,N_19170);
nand U19609 (N_19609,N_18342,N_18812);
nand U19610 (N_19610,N_18986,N_18134);
nand U19611 (N_19611,N_18563,N_18472);
or U19612 (N_19612,N_18705,N_18020);
xor U19613 (N_19613,N_18466,N_18926);
and U19614 (N_19614,N_18747,N_18161);
xnor U19615 (N_19615,N_19113,N_18222);
nand U19616 (N_19616,N_18956,N_18735);
nand U19617 (N_19617,N_18540,N_18827);
xor U19618 (N_19618,N_18873,N_18946);
and U19619 (N_19619,N_18364,N_18637);
nand U19620 (N_19620,N_19080,N_18917);
or U19621 (N_19621,N_19043,N_19041);
and U19622 (N_19622,N_18046,N_19066);
or U19623 (N_19623,N_18502,N_18083);
and U19624 (N_19624,N_18311,N_18632);
nor U19625 (N_19625,N_19027,N_18497);
xor U19626 (N_19626,N_18079,N_19016);
or U19627 (N_19627,N_18434,N_18853);
and U19628 (N_19628,N_19174,N_18512);
and U19629 (N_19629,N_18458,N_18010);
or U19630 (N_19630,N_18277,N_18336);
and U19631 (N_19631,N_19172,N_18933);
or U19632 (N_19632,N_19056,N_18517);
nand U19633 (N_19633,N_18295,N_19130);
nand U19634 (N_19634,N_18262,N_18856);
nand U19635 (N_19635,N_18422,N_19102);
nor U19636 (N_19636,N_18290,N_18894);
xnor U19637 (N_19637,N_18562,N_19092);
nor U19638 (N_19638,N_18742,N_18168);
xnor U19639 (N_19639,N_18130,N_19037);
xnor U19640 (N_19640,N_18580,N_18003);
xor U19641 (N_19641,N_18115,N_18146);
and U19642 (N_19642,N_18307,N_19031);
nand U19643 (N_19643,N_18367,N_18602);
and U19644 (N_19644,N_18491,N_18846);
xor U19645 (N_19645,N_18791,N_18838);
nand U19646 (N_19646,N_18104,N_18682);
nor U19647 (N_19647,N_18947,N_18958);
nor U19648 (N_19648,N_18107,N_18932);
and U19649 (N_19649,N_19004,N_19075);
and U19650 (N_19650,N_18937,N_18719);
and U19651 (N_19651,N_19053,N_18294);
nand U19652 (N_19652,N_18081,N_18310);
and U19653 (N_19653,N_18729,N_18347);
nor U19654 (N_19654,N_19074,N_18273);
or U19655 (N_19655,N_19058,N_18944);
nand U19656 (N_19656,N_19009,N_18453);
xnor U19657 (N_19657,N_18418,N_18192);
or U19658 (N_19658,N_18265,N_18506);
nor U19659 (N_19659,N_18226,N_19119);
xnor U19660 (N_19660,N_18898,N_19197);
nor U19661 (N_19661,N_19122,N_18147);
xor U19662 (N_19662,N_18427,N_19114);
or U19663 (N_19663,N_19063,N_18913);
nor U19664 (N_19664,N_18122,N_18531);
xnor U19665 (N_19665,N_18575,N_18581);
nand U19666 (N_19666,N_18437,N_18225);
or U19667 (N_19667,N_18060,N_18615);
nand U19668 (N_19668,N_18429,N_18813);
nor U19669 (N_19669,N_18985,N_18709);
or U19670 (N_19670,N_18135,N_18128);
nand U19671 (N_19671,N_19142,N_18039);
and U19672 (N_19672,N_18425,N_18406);
nor U19673 (N_19673,N_18394,N_19081);
nor U19674 (N_19674,N_18036,N_18816);
nand U19675 (N_19675,N_18195,N_18109);
nor U19676 (N_19676,N_18140,N_18999);
nor U19677 (N_19677,N_18283,N_19040);
xor U19678 (N_19678,N_18975,N_18366);
xor U19679 (N_19679,N_19127,N_18412);
nand U19680 (N_19680,N_18616,N_19153);
nor U19681 (N_19681,N_18111,N_18065);
and U19682 (N_19682,N_18462,N_18694);
nand U19683 (N_19683,N_18167,N_18905);
nor U19684 (N_19684,N_19048,N_18056);
or U19685 (N_19685,N_18464,N_18070);
and U19686 (N_19686,N_18738,N_18447);
nor U19687 (N_19687,N_19103,N_18490);
xor U19688 (N_19688,N_18316,N_18861);
or U19689 (N_19689,N_18442,N_18078);
xor U19690 (N_19690,N_18088,N_19128);
or U19691 (N_19691,N_18733,N_18533);
and U19692 (N_19692,N_18456,N_18091);
or U19693 (N_19693,N_19039,N_18218);
nor U19694 (N_19694,N_18815,N_19054);
and U19695 (N_19695,N_18173,N_18057);
and U19696 (N_19696,N_18545,N_18888);
nor U19697 (N_19697,N_18848,N_18251);
nor U19698 (N_19698,N_18624,N_18565);
xnor U19699 (N_19699,N_18242,N_18809);
xor U19700 (N_19700,N_18879,N_18871);
nor U19701 (N_19701,N_19157,N_18623);
xor U19702 (N_19702,N_18912,N_18741);
and U19703 (N_19703,N_18127,N_18642);
or U19704 (N_19704,N_18354,N_18546);
and U19705 (N_19705,N_18673,N_18667);
nand U19706 (N_19706,N_18960,N_18819);
and U19707 (N_19707,N_18778,N_18807);
and U19708 (N_19708,N_18976,N_18695);
xor U19709 (N_19709,N_18444,N_18371);
or U19710 (N_19710,N_19069,N_18043);
or U19711 (N_19711,N_18408,N_18329);
or U19712 (N_19712,N_19193,N_18528);
xnor U19713 (N_19713,N_18481,N_19094);
or U19714 (N_19714,N_18272,N_19078);
or U19715 (N_19715,N_18892,N_18679);
nand U19716 (N_19716,N_18865,N_19177);
nor U19717 (N_19717,N_18760,N_18169);
and U19718 (N_19718,N_18722,N_18971);
nor U19719 (N_19719,N_18897,N_19140);
nand U19720 (N_19720,N_18535,N_18558);
xnor U19721 (N_19721,N_18596,N_19087);
and U19722 (N_19722,N_18035,N_19020);
or U19723 (N_19723,N_19179,N_18802);
xor U19724 (N_19724,N_18952,N_19045);
nand U19725 (N_19725,N_18164,N_18938);
nor U19726 (N_19726,N_18178,N_18315);
and U19727 (N_19727,N_18858,N_18586);
xnor U19728 (N_19728,N_19163,N_19131);
nor U19729 (N_19729,N_18600,N_18326);
xor U19730 (N_19730,N_18527,N_18362);
or U19731 (N_19731,N_18559,N_18017);
xnor U19732 (N_19732,N_18358,N_18801);
xor U19733 (N_19733,N_18934,N_19033);
nand U19734 (N_19734,N_18607,N_18276);
and U19735 (N_19735,N_18567,N_18155);
and U19736 (N_19736,N_18113,N_18387);
or U19737 (N_19737,N_19077,N_18972);
or U19738 (N_19738,N_18578,N_18516);
and U19739 (N_19739,N_18710,N_18501);
nor U19740 (N_19740,N_18391,N_18492);
nor U19741 (N_19741,N_18731,N_18339);
nor U19742 (N_19742,N_19013,N_19180);
nor U19743 (N_19743,N_18380,N_18630);
xnor U19744 (N_19744,N_18101,N_18714);
and U19745 (N_19745,N_18419,N_18094);
nand U19746 (N_19746,N_18470,N_18635);
or U19747 (N_19747,N_18183,N_18724);
or U19748 (N_19748,N_18619,N_18468);
nand U19749 (N_19749,N_18145,N_18804);
nor U19750 (N_19750,N_18015,N_18334);
xnor U19751 (N_19751,N_18653,N_18313);
or U19752 (N_19752,N_18112,N_18031);
xnor U19753 (N_19753,N_18757,N_18209);
xor U19754 (N_19754,N_18703,N_18977);
nand U19755 (N_19755,N_18077,N_18271);
nand U19756 (N_19756,N_18194,N_18379);
nand U19757 (N_19757,N_18832,N_18847);
nor U19758 (N_19758,N_18166,N_18372);
or U19759 (N_19759,N_18614,N_18402);
nand U19760 (N_19760,N_18849,N_18864);
and U19761 (N_19761,N_19173,N_18318);
or U19762 (N_19762,N_18579,N_18246);
nor U19763 (N_19763,N_18477,N_18542);
xnor U19764 (N_19764,N_19099,N_19117);
nand U19765 (N_19765,N_18831,N_18042);
and U19766 (N_19766,N_18993,N_18158);
nand U19767 (N_19767,N_19176,N_18426);
and U19768 (N_19768,N_18851,N_18573);
nand U19769 (N_19769,N_18407,N_18736);
or U19770 (N_19770,N_18787,N_18890);
or U19771 (N_19771,N_18598,N_18355);
and U19772 (N_19772,N_18794,N_18197);
and U19773 (N_19773,N_19030,N_18144);
nand U19774 (N_19774,N_18680,N_18914);
xor U19775 (N_19775,N_18012,N_18920);
xor U19776 (N_19776,N_18129,N_18007);
xor U19777 (N_19777,N_19196,N_18300);
and U19778 (N_19778,N_18808,N_19052);
or U19779 (N_19779,N_18727,N_18095);
and U19780 (N_19780,N_19175,N_18998);
nand U19781 (N_19781,N_18368,N_18269);
nand U19782 (N_19782,N_18154,N_18016);
nand U19783 (N_19783,N_18485,N_18991);
nor U19784 (N_19784,N_19105,N_19186);
nor U19785 (N_19785,N_19044,N_18062);
nor U19786 (N_19786,N_19035,N_18302);
xnor U19787 (N_19787,N_18286,N_18038);
nand U19788 (N_19788,N_18836,N_18922);
nor U19789 (N_19789,N_18452,N_18494);
or U19790 (N_19790,N_19184,N_18027);
or U19791 (N_19791,N_18769,N_18384);
or U19792 (N_19792,N_18125,N_18215);
xnor U19793 (N_19793,N_18509,N_18654);
xor U19794 (N_19794,N_18806,N_18280);
or U19795 (N_19795,N_18252,N_18216);
nand U19796 (N_19796,N_18617,N_18597);
xnor U19797 (N_19797,N_18469,N_18117);
or U19798 (N_19798,N_18096,N_18638);
nand U19799 (N_19799,N_18170,N_18923);
nor U19800 (N_19800,N_18359,N_19075);
nor U19801 (N_19801,N_18972,N_18968);
nor U19802 (N_19802,N_18819,N_18633);
nand U19803 (N_19803,N_18123,N_18593);
and U19804 (N_19804,N_18870,N_18891);
nand U19805 (N_19805,N_18514,N_19033);
nor U19806 (N_19806,N_18671,N_18829);
nor U19807 (N_19807,N_18549,N_18300);
nor U19808 (N_19808,N_18536,N_18823);
nor U19809 (N_19809,N_18018,N_18861);
nor U19810 (N_19810,N_18498,N_19159);
or U19811 (N_19811,N_18103,N_18567);
nor U19812 (N_19812,N_18486,N_18336);
xnor U19813 (N_19813,N_18269,N_18843);
or U19814 (N_19814,N_18166,N_19159);
nor U19815 (N_19815,N_18314,N_18219);
nor U19816 (N_19816,N_18927,N_18296);
and U19817 (N_19817,N_18622,N_18903);
nand U19818 (N_19818,N_18986,N_18063);
or U19819 (N_19819,N_18586,N_18869);
xor U19820 (N_19820,N_18038,N_18606);
or U19821 (N_19821,N_18662,N_18877);
or U19822 (N_19822,N_18821,N_18080);
nor U19823 (N_19823,N_18668,N_18020);
nand U19824 (N_19824,N_18290,N_19187);
xor U19825 (N_19825,N_18428,N_19015);
and U19826 (N_19826,N_18075,N_18169);
nor U19827 (N_19827,N_18654,N_18397);
xnor U19828 (N_19828,N_18819,N_18731);
nor U19829 (N_19829,N_18278,N_18891);
nor U19830 (N_19830,N_19110,N_18610);
nand U19831 (N_19831,N_18978,N_18372);
and U19832 (N_19832,N_18648,N_18996);
and U19833 (N_19833,N_18344,N_18030);
xnor U19834 (N_19834,N_18630,N_19163);
xnor U19835 (N_19835,N_18601,N_18775);
nand U19836 (N_19836,N_19155,N_18785);
and U19837 (N_19837,N_18394,N_18525);
or U19838 (N_19838,N_18447,N_18441);
or U19839 (N_19839,N_18304,N_18949);
and U19840 (N_19840,N_18202,N_18355);
xor U19841 (N_19841,N_18973,N_18822);
xor U19842 (N_19842,N_18990,N_18306);
nand U19843 (N_19843,N_18606,N_19134);
nor U19844 (N_19844,N_19111,N_18812);
nand U19845 (N_19845,N_19132,N_18331);
xor U19846 (N_19846,N_19011,N_18417);
nor U19847 (N_19847,N_19007,N_19067);
nand U19848 (N_19848,N_18780,N_19186);
or U19849 (N_19849,N_18101,N_18594);
nor U19850 (N_19850,N_18116,N_18989);
or U19851 (N_19851,N_18568,N_18138);
nor U19852 (N_19852,N_18572,N_19138);
nand U19853 (N_19853,N_19188,N_18246);
or U19854 (N_19854,N_18885,N_18108);
or U19855 (N_19855,N_18296,N_19101);
nand U19856 (N_19856,N_19074,N_19166);
nand U19857 (N_19857,N_18633,N_18078);
xnor U19858 (N_19858,N_18288,N_18639);
nor U19859 (N_19859,N_18293,N_18549);
xor U19860 (N_19860,N_18414,N_18392);
xor U19861 (N_19861,N_18761,N_19130);
nor U19862 (N_19862,N_18337,N_18255);
nand U19863 (N_19863,N_18074,N_18403);
nand U19864 (N_19864,N_18787,N_19004);
nand U19865 (N_19865,N_19025,N_18254);
and U19866 (N_19866,N_18503,N_18991);
nor U19867 (N_19867,N_18816,N_18315);
nand U19868 (N_19868,N_19197,N_18883);
nor U19869 (N_19869,N_18150,N_18762);
xor U19870 (N_19870,N_18626,N_18326);
nor U19871 (N_19871,N_19144,N_19082);
or U19872 (N_19872,N_18984,N_19021);
and U19873 (N_19873,N_18562,N_18464);
xnor U19874 (N_19874,N_18962,N_19042);
nor U19875 (N_19875,N_18197,N_18974);
xnor U19876 (N_19876,N_19145,N_18587);
nand U19877 (N_19877,N_18695,N_18093);
and U19878 (N_19878,N_18867,N_18114);
xnor U19879 (N_19879,N_18911,N_18295);
nand U19880 (N_19880,N_18652,N_18639);
nand U19881 (N_19881,N_18521,N_18408);
or U19882 (N_19882,N_18116,N_18317);
nor U19883 (N_19883,N_18913,N_19184);
and U19884 (N_19884,N_18630,N_18880);
nor U19885 (N_19885,N_18438,N_18332);
xor U19886 (N_19886,N_18250,N_18505);
xnor U19887 (N_19887,N_18533,N_18138);
nor U19888 (N_19888,N_18032,N_18776);
nand U19889 (N_19889,N_18421,N_18466);
xnor U19890 (N_19890,N_18987,N_19067);
xnor U19891 (N_19891,N_19159,N_18819);
or U19892 (N_19892,N_19040,N_18809);
xor U19893 (N_19893,N_18528,N_18854);
xor U19894 (N_19894,N_18450,N_18347);
xnor U19895 (N_19895,N_18122,N_18325);
nand U19896 (N_19896,N_18176,N_18224);
or U19897 (N_19897,N_18798,N_19039);
xor U19898 (N_19898,N_18335,N_18738);
nor U19899 (N_19899,N_18007,N_18415);
and U19900 (N_19900,N_18735,N_18443);
nor U19901 (N_19901,N_18668,N_18191);
and U19902 (N_19902,N_18266,N_18621);
or U19903 (N_19903,N_18331,N_18434);
nor U19904 (N_19904,N_18775,N_18567);
nand U19905 (N_19905,N_18868,N_18657);
xnor U19906 (N_19906,N_18510,N_18150);
nor U19907 (N_19907,N_19048,N_19180);
xor U19908 (N_19908,N_18645,N_18938);
nor U19909 (N_19909,N_19111,N_18892);
xnor U19910 (N_19910,N_18756,N_18124);
or U19911 (N_19911,N_18579,N_18656);
or U19912 (N_19912,N_18714,N_18565);
and U19913 (N_19913,N_18961,N_18325);
and U19914 (N_19914,N_18099,N_18520);
nor U19915 (N_19915,N_18142,N_18127);
nand U19916 (N_19916,N_18527,N_19008);
or U19917 (N_19917,N_19136,N_18761);
nor U19918 (N_19918,N_18937,N_18265);
xor U19919 (N_19919,N_18819,N_18746);
nor U19920 (N_19920,N_18269,N_18530);
and U19921 (N_19921,N_18596,N_18198);
nor U19922 (N_19922,N_18351,N_18840);
or U19923 (N_19923,N_18265,N_19029);
and U19924 (N_19924,N_18138,N_18932);
xor U19925 (N_19925,N_18193,N_18115);
and U19926 (N_19926,N_18891,N_18242);
or U19927 (N_19927,N_18083,N_18642);
and U19928 (N_19928,N_18485,N_18327);
or U19929 (N_19929,N_19103,N_18500);
nor U19930 (N_19930,N_19057,N_18758);
or U19931 (N_19931,N_18313,N_19060);
nand U19932 (N_19932,N_18393,N_19140);
nor U19933 (N_19933,N_18607,N_18716);
xor U19934 (N_19934,N_18202,N_18418);
nand U19935 (N_19935,N_18367,N_18878);
nor U19936 (N_19936,N_18029,N_18757);
and U19937 (N_19937,N_18738,N_18140);
or U19938 (N_19938,N_18661,N_18867);
and U19939 (N_19939,N_18986,N_18152);
xnor U19940 (N_19940,N_18169,N_18293);
or U19941 (N_19941,N_18188,N_18786);
nor U19942 (N_19942,N_18205,N_18924);
and U19943 (N_19943,N_18145,N_18848);
nor U19944 (N_19944,N_18846,N_18696);
xnor U19945 (N_19945,N_18733,N_18893);
xnor U19946 (N_19946,N_18844,N_18379);
nor U19947 (N_19947,N_18572,N_19006);
xnor U19948 (N_19948,N_18637,N_18016);
or U19949 (N_19949,N_18141,N_18770);
xor U19950 (N_19950,N_18889,N_18846);
nor U19951 (N_19951,N_18156,N_18045);
and U19952 (N_19952,N_18212,N_18180);
nor U19953 (N_19953,N_18702,N_18094);
nor U19954 (N_19954,N_19034,N_18009);
and U19955 (N_19955,N_19185,N_18777);
or U19956 (N_19956,N_18292,N_18481);
nor U19957 (N_19957,N_18227,N_18105);
and U19958 (N_19958,N_19174,N_18182);
xor U19959 (N_19959,N_18817,N_18429);
and U19960 (N_19960,N_18108,N_18271);
and U19961 (N_19961,N_19020,N_18293);
xor U19962 (N_19962,N_18825,N_18188);
nand U19963 (N_19963,N_18709,N_18620);
and U19964 (N_19964,N_18880,N_18089);
xnor U19965 (N_19965,N_18019,N_18642);
xor U19966 (N_19966,N_18557,N_18507);
or U19967 (N_19967,N_18036,N_19078);
and U19968 (N_19968,N_18459,N_18715);
xnor U19969 (N_19969,N_19137,N_18709);
xnor U19970 (N_19970,N_18933,N_18448);
nor U19971 (N_19971,N_18178,N_18276);
xnor U19972 (N_19972,N_18537,N_18944);
xor U19973 (N_19973,N_18968,N_18639);
nand U19974 (N_19974,N_18294,N_18632);
nor U19975 (N_19975,N_18604,N_18389);
or U19976 (N_19976,N_18229,N_18368);
nor U19977 (N_19977,N_18916,N_18827);
xnor U19978 (N_19978,N_18045,N_18241);
nand U19979 (N_19979,N_18062,N_18942);
nand U19980 (N_19980,N_18339,N_18638);
and U19981 (N_19981,N_18338,N_18415);
or U19982 (N_19982,N_18370,N_18544);
and U19983 (N_19983,N_19150,N_18998);
and U19984 (N_19984,N_18110,N_18243);
nor U19985 (N_19985,N_18326,N_18450);
nand U19986 (N_19986,N_18561,N_19035);
and U19987 (N_19987,N_18392,N_18489);
xor U19988 (N_19988,N_18846,N_18374);
and U19989 (N_19989,N_19173,N_18768);
nand U19990 (N_19990,N_18400,N_19084);
or U19991 (N_19991,N_18500,N_18746);
and U19992 (N_19992,N_18838,N_18534);
nor U19993 (N_19993,N_18692,N_18319);
xnor U19994 (N_19994,N_18715,N_18404);
xor U19995 (N_19995,N_19113,N_18514);
nor U19996 (N_19996,N_18043,N_18046);
and U19997 (N_19997,N_18674,N_18546);
nand U19998 (N_19998,N_18966,N_18193);
nor U19999 (N_19999,N_18041,N_18223);
or U20000 (N_20000,N_19127,N_18077);
nand U20001 (N_20001,N_18668,N_18161);
and U20002 (N_20002,N_18594,N_18700);
or U20003 (N_20003,N_19191,N_19127);
xnor U20004 (N_20004,N_18164,N_18812);
nor U20005 (N_20005,N_18491,N_18328);
and U20006 (N_20006,N_19016,N_18655);
or U20007 (N_20007,N_18633,N_18436);
nand U20008 (N_20008,N_18882,N_18649);
xor U20009 (N_20009,N_18548,N_18192);
or U20010 (N_20010,N_18194,N_18034);
and U20011 (N_20011,N_18148,N_18542);
xor U20012 (N_20012,N_18772,N_18800);
or U20013 (N_20013,N_18031,N_18156);
xnor U20014 (N_20014,N_18911,N_18338);
or U20015 (N_20015,N_19161,N_18506);
or U20016 (N_20016,N_19137,N_19079);
xnor U20017 (N_20017,N_19196,N_18783);
and U20018 (N_20018,N_18711,N_18162);
and U20019 (N_20019,N_18232,N_18762);
nand U20020 (N_20020,N_18252,N_18046);
and U20021 (N_20021,N_18528,N_19082);
nor U20022 (N_20022,N_18165,N_19134);
and U20023 (N_20023,N_18957,N_18347);
xnor U20024 (N_20024,N_19151,N_18637);
and U20025 (N_20025,N_18372,N_18609);
and U20026 (N_20026,N_19196,N_18987);
xnor U20027 (N_20027,N_19196,N_18541);
nand U20028 (N_20028,N_18604,N_18988);
or U20029 (N_20029,N_19108,N_18637);
or U20030 (N_20030,N_18813,N_19149);
xnor U20031 (N_20031,N_18145,N_19046);
nand U20032 (N_20032,N_18328,N_18330);
or U20033 (N_20033,N_18787,N_18099);
nand U20034 (N_20034,N_19121,N_18819);
nand U20035 (N_20035,N_18302,N_18269);
or U20036 (N_20036,N_18683,N_18682);
and U20037 (N_20037,N_19179,N_18697);
xnor U20038 (N_20038,N_18051,N_18352);
nand U20039 (N_20039,N_18176,N_19147);
or U20040 (N_20040,N_18268,N_18548);
nand U20041 (N_20041,N_18878,N_18375);
xor U20042 (N_20042,N_19152,N_18764);
or U20043 (N_20043,N_18860,N_19063);
nand U20044 (N_20044,N_18345,N_18178);
nand U20045 (N_20045,N_18322,N_18253);
xnor U20046 (N_20046,N_18987,N_18095);
and U20047 (N_20047,N_18605,N_18492);
and U20048 (N_20048,N_18014,N_18589);
xnor U20049 (N_20049,N_18465,N_18830);
or U20050 (N_20050,N_18287,N_18005);
xor U20051 (N_20051,N_18314,N_18818);
nor U20052 (N_20052,N_18239,N_18328);
nor U20053 (N_20053,N_19004,N_18764);
and U20054 (N_20054,N_18659,N_18070);
xnor U20055 (N_20055,N_18147,N_18062);
and U20056 (N_20056,N_18820,N_18575);
or U20057 (N_20057,N_19039,N_18310);
nor U20058 (N_20058,N_18375,N_18750);
nor U20059 (N_20059,N_18589,N_18669);
or U20060 (N_20060,N_18998,N_19009);
and U20061 (N_20061,N_18657,N_18041);
or U20062 (N_20062,N_18916,N_18127);
nand U20063 (N_20063,N_18450,N_18311);
nand U20064 (N_20064,N_18194,N_19118);
nand U20065 (N_20065,N_18203,N_18670);
nand U20066 (N_20066,N_18247,N_19107);
nor U20067 (N_20067,N_18788,N_18467);
xnor U20068 (N_20068,N_18434,N_18296);
and U20069 (N_20069,N_18219,N_18012);
and U20070 (N_20070,N_18645,N_19069);
and U20071 (N_20071,N_19044,N_18277);
nor U20072 (N_20072,N_18080,N_19115);
or U20073 (N_20073,N_18328,N_18243);
nand U20074 (N_20074,N_18534,N_19124);
nor U20075 (N_20075,N_18619,N_18046);
xor U20076 (N_20076,N_18093,N_19050);
nand U20077 (N_20077,N_18522,N_18423);
and U20078 (N_20078,N_18526,N_18400);
xnor U20079 (N_20079,N_18888,N_18167);
nor U20080 (N_20080,N_18286,N_19167);
xor U20081 (N_20081,N_18749,N_18757);
or U20082 (N_20082,N_19149,N_18149);
and U20083 (N_20083,N_18537,N_19151);
nor U20084 (N_20084,N_18220,N_18954);
nand U20085 (N_20085,N_18795,N_18685);
nor U20086 (N_20086,N_18158,N_18086);
and U20087 (N_20087,N_18733,N_18646);
nor U20088 (N_20088,N_18298,N_18682);
and U20089 (N_20089,N_18623,N_18408);
xor U20090 (N_20090,N_18958,N_18206);
or U20091 (N_20091,N_18165,N_19082);
xor U20092 (N_20092,N_18820,N_18147);
xor U20093 (N_20093,N_18360,N_18794);
xor U20094 (N_20094,N_18329,N_19173);
and U20095 (N_20095,N_18408,N_18149);
and U20096 (N_20096,N_18440,N_19029);
or U20097 (N_20097,N_19130,N_19069);
nor U20098 (N_20098,N_19016,N_18679);
and U20099 (N_20099,N_19161,N_18232);
xor U20100 (N_20100,N_18365,N_18545);
or U20101 (N_20101,N_18569,N_18456);
or U20102 (N_20102,N_19138,N_18928);
xnor U20103 (N_20103,N_19134,N_18596);
xnor U20104 (N_20104,N_18276,N_18835);
and U20105 (N_20105,N_18336,N_18836);
and U20106 (N_20106,N_18357,N_19121);
or U20107 (N_20107,N_18042,N_18184);
or U20108 (N_20108,N_18178,N_18794);
nor U20109 (N_20109,N_18586,N_18949);
or U20110 (N_20110,N_18641,N_18999);
nand U20111 (N_20111,N_19172,N_18179);
nand U20112 (N_20112,N_19056,N_18301);
nor U20113 (N_20113,N_18131,N_19148);
and U20114 (N_20114,N_18169,N_18532);
nor U20115 (N_20115,N_18620,N_18009);
xor U20116 (N_20116,N_18584,N_18563);
and U20117 (N_20117,N_18450,N_18860);
nor U20118 (N_20118,N_18175,N_18733);
or U20119 (N_20119,N_18369,N_19051);
or U20120 (N_20120,N_18525,N_18820);
nor U20121 (N_20121,N_18431,N_18621);
and U20122 (N_20122,N_18281,N_18196);
xnor U20123 (N_20123,N_18152,N_19155);
or U20124 (N_20124,N_18893,N_18912);
nor U20125 (N_20125,N_18055,N_18783);
and U20126 (N_20126,N_19061,N_19000);
or U20127 (N_20127,N_18194,N_18025);
and U20128 (N_20128,N_18736,N_18875);
xnor U20129 (N_20129,N_18674,N_18757);
nand U20130 (N_20130,N_18036,N_18506);
nand U20131 (N_20131,N_18179,N_18457);
or U20132 (N_20132,N_18494,N_19078);
nand U20133 (N_20133,N_18323,N_19182);
or U20134 (N_20134,N_18676,N_19064);
nor U20135 (N_20135,N_19198,N_18815);
and U20136 (N_20136,N_18837,N_18389);
and U20137 (N_20137,N_18605,N_18445);
or U20138 (N_20138,N_18405,N_19166);
or U20139 (N_20139,N_18309,N_18826);
or U20140 (N_20140,N_19044,N_18918);
nor U20141 (N_20141,N_18826,N_18418);
or U20142 (N_20142,N_18758,N_18522);
or U20143 (N_20143,N_19151,N_19080);
and U20144 (N_20144,N_18390,N_18380);
nor U20145 (N_20145,N_18594,N_18538);
xor U20146 (N_20146,N_18757,N_18454);
nor U20147 (N_20147,N_19022,N_18021);
xor U20148 (N_20148,N_18540,N_18525);
xnor U20149 (N_20149,N_18448,N_18979);
or U20150 (N_20150,N_18421,N_19041);
nand U20151 (N_20151,N_18647,N_18652);
or U20152 (N_20152,N_18584,N_18678);
xnor U20153 (N_20153,N_18575,N_18883);
or U20154 (N_20154,N_18589,N_18181);
xnor U20155 (N_20155,N_18373,N_18969);
xor U20156 (N_20156,N_18573,N_18878);
nor U20157 (N_20157,N_19111,N_18322);
nor U20158 (N_20158,N_18754,N_18870);
nand U20159 (N_20159,N_18826,N_19081);
nor U20160 (N_20160,N_18946,N_19092);
nor U20161 (N_20161,N_18104,N_18331);
or U20162 (N_20162,N_18680,N_18737);
nor U20163 (N_20163,N_18121,N_18749);
nor U20164 (N_20164,N_18984,N_18353);
and U20165 (N_20165,N_18007,N_18936);
nor U20166 (N_20166,N_18340,N_18640);
nor U20167 (N_20167,N_18145,N_18750);
nand U20168 (N_20168,N_18158,N_18888);
nor U20169 (N_20169,N_18838,N_18482);
nand U20170 (N_20170,N_18667,N_18264);
xor U20171 (N_20171,N_18805,N_18342);
nand U20172 (N_20172,N_18250,N_18878);
or U20173 (N_20173,N_18795,N_18673);
nor U20174 (N_20174,N_18453,N_18348);
and U20175 (N_20175,N_19147,N_18114);
nand U20176 (N_20176,N_18502,N_18520);
and U20177 (N_20177,N_18903,N_18942);
xor U20178 (N_20178,N_18652,N_18324);
nor U20179 (N_20179,N_18082,N_18095);
nand U20180 (N_20180,N_18717,N_19155);
nor U20181 (N_20181,N_18298,N_18189);
xnor U20182 (N_20182,N_19005,N_18281);
and U20183 (N_20183,N_18980,N_18911);
and U20184 (N_20184,N_18955,N_18942);
nand U20185 (N_20185,N_18689,N_18525);
and U20186 (N_20186,N_18985,N_19102);
xnor U20187 (N_20187,N_18982,N_18585);
nor U20188 (N_20188,N_18646,N_18660);
or U20189 (N_20189,N_18942,N_18568);
nor U20190 (N_20190,N_18410,N_18094);
nor U20191 (N_20191,N_18780,N_18034);
nand U20192 (N_20192,N_18728,N_18974);
xor U20193 (N_20193,N_18738,N_18890);
nand U20194 (N_20194,N_18902,N_18525);
or U20195 (N_20195,N_18743,N_18541);
and U20196 (N_20196,N_18855,N_18847);
xnor U20197 (N_20197,N_18725,N_18540);
or U20198 (N_20198,N_19199,N_18842);
nand U20199 (N_20199,N_18399,N_19124);
nor U20200 (N_20200,N_19035,N_18704);
and U20201 (N_20201,N_18823,N_18715);
and U20202 (N_20202,N_18035,N_19103);
nand U20203 (N_20203,N_18826,N_18234);
nand U20204 (N_20204,N_19159,N_19057);
nand U20205 (N_20205,N_18301,N_18695);
nand U20206 (N_20206,N_18449,N_18595);
nand U20207 (N_20207,N_18773,N_18410);
or U20208 (N_20208,N_18701,N_18224);
nand U20209 (N_20209,N_19158,N_18804);
or U20210 (N_20210,N_18813,N_18239);
nor U20211 (N_20211,N_19025,N_18472);
or U20212 (N_20212,N_18559,N_18572);
and U20213 (N_20213,N_19140,N_18577);
and U20214 (N_20214,N_18055,N_18190);
nand U20215 (N_20215,N_18483,N_18094);
xor U20216 (N_20216,N_18808,N_18255);
or U20217 (N_20217,N_18519,N_18586);
xor U20218 (N_20218,N_18972,N_18910);
xor U20219 (N_20219,N_18605,N_18239);
or U20220 (N_20220,N_18054,N_18564);
xor U20221 (N_20221,N_18817,N_18464);
and U20222 (N_20222,N_18757,N_18873);
nor U20223 (N_20223,N_18530,N_18957);
or U20224 (N_20224,N_19001,N_18404);
and U20225 (N_20225,N_18392,N_19051);
nor U20226 (N_20226,N_18908,N_18851);
xnor U20227 (N_20227,N_18233,N_18750);
or U20228 (N_20228,N_18008,N_19057);
and U20229 (N_20229,N_18788,N_19028);
nand U20230 (N_20230,N_19073,N_18084);
nor U20231 (N_20231,N_18417,N_19196);
xnor U20232 (N_20232,N_19138,N_18805);
and U20233 (N_20233,N_19180,N_18620);
or U20234 (N_20234,N_18607,N_19031);
xor U20235 (N_20235,N_18028,N_19139);
nor U20236 (N_20236,N_19170,N_18838);
or U20237 (N_20237,N_18215,N_18475);
or U20238 (N_20238,N_18633,N_18014);
or U20239 (N_20239,N_18740,N_18149);
nor U20240 (N_20240,N_18461,N_18427);
nand U20241 (N_20241,N_18606,N_19120);
and U20242 (N_20242,N_18530,N_18366);
xor U20243 (N_20243,N_18103,N_18584);
and U20244 (N_20244,N_18024,N_18734);
nand U20245 (N_20245,N_18604,N_18241);
nor U20246 (N_20246,N_19084,N_18311);
xnor U20247 (N_20247,N_18793,N_18224);
nor U20248 (N_20248,N_18623,N_19000);
or U20249 (N_20249,N_18200,N_18209);
nor U20250 (N_20250,N_18770,N_18436);
xor U20251 (N_20251,N_19072,N_18256);
and U20252 (N_20252,N_18747,N_18472);
and U20253 (N_20253,N_18219,N_18691);
nand U20254 (N_20254,N_18849,N_18987);
nand U20255 (N_20255,N_19020,N_18889);
nand U20256 (N_20256,N_19166,N_18444);
nor U20257 (N_20257,N_18040,N_18424);
xnor U20258 (N_20258,N_19138,N_19022);
xor U20259 (N_20259,N_18943,N_18375);
nand U20260 (N_20260,N_18304,N_18849);
or U20261 (N_20261,N_18180,N_18730);
nand U20262 (N_20262,N_19125,N_18687);
nor U20263 (N_20263,N_18182,N_18115);
nor U20264 (N_20264,N_18528,N_18111);
or U20265 (N_20265,N_18036,N_18405);
nand U20266 (N_20266,N_19064,N_18876);
or U20267 (N_20267,N_18530,N_18759);
nand U20268 (N_20268,N_18243,N_18570);
and U20269 (N_20269,N_18030,N_18913);
and U20270 (N_20270,N_19029,N_19129);
or U20271 (N_20271,N_18200,N_18625);
xor U20272 (N_20272,N_18339,N_18808);
nand U20273 (N_20273,N_18567,N_19144);
nand U20274 (N_20274,N_18806,N_18300);
xor U20275 (N_20275,N_18802,N_18714);
nand U20276 (N_20276,N_18069,N_18013);
xnor U20277 (N_20277,N_18806,N_18421);
nor U20278 (N_20278,N_18429,N_18920);
nor U20279 (N_20279,N_19035,N_19069);
or U20280 (N_20280,N_18340,N_19104);
or U20281 (N_20281,N_18639,N_18287);
nand U20282 (N_20282,N_18491,N_18111);
nor U20283 (N_20283,N_18955,N_18821);
xnor U20284 (N_20284,N_18090,N_18918);
and U20285 (N_20285,N_19105,N_19081);
and U20286 (N_20286,N_18215,N_18556);
nand U20287 (N_20287,N_19128,N_18368);
xnor U20288 (N_20288,N_18062,N_18651);
and U20289 (N_20289,N_18251,N_18679);
nor U20290 (N_20290,N_18299,N_18804);
nor U20291 (N_20291,N_18741,N_19004);
nand U20292 (N_20292,N_18215,N_18484);
xor U20293 (N_20293,N_18927,N_18566);
nor U20294 (N_20294,N_18822,N_18729);
nand U20295 (N_20295,N_18479,N_18604);
nor U20296 (N_20296,N_18319,N_18991);
nand U20297 (N_20297,N_18770,N_19054);
and U20298 (N_20298,N_19111,N_18917);
nand U20299 (N_20299,N_18218,N_19137);
nor U20300 (N_20300,N_18206,N_18865);
and U20301 (N_20301,N_18483,N_18008);
and U20302 (N_20302,N_18461,N_18552);
xor U20303 (N_20303,N_19107,N_18442);
nor U20304 (N_20304,N_18866,N_18214);
and U20305 (N_20305,N_18222,N_19001);
nand U20306 (N_20306,N_19055,N_18845);
nor U20307 (N_20307,N_18413,N_18231);
and U20308 (N_20308,N_18452,N_18157);
nor U20309 (N_20309,N_18253,N_18398);
xnor U20310 (N_20310,N_19010,N_18392);
nand U20311 (N_20311,N_18788,N_18852);
nor U20312 (N_20312,N_18452,N_19076);
nor U20313 (N_20313,N_18498,N_18816);
and U20314 (N_20314,N_18388,N_18605);
xor U20315 (N_20315,N_18576,N_18975);
nor U20316 (N_20316,N_18617,N_18899);
nand U20317 (N_20317,N_18891,N_19072);
nand U20318 (N_20318,N_18568,N_18413);
nor U20319 (N_20319,N_19180,N_19027);
nand U20320 (N_20320,N_18825,N_18870);
nor U20321 (N_20321,N_18721,N_19002);
nand U20322 (N_20322,N_18866,N_18496);
nand U20323 (N_20323,N_18790,N_18529);
and U20324 (N_20324,N_19130,N_19029);
xor U20325 (N_20325,N_18138,N_18151);
nor U20326 (N_20326,N_18844,N_18111);
nor U20327 (N_20327,N_18595,N_18707);
nand U20328 (N_20328,N_18464,N_18720);
nor U20329 (N_20329,N_18324,N_18863);
nand U20330 (N_20330,N_18575,N_18767);
nand U20331 (N_20331,N_18419,N_18347);
nor U20332 (N_20332,N_18222,N_19095);
nand U20333 (N_20333,N_18627,N_18525);
xor U20334 (N_20334,N_18716,N_18916);
xnor U20335 (N_20335,N_18728,N_18802);
nor U20336 (N_20336,N_18272,N_19175);
and U20337 (N_20337,N_18075,N_18601);
or U20338 (N_20338,N_18095,N_18274);
and U20339 (N_20339,N_18390,N_18967);
nor U20340 (N_20340,N_18284,N_18765);
nand U20341 (N_20341,N_18274,N_18464);
nand U20342 (N_20342,N_18768,N_18555);
xor U20343 (N_20343,N_18972,N_18391);
and U20344 (N_20344,N_18161,N_18438);
nor U20345 (N_20345,N_19092,N_18176);
or U20346 (N_20346,N_18492,N_18871);
xnor U20347 (N_20347,N_19076,N_18966);
xor U20348 (N_20348,N_18365,N_18638);
nand U20349 (N_20349,N_18228,N_18762);
and U20350 (N_20350,N_18780,N_18091);
and U20351 (N_20351,N_18786,N_18587);
or U20352 (N_20352,N_18829,N_18541);
nand U20353 (N_20353,N_18371,N_18742);
xnor U20354 (N_20354,N_18850,N_18525);
xor U20355 (N_20355,N_18314,N_18061);
or U20356 (N_20356,N_19183,N_18655);
or U20357 (N_20357,N_18071,N_18178);
or U20358 (N_20358,N_19063,N_18856);
and U20359 (N_20359,N_18723,N_18385);
xor U20360 (N_20360,N_18290,N_18757);
nand U20361 (N_20361,N_18352,N_18095);
and U20362 (N_20362,N_18099,N_18730);
xnor U20363 (N_20363,N_18463,N_18106);
or U20364 (N_20364,N_18746,N_18497);
or U20365 (N_20365,N_18061,N_18741);
nand U20366 (N_20366,N_18141,N_18111);
xnor U20367 (N_20367,N_18218,N_18554);
nand U20368 (N_20368,N_19099,N_19048);
or U20369 (N_20369,N_18564,N_18728);
nand U20370 (N_20370,N_18915,N_18105);
xor U20371 (N_20371,N_18559,N_18001);
and U20372 (N_20372,N_19188,N_19094);
xor U20373 (N_20373,N_18688,N_19119);
or U20374 (N_20374,N_18969,N_18799);
nor U20375 (N_20375,N_18540,N_18634);
nand U20376 (N_20376,N_18780,N_18741);
nor U20377 (N_20377,N_18754,N_18433);
nand U20378 (N_20378,N_18773,N_18252);
xnor U20379 (N_20379,N_18776,N_18262);
and U20380 (N_20380,N_18862,N_18069);
and U20381 (N_20381,N_19016,N_18268);
nor U20382 (N_20382,N_18552,N_18192);
and U20383 (N_20383,N_18120,N_18850);
nor U20384 (N_20384,N_19088,N_18484);
xnor U20385 (N_20385,N_18512,N_18696);
and U20386 (N_20386,N_18310,N_18732);
nand U20387 (N_20387,N_18478,N_19088);
nand U20388 (N_20388,N_18264,N_18779);
nor U20389 (N_20389,N_18640,N_18721);
and U20390 (N_20390,N_18602,N_18658);
xor U20391 (N_20391,N_18672,N_18384);
nand U20392 (N_20392,N_18707,N_18810);
nor U20393 (N_20393,N_18316,N_19131);
xor U20394 (N_20394,N_18603,N_18874);
xnor U20395 (N_20395,N_18155,N_18995);
xor U20396 (N_20396,N_19121,N_18385);
or U20397 (N_20397,N_18594,N_18444);
xnor U20398 (N_20398,N_18304,N_18393);
and U20399 (N_20399,N_19118,N_18475);
nor U20400 (N_20400,N_19880,N_19670);
and U20401 (N_20401,N_19340,N_19626);
nand U20402 (N_20402,N_19360,N_19290);
xor U20403 (N_20403,N_20221,N_20259);
or U20404 (N_20404,N_19500,N_19968);
and U20405 (N_20405,N_19210,N_20143);
and U20406 (N_20406,N_19533,N_19767);
or U20407 (N_20407,N_19708,N_19939);
nand U20408 (N_20408,N_19996,N_19748);
xnor U20409 (N_20409,N_19927,N_19788);
xor U20410 (N_20410,N_20008,N_20305);
or U20411 (N_20411,N_19833,N_20041);
nand U20412 (N_20412,N_20165,N_20346);
xor U20413 (N_20413,N_19321,N_19588);
nand U20414 (N_20414,N_20397,N_19826);
or U20415 (N_20415,N_19717,N_20246);
or U20416 (N_20416,N_20016,N_19505);
and U20417 (N_20417,N_19575,N_20327);
xnor U20418 (N_20418,N_19657,N_19359);
nand U20419 (N_20419,N_19655,N_19902);
xor U20420 (N_20420,N_20058,N_19416);
or U20421 (N_20421,N_19664,N_19761);
or U20422 (N_20422,N_19335,N_19525);
and U20423 (N_20423,N_20337,N_20192);
nor U20424 (N_20424,N_20319,N_19355);
nand U20425 (N_20425,N_20236,N_19794);
xor U20426 (N_20426,N_20168,N_19994);
nor U20427 (N_20427,N_20055,N_19770);
xor U20428 (N_20428,N_19837,N_19244);
or U20429 (N_20429,N_19909,N_19564);
nor U20430 (N_20430,N_19225,N_20219);
or U20431 (N_20431,N_19487,N_20301);
nor U20432 (N_20432,N_19771,N_19822);
nor U20433 (N_20433,N_19637,N_19718);
nand U20434 (N_20434,N_20380,N_20211);
nand U20435 (N_20435,N_19255,N_20359);
nand U20436 (N_20436,N_19705,N_20112);
or U20437 (N_20437,N_19901,N_19323);
nor U20438 (N_20438,N_19916,N_19236);
xnor U20439 (N_20439,N_20132,N_20089);
and U20440 (N_20440,N_19773,N_19920);
and U20441 (N_20441,N_19517,N_19452);
nor U20442 (N_20442,N_20318,N_20097);
xor U20443 (N_20443,N_19246,N_19636);
and U20444 (N_20444,N_19490,N_19519);
and U20445 (N_20445,N_19904,N_20258);
and U20446 (N_20446,N_19877,N_20224);
and U20447 (N_20447,N_20169,N_19775);
nor U20448 (N_20448,N_20103,N_19923);
or U20449 (N_20449,N_19552,N_20051);
xor U20450 (N_20450,N_20060,N_19324);
nand U20451 (N_20451,N_20201,N_19211);
xor U20452 (N_20452,N_19958,N_20090);
nand U20453 (N_20453,N_19507,N_19991);
nor U20454 (N_20454,N_20394,N_19677);
or U20455 (N_20455,N_19806,N_20033);
or U20456 (N_20456,N_19689,N_19566);
nor U20457 (N_20457,N_20212,N_19387);
and U20458 (N_20458,N_20226,N_19337);
xor U20459 (N_20459,N_19855,N_19441);
or U20460 (N_20460,N_19493,N_19783);
xnor U20461 (N_20461,N_19478,N_20199);
or U20462 (N_20462,N_19873,N_19724);
nor U20463 (N_20463,N_19528,N_19814);
or U20464 (N_20464,N_20094,N_19680);
or U20465 (N_20465,N_19804,N_19266);
or U20466 (N_20466,N_20216,N_20036);
xor U20467 (N_20467,N_19895,N_19394);
nor U20468 (N_20468,N_19252,N_19456);
nand U20469 (N_20469,N_19473,N_19673);
xor U20470 (N_20470,N_20227,N_20292);
xnor U20471 (N_20471,N_19404,N_20367);
xor U20472 (N_20472,N_19903,N_20390);
nor U20473 (N_20473,N_20282,N_20023);
xnor U20474 (N_20474,N_20306,N_19737);
nor U20475 (N_20475,N_19922,N_19330);
and U20476 (N_20476,N_20348,N_19819);
nand U20477 (N_20477,N_19848,N_19972);
xor U20478 (N_20478,N_19897,N_20369);
nand U20479 (N_20479,N_20204,N_20198);
nor U20480 (N_20480,N_20277,N_19662);
nand U20481 (N_20481,N_19408,N_19406);
xor U20482 (N_20482,N_20045,N_20148);
and U20483 (N_20483,N_19397,N_19437);
or U20484 (N_20484,N_20106,N_20159);
xnor U20485 (N_20485,N_19440,N_20077);
or U20486 (N_20486,N_19450,N_20080);
nand U20487 (N_20487,N_20338,N_19774);
or U20488 (N_20488,N_20311,N_19691);
xor U20489 (N_20489,N_20186,N_19302);
nand U20490 (N_20490,N_19369,N_19600);
nand U20491 (N_20491,N_19562,N_19429);
and U20492 (N_20492,N_19975,N_20015);
and U20493 (N_20493,N_19784,N_19345);
nand U20494 (N_20494,N_20190,N_19545);
or U20495 (N_20495,N_20009,N_19215);
and U20496 (N_20496,N_19870,N_19257);
nand U20497 (N_20497,N_19858,N_19486);
and U20498 (N_20498,N_19216,N_20158);
nor U20499 (N_20499,N_19988,N_19831);
and U20500 (N_20500,N_20088,N_19872);
or U20501 (N_20501,N_19803,N_19596);
xor U20502 (N_20502,N_19746,N_20021);
or U20503 (N_20503,N_19300,N_19735);
or U20504 (N_20504,N_19849,N_19288);
xnor U20505 (N_20505,N_20303,N_19931);
or U20506 (N_20506,N_19581,N_19924);
and U20507 (N_20507,N_19845,N_19489);
nand U20508 (N_20508,N_19363,N_20296);
nand U20509 (N_20509,N_19523,N_19982);
and U20510 (N_20510,N_19801,N_20142);
nand U20511 (N_20511,N_19366,N_19889);
xnor U20512 (N_20512,N_19424,N_19379);
and U20513 (N_20513,N_20032,N_19319);
nor U20514 (N_20514,N_19462,N_19373);
and U20515 (N_20515,N_19910,N_19498);
nand U20516 (N_20516,N_19659,N_19568);
xnor U20517 (N_20517,N_19905,N_19827);
nor U20518 (N_20518,N_20161,N_19692);
nand U20519 (N_20519,N_19232,N_19892);
nor U20520 (N_20520,N_19740,N_20269);
nand U20521 (N_20521,N_20357,N_19840);
nand U20522 (N_20522,N_19479,N_19222);
xor U20523 (N_20523,N_19650,N_20107);
nor U20524 (N_20524,N_19956,N_19812);
nand U20525 (N_20525,N_19307,N_20095);
nor U20526 (N_20526,N_20257,N_19630);
nand U20527 (N_20527,N_19207,N_20233);
or U20528 (N_20528,N_19987,N_19412);
xor U20529 (N_20529,N_19457,N_19698);
xnor U20530 (N_20530,N_19325,N_20196);
and U20531 (N_20531,N_20262,N_20061);
or U20532 (N_20532,N_19926,N_20131);
nor U20533 (N_20533,N_19890,N_19550);
and U20534 (N_20534,N_19728,N_19654);
or U20535 (N_20535,N_19696,N_20118);
xnor U20536 (N_20536,N_20068,N_20162);
nand U20537 (N_20537,N_19648,N_19729);
xor U20538 (N_20538,N_19966,N_20184);
or U20539 (N_20539,N_19209,N_20149);
and U20540 (N_20540,N_19296,N_20175);
nand U20541 (N_20541,N_19713,N_19242);
or U20542 (N_20542,N_20027,N_19953);
nor U20543 (N_20543,N_19417,N_20345);
or U20544 (N_20544,N_20284,N_19834);
nand U20545 (N_20545,N_19221,N_19974);
and U20546 (N_20546,N_19825,N_20194);
nor U20547 (N_20547,N_19738,N_20232);
and U20548 (N_20548,N_20302,N_19992);
nand U20549 (N_20549,N_19886,N_19237);
and U20550 (N_20550,N_19269,N_20119);
xnor U20551 (N_20551,N_19248,N_19538);
or U20552 (N_20552,N_19732,N_19272);
nor U20553 (N_20553,N_20341,N_19639);
xor U20554 (N_20554,N_20156,N_20377);
or U20555 (N_20555,N_19426,N_19442);
or U20556 (N_20556,N_19863,N_20247);
and U20557 (N_20557,N_20020,N_19807);
or U20558 (N_20558,N_19374,N_19934);
nor U20559 (N_20559,N_20365,N_19343);
nor U20560 (N_20560,N_19841,N_19835);
nor U20561 (N_20561,N_20351,N_19929);
nand U20562 (N_20562,N_19560,N_20207);
or U20563 (N_20563,N_19380,N_19375);
or U20564 (N_20564,N_19569,N_20109);
and U20565 (N_20565,N_20239,N_19912);
or U20566 (N_20566,N_19331,N_19857);
nand U20567 (N_20567,N_20398,N_19496);
nand U20568 (N_20568,N_19629,N_19584);
or U20569 (N_20569,N_20382,N_19453);
nor U20570 (N_20570,N_19391,N_20343);
or U20571 (N_20571,N_20133,N_19888);
xor U20572 (N_20572,N_19401,N_20039);
nand U20573 (N_20573,N_19304,N_19970);
and U20574 (N_20574,N_20150,N_19219);
nor U20575 (N_20575,N_20388,N_20272);
and U20576 (N_20576,N_19853,N_19671);
or U20577 (N_20577,N_19646,N_19548);
or U20578 (N_20578,N_19764,N_19431);
nand U20579 (N_20579,N_20253,N_19410);
and U20580 (N_20580,N_19805,N_20163);
or U20581 (N_20581,N_19846,N_19781);
and U20582 (N_20582,N_19291,N_19610);
and U20583 (N_20583,N_20197,N_19963);
and U20584 (N_20584,N_20366,N_19942);
nor U20585 (N_20585,N_19995,N_19521);
xor U20586 (N_20586,N_20245,N_20129);
nand U20587 (N_20587,N_19509,N_19513);
nand U20588 (N_20588,N_19710,N_20145);
nand U20589 (N_20589,N_19537,N_19409);
nand U20590 (N_20590,N_19388,N_19235);
nand U20591 (N_20591,N_19264,N_19510);
and U20592 (N_20592,N_19503,N_19682);
nor U20593 (N_20593,N_19567,N_19754);
and U20594 (N_20594,N_20117,N_19420);
xnor U20595 (N_20595,N_20013,N_19859);
nand U20596 (N_20596,N_20048,N_19459);
xnor U20597 (N_20597,N_19400,N_19551);
and U20598 (N_20598,N_20304,N_19802);
and U20599 (N_20599,N_19669,N_19603);
nor U20600 (N_20600,N_19756,N_20123);
xor U20601 (N_20601,N_19516,N_19483);
nand U20602 (N_20602,N_19540,N_20278);
or U20603 (N_20603,N_20038,N_20276);
xor U20604 (N_20604,N_20116,N_19645);
or U20605 (N_20605,N_19351,N_20022);
nand U20606 (N_20606,N_19917,N_19549);
nand U20607 (N_20607,N_20326,N_19721);
or U20608 (N_20608,N_20260,N_19421);
or U20609 (N_20609,N_19475,N_20141);
and U20610 (N_20610,N_20115,N_19263);
xor U20611 (N_20611,N_19494,N_20354);
and U20612 (N_20612,N_19578,N_19425);
nor U20613 (N_20613,N_19285,N_19820);
nand U20614 (N_20614,N_19699,N_20137);
xor U20615 (N_20615,N_19776,N_20283);
nor U20616 (N_20616,N_20057,N_19709);
nor U20617 (N_20617,N_19874,N_19270);
and U20618 (N_20618,N_19249,N_19439);
nor U20619 (N_20619,N_20237,N_20268);
xor U20620 (N_20620,N_19392,N_19606);
xor U20621 (N_20621,N_19476,N_19875);
nand U20622 (N_20622,N_20087,N_20315);
and U20623 (N_20623,N_20099,N_20370);
nand U20624 (N_20624,N_20096,N_19915);
xnor U20625 (N_20625,N_19700,N_20358);
nor U20626 (N_20626,N_19579,N_20071);
and U20627 (N_20627,N_19668,N_19451);
nand U20628 (N_20628,N_19658,N_19900);
or U20629 (N_20629,N_20062,N_19573);
nor U20630 (N_20630,N_19866,N_19468);
nor U20631 (N_20631,N_19435,N_19438);
xnor U20632 (N_20632,N_19836,N_20085);
nand U20633 (N_20633,N_19543,N_19576);
nor U20634 (N_20634,N_20255,N_20130);
and U20635 (N_20635,N_19779,N_19260);
and U20636 (N_20636,N_19287,N_19960);
and U20637 (N_20637,N_20178,N_19697);
xnor U20638 (N_20638,N_19842,N_19719);
nor U20639 (N_20639,N_19217,N_20389);
nor U20640 (N_20640,N_20288,N_19577);
nand U20641 (N_20641,N_19554,N_19368);
nor U20642 (N_20642,N_19484,N_19372);
xnor U20643 (N_20643,N_20384,N_19928);
nand U20644 (N_20644,N_19301,N_19678);
nand U20645 (N_20645,N_20363,N_20004);
or U20646 (N_20646,N_19245,N_19470);
or U20647 (N_20647,N_19349,N_19843);
nand U20648 (N_20648,N_19862,N_19869);
nor U20649 (N_20649,N_19306,N_19907);
xnor U20650 (N_20650,N_19247,N_19883);
nand U20651 (N_20651,N_19649,N_20275);
nand U20652 (N_20652,N_19961,N_20313);
nor U20653 (N_20653,N_20267,N_20353);
nor U20654 (N_20654,N_20355,N_20360);
nor U20655 (N_20655,N_19204,N_19601);
xor U20656 (N_20656,N_20073,N_19633);
nor U20657 (N_20657,N_19641,N_20375);
xnor U20658 (N_20658,N_19485,N_19769);
nand U20659 (N_20659,N_19730,N_19943);
xnor U20660 (N_20660,N_19376,N_20074);
and U20661 (N_20661,N_19635,N_19711);
xnor U20662 (N_20662,N_20254,N_19386);
and U20663 (N_20663,N_19227,N_19497);
xor U20664 (N_20664,N_19282,N_20356);
nor U20665 (N_20665,N_19675,N_20063);
or U20666 (N_20666,N_19524,N_19419);
and U20667 (N_20667,N_19780,N_20378);
xor U20668 (N_20668,N_19334,N_19529);
or U20669 (N_20669,N_19587,N_19981);
and U20670 (N_20670,N_19320,N_19506);
or U20671 (N_20671,N_20105,N_19621);
nor U20672 (N_20672,N_19464,N_19712);
and U20673 (N_20673,N_20287,N_19983);
or U20674 (N_20674,N_19891,N_19449);
nand U20675 (N_20675,N_19213,N_19515);
nor U20676 (N_20676,N_19714,N_20195);
xor U20677 (N_20677,N_19930,N_20081);
nand U20678 (N_20678,N_19220,N_19458);
and U20679 (N_20679,N_19289,N_19684);
or U20680 (N_20680,N_20050,N_20271);
xnor U20681 (N_20681,N_19563,N_19407);
or U20682 (N_20682,N_20134,N_19925);
and U20683 (N_20683,N_19491,N_20135);
xor U20684 (N_20684,N_20188,N_19559);
nand U20685 (N_20685,N_19980,N_20209);
nand U20686 (N_20686,N_20368,N_20342);
xnor U20687 (N_20687,N_19514,N_19534);
and U20688 (N_20688,N_20230,N_20396);
and U20689 (N_20689,N_19203,N_20024);
nand U20690 (N_20690,N_19336,N_20298);
or U20691 (N_20691,N_20312,N_19879);
nor U20692 (N_20692,N_19526,N_19271);
and U20693 (N_20693,N_19949,N_19832);
or U20694 (N_20694,N_20054,N_19793);
or U20695 (N_20695,N_20011,N_19460);
nor U20696 (N_20696,N_19422,N_20249);
nor U20697 (N_20697,N_19597,N_19202);
and U20698 (N_20698,N_20231,N_19572);
xor U20699 (N_20699,N_20079,N_19893);
nand U20700 (N_20700,N_20206,N_19716);
nor U20701 (N_20701,N_20047,N_19950);
or U20702 (N_20702,N_20270,N_19962);
xor U20703 (N_20703,N_20025,N_20160);
nor U20704 (N_20704,N_20279,N_19502);
nor U20705 (N_20705,N_20222,N_19229);
and U20706 (N_20706,N_19999,N_20127);
nand U20707 (N_20707,N_19967,N_19653);
or U20708 (N_20708,N_19839,N_20281);
and U20709 (N_20709,N_19251,N_19495);
xor U20710 (N_20710,N_19815,N_20330);
nand U20711 (N_20711,N_19693,N_19353);
xnor U20712 (N_20712,N_20286,N_19741);
nand U20713 (N_20713,N_19444,N_19383);
xor U20714 (N_20714,N_20264,N_19796);
xor U20715 (N_20715,N_19243,N_19749);
nor U20716 (N_20716,N_20332,N_20002);
or U20717 (N_20717,N_19743,N_19685);
or U20718 (N_20718,N_19472,N_19683);
xor U20719 (N_20719,N_20046,N_19477);
and U20720 (N_20720,N_20387,N_19303);
xnor U20721 (N_20721,N_19955,N_19951);
and U20722 (N_20722,N_20034,N_19230);
xor U20723 (N_20723,N_20078,N_19396);
and U20724 (N_20724,N_19367,N_19241);
nand U20725 (N_20725,N_19763,N_19726);
nand U20726 (N_20726,N_19861,N_19256);
and U20727 (N_20727,N_19782,N_19766);
or U20728 (N_20728,N_19350,N_19667);
xnor U20729 (N_20729,N_20125,N_19617);
nand U20730 (N_20730,N_19703,N_19896);
nand U20731 (N_20731,N_19762,N_19964);
nand U20732 (N_20732,N_19817,N_19240);
xor U20733 (N_20733,N_19520,N_20294);
xor U20734 (N_20734,N_19413,N_19275);
or U20735 (N_20735,N_20100,N_19535);
nand U20736 (N_20736,N_19676,N_20086);
xnor U20737 (N_20737,N_19608,N_19226);
xnor U20738 (N_20738,N_20098,N_20191);
or U20739 (N_20739,N_19281,N_20347);
and U20740 (N_20740,N_19233,N_20126);
nand U20741 (N_20741,N_19454,N_19688);
nor U20742 (N_20742,N_19681,N_19279);
and U20743 (N_20743,N_20333,N_20029);
nor U20744 (N_20744,N_20273,N_19702);
and U20745 (N_20745,N_20364,N_19864);
or U20746 (N_20746,N_19398,N_19522);
xor U20747 (N_20747,N_20101,N_19298);
or U20748 (N_20748,N_20250,N_19979);
nor U20749 (N_20749,N_19616,N_20350);
or U20750 (N_20750,N_20323,N_19612);
xnor U20751 (N_20751,N_20220,N_20147);
xnor U20752 (N_20752,N_19358,N_19378);
xor U20753 (N_20753,N_20213,N_20166);
and U20754 (N_20754,N_20325,N_19679);
or U20755 (N_20755,N_20223,N_20049);
xnor U20756 (N_20756,N_19952,N_19354);
or U20757 (N_20757,N_20138,N_19214);
and U20758 (N_20758,N_20012,N_19259);
nor U20759 (N_20759,N_19382,N_20072);
and U20760 (N_20760,N_19619,N_20157);
xor U20761 (N_20761,N_19885,N_20018);
or U20762 (N_20762,N_20322,N_19274);
nor U20763 (N_20763,N_19973,N_20280);
and U20764 (N_20764,N_19989,N_19993);
xnor U20765 (N_20765,N_19583,N_19997);
nor U20766 (N_20766,N_19268,N_20385);
and U20767 (N_20767,N_19656,N_19432);
or U20768 (N_20768,N_20392,N_19377);
nor U20769 (N_20769,N_19823,N_19824);
nor U20770 (N_20770,N_19595,N_19948);
nor U20771 (N_20771,N_20177,N_19607);
xor U20772 (N_20772,N_19908,N_19365);
nand U20773 (N_20773,N_19415,N_19370);
xnor U20774 (N_20774,N_19791,N_19200);
xor U20775 (N_20775,N_19787,N_20122);
nand U20776 (N_20776,N_20361,N_19739);
or U20777 (N_20777,N_20181,N_19850);
and U20778 (N_20778,N_20113,N_19402);
nor U20779 (N_20779,N_20243,N_20093);
or U20780 (N_20780,N_19326,N_19720);
xor U20781 (N_20781,N_20308,N_19565);
nor U20782 (N_20782,N_19314,N_19561);
nand U20783 (N_20783,N_19239,N_19508);
nand U20784 (N_20784,N_19625,N_19556);
and U20785 (N_20785,N_20349,N_20179);
and U20786 (N_20786,N_20317,N_19297);
nor U20787 (N_20787,N_19620,N_20154);
and U20788 (N_20788,N_20014,N_19734);
nor U20789 (N_20789,N_20285,N_19986);
nand U20790 (N_20790,N_20146,N_20291);
nand U20791 (N_20791,N_19258,N_19797);
nand U20792 (N_20792,N_19944,N_19571);
nand U20793 (N_20793,N_19542,N_19574);
xnor U20794 (N_20794,N_19665,N_19267);
xnor U20795 (N_20795,N_20172,N_19254);
or U20796 (N_20796,N_20167,N_19844);
nand U20797 (N_20797,N_20121,N_19348);
nor U20798 (N_20798,N_19957,N_20263);
or U20799 (N_20799,N_20114,N_19466);
nor U20800 (N_20800,N_19580,N_20234);
xor U20801 (N_20801,N_19674,N_20261);
xnor U20802 (N_20802,N_20187,N_19310);
xnor U20803 (N_20803,N_19536,N_20056);
nand U20804 (N_20804,N_20208,N_19511);
or U20805 (N_20805,N_19602,N_19644);
and U20806 (N_20806,N_19628,N_20299);
xnor U20807 (N_20807,N_19854,N_19611);
nor U20808 (N_20808,N_19868,N_19932);
nor U20809 (N_20809,N_20235,N_20386);
xnor U20810 (N_20810,N_20030,N_19250);
nor U20811 (N_20811,N_19894,N_19615);
xor U20812 (N_20812,N_20314,N_19411);
and U20813 (N_20813,N_19231,N_19341);
nor U20814 (N_20814,N_20251,N_19609);
xnor U20815 (N_20815,N_20240,N_19218);
and U20816 (N_20816,N_19731,N_20336);
nor U20817 (N_20817,N_19744,N_20120);
nand U20818 (N_20818,N_19433,N_19261);
or U20819 (N_20819,N_19663,N_19467);
and U20820 (N_20820,N_19750,N_19294);
and U20821 (N_20821,N_20076,N_20110);
nand U20822 (N_20822,N_20102,N_19640);
nor U20823 (N_20823,N_19499,N_19329);
nand U20824 (N_20824,N_19501,N_19860);
nand U20825 (N_20825,N_19821,N_19760);
nand U20826 (N_20826,N_19638,N_19660);
nor U20827 (N_20827,N_19690,N_19936);
xor U20828 (N_20828,N_20152,N_20329);
nand U20829 (N_20829,N_20252,N_20044);
and U20830 (N_20830,N_20242,N_19882);
nand U20831 (N_20831,N_19755,N_19687);
nand U20832 (N_20832,N_20052,N_19434);
nand U20833 (N_20833,N_20339,N_19599);
xnor U20834 (N_20834,N_19758,N_19813);
or U20835 (N_20835,N_20218,N_19208);
nand U20836 (N_20836,N_19381,N_20241);
nand U20837 (N_20837,N_19772,N_20019);
nor U20838 (N_20838,N_20151,N_19701);
xor U20839 (N_20839,N_19911,N_19399);
nor U20840 (N_20840,N_19940,N_19480);
or U20841 (N_20841,N_19384,N_20324);
and U20842 (N_20842,N_19623,N_20017);
xnor U20843 (N_20843,N_19715,N_19742);
nand U20844 (N_20844,N_19867,N_19356);
and U20845 (N_20845,N_19295,N_20070);
nor U20846 (N_20846,N_19443,N_19828);
nor U20847 (N_20847,N_19547,N_20067);
or U20848 (N_20848,N_20104,N_19586);
nor U20849 (N_20849,N_19933,N_19809);
and U20850 (N_20850,N_19613,N_20393);
and U20851 (N_20851,N_20374,N_19338);
xor U20852 (N_20852,N_19747,N_19816);
or U20853 (N_20853,N_19642,N_19446);
or U20854 (N_20854,N_19634,N_19733);
and U20855 (N_20855,N_19292,N_20155);
nor U20856 (N_20856,N_19558,N_20031);
or U20857 (N_20857,N_19544,N_19403);
xor U20858 (N_20858,N_20108,N_20053);
and U20859 (N_20859,N_20391,N_19364);
xnor U20860 (N_20860,N_20007,N_19727);
and U20861 (N_20861,N_19531,N_19795);
nand U20862 (N_20862,N_20174,N_19971);
nand U20863 (N_20863,N_19959,N_20383);
or U20864 (N_20864,N_19643,N_19445);
nor U20865 (N_20865,N_20006,N_20310);
nor U20866 (N_20866,N_20010,N_20136);
and U20867 (N_20867,N_20092,N_19532);
or U20868 (N_20868,N_19921,N_20005);
xor U20869 (N_20869,N_19346,N_20265);
nand U20870 (N_20870,N_19313,N_19265);
xor U20871 (N_20871,N_20164,N_20328);
nor U20872 (N_20872,N_19605,N_20228);
or U20873 (N_20873,N_19312,N_19707);
xnor U20874 (N_20874,N_19622,N_19541);
nor U20875 (N_20875,N_20290,N_19347);
or U20876 (N_20876,N_19546,N_20180);
or U20877 (N_20877,N_20128,N_19539);
nor U20878 (N_20878,N_19852,N_19206);
or U20879 (N_20879,N_20215,N_19371);
nor U20880 (N_20880,N_20321,N_20170);
and U20881 (N_20881,N_19651,N_19228);
or U20882 (N_20882,N_19919,N_19488);
nand U20883 (N_20883,N_19876,N_19317);
or U20884 (N_20884,N_19278,N_19212);
and U20885 (N_20885,N_19593,N_19418);
or U20886 (N_20886,N_20139,N_20376);
nand U20887 (N_20887,N_19661,N_19253);
nand U20888 (N_20888,N_20171,N_19695);
xnor U20889 (N_20889,N_20225,N_19811);
and U20890 (N_20890,N_20091,N_20334);
xnor U20891 (N_20891,N_19280,N_19469);
nor U20892 (N_20892,N_19594,N_20300);
or U20893 (N_20893,N_19878,N_20352);
xnor U20894 (N_20894,N_19205,N_19332);
or U20895 (N_20895,N_20331,N_19706);
xor U20896 (N_20896,N_20210,N_19582);
or U20897 (N_20897,N_20173,N_19778);
or U20898 (N_20898,N_19808,N_20340);
and U20899 (N_20899,N_19759,N_20238);
or U20900 (N_20900,N_19591,N_20153);
or U20901 (N_20901,N_19765,N_20202);
and U20902 (N_20902,N_19757,N_19786);
and U20903 (N_20903,N_19914,N_19342);
and U20904 (N_20904,N_20185,N_19977);
xor U20905 (N_20905,N_20200,N_19482);
or U20906 (N_20906,N_19436,N_19627);
nor U20907 (N_20907,N_19277,N_19990);
nor U20908 (N_20908,N_20297,N_19652);
and U20909 (N_20909,N_20293,N_19423);
xnor U20910 (N_20910,N_20289,N_19585);
nand U20911 (N_20911,N_20244,N_20124);
and U20912 (N_20912,N_19427,N_19945);
and U20913 (N_20913,N_19352,N_19856);
or U20914 (N_20914,N_20064,N_20214);
nand U20915 (N_20915,N_20295,N_19322);
and U20916 (N_20916,N_19393,N_19969);
xor U20917 (N_20917,N_19598,N_19881);
and U20918 (N_20918,N_20229,N_20372);
or U20919 (N_20919,N_20320,N_19913);
nor U20920 (N_20920,N_19428,N_20037);
nand U20921 (N_20921,N_19604,N_19405);
nand U20922 (N_20922,N_19984,N_19851);
and U20923 (N_20923,N_19311,N_19899);
or U20924 (N_20924,N_20274,N_20248);
nor U20925 (N_20925,N_19555,N_19624);
nand U20926 (N_20926,N_20111,N_19318);
and U20927 (N_20927,N_20075,N_20026);
nand U20928 (N_20928,N_19471,N_19262);
or U20929 (N_20929,N_19518,N_19474);
nor U20930 (N_20930,N_19777,N_19327);
and U20931 (N_20931,N_19455,N_20335);
and U20932 (N_20932,N_20189,N_19725);
xnor U20933 (N_20933,N_19790,N_19753);
and U20934 (N_20934,N_19224,N_19333);
and U20935 (N_20935,N_19847,N_20140);
xnor U20936 (N_20936,N_19389,N_19316);
and U20937 (N_20937,N_19557,N_19527);
nand U20938 (N_20938,N_19799,N_19339);
nand U20939 (N_20939,N_20379,N_19273);
and U20940 (N_20940,N_19632,N_19284);
nand U20941 (N_20941,N_20028,N_20373);
or U20942 (N_20942,N_20043,N_20266);
nand U20943 (N_20943,N_19965,N_20082);
and U20944 (N_20944,N_19704,N_19830);
xnor U20945 (N_20945,N_19238,N_20395);
xnor U20946 (N_20946,N_19390,N_20256);
or U20947 (N_20947,N_20000,N_19589);
nand U20948 (N_20948,N_19631,N_19492);
and U20949 (N_20949,N_20001,N_19512);
and U20950 (N_20950,N_19385,N_19553);
xnor U20951 (N_20951,N_19570,N_20144);
and U20952 (N_20952,N_19357,N_19666);
and U20953 (N_20953,N_19686,N_19937);
or U20954 (N_20954,N_19463,N_19800);
nor U20955 (N_20955,N_19309,N_19308);
xnor U20956 (N_20956,N_20217,N_20371);
nor U20957 (N_20957,N_19299,N_19723);
or U20958 (N_20958,N_19447,N_19448);
xor U20959 (N_20959,N_19818,N_19798);
xnor U20960 (N_20960,N_19315,N_19941);
or U20961 (N_20961,N_19430,N_20399);
nand U20962 (N_20962,N_19286,N_19234);
xnor U20963 (N_20963,N_19906,N_19328);
or U20964 (N_20964,N_19751,N_19465);
nor U20965 (N_20965,N_20205,N_19672);
nand U20966 (N_20966,N_19810,N_19283);
nor U20967 (N_20967,N_19305,N_20176);
nand U20968 (N_20968,N_19362,N_19293);
xnor U20969 (N_20969,N_19976,N_20069);
or U20970 (N_20970,N_19918,N_19865);
and U20971 (N_20971,N_19361,N_20059);
and U20972 (N_20972,N_19592,N_19590);
nand U20973 (N_20973,N_20344,N_19829);
nor U20974 (N_20974,N_19871,N_19789);
nand U20975 (N_20975,N_19935,N_19414);
and U20976 (N_20976,N_19694,N_19461);
nor U20977 (N_20977,N_20183,N_20083);
xor U20978 (N_20978,N_20066,N_20307);
xor U20979 (N_20979,N_20042,N_19785);
nor U20980 (N_20980,N_19745,N_19947);
or U20981 (N_20981,N_20003,N_19647);
and U20982 (N_20982,N_20035,N_20193);
or U20983 (N_20983,N_19985,N_19201);
nand U20984 (N_20984,N_19344,N_19276);
and U20985 (N_20985,N_20316,N_19614);
xor U20986 (N_20986,N_19938,N_20362);
and U20987 (N_20987,N_20065,N_19978);
nor U20988 (N_20988,N_19998,N_19946);
xor U20989 (N_20989,N_20182,N_19768);
nand U20990 (N_20990,N_19898,N_20309);
nor U20991 (N_20991,N_20040,N_20381);
nand U20992 (N_20992,N_20084,N_20203);
xor U20993 (N_20993,N_19530,N_19884);
nor U20994 (N_20994,N_19954,N_19736);
or U20995 (N_20995,N_19223,N_19838);
and U20996 (N_20996,N_19722,N_19618);
and U20997 (N_20997,N_19752,N_19504);
nand U20998 (N_20998,N_19792,N_19887);
nor U20999 (N_20999,N_19395,N_19481);
or U21000 (N_21000,N_19879,N_19357);
or U21001 (N_21001,N_19781,N_19467);
and U21002 (N_21002,N_19596,N_19713);
xnor U21003 (N_21003,N_19411,N_20108);
xor U21004 (N_21004,N_20115,N_19524);
xor U21005 (N_21005,N_20248,N_19314);
or U21006 (N_21006,N_19619,N_19310);
or U21007 (N_21007,N_19858,N_19959);
nand U21008 (N_21008,N_19650,N_19889);
or U21009 (N_21009,N_19476,N_19660);
nor U21010 (N_21010,N_19491,N_19684);
nor U21011 (N_21011,N_19989,N_19555);
nor U21012 (N_21012,N_19966,N_20297);
or U21013 (N_21013,N_19854,N_19519);
or U21014 (N_21014,N_19668,N_19361);
and U21015 (N_21015,N_20255,N_19462);
nor U21016 (N_21016,N_19523,N_19295);
or U21017 (N_21017,N_19454,N_20025);
nor U21018 (N_21018,N_19706,N_19203);
xor U21019 (N_21019,N_20166,N_20080);
nor U21020 (N_21020,N_20254,N_20346);
or U21021 (N_21021,N_20037,N_19719);
nor U21022 (N_21022,N_20026,N_20223);
or U21023 (N_21023,N_19609,N_19790);
or U21024 (N_21024,N_19294,N_19409);
or U21025 (N_21025,N_19475,N_19586);
nor U21026 (N_21026,N_20132,N_19521);
nand U21027 (N_21027,N_19784,N_20046);
or U21028 (N_21028,N_20046,N_20190);
xor U21029 (N_21029,N_19961,N_19342);
and U21030 (N_21030,N_20178,N_19352);
or U21031 (N_21031,N_19861,N_20220);
xnor U21032 (N_21032,N_19963,N_19921);
nand U21033 (N_21033,N_19611,N_19381);
and U21034 (N_21034,N_19507,N_19971);
nand U21035 (N_21035,N_19753,N_19507);
nor U21036 (N_21036,N_19404,N_19466);
nor U21037 (N_21037,N_19473,N_19324);
nor U21038 (N_21038,N_20209,N_19649);
xor U21039 (N_21039,N_20204,N_19781);
nor U21040 (N_21040,N_20041,N_19967);
or U21041 (N_21041,N_19271,N_19857);
nor U21042 (N_21042,N_19839,N_20356);
nor U21043 (N_21043,N_20248,N_19429);
and U21044 (N_21044,N_19775,N_19785);
xor U21045 (N_21045,N_20355,N_19714);
xor U21046 (N_21046,N_19474,N_19972);
nand U21047 (N_21047,N_19405,N_20297);
nor U21048 (N_21048,N_20125,N_20367);
nor U21049 (N_21049,N_19786,N_20256);
or U21050 (N_21050,N_19339,N_20264);
nor U21051 (N_21051,N_19429,N_19523);
and U21052 (N_21052,N_20173,N_19711);
nor U21053 (N_21053,N_20113,N_19352);
nand U21054 (N_21054,N_20111,N_19233);
nor U21055 (N_21055,N_19662,N_20019);
xor U21056 (N_21056,N_20018,N_19575);
nor U21057 (N_21057,N_19373,N_19673);
nand U21058 (N_21058,N_20211,N_20236);
and U21059 (N_21059,N_19863,N_20180);
and U21060 (N_21060,N_19336,N_19911);
or U21061 (N_21061,N_19663,N_20056);
or U21062 (N_21062,N_19896,N_19672);
nand U21063 (N_21063,N_20166,N_20068);
xor U21064 (N_21064,N_19268,N_19254);
nand U21065 (N_21065,N_19942,N_19752);
or U21066 (N_21066,N_19725,N_19962);
or U21067 (N_21067,N_20229,N_19800);
and U21068 (N_21068,N_19911,N_20316);
or U21069 (N_21069,N_19279,N_20244);
nand U21070 (N_21070,N_19557,N_19491);
xor U21071 (N_21071,N_19366,N_20091);
nand U21072 (N_21072,N_20285,N_20066);
nand U21073 (N_21073,N_19329,N_19663);
nand U21074 (N_21074,N_19583,N_19585);
nor U21075 (N_21075,N_19389,N_19543);
nand U21076 (N_21076,N_20326,N_19858);
xnor U21077 (N_21077,N_19709,N_19252);
nor U21078 (N_21078,N_20156,N_19755);
xor U21079 (N_21079,N_20154,N_20155);
nor U21080 (N_21080,N_19314,N_19206);
or U21081 (N_21081,N_20072,N_19565);
xnor U21082 (N_21082,N_19775,N_19569);
xnor U21083 (N_21083,N_19805,N_20155);
nand U21084 (N_21084,N_19863,N_19554);
nor U21085 (N_21085,N_19715,N_19349);
xnor U21086 (N_21086,N_20276,N_19790);
xnor U21087 (N_21087,N_19811,N_20135);
and U21088 (N_21088,N_19951,N_19839);
and U21089 (N_21089,N_20034,N_19820);
or U21090 (N_21090,N_19773,N_19563);
and U21091 (N_21091,N_19480,N_19236);
xnor U21092 (N_21092,N_19696,N_19505);
nand U21093 (N_21093,N_20258,N_19458);
xor U21094 (N_21094,N_20211,N_19946);
nand U21095 (N_21095,N_19428,N_19750);
xnor U21096 (N_21096,N_19975,N_19255);
xnor U21097 (N_21097,N_19296,N_19827);
nand U21098 (N_21098,N_19459,N_20358);
or U21099 (N_21099,N_19581,N_19972);
nand U21100 (N_21100,N_19218,N_20290);
or U21101 (N_21101,N_19455,N_19948);
xor U21102 (N_21102,N_20202,N_19325);
nor U21103 (N_21103,N_19350,N_19808);
nor U21104 (N_21104,N_19654,N_20203);
or U21105 (N_21105,N_19368,N_20399);
nor U21106 (N_21106,N_19490,N_19917);
or U21107 (N_21107,N_19597,N_20145);
nor U21108 (N_21108,N_19500,N_20044);
or U21109 (N_21109,N_19781,N_20236);
or U21110 (N_21110,N_19766,N_19814);
nand U21111 (N_21111,N_19674,N_19847);
nor U21112 (N_21112,N_20385,N_19281);
nand U21113 (N_21113,N_19910,N_20335);
nor U21114 (N_21114,N_19208,N_19310);
nor U21115 (N_21115,N_20041,N_20190);
and U21116 (N_21116,N_19437,N_19252);
nand U21117 (N_21117,N_20164,N_19807);
nor U21118 (N_21118,N_19798,N_19312);
and U21119 (N_21119,N_19465,N_19951);
nor U21120 (N_21120,N_20312,N_20373);
xor U21121 (N_21121,N_20241,N_19373);
or U21122 (N_21122,N_19892,N_19297);
or U21123 (N_21123,N_19699,N_19287);
nor U21124 (N_21124,N_20278,N_19918);
nand U21125 (N_21125,N_20004,N_19304);
nand U21126 (N_21126,N_19786,N_19942);
nand U21127 (N_21127,N_20031,N_19464);
xor U21128 (N_21128,N_19815,N_19751);
nand U21129 (N_21129,N_19886,N_19379);
or U21130 (N_21130,N_19799,N_19593);
nor U21131 (N_21131,N_20301,N_20322);
and U21132 (N_21132,N_19293,N_19974);
nand U21133 (N_21133,N_19553,N_20222);
or U21134 (N_21134,N_19308,N_19376);
and U21135 (N_21135,N_19480,N_20041);
xnor U21136 (N_21136,N_19954,N_19680);
or U21137 (N_21137,N_19618,N_19988);
and U21138 (N_21138,N_20346,N_19990);
nand U21139 (N_21139,N_19423,N_19662);
or U21140 (N_21140,N_19340,N_19842);
nand U21141 (N_21141,N_19293,N_20253);
or U21142 (N_21142,N_20387,N_19838);
or U21143 (N_21143,N_19904,N_19378);
nand U21144 (N_21144,N_19323,N_19877);
or U21145 (N_21145,N_20034,N_19234);
nor U21146 (N_21146,N_20331,N_20200);
xnor U21147 (N_21147,N_19490,N_19764);
nand U21148 (N_21148,N_19237,N_20299);
nand U21149 (N_21149,N_19366,N_19683);
nor U21150 (N_21150,N_20130,N_19797);
or U21151 (N_21151,N_19431,N_20392);
nor U21152 (N_21152,N_20345,N_19533);
nor U21153 (N_21153,N_19940,N_19496);
xnor U21154 (N_21154,N_19404,N_19653);
and U21155 (N_21155,N_20101,N_19560);
nand U21156 (N_21156,N_20003,N_20135);
nor U21157 (N_21157,N_19698,N_19438);
or U21158 (N_21158,N_20188,N_19946);
or U21159 (N_21159,N_19315,N_19552);
or U21160 (N_21160,N_20190,N_20243);
nor U21161 (N_21161,N_19556,N_19690);
and U21162 (N_21162,N_19443,N_20052);
nor U21163 (N_21163,N_19215,N_19844);
xor U21164 (N_21164,N_19208,N_19746);
nand U21165 (N_21165,N_19283,N_20322);
xor U21166 (N_21166,N_20002,N_19776);
nand U21167 (N_21167,N_19313,N_19466);
or U21168 (N_21168,N_19349,N_20232);
nor U21169 (N_21169,N_20272,N_19280);
nor U21170 (N_21170,N_19684,N_19404);
or U21171 (N_21171,N_20102,N_19641);
or U21172 (N_21172,N_19579,N_20258);
nor U21173 (N_21173,N_19820,N_19936);
nand U21174 (N_21174,N_20188,N_20088);
nor U21175 (N_21175,N_19872,N_20025);
and U21176 (N_21176,N_19718,N_20301);
and U21177 (N_21177,N_19689,N_20146);
nand U21178 (N_21178,N_20277,N_19310);
xor U21179 (N_21179,N_19543,N_19209);
xnor U21180 (N_21180,N_19659,N_19613);
xnor U21181 (N_21181,N_19471,N_19559);
nor U21182 (N_21182,N_19326,N_20310);
or U21183 (N_21183,N_19524,N_20361);
or U21184 (N_21184,N_19485,N_19985);
xor U21185 (N_21185,N_19642,N_19958);
and U21186 (N_21186,N_19282,N_19579);
nor U21187 (N_21187,N_20220,N_19296);
and U21188 (N_21188,N_19424,N_19491);
or U21189 (N_21189,N_20355,N_19620);
nor U21190 (N_21190,N_19821,N_19959);
and U21191 (N_21191,N_19995,N_20214);
nand U21192 (N_21192,N_19386,N_19437);
nor U21193 (N_21193,N_19853,N_20227);
xor U21194 (N_21194,N_20130,N_19369);
and U21195 (N_21195,N_20253,N_19712);
and U21196 (N_21196,N_19326,N_20117);
nor U21197 (N_21197,N_20341,N_20135);
nand U21198 (N_21198,N_20132,N_19860);
nand U21199 (N_21199,N_19799,N_19970);
and U21200 (N_21200,N_20294,N_19230);
and U21201 (N_21201,N_19445,N_19258);
nand U21202 (N_21202,N_19699,N_20378);
xor U21203 (N_21203,N_20104,N_19421);
nor U21204 (N_21204,N_20383,N_19899);
or U21205 (N_21205,N_19477,N_20364);
xor U21206 (N_21206,N_19232,N_19721);
nor U21207 (N_21207,N_19604,N_19841);
nor U21208 (N_21208,N_20088,N_19865);
or U21209 (N_21209,N_19382,N_19201);
nor U21210 (N_21210,N_19458,N_19502);
or U21211 (N_21211,N_20025,N_19904);
nand U21212 (N_21212,N_20274,N_20035);
or U21213 (N_21213,N_19224,N_19278);
nor U21214 (N_21214,N_19638,N_19314);
nor U21215 (N_21215,N_19795,N_19472);
nor U21216 (N_21216,N_19827,N_19722);
and U21217 (N_21217,N_19975,N_20059);
xor U21218 (N_21218,N_19321,N_19943);
nor U21219 (N_21219,N_19408,N_20015);
nor U21220 (N_21220,N_19711,N_19889);
nor U21221 (N_21221,N_19301,N_19313);
and U21222 (N_21222,N_19999,N_20169);
or U21223 (N_21223,N_20037,N_19605);
nor U21224 (N_21224,N_19829,N_19589);
or U21225 (N_21225,N_19648,N_19419);
nor U21226 (N_21226,N_19539,N_19499);
nand U21227 (N_21227,N_19460,N_20317);
and U21228 (N_21228,N_20095,N_19803);
xnor U21229 (N_21229,N_19846,N_19409);
and U21230 (N_21230,N_19850,N_19838);
or U21231 (N_21231,N_19650,N_20308);
and U21232 (N_21232,N_19926,N_19876);
or U21233 (N_21233,N_19892,N_19601);
nor U21234 (N_21234,N_20274,N_19611);
xor U21235 (N_21235,N_20106,N_19500);
nor U21236 (N_21236,N_20334,N_19569);
nand U21237 (N_21237,N_20366,N_19609);
and U21238 (N_21238,N_19833,N_19284);
xnor U21239 (N_21239,N_19329,N_19551);
nand U21240 (N_21240,N_19498,N_20155);
nand U21241 (N_21241,N_19240,N_19617);
nor U21242 (N_21242,N_19395,N_19955);
or U21243 (N_21243,N_19957,N_19223);
or U21244 (N_21244,N_19608,N_19699);
and U21245 (N_21245,N_19941,N_19295);
xor U21246 (N_21246,N_19224,N_19272);
or U21247 (N_21247,N_19373,N_19279);
nand U21248 (N_21248,N_19421,N_19966);
nor U21249 (N_21249,N_20110,N_19684);
and U21250 (N_21250,N_19451,N_19884);
and U21251 (N_21251,N_19933,N_19449);
and U21252 (N_21252,N_19360,N_19361);
nand U21253 (N_21253,N_19809,N_19773);
and U21254 (N_21254,N_19430,N_19508);
and U21255 (N_21255,N_19937,N_19245);
and U21256 (N_21256,N_19653,N_19866);
nand U21257 (N_21257,N_20231,N_19500);
xor U21258 (N_21258,N_19588,N_19451);
nor U21259 (N_21259,N_19655,N_19861);
nand U21260 (N_21260,N_20063,N_20324);
and U21261 (N_21261,N_19732,N_19797);
nor U21262 (N_21262,N_20329,N_19875);
nand U21263 (N_21263,N_20309,N_20380);
xnor U21264 (N_21264,N_20399,N_19266);
or U21265 (N_21265,N_19532,N_20274);
and U21266 (N_21266,N_19385,N_20172);
nand U21267 (N_21267,N_19857,N_19563);
nand U21268 (N_21268,N_19512,N_20287);
and U21269 (N_21269,N_19439,N_20013);
and U21270 (N_21270,N_19268,N_19307);
xor U21271 (N_21271,N_19373,N_19226);
nor U21272 (N_21272,N_19376,N_19270);
or U21273 (N_21273,N_19935,N_20071);
xor U21274 (N_21274,N_20309,N_20032);
or U21275 (N_21275,N_19390,N_19961);
xnor U21276 (N_21276,N_20202,N_20324);
nand U21277 (N_21277,N_20381,N_20374);
nand U21278 (N_21278,N_20282,N_19531);
nand U21279 (N_21279,N_20296,N_19610);
and U21280 (N_21280,N_20376,N_20176);
xnor U21281 (N_21281,N_19289,N_19645);
nand U21282 (N_21282,N_20204,N_20271);
nor U21283 (N_21283,N_19991,N_20195);
nand U21284 (N_21284,N_20116,N_19570);
nor U21285 (N_21285,N_19982,N_19285);
and U21286 (N_21286,N_19971,N_19299);
or U21287 (N_21287,N_20055,N_19256);
nand U21288 (N_21288,N_19299,N_20243);
and U21289 (N_21289,N_19260,N_20076);
xnor U21290 (N_21290,N_19946,N_20344);
or U21291 (N_21291,N_19484,N_20217);
or U21292 (N_21292,N_19793,N_19789);
nand U21293 (N_21293,N_19443,N_20084);
xor U21294 (N_21294,N_19983,N_19809);
or U21295 (N_21295,N_20270,N_19352);
nand U21296 (N_21296,N_20390,N_19840);
and U21297 (N_21297,N_20041,N_20344);
or U21298 (N_21298,N_19261,N_19521);
and U21299 (N_21299,N_19589,N_19377);
and U21300 (N_21300,N_19973,N_20024);
and U21301 (N_21301,N_19843,N_19832);
or U21302 (N_21302,N_19605,N_19275);
nand U21303 (N_21303,N_19866,N_20218);
and U21304 (N_21304,N_19736,N_20193);
xnor U21305 (N_21305,N_19735,N_20197);
and U21306 (N_21306,N_19324,N_19954);
and U21307 (N_21307,N_20254,N_20050);
nand U21308 (N_21308,N_19742,N_19550);
xnor U21309 (N_21309,N_19233,N_19722);
xnor U21310 (N_21310,N_19552,N_19691);
and U21311 (N_21311,N_20045,N_19745);
nand U21312 (N_21312,N_20118,N_20197);
and U21313 (N_21313,N_19427,N_20376);
or U21314 (N_21314,N_20146,N_20069);
and U21315 (N_21315,N_20383,N_20123);
nand U21316 (N_21316,N_20179,N_19365);
or U21317 (N_21317,N_19589,N_20370);
and U21318 (N_21318,N_20155,N_19394);
and U21319 (N_21319,N_20128,N_19990);
or U21320 (N_21320,N_20314,N_19744);
nand U21321 (N_21321,N_20099,N_20345);
and U21322 (N_21322,N_19795,N_19742);
nor U21323 (N_21323,N_20265,N_19241);
nor U21324 (N_21324,N_19690,N_20252);
nand U21325 (N_21325,N_19507,N_20113);
xnor U21326 (N_21326,N_19790,N_20103);
or U21327 (N_21327,N_19677,N_19834);
xnor U21328 (N_21328,N_19762,N_19246);
xor U21329 (N_21329,N_19498,N_19973);
nand U21330 (N_21330,N_20026,N_19238);
xor U21331 (N_21331,N_19696,N_20098);
nand U21332 (N_21332,N_19420,N_19796);
xnor U21333 (N_21333,N_19202,N_19475);
nand U21334 (N_21334,N_19586,N_20292);
and U21335 (N_21335,N_19940,N_19931);
and U21336 (N_21336,N_19539,N_19483);
xnor U21337 (N_21337,N_19703,N_19408);
nand U21338 (N_21338,N_20315,N_19937);
xor U21339 (N_21339,N_20218,N_19941);
nand U21340 (N_21340,N_19910,N_19288);
xnor U21341 (N_21341,N_19233,N_19868);
or U21342 (N_21342,N_19262,N_19432);
nand U21343 (N_21343,N_19577,N_19307);
nor U21344 (N_21344,N_19993,N_19936);
and U21345 (N_21345,N_19209,N_19222);
and U21346 (N_21346,N_19364,N_19834);
and U21347 (N_21347,N_19352,N_20043);
and U21348 (N_21348,N_19506,N_19858);
nor U21349 (N_21349,N_19442,N_19627);
nor U21350 (N_21350,N_19647,N_20313);
and U21351 (N_21351,N_19838,N_20329);
or U21352 (N_21352,N_19583,N_19835);
nor U21353 (N_21353,N_19596,N_19361);
or U21354 (N_21354,N_20349,N_20105);
nand U21355 (N_21355,N_19996,N_20243);
nand U21356 (N_21356,N_20023,N_20168);
nand U21357 (N_21357,N_19870,N_19328);
nand U21358 (N_21358,N_19449,N_20390);
nor U21359 (N_21359,N_19668,N_19507);
nor U21360 (N_21360,N_19692,N_20242);
and U21361 (N_21361,N_20226,N_20302);
xnor U21362 (N_21362,N_19951,N_20340);
nor U21363 (N_21363,N_20135,N_19880);
and U21364 (N_21364,N_19215,N_19931);
xor U21365 (N_21365,N_19624,N_19232);
nor U21366 (N_21366,N_20388,N_20042);
and U21367 (N_21367,N_20092,N_20127);
nand U21368 (N_21368,N_20086,N_19981);
nand U21369 (N_21369,N_20073,N_19300);
nor U21370 (N_21370,N_19610,N_19200);
nand U21371 (N_21371,N_19526,N_19683);
and U21372 (N_21372,N_19440,N_20212);
xnor U21373 (N_21373,N_19488,N_19254);
nand U21374 (N_21374,N_20179,N_19473);
xnor U21375 (N_21375,N_20038,N_20383);
and U21376 (N_21376,N_19904,N_20343);
and U21377 (N_21377,N_19883,N_20392);
xor U21378 (N_21378,N_20229,N_20129);
or U21379 (N_21379,N_20147,N_19311);
or U21380 (N_21380,N_19235,N_20177);
xnor U21381 (N_21381,N_19965,N_20066);
nor U21382 (N_21382,N_19515,N_20096);
nor U21383 (N_21383,N_19472,N_19271);
nor U21384 (N_21384,N_19768,N_20195);
xnor U21385 (N_21385,N_19630,N_19289);
nand U21386 (N_21386,N_20396,N_20251);
xnor U21387 (N_21387,N_19944,N_19353);
or U21388 (N_21388,N_20364,N_19453);
xor U21389 (N_21389,N_19544,N_19491);
or U21390 (N_21390,N_20074,N_19789);
xor U21391 (N_21391,N_19481,N_20257);
or U21392 (N_21392,N_20315,N_19465);
or U21393 (N_21393,N_19825,N_20138);
xor U21394 (N_21394,N_19333,N_19853);
nand U21395 (N_21395,N_19894,N_19503);
nor U21396 (N_21396,N_19748,N_19749);
nor U21397 (N_21397,N_19999,N_19835);
xor U21398 (N_21398,N_19340,N_19876);
or U21399 (N_21399,N_20196,N_19481);
nand U21400 (N_21400,N_20249,N_19468);
or U21401 (N_21401,N_19852,N_19793);
nor U21402 (N_21402,N_20248,N_19517);
nor U21403 (N_21403,N_19716,N_20189);
nor U21404 (N_21404,N_19464,N_19828);
nor U21405 (N_21405,N_20389,N_19461);
xnor U21406 (N_21406,N_20084,N_19958);
nand U21407 (N_21407,N_19276,N_19380);
xor U21408 (N_21408,N_20274,N_19380);
and U21409 (N_21409,N_19660,N_19331);
or U21410 (N_21410,N_19496,N_19320);
nand U21411 (N_21411,N_19807,N_19961);
nor U21412 (N_21412,N_20233,N_19358);
and U21413 (N_21413,N_19819,N_20017);
and U21414 (N_21414,N_19546,N_20178);
and U21415 (N_21415,N_19330,N_19772);
or U21416 (N_21416,N_19678,N_19825);
or U21417 (N_21417,N_19332,N_20327);
nand U21418 (N_21418,N_20025,N_19635);
nand U21419 (N_21419,N_19306,N_19388);
or U21420 (N_21420,N_19316,N_19219);
nor U21421 (N_21421,N_19471,N_19661);
and U21422 (N_21422,N_19904,N_19301);
nor U21423 (N_21423,N_19474,N_19275);
xor U21424 (N_21424,N_19553,N_19426);
nand U21425 (N_21425,N_19396,N_19714);
xnor U21426 (N_21426,N_20315,N_19660);
nand U21427 (N_21427,N_20114,N_19974);
xor U21428 (N_21428,N_19240,N_19585);
and U21429 (N_21429,N_20339,N_19503);
nand U21430 (N_21430,N_20097,N_20194);
nor U21431 (N_21431,N_20181,N_19917);
and U21432 (N_21432,N_20327,N_19712);
nor U21433 (N_21433,N_19403,N_20263);
nor U21434 (N_21434,N_19698,N_19995);
nand U21435 (N_21435,N_19267,N_19999);
nor U21436 (N_21436,N_19640,N_19862);
and U21437 (N_21437,N_19653,N_19976);
nor U21438 (N_21438,N_19476,N_20283);
xor U21439 (N_21439,N_19496,N_20102);
and U21440 (N_21440,N_19334,N_19780);
xor U21441 (N_21441,N_19419,N_19265);
or U21442 (N_21442,N_19297,N_19320);
nor U21443 (N_21443,N_20305,N_20044);
nand U21444 (N_21444,N_19746,N_19401);
nand U21445 (N_21445,N_19815,N_19534);
and U21446 (N_21446,N_19759,N_19634);
xnor U21447 (N_21447,N_19935,N_19511);
nand U21448 (N_21448,N_19637,N_19651);
nor U21449 (N_21449,N_20026,N_19423);
nand U21450 (N_21450,N_19930,N_19769);
and U21451 (N_21451,N_19479,N_19817);
nand U21452 (N_21452,N_19540,N_19766);
and U21453 (N_21453,N_19395,N_19740);
nand U21454 (N_21454,N_19466,N_20202);
and U21455 (N_21455,N_19855,N_20109);
xor U21456 (N_21456,N_20150,N_19528);
or U21457 (N_21457,N_19493,N_20041);
xor U21458 (N_21458,N_19479,N_19596);
or U21459 (N_21459,N_19352,N_20126);
and U21460 (N_21460,N_20321,N_19998);
or U21461 (N_21461,N_19878,N_19673);
and U21462 (N_21462,N_20127,N_19352);
or U21463 (N_21463,N_19859,N_19338);
nor U21464 (N_21464,N_19281,N_19722);
or U21465 (N_21465,N_20256,N_19230);
xnor U21466 (N_21466,N_20007,N_19894);
or U21467 (N_21467,N_19919,N_19534);
nand U21468 (N_21468,N_19395,N_19418);
and U21469 (N_21469,N_20203,N_20362);
or U21470 (N_21470,N_20098,N_20111);
nor U21471 (N_21471,N_19572,N_19340);
nand U21472 (N_21472,N_19884,N_19528);
nand U21473 (N_21473,N_19937,N_19660);
or U21474 (N_21474,N_19280,N_19869);
xor U21475 (N_21475,N_19630,N_19299);
nor U21476 (N_21476,N_20257,N_20142);
nor U21477 (N_21477,N_19492,N_20298);
xor U21478 (N_21478,N_19307,N_19304);
nor U21479 (N_21479,N_20303,N_20244);
xnor U21480 (N_21480,N_20350,N_19735);
xor U21481 (N_21481,N_20129,N_19598);
nor U21482 (N_21482,N_19482,N_19943);
and U21483 (N_21483,N_20347,N_20338);
or U21484 (N_21484,N_19220,N_19353);
nand U21485 (N_21485,N_19899,N_20363);
xnor U21486 (N_21486,N_19613,N_20387);
nor U21487 (N_21487,N_20055,N_19547);
and U21488 (N_21488,N_19446,N_19430);
xor U21489 (N_21489,N_19406,N_20118);
and U21490 (N_21490,N_19846,N_19960);
and U21491 (N_21491,N_20106,N_19301);
or U21492 (N_21492,N_19504,N_19881);
nor U21493 (N_21493,N_19799,N_20001);
nand U21494 (N_21494,N_20129,N_19768);
nor U21495 (N_21495,N_19208,N_19965);
xnor U21496 (N_21496,N_19579,N_19665);
nand U21497 (N_21497,N_20326,N_20006);
and U21498 (N_21498,N_19900,N_19890);
and U21499 (N_21499,N_20335,N_20137);
nor U21500 (N_21500,N_19498,N_19638);
nand U21501 (N_21501,N_19480,N_20363);
nor U21502 (N_21502,N_19461,N_19649);
or U21503 (N_21503,N_20193,N_19273);
and U21504 (N_21504,N_19662,N_19452);
or U21505 (N_21505,N_19571,N_19323);
xnor U21506 (N_21506,N_19240,N_20317);
nand U21507 (N_21507,N_20393,N_20165);
and U21508 (N_21508,N_19572,N_19970);
nor U21509 (N_21509,N_20288,N_20178);
and U21510 (N_21510,N_20263,N_19345);
or U21511 (N_21511,N_19378,N_20107);
and U21512 (N_21512,N_19907,N_20085);
or U21513 (N_21513,N_19630,N_20333);
and U21514 (N_21514,N_19647,N_20008);
and U21515 (N_21515,N_20323,N_20322);
and U21516 (N_21516,N_19911,N_20345);
and U21517 (N_21517,N_19383,N_19937);
nand U21518 (N_21518,N_20245,N_19853);
nor U21519 (N_21519,N_19508,N_20172);
nand U21520 (N_21520,N_19427,N_19469);
or U21521 (N_21521,N_19674,N_19216);
xnor U21522 (N_21522,N_19928,N_20177);
nand U21523 (N_21523,N_19263,N_19612);
xor U21524 (N_21524,N_19620,N_20231);
nor U21525 (N_21525,N_20112,N_19740);
nand U21526 (N_21526,N_20390,N_19839);
nand U21527 (N_21527,N_19290,N_20213);
nor U21528 (N_21528,N_19990,N_19999);
nand U21529 (N_21529,N_19475,N_20222);
nor U21530 (N_21530,N_19480,N_20288);
nor U21531 (N_21531,N_20068,N_20143);
and U21532 (N_21532,N_19326,N_19615);
nor U21533 (N_21533,N_19804,N_19651);
nor U21534 (N_21534,N_20080,N_20353);
nand U21535 (N_21535,N_19286,N_19949);
xor U21536 (N_21536,N_19635,N_20044);
and U21537 (N_21537,N_19992,N_20335);
xor U21538 (N_21538,N_19930,N_19223);
and U21539 (N_21539,N_19420,N_19590);
xnor U21540 (N_21540,N_20180,N_19430);
nand U21541 (N_21541,N_19462,N_19293);
and U21542 (N_21542,N_20066,N_20036);
nor U21543 (N_21543,N_20332,N_20091);
xor U21544 (N_21544,N_19467,N_20275);
and U21545 (N_21545,N_20157,N_19965);
xnor U21546 (N_21546,N_19762,N_19852);
nor U21547 (N_21547,N_19406,N_19677);
xor U21548 (N_21548,N_19840,N_19485);
nor U21549 (N_21549,N_20040,N_19902);
nand U21550 (N_21550,N_19511,N_19267);
and U21551 (N_21551,N_19805,N_19742);
xnor U21552 (N_21552,N_19649,N_19257);
nor U21553 (N_21553,N_19475,N_20132);
nor U21554 (N_21554,N_19281,N_20026);
xnor U21555 (N_21555,N_20246,N_19658);
or U21556 (N_21556,N_20288,N_19508);
and U21557 (N_21557,N_19287,N_19670);
nor U21558 (N_21558,N_19915,N_19201);
and U21559 (N_21559,N_19602,N_19982);
and U21560 (N_21560,N_19644,N_19933);
nand U21561 (N_21561,N_20194,N_19552);
nor U21562 (N_21562,N_19291,N_19425);
nand U21563 (N_21563,N_19635,N_19911);
and U21564 (N_21564,N_19549,N_19709);
or U21565 (N_21565,N_19347,N_20297);
and U21566 (N_21566,N_19566,N_19621);
nor U21567 (N_21567,N_19528,N_20161);
or U21568 (N_21568,N_19763,N_19240);
xnor U21569 (N_21569,N_19250,N_20036);
nand U21570 (N_21570,N_19225,N_19421);
nor U21571 (N_21571,N_19866,N_19703);
or U21572 (N_21572,N_19366,N_19973);
nor U21573 (N_21573,N_19270,N_19509);
or U21574 (N_21574,N_20163,N_20052);
xnor U21575 (N_21575,N_19831,N_20034);
and U21576 (N_21576,N_20176,N_20058);
nor U21577 (N_21577,N_19368,N_19926);
xor U21578 (N_21578,N_19474,N_19750);
and U21579 (N_21579,N_20330,N_19905);
nand U21580 (N_21580,N_19860,N_19819);
nor U21581 (N_21581,N_19372,N_20392);
nor U21582 (N_21582,N_19981,N_19523);
nor U21583 (N_21583,N_20079,N_20265);
and U21584 (N_21584,N_19303,N_19636);
xor U21585 (N_21585,N_19938,N_19731);
nand U21586 (N_21586,N_19612,N_19668);
and U21587 (N_21587,N_19943,N_19743);
or U21588 (N_21588,N_19305,N_20204);
nand U21589 (N_21589,N_19840,N_20143);
nor U21590 (N_21590,N_19265,N_19902);
xor U21591 (N_21591,N_20385,N_20180);
and U21592 (N_21592,N_19971,N_20364);
nor U21593 (N_21593,N_19665,N_19349);
xnor U21594 (N_21594,N_19334,N_19591);
and U21595 (N_21595,N_19534,N_19351);
nand U21596 (N_21596,N_19697,N_20049);
nor U21597 (N_21597,N_19792,N_19884);
or U21598 (N_21598,N_20179,N_20019);
and U21599 (N_21599,N_20223,N_19673);
and U21600 (N_21600,N_20404,N_21224);
nand U21601 (N_21601,N_20801,N_20710);
xor U21602 (N_21602,N_21083,N_21547);
and U21603 (N_21603,N_20683,N_21414);
or U21604 (N_21604,N_21256,N_21361);
nor U21605 (N_21605,N_21472,N_20927);
xor U21606 (N_21606,N_21548,N_21596);
xor U21607 (N_21607,N_21282,N_20735);
or U21608 (N_21608,N_21305,N_20776);
or U21609 (N_21609,N_21303,N_20437);
xnor U21610 (N_21610,N_21258,N_20850);
xnor U21611 (N_21611,N_21501,N_21125);
and U21612 (N_21612,N_21434,N_21079);
nand U21613 (N_21613,N_20548,N_20601);
or U21614 (N_21614,N_21112,N_21477);
and U21615 (N_21615,N_21595,N_21337);
and U21616 (N_21616,N_21397,N_21494);
and U21617 (N_21617,N_21302,N_20986);
nand U21618 (N_21618,N_20874,N_21425);
nor U21619 (N_21619,N_21516,N_21463);
and U21620 (N_21620,N_21014,N_20833);
xor U21621 (N_21621,N_20894,N_21413);
xor U21622 (N_21622,N_21242,N_21149);
or U21623 (N_21623,N_21520,N_21571);
nand U21624 (N_21624,N_21190,N_20538);
xnor U21625 (N_21625,N_21288,N_20722);
nand U21626 (N_21626,N_21567,N_21390);
xor U21627 (N_21627,N_21357,N_21212);
or U21628 (N_21628,N_21591,N_21101);
and U21629 (N_21629,N_21121,N_20493);
and U21630 (N_21630,N_21369,N_21323);
xor U21631 (N_21631,N_21013,N_21515);
nor U21632 (N_21632,N_20803,N_21073);
or U21633 (N_21633,N_21445,N_21284);
and U21634 (N_21634,N_21245,N_20810);
xnor U21635 (N_21635,N_21575,N_20694);
and U21636 (N_21636,N_20889,N_21106);
nand U21637 (N_21637,N_21159,N_21485);
xor U21638 (N_21638,N_20549,N_21069);
and U21639 (N_21639,N_21329,N_21031);
xor U21640 (N_21640,N_20862,N_20996);
nand U21641 (N_21641,N_20408,N_21119);
and U21642 (N_21642,N_20854,N_20793);
nor U21643 (N_21643,N_20488,N_20650);
and U21644 (N_21644,N_21180,N_20730);
xnor U21645 (N_21645,N_21195,N_20899);
and U21646 (N_21646,N_20812,N_20980);
nand U21647 (N_21647,N_21133,N_20705);
xnor U21648 (N_21648,N_20435,N_20764);
or U21649 (N_21649,N_20753,N_21495);
nor U21650 (N_21650,N_20690,N_21569);
nor U21651 (N_21651,N_21071,N_20529);
xor U21652 (N_21652,N_21253,N_21024);
xnor U21653 (N_21653,N_20796,N_21410);
nand U21654 (N_21654,N_21111,N_20808);
or U21655 (N_21655,N_20841,N_21115);
nor U21656 (N_21656,N_20863,N_21244);
xnor U21657 (N_21657,N_21285,N_21401);
or U21658 (N_21658,N_21273,N_20798);
nor U21659 (N_21659,N_21298,N_21088);
nor U21660 (N_21660,N_20870,N_20684);
nor U21661 (N_21661,N_20733,N_20584);
nor U21662 (N_21662,N_21448,N_21034);
nor U21663 (N_21663,N_21093,N_21446);
nand U21664 (N_21664,N_20550,N_20706);
or U21665 (N_21665,N_21549,N_21469);
nand U21666 (N_21666,N_20979,N_20610);
nand U21667 (N_21667,N_21379,N_20726);
and U21668 (N_21668,N_20868,N_21082);
or U21669 (N_21669,N_21551,N_21312);
and U21670 (N_21670,N_21192,N_20648);
nor U21671 (N_21671,N_21290,N_21336);
nor U21672 (N_21672,N_21471,N_20483);
xor U21673 (N_21673,N_21233,N_21480);
nor U21674 (N_21674,N_21132,N_20989);
and U21675 (N_21675,N_20755,N_21009);
or U21676 (N_21676,N_20964,N_20900);
nand U21677 (N_21677,N_21230,N_20957);
nand U21678 (N_21678,N_20811,N_21051);
or U21679 (N_21679,N_21213,N_20615);
and U21680 (N_21680,N_21560,N_21412);
and U21681 (N_21681,N_20756,N_21206);
and U21682 (N_21682,N_20592,N_20595);
nor U21683 (N_21683,N_20525,N_20859);
and U21684 (N_21684,N_20959,N_21226);
nor U21685 (N_21685,N_21353,N_20649);
or U21686 (N_21686,N_20737,N_21175);
nor U21687 (N_21687,N_20939,N_20998);
nor U21688 (N_21688,N_21478,N_20541);
nor U21689 (N_21689,N_20774,N_20687);
nor U21690 (N_21690,N_20951,N_20586);
and U21691 (N_21691,N_21077,N_20406);
or U21692 (N_21692,N_21144,N_20976);
nor U21693 (N_21693,N_21450,N_21382);
nor U21694 (N_21694,N_21222,N_20689);
nor U21695 (N_21695,N_21442,N_21492);
or U21696 (N_21696,N_21097,N_21153);
and U21697 (N_21697,N_21439,N_20831);
nand U21698 (N_21698,N_21229,N_21393);
nand U21699 (N_21699,N_20955,N_20761);
nor U21700 (N_21700,N_20740,N_21210);
or U21701 (N_21701,N_20962,N_21040);
or U21702 (N_21702,N_20893,N_20558);
xor U21703 (N_21703,N_21043,N_21294);
xnor U21704 (N_21704,N_21186,N_20698);
and U21705 (N_21705,N_21044,N_20931);
xor U21706 (N_21706,N_20625,N_21377);
xnor U21707 (N_21707,N_20459,N_20975);
and U21708 (N_21708,N_21301,N_21191);
or U21709 (N_21709,N_20813,N_20999);
xor U21710 (N_21710,N_21510,N_21200);
and U21711 (N_21711,N_21334,N_21062);
xnor U21712 (N_21712,N_21588,N_20914);
and U21713 (N_21713,N_20457,N_20856);
nor U21714 (N_21714,N_21532,N_21565);
nand U21715 (N_21715,N_20709,N_20817);
nor U21716 (N_21716,N_21466,N_21372);
and U21717 (N_21717,N_21295,N_20703);
nor U21718 (N_21718,N_21537,N_21543);
xnor U21719 (N_21719,N_20575,N_21189);
nor U21720 (N_21720,N_21289,N_21100);
and U21721 (N_21721,N_20556,N_21579);
or U21722 (N_21722,N_20949,N_20510);
and U21723 (N_21723,N_21235,N_21590);
or U21724 (N_21724,N_21521,N_21061);
nand U21725 (N_21725,N_20947,N_20447);
or U21726 (N_21726,N_21032,N_20641);
nand U21727 (N_21727,N_21460,N_20554);
and U21728 (N_21728,N_20768,N_21286);
nor U21729 (N_21729,N_20477,N_20840);
nor U21730 (N_21730,N_21299,N_20659);
xor U21731 (N_21731,N_20664,N_20762);
xnor U21732 (N_21732,N_21259,N_21558);
nand U21733 (N_21733,N_21489,N_21020);
or U21734 (N_21734,N_21095,N_20436);
xnor U21735 (N_21735,N_20660,N_20861);
and U21736 (N_21736,N_20770,N_20898);
and U21737 (N_21737,N_21002,N_21239);
nor U21738 (N_21738,N_21534,N_20429);
or U21739 (N_21739,N_20852,N_20476);
xor U21740 (N_21740,N_21542,N_20973);
xor U21741 (N_21741,N_20466,N_21137);
xnor U21742 (N_21742,N_20462,N_21150);
nand U21743 (N_21743,N_21080,N_20587);
xnor U21744 (N_21744,N_20908,N_20750);
and U21745 (N_21745,N_21280,N_20555);
xor U21746 (N_21746,N_21432,N_21170);
or U21747 (N_21747,N_21296,N_20825);
and U21748 (N_21748,N_20410,N_20616);
and U21749 (N_21749,N_21261,N_20443);
nor U21750 (N_21750,N_21292,N_20430);
nor U21751 (N_21751,N_21103,N_20418);
xor U21752 (N_21752,N_21526,N_21060);
xnor U21753 (N_21753,N_21524,N_21072);
nand U21754 (N_21754,N_20469,N_21267);
nand U21755 (N_21755,N_20872,N_20456);
and U21756 (N_21756,N_20997,N_20982);
nand U21757 (N_21757,N_21525,N_21368);
and U21758 (N_21758,N_21386,N_21021);
nor U21759 (N_21759,N_20572,N_21152);
xor U21760 (N_21760,N_20468,N_21260);
nand U21761 (N_21761,N_20746,N_21523);
xnor U21762 (N_21762,N_21263,N_20552);
and U21763 (N_21763,N_21257,N_20569);
nand U21764 (N_21764,N_20452,N_21437);
or U21765 (N_21765,N_21171,N_21281);
and U21766 (N_21766,N_20417,N_20665);
xnor U21767 (N_21767,N_20857,N_20805);
or U21768 (N_21768,N_20952,N_20514);
nand U21769 (N_21769,N_21454,N_21362);
nand U21770 (N_21770,N_20919,N_20634);
nand U21771 (N_21771,N_21049,N_20645);
nor U21772 (N_21772,N_21160,N_21050);
xor U21773 (N_21773,N_20744,N_20467);
nor U21774 (N_21774,N_21384,N_21255);
or U21775 (N_21775,N_21507,N_20945);
and U21776 (N_21776,N_21586,N_21028);
nand U21777 (N_21777,N_21350,N_20930);
or U21778 (N_21778,N_20832,N_21208);
or U21779 (N_21779,N_20836,N_21004);
nor U21780 (N_21780,N_21554,N_20451);
or U21781 (N_21781,N_20557,N_20969);
nor U21782 (N_21782,N_21440,N_20935);
or U21783 (N_21783,N_21400,N_21254);
nand U21784 (N_21784,N_20699,N_20409);
nor U21785 (N_21785,N_21574,N_21158);
nor U21786 (N_21786,N_21127,N_20604);
nand U21787 (N_21787,N_21277,N_21402);
xor U21788 (N_21788,N_21056,N_20530);
and U21789 (N_21789,N_20714,N_21441);
nand U21790 (N_21790,N_20797,N_21395);
or U21791 (N_21791,N_21433,N_20482);
xnor U21792 (N_21792,N_20784,N_20772);
or U21793 (N_21793,N_20669,N_21529);
xor U21794 (N_21794,N_20666,N_20591);
nand U21795 (N_21795,N_20895,N_20523);
and U21796 (N_21796,N_20985,N_21539);
or U21797 (N_21797,N_20424,N_21573);
nor U21798 (N_21798,N_20734,N_20433);
nand U21799 (N_21799,N_21057,N_20759);
and U21800 (N_21800,N_20423,N_20745);
and U21801 (N_21801,N_20420,N_21317);
or U21802 (N_21802,N_21348,N_20782);
and U21803 (N_21803,N_20879,N_21135);
or U21804 (N_21804,N_20578,N_20495);
or U21805 (N_21805,N_21130,N_20606);
nand U21806 (N_21806,N_21066,N_21092);
nor U21807 (N_21807,N_20620,N_20932);
and U21808 (N_21808,N_20674,N_21346);
and U21809 (N_21809,N_20455,N_20594);
and U21810 (N_21810,N_20925,N_20583);
nor U21811 (N_21811,N_21145,N_21398);
nand U21812 (N_21812,N_20922,N_21283);
nor U21813 (N_21813,N_20504,N_21587);
nand U21814 (N_21814,N_20635,N_20501);
and U21815 (N_21815,N_21462,N_20695);
xor U21816 (N_21816,N_20512,N_20521);
nand U21817 (N_21817,N_20639,N_20403);
nor U21818 (N_21818,N_21594,N_20642);
or U21819 (N_21819,N_21376,N_20878);
nor U21820 (N_21820,N_21564,N_21107);
and U21821 (N_21821,N_20499,N_21287);
xor U21822 (N_21822,N_21085,N_20640);
nand U21823 (N_21823,N_21447,N_21332);
nor U21824 (N_21824,N_20562,N_20497);
or U21825 (N_21825,N_21123,N_20623);
nor U21826 (N_21826,N_21330,N_21355);
and U21827 (N_21827,N_21065,N_21250);
nor U21828 (N_21828,N_20763,N_21503);
nand U21829 (N_21829,N_21262,N_21363);
or U21830 (N_21830,N_21513,N_21344);
or U21831 (N_21831,N_20413,N_21530);
or U21832 (N_21832,N_20405,N_20799);
nor U21833 (N_21833,N_21165,N_21018);
or U21834 (N_21834,N_21220,N_21465);
or U21835 (N_21835,N_20540,N_21008);
or U21836 (N_21836,N_20771,N_20702);
and U21837 (N_21837,N_21010,N_21464);
or U21838 (N_21838,N_20445,N_21570);
or U21839 (N_21839,N_20789,N_20723);
and U21840 (N_21840,N_20685,N_21577);
and U21841 (N_21841,N_21509,N_20883);
xnor U21842 (N_21842,N_21197,N_20400);
and U21843 (N_21843,N_20524,N_21114);
nand U21844 (N_21844,N_21048,N_21426);
nor U21845 (N_21845,N_20897,N_21316);
xnor U21846 (N_21846,N_21248,N_21096);
nor U21847 (N_21847,N_21364,N_20605);
or U21848 (N_21848,N_20830,N_20614);
nand U21849 (N_21849,N_20478,N_21598);
xnor U21850 (N_21850,N_20672,N_20713);
or U21851 (N_21851,N_20630,N_21052);
or U21852 (N_21852,N_21185,N_20864);
nand U21853 (N_21853,N_21544,N_20663);
nor U21854 (N_21854,N_20688,N_21265);
nand U21855 (N_21855,N_20736,N_20580);
xor U21856 (N_21856,N_20600,N_20471);
xor U21857 (N_21857,N_20958,N_20570);
nor U21858 (N_21858,N_21205,N_21027);
nand U21859 (N_21859,N_21580,N_20566);
nor U21860 (N_21860,N_20779,N_20657);
nand U21861 (N_21861,N_21493,N_21428);
nand U21862 (N_21862,N_21394,N_21136);
nor U21863 (N_21863,N_20911,N_21467);
xor U21864 (N_21864,N_21309,N_21249);
nand U21865 (N_21865,N_21117,N_20511);
nor U21866 (N_21866,N_21340,N_20590);
and U21867 (N_21867,N_20896,N_21176);
or U21868 (N_21868,N_21418,N_21427);
xnor U21869 (N_21869,N_20778,N_20636);
xnor U21870 (N_21870,N_20754,N_20676);
and U21871 (N_21871,N_20967,N_21474);
and U21872 (N_21872,N_20553,N_20991);
and U21873 (N_21873,N_21169,N_21319);
or U21874 (N_21874,N_21475,N_21354);
xor U21875 (N_21875,N_21241,N_20576);
xnor U21876 (N_21876,N_20439,N_21108);
and U21877 (N_21877,N_20937,N_21396);
nor U21878 (N_21878,N_20970,N_20464);
nor U21879 (N_21879,N_20800,N_20823);
nor U21880 (N_21880,N_21487,N_20598);
and U21881 (N_21881,N_21499,N_21068);
xnor U21882 (N_21882,N_20682,N_21228);
and U21883 (N_21883,N_21279,N_20795);
nand U21884 (N_21884,N_21172,N_20419);
and U21885 (N_21885,N_20473,N_21552);
xnor U21886 (N_21886,N_20727,N_21154);
nand U21887 (N_21887,N_21511,N_20865);
or U21888 (N_21888,N_21023,N_21387);
nand U21889 (N_21889,N_21383,N_20520);
xnor U21890 (N_21890,N_20902,N_21408);
nand U21891 (N_21891,N_21436,N_21266);
nand U21892 (N_21892,N_20481,N_20757);
xor U21893 (N_21893,N_20882,N_21358);
and U21894 (N_21894,N_20426,N_20547);
and U21895 (N_21895,N_21124,N_20712);
and U21896 (N_21896,N_21029,N_20602);
and U21897 (N_21897,N_20559,N_21452);
nand U21898 (N_21898,N_21514,N_20974);
or U21899 (N_21899,N_20487,N_21360);
and U21900 (N_21900,N_21578,N_20928);
xnor U21901 (N_21901,N_20815,N_20758);
xor U21902 (N_21902,N_21270,N_20769);
and U21903 (N_21903,N_21519,N_21391);
nand U21904 (N_21904,N_21335,N_20934);
and U21905 (N_21905,N_20792,N_20608);
and U21906 (N_21906,N_21438,N_21128);
nand U21907 (N_21907,N_21063,N_21151);
or U21908 (N_21908,N_20638,N_20412);
nand U21909 (N_21909,N_20596,N_20916);
nand U21910 (N_21910,N_20573,N_21506);
or U21911 (N_21911,N_20866,N_20804);
xor U21912 (N_21912,N_20619,N_21225);
or U21913 (N_21913,N_21435,N_21297);
nand U21914 (N_21914,N_21484,N_21274);
xor U21915 (N_21915,N_20867,N_21392);
nor U21916 (N_21916,N_20993,N_20818);
nor U21917 (N_21917,N_20472,N_21424);
nand U21918 (N_21918,N_20599,N_21517);
and U21919 (N_21919,N_21352,N_20700);
or U21920 (N_21920,N_21174,N_21141);
or U21921 (N_21921,N_21099,N_21385);
xnor U21922 (N_21922,N_20936,N_21568);
or U21923 (N_21923,N_20858,N_20678);
and U21924 (N_21924,N_21268,N_20465);
nand U21925 (N_21925,N_20777,N_20905);
and U21926 (N_21926,N_21113,N_20903);
and U21927 (N_21927,N_21237,N_21247);
nand U21928 (N_21928,N_20906,N_21563);
nand U21929 (N_21929,N_20503,N_20446);
or U21930 (N_21930,N_21419,N_21498);
or U21931 (N_21931,N_21074,N_20438);
nand U21932 (N_21932,N_20942,N_21015);
and U21933 (N_21933,N_21118,N_20968);
or U21934 (N_21934,N_21000,N_20629);
or U21935 (N_21935,N_20593,N_21411);
nor U21936 (N_21936,N_21025,N_21047);
xor U21937 (N_21937,N_20536,N_20855);
nand U21938 (N_21938,N_21311,N_21444);
xor U21939 (N_21939,N_20621,N_20924);
xor U21940 (N_21940,N_21147,N_20581);
and U21941 (N_21941,N_21320,N_20577);
nand U21942 (N_21942,N_21199,N_20860);
or U21943 (N_21943,N_21177,N_21504);
and U21944 (N_21944,N_21420,N_20884);
or U21945 (N_21945,N_20627,N_20721);
nand U21946 (N_21946,N_21304,N_21219);
and U21947 (N_21947,N_20851,N_21349);
or U21948 (N_21948,N_20509,N_20507);
nand U21949 (N_21949,N_20474,N_21388);
nor U21950 (N_21950,N_20527,N_21518);
and U21951 (N_21951,N_21139,N_20885);
and U21952 (N_21952,N_21496,N_21318);
and U21953 (N_21953,N_21216,N_20532);
and U21954 (N_21954,N_20827,N_21059);
xnor U21955 (N_21955,N_21331,N_20546);
or U21956 (N_21956,N_20519,N_21203);
nand U21957 (N_21957,N_20652,N_20953);
or U21958 (N_21958,N_20416,N_20693);
nor U21959 (N_21959,N_20901,N_20613);
nand U21960 (N_21960,N_20506,N_20571);
or U21961 (N_21961,N_20644,N_21535);
nand U21962 (N_21962,N_20978,N_21202);
or U21963 (N_21963,N_20480,N_21581);
nand U21964 (N_21964,N_20835,N_21278);
and U21965 (N_21965,N_20876,N_21365);
nor U21966 (N_21966,N_20711,N_20491);
nand U21967 (N_21967,N_21035,N_20516);
or U21968 (N_21968,N_20539,N_20839);
nand U21969 (N_21969,N_20708,N_20407);
or U21970 (N_21970,N_20802,N_20425);
or U21971 (N_21971,N_21161,N_20716);
xnor U21972 (N_21972,N_21562,N_20496);
xor U21973 (N_21973,N_20749,N_20829);
nand U21974 (N_21974,N_20565,N_20984);
and U21975 (N_21975,N_21183,N_21491);
and U21976 (N_21976,N_20943,N_21561);
and U21977 (N_21977,N_20414,N_21264);
nand U21978 (N_21978,N_21131,N_21389);
nor U21979 (N_21979,N_21459,N_21538);
or U21980 (N_21980,N_20828,N_20441);
xnor U21981 (N_21981,N_21589,N_21553);
nor U21982 (N_21982,N_21019,N_21178);
nor U21983 (N_21983,N_20886,N_20461);
and U21984 (N_21984,N_21592,N_20513);
nor U21985 (N_21985,N_21307,N_21194);
or U21986 (N_21986,N_20428,N_20498);
and U21987 (N_21987,N_20637,N_21343);
xor U21988 (N_21988,N_20564,N_21227);
nor U21989 (N_21989,N_21033,N_20515);
nand U21990 (N_21990,N_20977,N_20574);
or U21991 (N_21991,N_21067,N_20551);
xor U21992 (N_21992,N_20500,N_21236);
and U21993 (N_21993,N_20545,N_20651);
nand U21994 (N_21994,N_21505,N_21490);
xor U21995 (N_21995,N_21276,N_20485);
xor U21996 (N_21996,N_21324,N_21234);
xnor U21997 (N_21997,N_21179,N_20579);
and U21998 (N_21998,N_20820,N_21423);
xor U21999 (N_21999,N_21039,N_21541);
nor U22000 (N_22000,N_20875,N_21315);
and U22001 (N_22001,N_21597,N_21163);
and U22002 (N_22002,N_21162,N_21356);
nand U22003 (N_22003,N_21546,N_21058);
or U22004 (N_22004,N_21181,N_20992);
or U22005 (N_22005,N_20508,N_21109);
nor U22006 (N_22006,N_20869,N_20624);
and U22007 (N_22007,N_21421,N_21173);
nor U22008 (N_22008,N_21007,N_21374);
xnor U22009 (N_22009,N_20728,N_21409);
nor U22010 (N_22010,N_21105,N_20449);
and U22011 (N_22011,N_21456,N_21457);
xnor U22012 (N_22012,N_21429,N_21143);
and U22013 (N_22013,N_20611,N_20788);
xor U22014 (N_22014,N_21218,N_20612);
nand U22015 (N_22015,N_20739,N_20486);
nand U22016 (N_22016,N_21306,N_20494);
and U22017 (N_22017,N_20790,N_20785);
nand U22018 (N_22018,N_20518,N_20718);
and U22019 (N_22019,N_21333,N_20568);
and U22020 (N_22020,N_21403,N_20888);
xnor U22021 (N_22021,N_21271,N_21221);
nor U22022 (N_22022,N_21599,N_20724);
nor U22023 (N_22023,N_20720,N_20563);
xor U22024 (N_22024,N_21157,N_21038);
or U22025 (N_22025,N_20950,N_20929);
and U22026 (N_22026,N_21006,N_21341);
xor U22027 (N_22027,N_21090,N_21572);
xnor U22028 (N_22028,N_21593,N_20582);
xor U22029 (N_22029,N_21187,N_20460);
xnor U22030 (N_22030,N_20921,N_20824);
nand U22031 (N_22031,N_21275,N_20912);
and U22032 (N_22032,N_21325,N_21016);
nor U22033 (N_22033,N_20892,N_20526);
and U22034 (N_22034,N_20738,N_20767);
or U22035 (N_22035,N_21373,N_20691);
xnor U22036 (N_22036,N_21375,N_21003);
xor U22037 (N_22037,N_20956,N_20490);
and U22038 (N_22038,N_20470,N_20656);
xor U22039 (N_22039,N_20809,N_21576);
and U22040 (N_22040,N_21217,N_20783);
xnor U22041 (N_22041,N_21468,N_20853);
nand U22042 (N_22042,N_20534,N_20673);
xor U22043 (N_22043,N_20444,N_21196);
xnor U22044 (N_22044,N_21326,N_21001);
and U22045 (N_22045,N_21070,N_21104);
or U22046 (N_22046,N_21555,N_20747);
nor U22047 (N_22047,N_20647,N_21321);
nand U22048 (N_22048,N_21076,N_20941);
xor U22049 (N_22049,N_20654,N_21167);
and U22050 (N_22050,N_20522,N_21528);
nand U22051 (N_22051,N_20458,N_21479);
xnor U22052 (N_22052,N_20775,N_21508);
nor U22053 (N_22053,N_20781,N_21240);
or U22054 (N_22054,N_20662,N_20628);
and U22055 (N_22055,N_21138,N_20401);
xor U22056 (N_22056,N_21458,N_20655);
nand U22057 (N_22057,N_21431,N_21556);
or U22058 (N_22058,N_20848,N_21146);
or U22059 (N_22059,N_21238,N_20528);
xnor U22060 (N_22060,N_21055,N_20432);
xnor U22061 (N_22061,N_20909,N_20692);
or U22062 (N_22062,N_20933,N_20675);
xor U22063 (N_22063,N_20972,N_21536);
xnor U22064 (N_22064,N_20963,N_21486);
or U22065 (N_22065,N_20732,N_21406);
nor U22066 (N_22066,N_21091,N_21322);
nor U22067 (N_22067,N_20983,N_20543);
or U22068 (N_22068,N_20729,N_21129);
xor U22069 (N_22069,N_21367,N_20697);
nor U22070 (N_22070,N_21443,N_20646);
nand U22071 (N_22071,N_20760,N_20881);
and U22072 (N_22072,N_21584,N_20434);
nand U22073 (N_22073,N_21084,N_20987);
and U22074 (N_22074,N_21209,N_20948);
xnor U22075 (N_22075,N_21045,N_21488);
nor U22076 (N_22076,N_21461,N_21211);
xnor U22077 (N_22077,N_21342,N_21300);
and U22078 (N_22078,N_21328,N_20752);
and U22079 (N_22079,N_21246,N_21313);
nor U22080 (N_22080,N_20411,N_20427);
and U22081 (N_22081,N_20585,N_20743);
nor U22082 (N_22082,N_21527,N_20965);
and U22083 (N_22083,N_20786,N_20742);
or U22084 (N_22084,N_20661,N_20535);
and U22085 (N_22085,N_21399,N_21011);
xnor U22086 (N_22086,N_21453,N_21030);
or U22087 (N_22087,N_21164,N_20431);
nand U22088 (N_22088,N_21451,N_20588);
and U22089 (N_22089,N_21232,N_20880);
and U22090 (N_22090,N_20807,N_21339);
or U22091 (N_22091,N_20845,N_20994);
and U22092 (N_22092,N_21404,N_20560);
nor U22093 (N_22093,N_20821,N_20960);
nor U22094 (N_22094,N_21381,N_20838);
nand U22095 (N_22095,N_20440,N_20773);
and U22096 (N_22096,N_21540,N_21188);
nor U22097 (N_22097,N_20981,N_21502);
nor U22098 (N_22098,N_20806,N_21291);
nor U22099 (N_22099,N_20653,N_21416);
nand U22100 (N_22100,N_20990,N_21378);
xor U22101 (N_22101,N_21148,N_21122);
nand U22102 (N_22102,N_21359,N_21351);
nand U22103 (N_22103,N_21422,N_21252);
or U22104 (N_22104,N_21345,N_21223);
xor U22105 (N_22105,N_21482,N_20940);
or U22106 (N_22106,N_20415,N_20834);
nand U22107 (N_22107,N_20537,N_20658);
and U22108 (N_22108,N_20910,N_21481);
nor U22109 (N_22109,N_21193,N_20696);
and U22110 (N_22110,N_21110,N_21582);
nand U22111 (N_22111,N_20816,N_21116);
or U22112 (N_22112,N_20609,N_21140);
nand U22113 (N_22113,N_21559,N_20918);
nor U22114 (N_22114,N_20589,N_20448);
nor U22115 (N_22115,N_20633,N_20741);
and U22116 (N_22116,N_21251,N_21455);
xnor U22117 (N_22117,N_20849,N_20463);
xor U22118 (N_22118,N_21415,N_21005);
nor U22119 (N_22119,N_21430,N_21583);
or U22120 (N_22120,N_20686,N_21545);
and U22121 (N_22121,N_21184,N_20725);
and U22122 (N_22122,N_20442,N_20681);
xor U22123 (N_22123,N_21046,N_20505);
nand U22124 (N_22124,N_20873,N_20622);
and U22125 (N_22125,N_20643,N_21198);
xnor U22126 (N_22126,N_20913,N_21533);
nor U22127 (N_22127,N_21272,N_20618);
nand U22128 (N_22128,N_20717,N_20707);
or U22129 (N_22129,N_21142,N_20748);
nor U22130 (N_22130,N_21347,N_21064);
xor U22131 (N_22131,N_20670,N_20961);
and U22132 (N_22132,N_21155,N_20479);
and U22133 (N_22133,N_20843,N_21017);
and U22134 (N_22134,N_20826,N_20787);
xnor U22135 (N_22135,N_20938,N_20475);
and U22136 (N_22136,N_21566,N_21166);
xor U22137 (N_22137,N_21120,N_20819);
or U22138 (N_22138,N_20715,N_21314);
or U22139 (N_22139,N_21098,N_20891);
and U22140 (N_22140,N_20907,N_20544);
xnor U22141 (N_22141,N_21585,N_20842);
or U22142 (N_22142,N_20917,N_21089);
xnor U22143 (N_22143,N_21042,N_20517);
or U22144 (N_22144,N_20780,N_21449);
nand U22145 (N_22145,N_21405,N_21366);
and U22146 (N_22146,N_20542,N_20453);
and U22147 (N_22147,N_20719,N_21026);
or U22148 (N_22148,N_20837,N_20607);
nand U22149 (N_22149,N_20680,N_21022);
or U22150 (N_22150,N_21134,N_21371);
or U22151 (N_22151,N_20844,N_21417);
or U22152 (N_22152,N_20631,N_20887);
nor U22153 (N_22153,N_20847,N_20926);
and U22154 (N_22154,N_20531,N_20731);
xor U22155 (N_22155,N_20671,N_21269);
nor U22156 (N_22156,N_21207,N_21086);
xor U22157 (N_22157,N_21470,N_21231);
and U22158 (N_22158,N_20890,N_20814);
and U22159 (N_22159,N_20422,N_20794);
xor U22160 (N_22160,N_20751,N_20421);
or U22161 (N_22161,N_21483,N_21037);
xor U22162 (N_22162,N_21012,N_21370);
xor U22163 (N_22163,N_20877,N_21476);
nand U22164 (N_22164,N_20450,N_20617);
xnor U22165 (N_22165,N_21407,N_20489);
nor U22166 (N_22166,N_21094,N_21168);
and U22167 (N_22167,N_21380,N_21327);
and U22168 (N_22168,N_20454,N_21182);
nor U22169 (N_22169,N_20626,N_20946);
and U22170 (N_22170,N_21214,N_21243);
xor U22171 (N_22171,N_21497,N_21531);
and U22172 (N_22172,N_21053,N_21081);
nand U22173 (N_22173,N_20871,N_20597);
xnor U22174 (N_22174,N_20920,N_21041);
nor U22175 (N_22175,N_21310,N_20904);
or U22176 (N_22176,N_20954,N_20603);
and U22177 (N_22177,N_20846,N_21550);
or U22178 (N_22178,N_21156,N_20704);
nor U22179 (N_22179,N_20995,N_21036);
nor U22180 (N_22180,N_20701,N_20944);
nand U22181 (N_22181,N_20567,N_21054);
and U22182 (N_22182,N_20533,N_21557);
nand U22183 (N_22183,N_20484,N_21338);
nand U22184 (N_22184,N_20766,N_21126);
nor U22185 (N_22185,N_20923,N_21512);
nor U22186 (N_22186,N_20677,N_20679);
or U22187 (N_22187,N_20502,N_21308);
nand U22188 (N_22188,N_20966,N_20492);
and U22189 (N_22189,N_20668,N_20915);
and U22190 (N_22190,N_21078,N_20667);
and U22191 (N_22191,N_21087,N_21102);
nand U22192 (N_22192,N_20561,N_20971);
and U22193 (N_22193,N_20632,N_21500);
and U22194 (N_22194,N_21473,N_21293);
nor U22195 (N_22195,N_21204,N_21201);
or U22196 (N_22196,N_21075,N_20822);
nor U22197 (N_22197,N_21522,N_21215);
nor U22198 (N_22198,N_20402,N_20765);
nand U22199 (N_22199,N_20988,N_20791);
nor U22200 (N_22200,N_20481,N_20812);
and U22201 (N_22201,N_20660,N_21109);
and U22202 (N_22202,N_20799,N_21421);
or U22203 (N_22203,N_21274,N_21082);
nand U22204 (N_22204,N_21497,N_21066);
xor U22205 (N_22205,N_20474,N_20629);
or U22206 (N_22206,N_20406,N_20796);
nand U22207 (N_22207,N_20450,N_21344);
and U22208 (N_22208,N_20643,N_20512);
xor U22209 (N_22209,N_21407,N_21421);
xnor U22210 (N_22210,N_21035,N_21340);
nand U22211 (N_22211,N_21155,N_20935);
nor U22212 (N_22212,N_20791,N_21306);
nand U22213 (N_22213,N_20418,N_21590);
nor U22214 (N_22214,N_20681,N_20778);
nor U22215 (N_22215,N_20811,N_21475);
xnor U22216 (N_22216,N_20535,N_21120);
and U22217 (N_22217,N_20876,N_21076);
and U22218 (N_22218,N_21163,N_20629);
and U22219 (N_22219,N_20510,N_21400);
nand U22220 (N_22220,N_21074,N_21035);
nand U22221 (N_22221,N_21067,N_21491);
xor U22222 (N_22222,N_20484,N_21185);
and U22223 (N_22223,N_20553,N_21138);
nor U22224 (N_22224,N_20980,N_20596);
nor U22225 (N_22225,N_20479,N_21348);
nand U22226 (N_22226,N_20769,N_20494);
or U22227 (N_22227,N_20474,N_20880);
or U22228 (N_22228,N_21233,N_20629);
xor U22229 (N_22229,N_20509,N_21174);
nand U22230 (N_22230,N_20501,N_20755);
and U22231 (N_22231,N_21449,N_20663);
nand U22232 (N_22232,N_20416,N_21158);
nand U22233 (N_22233,N_20602,N_21190);
nor U22234 (N_22234,N_21392,N_20721);
xnor U22235 (N_22235,N_20888,N_21549);
or U22236 (N_22236,N_21023,N_20897);
nor U22237 (N_22237,N_21035,N_21022);
nand U22238 (N_22238,N_21207,N_20860);
xor U22239 (N_22239,N_21471,N_20680);
xnor U22240 (N_22240,N_20877,N_20705);
and U22241 (N_22241,N_20739,N_21112);
or U22242 (N_22242,N_21195,N_21366);
nand U22243 (N_22243,N_21496,N_20813);
and U22244 (N_22244,N_20409,N_21284);
or U22245 (N_22245,N_21489,N_20820);
xor U22246 (N_22246,N_20661,N_20879);
nand U22247 (N_22247,N_20740,N_20862);
nand U22248 (N_22248,N_20409,N_20949);
nor U22249 (N_22249,N_20636,N_21418);
and U22250 (N_22250,N_21178,N_20497);
and U22251 (N_22251,N_20690,N_21136);
nor U22252 (N_22252,N_20743,N_21529);
xor U22253 (N_22253,N_21280,N_20489);
xor U22254 (N_22254,N_21522,N_20418);
or U22255 (N_22255,N_20870,N_20446);
nor U22256 (N_22256,N_20444,N_20517);
xor U22257 (N_22257,N_20746,N_20772);
nand U22258 (N_22258,N_20856,N_20525);
nand U22259 (N_22259,N_21438,N_21491);
or U22260 (N_22260,N_20694,N_20678);
nand U22261 (N_22261,N_20834,N_20815);
or U22262 (N_22262,N_20910,N_21302);
and U22263 (N_22263,N_21219,N_21309);
or U22264 (N_22264,N_20412,N_20728);
and U22265 (N_22265,N_21175,N_21123);
nor U22266 (N_22266,N_21152,N_20905);
nor U22267 (N_22267,N_20491,N_20547);
xor U22268 (N_22268,N_21347,N_21492);
and U22269 (N_22269,N_21591,N_20535);
nor U22270 (N_22270,N_20742,N_21478);
nor U22271 (N_22271,N_21349,N_20433);
and U22272 (N_22272,N_20625,N_20487);
or U22273 (N_22273,N_21169,N_20599);
nand U22274 (N_22274,N_20994,N_21329);
xor U22275 (N_22275,N_20864,N_21474);
nor U22276 (N_22276,N_21068,N_21332);
and U22277 (N_22277,N_20564,N_21169);
nor U22278 (N_22278,N_21501,N_21156);
or U22279 (N_22279,N_21051,N_20580);
or U22280 (N_22280,N_21466,N_21072);
nand U22281 (N_22281,N_21501,N_21040);
and U22282 (N_22282,N_21156,N_20749);
and U22283 (N_22283,N_20827,N_21340);
xnor U22284 (N_22284,N_21160,N_21549);
or U22285 (N_22285,N_21056,N_20988);
xor U22286 (N_22286,N_20888,N_20886);
nand U22287 (N_22287,N_20698,N_20726);
nand U22288 (N_22288,N_21352,N_20606);
nand U22289 (N_22289,N_21199,N_20941);
or U22290 (N_22290,N_21003,N_20619);
or U22291 (N_22291,N_21210,N_21585);
xnor U22292 (N_22292,N_20478,N_20528);
or U22293 (N_22293,N_20929,N_20873);
nor U22294 (N_22294,N_21429,N_21369);
or U22295 (N_22295,N_21405,N_21185);
and U22296 (N_22296,N_20632,N_21593);
xnor U22297 (N_22297,N_21382,N_21485);
and U22298 (N_22298,N_21585,N_20738);
or U22299 (N_22299,N_21245,N_20481);
and U22300 (N_22300,N_21328,N_20733);
or U22301 (N_22301,N_21261,N_20696);
and U22302 (N_22302,N_21152,N_20885);
or U22303 (N_22303,N_21195,N_20838);
or U22304 (N_22304,N_21323,N_20867);
nor U22305 (N_22305,N_20496,N_20438);
and U22306 (N_22306,N_21493,N_21020);
xor U22307 (N_22307,N_21300,N_20731);
xor U22308 (N_22308,N_21267,N_21350);
or U22309 (N_22309,N_20474,N_20941);
nor U22310 (N_22310,N_20789,N_21457);
nand U22311 (N_22311,N_21324,N_20820);
or U22312 (N_22312,N_20874,N_21471);
and U22313 (N_22313,N_21115,N_20951);
nor U22314 (N_22314,N_20794,N_20485);
and U22315 (N_22315,N_20455,N_20523);
xor U22316 (N_22316,N_20482,N_20652);
or U22317 (N_22317,N_21325,N_20752);
nor U22318 (N_22318,N_21157,N_21356);
xor U22319 (N_22319,N_20863,N_21494);
and U22320 (N_22320,N_20539,N_21076);
nor U22321 (N_22321,N_20482,N_21004);
nand U22322 (N_22322,N_20520,N_21208);
xor U22323 (N_22323,N_20739,N_21134);
nor U22324 (N_22324,N_21585,N_21356);
and U22325 (N_22325,N_21345,N_21158);
xor U22326 (N_22326,N_21165,N_21581);
nor U22327 (N_22327,N_20859,N_20986);
and U22328 (N_22328,N_20491,N_20593);
nand U22329 (N_22329,N_20975,N_21444);
or U22330 (N_22330,N_20463,N_20874);
nor U22331 (N_22331,N_21578,N_21428);
or U22332 (N_22332,N_20843,N_20737);
nor U22333 (N_22333,N_20486,N_20670);
nand U22334 (N_22334,N_21023,N_21599);
nor U22335 (N_22335,N_20966,N_21464);
and U22336 (N_22336,N_20709,N_20726);
nand U22337 (N_22337,N_21184,N_20762);
or U22338 (N_22338,N_21516,N_21525);
or U22339 (N_22339,N_21486,N_20696);
nor U22340 (N_22340,N_20785,N_21363);
or U22341 (N_22341,N_20634,N_21186);
or U22342 (N_22342,N_20528,N_20790);
xnor U22343 (N_22343,N_21410,N_21534);
or U22344 (N_22344,N_21266,N_20421);
or U22345 (N_22345,N_21056,N_21029);
nor U22346 (N_22346,N_20473,N_21342);
nor U22347 (N_22347,N_21544,N_20565);
nand U22348 (N_22348,N_21284,N_21467);
xor U22349 (N_22349,N_21346,N_21341);
and U22350 (N_22350,N_20981,N_21423);
nand U22351 (N_22351,N_20636,N_21318);
and U22352 (N_22352,N_21451,N_21148);
nor U22353 (N_22353,N_21347,N_21089);
nor U22354 (N_22354,N_21072,N_21376);
and U22355 (N_22355,N_20984,N_20545);
or U22356 (N_22356,N_21044,N_20478);
nor U22357 (N_22357,N_20615,N_20544);
nor U22358 (N_22358,N_20429,N_20704);
nor U22359 (N_22359,N_20473,N_20663);
or U22360 (N_22360,N_21234,N_21275);
nor U22361 (N_22361,N_21021,N_20639);
nor U22362 (N_22362,N_21387,N_21191);
xnor U22363 (N_22363,N_20729,N_20956);
xnor U22364 (N_22364,N_21263,N_21044);
nand U22365 (N_22365,N_21495,N_20639);
xor U22366 (N_22366,N_21016,N_20405);
or U22367 (N_22367,N_20725,N_21131);
nand U22368 (N_22368,N_20766,N_21533);
xor U22369 (N_22369,N_20518,N_21170);
and U22370 (N_22370,N_21073,N_21251);
nor U22371 (N_22371,N_20974,N_21182);
nand U22372 (N_22372,N_20495,N_21024);
nand U22373 (N_22373,N_20858,N_21364);
nor U22374 (N_22374,N_20782,N_20509);
xnor U22375 (N_22375,N_20686,N_21370);
nor U22376 (N_22376,N_20912,N_21520);
and U22377 (N_22377,N_20470,N_21371);
xor U22378 (N_22378,N_21242,N_21570);
xor U22379 (N_22379,N_20862,N_21449);
and U22380 (N_22380,N_20605,N_21051);
nor U22381 (N_22381,N_21140,N_21537);
or U22382 (N_22382,N_20882,N_20689);
nand U22383 (N_22383,N_20489,N_21380);
nor U22384 (N_22384,N_21589,N_21073);
xor U22385 (N_22385,N_21367,N_20786);
xor U22386 (N_22386,N_20641,N_21125);
nor U22387 (N_22387,N_21553,N_20567);
nand U22388 (N_22388,N_20704,N_20554);
nor U22389 (N_22389,N_21122,N_20861);
nand U22390 (N_22390,N_21122,N_21323);
xor U22391 (N_22391,N_21496,N_21088);
nor U22392 (N_22392,N_21360,N_20894);
or U22393 (N_22393,N_20933,N_20544);
or U22394 (N_22394,N_21194,N_21490);
nor U22395 (N_22395,N_20564,N_21216);
nor U22396 (N_22396,N_21183,N_20653);
or U22397 (N_22397,N_20402,N_21083);
nor U22398 (N_22398,N_21407,N_21293);
and U22399 (N_22399,N_21183,N_21105);
xnor U22400 (N_22400,N_21540,N_21468);
and U22401 (N_22401,N_20523,N_21075);
nor U22402 (N_22402,N_20894,N_20858);
xor U22403 (N_22403,N_20619,N_20838);
xnor U22404 (N_22404,N_21107,N_20450);
or U22405 (N_22405,N_21538,N_21278);
and U22406 (N_22406,N_21221,N_20896);
nor U22407 (N_22407,N_20799,N_21361);
or U22408 (N_22408,N_21106,N_20491);
and U22409 (N_22409,N_21119,N_20438);
nand U22410 (N_22410,N_20687,N_20670);
nor U22411 (N_22411,N_20605,N_20940);
xor U22412 (N_22412,N_21349,N_20861);
nand U22413 (N_22413,N_20482,N_21018);
xnor U22414 (N_22414,N_21172,N_20605);
and U22415 (N_22415,N_20761,N_21140);
or U22416 (N_22416,N_21282,N_21391);
nand U22417 (N_22417,N_20634,N_21126);
nor U22418 (N_22418,N_20692,N_21196);
nand U22419 (N_22419,N_21041,N_21452);
nand U22420 (N_22420,N_21295,N_20962);
or U22421 (N_22421,N_20448,N_21431);
nand U22422 (N_22422,N_21476,N_21336);
and U22423 (N_22423,N_20592,N_20622);
or U22424 (N_22424,N_21200,N_20945);
xor U22425 (N_22425,N_21002,N_21121);
nor U22426 (N_22426,N_20819,N_21121);
nand U22427 (N_22427,N_21475,N_21566);
nor U22428 (N_22428,N_21428,N_20569);
or U22429 (N_22429,N_20690,N_20436);
or U22430 (N_22430,N_21486,N_20700);
xnor U22431 (N_22431,N_21260,N_20817);
nor U22432 (N_22432,N_21237,N_20536);
xor U22433 (N_22433,N_20780,N_20491);
or U22434 (N_22434,N_21061,N_20852);
or U22435 (N_22435,N_20478,N_21272);
and U22436 (N_22436,N_21332,N_21248);
and U22437 (N_22437,N_20428,N_20647);
or U22438 (N_22438,N_20940,N_20955);
nor U22439 (N_22439,N_21318,N_20596);
xor U22440 (N_22440,N_21103,N_21167);
or U22441 (N_22441,N_21453,N_21442);
nand U22442 (N_22442,N_20702,N_20633);
nand U22443 (N_22443,N_21583,N_21396);
or U22444 (N_22444,N_21353,N_21410);
xnor U22445 (N_22445,N_21302,N_21351);
xnor U22446 (N_22446,N_21167,N_20816);
nor U22447 (N_22447,N_21310,N_21554);
or U22448 (N_22448,N_21469,N_21269);
nor U22449 (N_22449,N_21165,N_21431);
nand U22450 (N_22450,N_21420,N_20494);
or U22451 (N_22451,N_21110,N_21476);
nor U22452 (N_22452,N_21506,N_20540);
nand U22453 (N_22453,N_20697,N_21479);
nor U22454 (N_22454,N_21209,N_20702);
xnor U22455 (N_22455,N_21328,N_21584);
xor U22456 (N_22456,N_20435,N_21315);
and U22457 (N_22457,N_21540,N_20939);
or U22458 (N_22458,N_21002,N_20532);
nand U22459 (N_22459,N_20569,N_21390);
or U22460 (N_22460,N_20472,N_20660);
nor U22461 (N_22461,N_21589,N_20603);
nor U22462 (N_22462,N_20777,N_20798);
nor U22463 (N_22463,N_20555,N_21223);
nand U22464 (N_22464,N_20860,N_20674);
xnor U22465 (N_22465,N_21473,N_21291);
and U22466 (N_22466,N_21080,N_21504);
nand U22467 (N_22467,N_20560,N_21455);
and U22468 (N_22468,N_21092,N_21511);
nor U22469 (N_22469,N_20738,N_20475);
or U22470 (N_22470,N_20499,N_20516);
nor U22471 (N_22471,N_21151,N_20718);
nor U22472 (N_22472,N_20734,N_20591);
xor U22473 (N_22473,N_21271,N_20844);
nor U22474 (N_22474,N_20908,N_20767);
and U22475 (N_22475,N_20733,N_21200);
xnor U22476 (N_22476,N_21185,N_21011);
and U22477 (N_22477,N_20649,N_21388);
nor U22478 (N_22478,N_21498,N_21075);
nand U22479 (N_22479,N_21196,N_20559);
nor U22480 (N_22480,N_21533,N_20969);
nor U22481 (N_22481,N_21250,N_21567);
nand U22482 (N_22482,N_20986,N_20800);
nand U22483 (N_22483,N_21557,N_21206);
nor U22484 (N_22484,N_21116,N_20613);
and U22485 (N_22485,N_21125,N_20807);
or U22486 (N_22486,N_21049,N_20597);
nor U22487 (N_22487,N_20514,N_21314);
and U22488 (N_22488,N_20433,N_21469);
and U22489 (N_22489,N_20844,N_20826);
and U22490 (N_22490,N_20993,N_21112);
nand U22491 (N_22491,N_21401,N_21506);
and U22492 (N_22492,N_20625,N_21362);
and U22493 (N_22493,N_21193,N_21322);
xor U22494 (N_22494,N_20425,N_20840);
nor U22495 (N_22495,N_20671,N_20720);
or U22496 (N_22496,N_21071,N_21108);
xnor U22497 (N_22497,N_21054,N_20781);
nand U22498 (N_22498,N_21481,N_20647);
and U22499 (N_22499,N_20870,N_20832);
and U22500 (N_22500,N_20625,N_21572);
nor U22501 (N_22501,N_20574,N_21308);
nand U22502 (N_22502,N_21456,N_21391);
and U22503 (N_22503,N_21518,N_20494);
nor U22504 (N_22504,N_20999,N_20982);
nand U22505 (N_22505,N_21561,N_21264);
or U22506 (N_22506,N_21543,N_20519);
and U22507 (N_22507,N_21565,N_21150);
nor U22508 (N_22508,N_21588,N_20588);
nor U22509 (N_22509,N_20481,N_21120);
or U22510 (N_22510,N_21033,N_21065);
xnor U22511 (N_22511,N_20572,N_20868);
nor U22512 (N_22512,N_20423,N_21232);
xnor U22513 (N_22513,N_20844,N_21089);
nor U22514 (N_22514,N_20926,N_20764);
nor U22515 (N_22515,N_21187,N_20948);
nor U22516 (N_22516,N_21301,N_21400);
nor U22517 (N_22517,N_20482,N_21213);
or U22518 (N_22518,N_20484,N_21300);
or U22519 (N_22519,N_21203,N_20869);
and U22520 (N_22520,N_21581,N_21334);
nor U22521 (N_22521,N_21320,N_20903);
nand U22522 (N_22522,N_21515,N_21388);
nand U22523 (N_22523,N_21214,N_21330);
and U22524 (N_22524,N_21226,N_21558);
nand U22525 (N_22525,N_20973,N_20431);
or U22526 (N_22526,N_20414,N_21152);
nand U22527 (N_22527,N_21116,N_21319);
nand U22528 (N_22528,N_21515,N_20825);
and U22529 (N_22529,N_20691,N_21432);
and U22530 (N_22530,N_20535,N_20865);
nor U22531 (N_22531,N_21488,N_20760);
nor U22532 (N_22532,N_21503,N_21194);
nor U22533 (N_22533,N_21567,N_21409);
and U22534 (N_22534,N_20637,N_20711);
or U22535 (N_22535,N_21321,N_20777);
xor U22536 (N_22536,N_21482,N_20702);
or U22537 (N_22537,N_20998,N_20795);
nor U22538 (N_22538,N_21126,N_20998);
and U22539 (N_22539,N_20989,N_20981);
or U22540 (N_22540,N_20812,N_20702);
nor U22541 (N_22541,N_21591,N_20685);
and U22542 (N_22542,N_20964,N_21251);
xor U22543 (N_22543,N_20683,N_20964);
nand U22544 (N_22544,N_20899,N_21573);
and U22545 (N_22545,N_21502,N_21543);
and U22546 (N_22546,N_20423,N_21543);
xor U22547 (N_22547,N_21091,N_20867);
and U22548 (N_22548,N_21488,N_20505);
nor U22549 (N_22549,N_21096,N_21219);
xnor U22550 (N_22550,N_21548,N_21569);
and U22551 (N_22551,N_21012,N_20476);
or U22552 (N_22552,N_20931,N_21206);
and U22553 (N_22553,N_21097,N_20519);
and U22554 (N_22554,N_21431,N_20546);
and U22555 (N_22555,N_20506,N_21529);
and U22556 (N_22556,N_20698,N_21118);
and U22557 (N_22557,N_20986,N_20647);
or U22558 (N_22558,N_21421,N_21086);
nor U22559 (N_22559,N_21267,N_20554);
and U22560 (N_22560,N_21044,N_20606);
xnor U22561 (N_22561,N_21261,N_20448);
xnor U22562 (N_22562,N_20491,N_21539);
nand U22563 (N_22563,N_20809,N_21075);
xor U22564 (N_22564,N_20420,N_21258);
xor U22565 (N_22565,N_20903,N_20423);
or U22566 (N_22566,N_20621,N_21307);
nor U22567 (N_22567,N_20575,N_20842);
or U22568 (N_22568,N_21367,N_20576);
and U22569 (N_22569,N_21203,N_20512);
and U22570 (N_22570,N_21228,N_21365);
nor U22571 (N_22571,N_21162,N_20889);
and U22572 (N_22572,N_21364,N_20438);
and U22573 (N_22573,N_20612,N_20721);
nor U22574 (N_22574,N_21351,N_20654);
nor U22575 (N_22575,N_20822,N_20638);
nand U22576 (N_22576,N_20493,N_21077);
and U22577 (N_22577,N_21414,N_21097);
or U22578 (N_22578,N_21599,N_20748);
nor U22579 (N_22579,N_20616,N_20944);
xor U22580 (N_22580,N_20840,N_20675);
and U22581 (N_22581,N_20512,N_21126);
xnor U22582 (N_22582,N_20835,N_20558);
nor U22583 (N_22583,N_21113,N_21584);
nand U22584 (N_22584,N_20699,N_20849);
nand U22585 (N_22585,N_21218,N_20875);
nand U22586 (N_22586,N_20400,N_20443);
and U22587 (N_22587,N_21443,N_21140);
and U22588 (N_22588,N_21205,N_20491);
nor U22589 (N_22589,N_20980,N_20427);
or U22590 (N_22590,N_20811,N_21146);
or U22591 (N_22591,N_20705,N_21027);
and U22592 (N_22592,N_21363,N_20423);
xor U22593 (N_22593,N_21111,N_20909);
and U22594 (N_22594,N_20697,N_20741);
xor U22595 (N_22595,N_21398,N_20573);
xor U22596 (N_22596,N_20467,N_21239);
xnor U22597 (N_22597,N_21465,N_21287);
or U22598 (N_22598,N_21082,N_21276);
xor U22599 (N_22599,N_20934,N_21003);
nand U22600 (N_22600,N_21250,N_21115);
xnor U22601 (N_22601,N_20948,N_21212);
or U22602 (N_22602,N_21417,N_20625);
xor U22603 (N_22603,N_21415,N_20792);
nor U22604 (N_22604,N_20684,N_21441);
and U22605 (N_22605,N_21460,N_21018);
nand U22606 (N_22606,N_20767,N_20481);
and U22607 (N_22607,N_21287,N_20610);
xor U22608 (N_22608,N_21424,N_21563);
nand U22609 (N_22609,N_20719,N_20673);
nand U22610 (N_22610,N_21146,N_20940);
xor U22611 (N_22611,N_21327,N_20712);
xor U22612 (N_22612,N_20420,N_21043);
and U22613 (N_22613,N_20827,N_21529);
nor U22614 (N_22614,N_20505,N_20760);
xnor U22615 (N_22615,N_21521,N_21309);
nor U22616 (N_22616,N_21446,N_20610);
nand U22617 (N_22617,N_20944,N_20960);
nand U22618 (N_22618,N_21209,N_21335);
or U22619 (N_22619,N_21114,N_20566);
and U22620 (N_22620,N_21527,N_21004);
nor U22621 (N_22621,N_20727,N_20851);
nand U22622 (N_22622,N_21039,N_21460);
nand U22623 (N_22623,N_21182,N_21134);
xor U22624 (N_22624,N_21046,N_20407);
or U22625 (N_22625,N_21579,N_21341);
and U22626 (N_22626,N_21369,N_21121);
xnor U22627 (N_22627,N_20640,N_21425);
or U22628 (N_22628,N_21113,N_20708);
nand U22629 (N_22629,N_21294,N_21088);
and U22630 (N_22630,N_21197,N_20572);
and U22631 (N_22631,N_20476,N_21184);
nand U22632 (N_22632,N_21493,N_21316);
xnor U22633 (N_22633,N_21272,N_20719);
nand U22634 (N_22634,N_21518,N_21399);
or U22635 (N_22635,N_21099,N_21466);
nand U22636 (N_22636,N_20666,N_21384);
xnor U22637 (N_22637,N_21197,N_21412);
nor U22638 (N_22638,N_20440,N_21412);
nand U22639 (N_22639,N_20504,N_21500);
or U22640 (N_22640,N_20642,N_21143);
nand U22641 (N_22641,N_20894,N_20502);
and U22642 (N_22642,N_21371,N_21399);
and U22643 (N_22643,N_21115,N_20667);
and U22644 (N_22644,N_21147,N_20495);
and U22645 (N_22645,N_21394,N_21320);
nor U22646 (N_22646,N_20425,N_20974);
xnor U22647 (N_22647,N_20630,N_20430);
or U22648 (N_22648,N_20888,N_21444);
xnor U22649 (N_22649,N_21451,N_20772);
nand U22650 (N_22650,N_20836,N_21385);
xnor U22651 (N_22651,N_20591,N_21572);
nand U22652 (N_22652,N_21470,N_20897);
xor U22653 (N_22653,N_20663,N_21215);
xnor U22654 (N_22654,N_20823,N_20807);
or U22655 (N_22655,N_20823,N_20792);
nor U22656 (N_22656,N_20784,N_21167);
nor U22657 (N_22657,N_21051,N_20998);
xor U22658 (N_22658,N_20486,N_21005);
xnor U22659 (N_22659,N_20686,N_20442);
nand U22660 (N_22660,N_21089,N_20607);
xor U22661 (N_22661,N_20831,N_21547);
and U22662 (N_22662,N_20879,N_21378);
xnor U22663 (N_22663,N_20838,N_21587);
xnor U22664 (N_22664,N_21306,N_20956);
xnor U22665 (N_22665,N_21477,N_20640);
and U22666 (N_22666,N_21003,N_21459);
xor U22667 (N_22667,N_21350,N_20943);
nand U22668 (N_22668,N_20809,N_21546);
and U22669 (N_22669,N_21405,N_20445);
nor U22670 (N_22670,N_21424,N_21001);
and U22671 (N_22671,N_20499,N_20503);
nand U22672 (N_22672,N_21476,N_20927);
xor U22673 (N_22673,N_21219,N_21483);
xnor U22674 (N_22674,N_21357,N_21358);
and U22675 (N_22675,N_21478,N_21143);
xnor U22676 (N_22676,N_21055,N_20798);
nor U22677 (N_22677,N_20587,N_21525);
or U22678 (N_22678,N_20966,N_20829);
or U22679 (N_22679,N_21572,N_20658);
or U22680 (N_22680,N_21572,N_21023);
nor U22681 (N_22681,N_21474,N_21281);
xnor U22682 (N_22682,N_20493,N_21277);
nor U22683 (N_22683,N_20773,N_21527);
and U22684 (N_22684,N_20803,N_20780);
nor U22685 (N_22685,N_21376,N_20416);
or U22686 (N_22686,N_21392,N_20921);
nor U22687 (N_22687,N_21562,N_21592);
nand U22688 (N_22688,N_21464,N_20898);
or U22689 (N_22689,N_20515,N_20482);
nor U22690 (N_22690,N_21030,N_21479);
and U22691 (N_22691,N_20933,N_20511);
and U22692 (N_22692,N_20767,N_20742);
nand U22693 (N_22693,N_20791,N_21499);
xnor U22694 (N_22694,N_20817,N_20788);
or U22695 (N_22695,N_20786,N_21278);
nand U22696 (N_22696,N_20610,N_20694);
nor U22697 (N_22697,N_21234,N_20609);
and U22698 (N_22698,N_20562,N_20679);
or U22699 (N_22699,N_20562,N_20400);
or U22700 (N_22700,N_20864,N_20765);
and U22701 (N_22701,N_20659,N_20511);
nand U22702 (N_22702,N_20654,N_21079);
and U22703 (N_22703,N_20983,N_21174);
and U22704 (N_22704,N_20829,N_20649);
and U22705 (N_22705,N_20989,N_20785);
nor U22706 (N_22706,N_20970,N_21474);
nand U22707 (N_22707,N_21521,N_21382);
nor U22708 (N_22708,N_21420,N_20496);
nand U22709 (N_22709,N_21303,N_21454);
and U22710 (N_22710,N_20985,N_20931);
or U22711 (N_22711,N_21593,N_20955);
nor U22712 (N_22712,N_21230,N_21395);
xor U22713 (N_22713,N_20599,N_20657);
and U22714 (N_22714,N_21262,N_21137);
or U22715 (N_22715,N_20678,N_21485);
nor U22716 (N_22716,N_20874,N_20470);
or U22717 (N_22717,N_20736,N_21061);
or U22718 (N_22718,N_20424,N_21566);
nor U22719 (N_22719,N_20425,N_21259);
xor U22720 (N_22720,N_20835,N_20404);
and U22721 (N_22721,N_20518,N_21280);
nor U22722 (N_22722,N_21571,N_21030);
nor U22723 (N_22723,N_21560,N_20493);
nor U22724 (N_22724,N_21027,N_20874);
or U22725 (N_22725,N_20981,N_20735);
and U22726 (N_22726,N_20424,N_21405);
or U22727 (N_22727,N_20539,N_21585);
and U22728 (N_22728,N_21011,N_21462);
nand U22729 (N_22729,N_21106,N_20445);
or U22730 (N_22730,N_20880,N_21168);
nor U22731 (N_22731,N_20642,N_21392);
and U22732 (N_22732,N_20439,N_20531);
nor U22733 (N_22733,N_21599,N_21520);
or U22734 (N_22734,N_20489,N_21051);
nand U22735 (N_22735,N_21427,N_20909);
nand U22736 (N_22736,N_20693,N_21287);
nand U22737 (N_22737,N_21049,N_20709);
or U22738 (N_22738,N_20993,N_20439);
or U22739 (N_22739,N_21010,N_20442);
nor U22740 (N_22740,N_21433,N_20629);
nor U22741 (N_22741,N_21333,N_20417);
and U22742 (N_22742,N_20615,N_20400);
nand U22743 (N_22743,N_20424,N_20768);
nand U22744 (N_22744,N_21229,N_21141);
or U22745 (N_22745,N_20513,N_21263);
xnor U22746 (N_22746,N_21147,N_20762);
and U22747 (N_22747,N_20864,N_20576);
nand U22748 (N_22748,N_21112,N_20796);
xnor U22749 (N_22749,N_21055,N_21053);
xnor U22750 (N_22750,N_21556,N_20810);
xnor U22751 (N_22751,N_20880,N_20606);
nand U22752 (N_22752,N_20926,N_20851);
xnor U22753 (N_22753,N_20656,N_21243);
or U22754 (N_22754,N_20512,N_20974);
nor U22755 (N_22755,N_21438,N_21073);
nor U22756 (N_22756,N_20479,N_21106);
xor U22757 (N_22757,N_21154,N_21012);
and U22758 (N_22758,N_21057,N_21247);
or U22759 (N_22759,N_20927,N_21150);
and U22760 (N_22760,N_21492,N_20643);
nor U22761 (N_22761,N_21457,N_20694);
nand U22762 (N_22762,N_20730,N_20554);
xor U22763 (N_22763,N_20963,N_20962);
and U22764 (N_22764,N_21391,N_21233);
or U22765 (N_22765,N_21521,N_21345);
xor U22766 (N_22766,N_20675,N_21237);
and U22767 (N_22767,N_21023,N_21016);
xor U22768 (N_22768,N_20764,N_21250);
xnor U22769 (N_22769,N_20510,N_21456);
or U22770 (N_22770,N_21447,N_21190);
or U22771 (N_22771,N_20449,N_20697);
xnor U22772 (N_22772,N_20829,N_21561);
xnor U22773 (N_22773,N_20457,N_20735);
or U22774 (N_22774,N_21450,N_20564);
nor U22775 (N_22775,N_21218,N_21433);
xnor U22776 (N_22776,N_21499,N_20497);
xor U22777 (N_22777,N_21148,N_20882);
nand U22778 (N_22778,N_21351,N_21551);
nand U22779 (N_22779,N_20589,N_21304);
and U22780 (N_22780,N_21430,N_21074);
or U22781 (N_22781,N_20547,N_20751);
xnor U22782 (N_22782,N_20424,N_20665);
nand U22783 (N_22783,N_20441,N_21422);
and U22784 (N_22784,N_20768,N_20986);
xor U22785 (N_22785,N_21379,N_20618);
nand U22786 (N_22786,N_21246,N_20790);
or U22787 (N_22787,N_21147,N_20942);
nand U22788 (N_22788,N_20935,N_21104);
nand U22789 (N_22789,N_21575,N_20752);
and U22790 (N_22790,N_20846,N_20758);
nand U22791 (N_22791,N_21182,N_21458);
nor U22792 (N_22792,N_20586,N_20679);
nor U22793 (N_22793,N_21301,N_20496);
nand U22794 (N_22794,N_20864,N_21577);
xnor U22795 (N_22795,N_20716,N_20436);
xnor U22796 (N_22796,N_20409,N_20895);
and U22797 (N_22797,N_20979,N_21555);
or U22798 (N_22798,N_21539,N_20853);
xor U22799 (N_22799,N_21444,N_21505);
or U22800 (N_22800,N_22039,N_21605);
or U22801 (N_22801,N_22663,N_21721);
xnor U22802 (N_22802,N_21852,N_22376);
or U22803 (N_22803,N_22422,N_22233);
and U22804 (N_22804,N_22453,N_22547);
nor U22805 (N_22805,N_22249,N_22562);
nor U22806 (N_22806,N_22150,N_22049);
or U22807 (N_22807,N_22478,N_22045);
or U22808 (N_22808,N_21664,N_22630);
and U22809 (N_22809,N_21991,N_22671);
nand U22810 (N_22810,N_22207,N_22391);
nor U22811 (N_22811,N_22351,N_22483);
or U22812 (N_22812,N_22796,N_21633);
or U22813 (N_22813,N_22604,N_21672);
and U22814 (N_22814,N_22290,N_22579);
or U22815 (N_22815,N_22193,N_21900);
nand U22816 (N_22816,N_22423,N_22229);
nor U22817 (N_22817,N_22472,N_21988);
nand U22818 (N_22818,N_22775,N_21893);
nand U22819 (N_22819,N_21689,N_22757);
nand U22820 (N_22820,N_21654,N_22690);
and U22821 (N_22821,N_22582,N_22467);
xnor U22822 (N_22822,N_22257,N_21801);
nor U22823 (N_22823,N_22743,N_21744);
nand U22824 (N_22824,N_22642,N_22074);
or U22825 (N_22825,N_21833,N_22718);
nand U22826 (N_22826,N_22486,N_22747);
or U22827 (N_22827,N_21766,N_22541);
nand U22828 (N_22828,N_21824,N_21691);
or U22829 (N_22829,N_22023,N_21614);
or U22830 (N_22830,N_22687,N_21874);
nor U22831 (N_22831,N_21939,N_22659);
or U22832 (N_22832,N_22410,N_22355);
nor U22833 (N_22833,N_22738,N_22224);
and U22834 (N_22834,N_22250,N_22130);
and U22835 (N_22835,N_21945,N_22773);
xor U22836 (N_22836,N_22463,N_22251);
nor U22837 (N_22837,N_22360,N_22585);
nor U22838 (N_22838,N_21968,N_22199);
nor U22839 (N_22839,N_21918,N_21829);
nor U22840 (N_22840,N_22765,N_22634);
nand U22841 (N_22841,N_22037,N_22436);
or U22842 (N_22842,N_22756,N_22416);
or U22843 (N_22843,N_21869,N_22244);
or U22844 (N_22844,N_21867,N_22700);
xnor U22845 (N_22845,N_22245,N_21719);
or U22846 (N_22846,N_22689,N_22699);
and U22847 (N_22847,N_22401,N_22145);
nand U22848 (N_22848,N_22632,N_21944);
nor U22849 (N_22849,N_22396,N_22750);
nand U22850 (N_22850,N_21873,N_22214);
and U22851 (N_22851,N_21959,N_22383);
nand U22852 (N_22852,N_22415,N_22664);
nor U22853 (N_22853,N_22669,N_22397);
and U22854 (N_22854,N_21625,N_21982);
nor U22855 (N_22855,N_22452,N_22685);
nand U22856 (N_22856,N_22073,N_22313);
xor U22857 (N_22857,N_22650,N_22782);
nand U22858 (N_22858,N_22460,N_22378);
nand U22859 (N_22859,N_22029,N_21643);
nand U22860 (N_22860,N_22232,N_21679);
nor U22861 (N_22861,N_21804,N_21876);
nor U22862 (N_22862,N_22160,N_21717);
nor U22863 (N_22863,N_22456,N_22442);
nand U22864 (N_22864,N_22319,N_22169);
nor U22865 (N_22865,N_21805,N_22728);
xnor U22866 (N_22866,N_21899,N_21765);
nand U22867 (N_22867,N_22785,N_22361);
xor U22868 (N_22868,N_22783,N_22609);
nand U22869 (N_22869,N_22267,N_22119);
nand U22870 (N_22870,N_22139,N_21704);
and U22871 (N_22871,N_21619,N_22296);
xor U22872 (N_22872,N_22680,N_22051);
xor U22873 (N_22873,N_22474,N_21865);
nand U22874 (N_22874,N_22204,N_22525);
and U22875 (N_22875,N_22243,N_21888);
and U22876 (N_22876,N_21911,N_22166);
xor U22877 (N_22877,N_21973,N_22724);
or U22878 (N_22878,N_22753,N_21700);
nor U22879 (N_22879,N_22109,N_22485);
nand U22880 (N_22880,N_21610,N_22067);
nor U22881 (N_22881,N_21743,N_22034);
nor U22882 (N_22882,N_22187,N_22600);
nand U22883 (N_22883,N_22066,N_21661);
or U22884 (N_22884,N_22320,N_21795);
nor U22885 (N_22885,N_21769,N_22786);
nor U22886 (N_22886,N_21797,N_22056);
xnor U22887 (N_22887,N_22778,N_22352);
or U22888 (N_22888,N_22566,N_22613);
and U22889 (N_22889,N_21894,N_22789);
nor U22890 (N_22890,N_22674,N_22009);
nand U22891 (N_22891,N_21884,N_22437);
nand U22892 (N_22892,N_21861,N_22519);
and U22893 (N_22893,N_22333,N_22622);
and U22894 (N_22894,N_22236,N_22777);
xor U22895 (N_22895,N_22060,N_22105);
nor U22896 (N_22896,N_22758,N_22127);
nand U22897 (N_22897,N_22618,N_22683);
or U22898 (N_22898,N_21663,N_22400);
and U22899 (N_22899,N_22516,N_21849);
or U22900 (N_22900,N_22022,N_22253);
nand U22901 (N_22901,N_22714,N_21621);
or U22902 (N_22902,N_22768,N_22165);
nor U22903 (N_22903,N_21648,N_21832);
or U22904 (N_22904,N_22246,N_22476);
nand U22905 (N_22905,N_22480,N_21677);
or U22906 (N_22906,N_22503,N_22226);
or U22907 (N_22907,N_22210,N_22629);
and U22908 (N_22908,N_22247,N_22314);
or U22909 (N_22909,N_22504,N_21995);
nand U22910 (N_22910,N_22665,N_22784);
xnor U22911 (N_22911,N_21668,N_21822);
nand U22912 (N_22912,N_21601,N_21686);
or U22913 (N_22913,N_21741,N_22272);
or U22914 (N_22914,N_21620,N_22184);
nor U22915 (N_22915,N_21715,N_22543);
nand U22916 (N_22916,N_22538,N_22217);
and U22917 (N_22917,N_21688,N_22398);
xnor U22918 (N_22918,N_22046,N_21803);
or U22919 (N_22919,N_22451,N_22592);
and U22920 (N_22920,N_21738,N_21669);
nor U22921 (N_22921,N_22740,N_22495);
nor U22922 (N_22922,N_22473,N_21613);
nand U22923 (N_22923,N_22596,N_22106);
nand U22924 (N_22924,N_22752,N_22248);
and U22925 (N_22925,N_22524,N_21961);
nand U22926 (N_22926,N_21792,N_22156);
nand U22927 (N_22927,N_22438,N_21993);
nand U22928 (N_22928,N_21622,N_22318);
and U22929 (N_22929,N_21750,N_22481);
nand U22930 (N_22930,N_21752,N_21800);
or U22931 (N_22931,N_22194,N_22429);
or U22932 (N_22932,N_22667,N_21904);
and U22933 (N_22933,N_21952,N_22607);
nor U22934 (N_22934,N_22539,N_21720);
nor U22935 (N_22935,N_22470,N_21705);
or U22936 (N_22936,N_22697,N_22694);
or U22937 (N_22937,N_22307,N_22061);
nand U22938 (N_22938,N_22734,N_22557);
nor U22939 (N_22939,N_22168,N_22614);
or U22940 (N_22940,N_21971,N_21877);
and U22941 (N_22941,N_22354,N_22167);
xnor U22942 (N_22942,N_22334,N_22108);
xor U22943 (N_22943,N_22723,N_22731);
nand U22944 (N_22944,N_22588,N_22071);
and U22945 (N_22945,N_21838,N_22120);
or U22946 (N_22946,N_22366,N_22759);
and U22947 (N_22947,N_21799,N_22475);
or U22948 (N_22948,N_22534,N_22326);
nor U22949 (N_22949,N_22370,N_22129);
and U22950 (N_22950,N_22513,N_22624);
or U22951 (N_22951,N_22348,N_21645);
and U22952 (N_22952,N_22338,N_22392);
nand U22953 (N_22953,N_22294,N_22241);
nand U22954 (N_22954,N_21934,N_22793);
nand U22955 (N_22955,N_22344,N_22365);
xnor U22956 (N_22956,N_22692,N_21623);
nand U22957 (N_22957,N_22490,N_21889);
nand U22958 (N_22958,N_21665,N_21928);
and U22959 (N_22959,N_21810,N_22528);
nor U22960 (N_22960,N_22617,N_22568);
xnor U22961 (N_22961,N_21956,N_22556);
or U22962 (N_22962,N_21908,N_21975);
nand U22963 (N_22963,N_21747,N_22535);
and U22964 (N_22964,N_22761,N_22603);
xnor U22965 (N_22965,N_21785,N_21639);
and U22966 (N_22966,N_22181,N_21949);
nand U22967 (N_22967,N_21967,N_22576);
nor U22968 (N_22968,N_22271,N_21714);
or U22969 (N_22969,N_21909,N_22363);
nand U22970 (N_22970,N_21757,N_22620);
and U22971 (N_22971,N_22005,N_22339);
nand U22972 (N_22972,N_22626,N_22015);
nand U22973 (N_22973,N_22494,N_22517);
xor U22974 (N_22974,N_22335,N_22721);
or U22975 (N_22975,N_22175,N_22058);
xnor U22976 (N_22976,N_22610,N_22762);
nand U22977 (N_22977,N_22096,N_21969);
and U22978 (N_22978,N_22379,N_21722);
xor U22979 (N_22979,N_22703,N_22545);
or U22980 (N_22980,N_22084,N_22371);
xor U22981 (N_22981,N_22121,N_22792);
and U22982 (N_22982,N_22043,N_22040);
xnor U22983 (N_22983,N_22085,N_22446);
nand U22984 (N_22984,N_22716,N_22114);
xnor U22985 (N_22985,N_22563,N_22087);
and U22986 (N_22986,N_22135,N_22321);
xnor U22987 (N_22987,N_21895,N_22310);
nand U22988 (N_22988,N_21710,N_22183);
nand U22989 (N_22989,N_21606,N_21624);
or U22990 (N_22990,N_21989,N_22123);
or U22991 (N_22991,N_22107,N_22011);
nand U22992 (N_22992,N_22180,N_21657);
and U22993 (N_22993,N_22542,N_22044);
xor U22994 (N_22994,N_21842,N_22605);
or U22995 (N_22995,N_22502,N_21687);
and U22996 (N_22996,N_22515,N_22657);
or U22997 (N_22997,N_22308,N_22522);
nand U22998 (N_22998,N_21635,N_22197);
nor U22999 (N_22999,N_22035,N_22449);
and U23000 (N_23000,N_21641,N_21859);
nor U23001 (N_23001,N_21812,N_21948);
or U23002 (N_23002,N_21727,N_22748);
xor U23003 (N_23003,N_21807,N_22551);
nor U23004 (N_23004,N_22010,N_21607);
and U23005 (N_23005,N_22678,N_21731);
or U23006 (N_23006,N_22098,N_22076);
xnor U23007 (N_23007,N_21789,N_22091);
nand U23008 (N_23008,N_21777,N_21706);
or U23009 (N_23009,N_21760,N_22162);
xor U23010 (N_23010,N_22727,N_22549);
or U23011 (N_23011,N_21951,N_22275);
nor U23012 (N_23012,N_22128,N_21782);
nand U23013 (N_23013,N_22277,N_22345);
nor U23014 (N_23014,N_22564,N_22599);
and U23015 (N_23015,N_21942,N_22681);
nand U23016 (N_23016,N_21612,N_22403);
nor U23017 (N_23017,N_22203,N_22636);
nand U23018 (N_23018,N_21881,N_21604);
nand U23019 (N_23019,N_22050,N_22769);
xnor U23020 (N_23020,N_22269,N_21667);
or U23021 (N_23021,N_22325,N_21977);
xor U23022 (N_23022,N_22394,N_22698);
nor U23023 (N_23023,N_21675,N_22368);
or U23024 (N_23024,N_21848,N_22342);
xnor U23025 (N_23025,N_22033,N_21809);
and U23026 (N_23026,N_21902,N_21755);
or U23027 (N_23027,N_21966,N_21781);
nor U23028 (N_23028,N_22788,N_21768);
nand U23029 (N_23029,N_22302,N_22695);
and U23030 (N_23030,N_21846,N_21814);
and U23031 (N_23031,N_22118,N_21646);
or U23032 (N_23032,N_22216,N_22508);
nand U23033 (N_23033,N_22266,N_21980);
xor U23034 (N_23034,N_22791,N_21671);
xor U23035 (N_23035,N_21882,N_22159);
nor U23036 (N_23036,N_21767,N_22565);
or U23037 (N_23037,N_22670,N_22461);
and U23038 (N_23038,N_21746,N_22493);
nand U23039 (N_23039,N_21910,N_22751);
and U23040 (N_23040,N_22151,N_21868);
and U23041 (N_23041,N_22003,N_21616);
nor U23042 (N_23042,N_21924,N_22025);
or U23043 (N_23043,N_22016,N_21730);
and U23044 (N_23044,N_22041,N_22268);
nand U23045 (N_23045,N_22763,N_22309);
nand U23046 (N_23046,N_22717,N_22691);
nor U23047 (N_23047,N_21745,N_21608);
xor U23048 (N_23048,N_21630,N_22036);
xnor U23049 (N_23049,N_21703,N_22640);
nand U23050 (N_23050,N_22125,N_22627);
nor U23051 (N_23051,N_21775,N_21855);
or U23052 (N_23052,N_22772,N_21783);
nor U23053 (N_23053,N_22395,N_22255);
nand U23054 (N_23054,N_21923,N_22350);
and U23055 (N_23055,N_22643,N_21990);
nand U23056 (N_23056,N_21913,N_22090);
xnor U23057 (N_23057,N_22787,N_22346);
nand U23058 (N_23058,N_22002,N_22509);
or U23059 (N_23059,N_22725,N_22293);
or U23060 (N_23060,N_21798,N_22137);
or U23061 (N_23061,N_22340,N_22225);
nand U23062 (N_23062,N_21866,N_22089);
xnor U23063 (N_23063,N_22052,N_21695);
nand U23064 (N_23064,N_22559,N_22735);
and U23065 (N_23065,N_22567,N_22021);
nor U23066 (N_23066,N_21762,N_22206);
nor U23067 (N_23067,N_22676,N_22651);
xor U23068 (N_23068,N_22209,N_22615);
xor U23069 (N_23069,N_22235,N_21753);
and U23070 (N_23070,N_21826,N_22256);
nand U23071 (N_23071,N_21841,N_22072);
and U23072 (N_23072,N_22679,N_22649);
and U23073 (N_23073,N_21958,N_22575);
and U23074 (N_23074,N_21656,N_22274);
and U23075 (N_23075,N_22215,N_22497);
xor U23076 (N_23076,N_21659,N_22202);
or U23077 (N_23077,N_21938,N_21627);
nand U23078 (N_23078,N_21883,N_22311);
or U23079 (N_23079,N_22148,N_21864);
nand U23080 (N_23080,N_21886,N_22544);
nor U23081 (N_23081,N_22668,N_21817);
xnor U23082 (N_23082,N_22656,N_22420);
nor U23083 (N_23083,N_22279,N_22693);
and U23084 (N_23084,N_21907,N_21839);
or U23085 (N_23085,N_22413,N_21778);
nand U23086 (N_23086,N_22100,N_22583);
or U23087 (N_23087,N_21850,N_22315);
xnor U23088 (N_23088,N_22264,N_21712);
and U23089 (N_23089,N_22144,N_21749);
nor U23090 (N_23090,N_22064,N_22295);
or U23091 (N_23091,N_22459,N_21739);
and U23092 (N_23092,N_22684,N_22434);
nor U23093 (N_23093,N_22349,N_22462);
nand U23094 (N_23094,N_22358,N_22428);
and U23095 (N_23095,N_22492,N_22702);
xnor U23096 (N_23096,N_22377,N_21825);
and U23097 (N_23097,N_22570,N_22292);
or U23098 (N_23098,N_22682,N_22688);
and U23099 (N_23099,N_22387,N_22755);
nand U23100 (N_23100,N_22482,N_22327);
nor U23101 (N_23101,N_22399,N_22157);
nand U23102 (N_23102,N_21770,N_22238);
nor U23103 (N_23103,N_22218,N_21920);
nand U23104 (N_23104,N_22794,N_21964);
nor U23105 (N_23105,N_22031,N_22468);
or U23106 (N_23106,N_22448,N_22343);
xor U23107 (N_23107,N_22324,N_22514);
and U23108 (N_23108,N_22303,N_21733);
or U23109 (N_23109,N_21985,N_22178);
xnor U23110 (N_23110,N_21835,N_22195);
or U23111 (N_23111,N_22196,N_21957);
xor U23112 (N_23112,N_21912,N_21981);
nand U23113 (N_23113,N_22301,N_22337);
and U23114 (N_23114,N_22057,N_22484);
and U23115 (N_23115,N_22405,N_22116);
and U23116 (N_23116,N_21734,N_21729);
nor U23117 (N_23117,N_22357,N_22297);
nor U23118 (N_23118,N_22540,N_22404);
nor U23119 (N_23119,N_22347,N_22637);
nand U23120 (N_23120,N_21611,N_22639);
xor U23121 (N_23121,N_22533,N_22465);
nor U23122 (N_23122,N_22097,N_22790);
xnor U23123 (N_23123,N_22553,N_22648);
xor U23124 (N_23124,N_22173,N_22631);
and U23125 (N_23125,N_21987,N_21644);
or U23126 (N_23126,N_22536,N_22720);
xor U23127 (N_23127,N_22131,N_21954);
xor U23128 (N_23128,N_22198,N_22781);
and U23129 (N_23129,N_21806,N_21692);
nand U23130 (N_23130,N_22208,N_21940);
and U23131 (N_23131,N_21662,N_22708);
and U23132 (N_23132,N_21640,N_22587);
xnor U23133 (N_23133,N_22414,N_22185);
or U23134 (N_23134,N_22580,N_22088);
and U23135 (N_23135,N_21955,N_21693);
xnor U23136 (N_23136,N_22287,N_22007);
nor U23137 (N_23137,N_22407,N_22126);
xor U23138 (N_23138,N_22571,N_22261);
nand U23139 (N_23139,N_22730,N_21784);
and U23140 (N_23140,N_22767,N_22799);
xor U23141 (N_23141,N_22000,N_22093);
and U23142 (N_23142,N_22645,N_22715);
xor U23143 (N_23143,N_22662,N_22602);
nor U23144 (N_23144,N_22555,N_22589);
and U23145 (N_23145,N_22739,N_21701);
nor U23146 (N_23146,N_21709,N_22273);
xor U23147 (N_23147,N_22498,N_22099);
xnor U23148 (N_23148,N_22189,N_21631);
and U23149 (N_23149,N_22179,N_22026);
and U23150 (N_23150,N_22006,N_21921);
xor U23151 (N_23151,N_22477,N_21647);
or U23152 (N_23152,N_21694,N_22286);
nand U23153 (N_23153,N_22223,N_22328);
nor U23154 (N_23154,N_22265,N_22155);
nor U23155 (N_23155,N_22496,N_22149);
nand U23156 (N_23156,N_21754,N_21698);
xnor U23157 (N_23157,N_22635,N_22445);
xnor U23158 (N_23158,N_21723,N_22393);
and U23159 (N_23159,N_22323,N_22263);
nor U23160 (N_23160,N_22406,N_22242);
xor U23161 (N_23161,N_22611,N_22234);
nand U23162 (N_23162,N_22625,N_22369);
or U23163 (N_23163,N_21690,N_21699);
and U23164 (N_23164,N_22075,N_21793);
and U23165 (N_23165,N_21779,N_21780);
xnor U23166 (N_23166,N_22054,N_22638);
or U23167 (N_23167,N_22278,N_22227);
xnor U23168 (N_23168,N_21890,N_22707);
or U23169 (N_23169,N_22499,N_22312);
or U23170 (N_23170,N_22221,N_22288);
and U23171 (N_23171,N_22136,N_21843);
nand U23172 (N_23172,N_22222,N_22464);
or U23173 (N_23173,N_21929,N_22647);
nor U23174 (N_23174,N_21636,N_22101);
nand U23175 (N_23175,N_22726,N_21925);
nand U23176 (N_23176,N_21953,N_22212);
nor U23177 (N_23177,N_21684,N_22048);
nor U23178 (N_23178,N_21965,N_21653);
nor U23179 (N_23179,N_22586,N_22431);
xor U23180 (N_23180,N_22706,N_22741);
or U23181 (N_23181,N_22518,N_21628);
xor U23182 (N_23182,N_21634,N_22488);
xnor U23183 (N_23183,N_21974,N_22133);
and U23184 (N_23184,N_22746,N_22736);
nand U23185 (N_23185,N_22594,N_22163);
nand U23186 (N_23186,N_22381,N_22412);
nand U23187 (N_23187,N_21936,N_22779);
or U23188 (N_23188,N_22471,N_22170);
nand U23189 (N_23189,N_22001,N_21816);
nand U23190 (N_23190,N_21742,N_21851);
or U23191 (N_23191,N_22623,N_22030);
xor U23192 (N_23192,N_21823,N_22749);
nor U23193 (N_23193,N_22455,N_22182);
nor U23194 (N_23194,N_22068,N_21708);
xor U23195 (N_23195,N_21702,N_21676);
nor U23196 (N_23196,N_22220,N_22063);
and U23197 (N_23197,N_22329,N_22548);
and U23198 (N_23198,N_21711,N_21748);
xor U23199 (N_23199,N_22158,N_21856);
nand U23200 (N_23200,N_22004,N_21994);
nor U23201 (N_23201,N_22171,N_22299);
xor U23202 (N_23202,N_22284,N_21932);
nor U23203 (N_23203,N_22032,N_21901);
or U23204 (N_23204,N_22188,N_22439);
nand U23205 (N_23205,N_22373,N_21802);
nor U23206 (N_23206,N_22316,N_22134);
and U23207 (N_23207,N_21916,N_22262);
nand U23208 (N_23208,N_22776,N_22505);
or U23209 (N_23209,N_22584,N_22027);
nor U23210 (N_23210,N_21682,N_22597);
and U23211 (N_23211,N_22142,N_22069);
xor U23212 (N_23212,N_22491,N_22201);
nor U23213 (N_23213,N_22177,N_21600);
nand U23214 (N_23214,N_22704,N_22095);
xnor U23215 (N_23215,N_22024,N_22132);
or U23216 (N_23216,N_22709,N_22191);
nor U23217 (N_23217,N_22621,N_22729);
or U23218 (N_23218,N_22102,N_21853);
nor U23219 (N_23219,N_22259,N_21903);
nor U23220 (N_23220,N_21724,N_21976);
and U23221 (N_23221,N_22280,N_22424);
xor U23222 (N_23222,N_22047,N_22577);
nand U23223 (N_23223,N_22590,N_22013);
and U23224 (N_23224,N_22795,N_22192);
and U23225 (N_23225,N_22552,N_21808);
or U23226 (N_23226,N_22432,N_21602);
nand U23227 (N_23227,N_21773,N_21642);
xor U23228 (N_23228,N_22719,N_22537);
nand U23229 (N_23229,N_22331,N_21854);
and U23230 (N_23230,N_22053,N_22304);
nand U23231 (N_23231,N_22532,N_22506);
xor U23232 (N_23232,N_22332,N_21898);
nor U23233 (N_23233,N_22745,N_21840);
or U23234 (N_23234,N_21674,N_22382);
nand U23235 (N_23235,N_21919,N_22660);
nand U23236 (N_23236,N_22384,N_21764);
xnor U23237 (N_23237,N_22487,N_21986);
xor U23238 (N_23238,N_22140,N_22283);
nor U23239 (N_23239,N_21906,N_22143);
and U23240 (N_23240,N_22601,N_22305);
nand U23241 (N_23241,N_21872,N_22526);
and U23242 (N_23242,N_21790,N_22231);
nor U23243 (N_23243,N_22572,N_22141);
and U23244 (N_23244,N_22385,N_21998);
nand U23245 (N_23245,N_22153,N_22115);
nand U23246 (N_23246,N_22426,N_21943);
xor U23247 (N_23247,N_21941,N_22042);
nor U23248 (N_23248,N_21651,N_22529);
nor U23249 (N_23249,N_22070,N_21962);
or U23250 (N_23250,N_22531,N_21649);
nor U23251 (N_23251,N_22458,N_22443);
xnor U23252 (N_23252,N_21847,N_22644);
nand U23253 (N_23253,N_22078,N_22213);
or U23254 (N_23254,N_21796,N_21891);
and U23255 (N_23255,N_22172,N_22174);
and U23256 (N_23256,N_21845,N_22317);
nor U23257 (N_23257,N_22560,N_22595);
and U23258 (N_23258,N_22417,N_22230);
nor U23259 (N_23259,N_22079,N_21758);
xnor U23260 (N_23260,N_22359,N_22673);
or U23261 (N_23261,N_22388,N_21858);
xnor U23262 (N_23262,N_22489,N_21819);
xor U23263 (N_23263,N_22512,N_21972);
or U23264 (N_23264,N_21946,N_22390);
or U23265 (N_23265,N_22457,N_22122);
xnor U23266 (N_23266,N_21950,N_22356);
nor U23267 (N_23267,N_22421,N_22270);
nand U23268 (N_23268,N_21897,N_22652);
xor U23269 (N_23269,N_21834,N_21818);
nand U23270 (N_23270,N_22375,N_22374);
nand U23271 (N_23271,N_22675,N_22111);
xnor U23272 (N_23272,N_22510,N_21629);
and U23273 (N_23273,N_21857,N_22012);
nand U23274 (N_23274,N_22710,N_22732);
nor U23275 (N_23275,N_21992,N_22770);
nand U23276 (N_23276,N_21771,N_22190);
or U23277 (N_23277,N_22402,N_21736);
nand U23278 (N_23278,N_22367,N_22501);
nand U23279 (N_23279,N_22646,N_22658);
and U23280 (N_23280,N_22086,N_22554);
nor U23281 (N_23281,N_21759,N_21860);
nor U23282 (N_23282,N_22330,N_22441);
and U23283 (N_23283,N_22094,N_22124);
xnor U23284 (N_23284,N_22633,N_22578);
xnor U23285 (N_23285,N_22154,N_21947);
nor U23286 (N_23286,N_22591,N_22276);
xnor U23287 (N_23287,N_22558,N_21707);
or U23288 (N_23288,N_21680,N_22017);
or U23289 (N_23289,N_22523,N_22696);
nand U23290 (N_23290,N_21732,N_22569);
xor U23291 (N_23291,N_22038,N_21905);
nor U23292 (N_23292,N_21666,N_21815);
nand U23293 (N_23293,N_21681,N_21878);
nor U23294 (N_23294,N_22705,N_22380);
nor U23295 (N_23295,N_22500,N_21879);
or U23296 (N_23296,N_22147,N_22764);
or U23297 (N_23297,N_22479,N_22530);
or U23298 (N_23298,N_22447,N_21880);
and U23299 (N_23299,N_22593,N_22336);
or U23300 (N_23300,N_22306,N_22418);
nor U23301 (N_23301,N_21791,N_22733);
xor U23302 (N_23302,N_21885,N_22573);
xnor U23303 (N_23303,N_21978,N_21931);
nor U23304 (N_23304,N_22774,N_22103);
nor U23305 (N_23305,N_21756,N_21776);
xnor U23306 (N_23306,N_21617,N_21660);
nor U23307 (N_23307,N_22092,N_21786);
nand U23308 (N_23308,N_22186,N_21696);
nor U23309 (N_23309,N_21763,N_22055);
or U23310 (N_23310,N_22527,N_22444);
nand U23311 (N_23311,N_22430,N_22771);
nand U23312 (N_23312,N_21632,N_21737);
nor U23313 (N_23313,N_22200,N_21821);
nand U23314 (N_23314,N_21937,N_22561);
and U23315 (N_23315,N_22065,N_22353);
and U23316 (N_23316,N_21718,N_21837);
xor U23317 (N_23317,N_22110,N_21922);
or U23318 (N_23318,N_21896,N_21740);
xnor U23319 (N_23319,N_21788,N_21915);
or U23320 (N_23320,N_22372,N_21761);
and U23321 (N_23321,N_22511,N_22300);
nor U23322 (N_23322,N_21935,N_22239);
nand U23323 (N_23323,N_22152,N_22433);
nor U23324 (N_23324,N_22059,N_21863);
xnor U23325 (N_23325,N_22606,N_22258);
nor U23326 (N_23326,N_21887,N_21831);
xor U23327 (N_23327,N_22322,N_22711);
nand U23328 (N_23328,N_21970,N_22228);
xor U23329 (N_23329,N_22364,N_21960);
and U23330 (N_23330,N_22581,N_21830);
or U23331 (N_23331,N_22281,N_22598);
or U23332 (N_23332,N_22008,N_22219);
nor U23333 (N_23333,N_22211,N_22616);
or U23334 (N_23334,N_21927,N_22386);
xor U23335 (N_23335,N_21983,N_21827);
xor U23336 (N_23336,N_21638,N_21926);
and U23337 (N_23337,N_22419,N_22737);
nor U23338 (N_23338,N_21726,N_21683);
or U23339 (N_23339,N_21655,N_21996);
nand U23340 (N_23340,N_21862,N_22655);
nor U23341 (N_23341,N_21728,N_22291);
nor U23342 (N_23342,N_21813,N_22408);
or U23343 (N_23343,N_21871,N_21892);
nand U23344 (N_23344,N_22411,N_22254);
nor U23345 (N_23345,N_21697,N_22520);
nor U23346 (N_23346,N_22754,N_21626);
xnor U23347 (N_23347,N_22521,N_22440);
and U23348 (N_23348,N_22798,N_22435);
nor U23349 (N_23349,N_22298,N_21930);
nand U23350 (N_23350,N_22450,N_22797);
nand U23351 (N_23351,N_21650,N_22341);
and U23352 (N_23352,N_21673,N_22409);
and U23353 (N_23353,N_21979,N_21997);
xnor U23354 (N_23354,N_21685,N_22020);
nor U23355 (N_23355,N_22082,N_21652);
nor U23356 (N_23356,N_22653,N_21603);
nand U23357 (N_23357,N_21751,N_22176);
and U23358 (N_23358,N_22612,N_22237);
xnor U23359 (N_23359,N_22641,N_22742);
or U23360 (N_23360,N_22014,N_21658);
or U23361 (N_23361,N_22661,N_21772);
nor U23362 (N_23362,N_22081,N_21725);
and U23363 (N_23363,N_22713,N_22164);
nand U23364 (N_23364,N_22138,N_21670);
or U23365 (N_23365,N_22083,N_22686);
nor U23366 (N_23366,N_21618,N_22028);
or U23367 (N_23367,N_22469,N_21716);
or U23368 (N_23368,N_22608,N_22260);
nor U23369 (N_23369,N_21820,N_22712);
nand U23370 (N_23370,N_22146,N_21615);
and U23371 (N_23371,N_22628,N_21609);
nor U23372 (N_23372,N_22654,N_22018);
nor U23373 (N_23373,N_22744,N_21713);
nor U23374 (N_23374,N_21999,N_22550);
nor U23375 (N_23375,N_22104,N_22362);
or U23376 (N_23376,N_22701,N_22289);
nand U23377 (N_23377,N_22666,N_21774);
nor U23378 (N_23378,N_22466,N_22507);
and U23379 (N_23379,N_22722,N_22117);
and U23380 (N_23380,N_21917,N_21735);
and U23381 (N_23381,N_22619,N_22780);
nor U23382 (N_23382,N_22546,N_22240);
nand U23383 (N_23383,N_22112,N_21984);
xnor U23384 (N_23384,N_22062,N_21828);
xnor U23385 (N_23385,N_22574,N_22161);
and U23386 (N_23386,N_22252,N_21844);
nand U23387 (N_23387,N_22285,N_22672);
nor U23388 (N_23388,N_22077,N_22766);
and U23389 (N_23389,N_21794,N_22205);
nor U23390 (N_23390,N_21811,N_21637);
nand U23391 (N_23391,N_21787,N_22454);
nand U23392 (N_23392,N_22677,N_21963);
or U23393 (N_23393,N_21870,N_21933);
xnor U23394 (N_23394,N_22113,N_22389);
nor U23395 (N_23395,N_22019,N_22427);
xnor U23396 (N_23396,N_21836,N_22282);
xnor U23397 (N_23397,N_21914,N_21678);
or U23398 (N_23398,N_22760,N_22425);
nor U23399 (N_23399,N_22080,N_21875);
nand U23400 (N_23400,N_22583,N_21845);
nor U23401 (N_23401,N_21644,N_22652);
xor U23402 (N_23402,N_22441,N_21851);
and U23403 (N_23403,N_22554,N_22387);
nand U23404 (N_23404,N_22455,N_22612);
nand U23405 (N_23405,N_22757,N_21633);
nand U23406 (N_23406,N_22097,N_22247);
or U23407 (N_23407,N_21732,N_22280);
or U23408 (N_23408,N_22027,N_22236);
or U23409 (N_23409,N_22390,N_22047);
nand U23410 (N_23410,N_21967,N_22603);
and U23411 (N_23411,N_21693,N_22178);
nand U23412 (N_23412,N_21627,N_21879);
and U23413 (N_23413,N_22195,N_22374);
xnor U23414 (N_23414,N_22648,N_21827);
or U23415 (N_23415,N_22796,N_21978);
and U23416 (N_23416,N_22179,N_22091);
and U23417 (N_23417,N_22294,N_21778);
and U23418 (N_23418,N_22488,N_21717);
nor U23419 (N_23419,N_21895,N_21660);
nand U23420 (N_23420,N_22312,N_22286);
xor U23421 (N_23421,N_22369,N_22173);
and U23422 (N_23422,N_22282,N_21831);
and U23423 (N_23423,N_22309,N_22259);
nor U23424 (N_23424,N_21806,N_22516);
and U23425 (N_23425,N_22732,N_22316);
nor U23426 (N_23426,N_21855,N_22104);
and U23427 (N_23427,N_21900,N_22354);
xnor U23428 (N_23428,N_22632,N_22535);
nand U23429 (N_23429,N_22253,N_22351);
nand U23430 (N_23430,N_22265,N_22126);
and U23431 (N_23431,N_21789,N_22518);
xor U23432 (N_23432,N_22216,N_21937);
and U23433 (N_23433,N_21738,N_22528);
xnor U23434 (N_23434,N_22466,N_22234);
and U23435 (N_23435,N_22238,N_22193);
nor U23436 (N_23436,N_21796,N_21931);
and U23437 (N_23437,N_21954,N_21792);
and U23438 (N_23438,N_22539,N_22767);
nand U23439 (N_23439,N_22398,N_21615);
and U23440 (N_23440,N_22753,N_21891);
nor U23441 (N_23441,N_22583,N_21998);
or U23442 (N_23442,N_21631,N_21806);
and U23443 (N_23443,N_22495,N_22531);
or U23444 (N_23444,N_22502,N_22620);
nand U23445 (N_23445,N_21999,N_22383);
nor U23446 (N_23446,N_22205,N_22704);
xor U23447 (N_23447,N_21888,N_21944);
nand U23448 (N_23448,N_22583,N_22215);
nor U23449 (N_23449,N_22237,N_22731);
nor U23450 (N_23450,N_22155,N_22383);
or U23451 (N_23451,N_22150,N_22015);
nor U23452 (N_23452,N_21995,N_21639);
and U23453 (N_23453,N_21914,N_21853);
or U23454 (N_23454,N_22018,N_21959);
xnor U23455 (N_23455,N_22306,N_21732);
nor U23456 (N_23456,N_22052,N_21697);
and U23457 (N_23457,N_22048,N_21705);
or U23458 (N_23458,N_22496,N_22375);
and U23459 (N_23459,N_22242,N_22374);
xnor U23460 (N_23460,N_21985,N_22207);
and U23461 (N_23461,N_21915,N_21625);
nand U23462 (N_23462,N_22148,N_21964);
or U23463 (N_23463,N_22748,N_22252);
and U23464 (N_23464,N_22722,N_21773);
and U23465 (N_23465,N_21928,N_21676);
nor U23466 (N_23466,N_21776,N_22718);
or U23467 (N_23467,N_22174,N_22642);
xnor U23468 (N_23468,N_22416,N_21992);
nor U23469 (N_23469,N_21670,N_22669);
nor U23470 (N_23470,N_21821,N_22475);
and U23471 (N_23471,N_22614,N_22524);
xnor U23472 (N_23472,N_22034,N_22632);
or U23473 (N_23473,N_21712,N_21625);
nor U23474 (N_23474,N_21908,N_22313);
and U23475 (N_23475,N_21865,N_22230);
nand U23476 (N_23476,N_22059,N_22123);
and U23477 (N_23477,N_22411,N_22550);
or U23478 (N_23478,N_22510,N_22101);
xor U23479 (N_23479,N_22280,N_21972);
nand U23480 (N_23480,N_21779,N_22431);
nor U23481 (N_23481,N_22299,N_21968);
nor U23482 (N_23482,N_22490,N_22414);
xnor U23483 (N_23483,N_21773,N_21742);
or U23484 (N_23484,N_22414,N_21880);
nand U23485 (N_23485,N_22024,N_22793);
nor U23486 (N_23486,N_22328,N_22568);
nor U23487 (N_23487,N_22017,N_22743);
or U23488 (N_23488,N_22012,N_22671);
xor U23489 (N_23489,N_22321,N_21637);
nor U23490 (N_23490,N_22032,N_22708);
nand U23491 (N_23491,N_21631,N_22343);
xnor U23492 (N_23492,N_22100,N_22243);
or U23493 (N_23493,N_22441,N_21629);
or U23494 (N_23494,N_22036,N_22201);
nand U23495 (N_23495,N_22388,N_22658);
xnor U23496 (N_23496,N_21887,N_22783);
xor U23497 (N_23497,N_22062,N_22176);
and U23498 (N_23498,N_21817,N_22559);
and U23499 (N_23499,N_22466,N_22530);
nand U23500 (N_23500,N_22065,N_22467);
or U23501 (N_23501,N_22724,N_21921);
nor U23502 (N_23502,N_22782,N_21793);
and U23503 (N_23503,N_22103,N_22390);
and U23504 (N_23504,N_22744,N_22796);
nand U23505 (N_23505,N_22431,N_21850);
and U23506 (N_23506,N_22748,N_21815);
xnor U23507 (N_23507,N_21693,N_22741);
xor U23508 (N_23508,N_22235,N_22533);
nor U23509 (N_23509,N_22499,N_22342);
nand U23510 (N_23510,N_21686,N_22017);
nor U23511 (N_23511,N_21964,N_22670);
or U23512 (N_23512,N_21971,N_22395);
and U23513 (N_23513,N_22720,N_22278);
nand U23514 (N_23514,N_22235,N_22657);
or U23515 (N_23515,N_22794,N_22769);
xnor U23516 (N_23516,N_22200,N_22641);
and U23517 (N_23517,N_21729,N_22350);
nand U23518 (N_23518,N_22218,N_22061);
nor U23519 (N_23519,N_21978,N_21761);
or U23520 (N_23520,N_22019,N_22658);
or U23521 (N_23521,N_21856,N_21795);
nand U23522 (N_23522,N_22596,N_21960);
nor U23523 (N_23523,N_22672,N_22102);
xnor U23524 (N_23524,N_22484,N_22411);
nor U23525 (N_23525,N_22560,N_22315);
nor U23526 (N_23526,N_22505,N_22111);
or U23527 (N_23527,N_22299,N_22504);
and U23528 (N_23528,N_22798,N_21844);
or U23529 (N_23529,N_21851,N_22041);
or U23530 (N_23530,N_22538,N_22432);
xor U23531 (N_23531,N_21809,N_22590);
xor U23532 (N_23532,N_22179,N_22244);
or U23533 (N_23533,N_22666,N_21741);
or U23534 (N_23534,N_22164,N_21802);
xnor U23535 (N_23535,N_22582,N_22702);
nor U23536 (N_23536,N_21942,N_22494);
nand U23537 (N_23537,N_22683,N_22445);
or U23538 (N_23538,N_22008,N_21998);
and U23539 (N_23539,N_22761,N_22419);
and U23540 (N_23540,N_22499,N_21802);
nand U23541 (N_23541,N_22751,N_21644);
and U23542 (N_23542,N_22684,N_21788);
nor U23543 (N_23543,N_21970,N_22627);
or U23544 (N_23544,N_22294,N_22522);
nand U23545 (N_23545,N_22773,N_21852);
and U23546 (N_23546,N_22373,N_22027);
nand U23547 (N_23547,N_22494,N_21974);
and U23548 (N_23548,N_22561,N_22471);
nand U23549 (N_23549,N_22669,N_22066);
or U23550 (N_23550,N_21605,N_22114);
xor U23551 (N_23551,N_22192,N_22554);
and U23552 (N_23552,N_22148,N_22683);
nor U23553 (N_23553,N_22303,N_21986);
and U23554 (N_23554,N_22486,N_22439);
and U23555 (N_23555,N_21988,N_22750);
or U23556 (N_23556,N_21961,N_22188);
nor U23557 (N_23557,N_22763,N_21754);
nor U23558 (N_23558,N_22004,N_21781);
and U23559 (N_23559,N_21964,N_21904);
xnor U23560 (N_23560,N_22448,N_21866);
xnor U23561 (N_23561,N_22532,N_22611);
nor U23562 (N_23562,N_22465,N_22725);
xnor U23563 (N_23563,N_22172,N_22088);
and U23564 (N_23564,N_22715,N_22785);
nor U23565 (N_23565,N_22406,N_22212);
or U23566 (N_23566,N_22290,N_21688);
nand U23567 (N_23567,N_22793,N_22372);
nand U23568 (N_23568,N_22765,N_21805);
xnor U23569 (N_23569,N_22523,N_22716);
and U23570 (N_23570,N_21910,N_22400);
xnor U23571 (N_23571,N_22462,N_21901);
nor U23572 (N_23572,N_21696,N_22413);
xnor U23573 (N_23573,N_22045,N_21829);
xnor U23574 (N_23574,N_22187,N_22580);
xor U23575 (N_23575,N_22546,N_22234);
or U23576 (N_23576,N_22391,N_22444);
nand U23577 (N_23577,N_22574,N_22630);
nand U23578 (N_23578,N_22553,N_21749);
nand U23579 (N_23579,N_22355,N_21998);
and U23580 (N_23580,N_22560,N_22333);
and U23581 (N_23581,N_22355,N_22552);
or U23582 (N_23582,N_22766,N_21805);
and U23583 (N_23583,N_22657,N_22591);
and U23584 (N_23584,N_22078,N_22646);
nand U23585 (N_23585,N_22274,N_22788);
xnor U23586 (N_23586,N_22493,N_22464);
or U23587 (N_23587,N_22328,N_22322);
or U23588 (N_23588,N_22724,N_22513);
and U23589 (N_23589,N_21887,N_21600);
and U23590 (N_23590,N_21841,N_22107);
nor U23591 (N_23591,N_22446,N_22518);
nor U23592 (N_23592,N_22606,N_22687);
and U23593 (N_23593,N_21662,N_21911);
nand U23594 (N_23594,N_21765,N_22638);
nand U23595 (N_23595,N_22560,N_21823);
and U23596 (N_23596,N_22587,N_21957);
xnor U23597 (N_23597,N_22285,N_21939);
and U23598 (N_23598,N_21902,N_22226);
nor U23599 (N_23599,N_22149,N_21914);
or U23600 (N_23600,N_22266,N_21893);
nor U23601 (N_23601,N_22486,N_21720);
or U23602 (N_23602,N_22721,N_22659);
or U23603 (N_23603,N_22299,N_22627);
and U23604 (N_23604,N_22319,N_21974);
nor U23605 (N_23605,N_21679,N_22356);
nor U23606 (N_23606,N_21655,N_22598);
nand U23607 (N_23607,N_21720,N_22124);
nor U23608 (N_23608,N_22422,N_21637);
xor U23609 (N_23609,N_21992,N_22338);
and U23610 (N_23610,N_21951,N_22628);
and U23611 (N_23611,N_21895,N_21996);
nor U23612 (N_23612,N_21819,N_21917);
nand U23613 (N_23613,N_21661,N_22038);
nand U23614 (N_23614,N_22442,N_21985);
nand U23615 (N_23615,N_22537,N_22315);
xnor U23616 (N_23616,N_22646,N_21782);
and U23617 (N_23617,N_22026,N_22535);
or U23618 (N_23618,N_22084,N_22511);
or U23619 (N_23619,N_22747,N_22601);
and U23620 (N_23620,N_22323,N_21833);
xnor U23621 (N_23621,N_21779,N_22352);
and U23622 (N_23622,N_22062,N_22043);
xor U23623 (N_23623,N_22681,N_22196);
and U23624 (N_23624,N_21708,N_21768);
nand U23625 (N_23625,N_22444,N_21624);
and U23626 (N_23626,N_22669,N_22429);
nand U23627 (N_23627,N_21834,N_22043);
nand U23628 (N_23628,N_22270,N_22652);
nand U23629 (N_23629,N_22035,N_22371);
xor U23630 (N_23630,N_22737,N_22544);
and U23631 (N_23631,N_21610,N_22349);
or U23632 (N_23632,N_22153,N_21679);
xnor U23633 (N_23633,N_22212,N_22126);
nand U23634 (N_23634,N_22410,N_21604);
and U23635 (N_23635,N_22394,N_21854);
and U23636 (N_23636,N_22426,N_22772);
and U23637 (N_23637,N_22783,N_21774);
xnor U23638 (N_23638,N_21976,N_22423);
nor U23639 (N_23639,N_22521,N_22003);
and U23640 (N_23640,N_22529,N_22515);
nand U23641 (N_23641,N_22095,N_22085);
nand U23642 (N_23642,N_22469,N_22122);
xor U23643 (N_23643,N_21668,N_22362);
and U23644 (N_23644,N_22785,N_21852);
nor U23645 (N_23645,N_21898,N_22517);
or U23646 (N_23646,N_22748,N_22454);
and U23647 (N_23647,N_22372,N_22649);
nand U23648 (N_23648,N_22311,N_22609);
xor U23649 (N_23649,N_21737,N_21861);
nand U23650 (N_23650,N_21845,N_22229);
nand U23651 (N_23651,N_22490,N_22253);
or U23652 (N_23652,N_22759,N_21869);
xor U23653 (N_23653,N_22013,N_22073);
and U23654 (N_23654,N_21647,N_22382);
nand U23655 (N_23655,N_22064,N_21879);
or U23656 (N_23656,N_22796,N_22281);
nand U23657 (N_23657,N_22556,N_21914);
nand U23658 (N_23658,N_21797,N_21988);
or U23659 (N_23659,N_22312,N_21869);
and U23660 (N_23660,N_21732,N_22557);
and U23661 (N_23661,N_22114,N_21945);
or U23662 (N_23662,N_22774,N_22301);
nor U23663 (N_23663,N_22644,N_21905);
and U23664 (N_23664,N_21648,N_21841);
or U23665 (N_23665,N_21928,N_22780);
and U23666 (N_23666,N_21890,N_21813);
nor U23667 (N_23667,N_21675,N_21823);
nand U23668 (N_23668,N_22468,N_21703);
or U23669 (N_23669,N_22405,N_21696);
and U23670 (N_23670,N_21678,N_21849);
nand U23671 (N_23671,N_22232,N_21749);
nor U23672 (N_23672,N_22684,N_22751);
nand U23673 (N_23673,N_21841,N_21926);
nor U23674 (N_23674,N_22710,N_22180);
nand U23675 (N_23675,N_22245,N_22416);
nor U23676 (N_23676,N_22725,N_22267);
nor U23677 (N_23677,N_22777,N_22160);
nor U23678 (N_23678,N_22056,N_22372);
and U23679 (N_23679,N_22342,N_22259);
and U23680 (N_23680,N_21971,N_22139);
xnor U23681 (N_23681,N_22325,N_22669);
nor U23682 (N_23682,N_22706,N_22368);
or U23683 (N_23683,N_22113,N_21899);
xnor U23684 (N_23684,N_21904,N_22411);
and U23685 (N_23685,N_22283,N_22659);
nor U23686 (N_23686,N_22750,N_22258);
and U23687 (N_23687,N_22569,N_22214);
or U23688 (N_23688,N_22710,N_22137);
nor U23689 (N_23689,N_22463,N_22036);
nor U23690 (N_23690,N_22430,N_21855);
or U23691 (N_23691,N_21908,N_21827);
nor U23692 (N_23692,N_21757,N_22766);
and U23693 (N_23693,N_22016,N_21720);
or U23694 (N_23694,N_22166,N_21724);
nor U23695 (N_23695,N_22750,N_21727);
xnor U23696 (N_23696,N_21784,N_22352);
nand U23697 (N_23697,N_22531,N_22693);
or U23698 (N_23698,N_21816,N_21863);
xor U23699 (N_23699,N_22223,N_22157);
xor U23700 (N_23700,N_22652,N_22412);
or U23701 (N_23701,N_22522,N_22444);
nand U23702 (N_23702,N_22152,N_21847);
nand U23703 (N_23703,N_22276,N_22051);
xnor U23704 (N_23704,N_22164,N_22084);
and U23705 (N_23705,N_22328,N_22669);
nand U23706 (N_23706,N_22520,N_21621);
nor U23707 (N_23707,N_22598,N_22233);
or U23708 (N_23708,N_22564,N_21761);
nor U23709 (N_23709,N_22666,N_21978);
nand U23710 (N_23710,N_21861,N_22640);
and U23711 (N_23711,N_21740,N_21624);
xor U23712 (N_23712,N_21679,N_22791);
nand U23713 (N_23713,N_21640,N_22251);
nor U23714 (N_23714,N_21768,N_21983);
nand U23715 (N_23715,N_22035,N_22483);
xnor U23716 (N_23716,N_22203,N_22088);
xor U23717 (N_23717,N_22446,N_22521);
nor U23718 (N_23718,N_21796,N_21949);
nand U23719 (N_23719,N_22115,N_22314);
nor U23720 (N_23720,N_22218,N_22682);
or U23721 (N_23721,N_22399,N_21957);
or U23722 (N_23722,N_22378,N_22653);
xnor U23723 (N_23723,N_22609,N_21891);
xnor U23724 (N_23724,N_21856,N_22476);
nor U23725 (N_23725,N_21860,N_21863);
xnor U23726 (N_23726,N_22515,N_22474);
xnor U23727 (N_23727,N_22740,N_22034);
nand U23728 (N_23728,N_22079,N_22403);
nand U23729 (N_23729,N_21758,N_22349);
xor U23730 (N_23730,N_21865,N_21611);
nor U23731 (N_23731,N_22522,N_22756);
xor U23732 (N_23732,N_21939,N_21839);
or U23733 (N_23733,N_22768,N_22095);
nand U23734 (N_23734,N_21695,N_22791);
and U23735 (N_23735,N_22125,N_22508);
nand U23736 (N_23736,N_22651,N_22129);
nand U23737 (N_23737,N_22712,N_22067);
nand U23738 (N_23738,N_22364,N_21912);
and U23739 (N_23739,N_22018,N_21854);
nor U23740 (N_23740,N_22508,N_22592);
xnor U23741 (N_23741,N_21752,N_22451);
nor U23742 (N_23742,N_22708,N_21738);
and U23743 (N_23743,N_21929,N_22320);
nor U23744 (N_23744,N_22780,N_22715);
xnor U23745 (N_23745,N_22765,N_22318);
and U23746 (N_23746,N_22295,N_22684);
nand U23747 (N_23747,N_21702,N_22190);
and U23748 (N_23748,N_22518,N_21602);
nand U23749 (N_23749,N_22480,N_22489);
xor U23750 (N_23750,N_22799,N_22183);
and U23751 (N_23751,N_21995,N_22302);
and U23752 (N_23752,N_21786,N_22341);
and U23753 (N_23753,N_22105,N_22174);
and U23754 (N_23754,N_22278,N_22559);
or U23755 (N_23755,N_22159,N_21661);
and U23756 (N_23756,N_22608,N_22436);
or U23757 (N_23757,N_21754,N_22748);
xor U23758 (N_23758,N_22063,N_22048);
xnor U23759 (N_23759,N_22472,N_21877);
and U23760 (N_23760,N_21617,N_21750);
or U23761 (N_23761,N_21996,N_21612);
and U23762 (N_23762,N_22767,N_22148);
and U23763 (N_23763,N_22744,N_21791);
nand U23764 (N_23764,N_22527,N_22242);
nand U23765 (N_23765,N_21808,N_22087);
or U23766 (N_23766,N_22016,N_22076);
nand U23767 (N_23767,N_22432,N_22412);
nor U23768 (N_23768,N_22231,N_21673);
or U23769 (N_23769,N_22543,N_21926);
xnor U23770 (N_23770,N_22323,N_21850);
nand U23771 (N_23771,N_22201,N_21742);
nand U23772 (N_23772,N_22113,N_21735);
and U23773 (N_23773,N_22168,N_21897);
xor U23774 (N_23774,N_22583,N_22408);
xnor U23775 (N_23775,N_22546,N_21920);
and U23776 (N_23776,N_22100,N_21735);
nor U23777 (N_23777,N_21782,N_22566);
xnor U23778 (N_23778,N_21877,N_22617);
nor U23779 (N_23779,N_22105,N_22267);
nand U23780 (N_23780,N_22286,N_22402);
and U23781 (N_23781,N_21987,N_22156);
and U23782 (N_23782,N_22186,N_22484);
nand U23783 (N_23783,N_22770,N_22341);
nand U23784 (N_23784,N_21724,N_22218);
nor U23785 (N_23785,N_21957,N_22288);
xor U23786 (N_23786,N_22232,N_21625);
and U23787 (N_23787,N_21755,N_21799);
or U23788 (N_23788,N_22267,N_21804);
nor U23789 (N_23789,N_21741,N_22061);
or U23790 (N_23790,N_21887,N_22023);
xor U23791 (N_23791,N_22010,N_22640);
and U23792 (N_23792,N_22757,N_22508);
nand U23793 (N_23793,N_22372,N_22433);
or U23794 (N_23794,N_22310,N_22142);
nor U23795 (N_23795,N_21936,N_22511);
nand U23796 (N_23796,N_21657,N_22144);
xor U23797 (N_23797,N_21904,N_21804);
nor U23798 (N_23798,N_22578,N_22237);
or U23799 (N_23799,N_22067,N_22718);
nand U23800 (N_23800,N_21787,N_22715);
xor U23801 (N_23801,N_22626,N_21777);
nor U23802 (N_23802,N_21756,N_22324);
or U23803 (N_23803,N_22652,N_22087);
and U23804 (N_23804,N_21609,N_21962);
nand U23805 (N_23805,N_21791,N_21976);
xor U23806 (N_23806,N_22230,N_21819);
nor U23807 (N_23807,N_22484,N_21616);
nand U23808 (N_23808,N_21822,N_22766);
nand U23809 (N_23809,N_21821,N_22343);
or U23810 (N_23810,N_22113,N_22551);
and U23811 (N_23811,N_22109,N_21960);
nor U23812 (N_23812,N_22366,N_21995);
nand U23813 (N_23813,N_22631,N_22178);
nand U23814 (N_23814,N_21632,N_22758);
xor U23815 (N_23815,N_22750,N_22797);
and U23816 (N_23816,N_21862,N_22248);
or U23817 (N_23817,N_21951,N_21862);
xor U23818 (N_23818,N_22658,N_22601);
and U23819 (N_23819,N_21973,N_21791);
nand U23820 (N_23820,N_22411,N_22346);
xnor U23821 (N_23821,N_22756,N_21823);
nor U23822 (N_23822,N_22133,N_21669);
nand U23823 (N_23823,N_21720,N_21743);
nand U23824 (N_23824,N_22249,N_21818);
and U23825 (N_23825,N_22516,N_22590);
xnor U23826 (N_23826,N_22534,N_21784);
xnor U23827 (N_23827,N_21736,N_21827);
xor U23828 (N_23828,N_22621,N_21778);
or U23829 (N_23829,N_21910,N_21701);
and U23830 (N_23830,N_22691,N_22336);
xor U23831 (N_23831,N_22777,N_22454);
nor U23832 (N_23832,N_22652,N_22517);
or U23833 (N_23833,N_21732,N_21959);
and U23834 (N_23834,N_22387,N_21701);
or U23835 (N_23835,N_22100,N_21846);
nor U23836 (N_23836,N_21877,N_22297);
or U23837 (N_23837,N_22229,N_22593);
and U23838 (N_23838,N_22505,N_22561);
or U23839 (N_23839,N_22102,N_21854);
nor U23840 (N_23840,N_21745,N_22632);
and U23841 (N_23841,N_22557,N_22056);
and U23842 (N_23842,N_22262,N_22019);
nor U23843 (N_23843,N_22694,N_22155);
nor U23844 (N_23844,N_22753,N_22589);
nor U23845 (N_23845,N_22092,N_22396);
and U23846 (N_23846,N_22473,N_22065);
or U23847 (N_23847,N_22507,N_22617);
nand U23848 (N_23848,N_22499,N_22272);
or U23849 (N_23849,N_21653,N_21619);
nor U23850 (N_23850,N_21716,N_22144);
xnor U23851 (N_23851,N_22600,N_21680);
nand U23852 (N_23852,N_22175,N_22211);
xor U23853 (N_23853,N_21748,N_21635);
nor U23854 (N_23854,N_22125,N_22589);
or U23855 (N_23855,N_21675,N_21741);
and U23856 (N_23856,N_22269,N_22197);
or U23857 (N_23857,N_21981,N_21856);
xnor U23858 (N_23858,N_22666,N_22245);
nand U23859 (N_23859,N_21720,N_22243);
nor U23860 (N_23860,N_22214,N_22357);
and U23861 (N_23861,N_22584,N_22680);
nor U23862 (N_23862,N_22018,N_21695);
nand U23863 (N_23863,N_22619,N_21908);
xor U23864 (N_23864,N_21905,N_21627);
or U23865 (N_23865,N_21676,N_21846);
and U23866 (N_23866,N_22019,N_21980);
and U23867 (N_23867,N_21620,N_22080);
nand U23868 (N_23868,N_22492,N_22675);
and U23869 (N_23869,N_22477,N_21706);
nor U23870 (N_23870,N_22204,N_21780);
nand U23871 (N_23871,N_22305,N_21770);
nand U23872 (N_23872,N_22489,N_22407);
nand U23873 (N_23873,N_22508,N_22416);
nor U23874 (N_23874,N_22438,N_21782);
xor U23875 (N_23875,N_22488,N_22537);
nand U23876 (N_23876,N_22002,N_22260);
nor U23877 (N_23877,N_22754,N_21624);
xor U23878 (N_23878,N_22731,N_22428);
or U23879 (N_23879,N_21734,N_22114);
xnor U23880 (N_23880,N_22063,N_21688);
xnor U23881 (N_23881,N_21865,N_22497);
or U23882 (N_23882,N_22793,N_22515);
or U23883 (N_23883,N_22133,N_22062);
nand U23884 (N_23884,N_22124,N_21711);
nand U23885 (N_23885,N_22128,N_21947);
nor U23886 (N_23886,N_22059,N_22313);
nor U23887 (N_23887,N_22200,N_21949);
nand U23888 (N_23888,N_22002,N_21744);
xnor U23889 (N_23889,N_21855,N_21965);
or U23890 (N_23890,N_21736,N_21708);
or U23891 (N_23891,N_21972,N_22403);
or U23892 (N_23892,N_22577,N_22570);
or U23893 (N_23893,N_21708,N_22024);
nor U23894 (N_23894,N_21966,N_22270);
or U23895 (N_23895,N_22451,N_21719);
and U23896 (N_23896,N_22072,N_21989);
xor U23897 (N_23897,N_21786,N_21794);
or U23898 (N_23898,N_21706,N_21613);
nor U23899 (N_23899,N_21601,N_22135);
nand U23900 (N_23900,N_21984,N_22050);
nor U23901 (N_23901,N_21811,N_22369);
nand U23902 (N_23902,N_21881,N_21993);
nand U23903 (N_23903,N_22596,N_22590);
xor U23904 (N_23904,N_22112,N_22383);
nand U23905 (N_23905,N_22778,N_22586);
and U23906 (N_23906,N_22601,N_21909);
nor U23907 (N_23907,N_21796,N_22112);
nand U23908 (N_23908,N_22278,N_21918);
nor U23909 (N_23909,N_22527,N_22449);
or U23910 (N_23910,N_22433,N_22317);
nor U23911 (N_23911,N_22221,N_21670);
nor U23912 (N_23912,N_22352,N_22126);
nand U23913 (N_23913,N_22730,N_22005);
or U23914 (N_23914,N_21939,N_22032);
xor U23915 (N_23915,N_22067,N_22324);
xor U23916 (N_23916,N_22641,N_22749);
nor U23917 (N_23917,N_21977,N_22035);
nand U23918 (N_23918,N_22152,N_22067);
and U23919 (N_23919,N_21798,N_22467);
xnor U23920 (N_23920,N_22496,N_21628);
nand U23921 (N_23921,N_21872,N_22234);
or U23922 (N_23922,N_22670,N_22013);
xor U23923 (N_23923,N_21706,N_21773);
nor U23924 (N_23924,N_22724,N_22090);
and U23925 (N_23925,N_22326,N_22001);
nor U23926 (N_23926,N_22044,N_22759);
nor U23927 (N_23927,N_22078,N_22133);
or U23928 (N_23928,N_22597,N_22082);
nor U23929 (N_23929,N_22691,N_21900);
nand U23930 (N_23930,N_22653,N_22389);
nor U23931 (N_23931,N_22783,N_22400);
nand U23932 (N_23932,N_22052,N_22267);
xor U23933 (N_23933,N_22462,N_21716);
xnor U23934 (N_23934,N_21602,N_22401);
nor U23935 (N_23935,N_22505,N_21842);
xnor U23936 (N_23936,N_21773,N_21615);
or U23937 (N_23937,N_21673,N_22191);
and U23938 (N_23938,N_21885,N_22559);
nor U23939 (N_23939,N_22134,N_21766);
or U23940 (N_23940,N_22292,N_22025);
nand U23941 (N_23941,N_22488,N_22225);
nand U23942 (N_23942,N_21975,N_22018);
nor U23943 (N_23943,N_22337,N_22457);
nor U23944 (N_23944,N_22382,N_21746);
and U23945 (N_23945,N_22735,N_21923);
nor U23946 (N_23946,N_22453,N_21680);
xor U23947 (N_23947,N_21716,N_22506);
and U23948 (N_23948,N_22300,N_21742);
nand U23949 (N_23949,N_22492,N_22149);
or U23950 (N_23950,N_22336,N_22218);
nor U23951 (N_23951,N_22784,N_22739);
or U23952 (N_23952,N_22347,N_21934);
and U23953 (N_23953,N_22278,N_21748);
and U23954 (N_23954,N_22334,N_22195);
or U23955 (N_23955,N_21952,N_22066);
xnor U23956 (N_23956,N_22249,N_22623);
and U23957 (N_23957,N_22171,N_21932);
xor U23958 (N_23958,N_22289,N_22494);
and U23959 (N_23959,N_22685,N_22536);
nor U23960 (N_23960,N_22744,N_21892);
xor U23961 (N_23961,N_22502,N_21614);
xnor U23962 (N_23962,N_22657,N_22583);
nand U23963 (N_23963,N_22631,N_21916);
and U23964 (N_23964,N_22568,N_21734);
xor U23965 (N_23965,N_22252,N_22562);
and U23966 (N_23966,N_22030,N_22483);
nor U23967 (N_23967,N_22453,N_21854);
xnor U23968 (N_23968,N_21755,N_22637);
nand U23969 (N_23969,N_22608,N_21693);
or U23970 (N_23970,N_21936,N_22252);
and U23971 (N_23971,N_22282,N_22527);
xor U23972 (N_23972,N_22095,N_22665);
or U23973 (N_23973,N_22753,N_22479);
and U23974 (N_23974,N_22755,N_22633);
xor U23975 (N_23975,N_22767,N_22577);
xor U23976 (N_23976,N_22305,N_22739);
nand U23977 (N_23977,N_22454,N_21834);
nor U23978 (N_23978,N_22628,N_21636);
nor U23979 (N_23979,N_21875,N_22567);
xnor U23980 (N_23980,N_22098,N_21757);
or U23981 (N_23981,N_22421,N_21982);
xor U23982 (N_23982,N_21661,N_22748);
or U23983 (N_23983,N_21613,N_22245);
and U23984 (N_23984,N_21838,N_22535);
xnor U23985 (N_23985,N_22100,N_22752);
nor U23986 (N_23986,N_21712,N_22241);
nand U23987 (N_23987,N_22436,N_21775);
nand U23988 (N_23988,N_22691,N_22510);
nand U23989 (N_23989,N_22693,N_21684);
xor U23990 (N_23990,N_21695,N_22113);
nand U23991 (N_23991,N_22096,N_22565);
nand U23992 (N_23992,N_22269,N_22566);
nand U23993 (N_23993,N_21867,N_22015);
xor U23994 (N_23994,N_22450,N_21874);
nand U23995 (N_23995,N_22196,N_21987);
or U23996 (N_23996,N_22067,N_21629);
and U23997 (N_23997,N_22301,N_22053);
nand U23998 (N_23998,N_22496,N_22644);
xnor U23999 (N_23999,N_22116,N_22646);
and U24000 (N_24000,N_23569,N_23834);
xor U24001 (N_24001,N_23731,N_23232);
or U24002 (N_24002,N_23698,N_22991);
and U24003 (N_24003,N_23587,N_23685);
or U24004 (N_24004,N_23175,N_23634);
and U24005 (N_24005,N_22977,N_23292);
or U24006 (N_24006,N_22829,N_23545);
nand U24007 (N_24007,N_23517,N_22812);
nor U24008 (N_24008,N_22915,N_23049);
and U24009 (N_24009,N_23404,N_23480);
and U24010 (N_24010,N_23307,N_23219);
xor U24011 (N_24011,N_23181,N_23191);
and U24012 (N_24012,N_23659,N_22850);
nand U24013 (N_24013,N_23646,N_23141);
or U24014 (N_24014,N_23625,N_23788);
nand U24015 (N_24015,N_23862,N_23154);
nor U24016 (N_24016,N_23257,N_22896);
nor U24017 (N_24017,N_23782,N_23763);
nand U24018 (N_24018,N_22807,N_23573);
or U24019 (N_24019,N_23362,N_23614);
or U24020 (N_24020,N_22937,N_22941);
xnor U24021 (N_24021,N_23906,N_23789);
nand U24022 (N_24022,N_23543,N_23740);
xnor U24023 (N_24023,N_22943,N_23687);
xor U24024 (N_24024,N_23928,N_23552);
and U24025 (N_24025,N_23145,N_23468);
xnor U24026 (N_24026,N_23952,N_22962);
or U24027 (N_24027,N_23550,N_23341);
nor U24028 (N_24028,N_23123,N_23994);
nand U24029 (N_24029,N_22847,N_22894);
and U24030 (N_24030,N_23412,N_23287);
and U24031 (N_24031,N_23559,N_23425);
nand U24032 (N_24032,N_22806,N_22944);
nor U24033 (N_24033,N_23302,N_23147);
and U24034 (N_24034,N_22920,N_23028);
nor U24035 (N_24035,N_22947,N_23456);
and U24036 (N_24036,N_23273,N_23156);
nand U24037 (N_24037,N_23907,N_23411);
and U24038 (N_24038,N_23690,N_23136);
and U24039 (N_24039,N_23865,N_23567);
and U24040 (N_24040,N_23955,N_23976);
nand U24041 (N_24041,N_23266,N_23553);
xnor U24042 (N_24042,N_23716,N_23923);
xor U24043 (N_24043,N_22934,N_23329);
xor U24044 (N_24044,N_23605,N_23324);
nand U24045 (N_24045,N_22816,N_23762);
or U24046 (N_24046,N_23124,N_23854);
and U24047 (N_24047,N_23713,N_23968);
or U24048 (N_24048,N_22957,N_23382);
nand U24049 (N_24049,N_23228,N_23889);
and U24050 (N_24050,N_23664,N_23325);
nand U24051 (N_24051,N_22830,N_23348);
nor U24052 (N_24052,N_22835,N_23381);
and U24053 (N_24053,N_23594,N_23650);
xor U24054 (N_24054,N_23338,N_23901);
nor U24055 (N_24055,N_22895,N_23128);
nor U24056 (N_24056,N_23784,N_23490);
or U24057 (N_24057,N_23327,N_23530);
or U24058 (N_24058,N_23422,N_23774);
nand U24059 (N_24059,N_23632,N_23830);
nor U24060 (N_24060,N_23921,N_23790);
nand U24061 (N_24061,N_23982,N_23286);
nor U24062 (N_24062,N_23804,N_23355);
nand U24063 (N_24063,N_23255,N_22903);
xnor U24064 (N_24064,N_23139,N_22888);
and U24065 (N_24065,N_23610,N_23019);
nand U24066 (N_24066,N_23903,N_23845);
or U24067 (N_24067,N_23958,N_23132);
xor U24068 (N_24068,N_23729,N_23322);
and U24069 (N_24069,N_23462,N_23225);
nand U24070 (N_24070,N_23236,N_22993);
or U24071 (N_24071,N_23583,N_23313);
or U24072 (N_24072,N_23663,N_23146);
or U24073 (N_24073,N_23829,N_23205);
xnor U24074 (N_24074,N_22839,N_23498);
xnor U24075 (N_24075,N_23764,N_23642);
nor U24076 (N_24076,N_23083,N_22908);
nor U24077 (N_24077,N_23344,N_23105);
nand U24078 (N_24078,N_22838,N_23542);
nand U24079 (N_24079,N_22971,N_23566);
xnor U24080 (N_24080,N_23768,N_22906);
nand U24081 (N_24081,N_23844,N_22942);
nor U24082 (N_24082,N_23990,N_23004);
xnor U24083 (N_24083,N_23176,N_23673);
xnor U24084 (N_24084,N_23372,N_23174);
or U24085 (N_24085,N_23524,N_23827);
and U24086 (N_24086,N_23905,N_23821);
and U24087 (N_24087,N_23479,N_23656);
nand U24088 (N_24088,N_23939,N_23218);
nor U24089 (N_24089,N_23051,N_22960);
xor U24090 (N_24090,N_23024,N_23691);
xnor U24091 (N_24091,N_23860,N_23935);
nor U24092 (N_24092,N_23626,N_23967);
nor U24093 (N_24093,N_23592,N_23651);
or U24094 (N_24094,N_23135,N_23604);
or U24095 (N_24095,N_23560,N_23746);
xnor U24096 (N_24096,N_23142,N_22998);
and U24097 (N_24097,N_23018,N_23442);
nand U24098 (N_24098,N_23308,N_23525);
nand U24099 (N_24099,N_23930,N_22911);
nor U24100 (N_24100,N_23234,N_23109);
xor U24101 (N_24101,N_23365,N_23636);
or U24102 (N_24102,N_23577,N_23808);
nand U24103 (N_24103,N_23861,N_23361);
and U24104 (N_24104,N_23783,N_23470);
xor U24105 (N_24105,N_23532,N_23943);
nor U24106 (N_24106,N_23813,N_23516);
and U24107 (N_24107,N_23162,N_23841);
xor U24108 (N_24108,N_23239,N_23495);
xnor U24109 (N_24109,N_23483,N_23544);
nor U24110 (N_24110,N_23346,N_23256);
nand U24111 (N_24111,N_23669,N_23373);
and U24112 (N_24112,N_23333,N_23631);
and U24113 (N_24113,N_23590,N_22930);
xnor U24114 (N_24114,N_23416,N_23714);
and U24115 (N_24115,N_23364,N_23948);
and U24116 (N_24116,N_23817,N_23866);
nor U24117 (N_24117,N_23536,N_23117);
xnor U24118 (N_24118,N_23877,N_23771);
nand U24119 (N_24119,N_23607,N_23407);
nor U24120 (N_24120,N_23087,N_23814);
nand U24121 (N_24121,N_23765,N_22865);
or U24122 (N_24122,N_22872,N_23189);
nor U24123 (N_24123,N_23144,N_23250);
nand U24124 (N_24124,N_23600,N_23337);
nor U24125 (N_24125,N_23437,N_23689);
and U24126 (N_24126,N_23017,N_23005);
xor U24127 (N_24127,N_23606,N_23944);
nor U24128 (N_24128,N_23751,N_23535);
and U24129 (N_24129,N_23737,N_23091);
nor U24130 (N_24130,N_23027,N_23107);
or U24131 (N_24131,N_23114,N_23227);
and U24132 (N_24132,N_23038,N_23041);
or U24133 (N_24133,N_23248,N_23247);
xor U24134 (N_24134,N_23125,N_23163);
or U24135 (N_24135,N_23196,N_23067);
nor U24136 (N_24136,N_23528,N_23056);
or U24137 (N_24137,N_23747,N_23439);
nor U24138 (N_24138,N_23133,N_22926);
xor U24139 (N_24139,N_23658,N_22973);
or U24140 (N_24140,N_23812,N_23207);
xnor U24141 (N_24141,N_23303,N_23305);
or U24142 (N_24142,N_23596,N_23068);
or U24143 (N_24143,N_23758,N_23561);
nor U24144 (N_24144,N_22965,N_23756);
nor U24145 (N_24145,N_23319,N_22883);
nor U24146 (N_24146,N_22881,N_23203);
or U24147 (N_24147,N_22999,N_23315);
or U24148 (N_24148,N_23786,N_23356);
or U24149 (N_24149,N_23261,N_23281);
xor U24150 (N_24150,N_23855,N_23720);
or U24151 (N_24151,N_23167,N_22952);
nand U24152 (N_24152,N_22876,N_23274);
nor U24153 (N_24153,N_23973,N_23643);
and U24154 (N_24154,N_23288,N_23321);
and U24155 (N_24155,N_23276,N_22870);
xor U24156 (N_24156,N_23182,N_23795);
and U24157 (N_24157,N_23127,N_23892);
or U24158 (N_24158,N_23800,N_23179);
nor U24159 (N_24159,N_23157,N_23031);
and U24160 (N_24160,N_23963,N_23194);
nor U24161 (N_24161,N_23421,N_23195);
and U24162 (N_24162,N_23826,N_22842);
xor U24163 (N_24163,N_22904,N_22938);
nor U24164 (N_24164,N_23260,N_22820);
xnor U24165 (N_24165,N_23020,N_23742);
nor U24166 (N_24166,N_23897,N_23187);
and U24167 (N_24167,N_22809,N_23847);
or U24168 (N_24168,N_23832,N_22992);
nor U24169 (N_24169,N_23956,N_23471);
nand U24170 (N_24170,N_23200,N_23204);
or U24171 (N_24171,N_23211,N_23933);
nand U24172 (N_24172,N_23766,N_23754);
nand U24173 (N_24173,N_23100,N_23042);
and U24174 (N_24174,N_23738,N_23909);
nor U24175 (N_24175,N_23574,N_23352);
and U24176 (N_24176,N_23870,N_22914);
xnor U24177 (N_24177,N_23715,N_23620);
nor U24178 (N_24178,N_22929,N_23655);
or U24179 (N_24179,N_23730,N_23971);
and U24180 (N_24180,N_23780,N_23989);
or U24181 (N_24181,N_22893,N_23104);
and U24182 (N_24182,N_23012,N_23022);
nor U24183 (N_24183,N_23705,N_23445);
nor U24184 (N_24184,N_23824,N_22964);
nor U24185 (N_24185,N_23876,N_23394);
nand U24186 (N_24186,N_23076,N_23032);
nand U24187 (N_24187,N_22860,N_23945);
nor U24188 (N_24188,N_23568,N_23190);
xor U24189 (N_24189,N_23084,N_23922);
nand U24190 (N_24190,N_23541,N_23192);
or U24191 (N_24191,N_23527,N_23521);
xnor U24192 (N_24192,N_22846,N_22863);
or U24193 (N_24193,N_23092,N_23660);
or U24194 (N_24194,N_22931,N_23781);
or U24195 (N_24195,N_23972,N_23458);
and U24196 (N_24196,N_23297,N_23229);
xnor U24197 (N_24197,N_23061,N_23953);
nor U24198 (N_24198,N_22825,N_23271);
or U24199 (N_24199,N_23052,N_23172);
nor U24200 (N_24200,N_23551,N_22844);
and U24201 (N_24201,N_23682,N_23898);
xor U24202 (N_24202,N_23666,N_22880);
nor U24203 (N_24203,N_23074,N_23579);
and U24204 (N_24204,N_23243,N_22967);
xnor U24205 (N_24205,N_23453,N_23602);
or U24206 (N_24206,N_23010,N_23883);
and U24207 (N_24207,N_23961,N_23785);
nand U24208 (N_24208,N_23799,N_23881);
xor U24209 (N_24209,N_22921,N_23252);
nor U24210 (N_24210,N_23908,N_23148);
and U24211 (N_24211,N_22961,N_23809);
xnor U24212 (N_24212,N_23098,N_23197);
nand U24213 (N_24213,N_23949,N_23102);
xnor U24214 (N_24214,N_23289,N_22946);
or U24215 (N_24215,N_22955,N_22995);
xnor U24216 (N_24216,N_23978,N_23853);
nand U24217 (N_24217,N_23485,N_22935);
xnor U24218 (N_24218,N_23149,N_23431);
nor U24219 (N_24219,N_23680,N_23222);
and U24220 (N_24220,N_23003,N_23641);
or U24221 (N_24221,N_23937,N_23695);
nand U24222 (N_24222,N_23522,N_23706);
nand U24223 (N_24223,N_23753,N_23053);
or U24224 (N_24224,N_23242,N_23093);
or U24225 (N_24225,N_22912,N_23246);
and U24226 (N_24226,N_23387,N_23184);
and U24227 (N_24227,N_23318,N_23259);
and U24228 (N_24228,N_22933,N_23671);
nand U24229 (N_24229,N_23931,N_23419);
or U24230 (N_24230,N_22916,N_23386);
and U24231 (N_24231,N_23688,N_23777);
nor U24232 (N_24232,N_23513,N_23088);
nand U24233 (N_24233,N_23489,N_23836);
and U24234 (N_24234,N_22875,N_23349);
nand U24235 (N_24235,N_23538,N_22808);
and U24236 (N_24236,N_22997,N_23393);
nand U24237 (N_24237,N_23484,N_23755);
nand U24238 (N_24238,N_23492,N_23794);
nand U24239 (N_24239,N_22856,N_23741);
nand U24240 (N_24240,N_23676,N_23622);
nand U24241 (N_24241,N_22976,N_23558);
nor U24242 (N_24242,N_22840,N_23153);
nand U24243 (N_24243,N_22919,N_22996);
and U24244 (N_24244,N_23472,N_23661);
xor U24245 (N_24245,N_23769,N_23383);
and U24246 (N_24246,N_23959,N_23725);
nand U24247 (N_24247,N_23727,N_23748);
or U24248 (N_24248,N_23993,N_23301);
xor U24249 (N_24249,N_23385,N_23299);
nand U24250 (N_24250,N_22887,N_23418);
nor U24251 (N_24251,N_23612,N_23166);
xor U24252 (N_24252,N_23262,N_23708);
or U24253 (N_24253,N_23206,N_22864);
and U24254 (N_24254,N_23406,N_23090);
nand U24255 (N_24255,N_23185,N_23593);
and U24256 (N_24256,N_23752,N_23272);
xnor U24257 (N_24257,N_23793,N_23050);
or U24258 (N_24258,N_23835,N_23035);
xor U24259 (N_24259,N_23168,N_23888);
nor U24260 (N_24260,N_23183,N_23328);
nor U24261 (N_24261,N_23169,N_23571);
or U24262 (N_24262,N_23849,N_23595);
xor U24263 (N_24263,N_23900,N_23432);
and U24264 (N_24264,N_23890,N_23662);
or U24265 (N_24265,N_23389,N_22802);
nor U24266 (N_24266,N_23778,N_23858);
or U24267 (N_24267,N_22824,N_23792);
or U24268 (N_24268,N_22974,N_23693);
nand U24269 (N_24269,N_23405,N_22994);
xor U24270 (N_24270,N_23438,N_22859);
xnor U24271 (N_24271,N_23801,N_23354);
nand U24272 (N_24272,N_23697,N_23351);
or U24273 (N_24273,N_22956,N_23488);
nand U24274 (N_24274,N_23036,N_22862);
nor U24275 (N_24275,N_23531,N_23224);
nor U24276 (N_24276,N_22833,N_23268);
xor U24277 (N_24277,N_23216,N_23506);
nor U24278 (N_24278,N_23529,N_23429);
or U24279 (N_24279,N_23282,N_23370);
nor U24280 (N_24280,N_23657,N_23369);
nor U24281 (N_24281,N_23350,N_23494);
nor U24282 (N_24282,N_23734,N_22918);
nor U24283 (N_24283,N_23767,N_23095);
xnor U24284 (N_24284,N_23649,N_23712);
xnor U24285 (N_24285,N_23624,N_23859);
xor U24286 (N_24286,N_23565,N_23611);
or U24287 (N_24287,N_23724,N_22985);
or U24288 (N_24288,N_23681,N_23415);
xnor U24289 (N_24289,N_23121,N_23178);
and U24290 (N_24290,N_23408,N_23508);
nor U24291 (N_24291,N_23015,N_23704);
or U24292 (N_24292,N_23291,N_23384);
or U24293 (N_24293,N_23233,N_23628);
xnor U24294 (N_24294,N_23796,N_23444);
and U24295 (N_24295,N_23000,N_23465);
nand U24296 (N_24296,N_23214,N_23913);
or U24297 (N_24297,N_23016,N_23891);
xor U24298 (N_24298,N_23736,N_23810);
and U24299 (N_24299,N_22923,N_23115);
or U24300 (N_24300,N_23779,N_23576);
xor U24301 (N_24301,N_23300,N_22886);
nand U24302 (N_24302,N_22917,N_23330);
xnor U24303 (N_24303,N_23879,N_23077);
and U24304 (N_24304,N_23629,N_23221);
xnor U24305 (N_24305,N_23791,N_23509);
nand U24306 (N_24306,N_22907,N_22814);
or U24307 (N_24307,N_23451,N_23507);
nor U24308 (N_24308,N_22925,N_23505);
and U24309 (N_24309,N_23882,N_23639);
nand U24310 (N_24310,N_22975,N_22803);
nor U24311 (N_24311,N_23520,N_22811);
or U24312 (N_24312,N_23874,N_23208);
nor U24313 (N_24313,N_23343,N_23433);
or U24314 (N_24314,N_23820,N_23633);
or U24315 (N_24315,N_23414,N_23150);
nand U24316 (N_24316,N_22854,N_23430);
nand U24317 (N_24317,N_22902,N_23304);
nor U24318 (N_24318,N_23001,N_23951);
xnor U24319 (N_24319,N_23034,N_23376);
nor U24320 (N_24320,N_23924,N_23375);
nand U24321 (N_24321,N_22804,N_23739);
nand U24322 (N_24322,N_23549,N_23267);
xor U24323 (N_24323,N_23895,N_23991);
xor U24324 (N_24324,N_23914,N_23811);
or U24325 (N_24325,N_23173,N_22932);
xor U24326 (N_24326,N_22892,N_23409);
xnor U24327 (N_24327,N_23040,N_23140);
and U24328 (N_24328,N_23526,N_23942);
and U24329 (N_24329,N_22986,N_23899);
nand U24330 (N_24330,N_23210,N_23202);
xor U24331 (N_24331,N_23188,N_22866);
nand U24332 (N_24332,N_23608,N_22936);
or U24333 (N_24333,N_23402,N_23058);
and U24334 (N_24334,N_23496,N_23932);
xnor U24335 (N_24335,N_23316,N_23692);
and U24336 (N_24336,N_22905,N_23744);
xnor U24337 (N_24337,N_23047,N_22951);
or U24338 (N_24338,N_23941,N_23966);
nor U24339 (N_24339,N_23699,N_23723);
nand U24340 (N_24340,N_22899,N_22900);
xor U24341 (N_24341,N_22948,N_23078);
or U24342 (N_24342,N_23648,N_23613);
nor U24343 (N_24343,N_23245,N_22877);
nand U24344 (N_24344,N_23554,N_23589);
and U24345 (N_24345,N_23735,N_22958);
or U24346 (N_24346,N_23452,N_23390);
nand U24347 (N_24347,N_23395,N_23293);
nand U24348 (N_24348,N_23819,N_22874);
and U24349 (N_24349,N_23749,N_23701);
and U24350 (N_24350,N_23597,N_23802);
nand U24351 (N_24351,N_23223,N_23435);
nor U24352 (N_24352,N_22982,N_23118);
or U24353 (N_24353,N_23843,N_23391);
nand U24354 (N_24354,N_23326,N_23013);
and U24355 (N_24355,N_22970,N_23379);
and U24356 (N_24356,N_23073,N_22909);
or U24357 (N_24357,N_23129,N_23339);
nor U24358 (N_24358,N_23677,N_23424);
nand U24359 (N_24359,N_23071,N_23938);
nor U24360 (N_24360,N_23099,N_23220);
xnor U24361 (N_24361,N_23537,N_23198);
nand U24362 (N_24362,N_23707,N_23918);
nand U24363 (N_24363,N_23872,N_23226);
nand U24364 (N_24364,N_23732,N_22805);
or U24365 (N_24365,N_23066,N_23059);
nand U24366 (N_24366,N_23464,N_22858);
nand U24367 (N_24367,N_22949,N_23534);
nand U24368 (N_24368,N_23467,N_23331);
or U24369 (N_24369,N_22836,N_23743);
xnor U24370 (N_24370,N_23884,N_23992);
and U24371 (N_24371,N_23413,N_23335);
xnor U24372 (N_24372,N_22940,N_23652);
or U24373 (N_24373,N_23591,N_23665);
xor U24374 (N_24374,N_23647,N_23023);
and U24375 (N_24375,N_23045,N_23450);
nor U24376 (N_24376,N_23640,N_23987);
or U24377 (N_24377,N_23670,N_23251);
nor U24378 (N_24378,N_23816,N_23598);
nand U24379 (N_24379,N_23722,N_23919);
or U24380 (N_24380,N_22924,N_23998);
or U24381 (N_24381,N_23025,N_23295);
or U24382 (N_24382,N_23773,N_23249);
and U24383 (N_24383,N_23116,N_23500);
xor U24384 (N_24384,N_22978,N_23885);
xor U24385 (N_24385,N_23621,N_23950);
nor U24386 (N_24386,N_23635,N_23380);
or U24387 (N_24387,N_23999,N_23546);
nand U24388 (N_24388,N_23065,N_23772);
nand U24389 (N_24389,N_23986,N_23101);
nor U24390 (N_24390,N_22968,N_23235);
and U24391 (N_24391,N_23616,N_23455);
or U24392 (N_24392,N_23392,N_23401);
xor U24393 (N_24393,N_23336,N_22801);
xor U24394 (N_24394,N_23615,N_23254);
and U24395 (N_24395,N_23447,N_22966);
and U24396 (N_24396,N_23868,N_23097);
nor U24397 (N_24397,N_23152,N_23353);
or U24398 (N_24398,N_23902,N_23481);
or U24399 (N_24399,N_23709,N_23925);
nand U24400 (N_24400,N_23213,N_23582);
nor U24401 (N_24401,N_23367,N_23996);
xor U24402 (N_24402,N_23283,N_23703);
or U24403 (N_24403,N_23403,N_23603);
nand U24404 (N_24404,N_23463,N_23686);
or U24405 (N_24405,N_22984,N_22823);
or U24406 (N_24406,N_23911,N_23563);
xor U24407 (N_24407,N_23296,N_23497);
xor U24408 (N_24408,N_23103,N_23122);
nor U24409 (N_24409,N_23428,N_22927);
or U24410 (N_24410,N_23985,N_23570);
nor U24411 (N_24411,N_22822,N_23201);
nor U24412 (N_24412,N_23037,N_23504);
and U24413 (N_24413,N_23055,N_23426);
or U24414 (N_24414,N_23159,N_23309);
nor U24415 (N_24415,N_23653,N_23873);
nor U24416 (N_24416,N_23069,N_23347);
nor U24417 (N_24417,N_23674,N_22821);
and U24418 (N_24418,N_22828,N_23964);
and U24419 (N_24419,N_23838,N_23618);
and U24420 (N_24420,N_23311,N_23270);
or U24421 (N_24421,N_23927,N_23975);
nor U24422 (N_24422,N_23700,N_23871);
and U24423 (N_24423,N_23137,N_23161);
xor U24424 (N_24424,N_22891,N_22810);
nand U24425 (N_24425,N_23575,N_23113);
xnor U24426 (N_24426,N_23106,N_22901);
nor U24427 (N_24427,N_23947,N_23062);
xor U24428 (N_24428,N_23436,N_22857);
xor U24429 (N_24429,N_23171,N_23126);
nor U24430 (N_24430,N_22834,N_23454);
nand U24431 (N_24431,N_23601,N_23230);
nand U24432 (N_24432,N_23564,N_23981);
xnor U24433 (N_24433,N_23837,N_22939);
nor U24434 (N_24434,N_23177,N_23217);
xor U24435 (N_24435,N_23314,N_23887);
nor U24436 (N_24436,N_23623,N_23533);
and U24437 (N_24437,N_22969,N_23798);
or U24438 (N_24438,N_23578,N_23366);
or U24439 (N_24439,N_23063,N_23675);
or U24440 (N_24440,N_23761,N_23776);
nor U24441 (N_24441,N_22800,N_23459);
nor U24442 (N_24442,N_23912,N_23278);
nand U24443 (N_24443,N_23857,N_23108);
and U24444 (N_24444,N_23060,N_23007);
and U24445 (N_24445,N_23886,N_23134);
nand U24446 (N_24446,N_23342,N_23180);
nor U24447 (N_24447,N_23678,N_23717);
nor U24448 (N_24448,N_23852,N_23721);
and U24449 (N_24449,N_23006,N_23644);
xnor U24450 (N_24450,N_23683,N_23193);
xor U24451 (N_24451,N_23212,N_23119);
nand U24452 (N_24452,N_22843,N_23547);
and U24453 (N_24453,N_23086,N_23264);
or U24454 (N_24454,N_23916,N_23340);
or U24455 (N_24455,N_23957,N_23284);
nor U24456 (N_24456,N_23427,N_22954);
and U24457 (N_24457,N_23280,N_23915);
and U24458 (N_24458,N_23279,N_23515);
xor U24459 (N_24459,N_23158,N_23867);
nand U24460 (N_24460,N_23940,N_22945);
nand U24461 (N_24461,N_22848,N_23926);
or U24462 (N_24462,N_23936,N_23745);
or U24463 (N_24463,N_23449,N_23482);
and U24464 (N_24464,N_23096,N_23842);
and U24465 (N_24465,N_23323,N_23977);
xor U24466 (N_24466,N_22832,N_23828);
nor U24467 (N_24467,N_23475,N_23718);
and U24468 (N_24468,N_23954,N_23770);
and U24469 (N_24469,N_23850,N_23317);
xnor U24470 (N_24470,N_23014,N_23009);
nor U24471 (N_24471,N_23269,N_23277);
nor U24472 (N_24472,N_23983,N_23011);
or U24473 (N_24473,N_22884,N_23215);
xor U24474 (N_24474,N_23360,N_23186);
and U24475 (N_24475,N_23728,N_22885);
or U24476 (N_24476,N_23580,N_23469);
nor U24477 (N_24477,N_23540,N_22819);
xor U24478 (N_24478,N_22845,N_23491);
and U24479 (N_24479,N_23240,N_22861);
or U24480 (N_24480,N_23586,N_23572);
nor U24481 (N_24481,N_23499,N_23864);
and U24482 (N_24482,N_23143,N_23440);
nor U24483 (N_24483,N_23493,N_23397);
or U24484 (N_24484,N_23048,N_23803);
and U24485 (N_24485,N_23477,N_23237);
nand U24486 (N_24486,N_22889,N_22813);
nor U24487 (N_24487,N_23960,N_23054);
nand U24488 (N_24488,N_23473,N_23263);
xnor U24489 (N_24489,N_22849,N_23461);
nor U24490 (N_24490,N_23241,N_23759);
xor U24491 (N_24491,N_23079,N_23021);
and U24492 (N_24492,N_23388,N_23165);
nand U24493 (N_24493,N_23518,N_23238);
and U24494 (N_24494,N_22827,N_23974);
xor U24495 (N_24495,N_23033,N_23863);
nand U24496 (N_24496,N_23609,N_23443);
xor U24497 (N_24497,N_23787,N_23501);
and U24498 (N_24498,N_23733,N_23357);
or U24499 (N_24499,N_23075,N_23893);
xor U24500 (N_24500,N_23130,N_23815);
nand U24501 (N_24501,N_23294,N_23064);
nand U24502 (N_24502,N_23072,N_23917);
nand U24503 (N_24503,N_22983,N_23120);
xor U24504 (N_24504,N_23818,N_23719);
xnor U24505 (N_24505,N_23039,N_22989);
nand U24506 (N_24506,N_23846,N_22972);
xnor U24507 (N_24507,N_23920,N_22851);
xor U24508 (N_24508,N_23584,N_23510);
nand U24509 (N_24509,N_23757,N_23112);
xnor U24510 (N_24510,N_23760,N_23679);
nor U24511 (N_24511,N_23672,N_23512);
nor U24512 (N_24512,N_23487,N_23946);
nor U24513 (N_24513,N_23400,N_23667);
or U24514 (N_24514,N_23244,N_23081);
nand U24515 (N_24515,N_23599,N_23654);
nor U24516 (N_24516,N_23082,N_23420);
or U24517 (N_24517,N_23258,N_23910);
nand U24518 (N_24518,N_22990,N_23002);
nor U24519 (N_24519,N_23562,N_22950);
and U24520 (N_24520,N_23581,N_23995);
nor U24521 (N_24521,N_23070,N_23476);
and U24522 (N_24522,N_23298,N_22882);
nor U24523 (N_24523,N_23448,N_23619);
nor U24524 (N_24524,N_23446,N_23997);
nor U24525 (N_24525,N_23199,N_23378);
nand U24526 (N_24526,N_22988,N_23750);
and U24527 (N_24527,N_23694,N_23345);
and U24528 (N_24528,N_23371,N_23231);
nor U24529 (N_24529,N_23368,N_23806);
and U24530 (N_24530,N_23460,N_23969);
nor U24531 (N_24531,N_23310,N_23466);
or U24532 (N_24532,N_22913,N_23164);
xor U24533 (N_24533,N_22815,N_22953);
nor U24534 (N_24534,N_23585,N_23155);
or U24535 (N_24535,N_22897,N_22817);
and U24536 (N_24536,N_23851,N_23265);
nor U24537 (N_24537,N_22831,N_22837);
xor U24538 (N_24538,N_23417,N_23848);
nor U24539 (N_24539,N_23822,N_23358);
or U24540 (N_24540,N_23638,N_23617);
and U24541 (N_24541,N_23839,N_23511);
xnor U24542 (N_24542,N_23929,N_23823);
xor U24543 (N_24543,N_23209,N_23637);
nor U24544 (N_24544,N_23805,N_23710);
and U24545 (N_24545,N_23457,N_23486);
or U24546 (N_24546,N_23275,N_23008);
or U24547 (N_24547,N_22852,N_23539);
xnor U24548 (N_24548,N_23290,N_23399);
and U24549 (N_24549,N_23684,N_23962);
nor U24550 (N_24550,N_22963,N_23588);
nand U24551 (N_24551,N_23285,N_23253);
nor U24552 (N_24552,N_23934,N_23555);
xor U24553 (N_24553,N_23044,N_23085);
nor U24554 (N_24554,N_23896,N_23523);
xnor U24555 (N_24555,N_22922,N_23711);
xor U24556 (N_24556,N_23797,N_22890);
nor U24557 (N_24557,N_23434,N_23138);
nand U24558 (N_24558,N_23170,N_23160);
nand U24559 (N_24559,N_23630,N_22873);
xor U24560 (N_24560,N_23478,N_22928);
xnor U24561 (N_24561,N_23645,N_23029);
xor U24562 (N_24562,N_23556,N_23557);
nand U24563 (N_24563,N_23807,N_23979);
nand U24564 (N_24564,N_23111,N_23775);
xor U24565 (N_24565,N_23696,N_22818);
nor U24566 (N_24566,N_22871,N_23702);
and U24567 (N_24567,N_22959,N_23089);
xnor U24568 (N_24568,N_23869,N_22979);
xor U24569 (N_24569,N_23514,N_23046);
nand U24570 (N_24570,N_22987,N_22853);
nor U24571 (N_24571,N_23668,N_23334);
and U24572 (N_24572,N_23026,N_23726);
nand U24573 (N_24573,N_23965,N_23131);
xor U24574 (N_24574,N_23833,N_22869);
and U24575 (N_24575,N_23377,N_23988);
or U24576 (N_24576,N_23825,N_23548);
and U24577 (N_24577,N_22841,N_23359);
nor U24578 (N_24578,N_23094,N_23980);
nor U24579 (N_24579,N_23151,N_23080);
xor U24580 (N_24580,N_23320,N_23374);
or U24581 (N_24581,N_23831,N_23030);
and U24582 (N_24582,N_23894,N_23875);
nor U24583 (N_24583,N_23057,N_22855);
nand U24584 (N_24584,N_23043,N_23312);
and U24585 (N_24585,N_23441,N_23856);
or U24586 (N_24586,N_23984,N_23904);
xnor U24587 (N_24587,N_23332,N_23502);
nor U24588 (N_24588,N_23519,N_23880);
nor U24589 (N_24589,N_22898,N_22878);
nor U24590 (N_24590,N_23627,N_22868);
nand U24591 (N_24591,N_23970,N_22910);
nand U24592 (N_24592,N_23396,N_23840);
and U24593 (N_24593,N_23306,N_23398);
xnor U24594 (N_24594,N_22826,N_23474);
xor U24595 (N_24595,N_23878,N_22981);
nor U24596 (N_24596,N_22867,N_22980);
or U24597 (N_24597,N_23503,N_23423);
and U24598 (N_24598,N_23110,N_23363);
or U24599 (N_24599,N_23410,N_22879);
nor U24600 (N_24600,N_23066,N_23172);
nor U24601 (N_24601,N_23060,N_23159);
and U24602 (N_24602,N_23598,N_23060);
nand U24603 (N_24603,N_22982,N_23082);
nand U24604 (N_24604,N_23368,N_23381);
xnor U24605 (N_24605,N_23670,N_23331);
nand U24606 (N_24606,N_23318,N_23569);
nor U24607 (N_24607,N_23233,N_23151);
nand U24608 (N_24608,N_23216,N_23622);
or U24609 (N_24609,N_23785,N_22830);
and U24610 (N_24610,N_22987,N_23703);
or U24611 (N_24611,N_23329,N_23410);
nor U24612 (N_24612,N_23853,N_23316);
xor U24613 (N_24613,N_23182,N_23307);
or U24614 (N_24614,N_23591,N_23240);
or U24615 (N_24615,N_22856,N_23473);
xor U24616 (N_24616,N_23310,N_23607);
xnor U24617 (N_24617,N_23560,N_22907);
xnor U24618 (N_24618,N_23274,N_23561);
and U24619 (N_24619,N_23574,N_23000);
and U24620 (N_24620,N_23057,N_23507);
and U24621 (N_24621,N_23703,N_23178);
and U24622 (N_24622,N_22813,N_23757);
and U24623 (N_24623,N_23666,N_23211);
or U24624 (N_24624,N_23030,N_23754);
xor U24625 (N_24625,N_23105,N_23994);
nand U24626 (N_24626,N_23564,N_23468);
nand U24627 (N_24627,N_23672,N_22944);
xnor U24628 (N_24628,N_23082,N_23660);
or U24629 (N_24629,N_22954,N_22870);
nor U24630 (N_24630,N_23333,N_23427);
and U24631 (N_24631,N_23360,N_23855);
and U24632 (N_24632,N_23337,N_22863);
nor U24633 (N_24633,N_23149,N_23326);
nor U24634 (N_24634,N_23878,N_23480);
and U24635 (N_24635,N_23683,N_23673);
or U24636 (N_24636,N_23703,N_23177);
or U24637 (N_24637,N_23909,N_23694);
xor U24638 (N_24638,N_23212,N_22872);
and U24639 (N_24639,N_23935,N_23405);
xor U24640 (N_24640,N_23610,N_23237);
and U24641 (N_24641,N_23611,N_23262);
nor U24642 (N_24642,N_23213,N_23987);
and U24643 (N_24643,N_23708,N_23173);
nand U24644 (N_24644,N_22942,N_23199);
and U24645 (N_24645,N_23260,N_23548);
and U24646 (N_24646,N_23385,N_23420);
and U24647 (N_24647,N_23571,N_23243);
and U24648 (N_24648,N_23441,N_23954);
nand U24649 (N_24649,N_23161,N_23090);
and U24650 (N_24650,N_23498,N_23825);
and U24651 (N_24651,N_22989,N_23947);
nand U24652 (N_24652,N_23474,N_23156);
and U24653 (N_24653,N_23343,N_23761);
xnor U24654 (N_24654,N_23409,N_23552);
nand U24655 (N_24655,N_23961,N_22874);
or U24656 (N_24656,N_23625,N_23374);
and U24657 (N_24657,N_23247,N_23616);
and U24658 (N_24658,N_23594,N_23167);
and U24659 (N_24659,N_23888,N_22984);
nor U24660 (N_24660,N_22829,N_23136);
and U24661 (N_24661,N_22833,N_22844);
or U24662 (N_24662,N_22845,N_23458);
and U24663 (N_24663,N_23042,N_22896);
or U24664 (N_24664,N_23799,N_22803);
and U24665 (N_24665,N_23001,N_23851);
nor U24666 (N_24666,N_23223,N_23532);
nand U24667 (N_24667,N_22956,N_23040);
nand U24668 (N_24668,N_23449,N_23689);
or U24669 (N_24669,N_23704,N_23249);
or U24670 (N_24670,N_23342,N_23754);
nor U24671 (N_24671,N_22967,N_23903);
and U24672 (N_24672,N_23770,N_22919);
or U24673 (N_24673,N_23342,N_22847);
nor U24674 (N_24674,N_23726,N_23062);
xor U24675 (N_24675,N_23549,N_23640);
xnor U24676 (N_24676,N_23504,N_23613);
nor U24677 (N_24677,N_23279,N_23817);
xnor U24678 (N_24678,N_23105,N_23828);
and U24679 (N_24679,N_23675,N_23140);
nor U24680 (N_24680,N_23129,N_23576);
nor U24681 (N_24681,N_23699,N_23718);
xnor U24682 (N_24682,N_23501,N_23863);
nand U24683 (N_24683,N_23098,N_22877);
nor U24684 (N_24684,N_23026,N_22901);
nand U24685 (N_24685,N_23838,N_23685);
and U24686 (N_24686,N_23581,N_23141);
nor U24687 (N_24687,N_23288,N_23666);
xor U24688 (N_24688,N_23294,N_23991);
xor U24689 (N_24689,N_23492,N_23560);
or U24690 (N_24690,N_23082,N_23481);
xor U24691 (N_24691,N_23013,N_23704);
nor U24692 (N_24692,N_23244,N_23052);
nand U24693 (N_24693,N_23709,N_23216);
or U24694 (N_24694,N_22952,N_23184);
or U24695 (N_24695,N_23046,N_23293);
nand U24696 (N_24696,N_22806,N_22960);
nor U24697 (N_24697,N_23998,N_23501);
or U24698 (N_24698,N_23382,N_22931);
nand U24699 (N_24699,N_23111,N_23828);
and U24700 (N_24700,N_23395,N_23475);
nand U24701 (N_24701,N_23064,N_22864);
and U24702 (N_24702,N_23301,N_22982);
nor U24703 (N_24703,N_23036,N_22984);
or U24704 (N_24704,N_23627,N_23664);
nand U24705 (N_24705,N_23859,N_23372);
nor U24706 (N_24706,N_22834,N_23092);
nor U24707 (N_24707,N_23406,N_23576);
or U24708 (N_24708,N_23151,N_23411);
or U24709 (N_24709,N_22972,N_23643);
nand U24710 (N_24710,N_23557,N_23129);
and U24711 (N_24711,N_23409,N_23807);
nor U24712 (N_24712,N_22843,N_23320);
nand U24713 (N_24713,N_23449,N_22892);
nor U24714 (N_24714,N_22984,N_23711);
xor U24715 (N_24715,N_22804,N_23197);
xnor U24716 (N_24716,N_23260,N_23442);
nor U24717 (N_24717,N_23038,N_23405);
xor U24718 (N_24718,N_22946,N_23028);
and U24719 (N_24719,N_23363,N_23911);
nor U24720 (N_24720,N_23145,N_23492);
xnor U24721 (N_24721,N_23727,N_23359);
nor U24722 (N_24722,N_23632,N_23756);
and U24723 (N_24723,N_22812,N_23462);
xnor U24724 (N_24724,N_23408,N_23434);
xnor U24725 (N_24725,N_23832,N_23384);
xor U24726 (N_24726,N_23804,N_23995);
xnor U24727 (N_24727,N_23577,N_22884);
xnor U24728 (N_24728,N_23074,N_23000);
xnor U24729 (N_24729,N_23819,N_23283);
nand U24730 (N_24730,N_23269,N_22955);
and U24731 (N_24731,N_23529,N_23330);
nand U24732 (N_24732,N_23820,N_23248);
nand U24733 (N_24733,N_23133,N_22838);
and U24734 (N_24734,N_23085,N_23501);
or U24735 (N_24735,N_23929,N_23192);
xor U24736 (N_24736,N_23836,N_23264);
nor U24737 (N_24737,N_23578,N_23523);
or U24738 (N_24738,N_23188,N_23631);
and U24739 (N_24739,N_23965,N_23002);
and U24740 (N_24740,N_23882,N_23923);
nor U24741 (N_24741,N_23923,N_23772);
and U24742 (N_24742,N_23413,N_23613);
or U24743 (N_24743,N_23268,N_23869);
xor U24744 (N_24744,N_23135,N_22964);
or U24745 (N_24745,N_22850,N_23707);
nand U24746 (N_24746,N_22832,N_23561);
or U24747 (N_24747,N_23493,N_23519);
nand U24748 (N_24748,N_22872,N_22863);
and U24749 (N_24749,N_23438,N_22818);
and U24750 (N_24750,N_22824,N_23539);
nor U24751 (N_24751,N_23917,N_22816);
nand U24752 (N_24752,N_23128,N_23924);
or U24753 (N_24753,N_22877,N_23424);
xnor U24754 (N_24754,N_23975,N_23089);
or U24755 (N_24755,N_22828,N_23838);
nand U24756 (N_24756,N_23462,N_23640);
or U24757 (N_24757,N_23796,N_23854);
xnor U24758 (N_24758,N_23282,N_23671);
nor U24759 (N_24759,N_23898,N_22892);
xnor U24760 (N_24760,N_22812,N_22809);
nor U24761 (N_24761,N_23652,N_23584);
and U24762 (N_24762,N_23801,N_23042);
xor U24763 (N_24763,N_23383,N_23195);
nand U24764 (N_24764,N_23099,N_23933);
xor U24765 (N_24765,N_23086,N_23224);
or U24766 (N_24766,N_22925,N_23563);
or U24767 (N_24767,N_22878,N_23850);
and U24768 (N_24768,N_22897,N_23328);
nand U24769 (N_24769,N_23823,N_23147);
nor U24770 (N_24770,N_23706,N_23570);
or U24771 (N_24771,N_23743,N_23255);
nand U24772 (N_24772,N_22891,N_22873);
xor U24773 (N_24773,N_22854,N_23733);
or U24774 (N_24774,N_22990,N_23992);
xor U24775 (N_24775,N_23474,N_23339);
nand U24776 (N_24776,N_23680,N_22923);
nand U24777 (N_24777,N_23703,N_23896);
nand U24778 (N_24778,N_23546,N_23720);
nand U24779 (N_24779,N_23572,N_23396);
nor U24780 (N_24780,N_23755,N_23560);
or U24781 (N_24781,N_23716,N_23282);
xnor U24782 (N_24782,N_23685,N_23761);
and U24783 (N_24783,N_23186,N_23393);
nand U24784 (N_24784,N_23368,N_23463);
and U24785 (N_24785,N_23169,N_23742);
nand U24786 (N_24786,N_23770,N_23861);
nor U24787 (N_24787,N_23244,N_23798);
or U24788 (N_24788,N_23192,N_23620);
or U24789 (N_24789,N_23825,N_22880);
and U24790 (N_24790,N_23806,N_23525);
xor U24791 (N_24791,N_23909,N_22850);
xor U24792 (N_24792,N_23745,N_23353);
xnor U24793 (N_24793,N_23616,N_22802);
or U24794 (N_24794,N_23052,N_23042);
nor U24795 (N_24795,N_23540,N_23189);
nand U24796 (N_24796,N_23122,N_22830);
nor U24797 (N_24797,N_23428,N_22887);
and U24798 (N_24798,N_23217,N_23653);
xor U24799 (N_24799,N_23274,N_22971);
nor U24800 (N_24800,N_23196,N_23271);
nor U24801 (N_24801,N_23472,N_23479);
and U24802 (N_24802,N_23426,N_22920);
and U24803 (N_24803,N_23672,N_23674);
or U24804 (N_24804,N_23602,N_23078);
or U24805 (N_24805,N_23258,N_22936);
xnor U24806 (N_24806,N_23289,N_23579);
xor U24807 (N_24807,N_23103,N_22966);
and U24808 (N_24808,N_23488,N_23698);
and U24809 (N_24809,N_22915,N_23917);
and U24810 (N_24810,N_23987,N_23026);
nand U24811 (N_24811,N_23304,N_23542);
nor U24812 (N_24812,N_23565,N_23591);
nor U24813 (N_24813,N_23571,N_22847);
xor U24814 (N_24814,N_22851,N_23717);
xnor U24815 (N_24815,N_23588,N_23913);
and U24816 (N_24816,N_22913,N_22956);
nor U24817 (N_24817,N_23878,N_23668);
nor U24818 (N_24818,N_23580,N_23963);
nand U24819 (N_24819,N_23967,N_23496);
or U24820 (N_24820,N_23506,N_23966);
xor U24821 (N_24821,N_23237,N_23649);
and U24822 (N_24822,N_23327,N_23047);
nor U24823 (N_24823,N_23661,N_23982);
nor U24824 (N_24824,N_23230,N_23909);
xor U24825 (N_24825,N_23530,N_22863);
and U24826 (N_24826,N_23573,N_22898);
and U24827 (N_24827,N_23134,N_23267);
nand U24828 (N_24828,N_23560,N_23086);
xnor U24829 (N_24829,N_23226,N_23775);
nor U24830 (N_24830,N_22806,N_23687);
or U24831 (N_24831,N_23446,N_22995);
and U24832 (N_24832,N_23527,N_23835);
xor U24833 (N_24833,N_23522,N_23118);
and U24834 (N_24834,N_23029,N_22983);
or U24835 (N_24835,N_22901,N_23884);
and U24836 (N_24836,N_23982,N_23857);
nand U24837 (N_24837,N_23254,N_23945);
or U24838 (N_24838,N_23568,N_22853);
xnor U24839 (N_24839,N_23651,N_23380);
and U24840 (N_24840,N_23473,N_23842);
xor U24841 (N_24841,N_23208,N_23245);
nor U24842 (N_24842,N_23447,N_23685);
xor U24843 (N_24843,N_23053,N_23670);
or U24844 (N_24844,N_23143,N_23756);
and U24845 (N_24845,N_23663,N_23326);
nor U24846 (N_24846,N_22858,N_23321);
and U24847 (N_24847,N_23291,N_23028);
and U24848 (N_24848,N_23320,N_23618);
or U24849 (N_24849,N_22926,N_23487);
xnor U24850 (N_24850,N_23262,N_23141);
nor U24851 (N_24851,N_23100,N_23886);
nand U24852 (N_24852,N_22830,N_22938);
or U24853 (N_24853,N_23799,N_23163);
or U24854 (N_24854,N_23694,N_23786);
and U24855 (N_24855,N_23670,N_23123);
or U24856 (N_24856,N_23057,N_23989);
nor U24857 (N_24857,N_23751,N_23230);
nor U24858 (N_24858,N_23301,N_22889);
nand U24859 (N_24859,N_23746,N_22902);
nor U24860 (N_24860,N_22951,N_23465);
or U24861 (N_24861,N_23442,N_23084);
nor U24862 (N_24862,N_23603,N_23640);
xnor U24863 (N_24863,N_23028,N_23334);
or U24864 (N_24864,N_23834,N_23199);
nor U24865 (N_24865,N_23293,N_23248);
xor U24866 (N_24866,N_23362,N_23433);
or U24867 (N_24867,N_23304,N_22817);
and U24868 (N_24868,N_23142,N_23429);
nand U24869 (N_24869,N_23002,N_22839);
nand U24870 (N_24870,N_23953,N_23975);
nand U24871 (N_24871,N_23661,N_23774);
and U24872 (N_24872,N_23713,N_23969);
and U24873 (N_24873,N_23569,N_23028);
nand U24874 (N_24874,N_23024,N_23675);
nor U24875 (N_24875,N_22804,N_23261);
xnor U24876 (N_24876,N_23909,N_22912);
or U24877 (N_24877,N_23544,N_22942);
and U24878 (N_24878,N_23261,N_23583);
nor U24879 (N_24879,N_23937,N_23998);
nand U24880 (N_24880,N_23361,N_23632);
nand U24881 (N_24881,N_23836,N_22939);
and U24882 (N_24882,N_22998,N_23307);
nand U24883 (N_24883,N_23688,N_23433);
or U24884 (N_24884,N_23440,N_23257);
or U24885 (N_24885,N_23581,N_22944);
and U24886 (N_24886,N_23556,N_23402);
nor U24887 (N_24887,N_23567,N_22891);
or U24888 (N_24888,N_23973,N_23681);
and U24889 (N_24889,N_23646,N_23352);
nand U24890 (N_24890,N_23408,N_23973);
xnor U24891 (N_24891,N_23649,N_22833);
xnor U24892 (N_24892,N_23217,N_23070);
xnor U24893 (N_24893,N_23060,N_23155);
nand U24894 (N_24894,N_23570,N_23024);
and U24895 (N_24895,N_23387,N_23952);
and U24896 (N_24896,N_22983,N_22842);
xor U24897 (N_24897,N_23223,N_23796);
nor U24898 (N_24898,N_23976,N_23407);
or U24899 (N_24899,N_22861,N_23466);
or U24900 (N_24900,N_22927,N_23338);
and U24901 (N_24901,N_23905,N_22979);
and U24902 (N_24902,N_23027,N_23196);
or U24903 (N_24903,N_23874,N_23350);
or U24904 (N_24904,N_23820,N_23591);
nand U24905 (N_24905,N_23465,N_23081);
and U24906 (N_24906,N_23368,N_22913);
nand U24907 (N_24907,N_23591,N_23070);
and U24908 (N_24908,N_22909,N_23998);
xnor U24909 (N_24909,N_23495,N_23544);
or U24910 (N_24910,N_23573,N_23899);
nor U24911 (N_24911,N_23098,N_23028);
xor U24912 (N_24912,N_23932,N_23616);
or U24913 (N_24913,N_23916,N_23472);
or U24914 (N_24914,N_23972,N_23926);
xor U24915 (N_24915,N_23278,N_23029);
xor U24916 (N_24916,N_23792,N_23796);
or U24917 (N_24917,N_22858,N_23505);
or U24918 (N_24918,N_23863,N_22803);
and U24919 (N_24919,N_23378,N_23669);
nor U24920 (N_24920,N_23536,N_23040);
xor U24921 (N_24921,N_23719,N_23542);
or U24922 (N_24922,N_23610,N_22826);
xor U24923 (N_24923,N_23661,N_23262);
xnor U24924 (N_24924,N_23871,N_23959);
nor U24925 (N_24925,N_23673,N_23607);
or U24926 (N_24926,N_23608,N_23522);
and U24927 (N_24927,N_23723,N_23366);
xor U24928 (N_24928,N_23078,N_23633);
nor U24929 (N_24929,N_23145,N_22855);
and U24930 (N_24930,N_23017,N_23216);
and U24931 (N_24931,N_23138,N_23690);
xnor U24932 (N_24932,N_23542,N_23802);
nor U24933 (N_24933,N_23643,N_22843);
and U24934 (N_24934,N_23414,N_23843);
nor U24935 (N_24935,N_23124,N_23493);
or U24936 (N_24936,N_23992,N_23256);
xnor U24937 (N_24937,N_23725,N_22861);
nor U24938 (N_24938,N_23311,N_23038);
and U24939 (N_24939,N_23590,N_23905);
nor U24940 (N_24940,N_22827,N_22993);
nor U24941 (N_24941,N_22856,N_23810);
nor U24942 (N_24942,N_23077,N_23946);
nand U24943 (N_24943,N_23934,N_23718);
xnor U24944 (N_24944,N_23729,N_23287);
xor U24945 (N_24945,N_23661,N_23288);
nor U24946 (N_24946,N_23670,N_23691);
or U24947 (N_24947,N_23559,N_23708);
xor U24948 (N_24948,N_23550,N_23023);
nor U24949 (N_24949,N_23903,N_23449);
or U24950 (N_24950,N_22864,N_23255);
and U24951 (N_24951,N_23297,N_22908);
and U24952 (N_24952,N_23864,N_23231);
nor U24953 (N_24953,N_23466,N_23990);
xnor U24954 (N_24954,N_23317,N_23692);
or U24955 (N_24955,N_23317,N_23107);
nor U24956 (N_24956,N_22903,N_23488);
xnor U24957 (N_24957,N_23093,N_23583);
nor U24958 (N_24958,N_23484,N_23901);
xnor U24959 (N_24959,N_23230,N_23572);
or U24960 (N_24960,N_22959,N_23831);
xor U24961 (N_24961,N_23717,N_23949);
and U24962 (N_24962,N_23477,N_23894);
and U24963 (N_24963,N_22870,N_23821);
nor U24964 (N_24964,N_23459,N_23105);
xor U24965 (N_24965,N_23793,N_22943);
or U24966 (N_24966,N_23884,N_23856);
nor U24967 (N_24967,N_22933,N_23073);
nand U24968 (N_24968,N_22802,N_23737);
nand U24969 (N_24969,N_23324,N_23152);
or U24970 (N_24970,N_23467,N_23325);
and U24971 (N_24971,N_23401,N_23037);
nor U24972 (N_24972,N_23478,N_23069);
nand U24973 (N_24973,N_23046,N_23472);
nand U24974 (N_24974,N_23663,N_23872);
nand U24975 (N_24975,N_23214,N_22835);
xnor U24976 (N_24976,N_23230,N_23849);
nand U24977 (N_24977,N_23686,N_23731);
or U24978 (N_24978,N_23649,N_23270);
xor U24979 (N_24979,N_23736,N_23647);
nor U24980 (N_24980,N_23317,N_23104);
nand U24981 (N_24981,N_23080,N_23960);
nor U24982 (N_24982,N_23753,N_23944);
xor U24983 (N_24983,N_23950,N_23622);
nand U24984 (N_24984,N_23299,N_22990);
or U24985 (N_24985,N_23355,N_23925);
nand U24986 (N_24986,N_23692,N_23084);
or U24987 (N_24987,N_23178,N_23441);
and U24988 (N_24988,N_23768,N_23468);
or U24989 (N_24989,N_23637,N_22920);
xor U24990 (N_24990,N_23609,N_23391);
nor U24991 (N_24991,N_23301,N_23529);
or U24992 (N_24992,N_23366,N_23973);
and U24993 (N_24993,N_23650,N_23812);
and U24994 (N_24994,N_23441,N_23047);
or U24995 (N_24995,N_22828,N_23588);
xnor U24996 (N_24996,N_23934,N_22979);
nor U24997 (N_24997,N_23336,N_22999);
and U24998 (N_24998,N_23819,N_23738);
or U24999 (N_24999,N_23496,N_23551);
nand U25000 (N_25000,N_22895,N_22875);
nor U25001 (N_25001,N_23438,N_22832);
or U25002 (N_25002,N_22901,N_23626);
nand U25003 (N_25003,N_22809,N_23875);
nor U25004 (N_25004,N_23006,N_23994);
nor U25005 (N_25005,N_23354,N_23000);
xnor U25006 (N_25006,N_23420,N_23390);
xnor U25007 (N_25007,N_23378,N_22896);
xnor U25008 (N_25008,N_23589,N_23390);
xnor U25009 (N_25009,N_23826,N_23271);
nand U25010 (N_25010,N_22817,N_23805);
nor U25011 (N_25011,N_23474,N_23510);
or U25012 (N_25012,N_22805,N_23612);
or U25013 (N_25013,N_23197,N_23005);
nand U25014 (N_25014,N_22829,N_23487);
and U25015 (N_25015,N_23637,N_23217);
nand U25016 (N_25016,N_22961,N_23046);
or U25017 (N_25017,N_23940,N_23830);
and U25018 (N_25018,N_23227,N_23841);
nand U25019 (N_25019,N_23007,N_22933);
and U25020 (N_25020,N_23785,N_22961);
xor U25021 (N_25021,N_23768,N_23676);
nand U25022 (N_25022,N_23143,N_23033);
nor U25023 (N_25023,N_22864,N_23296);
xor U25024 (N_25024,N_23282,N_23737);
and U25025 (N_25025,N_23372,N_23447);
nand U25026 (N_25026,N_23105,N_23872);
nand U25027 (N_25027,N_23423,N_23946);
nor U25028 (N_25028,N_23651,N_23282);
and U25029 (N_25029,N_23569,N_23936);
and U25030 (N_25030,N_23855,N_23999);
xor U25031 (N_25031,N_23120,N_23505);
nand U25032 (N_25032,N_23987,N_23019);
nand U25033 (N_25033,N_23661,N_23449);
and U25034 (N_25034,N_23151,N_22815);
nor U25035 (N_25035,N_23664,N_22908);
xnor U25036 (N_25036,N_23836,N_23160);
xnor U25037 (N_25037,N_23776,N_23295);
nand U25038 (N_25038,N_23272,N_23560);
nor U25039 (N_25039,N_22912,N_23463);
xnor U25040 (N_25040,N_23725,N_22997);
xor U25041 (N_25041,N_23829,N_23146);
xor U25042 (N_25042,N_23888,N_23382);
xor U25043 (N_25043,N_23293,N_23186);
xor U25044 (N_25044,N_23823,N_23927);
xnor U25045 (N_25045,N_23294,N_22848);
xor U25046 (N_25046,N_23483,N_22980);
nand U25047 (N_25047,N_22814,N_23605);
nand U25048 (N_25048,N_22868,N_23097);
xnor U25049 (N_25049,N_23931,N_23336);
xor U25050 (N_25050,N_23156,N_23106);
and U25051 (N_25051,N_23075,N_23514);
and U25052 (N_25052,N_23500,N_23597);
or U25053 (N_25053,N_23096,N_23338);
and U25054 (N_25054,N_23064,N_23623);
nand U25055 (N_25055,N_23039,N_22884);
and U25056 (N_25056,N_23111,N_23175);
and U25057 (N_25057,N_23545,N_23790);
or U25058 (N_25058,N_22971,N_23173);
nor U25059 (N_25059,N_23354,N_23123);
xnor U25060 (N_25060,N_23431,N_23605);
and U25061 (N_25061,N_23808,N_23781);
nor U25062 (N_25062,N_23626,N_23404);
or U25063 (N_25063,N_23472,N_23281);
nand U25064 (N_25064,N_23163,N_23244);
and U25065 (N_25065,N_23329,N_23516);
nor U25066 (N_25066,N_23565,N_22993);
nor U25067 (N_25067,N_23268,N_23827);
xor U25068 (N_25068,N_23054,N_23706);
and U25069 (N_25069,N_22801,N_23517);
nand U25070 (N_25070,N_23386,N_23107);
or U25071 (N_25071,N_22852,N_23873);
and U25072 (N_25072,N_22997,N_23898);
and U25073 (N_25073,N_23495,N_23587);
nor U25074 (N_25074,N_22814,N_23940);
nor U25075 (N_25075,N_23748,N_22860);
nor U25076 (N_25076,N_23081,N_23748);
or U25077 (N_25077,N_23779,N_23766);
or U25078 (N_25078,N_23249,N_23499);
nand U25079 (N_25079,N_23940,N_23368);
and U25080 (N_25080,N_23842,N_23777);
or U25081 (N_25081,N_23759,N_23533);
and U25082 (N_25082,N_23085,N_23311);
nand U25083 (N_25083,N_23032,N_23523);
nand U25084 (N_25084,N_23723,N_23345);
nor U25085 (N_25085,N_22900,N_23783);
and U25086 (N_25086,N_22898,N_23346);
and U25087 (N_25087,N_22960,N_23930);
or U25088 (N_25088,N_23709,N_23783);
or U25089 (N_25089,N_23514,N_23685);
and U25090 (N_25090,N_23318,N_23791);
or U25091 (N_25091,N_23321,N_23056);
xnor U25092 (N_25092,N_23006,N_23649);
and U25093 (N_25093,N_23484,N_22988);
xor U25094 (N_25094,N_22982,N_23776);
nand U25095 (N_25095,N_23906,N_23718);
or U25096 (N_25096,N_22916,N_23201);
or U25097 (N_25097,N_23107,N_22930);
or U25098 (N_25098,N_23140,N_23458);
or U25099 (N_25099,N_23600,N_23699);
and U25100 (N_25100,N_22868,N_22958);
and U25101 (N_25101,N_23744,N_23806);
or U25102 (N_25102,N_22868,N_23692);
or U25103 (N_25103,N_22952,N_23749);
nand U25104 (N_25104,N_23768,N_23379);
and U25105 (N_25105,N_22906,N_23834);
xor U25106 (N_25106,N_23633,N_23207);
or U25107 (N_25107,N_23371,N_22921);
nor U25108 (N_25108,N_23426,N_23765);
nor U25109 (N_25109,N_23934,N_23974);
nand U25110 (N_25110,N_23296,N_22822);
nand U25111 (N_25111,N_23545,N_23945);
or U25112 (N_25112,N_23968,N_23196);
or U25113 (N_25113,N_23253,N_23773);
or U25114 (N_25114,N_23381,N_23412);
or U25115 (N_25115,N_23645,N_23713);
nand U25116 (N_25116,N_23404,N_22869);
or U25117 (N_25117,N_22844,N_23052);
or U25118 (N_25118,N_23613,N_22947);
nor U25119 (N_25119,N_23400,N_23005);
and U25120 (N_25120,N_22898,N_23215);
or U25121 (N_25121,N_23570,N_23701);
xnor U25122 (N_25122,N_23579,N_23809);
and U25123 (N_25123,N_23118,N_23944);
nand U25124 (N_25124,N_23134,N_23212);
xnor U25125 (N_25125,N_23812,N_22891);
nand U25126 (N_25126,N_22962,N_23319);
and U25127 (N_25127,N_23133,N_23524);
xor U25128 (N_25128,N_23254,N_23971);
nand U25129 (N_25129,N_22889,N_23584);
nand U25130 (N_25130,N_23783,N_23403);
nand U25131 (N_25131,N_23454,N_23144);
nand U25132 (N_25132,N_23978,N_23402);
xnor U25133 (N_25133,N_22897,N_23872);
or U25134 (N_25134,N_23716,N_22907);
nor U25135 (N_25135,N_23797,N_23382);
and U25136 (N_25136,N_23543,N_23556);
xnor U25137 (N_25137,N_22854,N_23688);
xnor U25138 (N_25138,N_22906,N_23013);
nor U25139 (N_25139,N_23272,N_23311);
nor U25140 (N_25140,N_23303,N_23873);
nor U25141 (N_25141,N_22948,N_23580);
xnor U25142 (N_25142,N_22877,N_23521);
and U25143 (N_25143,N_23251,N_23861);
xnor U25144 (N_25144,N_23085,N_23535);
xor U25145 (N_25145,N_23059,N_23474);
xor U25146 (N_25146,N_23253,N_23330);
nor U25147 (N_25147,N_23371,N_23956);
or U25148 (N_25148,N_23661,N_23241);
or U25149 (N_25149,N_23234,N_23396);
nor U25150 (N_25150,N_23290,N_23074);
nand U25151 (N_25151,N_23781,N_23377);
xnor U25152 (N_25152,N_23212,N_23453);
nor U25153 (N_25153,N_23492,N_23747);
xor U25154 (N_25154,N_23242,N_23133);
and U25155 (N_25155,N_23214,N_23126);
xor U25156 (N_25156,N_22828,N_23039);
nor U25157 (N_25157,N_23953,N_23071);
xnor U25158 (N_25158,N_23888,N_23068);
xor U25159 (N_25159,N_22804,N_22967);
or U25160 (N_25160,N_23606,N_22834);
nor U25161 (N_25161,N_23862,N_23088);
xor U25162 (N_25162,N_23486,N_23761);
nand U25163 (N_25163,N_23153,N_23513);
nor U25164 (N_25164,N_22815,N_23251);
nand U25165 (N_25165,N_23648,N_23692);
nand U25166 (N_25166,N_23251,N_23785);
nor U25167 (N_25167,N_23445,N_23752);
and U25168 (N_25168,N_23035,N_22983);
nand U25169 (N_25169,N_23570,N_23573);
nor U25170 (N_25170,N_23710,N_23054);
or U25171 (N_25171,N_23945,N_23970);
nand U25172 (N_25172,N_23891,N_23149);
xnor U25173 (N_25173,N_23605,N_23128);
nand U25174 (N_25174,N_22982,N_23809);
or U25175 (N_25175,N_23264,N_22878);
and U25176 (N_25176,N_23898,N_22990);
nand U25177 (N_25177,N_23160,N_22964);
nand U25178 (N_25178,N_23437,N_23114);
and U25179 (N_25179,N_22954,N_22887);
or U25180 (N_25180,N_22995,N_23652);
nor U25181 (N_25181,N_23603,N_23192);
nand U25182 (N_25182,N_23302,N_23474);
xor U25183 (N_25183,N_23274,N_23441);
and U25184 (N_25184,N_23718,N_22972);
and U25185 (N_25185,N_23242,N_23083);
xor U25186 (N_25186,N_23120,N_23005);
or U25187 (N_25187,N_23739,N_23254);
or U25188 (N_25188,N_22962,N_22858);
nor U25189 (N_25189,N_23946,N_23517);
or U25190 (N_25190,N_23971,N_22861);
nand U25191 (N_25191,N_23886,N_23691);
or U25192 (N_25192,N_22821,N_23941);
and U25193 (N_25193,N_23641,N_23375);
nor U25194 (N_25194,N_23797,N_22932);
nand U25195 (N_25195,N_23206,N_23145);
nand U25196 (N_25196,N_23711,N_23331);
nand U25197 (N_25197,N_23144,N_23937);
nor U25198 (N_25198,N_23175,N_23493);
or U25199 (N_25199,N_22955,N_23396);
or U25200 (N_25200,N_24558,N_24319);
and U25201 (N_25201,N_24867,N_24226);
nand U25202 (N_25202,N_24931,N_24722);
and U25203 (N_25203,N_24087,N_24136);
xor U25204 (N_25204,N_24238,N_24749);
nand U25205 (N_25205,N_25044,N_24107);
xor U25206 (N_25206,N_24383,N_25138);
nor U25207 (N_25207,N_24428,N_24381);
or U25208 (N_25208,N_24316,N_24103);
xor U25209 (N_25209,N_24727,N_24811);
nand U25210 (N_25210,N_24273,N_24862);
and U25211 (N_25211,N_24992,N_24050);
nand U25212 (N_25212,N_24790,N_24349);
nor U25213 (N_25213,N_24212,N_25047);
and U25214 (N_25214,N_25096,N_24698);
or U25215 (N_25215,N_24938,N_24630);
and U25216 (N_25216,N_24803,N_25107);
nor U25217 (N_25217,N_24982,N_24371);
nand U25218 (N_25218,N_24486,N_24051);
nand U25219 (N_25219,N_25065,N_25051);
nor U25220 (N_25220,N_24220,N_24490);
nor U25221 (N_25221,N_24792,N_24951);
xnor U25222 (N_25222,N_24510,N_24824);
and U25223 (N_25223,N_24621,N_25015);
or U25224 (N_25224,N_24866,N_24329);
and U25225 (N_25225,N_24146,N_24755);
or U25226 (N_25226,N_24833,N_24855);
or U25227 (N_25227,N_24148,N_25063);
or U25228 (N_25228,N_24019,N_24828);
xnor U25229 (N_25229,N_24234,N_24441);
xor U25230 (N_25230,N_24820,N_24406);
nand U25231 (N_25231,N_24467,N_25185);
nor U25232 (N_25232,N_24607,N_25112);
xor U25233 (N_25233,N_24491,N_24239);
nand U25234 (N_25234,N_25105,N_24493);
xnor U25235 (N_25235,N_24043,N_25148);
nand U25236 (N_25236,N_24813,N_25177);
nor U25237 (N_25237,N_24993,N_24771);
nor U25238 (N_25238,N_25070,N_25145);
xnor U25239 (N_25239,N_24795,N_25073);
or U25240 (N_25240,N_24044,N_24396);
nor U25241 (N_25241,N_24819,N_25032);
nand U25242 (N_25242,N_24070,N_24458);
and U25243 (N_25243,N_24508,N_24207);
nand U25244 (N_25244,N_24169,N_24487);
or U25245 (N_25245,N_25199,N_24586);
and U25246 (N_25246,N_24193,N_24845);
and U25247 (N_25247,N_24142,N_24957);
and U25248 (N_25248,N_24304,N_25193);
xor U25249 (N_25249,N_24906,N_25014);
nor U25250 (N_25250,N_24449,N_24633);
nor U25251 (N_25251,N_24699,N_24466);
nand U25252 (N_25252,N_25027,N_24187);
nor U25253 (N_25253,N_24286,N_25017);
nand U25254 (N_25254,N_24900,N_24553);
nor U25255 (N_25255,N_25159,N_24414);
and U25256 (N_25256,N_24001,N_24147);
nand U25257 (N_25257,N_24770,N_24579);
xor U25258 (N_25258,N_24397,N_24981);
nand U25259 (N_25259,N_24005,N_24988);
nand U25260 (N_25260,N_24036,N_24884);
nand U25261 (N_25261,N_25154,N_24965);
or U25262 (N_25262,N_24057,N_24445);
nor U25263 (N_25263,N_24126,N_24111);
nor U25264 (N_25264,N_24378,N_24963);
or U25265 (N_25265,N_24958,N_24846);
xor U25266 (N_25266,N_24604,N_24509);
or U25267 (N_25267,N_24806,N_24578);
and U25268 (N_25268,N_24264,N_25198);
nor U25269 (N_25269,N_24455,N_24045);
xnor U25270 (N_25270,N_25092,N_24011);
nand U25271 (N_25271,N_24496,N_24893);
nor U25272 (N_25272,N_24452,N_24394);
nand U25273 (N_25273,N_24164,N_24878);
nand U25274 (N_25274,N_24966,N_24088);
or U25275 (N_25275,N_24544,N_24268);
or U25276 (N_25276,N_24315,N_25166);
nand U25277 (N_25277,N_24980,N_24106);
nand U25278 (N_25278,N_25192,N_24214);
or U25279 (N_25279,N_25039,N_24099);
nand U25280 (N_25280,N_25187,N_24233);
and U25281 (N_25281,N_24040,N_24404);
nand U25282 (N_25282,N_24355,N_24461);
or U25283 (N_25283,N_24912,N_25064);
and U25284 (N_25284,N_25012,N_24017);
nand U25285 (N_25285,N_24280,N_24779);
or U25286 (N_25286,N_24200,N_24506);
or U25287 (N_25287,N_24376,N_24556);
xnor U25288 (N_25288,N_24521,N_25061);
and U25289 (N_25289,N_24703,N_24113);
xor U25290 (N_25290,N_24868,N_25147);
nand U25291 (N_25291,N_24129,N_24520);
or U25292 (N_25292,N_24185,N_24390);
nor U25293 (N_25293,N_24027,N_24047);
and U25294 (N_25294,N_24503,N_24822);
or U25295 (N_25295,N_24116,N_24014);
nand U25296 (N_25296,N_24525,N_24393);
nand U25297 (N_25297,N_24901,N_24231);
or U25298 (N_25298,N_24171,N_25010);
nand U25299 (N_25299,N_24384,N_24844);
xor U25300 (N_25300,N_24317,N_24661);
nor U25301 (N_25301,N_24863,N_24530);
nor U25302 (N_25302,N_24569,N_24538);
xor U25303 (N_25303,N_24737,N_24590);
and U25304 (N_25304,N_24004,N_24723);
nor U25305 (N_25305,N_24624,N_24483);
nor U25306 (N_25306,N_24724,N_25068);
nand U25307 (N_25307,N_24972,N_24697);
or U25308 (N_25308,N_25006,N_24096);
nand U25309 (N_25309,N_24746,N_24761);
and U25310 (N_25310,N_25158,N_24130);
and U25311 (N_25311,N_24913,N_24476);
and U25312 (N_25312,N_24548,N_24440);
nor U25313 (N_25313,N_25135,N_24612);
or U25314 (N_25314,N_24533,N_24944);
nand U25315 (N_25315,N_24758,N_24137);
nand U25316 (N_25316,N_24772,N_25018);
nor U25317 (N_25317,N_25082,N_24998);
xnor U25318 (N_25318,N_24481,N_24660);
and U25319 (N_25319,N_24252,N_25060);
nand U25320 (N_25320,N_24805,N_25028);
and U25321 (N_25321,N_24898,N_24917);
and U25322 (N_25322,N_25109,N_24567);
nor U25323 (N_25323,N_25155,N_24768);
nand U25324 (N_25324,N_24265,N_24872);
xnor U25325 (N_25325,N_25183,N_24856);
or U25326 (N_25326,N_25072,N_24289);
and U25327 (N_25327,N_24780,N_24583);
xnor U25328 (N_25328,N_24743,N_24323);
nand U25329 (N_25329,N_24996,N_24092);
and U25330 (N_25330,N_24402,N_24584);
xor U25331 (N_25331,N_24350,N_24653);
xor U25332 (N_25332,N_25176,N_24124);
nand U25333 (N_25333,N_24705,N_24830);
or U25334 (N_25334,N_24831,N_25055);
and U25335 (N_25335,N_24240,N_24769);
xor U25336 (N_25336,N_24658,N_24628);
or U25337 (N_25337,N_24482,N_24232);
and U25338 (N_25338,N_25162,N_24299);
nand U25339 (N_25339,N_24462,N_24589);
nor U25340 (N_25340,N_24374,N_24451);
or U25341 (N_25341,N_24165,N_24694);
nor U25342 (N_25342,N_24748,N_24970);
or U25343 (N_25343,N_24915,N_24243);
nor U25344 (N_25344,N_24310,N_24942);
and U25345 (N_25345,N_24939,N_24563);
nor U25346 (N_25346,N_24030,N_24741);
and U25347 (N_25347,N_24881,N_24277);
xnor U25348 (N_25348,N_24385,N_25119);
xnor U25349 (N_25349,N_25124,N_24804);
nand U25350 (N_25350,N_24361,N_24158);
nand U25351 (N_25351,N_24926,N_24680);
or U25352 (N_25352,N_25165,N_24275);
and U25353 (N_25353,N_24313,N_24135);
xnor U25354 (N_25354,N_24084,N_24353);
nand U25355 (N_25355,N_24272,N_24848);
nor U25356 (N_25356,N_24500,N_24184);
nand U25357 (N_25357,N_24478,N_24306);
and U25358 (N_25358,N_24295,N_24796);
nand U25359 (N_25359,N_24561,N_24387);
nor U25360 (N_25360,N_24377,N_25023);
nand U25361 (N_25361,N_24916,N_24488);
nand U25362 (N_25362,N_24357,N_24489);
nor U25363 (N_25363,N_24358,N_24439);
xor U25364 (N_25364,N_24150,N_24246);
nand U25365 (N_25365,N_24688,N_24026);
nand U25366 (N_25366,N_24128,N_24664);
nor U25367 (N_25367,N_24679,N_25108);
nand U25368 (N_25368,N_24587,N_24549);
nor U25369 (N_25369,N_24719,N_24687);
or U25370 (N_25370,N_24386,N_24740);
xnor U25371 (N_25371,N_24983,N_24438);
nor U25372 (N_25372,N_24035,N_25146);
or U25373 (N_25373,N_24949,N_24566);
nand U25374 (N_25374,N_25160,N_24954);
and U25375 (N_25375,N_24843,N_24340);
or U25376 (N_25376,N_24009,N_24849);
nor U25377 (N_25377,N_24464,N_25102);
nor U25378 (N_25378,N_24157,N_24101);
nor U25379 (N_25379,N_24000,N_24710);
or U25380 (N_25380,N_25003,N_24261);
nand U25381 (N_25381,N_24656,N_24826);
or U25382 (N_25382,N_25000,N_24716);
or U25383 (N_25383,N_24497,N_24153);
nor U25384 (N_25384,N_24175,N_24149);
xnor U25385 (N_25385,N_24852,N_25048);
and U25386 (N_25386,N_24692,N_25141);
xnor U25387 (N_25387,N_24339,N_24457);
nor U25388 (N_25388,N_24421,N_24899);
nor U25389 (N_25389,N_24696,N_24707);
nand U25390 (N_25390,N_24943,N_24896);
xor U25391 (N_25391,N_24933,N_24978);
xor U25392 (N_25392,N_24351,N_24061);
nor U25393 (N_25393,N_24251,N_24155);
nand U25394 (N_25394,N_24642,N_24599);
and U25395 (N_25395,N_24392,N_25019);
xnor U25396 (N_25396,N_25033,N_24266);
nor U25397 (N_25397,N_24605,N_24889);
and U25398 (N_25398,N_24325,N_24422);
xnor U25399 (N_25399,N_25090,N_24423);
or U25400 (N_25400,N_24643,N_24514);
and U25401 (N_25401,N_25151,N_24647);
and U25402 (N_25402,N_25091,N_24616);
nand U25403 (N_25403,N_24783,N_25050);
or U25404 (N_25404,N_24593,N_24577);
nor U25405 (N_25405,N_25182,N_24269);
xor U25406 (N_25406,N_24190,N_25007);
nor U25407 (N_25407,N_24834,N_24219);
nor U25408 (N_25408,N_24847,N_24735);
or U25409 (N_25409,N_24728,N_24902);
xnor U25410 (N_25410,N_24559,N_24039);
or U25411 (N_25411,N_24560,N_24870);
xor U25412 (N_25412,N_25069,N_24104);
nand U25413 (N_25413,N_24542,N_24110);
and U25414 (N_25414,N_24839,N_24504);
xnor U25415 (N_25415,N_24032,N_24048);
nand U25416 (N_25416,N_24940,N_24573);
or U25417 (N_25417,N_24681,N_24652);
nor U25418 (N_25418,N_24536,N_25083);
and U25419 (N_25419,N_24888,N_24882);
or U25420 (N_25420,N_24763,N_24989);
xor U25421 (N_25421,N_24934,N_24701);
xnor U25422 (N_25422,N_24927,N_24920);
and U25423 (N_25423,N_24572,N_24140);
or U25424 (N_25424,N_25053,N_24754);
nand U25425 (N_25425,N_24021,N_24494);
xnor U25426 (N_25426,N_24418,N_24615);
or U25427 (N_25427,N_25034,N_25179);
nor U25428 (N_25428,N_24401,N_24132);
nand U25429 (N_25429,N_24279,N_24627);
and U25430 (N_25430,N_24886,N_24959);
or U25431 (N_25431,N_24591,N_24990);
or U25432 (N_25432,N_24756,N_24961);
or U25433 (N_25433,N_24670,N_24145);
xor U25434 (N_25434,N_25020,N_24354);
or U25435 (N_25435,N_24617,N_24619);
and U25436 (N_25436,N_24336,N_24880);
xnor U25437 (N_25437,N_24837,N_25004);
nor U25438 (N_25438,N_24760,N_24960);
xnor U25439 (N_25439,N_24767,N_25157);
nand U25440 (N_25440,N_24539,N_24236);
and U25441 (N_25441,N_24256,N_24100);
nor U25442 (N_25442,N_24292,N_24108);
nand U25443 (N_25443,N_24257,N_24524);
nor U25444 (N_25444,N_24874,N_24413);
nand U25445 (N_25445,N_24332,N_24320);
or U25446 (N_25446,N_24301,N_24076);
and U25447 (N_25447,N_24684,N_24971);
and U25448 (N_25448,N_25085,N_24033);
and U25449 (N_25449,N_24131,N_24006);
nand U25450 (N_25450,N_25024,N_25076);
nand U25451 (N_25451,N_24079,N_24237);
xnor U25452 (N_25452,N_24197,N_24063);
nor U25453 (N_25453,N_25115,N_24693);
nand U25454 (N_25454,N_24668,N_24527);
or U25455 (N_25455,N_25178,N_25169);
nor U25456 (N_25456,N_25080,N_24713);
or U25457 (N_25457,N_24750,N_24170);
nor U25458 (N_25458,N_24673,N_24141);
xor U25459 (N_25459,N_24571,N_25041);
xnor U25460 (N_25460,N_24969,N_24946);
nor U25461 (N_25461,N_24024,N_24194);
nand U25462 (N_25462,N_24055,N_24736);
nand U25463 (N_25463,N_24498,N_24651);
nor U25464 (N_25464,N_24662,N_25079);
xor U25465 (N_25465,N_24608,N_24534);
nand U25466 (N_25466,N_25180,N_24799);
and U25467 (N_25467,N_24911,N_24159);
xor U25468 (N_25468,N_25089,N_24102);
or U25469 (N_25469,N_24072,N_24363);
nand U25470 (N_25470,N_24168,N_25008);
nor U25471 (N_25471,N_24198,N_25186);
nor U25472 (N_25472,N_24068,N_24787);
nand U25473 (N_25473,N_25066,N_24672);
xnor U25474 (N_25474,N_24667,N_24683);
xor U25475 (N_25475,N_24775,N_24766);
and U25476 (N_25476,N_24835,N_24582);
and U25477 (N_25477,N_24201,N_24816);
or U25478 (N_25478,N_24119,N_24495);
xor U25479 (N_25479,N_24641,N_25059);
nand U25480 (N_25480,N_24267,N_25111);
nor U25481 (N_25481,N_24784,N_24156);
xnor U25482 (N_25482,N_25163,N_24109);
or U25483 (N_25483,N_24984,N_24877);
nand U25484 (N_25484,N_24535,N_24352);
nand U25485 (N_25485,N_24777,N_24574);
or U25486 (N_25486,N_24655,N_24025);
or U25487 (N_25487,N_24064,N_25088);
and U25488 (N_25488,N_24738,N_25194);
and U25489 (N_25489,N_24012,N_24808);
xnor U25490 (N_25490,N_24714,N_24208);
or U25491 (N_25491,N_24059,N_24085);
nor U25492 (N_25492,N_24176,N_24985);
nand U25493 (N_25493,N_24327,N_25116);
or U25494 (N_25494,N_24968,N_24832);
and U25495 (N_25495,N_24375,N_24928);
xor U25496 (N_25496,N_25071,N_24007);
nor U25497 (N_25497,N_24543,N_24245);
nand U25498 (N_25498,N_24597,N_25129);
nor U25499 (N_25499,N_24318,N_25009);
nand U25500 (N_25500,N_24986,N_24859);
xor U25501 (N_25501,N_25078,N_25103);
nor U25502 (N_25502,N_24058,N_24093);
nand U25503 (N_25503,N_24342,N_24424);
nand U25504 (N_25504,N_24409,N_25042);
or U25505 (N_25505,N_24356,N_24362);
nand U25506 (N_25506,N_25142,N_24388);
or U25507 (N_25507,N_25013,N_25171);
and U25508 (N_25508,N_25168,N_24105);
and U25509 (N_25509,N_24213,N_24298);
or U25510 (N_25510,N_24869,N_25101);
nor U25511 (N_25511,N_24999,N_24437);
nor U25512 (N_25512,N_24403,N_24345);
or U25513 (N_25513,N_24365,N_24618);
nor U25514 (N_25514,N_24436,N_24241);
nand U25515 (N_25515,N_24479,N_24174);
and U25516 (N_25516,N_24042,N_24178);
and U25517 (N_25517,N_24013,N_24551);
nand U25518 (N_25518,N_24098,N_24603);
nor U25519 (N_25519,N_24663,N_24062);
nand U25520 (N_25520,N_24067,N_24229);
nand U25521 (N_25521,N_24979,N_24759);
nand U25522 (N_25522,N_25132,N_24629);
nand U25523 (N_25523,N_24282,N_25189);
nor U25524 (N_25524,N_25173,N_24676);
or U25525 (N_25525,N_25127,N_25149);
xnor U25526 (N_25526,N_24263,N_24471);
xnor U25527 (N_25527,N_24887,N_24188);
xor U25528 (N_25528,N_25093,N_24465);
nand U25529 (N_25529,N_24416,N_24975);
nand U25530 (N_25530,N_24432,N_24260);
xnor U25531 (N_25531,N_25175,N_24891);
and U25532 (N_25532,N_24858,N_24879);
and U25533 (N_25533,N_25002,N_24815);
nand U25534 (N_25534,N_24782,N_24281);
xnor U25535 (N_25535,N_24020,N_25143);
and U25536 (N_25536,N_24519,N_24793);
and U25537 (N_25537,N_24950,N_24634);
and U25538 (N_25538,N_25049,N_24459);
or U25539 (N_25539,N_25029,N_24595);
and U25540 (N_25540,N_24060,N_25184);
and U25541 (N_25541,N_24221,N_25161);
or U25542 (N_25542,N_24623,N_24463);
and U25543 (N_25543,N_24690,N_25038);
nand U25544 (N_25544,N_24895,N_25094);
and U25545 (N_25545,N_24700,N_24065);
and U25546 (N_25546,N_24925,N_24094);
nand U25547 (N_25547,N_24429,N_24638);
or U25548 (N_25548,N_24431,N_24196);
xor U25549 (N_25549,N_24733,N_25052);
nor U25550 (N_25550,N_24581,N_24751);
and U25551 (N_25551,N_24704,N_24302);
nand U25552 (N_25552,N_24914,N_24936);
xnor U25553 (N_25553,N_24294,N_24541);
nand U25554 (N_25554,N_25152,N_24154);
and U25555 (N_25555,N_24337,N_25084);
or U25556 (N_25556,N_24614,N_25005);
or U25557 (N_25557,N_24976,N_24179);
or U25558 (N_25558,N_24312,N_24434);
and U25559 (N_25559,N_24333,N_24120);
xor U25560 (N_25560,N_24300,N_24776);
or U25561 (N_25561,N_24372,N_25011);
xnor U25562 (N_25562,N_24427,N_24370);
nor U25563 (N_25563,N_24182,N_24121);
xor U25564 (N_25564,N_24262,N_24308);
nor U25565 (N_25565,N_24097,N_24801);
nand U25566 (N_25566,N_24507,N_24601);
nand U25567 (N_25567,N_24709,N_25190);
and U25568 (N_25568,N_24225,N_25067);
nor U25569 (N_25569,N_25188,N_25025);
and U25570 (N_25570,N_24250,N_24450);
or U25571 (N_25571,N_24725,N_24991);
nor U25572 (N_25572,N_24364,N_24433);
nor U25573 (N_25573,N_25097,N_24677);
nor U25574 (N_25574,N_24841,N_25167);
nor U25575 (N_25575,N_24718,N_24475);
nor U25576 (N_25576,N_24411,N_24626);
or U25577 (N_25577,N_25140,N_24249);
nor U25578 (N_25578,N_25114,N_25139);
or U25579 (N_25579,N_24649,N_24328);
nor U25580 (N_25580,N_25037,N_24369);
nor U25581 (N_25581,N_24995,N_24379);
xor U25582 (N_25582,N_24860,N_24191);
nand U25583 (N_25583,N_24666,N_25054);
and U25584 (N_25584,N_24288,N_24752);
and U25585 (N_25585,N_25043,N_24788);
xor U25586 (N_25586,N_24910,N_25031);
and U25587 (N_25587,N_24125,N_24810);
nor U25588 (N_25588,N_24053,N_24114);
nand U25589 (N_25589,N_24781,N_24081);
and U25590 (N_25590,N_24646,N_24570);
and U25591 (N_25591,N_24089,N_24468);
nand U25592 (N_25592,N_24720,N_24948);
nand U25593 (N_25593,N_25137,N_24138);
or U25594 (N_25594,N_24631,N_24163);
nand U25595 (N_25595,N_24453,N_24648);
and U25596 (N_25596,N_24675,N_24620);
xnor U25597 (N_25597,N_24258,N_25130);
nor U25598 (N_25598,N_24338,N_24919);
and U25599 (N_25599,N_25121,N_24937);
nand U25600 (N_25600,N_24090,N_24472);
nand U25601 (N_25601,N_25181,N_24512);
nand U25602 (N_25602,N_24523,N_24774);
nor U25603 (N_25603,N_24054,N_24838);
nand U25604 (N_25604,N_24945,N_24923);
and U25605 (N_25605,N_24227,N_24334);
nand U25606 (N_25606,N_24348,N_24918);
xor U25607 (N_25607,N_24470,N_25086);
and U25608 (N_25608,N_24773,N_24765);
or U25609 (N_25609,N_24492,N_24594);
nand U25610 (N_25610,N_24415,N_24123);
xor U25611 (N_25611,N_24904,N_24082);
nor U25612 (N_25612,N_24454,N_24161);
xor U25613 (N_25613,N_25122,N_24930);
and U25614 (N_25614,N_24526,N_24739);
nand U25615 (N_25615,N_24729,N_25123);
xor U25616 (N_25616,N_24678,N_24407);
or U25617 (N_25617,N_24861,N_24066);
or U25618 (N_25618,N_24691,N_24271);
nand U25619 (N_25619,N_24218,N_24596);
xor U25620 (N_25620,N_24410,N_25074);
xnor U25621 (N_25621,N_24797,N_24077);
or U25622 (N_25622,N_24785,N_24622);
and U25623 (N_25623,N_24818,N_24167);
nand U25624 (N_25624,N_24903,N_24217);
xor U25625 (N_25625,N_24659,N_24865);
nor U25626 (N_25626,N_24964,N_25022);
or U25627 (N_25627,N_24180,N_24956);
nor U25628 (N_25628,N_24762,N_24518);
or U25629 (N_25629,N_25095,N_25077);
and U25630 (N_25630,N_24734,N_24477);
nand U25631 (N_25631,N_25172,N_25170);
xor U25632 (N_25632,N_25100,N_24532);
or U25633 (N_25633,N_25026,N_24823);
and U25634 (N_25634,N_25110,N_24069);
xnor U25635 (N_25635,N_24448,N_24430);
nand U25636 (N_25636,N_24613,N_24028);
or U25637 (N_25637,N_24419,N_25125);
nand U25638 (N_25638,N_24049,N_24380);
nand U25639 (N_25639,N_24307,N_25174);
and U25640 (N_25640,N_24420,N_24003);
and U25641 (N_25641,N_24160,N_25040);
or U25642 (N_25642,N_24324,N_24223);
xnor U25643 (N_25643,N_24244,N_24366);
nand U25644 (N_25644,N_24399,N_24322);
nor U25645 (N_25645,N_24254,N_24731);
and U25646 (N_25646,N_24669,N_24412);
or U25647 (N_25647,N_24997,N_25195);
xnor U25648 (N_25648,N_24080,N_24941);
nor U25649 (N_25649,N_24215,N_24144);
or U25650 (N_25650,N_24654,N_24029);
nand U25651 (N_25651,N_24682,N_24545);
and U25652 (N_25652,N_24764,N_24686);
nor U25653 (N_25653,N_24206,N_25128);
nand U25654 (N_25654,N_24505,N_25106);
and U25655 (N_25655,N_25098,N_24347);
and U25656 (N_25656,N_24398,N_24031);
and U25657 (N_25657,N_25118,N_24202);
nor U25658 (N_25658,N_24890,N_24270);
nor U25659 (N_25659,N_24554,N_24480);
nor U25660 (N_25660,N_24602,N_24253);
nor U25661 (N_25661,N_24255,N_24550);
or U25662 (N_25662,N_24425,N_24166);
nand U25663 (N_25663,N_24210,N_24537);
or U25664 (N_25664,N_24311,N_24908);
xor U25665 (N_25665,N_24562,N_24598);
xnor U25666 (N_25666,N_24274,N_24851);
xor U25667 (N_25667,N_24635,N_24611);
xnor U25668 (N_25668,N_24474,N_24285);
nor U25669 (N_25669,N_24181,N_24195);
or U25670 (N_25670,N_24034,N_24610);
or U25671 (N_25671,N_24665,N_24657);
nand U25672 (N_25672,N_25062,N_24341);
xnor U25673 (N_25673,N_24052,N_24235);
xnor U25674 (N_25674,N_24953,N_24513);
and U25675 (N_25675,N_24230,N_24484);
nor U25676 (N_25676,N_24640,N_24671);
nor U25677 (N_25677,N_24637,N_24293);
and U25678 (N_25678,N_24199,N_24134);
and U25679 (N_25679,N_24836,N_24929);
or U25680 (N_25680,N_24600,N_24753);
xnor U25681 (N_25681,N_24973,N_24010);
or U25682 (N_25682,N_24564,N_24726);
xnor U25683 (N_25683,N_24922,N_24744);
nand U25684 (N_25684,N_24522,N_24075);
xnor U25685 (N_25685,N_24547,N_25099);
or U25686 (N_25686,N_25126,N_24444);
or U25687 (N_25687,N_25045,N_24177);
nand U25688 (N_25688,N_25001,N_24892);
nand U25689 (N_25689,N_24576,N_24321);
or U25690 (N_25690,N_24248,N_24932);
or U25691 (N_25691,N_24967,N_24609);
xnor U25692 (N_25692,N_24127,N_24565);
xor U25693 (N_25693,N_24205,N_24632);
nor U25694 (N_25694,N_24531,N_24712);
nor U25695 (N_25695,N_24935,N_24568);
and U25696 (N_25696,N_24417,N_24343);
nor U25697 (N_25697,N_24095,N_25117);
nand U25698 (N_25698,N_24732,N_24786);
nor U25699 (N_25699,N_24994,N_24987);
and U25700 (N_25700,N_24730,N_24825);
nor U25701 (N_25701,N_24745,N_25134);
or U25702 (N_25702,N_24247,N_25081);
and U25703 (N_25703,N_24606,N_24747);
xor U25704 (N_25704,N_24073,N_24715);
and U25705 (N_25705,N_25150,N_25035);
nand U25706 (N_25706,N_24875,N_24326);
or U25707 (N_25707,N_24644,N_24373);
nand U25708 (N_25708,N_24695,N_24515);
nor U25709 (N_25709,N_24183,N_24636);
nand U25710 (N_25710,N_24078,N_24469);
or U25711 (N_25711,N_24216,N_24408);
or U25712 (N_25712,N_25144,N_25133);
nand U25713 (N_25713,N_24360,N_24405);
xor U25714 (N_25714,N_24086,N_24829);
nor U25715 (N_25715,N_25197,N_24344);
or U25716 (N_25716,N_25030,N_24151);
nor U25717 (N_25717,N_24809,N_24689);
nand U25718 (N_25718,N_24446,N_24907);
and U25719 (N_25719,N_24152,N_24529);
nor U25720 (N_25720,N_24962,N_24211);
xor U25721 (N_25721,N_24122,N_24789);
or U25722 (N_25722,N_24038,N_24817);
nor U25723 (N_25723,N_24228,N_25136);
or U25724 (N_25724,N_24117,N_24278);
xnor U25725 (N_25725,N_24557,N_24389);
and U25726 (N_25726,N_24807,N_24885);
xor U25727 (N_25727,N_24585,N_24864);
or U25728 (N_25728,N_25164,N_24708);
xor U25729 (N_25729,N_24368,N_24592);
or U25730 (N_25730,N_24143,N_24540);
or U25731 (N_25731,N_24905,N_24742);
and U25732 (N_25732,N_24721,N_24706);
nand U25733 (N_25733,N_24022,N_24209);
and U25734 (N_25734,N_24473,N_25058);
and U25735 (N_25735,N_25016,N_24924);
or U25736 (N_25736,N_24346,N_25057);
and U25737 (N_25737,N_24650,N_25196);
nor U25738 (N_25738,N_24791,N_25120);
or U25739 (N_25739,N_24083,N_24842);
xor U25740 (N_25740,N_24359,N_24517);
nand U25741 (N_25741,N_24222,N_24821);
and U25742 (N_25742,N_24685,N_24485);
xnor U25743 (N_25743,N_24002,N_24802);
or U25744 (N_25744,N_24909,N_24426);
and U25745 (N_25745,N_24814,N_24588);
and U25746 (N_25746,N_24812,N_24717);
and U25747 (N_25747,N_24625,N_24501);
nor U25748 (N_25748,N_24118,N_24074);
nor U25749 (N_25749,N_24854,N_24023);
xor U25750 (N_25750,N_24071,N_24827);
or U25751 (N_25751,N_24580,N_25036);
xor U25752 (N_25752,N_24499,N_24296);
nor U25753 (N_25753,N_24008,N_24977);
xnor U25754 (N_25754,N_24162,N_25191);
and U25755 (N_25755,N_24303,N_24853);
nor U25756 (N_25756,N_24460,N_24952);
nor U25757 (N_25757,N_24297,N_24091);
nand U25758 (N_25758,N_24400,N_24876);
nor U25759 (N_25759,N_24552,N_25156);
xnor U25760 (N_25760,N_24172,N_24016);
xor U25761 (N_25761,N_25104,N_24511);
nand U25762 (N_25762,N_24674,N_24883);
nor U25763 (N_25763,N_24314,N_24894);
or U25764 (N_25764,N_25075,N_25153);
nor U25765 (N_25765,N_24794,N_24711);
or U25766 (N_25766,N_24871,N_25021);
nor U25767 (N_25767,N_24330,N_24435);
nor U25768 (N_25768,N_24309,N_24037);
or U25769 (N_25769,N_25113,N_24276);
or U25770 (N_25770,N_24186,N_24291);
and U25771 (N_25771,N_24798,N_24702);
nand U25772 (N_25772,N_24284,N_24447);
and U25773 (N_25773,N_24516,N_24955);
nand U25774 (N_25774,N_24840,N_24015);
xnor U25775 (N_25775,N_24443,N_24528);
nor U25776 (N_25776,N_24287,N_24947);
nor U25777 (N_25777,N_24192,N_25056);
nor U25778 (N_25778,N_24757,N_24800);
xnor U25779 (N_25779,N_24041,N_25131);
nor U25780 (N_25780,N_24283,N_25087);
xnor U25781 (N_25781,N_24546,N_24502);
nand U25782 (N_25782,N_24442,N_24203);
and U25783 (N_25783,N_24921,N_24290);
nand U25784 (N_25784,N_24133,N_24018);
or U25785 (N_25785,N_24139,N_24173);
nand U25786 (N_25786,N_24204,N_24645);
xnor U25787 (N_25787,N_24639,N_25046);
nor U25788 (N_25788,N_24974,N_24850);
xnor U25789 (N_25789,N_24305,N_24778);
nand U25790 (N_25790,N_24456,N_24046);
nand U25791 (N_25791,N_24056,N_24575);
nand U25792 (N_25792,N_24224,N_24115);
nand U25793 (N_25793,N_24367,N_24189);
xor U25794 (N_25794,N_24391,N_24382);
nand U25795 (N_25795,N_24259,N_24857);
and U25796 (N_25796,N_24873,N_24335);
or U25797 (N_25797,N_24112,N_24395);
and U25798 (N_25798,N_24331,N_24897);
or U25799 (N_25799,N_24555,N_24242);
nor U25800 (N_25800,N_24576,N_25082);
and U25801 (N_25801,N_24154,N_24771);
and U25802 (N_25802,N_24774,N_25121);
nor U25803 (N_25803,N_24286,N_24524);
nand U25804 (N_25804,N_24969,N_24466);
and U25805 (N_25805,N_24281,N_24875);
or U25806 (N_25806,N_24953,N_24256);
nor U25807 (N_25807,N_24512,N_24158);
and U25808 (N_25808,N_24140,N_25020);
xor U25809 (N_25809,N_24408,N_24514);
and U25810 (N_25810,N_25165,N_24130);
xnor U25811 (N_25811,N_24398,N_24096);
nor U25812 (N_25812,N_24531,N_24664);
nor U25813 (N_25813,N_24733,N_24785);
and U25814 (N_25814,N_25148,N_24104);
xor U25815 (N_25815,N_25194,N_24647);
or U25816 (N_25816,N_25177,N_24837);
xnor U25817 (N_25817,N_24597,N_24384);
or U25818 (N_25818,N_24506,N_24473);
xnor U25819 (N_25819,N_24720,N_24911);
and U25820 (N_25820,N_25019,N_24882);
nor U25821 (N_25821,N_24370,N_25186);
and U25822 (N_25822,N_24666,N_24989);
nand U25823 (N_25823,N_24639,N_24277);
and U25824 (N_25824,N_24259,N_25198);
nand U25825 (N_25825,N_24951,N_24451);
or U25826 (N_25826,N_25072,N_24737);
nor U25827 (N_25827,N_24168,N_25089);
nor U25828 (N_25828,N_24590,N_24583);
or U25829 (N_25829,N_24845,N_24642);
and U25830 (N_25830,N_25198,N_25187);
nor U25831 (N_25831,N_24096,N_24754);
xor U25832 (N_25832,N_25179,N_24746);
xor U25833 (N_25833,N_25091,N_24409);
or U25834 (N_25834,N_24649,N_24499);
or U25835 (N_25835,N_24645,N_24800);
nor U25836 (N_25836,N_24115,N_24355);
and U25837 (N_25837,N_24252,N_24284);
nand U25838 (N_25838,N_24305,N_24164);
nor U25839 (N_25839,N_24779,N_24751);
and U25840 (N_25840,N_24850,N_24900);
nand U25841 (N_25841,N_25067,N_24768);
xor U25842 (N_25842,N_25125,N_24570);
xor U25843 (N_25843,N_24892,N_24274);
nand U25844 (N_25844,N_24680,N_24712);
nor U25845 (N_25845,N_24721,N_24845);
nor U25846 (N_25846,N_24512,N_24290);
or U25847 (N_25847,N_24409,N_25013);
nor U25848 (N_25848,N_24218,N_24275);
nor U25849 (N_25849,N_24421,N_24210);
nor U25850 (N_25850,N_24556,N_24780);
and U25851 (N_25851,N_24938,N_24180);
nor U25852 (N_25852,N_24554,N_24519);
xor U25853 (N_25853,N_24020,N_24304);
and U25854 (N_25854,N_24513,N_25157);
nor U25855 (N_25855,N_24160,N_24262);
nand U25856 (N_25856,N_24760,N_24204);
and U25857 (N_25857,N_24527,N_25115);
xnor U25858 (N_25858,N_24728,N_25069);
nand U25859 (N_25859,N_24227,N_24125);
and U25860 (N_25860,N_24250,N_24983);
nor U25861 (N_25861,N_25139,N_24143);
or U25862 (N_25862,N_24638,N_24531);
nand U25863 (N_25863,N_24105,N_24027);
xnor U25864 (N_25864,N_24961,N_24060);
and U25865 (N_25865,N_24833,N_25022);
and U25866 (N_25866,N_25193,N_24133);
or U25867 (N_25867,N_24433,N_25115);
or U25868 (N_25868,N_25159,N_24946);
nand U25869 (N_25869,N_24464,N_24754);
and U25870 (N_25870,N_25199,N_24755);
nand U25871 (N_25871,N_24721,N_24066);
nor U25872 (N_25872,N_24538,N_24009);
nand U25873 (N_25873,N_24073,N_25053);
nand U25874 (N_25874,N_24088,N_24712);
nor U25875 (N_25875,N_25189,N_24734);
nand U25876 (N_25876,N_25013,N_24197);
or U25877 (N_25877,N_24784,N_25108);
and U25878 (N_25878,N_24569,N_24752);
xnor U25879 (N_25879,N_25063,N_25131);
nand U25880 (N_25880,N_24859,N_24210);
and U25881 (N_25881,N_24176,N_25071);
or U25882 (N_25882,N_24254,N_25075);
and U25883 (N_25883,N_25058,N_24199);
nand U25884 (N_25884,N_24311,N_24858);
nor U25885 (N_25885,N_24049,N_24464);
or U25886 (N_25886,N_24408,N_24351);
xnor U25887 (N_25887,N_25033,N_25073);
and U25888 (N_25888,N_24872,N_24645);
or U25889 (N_25889,N_24634,N_24159);
and U25890 (N_25890,N_24062,N_24043);
or U25891 (N_25891,N_24136,N_24488);
and U25892 (N_25892,N_24325,N_24085);
nand U25893 (N_25893,N_24681,N_24644);
or U25894 (N_25894,N_24128,N_24652);
nand U25895 (N_25895,N_24949,N_24347);
xnor U25896 (N_25896,N_24877,N_24132);
nor U25897 (N_25897,N_25088,N_24845);
or U25898 (N_25898,N_24417,N_24427);
or U25899 (N_25899,N_24772,N_24744);
or U25900 (N_25900,N_24684,N_24909);
xnor U25901 (N_25901,N_24579,N_24264);
nand U25902 (N_25902,N_24729,N_24471);
or U25903 (N_25903,N_24234,N_24836);
xor U25904 (N_25904,N_24870,N_24256);
nor U25905 (N_25905,N_24158,N_25167);
nor U25906 (N_25906,N_24833,N_24672);
and U25907 (N_25907,N_24987,N_24677);
nor U25908 (N_25908,N_24020,N_24920);
or U25909 (N_25909,N_24200,N_25158);
xor U25910 (N_25910,N_24375,N_24911);
and U25911 (N_25911,N_24296,N_24431);
or U25912 (N_25912,N_25185,N_24139);
and U25913 (N_25913,N_24610,N_25198);
or U25914 (N_25914,N_24632,N_24617);
or U25915 (N_25915,N_24393,N_24100);
or U25916 (N_25916,N_25024,N_24616);
nor U25917 (N_25917,N_24931,N_24657);
and U25918 (N_25918,N_24538,N_25146);
xnor U25919 (N_25919,N_24639,N_25165);
xor U25920 (N_25920,N_24601,N_24864);
xor U25921 (N_25921,N_24009,N_24795);
xnor U25922 (N_25922,N_24969,N_24226);
nand U25923 (N_25923,N_24446,N_24974);
xnor U25924 (N_25924,N_24145,N_24236);
or U25925 (N_25925,N_24444,N_25013);
nor U25926 (N_25926,N_24519,N_24227);
and U25927 (N_25927,N_24582,N_25141);
nand U25928 (N_25928,N_24858,N_24722);
or U25929 (N_25929,N_24849,N_25029);
or U25930 (N_25930,N_24356,N_24678);
nor U25931 (N_25931,N_24592,N_24717);
xnor U25932 (N_25932,N_24693,N_24406);
nand U25933 (N_25933,N_24345,N_24084);
or U25934 (N_25934,N_24662,N_24597);
nor U25935 (N_25935,N_24019,N_24087);
nand U25936 (N_25936,N_24927,N_24905);
or U25937 (N_25937,N_24797,N_24240);
nor U25938 (N_25938,N_25145,N_24209);
nand U25939 (N_25939,N_24807,N_24631);
xor U25940 (N_25940,N_24880,N_25096);
nand U25941 (N_25941,N_25098,N_25174);
nand U25942 (N_25942,N_24416,N_24862);
nand U25943 (N_25943,N_24035,N_25175);
nand U25944 (N_25944,N_24582,N_24328);
xnor U25945 (N_25945,N_24679,N_24694);
or U25946 (N_25946,N_24049,N_24017);
or U25947 (N_25947,N_24606,N_24835);
xor U25948 (N_25948,N_24223,N_24494);
xor U25949 (N_25949,N_25148,N_24350);
or U25950 (N_25950,N_24286,N_24000);
or U25951 (N_25951,N_25148,N_24452);
nand U25952 (N_25952,N_24222,N_24754);
nand U25953 (N_25953,N_24885,N_24456);
xor U25954 (N_25954,N_24137,N_24535);
and U25955 (N_25955,N_24946,N_24631);
nand U25956 (N_25956,N_24940,N_24477);
xor U25957 (N_25957,N_24868,N_24557);
nor U25958 (N_25958,N_24523,N_24400);
nor U25959 (N_25959,N_24850,N_24735);
or U25960 (N_25960,N_24092,N_24829);
nand U25961 (N_25961,N_25104,N_25137);
nor U25962 (N_25962,N_25127,N_24473);
xor U25963 (N_25963,N_24109,N_24343);
xor U25964 (N_25964,N_24087,N_24131);
and U25965 (N_25965,N_24435,N_24761);
and U25966 (N_25966,N_25132,N_25073);
nor U25967 (N_25967,N_24580,N_24218);
xor U25968 (N_25968,N_24984,N_24614);
and U25969 (N_25969,N_24802,N_25049);
xnor U25970 (N_25970,N_24460,N_24919);
xor U25971 (N_25971,N_24959,N_24183);
and U25972 (N_25972,N_24080,N_24804);
nand U25973 (N_25973,N_24009,N_24575);
nor U25974 (N_25974,N_24144,N_24890);
or U25975 (N_25975,N_24941,N_24940);
and U25976 (N_25976,N_25148,N_24225);
xnor U25977 (N_25977,N_24355,N_24479);
nor U25978 (N_25978,N_25115,N_25110);
or U25979 (N_25979,N_24441,N_24137);
nor U25980 (N_25980,N_24755,N_24332);
xnor U25981 (N_25981,N_24266,N_24301);
nor U25982 (N_25982,N_25084,N_24028);
or U25983 (N_25983,N_24696,N_24327);
nor U25984 (N_25984,N_24689,N_24968);
or U25985 (N_25985,N_24663,N_24329);
nor U25986 (N_25986,N_24221,N_24934);
and U25987 (N_25987,N_24358,N_24836);
or U25988 (N_25988,N_24131,N_25199);
and U25989 (N_25989,N_25014,N_24419);
or U25990 (N_25990,N_24552,N_24487);
or U25991 (N_25991,N_24637,N_24378);
xnor U25992 (N_25992,N_24651,N_24546);
nand U25993 (N_25993,N_24927,N_24286);
or U25994 (N_25994,N_25085,N_25051);
or U25995 (N_25995,N_25181,N_24058);
nor U25996 (N_25996,N_24158,N_25007);
nor U25997 (N_25997,N_24952,N_24734);
or U25998 (N_25998,N_24750,N_24040);
nor U25999 (N_25999,N_24704,N_24715);
nor U26000 (N_26000,N_24026,N_24638);
nor U26001 (N_26001,N_25069,N_25098);
nor U26002 (N_26002,N_24390,N_24935);
nand U26003 (N_26003,N_24754,N_24187);
or U26004 (N_26004,N_24386,N_24047);
nand U26005 (N_26005,N_24728,N_24218);
nand U26006 (N_26006,N_25070,N_24078);
or U26007 (N_26007,N_24991,N_24538);
xnor U26008 (N_26008,N_24381,N_24028);
nor U26009 (N_26009,N_24411,N_24468);
xnor U26010 (N_26010,N_25124,N_24207);
nand U26011 (N_26011,N_25196,N_24606);
nand U26012 (N_26012,N_24235,N_24702);
xor U26013 (N_26013,N_24507,N_24619);
xor U26014 (N_26014,N_24676,N_24135);
and U26015 (N_26015,N_24003,N_24380);
nor U26016 (N_26016,N_24207,N_25150);
nand U26017 (N_26017,N_24022,N_24918);
nand U26018 (N_26018,N_24170,N_24662);
or U26019 (N_26019,N_24611,N_24551);
xnor U26020 (N_26020,N_24088,N_24010);
nor U26021 (N_26021,N_24039,N_25140);
nand U26022 (N_26022,N_25159,N_24407);
nor U26023 (N_26023,N_24927,N_24586);
nor U26024 (N_26024,N_24098,N_24233);
and U26025 (N_26025,N_25168,N_24212);
xor U26026 (N_26026,N_24915,N_24563);
or U26027 (N_26027,N_24674,N_25112);
and U26028 (N_26028,N_24176,N_24944);
or U26029 (N_26029,N_25105,N_24818);
and U26030 (N_26030,N_24275,N_24637);
or U26031 (N_26031,N_24591,N_24746);
nand U26032 (N_26032,N_25087,N_24928);
nand U26033 (N_26033,N_24157,N_24944);
or U26034 (N_26034,N_24202,N_24734);
nor U26035 (N_26035,N_24197,N_24409);
nor U26036 (N_26036,N_24293,N_25174);
xnor U26037 (N_26037,N_24541,N_24767);
or U26038 (N_26038,N_24113,N_24538);
xnor U26039 (N_26039,N_24818,N_24170);
and U26040 (N_26040,N_24278,N_24172);
xnor U26041 (N_26041,N_25020,N_24432);
nor U26042 (N_26042,N_24658,N_24994);
nand U26043 (N_26043,N_24120,N_24191);
or U26044 (N_26044,N_24477,N_24950);
nor U26045 (N_26045,N_24117,N_25055);
xnor U26046 (N_26046,N_25014,N_25031);
xor U26047 (N_26047,N_25058,N_24854);
or U26048 (N_26048,N_24871,N_25085);
or U26049 (N_26049,N_24203,N_24634);
nand U26050 (N_26050,N_24445,N_24841);
nor U26051 (N_26051,N_24318,N_24817);
and U26052 (N_26052,N_24540,N_24573);
xor U26053 (N_26053,N_24314,N_24328);
or U26054 (N_26054,N_24394,N_25094);
nor U26055 (N_26055,N_24600,N_24155);
xnor U26056 (N_26056,N_24862,N_24444);
xor U26057 (N_26057,N_24172,N_25025);
nand U26058 (N_26058,N_24301,N_25174);
nand U26059 (N_26059,N_24753,N_24929);
nand U26060 (N_26060,N_24230,N_24652);
nor U26061 (N_26061,N_24555,N_24939);
nor U26062 (N_26062,N_24642,N_25001);
or U26063 (N_26063,N_24667,N_24044);
nand U26064 (N_26064,N_25017,N_24969);
nor U26065 (N_26065,N_24671,N_24025);
or U26066 (N_26066,N_25080,N_24418);
nand U26067 (N_26067,N_24099,N_24285);
xor U26068 (N_26068,N_24642,N_24310);
and U26069 (N_26069,N_24293,N_24903);
and U26070 (N_26070,N_24981,N_24219);
and U26071 (N_26071,N_24543,N_24105);
or U26072 (N_26072,N_24805,N_24070);
nand U26073 (N_26073,N_24380,N_24755);
nor U26074 (N_26074,N_24797,N_25097);
nand U26075 (N_26075,N_24573,N_24719);
nand U26076 (N_26076,N_24691,N_25074);
nand U26077 (N_26077,N_24522,N_24940);
nor U26078 (N_26078,N_24904,N_24878);
nor U26079 (N_26079,N_24202,N_24707);
or U26080 (N_26080,N_24371,N_25134);
and U26081 (N_26081,N_24199,N_24818);
nor U26082 (N_26082,N_24931,N_24354);
xnor U26083 (N_26083,N_24581,N_24454);
nor U26084 (N_26084,N_24735,N_24105);
nor U26085 (N_26085,N_24491,N_24985);
and U26086 (N_26086,N_24229,N_24594);
or U26087 (N_26087,N_24048,N_24617);
nor U26088 (N_26088,N_24037,N_24064);
or U26089 (N_26089,N_24992,N_24076);
nor U26090 (N_26090,N_24693,N_24850);
nand U26091 (N_26091,N_24125,N_25148);
xnor U26092 (N_26092,N_25153,N_24973);
xor U26093 (N_26093,N_24204,N_24737);
xor U26094 (N_26094,N_24413,N_24409);
nor U26095 (N_26095,N_25080,N_24064);
or U26096 (N_26096,N_24513,N_24064);
nor U26097 (N_26097,N_24195,N_24631);
or U26098 (N_26098,N_24569,N_24759);
nand U26099 (N_26099,N_24166,N_24157);
and U26100 (N_26100,N_24166,N_24273);
nand U26101 (N_26101,N_24316,N_24875);
nand U26102 (N_26102,N_24157,N_24126);
nor U26103 (N_26103,N_24300,N_24360);
nand U26104 (N_26104,N_24733,N_24892);
nor U26105 (N_26105,N_24971,N_24182);
xor U26106 (N_26106,N_25144,N_24420);
nor U26107 (N_26107,N_24717,N_25196);
xor U26108 (N_26108,N_25197,N_24788);
xnor U26109 (N_26109,N_24838,N_24176);
xnor U26110 (N_26110,N_25108,N_24522);
nand U26111 (N_26111,N_24012,N_24980);
xnor U26112 (N_26112,N_24619,N_24939);
nand U26113 (N_26113,N_24414,N_24804);
nand U26114 (N_26114,N_25181,N_24572);
nor U26115 (N_26115,N_24210,N_25054);
and U26116 (N_26116,N_24957,N_24784);
and U26117 (N_26117,N_24619,N_24260);
xor U26118 (N_26118,N_24154,N_24201);
and U26119 (N_26119,N_25132,N_24077);
nand U26120 (N_26120,N_24838,N_25198);
xnor U26121 (N_26121,N_24361,N_25071);
or U26122 (N_26122,N_24976,N_24451);
or U26123 (N_26123,N_24273,N_25028);
nand U26124 (N_26124,N_24661,N_24329);
nor U26125 (N_26125,N_24232,N_25123);
nand U26126 (N_26126,N_24414,N_24562);
nor U26127 (N_26127,N_24677,N_24869);
nand U26128 (N_26128,N_25053,N_24818);
nor U26129 (N_26129,N_24105,N_24091);
nand U26130 (N_26130,N_24408,N_25012);
xnor U26131 (N_26131,N_24466,N_24154);
nor U26132 (N_26132,N_24492,N_24558);
nand U26133 (N_26133,N_24086,N_24853);
nor U26134 (N_26134,N_24352,N_25068);
nor U26135 (N_26135,N_24789,N_24232);
xnor U26136 (N_26136,N_25152,N_24739);
or U26137 (N_26137,N_24056,N_24267);
nor U26138 (N_26138,N_24731,N_25050);
xor U26139 (N_26139,N_24101,N_24413);
nor U26140 (N_26140,N_24798,N_24988);
and U26141 (N_26141,N_24094,N_25054);
and U26142 (N_26142,N_25010,N_24121);
xnor U26143 (N_26143,N_24555,N_24835);
and U26144 (N_26144,N_24116,N_24150);
xnor U26145 (N_26145,N_24264,N_25067);
xnor U26146 (N_26146,N_24030,N_25049);
nand U26147 (N_26147,N_24804,N_24152);
or U26148 (N_26148,N_25124,N_24199);
or U26149 (N_26149,N_25095,N_24017);
xnor U26150 (N_26150,N_24233,N_25190);
nand U26151 (N_26151,N_25151,N_24739);
or U26152 (N_26152,N_25052,N_24602);
nand U26153 (N_26153,N_24550,N_24858);
nor U26154 (N_26154,N_24832,N_25154);
nor U26155 (N_26155,N_24710,N_24874);
nand U26156 (N_26156,N_25014,N_24188);
or U26157 (N_26157,N_25196,N_24085);
or U26158 (N_26158,N_24912,N_24147);
and U26159 (N_26159,N_24186,N_24518);
nor U26160 (N_26160,N_24913,N_24962);
and U26161 (N_26161,N_24297,N_24380);
nand U26162 (N_26162,N_25089,N_24982);
nand U26163 (N_26163,N_24306,N_24335);
nor U26164 (N_26164,N_24109,N_25138);
xor U26165 (N_26165,N_24610,N_24111);
and U26166 (N_26166,N_24535,N_24806);
nand U26167 (N_26167,N_24408,N_25053);
and U26168 (N_26168,N_25045,N_24925);
nor U26169 (N_26169,N_24126,N_24823);
xor U26170 (N_26170,N_24973,N_24247);
and U26171 (N_26171,N_24666,N_24723);
and U26172 (N_26172,N_24203,N_24643);
nand U26173 (N_26173,N_24132,N_24527);
xnor U26174 (N_26174,N_24822,N_24331);
nor U26175 (N_26175,N_24556,N_24148);
xnor U26176 (N_26176,N_24533,N_24215);
xnor U26177 (N_26177,N_25093,N_24642);
nor U26178 (N_26178,N_25004,N_24851);
nand U26179 (N_26179,N_24546,N_24904);
nand U26180 (N_26180,N_24935,N_24238);
nand U26181 (N_26181,N_24408,N_25191);
nor U26182 (N_26182,N_24324,N_25046);
or U26183 (N_26183,N_24091,N_24988);
xnor U26184 (N_26184,N_24473,N_24866);
nor U26185 (N_26185,N_24779,N_24193);
xnor U26186 (N_26186,N_24124,N_24826);
or U26187 (N_26187,N_24220,N_24611);
or U26188 (N_26188,N_24337,N_25095);
nand U26189 (N_26189,N_24765,N_24856);
and U26190 (N_26190,N_25007,N_24690);
xor U26191 (N_26191,N_24202,N_24478);
nor U26192 (N_26192,N_24300,N_24790);
xnor U26193 (N_26193,N_24491,N_25039);
xor U26194 (N_26194,N_24155,N_24364);
and U26195 (N_26195,N_24009,N_25087);
nor U26196 (N_26196,N_24791,N_24896);
xnor U26197 (N_26197,N_24304,N_25049);
or U26198 (N_26198,N_24896,N_24834);
and U26199 (N_26199,N_24538,N_24038);
nand U26200 (N_26200,N_24146,N_24351);
nor U26201 (N_26201,N_24174,N_24170);
xnor U26202 (N_26202,N_24473,N_24362);
xor U26203 (N_26203,N_24625,N_24715);
and U26204 (N_26204,N_24093,N_24735);
or U26205 (N_26205,N_24761,N_24710);
nand U26206 (N_26206,N_24717,N_24111);
xor U26207 (N_26207,N_24592,N_24117);
and U26208 (N_26208,N_24011,N_24984);
and U26209 (N_26209,N_24217,N_24373);
xor U26210 (N_26210,N_24318,N_25175);
nor U26211 (N_26211,N_24762,N_24744);
xnor U26212 (N_26212,N_24839,N_24922);
nor U26213 (N_26213,N_24226,N_24024);
nor U26214 (N_26214,N_25020,N_24301);
nand U26215 (N_26215,N_24492,N_24777);
nor U26216 (N_26216,N_24987,N_25168);
nor U26217 (N_26217,N_24229,N_25184);
or U26218 (N_26218,N_24658,N_24627);
xnor U26219 (N_26219,N_24351,N_24341);
nand U26220 (N_26220,N_25034,N_24064);
nand U26221 (N_26221,N_24450,N_24577);
and U26222 (N_26222,N_24158,N_24080);
or U26223 (N_26223,N_25061,N_24509);
and U26224 (N_26224,N_24471,N_24940);
or U26225 (N_26225,N_24634,N_24606);
and U26226 (N_26226,N_24803,N_24597);
and U26227 (N_26227,N_24177,N_24606);
nand U26228 (N_26228,N_24140,N_24184);
xor U26229 (N_26229,N_24318,N_24874);
nor U26230 (N_26230,N_25076,N_24140);
xor U26231 (N_26231,N_24890,N_25077);
and U26232 (N_26232,N_24926,N_24786);
nand U26233 (N_26233,N_24369,N_25002);
xnor U26234 (N_26234,N_24738,N_24074);
and U26235 (N_26235,N_24687,N_24101);
xnor U26236 (N_26236,N_24062,N_25173);
nor U26237 (N_26237,N_24673,N_24822);
nor U26238 (N_26238,N_24899,N_24580);
nand U26239 (N_26239,N_24133,N_24775);
nor U26240 (N_26240,N_24040,N_24432);
or U26241 (N_26241,N_24708,N_25182);
and U26242 (N_26242,N_25131,N_24829);
or U26243 (N_26243,N_25117,N_24212);
and U26244 (N_26244,N_24584,N_24224);
nand U26245 (N_26245,N_24421,N_24463);
nand U26246 (N_26246,N_24926,N_24862);
nor U26247 (N_26247,N_24517,N_24449);
and U26248 (N_26248,N_24312,N_24143);
nor U26249 (N_26249,N_24291,N_25027);
and U26250 (N_26250,N_24466,N_24845);
nor U26251 (N_26251,N_24547,N_24189);
nor U26252 (N_26252,N_24843,N_24625);
xnor U26253 (N_26253,N_24890,N_24068);
nor U26254 (N_26254,N_25184,N_25056);
and U26255 (N_26255,N_24534,N_24762);
nor U26256 (N_26256,N_24952,N_25031);
nand U26257 (N_26257,N_24986,N_25021);
nand U26258 (N_26258,N_24358,N_24600);
xor U26259 (N_26259,N_24105,N_25192);
nor U26260 (N_26260,N_24828,N_24211);
and U26261 (N_26261,N_24877,N_25050);
nand U26262 (N_26262,N_24702,N_24957);
nor U26263 (N_26263,N_24002,N_25054);
and U26264 (N_26264,N_24735,N_24904);
or U26265 (N_26265,N_24380,N_24861);
nand U26266 (N_26266,N_24493,N_24293);
nor U26267 (N_26267,N_24529,N_24616);
and U26268 (N_26268,N_24049,N_24835);
nand U26269 (N_26269,N_24050,N_24761);
nor U26270 (N_26270,N_24895,N_24222);
xnor U26271 (N_26271,N_24508,N_25111);
and U26272 (N_26272,N_24747,N_24668);
and U26273 (N_26273,N_24536,N_24288);
or U26274 (N_26274,N_25135,N_24458);
or U26275 (N_26275,N_24043,N_25182);
and U26276 (N_26276,N_24984,N_24847);
and U26277 (N_26277,N_24818,N_24782);
or U26278 (N_26278,N_25049,N_24833);
nor U26279 (N_26279,N_24044,N_25148);
and U26280 (N_26280,N_24181,N_25008);
nor U26281 (N_26281,N_24998,N_24062);
nand U26282 (N_26282,N_25025,N_24251);
xnor U26283 (N_26283,N_24750,N_25030);
and U26284 (N_26284,N_24758,N_24347);
nor U26285 (N_26285,N_24434,N_24394);
nor U26286 (N_26286,N_25019,N_25089);
nor U26287 (N_26287,N_24496,N_24089);
and U26288 (N_26288,N_24950,N_24359);
nand U26289 (N_26289,N_24166,N_25081);
and U26290 (N_26290,N_25078,N_25026);
nand U26291 (N_26291,N_24871,N_25099);
and U26292 (N_26292,N_24491,N_24652);
or U26293 (N_26293,N_24719,N_25017);
nand U26294 (N_26294,N_24563,N_24252);
xor U26295 (N_26295,N_24939,N_24474);
xor U26296 (N_26296,N_24784,N_24924);
nand U26297 (N_26297,N_24004,N_24255);
nand U26298 (N_26298,N_24002,N_24135);
and U26299 (N_26299,N_24423,N_24455);
and U26300 (N_26300,N_24280,N_24831);
nand U26301 (N_26301,N_25055,N_24747);
and U26302 (N_26302,N_25117,N_24162);
or U26303 (N_26303,N_24993,N_24301);
or U26304 (N_26304,N_24800,N_24780);
xor U26305 (N_26305,N_24917,N_24962);
and U26306 (N_26306,N_24667,N_24839);
xor U26307 (N_26307,N_24801,N_24107);
nor U26308 (N_26308,N_24041,N_24279);
xor U26309 (N_26309,N_24488,N_25120);
nand U26310 (N_26310,N_24236,N_24700);
nor U26311 (N_26311,N_24283,N_24385);
and U26312 (N_26312,N_24536,N_25196);
nor U26313 (N_26313,N_24933,N_24287);
and U26314 (N_26314,N_25195,N_24780);
nand U26315 (N_26315,N_24777,N_24824);
and U26316 (N_26316,N_24631,N_24010);
or U26317 (N_26317,N_25064,N_24342);
or U26318 (N_26318,N_24460,N_25160);
xnor U26319 (N_26319,N_24133,N_24683);
nand U26320 (N_26320,N_24682,N_24275);
xnor U26321 (N_26321,N_25181,N_24465);
xor U26322 (N_26322,N_24748,N_25075);
nor U26323 (N_26323,N_24765,N_25111);
xor U26324 (N_26324,N_24971,N_25057);
or U26325 (N_26325,N_24127,N_24460);
nand U26326 (N_26326,N_24750,N_24108);
nor U26327 (N_26327,N_25007,N_24548);
or U26328 (N_26328,N_24799,N_24726);
or U26329 (N_26329,N_24618,N_24547);
or U26330 (N_26330,N_24925,N_24096);
nand U26331 (N_26331,N_24113,N_24874);
and U26332 (N_26332,N_25024,N_24470);
xnor U26333 (N_26333,N_24298,N_24230);
and U26334 (N_26334,N_24300,N_24584);
nand U26335 (N_26335,N_25066,N_24462);
nor U26336 (N_26336,N_25014,N_24183);
and U26337 (N_26337,N_25000,N_24634);
or U26338 (N_26338,N_24952,N_24788);
and U26339 (N_26339,N_24443,N_24332);
xnor U26340 (N_26340,N_24713,N_24345);
or U26341 (N_26341,N_24677,N_25018);
nand U26342 (N_26342,N_24274,N_24292);
or U26343 (N_26343,N_24586,N_24089);
xnor U26344 (N_26344,N_24605,N_24933);
nand U26345 (N_26345,N_24389,N_24569);
nor U26346 (N_26346,N_24818,N_24872);
nor U26347 (N_26347,N_25196,N_24477);
or U26348 (N_26348,N_24862,N_25194);
and U26349 (N_26349,N_24162,N_24349);
xnor U26350 (N_26350,N_24780,N_24099);
nor U26351 (N_26351,N_24606,N_24215);
xnor U26352 (N_26352,N_24003,N_25004);
nand U26353 (N_26353,N_24286,N_24409);
or U26354 (N_26354,N_24500,N_24789);
nand U26355 (N_26355,N_24287,N_24559);
and U26356 (N_26356,N_24743,N_25145);
or U26357 (N_26357,N_24673,N_24801);
nor U26358 (N_26358,N_24330,N_24121);
or U26359 (N_26359,N_24536,N_24887);
nand U26360 (N_26360,N_24061,N_24555);
nand U26361 (N_26361,N_24730,N_24479);
and U26362 (N_26362,N_25159,N_24045);
nor U26363 (N_26363,N_24674,N_24227);
xnor U26364 (N_26364,N_24843,N_24648);
or U26365 (N_26365,N_25063,N_24911);
nand U26366 (N_26366,N_24075,N_24238);
or U26367 (N_26367,N_24238,N_24995);
xor U26368 (N_26368,N_25069,N_24317);
or U26369 (N_26369,N_24481,N_24773);
xnor U26370 (N_26370,N_24053,N_24668);
and U26371 (N_26371,N_24862,N_24178);
nand U26372 (N_26372,N_24456,N_24780);
xor U26373 (N_26373,N_24894,N_24380);
xor U26374 (N_26374,N_24660,N_25177);
nor U26375 (N_26375,N_24668,N_24786);
and U26376 (N_26376,N_24057,N_24490);
nor U26377 (N_26377,N_24551,N_24882);
xnor U26378 (N_26378,N_25156,N_24976);
or U26379 (N_26379,N_25168,N_24307);
xnor U26380 (N_26380,N_24399,N_24914);
and U26381 (N_26381,N_24634,N_24593);
or U26382 (N_26382,N_24770,N_24079);
or U26383 (N_26383,N_24495,N_25177);
and U26384 (N_26384,N_25112,N_24898);
and U26385 (N_26385,N_24288,N_24755);
nor U26386 (N_26386,N_25074,N_24065);
and U26387 (N_26387,N_24483,N_24135);
nand U26388 (N_26388,N_24301,N_24351);
nor U26389 (N_26389,N_24184,N_24792);
nand U26390 (N_26390,N_25196,N_24227);
and U26391 (N_26391,N_24008,N_24126);
and U26392 (N_26392,N_24458,N_24131);
nor U26393 (N_26393,N_24383,N_25195);
nand U26394 (N_26394,N_24789,N_25119);
nand U26395 (N_26395,N_24332,N_24739);
nand U26396 (N_26396,N_24130,N_24027);
and U26397 (N_26397,N_24018,N_24323);
nand U26398 (N_26398,N_24918,N_24189);
nand U26399 (N_26399,N_24075,N_24953);
and U26400 (N_26400,N_25368,N_26332);
nand U26401 (N_26401,N_25343,N_25875);
xnor U26402 (N_26402,N_25246,N_26174);
xor U26403 (N_26403,N_26147,N_25876);
nor U26404 (N_26404,N_25399,N_25581);
or U26405 (N_26405,N_25723,N_25441);
and U26406 (N_26406,N_25854,N_26200);
xnor U26407 (N_26407,N_25228,N_25743);
xor U26408 (N_26408,N_25548,N_25408);
and U26409 (N_26409,N_25921,N_25223);
and U26410 (N_26410,N_25862,N_25387);
or U26411 (N_26411,N_25637,N_25430);
nand U26412 (N_26412,N_26366,N_25473);
or U26413 (N_26413,N_25766,N_26377);
nand U26414 (N_26414,N_25678,N_26273);
and U26415 (N_26415,N_25322,N_25493);
nand U26416 (N_26416,N_25376,N_25627);
and U26417 (N_26417,N_26322,N_25331);
and U26418 (N_26418,N_25730,N_25792);
nor U26419 (N_26419,N_25756,N_25964);
nor U26420 (N_26420,N_25934,N_25729);
or U26421 (N_26421,N_25489,N_25334);
and U26422 (N_26422,N_25931,N_26348);
nor U26423 (N_26423,N_25825,N_25380);
and U26424 (N_26424,N_26091,N_25918);
nand U26425 (N_26425,N_25667,N_25783);
and U26426 (N_26426,N_26110,N_25971);
or U26427 (N_26427,N_26098,N_25495);
and U26428 (N_26428,N_25497,N_26338);
xor U26429 (N_26429,N_25390,N_26001);
nand U26430 (N_26430,N_25919,N_26151);
nand U26431 (N_26431,N_25311,N_25313);
nor U26432 (N_26432,N_26025,N_26029);
nand U26433 (N_26433,N_25321,N_26240);
nor U26434 (N_26434,N_25680,N_26372);
nor U26435 (N_26435,N_26284,N_25274);
xnor U26436 (N_26436,N_26289,N_25780);
and U26437 (N_26437,N_26282,N_25453);
nor U26438 (N_26438,N_25612,N_25328);
nor U26439 (N_26439,N_25538,N_25438);
or U26440 (N_26440,N_26249,N_25784);
nand U26441 (N_26441,N_25840,N_25398);
nand U26442 (N_26442,N_25270,N_25734);
nand U26443 (N_26443,N_25735,N_25536);
or U26444 (N_26444,N_25496,N_25686);
or U26445 (N_26445,N_25363,N_26012);
xor U26446 (N_26446,N_26335,N_26350);
nor U26447 (N_26447,N_25448,N_25556);
nor U26448 (N_26448,N_25700,N_25597);
nor U26449 (N_26449,N_26055,N_26078);
xor U26450 (N_26450,N_25268,N_26311);
and U26451 (N_26451,N_25927,N_26167);
xor U26452 (N_26452,N_25300,N_25367);
or U26453 (N_26453,N_25318,N_26255);
nand U26454 (N_26454,N_25582,N_26058);
and U26455 (N_26455,N_25744,N_26155);
xnor U26456 (N_26456,N_26220,N_25365);
nand U26457 (N_26457,N_25263,N_26076);
and U26458 (N_26458,N_25392,N_25447);
or U26459 (N_26459,N_26008,N_25323);
or U26460 (N_26460,N_25381,N_26238);
xor U26461 (N_26461,N_25939,N_25911);
xor U26462 (N_26462,N_26139,N_25917);
nand U26463 (N_26463,N_26048,N_26169);
nor U26464 (N_26464,N_26140,N_25809);
nor U26465 (N_26465,N_26072,N_25736);
or U26466 (N_26466,N_25775,N_25748);
and U26467 (N_26467,N_25511,N_25599);
nor U26468 (N_26468,N_26132,N_25632);
or U26469 (N_26469,N_25433,N_26117);
nand U26470 (N_26470,N_25781,N_25440);
or U26471 (N_26471,N_25633,N_25965);
and U26472 (N_26472,N_25431,N_25636);
xor U26473 (N_26473,N_25685,N_25845);
or U26474 (N_26474,N_26198,N_26188);
nor U26475 (N_26475,N_25993,N_25446);
nand U26476 (N_26476,N_25335,N_25578);
xnor U26477 (N_26477,N_25655,N_26297);
nor U26478 (N_26478,N_26083,N_25576);
nor U26479 (N_26479,N_25491,N_25292);
and U26480 (N_26480,N_25929,N_25925);
nand U26481 (N_26481,N_25656,N_26223);
or U26482 (N_26482,N_25979,N_25371);
xnor U26483 (N_26483,N_25240,N_25315);
xnor U26484 (N_26484,N_26340,N_25805);
or U26485 (N_26485,N_25624,N_26288);
and U26486 (N_26486,N_25378,N_26396);
nor U26487 (N_26487,N_25435,N_25217);
nand U26488 (N_26488,N_26006,N_25853);
and U26489 (N_26489,N_25722,N_25705);
nor U26490 (N_26490,N_25520,N_26218);
xnor U26491 (N_26491,N_26214,N_25967);
nand U26492 (N_26492,N_25510,N_25940);
nor U26493 (N_26493,N_25557,N_26114);
or U26494 (N_26494,N_26266,N_25949);
and U26495 (N_26495,N_25806,N_25838);
nand U26496 (N_26496,N_26180,N_26034);
and U26497 (N_26497,N_25475,N_25513);
or U26498 (N_26498,N_26233,N_25420);
xor U26499 (N_26499,N_25721,N_25471);
or U26500 (N_26500,N_25824,N_26106);
xor U26501 (N_26501,N_26305,N_26073);
and U26502 (N_26502,N_26392,N_25972);
or U26503 (N_26503,N_26056,N_25203);
nor U26504 (N_26504,N_26370,N_25570);
and U26505 (N_26505,N_25974,N_25621);
nand U26506 (N_26506,N_25865,N_25290);
nand U26507 (N_26507,N_25259,N_26391);
nand U26508 (N_26508,N_25754,N_26261);
or U26509 (N_26509,N_25807,N_25373);
and U26510 (N_26510,N_25858,N_25753);
and U26511 (N_26511,N_25885,N_25479);
xor U26512 (N_26512,N_26315,N_25200);
and U26513 (N_26513,N_25878,N_25232);
nor U26514 (N_26514,N_26224,N_25567);
and U26515 (N_26515,N_26146,N_25695);
or U26516 (N_26516,N_26028,N_25630);
xnor U26517 (N_26517,N_26150,N_25568);
nand U26518 (N_26518,N_25924,N_26386);
and U26519 (N_26519,N_26361,N_25469);
or U26520 (N_26520,N_25985,N_25450);
nand U26521 (N_26521,N_26022,N_25830);
or U26522 (N_26522,N_25863,N_25666);
nor U26523 (N_26523,N_25711,N_25498);
nand U26524 (N_26524,N_26172,N_25620);
nor U26525 (N_26525,N_25522,N_26381);
nand U26526 (N_26526,N_26164,N_26328);
nand U26527 (N_26527,N_25826,N_25291);
xor U26528 (N_26528,N_25451,N_26161);
or U26529 (N_26529,N_25276,N_25280);
or U26530 (N_26530,N_25418,N_26339);
and U26531 (N_26531,N_26144,N_26069);
nand U26532 (N_26532,N_25740,N_26199);
xnor U26533 (N_26533,N_26079,N_25848);
nor U26534 (N_26534,N_26157,N_25909);
nor U26535 (N_26535,N_25768,N_25801);
or U26536 (N_26536,N_25364,N_25560);
nor U26537 (N_26537,N_25247,N_25688);
xnor U26538 (N_26538,N_26120,N_26124);
and U26539 (N_26539,N_25713,N_25530);
or U26540 (N_26540,N_25998,N_26088);
xor U26541 (N_26541,N_26082,N_26389);
and U26542 (N_26542,N_26211,N_25693);
xor U26543 (N_26543,N_25478,N_25641);
and U26544 (N_26544,N_25235,N_26057);
nor U26545 (N_26545,N_26229,N_25906);
and U26546 (N_26546,N_25728,N_25608);
nand U26547 (N_26547,N_26321,N_26152);
or U26548 (N_26548,N_25997,N_25609);
nand U26549 (N_26549,N_25773,N_25675);
nor U26550 (N_26550,N_26045,N_25847);
and U26551 (N_26551,N_25304,N_25355);
or U26552 (N_26552,N_25370,N_26221);
xor U26553 (N_26553,N_25674,N_25654);
and U26554 (N_26554,N_26026,N_25209);
and U26555 (N_26555,N_26018,N_26253);
xor U26556 (N_26556,N_25910,N_26175);
nor U26557 (N_26557,N_26235,N_25629);
and U26558 (N_26558,N_25254,N_25938);
nand U26559 (N_26559,N_25220,N_25887);
xor U26560 (N_26560,N_25725,N_25540);
or U26561 (N_26561,N_25233,N_25466);
nand U26562 (N_26562,N_25851,N_25248);
nand U26563 (N_26563,N_26177,N_25782);
nor U26564 (N_26564,N_26208,N_26382);
xnor U26565 (N_26565,N_26101,N_26259);
and U26566 (N_26566,N_25698,N_26103);
and U26567 (N_26567,N_26104,N_25750);
xnor U26568 (N_26568,N_25996,N_26168);
nand U26569 (N_26569,N_26000,N_25841);
nor U26570 (N_26570,N_26325,N_25461);
xnor U26571 (N_26571,N_25661,N_26216);
nand U26572 (N_26572,N_25944,N_25360);
nor U26573 (N_26573,N_25712,N_26064);
or U26574 (N_26574,N_25341,N_26279);
xnor U26575 (N_26575,N_25211,N_25747);
nor U26576 (N_26576,N_26228,N_25542);
xnor U26577 (N_26577,N_25422,N_25720);
nand U26578 (N_26578,N_25553,N_25262);
xnor U26579 (N_26579,N_25600,N_25517);
nor U26580 (N_26580,N_25663,N_25879);
and U26581 (N_26581,N_25201,N_25755);
xor U26582 (N_26582,N_25294,N_25610);
or U26583 (N_26583,N_25970,N_25273);
nand U26584 (N_26584,N_25514,N_25385);
xor U26585 (N_26585,N_25386,N_26243);
or U26586 (N_26586,N_25896,N_26096);
xor U26587 (N_26587,N_25758,N_25257);
nand U26588 (N_26588,N_25877,N_25357);
xor U26589 (N_26589,N_26384,N_26318);
xnor U26590 (N_26590,N_26052,N_25884);
xor U26591 (N_26591,N_25669,N_25359);
and U26592 (N_26592,N_25615,N_25842);
nand U26593 (N_26593,N_25593,N_26272);
nor U26594 (N_26594,N_25963,N_26066);
nor U26595 (N_26595,N_25855,N_26360);
or U26596 (N_26596,N_25481,N_25810);
and U26597 (N_26597,N_25908,N_25554);
xor U26598 (N_26598,N_25774,N_25445);
nand U26599 (N_26599,N_25856,N_25777);
xnor U26600 (N_26600,N_26252,N_26383);
nor U26601 (N_26601,N_26262,N_26369);
xnor U26602 (N_26602,N_25933,N_25690);
xor U26603 (N_26603,N_26201,N_26239);
or U26604 (N_26604,N_25250,N_25509);
xnor U26605 (N_26605,N_26271,N_25353);
nand U26606 (N_26606,N_25739,N_25527);
or U26607 (N_26607,N_25326,N_25617);
and U26608 (N_26608,N_25697,N_25822);
or U26609 (N_26609,N_25799,N_25213);
and U26610 (N_26610,N_26142,N_25427);
and U26611 (N_26611,N_25699,N_25715);
xor U26612 (N_26612,N_26317,N_25891);
nand U26613 (N_26613,N_25763,N_26075);
xor U26614 (N_26614,N_25658,N_25339);
nor U26615 (N_26615,N_25868,N_25260);
nand U26616 (N_26616,N_25229,N_26038);
and U26617 (N_26617,N_26290,N_26246);
xnor U26618 (N_26618,N_25231,N_25245);
xor U26619 (N_26619,N_25831,N_25265);
nand U26620 (N_26620,N_25467,N_25936);
nor U26621 (N_26621,N_25237,N_25572);
nor U26622 (N_26622,N_26387,N_25415);
or U26623 (N_26623,N_26306,N_26368);
nor U26624 (N_26624,N_26293,N_26092);
or U26625 (N_26625,N_26373,N_25652);
xnor U26626 (N_26626,N_26226,N_25534);
xor U26627 (N_26627,N_25459,N_25569);
or U26628 (N_26628,N_25913,N_25616);
or U26629 (N_26629,N_25827,N_26270);
xnor U26630 (N_26630,N_25407,N_26195);
nor U26631 (N_26631,N_26053,N_25350);
xnor U26632 (N_26632,N_25874,N_26123);
nor U26633 (N_26633,N_25295,N_25508);
or U26634 (N_26634,N_26100,N_26397);
nand U26635 (N_26635,N_26021,N_25872);
nor U26636 (N_26636,N_26244,N_25990);
nand U26637 (N_26637,N_26268,N_26047);
xnor U26638 (N_26638,N_26042,N_25314);
or U26639 (N_26639,N_25577,N_25639);
xor U26640 (N_26640,N_26080,N_25396);
or U26641 (N_26641,N_25436,N_25892);
or U26642 (N_26642,N_26388,N_25764);
nand U26643 (N_26643,N_25428,N_25210);
and U26644 (N_26644,N_26269,N_25474);
xor U26645 (N_26645,N_26217,N_25258);
or U26646 (N_26646,N_26213,N_25980);
nor U26647 (N_26647,N_25829,N_25531);
xor U26648 (N_26648,N_26125,N_25626);
nor U26649 (N_26649,N_26116,N_26085);
xnor U26650 (N_26650,N_25643,N_26171);
and U26651 (N_26651,N_25494,N_26099);
nor U26652 (N_26652,N_26181,N_26015);
and U26653 (N_26653,N_26044,N_26046);
or U26654 (N_26654,N_25999,N_26062);
nor U26655 (N_26655,N_26179,N_25802);
and U26656 (N_26656,N_25293,N_25760);
and U26657 (N_26657,N_25953,N_26019);
xnor U26658 (N_26658,N_26153,N_26093);
and U26659 (N_26659,N_25717,N_26359);
and U26660 (N_26660,N_26063,N_26254);
nand U26661 (N_26661,N_25490,N_25969);
nor U26662 (N_26662,N_26385,N_25562);
xnor U26663 (N_26663,N_25545,N_25454);
nand U26664 (N_26664,N_25272,N_25316);
nor U26665 (N_26665,N_25342,N_25579);
and U26666 (N_26666,N_25589,N_26394);
nor U26667 (N_26667,N_26010,N_25285);
or U26668 (N_26668,N_25628,N_25791);
nor U26669 (N_26669,N_26294,N_26310);
or U26670 (N_26670,N_25216,N_26009);
and U26671 (N_26671,N_26260,N_26128);
xor U26672 (N_26672,N_25945,N_25382);
xor U26673 (N_26673,N_25895,N_26237);
xor U26674 (N_26674,N_25372,N_26030);
xor U26675 (N_26675,N_25236,N_25707);
xor U26676 (N_26676,N_26206,N_25411);
nand U26677 (N_26677,N_25279,N_25312);
nand U26678 (N_26678,N_25903,N_26300);
or U26679 (N_26679,N_26241,N_26267);
and U26680 (N_26680,N_26283,N_25389);
or U26681 (N_26681,N_25348,N_25253);
nor U26682 (N_26682,N_25470,N_25587);
and U26683 (N_26683,N_25866,N_25737);
nor U26684 (N_26684,N_25741,N_25611);
nand U26685 (N_26685,N_25890,N_25871);
or U26686 (N_26686,N_25835,N_25330);
xnor U26687 (N_26687,N_25591,N_26133);
xor U26688 (N_26688,N_25779,N_26035);
and U26689 (N_26689,N_25369,N_26251);
xnor U26690 (N_26690,N_25846,N_25504);
xor U26691 (N_26691,N_25391,N_26326);
or U26692 (N_26692,N_25535,N_26059);
or U26693 (N_26693,N_25329,N_25573);
and U26694 (N_26694,N_25930,N_25477);
nand U26695 (N_26695,N_25942,N_26286);
and U26696 (N_26696,N_26135,N_25524);
and U26697 (N_26697,N_25225,N_25923);
nand U26698 (N_26698,N_25640,N_25813);
nor U26699 (N_26699,N_25772,N_26129);
nand U26700 (N_26700,N_25307,N_25823);
and U26701 (N_26701,N_25586,N_25442);
or U26702 (N_26702,N_25687,N_26192);
xnor U26703 (N_26703,N_25425,N_25397);
nor U26704 (N_26704,N_26051,N_25409);
nand U26705 (N_26705,N_26024,N_26145);
or U26706 (N_26706,N_25836,N_25563);
nand U26707 (N_26707,N_26004,N_25959);
or U26708 (N_26708,N_25837,N_26166);
and U26709 (N_26709,N_26302,N_25602);
or U26710 (N_26710,N_25850,N_26067);
or U26711 (N_26711,N_25374,N_26111);
or U26712 (N_26712,N_26277,N_25673);
nor U26713 (N_26713,N_26027,N_26336);
or U26714 (N_26714,N_25812,N_25521);
or U26715 (N_26715,N_26301,N_26138);
nand U26716 (N_26716,N_26207,N_26303);
or U26717 (N_26717,N_26143,N_26095);
nand U26718 (N_26718,N_25310,N_25532);
nor U26719 (N_26719,N_25671,N_25710);
nand U26720 (N_26720,N_25893,N_26122);
xor U26721 (N_26721,N_26250,N_26355);
and U26722 (N_26722,N_26020,N_25219);
nor U26723 (N_26723,N_25682,N_25468);
and U26724 (N_26724,N_26256,N_25894);
and U26725 (N_26725,N_25981,N_26334);
and U26726 (N_26726,N_25653,N_25590);
or U26727 (N_26727,N_25218,N_26194);
nand U26728 (N_26728,N_25946,N_26347);
or U26729 (N_26729,N_26299,N_25790);
nand U26730 (N_26730,N_26173,N_25650);
or U26731 (N_26731,N_25583,N_26236);
or U26732 (N_26732,N_25649,N_26170);
and U26733 (N_26733,N_25302,N_25907);
xor U26734 (N_26734,N_25767,N_25828);
nand U26735 (N_26735,N_26324,N_26112);
nor U26736 (N_26736,N_26137,N_26222);
nor U26737 (N_26737,N_25769,N_25516);
nand U26738 (N_26738,N_26230,N_25708);
and U26739 (N_26739,N_25224,N_26314);
nand U26740 (N_26740,N_26304,N_26323);
xor U26741 (N_26741,N_26033,N_25539);
xnor U26742 (N_26742,N_25955,N_26219);
and U26743 (N_26743,N_25795,N_25487);
nand U26744 (N_26744,N_25269,N_25559);
or U26745 (N_26745,N_25306,N_25668);
nor U26746 (N_26746,N_25752,N_25241);
nor U26747 (N_26747,N_26023,N_25915);
nor U26748 (N_26748,N_25502,N_26165);
and U26749 (N_26749,N_25512,N_26362);
and U26750 (N_26750,N_26182,N_25659);
nand U26751 (N_26751,N_26071,N_26127);
xor U26752 (N_26752,N_25920,N_26320);
nor U26753 (N_26753,N_25883,N_25485);
nand U26754 (N_26754,N_26276,N_25765);
nor U26755 (N_26755,N_25948,N_25506);
and U26756 (N_26756,N_26327,N_25983);
and U26757 (N_26757,N_26365,N_25401);
and U26758 (N_26758,N_26105,N_26005);
xor U26759 (N_26759,N_25277,N_26065);
xnor U26760 (N_26760,N_25648,N_26037);
and U26761 (N_26761,N_25480,N_25308);
and U26762 (N_26762,N_25443,N_25215);
or U26763 (N_26763,N_26089,N_26390);
nand U26764 (N_26764,N_25995,N_25950);
or U26765 (N_26765,N_25657,N_26154);
nor U26766 (N_26766,N_25961,N_25800);
nand U26767 (N_26767,N_25332,N_25388);
nand U26768 (N_26768,N_25821,N_26285);
or U26769 (N_26769,N_26247,N_26274);
nor U26770 (N_26770,N_25361,N_25456);
nand U26771 (N_26771,N_25482,N_26108);
nand U26772 (N_26772,N_25281,N_25598);
nor U26773 (N_26773,N_25358,N_26013);
and U26774 (N_26774,N_25709,N_25882);
or U26775 (N_26775,N_25356,N_25226);
or U26776 (N_26776,N_25619,N_25749);
nand U26777 (N_26777,N_26159,N_26398);
and U26778 (N_26778,N_25202,N_26148);
nor U26779 (N_26779,N_26395,N_25499);
xor U26780 (N_26780,N_25421,N_25457);
and U26781 (N_26781,N_26002,N_25472);
nand U26782 (N_26782,N_25566,N_26131);
or U26783 (N_26783,N_26187,N_26352);
xnor U26784 (N_26784,N_25704,N_25444);
nor U26785 (N_26785,N_25904,N_25726);
and U26786 (N_26786,N_26049,N_25819);
nor U26787 (N_26787,N_25796,N_26014);
nor U26788 (N_26788,N_25564,N_25525);
nand U26789 (N_26789,N_26094,N_25664);
nor U26790 (N_26790,N_25452,N_25834);
or U26791 (N_26791,N_25958,N_25375);
nand U26792 (N_26792,N_25251,N_25596);
xor U26793 (N_26793,N_26086,N_25701);
or U26794 (N_26794,N_25941,N_25622);
and U26795 (N_26795,N_25537,N_25860);
nand U26796 (N_26796,N_25503,N_25413);
xor U26797 (N_26797,N_25761,N_25234);
or U26798 (N_26798,N_25681,N_25793);
nor U26799 (N_26799,N_26158,N_25975);
and U26800 (N_26800,N_25337,N_25244);
and U26801 (N_26801,N_26003,N_26231);
or U26802 (N_26802,N_25393,N_25249);
xnor U26803 (N_26803,N_25683,N_26097);
or U26804 (N_26804,N_25808,N_26227);
nor U26805 (N_26805,N_25432,N_25703);
or U26806 (N_26806,N_25286,N_25261);
and U26807 (N_26807,N_26313,N_26130);
or U26808 (N_26808,N_25968,N_25301);
or U26809 (N_26809,N_25205,N_25212);
or U26810 (N_26810,N_25787,N_25297);
nand U26811 (N_26811,N_26178,N_25719);
nor U26812 (N_26812,N_25552,N_25943);
xor U26813 (N_26813,N_25575,N_25679);
and U26814 (N_26814,N_26087,N_25419);
nor U26815 (N_26815,N_26205,N_25298);
and U26816 (N_26816,N_25325,N_25994);
xnor U26817 (N_26817,N_26376,N_25914);
nor U26818 (N_26818,N_25880,N_25327);
or U26819 (N_26819,N_26265,N_26189);
or U26820 (N_26820,N_25778,N_25922);
nand U26821 (N_26821,N_26309,N_26344);
nor U26822 (N_26822,N_25439,N_25476);
xor U26823 (N_26823,N_26121,N_25642);
or U26824 (N_26824,N_25287,N_25405);
and U26825 (N_26825,N_26281,N_26364);
xor U26826 (N_26826,N_25299,N_25746);
nand U26827 (N_26827,N_26134,N_25935);
nor U26828 (N_26828,N_25776,N_25757);
nand U26829 (N_26829,N_25515,N_26163);
and U26830 (N_26830,N_25956,N_25347);
and U26831 (N_26831,N_25584,N_25222);
and U26832 (N_26832,N_25604,N_25900);
nand U26833 (N_26833,N_25870,N_25242);
nor U26834 (N_26834,N_25954,N_25646);
and U26835 (N_26835,N_25346,N_26354);
xor U26836 (N_26836,N_25377,N_25987);
and U26837 (N_26837,N_25984,N_26204);
xor U26838 (N_26838,N_25864,N_25798);
and U26839 (N_26839,N_25797,N_25960);
or U26840 (N_26840,N_26341,N_25338);
xnor U26841 (N_26841,N_25458,N_25271);
xor U26842 (N_26842,N_25672,N_25501);
nor U26843 (N_26843,N_25283,N_25434);
nor U26844 (N_26844,N_26295,N_26337);
nor U26845 (N_26845,N_25354,N_25651);
nand U26846 (N_26846,N_25558,N_25256);
xor U26847 (N_26847,N_25976,N_25403);
or U26848 (N_26848,N_25873,N_26183);
and U26849 (N_26849,N_26308,N_25859);
nor U26850 (N_26850,N_26007,N_25843);
nor U26851 (N_26851,N_25465,N_25488);
xnor U26852 (N_26852,N_26393,N_25833);
nor U26853 (N_26853,N_26115,N_26060);
or U26854 (N_26854,N_25966,N_25518);
or U26855 (N_26855,N_25264,N_25282);
nand U26856 (N_26856,N_25815,N_26215);
nand U26857 (N_26857,N_25336,N_26242);
and U26858 (N_26858,N_26054,N_25786);
xnor U26859 (N_26859,N_26280,N_25410);
and U26860 (N_26860,N_26356,N_25691);
nand U26861 (N_26861,N_26070,N_25585);
or U26862 (N_26862,N_25533,N_25881);
or U26863 (N_26863,N_25901,N_25647);
or U26864 (N_26864,N_25952,N_26333);
nand U26865 (N_26865,N_25771,N_25541);
nand U26866 (N_26866,N_25716,N_25252);
or U26867 (N_26867,N_25345,N_25888);
nand U26868 (N_26868,N_25402,N_25255);
nand U26869 (N_26869,N_25449,N_26162);
xor U26870 (N_26870,N_25423,N_25207);
nand U26871 (N_26871,N_25644,N_25912);
xor U26872 (N_26872,N_26191,N_25319);
and U26873 (N_26873,N_26351,N_25519);
or U26874 (N_26874,N_25404,N_26081);
nand U26875 (N_26875,N_26263,N_26380);
xnor U26876 (N_26876,N_26210,N_25275);
or U26877 (N_26877,N_26346,N_26061);
nand U26878 (N_26878,N_25978,N_26050);
or U26879 (N_26879,N_26074,N_25662);
and U26880 (N_26880,N_25852,N_25804);
or U26881 (N_26881,N_26378,N_25592);
xor U26882 (N_26882,N_25614,N_26185);
or U26883 (N_26883,N_26156,N_25788);
or U26884 (N_26884,N_25594,N_25794);
and U26885 (N_26885,N_25351,N_25817);
xnor U26886 (N_26886,N_25732,N_26374);
or U26887 (N_26887,N_25574,N_25320);
nor U26888 (N_26888,N_26017,N_25333);
or U26889 (N_26889,N_26245,N_25899);
and U26890 (N_26890,N_25544,N_25937);
and U26891 (N_26891,N_25266,N_25785);
and U26892 (N_26892,N_25696,N_26041);
or U26893 (N_26893,N_25962,N_25947);
and U26894 (N_26894,N_26032,N_25762);
xor U26895 (N_26895,N_25239,N_25745);
and U26896 (N_26896,N_25529,N_25660);
xor U26897 (N_26897,N_25221,N_25605);
or U26898 (N_26898,N_26264,N_26043);
or U26899 (N_26899,N_25208,N_26367);
nand U26900 (N_26900,N_25417,N_25400);
nor U26901 (N_26901,N_26296,N_25818);
nand U26902 (N_26902,N_25463,N_25565);
and U26903 (N_26903,N_25625,N_25635);
and U26904 (N_26904,N_25898,N_25379);
nand U26905 (N_26905,N_25742,N_26141);
nor U26906 (N_26906,N_25344,N_25349);
nand U26907 (N_26907,N_26307,N_26225);
xnor U26908 (N_26908,N_25844,N_25547);
or U26909 (N_26909,N_25803,N_25414);
nand U26910 (N_26910,N_25340,N_25733);
nand U26911 (N_26911,N_26371,N_26349);
and U26912 (N_26912,N_25770,N_25977);
nor U26913 (N_26913,N_25814,N_25738);
or U26914 (N_26914,N_25507,N_26113);
xor U26915 (N_26915,N_25551,N_25429);
and U26916 (N_26916,N_26149,N_25206);
and U26917 (N_26917,N_25549,N_26039);
xnor U26918 (N_26918,N_26036,N_25982);
nand U26919 (N_26919,N_25718,N_25406);
nor U26920 (N_26920,N_26278,N_25613);
or U26921 (N_26921,N_25523,N_25238);
and U26922 (N_26922,N_25816,N_25706);
nand U26923 (N_26923,N_25867,N_25426);
xnor U26924 (N_26924,N_25486,N_25305);
nor U26925 (N_26925,N_25905,N_25500);
nor U26926 (N_26926,N_26190,N_25832);
nand U26927 (N_26927,N_25684,N_25623);
nor U26928 (N_26928,N_26068,N_25714);
and U26929 (N_26929,N_25861,N_25702);
nor U26930 (N_26930,N_25505,N_26209);
or U26931 (N_26931,N_26202,N_25603);
xnor U26932 (N_26932,N_26176,N_25957);
nor U26933 (N_26933,N_25267,N_25986);
or U26934 (N_26934,N_26107,N_25869);
nand U26935 (N_26935,N_25384,N_25366);
or U26936 (N_26936,N_26196,N_26329);
xor U26937 (N_26937,N_25932,N_25464);
or U26938 (N_26938,N_26109,N_26343);
or U26939 (N_26939,N_25689,N_25897);
nor U26940 (N_26940,N_26084,N_26160);
or U26941 (N_26941,N_25631,N_25455);
nand U26942 (N_26942,N_25492,N_25571);
xnor U26943 (N_26943,N_25849,N_25606);
xor U26944 (N_26944,N_26011,N_25204);
and U26945 (N_26945,N_25424,N_26379);
or U26946 (N_26946,N_26316,N_25303);
xnor U26947 (N_26947,N_26319,N_25916);
and U26948 (N_26948,N_25412,N_25462);
nand U26949 (N_26949,N_26331,N_25588);
and U26950 (N_26950,N_25634,N_26342);
nor U26951 (N_26951,N_25580,N_25437);
nand U26952 (N_26952,N_25926,N_25991);
and U26953 (N_26953,N_26358,N_25352);
nand U26954 (N_26954,N_25546,N_25278);
nor U26955 (N_26955,N_25992,N_26197);
or U26956 (N_26956,N_25789,N_26248);
or U26957 (N_26957,N_26203,N_25751);
nand U26958 (N_26958,N_25483,N_26184);
or U26959 (N_26959,N_26287,N_26232);
nor U26960 (N_26960,N_25902,N_26212);
and U26961 (N_26961,N_26330,N_25665);
or U26962 (N_26962,N_25324,N_25289);
and U26963 (N_26963,N_25230,N_25724);
and U26964 (N_26964,N_25595,N_25284);
or U26965 (N_26965,N_26275,N_25973);
or U26966 (N_26966,N_26292,N_26136);
and U26967 (N_26967,N_25676,N_25989);
and U26968 (N_26968,N_25638,N_25317);
and U26969 (N_26969,N_25561,N_25543);
nor U26970 (N_26970,N_25296,N_26357);
nor U26971 (N_26971,N_25416,N_25555);
and U26972 (N_26972,N_25727,N_25214);
nor U26973 (N_26973,N_26193,N_25857);
or U26974 (N_26974,N_26016,N_26090);
or U26975 (N_26975,N_25839,N_25484);
nand U26976 (N_26976,N_26312,N_26102);
nor U26977 (N_26977,N_25759,N_25362);
nand U26978 (N_26978,N_25677,N_26118);
or U26979 (N_26979,N_25526,N_25928);
nor U26980 (N_26980,N_25227,N_26298);
and U26981 (N_26981,N_25670,N_25694);
xnor U26982 (N_26982,N_25692,N_25550);
and U26983 (N_26983,N_26257,N_25645);
nor U26984 (N_26984,N_25288,N_25618);
or U26985 (N_26985,N_26077,N_26375);
or U26986 (N_26986,N_25886,N_25394);
and U26987 (N_26987,N_25528,N_26126);
xor U26988 (N_26988,N_25395,N_26363);
and U26989 (N_26989,N_25951,N_26119);
and U26990 (N_26990,N_25309,N_25383);
and U26991 (N_26991,N_26040,N_25731);
xnor U26992 (N_26992,N_26345,N_26291);
or U26993 (N_26993,N_25601,N_26258);
xor U26994 (N_26994,N_26234,N_25820);
or U26995 (N_26995,N_25607,N_25243);
xor U26996 (N_26996,N_26031,N_26399);
and U26997 (N_26997,N_26186,N_26353);
xor U26998 (N_26998,N_25811,N_25460);
xor U26999 (N_26999,N_25889,N_25988);
nor U27000 (N_27000,N_25769,N_25340);
or U27001 (N_27001,N_25654,N_25839);
nand U27002 (N_27002,N_25856,N_25302);
and U27003 (N_27003,N_26371,N_25914);
or U27004 (N_27004,N_26196,N_26200);
or U27005 (N_27005,N_25204,N_26046);
nor U27006 (N_27006,N_26046,N_25829);
nor U27007 (N_27007,N_26063,N_25304);
and U27008 (N_27008,N_25778,N_25689);
or U27009 (N_27009,N_25243,N_26336);
xnor U27010 (N_27010,N_26191,N_25407);
nand U27011 (N_27011,N_25875,N_25405);
nor U27012 (N_27012,N_26089,N_26331);
xnor U27013 (N_27013,N_25894,N_25621);
and U27014 (N_27014,N_25295,N_25621);
nand U27015 (N_27015,N_25793,N_26371);
nand U27016 (N_27016,N_26140,N_25921);
nand U27017 (N_27017,N_26055,N_25602);
nor U27018 (N_27018,N_25583,N_25732);
nand U27019 (N_27019,N_25259,N_26309);
or U27020 (N_27020,N_25470,N_25969);
or U27021 (N_27021,N_26310,N_25416);
nor U27022 (N_27022,N_26362,N_25290);
xor U27023 (N_27023,N_25745,N_25223);
nor U27024 (N_27024,N_26330,N_25421);
nand U27025 (N_27025,N_25739,N_25310);
nor U27026 (N_27026,N_25903,N_26326);
and U27027 (N_27027,N_25542,N_26276);
nand U27028 (N_27028,N_26192,N_25488);
xnor U27029 (N_27029,N_25568,N_25267);
xnor U27030 (N_27030,N_25987,N_26147);
xor U27031 (N_27031,N_26379,N_25789);
and U27032 (N_27032,N_25642,N_25775);
nand U27033 (N_27033,N_25885,N_25658);
nor U27034 (N_27034,N_25493,N_25750);
and U27035 (N_27035,N_26388,N_25873);
and U27036 (N_27036,N_25940,N_25362);
or U27037 (N_27037,N_25213,N_26166);
nor U27038 (N_27038,N_26340,N_25440);
nor U27039 (N_27039,N_25324,N_25789);
nand U27040 (N_27040,N_25747,N_26340);
or U27041 (N_27041,N_25484,N_25314);
nor U27042 (N_27042,N_25669,N_26102);
nand U27043 (N_27043,N_26358,N_25233);
or U27044 (N_27044,N_26151,N_26176);
and U27045 (N_27045,N_25236,N_25552);
nor U27046 (N_27046,N_25825,N_25393);
nor U27047 (N_27047,N_26120,N_26321);
nand U27048 (N_27048,N_25869,N_25933);
nor U27049 (N_27049,N_26049,N_25477);
xnor U27050 (N_27050,N_25736,N_26157);
nor U27051 (N_27051,N_25475,N_25701);
nand U27052 (N_27052,N_25941,N_25384);
and U27053 (N_27053,N_25968,N_25738);
xor U27054 (N_27054,N_25876,N_25654);
nor U27055 (N_27055,N_25646,N_26257);
and U27056 (N_27056,N_25582,N_25888);
nand U27057 (N_27057,N_25801,N_25649);
and U27058 (N_27058,N_25769,N_25309);
nor U27059 (N_27059,N_26376,N_25416);
nand U27060 (N_27060,N_26259,N_25230);
nand U27061 (N_27061,N_26086,N_26254);
xor U27062 (N_27062,N_25711,N_26249);
nor U27063 (N_27063,N_25805,N_26062);
nand U27064 (N_27064,N_26304,N_26277);
or U27065 (N_27065,N_25360,N_25322);
xnor U27066 (N_27066,N_25629,N_25814);
nand U27067 (N_27067,N_25827,N_26043);
nand U27068 (N_27068,N_25504,N_25854);
or U27069 (N_27069,N_25376,N_26298);
xnor U27070 (N_27070,N_25416,N_25418);
nand U27071 (N_27071,N_25621,N_25294);
and U27072 (N_27072,N_25930,N_25245);
or U27073 (N_27073,N_25387,N_26056);
or U27074 (N_27074,N_25337,N_26365);
xor U27075 (N_27075,N_26081,N_25987);
xnor U27076 (N_27076,N_26173,N_25989);
or U27077 (N_27077,N_26322,N_25906);
nand U27078 (N_27078,N_25613,N_25345);
or U27079 (N_27079,N_25398,N_26264);
nor U27080 (N_27080,N_25236,N_26041);
nor U27081 (N_27081,N_25509,N_25501);
xor U27082 (N_27082,N_25493,N_25628);
or U27083 (N_27083,N_25938,N_25350);
and U27084 (N_27084,N_25933,N_26202);
nor U27085 (N_27085,N_25513,N_26015);
and U27086 (N_27086,N_26055,N_25252);
xor U27087 (N_27087,N_25895,N_26025);
xnor U27088 (N_27088,N_25600,N_25389);
nor U27089 (N_27089,N_25566,N_25311);
and U27090 (N_27090,N_25524,N_25212);
or U27091 (N_27091,N_25983,N_25383);
and U27092 (N_27092,N_25772,N_25524);
nand U27093 (N_27093,N_25407,N_25926);
xnor U27094 (N_27094,N_25661,N_25858);
xor U27095 (N_27095,N_25768,N_26029);
xor U27096 (N_27096,N_25251,N_25479);
or U27097 (N_27097,N_25839,N_25709);
nor U27098 (N_27098,N_26133,N_26074);
xnor U27099 (N_27099,N_25543,N_26134);
xnor U27100 (N_27100,N_25224,N_25738);
or U27101 (N_27101,N_25500,N_25339);
nor U27102 (N_27102,N_26221,N_26025);
nand U27103 (N_27103,N_25451,N_25621);
xor U27104 (N_27104,N_26094,N_26280);
or U27105 (N_27105,N_26316,N_26128);
xnor U27106 (N_27106,N_25618,N_25423);
or U27107 (N_27107,N_25324,N_25902);
or U27108 (N_27108,N_26296,N_26366);
nand U27109 (N_27109,N_26300,N_26293);
and U27110 (N_27110,N_26167,N_25602);
or U27111 (N_27111,N_25779,N_25528);
nand U27112 (N_27112,N_26333,N_25403);
nand U27113 (N_27113,N_26142,N_25422);
or U27114 (N_27114,N_26343,N_26121);
nand U27115 (N_27115,N_25209,N_26171);
and U27116 (N_27116,N_26178,N_25797);
or U27117 (N_27117,N_26025,N_26227);
and U27118 (N_27118,N_25991,N_25230);
xor U27119 (N_27119,N_25808,N_25771);
and U27120 (N_27120,N_25348,N_25206);
and U27121 (N_27121,N_26166,N_25231);
or U27122 (N_27122,N_26356,N_25279);
xor U27123 (N_27123,N_26379,N_25276);
xor U27124 (N_27124,N_25373,N_25530);
nand U27125 (N_27125,N_26215,N_25943);
or U27126 (N_27126,N_25781,N_25478);
nor U27127 (N_27127,N_26019,N_25201);
and U27128 (N_27128,N_25296,N_25758);
xor U27129 (N_27129,N_25214,N_26094);
nor U27130 (N_27130,N_26284,N_25663);
and U27131 (N_27131,N_25473,N_25905);
xnor U27132 (N_27132,N_25214,N_25280);
nand U27133 (N_27133,N_25824,N_26210);
and U27134 (N_27134,N_25564,N_25844);
nand U27135 (N_27135,N_25420,N_25825);
nand U27136 (N_27136,N_25583,N_26215);
nor U27137 (N_27137,N_25636,N_25510);
and U27138 (N_27138,N_25427,N_26261);
nand U27139 (N_27139,N_25882,N_25584);
and U27140 (N_27140,N_25552,N_26066);
nor U27141 (N_27141,N_25315,N_26287);
xnor U27142 (N_27142,N_25879,N_25824);
xnor U27143 (N_27143,N_25410,N_25790);
xor U27144 (N_27144,N_25632,N_26015);
xnor U27145 (N_27145,N_26326,N_26053);
xnor U27146 (N_27146,N_25955,N_25621);
or U27147 (N_27147,N_26135,N_26366);
nor U27148 (N_27148,N_25554,N_25449);
nand U27149 (N_27149,N_25485,N_25204);
xnor U27150 (N_27150,N_25755,N_25536);
nand U27151 (N_27151,N_25427,N_26175);
nand U27152 (N_27152,N_26146,N_25364);
xnor U27153 (N_27153,N_25932,N_25754);
or U27154 (N_27154,N_26022,N_25927);
xor U27155 (N_27155,N_26115,N_25237);
xnor U27156 (N_27156,N_26175,N_26261);
nor U27157 (N_27157,N_25237,N_25302);
xnor U27158 (N_27158,N_25862,N_25603);
and U27159 (N_27159,N_25917,N_26379);
xnor U27160 (N_27160,N_26378,N_25530);
xor U27161 (N_27161,N_25759,N_25882);
xor U27162 (N_27162,N_26388,N_25561);
nand U27163 (N_27163,N_25843,N_25763);
nor U27164 (N_27164,N_25428,N_25751);
and U27165 (N_27165,N_26326,N_25548);
and U27166 (N_27166,N_26173,N_26295);
xnor U27167 (N_27167,N_26055,N_25376);
nor U27168 (N_27168,N_25668,N_26124);
nor U27169 (N_27169,N_25986,N_25215);
nand U27170 (N_27170,N_25832,N_25681);
or U27171 (N_27171,N_25307,N_25700);
nor U27172 (N_27172,N_25741,N_25239);
xor U27173 (N_27173,N_26302,N_25560);
nand U27174 (N_27174,N_25262,N_26361);
nor U27175 (N_27175,N_25894,N_26241);
and U27176 (N_27176,N_25646,N_25824);
or U27177 (N_27177,N_25787,N_25489);
or U27178 (N_27178,N_25734,N_26185);
or U27179 (N_27179,N_25296,N_26121);
nand U27180 (N_27180,N_25826,N_25380);
xor U27181 (N_27181,N_25685,N_26009);
nand U27182 (N_27182,N_25844,N_25744);
or U27183 (N_27183,N_25242,N_25438);
and U27184 (N_27184,N_25262,N_25479);
and U27185 (N_27185,N_26021,N_25567);
nor U27186 (N_27186,N_25974,N_25445);
xor U27187 (N_27187,N_26030,N_25917);
nand U27188 (N_27188,N_25304,N_25567);
or U27189 (N_27189,N_26126,N_25442);
or U27190 (N_27190,N_25466,N_26185);
xnor U27191 (N_27191,N_26184,N_26063);
xnor U27192 (N_27192,N_26340,N_26394);
nand U27193 (N_27193,N_25939,N_25414);
or U27194 (N_27194,N_25880,N_25624);
xor U27195 (N_27195,N_25455,N_25530);
nor U27196 (N_27196,N_26365,N_26362);
and U27197 (N_27197,N_26266,N_26132);
xnor U27198 (N_27198,N_25834,N_26331);
nor U27199 (N_27199,N_25899,N_26371);
nor U27200 (N_27200,N_25855,N_25738);
xnor U27201 (N_27201,N_26350,N_25374);
nor U27202 (N_27202,N_25752,N_26393);
nand U27203 (N_27203,N_26160,N_26177);
nand U27204 (N_27204,N_26080,N_26249);
and U27205 (N_27205,N_26179,N_26320);
and U27206 (N_27206,N_26133,N_26008);
xnor U27207 (N_27207,N_25642,N_26146);
nor U27208 (N_27208,N_26255,N_25643);
nor U27209 (N_27209,N_25262,N_26091);
nor U27210 (N_27210,N_25958,N_25880);
xor U27211 (N_27211,N_25201,N_25968);
and U27212 (N_27212,N_25389,N_26282);
and U27213 (N_27213,N_26067,N_25961);
or U27214 (N_27214,N_25739,N_26023);
xor U27215 (N_27215,N_25702,N_25886);
and U27216 (N_27216,N_26095,N_25338);
or U27217 (N_27217,N_25406,N_25721);
nor U27218 (N_27218,N_26197,N_25878);
nand U27219 (N_27219,N_26229,N_25515);
or U27220 (N_27220,N_25411,N_25807);
and U27221 (N_27221,N_26177,N_25413);
and U27222 (N_27222,N_25269,N_26152);
and U27223 (N_27223,N_25527,N_25341);
and U27224 (N_27224,N_26176,N_25499);
nor U27225 (N_27225,N_26056,N_25399);
xnor U27226 (N_27226,N_25599,N_25636);
and U27227 (N_27227,N_26313,N_25669);
nor U27228 (N_27228,N_26048,N_25413);
xor U27229 (N_27229,N_25489,N_25432);
nand U27230 (N_27230,N_25932,N_25443);
xnor U27231 (N_27231,N_25517,N_26117);
and U27232 (N_27232,N_25212,N_25624);
nand U27233 (N_27233,N_25767,N_26190);
xor U27234 (N_27234,N_25281,N_25973);
xor U27235 (N_27235,N_26339,N_26210);
nand U27236 (N_27236,N_26173,N_25294);
nand U27237 (N_27237,N_25205,N_26226);
and U27238 (N_27238,N_25346,N_25893);
nor U27239 (N_27239,N_26327,N_25753);
and U27240 (N_27240,N_25987,N_25945);
nor U27241 (N_27241,N_25819,N_25775);
and U27242 (N_27242,N_25679,N_25762);
and U27243 (N_27243,N_25413,N_25494);
nand U27244 (N_27244,N_25527,N_26334);
xor U27245 (N_27245,N_25367,N_26194);
nand U27246 (N_27246,N_25650,N_26122);
and U27247 (N_27247,N_25595,N_26024);
nor U27248 (N_27248,N_25393,N_25391);
or U27249 (N_27249,N_25559,N_25983);
nor U27250 (N_27250,N_26161,N_25677);
and U27251 (N_27251,N_26338,N_26110);
or U27252 (N_27252,N_25635,N_25857);
nor U27253 (N_27253,N_25351,N_25837);
nor U27254 (N_27254,N_26106,N_25957);
or U27255 (N_27255,N_26137,N_25392);
nor U27256 (N_27256,N_25527,N_25311);
xor U27257 (N_27257,N_26048,N_26288);
nor U27258 (N_27258,N_25974,N_26065);
and U27259 (N_27259,N_25437,N_26021);
nand U27260 (N_27260,N_26250,N_25977);
or U27261 (N_27261,N_26126,N_25244);
nand U27262 (N_27262,N_25310,N_25737);
xor U27263 (N_27263,N_25610,N_25879);
xnor U27264 (N_27264,N_25758,N_25590);
nor U27265 (N_27265,N_25468,N_26370);
and U27266 (N_27266,N_26318,N_25808);
nor U27267 (N_27267,N_25204,N_25931);
xnor U27268 (N_27268,N_25878,N_25731);
and U27269 (N_27269,N_26388,N_25830);
nand U27270 (N_27270,N_26155,N_26125);
nor U27271 (N_27271,N_25966,N_26022);
nor U27272 (N_27272,N_25389,N_25331);
xor U27273 (N_27273,N_26237,N_25768);
nor U27274 (N_27274,N_25436,N_25353);
nor U27275 (N_27275,N_25709,N_25577);
nand U27276 (N_27276,N_25369,N_25400);
xor U27277 (N_27277,N_25506,N_25263);
nand U27278 (N_27278,N_26062,N_25532);
xnor U27279 (N_27279,N_26363,N_25955);
nand U27280 (N_27280,N_25257,N_25815);
nand U27281 (N_27281,N_25992,N_25311);
or U27282 (N_27282,N_25666,N_25970);
or U27283 (N_27283,N_26312,N_25346);
xor U27284 (N_27284,N_26293,N_25734);
and U27285 (N_27285,N_25592,N_26327);
nor U27286 (N_27286,N_25921,N_26344);
and U27287 (N_27287,N_25652,N_25829);
or U27288 (N_27288,N_25651,N_26186);
and U27289 (N_27289,N_25701,N_25638);
and U27290 (N_27290,N_26012,N_26117);
nand U27291 (N_27291,N_25561,N_25715);
or U27292 (N_27292,N_26278,N_25924);
or U27293 (N_27293,N_25758,N_25219);
and U27294 (N_27294,N_25670,N_25223);
xnor U27295 (N_27295,N_25967,N_26286);
nor U27296 (N_27296,N_26161,N_25816);
nor U27297 (N_27297,N_25351,N_25885);
xor U27298 (N_27298,N_26262,N_26236);
nand U27299 (N_27299,N_25201,N_26280);
or U27300 (N_27300,N_26281,N_25553);
xnor U27301 (N_27301,N_25365,N_26180);
nand U27302 (N_27302,N_25653,N_25487);
nand U27303 (N_27303,N_25506,N_25378);
nand U27304 (N_27304,N_25332,N_26012);
or U27305 (N_27305,N_26138,N_26126);
xnor U27306 (N_27306,N_25473,N_26367);
or U27307 (N_27307,N_26352,N_25343);
and U27308 (N_27308,N_25720,N_25514);
nor U27309 (N_27309,N_25479,N_25600);
xor U27310 (N_27310,N_25262,N_25647);
xnor U27311 (N_27311,N_26162,N_25271);
or U27312 (N_27312,N_25298,N_26034);
nand U27313 (N_27313,N_26214,N_25279);
nand U27314 (N_27314,N_26078,N_25420);
xor U27315 (N_27315,N_25759,N_25781);
or U27316 (N_27316,N_25560,N_25643);
nand U27317 (N_27317,N_25553,N_26060);
nor U27318 (N_27318,N_25388,N_25561);
and U27319 (N_27319,N_25479,N_25456);
nor U27320 (N_27320,N_25768,N_25453);
and U27321 (N_27321,N_25596,N_26168);
nor U27322 (N_27322,N_25849,N_25675);
xnor U27323 (N_27323,N_25948,N_26104);
nand U27324 (N_27324,N_25994,N_26155);
or U27325 (N_27325,N_25352,N_25950);
nor U27326 (N_27326,N_26123,N_25818);
xor U27327 (N_27327,N_25568,N_25805);
xnor U27328 (N_27328,N_26123,N_26135);
nor U27329 (N_27329,N_26212,N_25428);
or U27330 (N_27330,N_25271,N_26000);
nor U27331 (N_27331,N_26319,N_25659);
and U27332 (N_27332,N_25822,N_25878);
and U27333 (N_27333,N_25836,N_25300);
and U27334 (N_27334,N_26202,N_25610);
nor U27335 (N_27335,N_26225,N_25712);
or U27336 (N_27336,N_25461,N_25346);
xor U27337 (N_27337,N_25217,N_26351);
nand U27338 (N_27338,N_25525,N_25717);
or U27339 (N_27339,N_26181,N_25891);
and U27340 (N_27340,N_25993,N_25308);
nand U27341 (N_27341,N_26290,N_25621);
and U27342 (N_27342,N_26184,N_25562);
or U27343 (N_27343,N_25518,N_26121);
or U27344 (N_27344,N_25948,N_25244);
and U27345 (N_27345,N_25587,N_25630);
and U27346 (N_27346,N_26261,N_25362);
and U27347 (N_27347,N_26111,N_25902);
nand U27348 (N_27348,N_25760,N_25217);
nand U27349 (N_27349,N_25844,N_26066);
xor U27350 (N_27350,N_25797,N_25599);
and U27351 (N_27351,N_25623,N_25759);
nor U27352 (N_27352,N_25714,N_25302);
and U27353 (N_27353,N_25483,N_26388);
xor U27354 (N_27354,N_25519,N_25545);
xnor U27355 (N_27355,N_25925,N_25264);
nor U27356 (N_27356,N_26346,N_26229);
xnor U27357 (N_27357,N_25578,N_25500);
or U27358 (N_27358,N_26071,N_25909);
xnor U27359 (N_27359,N_26027,N_26048);
or U27360 (N_27360,N_26139,N_26122);
nand U27361 (N_27361,N_25241,N_25975);
xnor U27362 (N_27362,N_26110,N_25458);
nand U27363 (N_27363,N_25887,N_26238);
and U27364 (N_27364,N_25245,N_26295);
nor U27365 (N_27365,N_25970,N_25688);
or U27366 (N_27366,N_25645,N_26245);
nor U27367 (N_27367,N_26061,N_25390);
nand U27368 (N_27368,N_25424,N_25466);
nand U27369 (N_27369,N_25349,N_26329);
nand U27370 (N_27370,N_25649,N_25273);
nand U27371 (N_27371,N_26212,N_26072);
nand U27372 (N_27372,N_25752,N_26234);
nor U27373 (N_27373,N_25336,N_26259);
or U27374 (N_27374,N_25975,N_26173);
nor U27375 (N_27375,N_25400,N_26322);
nand U27376 (N_27376,N_25491,N_26233);
xnor U27377 (N_27377,N_25489,N_25869);
and U27378 (N_27378,N_26349,N_25499);
nor U27379 (N_27379,N_25742,N_26021);
or U27380 (N_27380,N_25928,N_25650);
nor U27381 (N_27381,N_25745,N_25684);
xor U27382 (N_27382,N_25704,N_25903);
nand U27383 (N_27383,N_25909,N_25503);
xor U27384 (N_27384,N_25994,N_25827);
xnor U27385 (N_27385,N_26369,N_25880);
xor U27386 (N_27386,N_25833,N_25677);
and U27387 (N_27387,N_25643,N_25263);
nand U27388 (N_27388,N_25510,N_25607);
or U27389 (N_27389,N_26281,N_25930);
or U27390 (N_27390,N_25765,N_26362);
or U27391 (N_27391,N_26198,N_25648);
nor U27392 (N_27392,N_25665,N_26014);
and U27393 (N_27393,N_25341,N_25954);
xnor U27394 (N_27394,N_26339,N_26022);
xnor U27395 (N_27395,N_26141,N_26262);
or U27396 (N_27396,N_25328,N_25832);
or U27397 (N_27397,N_25740,N_25563);
or U27398 (N_27398,N_26131,N_26112);
and U27399 (N_27399,N_25916,N_26014);
nand U27400 (N_27400,N_26147,N_26103);
and U27401 (N_27401,N_25710,N_25691);
nand U27402 (N_27402,N_26012,N_26388);
or U27403 (N_27403,N_26205,N_25473);
nor U27404 (N_27404,N_26100,N_25487);
nor U27405 (N_27405,N_25334,N_26127);
nor U27406 (N_27406,N_25676,N_25340);
nand U27407 (N_27407,N_25993,N_25665);
nor U27408 (N_27408,N_25930,N_25683);
nor U27409 (N_27409,N_25328,N_25947);
xor U27410 (N_27410,N_25813,N_26394);
and U27411 (N_27411,N_25780,N_26385);
nand U27412 (N_27412,N_26328,N_25691);
nand U27413 (N_27413,N_26244,N_26073);
nor U27414 (N_27414,N_26333,N_25315);
or U27415 (N_27415,N_25733,N_25549);
and U27416 (N_27416,N_25483,N_25392);
and U27417 (N_27417,N_26068,N_25552);
nand U27418 (N_27418,N_25786,N_26045);
and U27419 (N_27419,N_25759,N_26368);
nand U27420 (N_27420,N_25242,N_26241);
nor U27421 (N_27421,N_25391,N_26392);
nand U27422 (N_27422,N_25238,N_25379);
nor U27423 (N_27423,N_25789,N_25862);
xnor U27424 (N_27424,N_25753,N_26185);
nand U27425 (N_27425,N_25253,N_26154);
nand U27426 (N_27426,N_25216,N_25595);
nand U27427 (N_27427,N_26384,N_26167);
and U27428 (N_27428,N_25730,N_26192);
xnor U27429 (N_27429,N_26089,N_25861);
nor U27430 (N_27430,N_25892,N_26012);
or U27431 (N_27431,N_26255,N_25637);
or U27432 (N_27432,N_25330,N_25905);
or U27433 (N_27433,N_25305,N_26202);
nand U27434 (N_27434,N_26002,N_26232);
xor U27435 (N_27435,N_26130,N_25946);
or U27436 (N_27436,N_26142,N_25343);
or U27437 (N_27437,N_26251,N_25658);
nand U27438 (N_27438,N_25203,N_26066);
and U27439 (N_27439,N_26189,N_25211);
or U27440 (N_27440,N_25515,N_26013);
nor U27441 (N_27441,N_25976,N_25522);
xor U27442 (N_27442,N_26338,N_26107);
xnor U27443 (N_27443,N_25677,N_25413);
or U27444 (N_27444,N_25522,N_25836);
nand U27445 (N_27445,N_26149,N_26094);
or U27446 (N_27446,N_25467,N_25801);
or U27447 (N_27447,N_26103,N_26129);
xnor U27448 (N_27448,N_25829,N_25884);
or U27449 (N_27449,N_26174,N_25568);
xor U27450 (N_27450,N_26265,N_26178);
nor U27451 (N_27451,N_26124,N_25522);
nand U27452 (N_27452,N_26043,N_25488);
nor U27453 (N_27453,N_25800,N_25256);
and U27454 (N_27454,N_26001,N_25419);
and U27455 (N_27455,N_25204,N_25605);
and U27456 (N_27456,N_26081,N_25765);
and U27457 (N_27457,N_25544,N_25542);
nor U27458 (N_27458,N_26086,N_26257);
nand U27459 (N_27459,N_26157,N_26082);
xnor U27460 (N_27460,N_25632,N_26064);
nand U27461 (N_27461,N_26366,N_25857);
or U27462 (N_27462,N_25332,N_26176);
or U27463 (N_27463,N_25659,N_26267);
and U27464 (N_27464,N_26116,N_25430);
or U27465 (N_27465,N_25839,N_25331);
xnor U27466 (N_27466,N_25780,N_26132);
xor U27467 (N_27467,N_25496,N_26338);
and U27468 (N_27468,N_26297,N_26371);
nor U27469 (N_27469,N_26365,N_25654);
nor U27470 (N_27470,N_25656,N_25970);
or U27471 (N_27471,N_25897,N_25919);
xor U27472 (N_27472,N_25281,N_25835);
and U27473 (N_27473,N_25730,N_25791);
xnor U27474 (N_27474,N_26277,N_25429);
and U27475 (N_27475,N_25547,N_25406);
nor U27476 (N_27476,N_25375,N_25486);
and U27477 (N_27477,N_26069,N_25842);
nand U27478 (N_27478,N_25581,N_26238);
nand U27479 (N_27479,N_26222,N_25294);
and U27480 (N_27480,N_25486,N_25405);
nand U27481 (N_27481,N_25881,N_25205);
xor U27482 (N_27482,N_26025,N_26347);
or U27483 (N_27483,N_25294,N_25897);
and U27484 (N_27484,N_25539,N_25387);
nor U27485 (N_27485,N_25371,N_25555);
nand U27486 (N_27486,N_25999,N_26290);
nor U27487 (N_27487,N_25944,N_25357);
nand U27488 (N_27488,N_25355,N_25533);
nand U27489 (N_27489,N_25435,N_25486);
nor U27490 (N_27490,N_25480,N_26161);
nor U27491 (N_27491,N_25713,N_25978);
and U27492 (N_27492,N_25818,N_26305);
nor U27493 (N_27493,N_25369,N_25945);
and U27494 (N_27494,N_25255,N_25440);
nor U27495 (N_27495,N_25910,N_25933);
nor U27496 (N_27496,N_26168,N_26193);
nand U27497 (N_27497,N_25236,N_25803);
nor U27498 (N_27498,N_25786,N_25317);
nor U27499 (N_27499,N_25275,N_25924);
or U27500 (N_27500,N_25900,N_25269);
or U27501 (N_27501,N_26082,N_25312);
nor U27502 (N_27502,N_26198,N_25905);
nor U27503 (N_27503,N_25444,N_26127);
nor U27504 (N_27504,N_26334,N_25747);
xnor U27505 (N_27505,N_25854,N_25911);
and U27506 (N_27506,N_25813,N_25477);
xor U27507 (N_27507,N_25547,N_25403);
xor U27508 (N_27508,N_26359,N_25512);
nor U27509 (N_27509,N_26147,N_25553);
or U27510 (N_27510,N_25829,N_25897);
nor U27511 (N_27511,N_25911,N_25278);
nand U27512 (N_27512,N_25714,N_25410);
nand U27513 (N_27513,N_25963,N_26134);
xnor U27514 (N_27514,N_25736,N_25512);
nand U27515 (N_27515,N_25286,N_25288);
or U27516 (N_27516,N_25205,N_25741);
and U27517 (N_27517,N_26148,N_25618);
nor U27518 (N_27518,N_26277,N_25224);
xor U27519 (N_27519,N_25593,N_25617);
nor U27520 (N_27520,N_25659,N_26339);
and U27521 (N_27521,N_25292,N_25912);
or U27522 (N_27522,N_25514,N_25386);
xnor U27523 (N_27523,N_25763,N_25574);
or U27524 (N_27524,N_26261,N_26390);
nor U27525 (N_27525,N_25751,N_25683);
xor U27526 (N_27526,N_25862,N_25631);
xor U27527 (N_27527,N_26030,N_25658);
nor U27528 (N_27528,N_25685,N_25696);
or U27529 (N_27529,N_26276,N_26310);
nand U27530 (N_27530,N_25918,N_26131);
or U27531 (N_27531,N_25961,N_25322);
xnor U27532 (N_27532,N_25613,N_25508);
nand U27533 (N_27533,N_26393,N_25868);
nor U27534 (N_27534,N_25844,N_25492);
xor U27535 (N_27535,N_25955,N_26202);
nand U27536 (N_27536,N_26160,N_25448);
nand U27537 (N_27537,N_26140,N_26377);
and U27538 (N_27538,N_25800,N_25989);
nor U27539 (N_27539,N_26328,N_25515);
xnor U27540 (N_27540,N_25451,N_26313);
or U27541 (N_27541,N_25672,N_26304);
xnor U27542 (N_27542,N_26245,N_25539);
nand U27543 (N_27543,N_25417,N_25386);
xor U27544 (N_27544,N_26168,N_25250);
and U27545 (N_27545,N_25927,N_26111);
nand U27546 (N_27546,N_26079,N_25352);
xnor U27547 (N_27547,N_25204,N_25316);
xnor U27548 (N_27548,N_25232,N_26073);
nand U27549 (N_27549,N_25258,N_25839);
nor U27550 (N_27550,N_25803,N_26058);
nor U27551 (N_27551,N_25425,N_25974);
or U27552 (N_27552,N_25305,N_25263);
nand U27553 (N_27553,N_26115,N_26281);
nand U27554 (N_27554,N_25629,N_25648);
and U27555 (N_27555,N_25860,N_25680);
nor U27556 (N_27556,N_26034,N_26050);
nor U27557 (N_27557,N_25898,N_25465);
xnor U27558 (N_27558,N_25440,N_26315);
nand U27559 (N_27559,N_25717,N_25303);
nor U27560 (N_27560,N_26179,N_25464);
xor U27561 (N_27561,N_26262,N_26264);
and U27562 (N_27562,N_25870,N_25797);
xor U27563 (N_27563,N_26221,N_25425);
xnor U27564 (N_27564,N_25815,N_26061);
or U27565 (N_27565,N_25828,N_25724);
and U27566 (N_27566,N_25302,N_25711);
nand U27567 (N_27567,N_25485,N_25454);
nor U27568 (N_27568,N_25945,N_25341);
nor U27569 (N_27569,N_26027,N_26294);
and U27570 (N_27570,N_25923,N_26311);
xnor U27571 (N_27571,N_25400,N_25721);
nor U27572 (N_27572,N_26098,N_26386);
or U27573 (N_27573,N_26047,N_26191);
and U27574 (N_27574,N_25799,N_26275);
nor U27575 (N_27575,N_25563,N_25277);
nand U27576 (N_27576,N_26134,N_25308);
and U27577 (N_27577,N_25843,N_25271);
xor U27578 (N_27578,N_25484,N_26135);
xor U27579 (N_27579,N_25270,N_25783);
xnor U27580 (N_27580,N_25965,N_26109);
xor U27581 (N_27581,N_26214,N_26026);
nor U27582 (N_27582,N_26336,N_25851);
or U27583 (N_27583,N_25788,N_25607);
nand U27584 (N_27584,N_25763,N_26154);
or U27585 (N_27585,N_25995,N_26076);
and U27586 (N_27586,N_25364,N_25392);
nand U27587 (N_27587,N_25566,N_26364);
nand U27588 (N_27588,N_26231,N_26276);
nor U27589 (N_27589,N_26093,N_26269);
and U27590 (N_27590,N_25699,N_26178);
and U27591 (N_27591,N_25441,N_25419);
nand U27592 (N_27592,N_25643,N_25830);
nand U27593 (N_27593,N_25946,N_25293);
nor U27594 (N_27594,N_26360,N_26298);
nor U27595 (N_27595,N_25236,N_26026);
nand U27596 (N_27596,N_25395,N_26119);
or U27597 (N_27597,N_25823,N_26035);
nand U27598 (N_27598,N_25860,N_25681);
nand U27599 (N_27599,N_26347,N_25792);
nor U27600 (N_27600,N_27286,N_26943);
nor U27601 (N_27601,N_26950,N_26913);
nand U27602 (N_27602,N_26909,N_26442);
or U27603 (N_27603,N_27350,N_26414);
nand U27604 (N_27604,N_27320,N_27386);
and U27605 (N_27605,N_26593,N_27497);
nor U27606 (N_27606,N_27063,N_26476);
or U27607 (N_27607,N_27112,N_26878);
or U27608 (N_27608,N_27029,N_26632);
or U27609 (N_27609,N_26844,N_27263);
nand U27610 (N_27610,N_27389,N_27444);
nand U27611 (N_27611,N_26885,N_26748);
or U27612 (N_27612,N_26852,N_26608);
or U27613 (N_27613,N_27394,N_26952);
nor U27614 (N_27614,N_26437,N_26827);
nor U27615 (N_27615,N_27363,N_26480);
and U27616 (N_27616,N_27473,N_26758);
xor U27617 (N_27617,N_26900,N_26911);
nand U27618 (N_27618,N_26497,N_26612);
and U27619 (N_27619,N_27194,N_27367);
xor U27620 (N_27620,N_27044,N_27231);
nand U27621 (N_27621,N_26797,N_26423);
nor U27622 (N_27622,N_26479,N_26542);
and U27623 (N_27623,N_26412,N_26435);
xor U27624 (N_27624,N_27448,N_26715);
nand U27625 (N_27625,N_27421,N_26651);
or U27626 (N_27626,N_27041,N_26471);
or U27627 (N_27627,N_26650,N_26594);
nand U27628 (N_27628,N_27519,N_26935);
or U27629 (N_27629,N_27494,N_26928);
nand U27630 (N_27630,N_27260,N_27356);
xor U27631 (N_27631,N_26982,N_26947);
and U27632 (N_27632,N_26857,N_27365);
or U27633 (N_27633,N_27294,N_27193);
nand U27634 (N_27634,N_26995,N_26426);
xor U27635 (N_27635,N_27304,N_27095);
or U27636 (N_27636,N_27065,N_26902);
and U27637 (N_27637,N_27078,N_26808);
xnor U27638 (N_27638,N_27317,N_26884);
nor U27639 (N_27639,N_26686,N_26417);
nand U27640 (N_27640,N_26996,N_26887);
and U27641 (N_27641,N_26907,N_27042);
xor U27642 (N_27642,N_26915,N_27300);
nand U27643 (N_27643,N_27007,N_27155);
and U27644 (N_27644,N_26820,N_27462);
or U27645 (N_27645,N_26851,N_26999);
and U27646 (N_27646,N_26755,N_26643);
xor U27647 (N_27647,N_26642,N_26511);
xnor U27648 (N_27648,N_27189,N_27414);
nor U27649 (N_27649,N_27434,N_26925);
and U27650 (N_27650,N_26464,N_26691);
and U27651 (N_27651,N_27293,N_26898);
xnor U27652 (N_27652,N_26545,N_26937);
nand U27653 (N_27653,N_26517,N_27492);
or U27654 (N_27654,N_26839,N_26421);
and U27655 (N_27655,N_27250,N_26795);
nand U27656 (N_27656,N_26835,N_27046);
xor U27657 (N_27657,N_26430,N_26836);
xor U27658 (N_27658,N_27113,N_27247);
or U27659 (N_27659,N_26550,N_27534);
or U27660 (N_27660,N_26962,N_26562);
nor U27661 (N_27661,N_26449,N_26949);
or U27662 (N_27662,N_27176,N_26726);
or U27663 (N_27663,N_26854,N_27028);
and U27664 (N_27664,N_26858,N_26527);
and U27665 (N_27665,N_26791,N_26829);
or U27666 (N_27666,N_26730,N_26802);
nor U27667 (N_27667,N_26655,N_26942);
nor U27668 (N_27668,N_26960,N_26500);
xor U27669 (N_27669,N_27117,N_27480);
xor U27670 (N_27670,N_27542,N_27520);
and U27671 (N_27671,N_26894,N_27005);
and U27672 (N_27672,N_26861,N_26514);
nor U27673 (N_27673,N_26618,N_26485);
or U27674 (N_27674,N_27200,N_26927);
xnor U27675 (N_27675,N_26600,N_26656);
nor U27676 (N_27676,N_27008,N_26638);
nand U27677 (N_27677,N_27119,N_26977);
or U27678 (N_27678,N_27285,N_26936);
xor U27679 (N_27679,N_27013,N_27171);
or U27680 (N_27680,N_27023,N_27220);
and U27681 (N_27681,N_27417,N_27196);
nor U27682 (N_27682,N_26867,N_27333);
xnor U27683 (N_27683,N_26870,N_26899);
and U27684 (N_27684,N_27488,N_26721);
or U27685 (N_27685,N_27128,N_27212);
or U27686 (N_27686,N_27526,N_27219);
nand U27687 (N_27687,N_26487,N_27390);
or U27688 (N_27688,N_27229,N_26871);
and U27689 (N_27689,N_27197,N_27207);
and U27690 (N_27690,N_27308,N_27109);
xnor U27691 (N_27691,N_27543,N_27545);
nand U27692 (N_27692,N_27116,N_26434);
nor U27693 (N_27693,N_26420,N_26664);
nor U27694 (N_27694,N_27129,N_27024);
and U27695 (N_27695,N_26742,N_27517);
and U27696 (N_27696,N_27156,N_27105);
xor U27697 (N_27697,N_27524,N_27221);
or U27698 (N_27698,N_27205,N_26645);
or U27699 (N_27699,N_27050,N_26780);
and U27700 (N_27700,N_26776,N_26408);
nor U27701 (N_27701,N_26714,N_26720);
nand U27702 (N_27702,N_27079,N_26483);
xnor U27703 (N_27703,N_27459,N_26616);
and U27704 (N_27704,N_27382,N_27596);
nand U27705 (N_27705,N_26433,N_26666);
nor U27706 (N_27706,N_26980,N_27073);
nor U27707 (N_27707,N_26478,N_26525);
or U27708 (N_27708,N_27115,N_26901);
or U27709 (N_27709,N_26892,N_27319);
and U27710 (N_27710,N_27407,N_26668);
nor U27711 (N_27711,N_26880,N_26706);
xnor U27712 (N_27712,N_27296,N_26559);
xor U27713 (N_27713,N_26577,N_26790);
nand U27714 (N_27714,N_26569,N_26971);
nor U27715 (N_27715,N_27477,N_27239);
xnor U27716 (N_27716,N_27233,N_27225);
and U27717 (N_27717,N_26964,N_27393);
nand U27718 (N_27718,N_27295,N_26912);
and U27719 (N_27719,N_26652,N_26516);
or U27720 (N_27720,N_27410,N_26474);
or U27721 (N_27721,N_27154,N_26922);
or U27722 (N_27722,N_26769,N_27489);
or U27723 (N_27723,N_27134,N_27313);
or U27724 (N_27724,N_26428,N_27476);
nand U27725 (N_27725,N_27080,N_27411);
nor U27726 (N_27726,N_27478,N_27159);
nand U27727 (N_27727,N_26419,N_26440);
xnor U27728 (N_27728,N_26853,N_26701);
or U27729 (N_27729,N_27375,N_26453);
nor U27730 (N_27730,N_27575,N_26679);
nand U27731 (N_27731,N_27438,N_27150);
xnor U27732 (N_27732,N_26764,N_27100);
and U27733 (N_27733,N_27589,N_27133);
or U27734 (N_27734,N_26567,N_27570);
nor U27735 (N_27735,N_26934,N_26498);
xor U27736 (N_27736,N_27351,N_26591);
xnor U27737 (N_27737,N_26708,N_27323);
nor U27738 (N_27738,N_27242,N_26573);
or U27739 (N_27739,N_27235,N_26889);
and U27740 (N_27740,N_27408,N_26495);
nand U27741 (N_27741,N_27036,N_27368);
and U27742 (N_27742,N_26817,N_26605);
nor U27743 (N_27743,N_26663,N_27214);
and U27744 (N_27744,N_27180,N_27525);
and U27745 (N_27745,N_26874,N_27572);
and U27746 (N_27746,N_27092,N_27192);
nor U27747 (N_27747,N_26452,N_27090);
xor U27748 (N_27748,N_27082,N_26418);
and U27749 (N_27749,N_26771,N_27465);
or U27750 (N_27750,N_26654,N_27051);
xor U27751 (N_27751,N_26546,N_27349);
and U27752 (N_27752,N_27172,N_27206);
xnor U27753 (N_27753,N_26634,N_26539);
nor U27754 (N_27754,N_27139,N_26717);
nand U27755 (N_27755,N_27198,N_26619);
or U27756 (N_27756,N_26929,N_26811);
xor U27757 (N_27757,N_27581,N_26403);
nor U27758 (N_27758,N_27508,N_26838);
nor U27759 (N_27759,N_26891,N_27157);
nand U27760 (N_27760,N_27290,N_27595);
nor U27761 (N_27761,N_27597,N_27321);
and U27762 (N_27762,N_27387,N_26905);
or U27763 (N_27763,N_26629,N_26568);
and U27764 (N_27764,N_27472,N_26683);
or U27765 (N_27765,N_26454,N_27280);
nand U27766 (N_27766,N_27305,N_26560);
or U27767 (N_27767,N_27071,N_26747);
nand U27768 (N_27768,N_26447,N_26917);
nor U27769 (N_27769,N_27096,N_26443);
nor U27770 (N_27770,N_26699,N_27467);
and U27771 (N_27771,N_27269,N_26985);
or U27772 (N_27772,N_27136,N_27289);
xnor U27773 (N_27773,N_27087,N_27377);
and U27774 (N_27774,N_27359,N_27422);
nor U27775 (N_27775,N_26620,N_27033);
and U27776 (N_27776,N_26866,N_27084);
xor U27777 (N_27777,N_26951,N_26675);
xor U27778 (N_27778,N_26722,N_26624);
nor U27779 (N_27779,N_27312,N_27215);
and U27780 (N_27780,N_27178,N_26723);
or U27781 (N_27781,N_27017,N_26680);
nor U27782 (N_27782,N_26636,N_27493);
nor U27783 (N_27783,N_26413,N_26606);
or U27784 (N_27784,N_26930,N_27236);
and U27785 (N_27785,N_27123,N_27164);
nand U27786 (N_27786,N_27506,N_27318);
or U27787 (N_27787,N_26875,N_26842);
nand U27788 (N_27788,N_27405,N_26639);
xor U27789 (N_27789,N_26596,N_26460);
and U27790 (N_27790,N_26425,N_27355);
xor U27791 (N_27791,N_26843,N_27152);
xnor U27792 (N_27792,N_26475,N_27412);
nor U27793 (N_27793,N_27081,N_26918);
xor U27794 (N_27794,N_27222,N_27259);
xnor U27795 (N_27795,N_27244,N_26993);
nor U27796 (N_27796,N_26767,N_26966);
or U27797 (N_27797,N_26580,N_27103);
and U27798 (N_27798,N_27107,N_27165);
and U27799 (N_27799,N_26729,N_27426);
nand U27800 (N_27800,N_26992,N_27279);
or U27801 (N_27801,N_26599,N_27429);
nor U27802 (N_27802,N_27151,N_26557);
nor U27803 (N_27803,N_27338,N_27076);
nor U27804 (N_27804,N_26973,N_27177);
or U27805 (N_27805,N_26762,N_27122);
or U27806 (N_27806,N_27565,N_26716);
or U27807 (N_27807,N_26646,N_26846);
or U27808 (N_27808,N_27278,N_26519);
nand U27809 (N_27809,N_27306,N_27070);
and U27810 (N_27810,N_27458,N_26965);
or U27811 (N_27811,N_26712,N_26731);
nor U27812 (N_27812,N_27077,N_26744);
xnor U27813 (N_27813,N_26696,N_27486);
or U27814 (N_27814,N_27550,N_26515);
or U27815 (N_27815,N_26728,N_26872);
or U27816 (N_27816,N_27471,N_27568);
xor U27817 (N_27817,N_26718,N_26556);
or U27818 (N_27818,N_27056,N_26969);
or U27819 (N_27819,N_27224,N_26687);
nor U27820 (N_27820,N_27153,N_27031);
and U27821 (N_27821,N_26526,N_27454);
nand U27822 (N_27822,N_27487,N_27371);
xnor U27823 (N_27823,N_27424,N_26578);
and U27824 (N_27824,N_27237,N_27327);
nor U27825 (N_27825,N_27252,N_27329);
nand U27826 (N_27826,N_27035,N_26761);
and U27827 (N_27827,N_26920,N_26828);
nor U27828 (N_27828,N_27413,N_27011);
or U27829 (N_27829,N_26725,N_26653);
nand U27830 (N_27830,N_26738,N_27549);
or U27831 (N_27831,N_26461,N_26532);
xor U27832 (N_27832,N_27284,N_26533);
nand U27833 (N_27833,N_27020,N_26782);
or U27834 (N_27834,N_27594,N_27001);
nand U27835 (N_27835,N_27039,N_27441);
nor U27836 (N_27836,N_27427,N_26753);
or U27837 (N_27837,N_27528,N_27273);
nor U27838 (N_27838,N_26484,N_27468);
nor U27839 (N_27839,N_27498,N_27240);
nor U27840 (N_27840,N_27253,N_26904);
nor U27841 (N_27841,N_26496,N_27199);
xor U27842 (N_27842,N_26531,N_26876);
and U27843 (N_27843,N_27057,N_26954);
nor U27844 (N_27844,N_26957,N_26592);
nor U27845 (N_27845,N_26908,N_26501);
xnor U27846 (N_27846,N_26416,N_26970);
nor U27847 (N_27847,N_26561,N_27110);
or U27848 (N_27848,N_27354,N_27243);
xor U27849 (N_27849,N_27352,N_26673);
nor U27850 (N_27850,N_27169,N_26575);
nor U27851 (N_27851,N_27392,N_26809);
xnor U27852 (N_27852,N_27264,N_26587);
and U27853 (N_27853,N_27014,N_26628);
nor U27854 (N_27854,N_26401,N_26963);
nor U27855 (N_27855,N_27012,N_27416);
and U27856 (N_27856,N_27055,N_26441);
and U27857 (N_27857,N_27288,N_27348);
nor U27858 (N_27858,N_26774,N_27030);
nor U27859 (N_27859,N_27353,N_27108);
nand U27860 (N_27860,N_26834,N_27188);
nor U27861 (N_27861,N_26850,N_26988);
nor U27862 (N_27862,N_26488,N_26648);
nand U27863 (N_27863,N_26490,N_26849);
or U27864 (N_27864,N_27579,N_26513);
nor U27865 (N_27865,N_27456,N_27464);
xor U27866 (N_27866,N_27381,N_27183);
or U27867 (N_27867,N_26446,N_26544);
xnor U27868 (N_27868,N_27201,N_26750);
or U27869 (N_27869,N_27432,N_27270);
xor U27870 (N_27870,N_27343,N_27450);
or U27871 (N_27871,N_26554,N_27587);
and U27872 (N_27872,N_26631,N_27578);
xnor U27873 (N_27873,N_27257,N_26611);
and U27874 (N_27874,N_27021,N_26644);
nand U27875 (N_27875,N_27449,N_26689);
or U27876 (N_27876,N_26543,N_27567);
xor U27877 (N_27877,N_26482,N_27086);
nand U27878 (N_27878,N_27258,N_26660);
or U27879 (N_27879,N_26402,N_27510);
or U27880 (N_27880,N_26800,N_26469);
xnor U27881 (N_27881,N_27435,N_26924);
nor U27882 (N_27882,N_26429,N_27527);
nor U27883 (N_27883,N_27255,N_27388);
and U27884 (N_27884,N_27370,N_26489);
or U27885 (N_27885,N_26986,N_27357);
xnor U27886 (N_27886,N_27060,N_26563);
xor U27887 (N_27887,N_27559,N_27563);
and U27888 (N_27888,N_27561,N_27218);
or U27889 (N_27889,N_26910,N_26504);
and U27890 (N_27890,N_26665,N_26535);
and U27891 (N_27891,N_27583,N_27554);
and U27892 (N_27892,N_27588,N_27453);
nor U27893 (N_27893,N_26404,N_26859);
nand U27894 (N_27894,N_27187,N_26953);
and U27895 (N_27895,N_27310,N_27470);
or U27896 (N_27896,N_26669,N_26868);
nand U27897 (N_27897,N_26522,N_27034);
nor U27898 (N_27898,N_26890,N_27491);
nor U27899 (N_27899,N_27261,N_27026);
or U27900 (N_27900,N_26555,N_27409);
or U27901 (N_27901,N_26760,N_27332);
xor U27902 (N_27902,N_26574,N_27141);
nand U27903 (N_27903,N_26819,N_26589);
nand U27904 (N_27904,N_26932,N_27400);
xnor U27905 (N_27905,N_26788,N_27292);
xor U27906 (N_27906,N_26524,N_27430);
or U27907 (N_27907,N_27303,N_27558);
and U27908 (N_27908,N_27437,N_26830);
xor U27909 (N_27909,N_27495,N_26987);
nand U27910 (N_27910,N_27170,N_27027);
or U27911 (N_27911,N_27521,N_27101);
xnor U27912 (N_27912,N_27420,N_27585);
xnor U27913 (N_27913,N_26815,N_27566);
and U27914 (N_27914,N_27158,N_26505);
nand U27915 (N_27915,N_26549,N_26812);
nor U27916 (N_27916,N_26837,N_26521);
or U27917 (N_27917,N_26778,N_27484);
and U27918 (N_27918,N_26923,N_27440);
and U27919 (N_27919,N_27537,N_26707);
or U27920 (N_27920,N_26822,N_26570);
and U27921 (N_27921,N_27513,N_26739);
xnor U27922 (N_27922,N_27569,N_26978);
or U27923 (N_27923,N_26450,N_26719);
nor U27924 (N_27924,N_27093,N_26407);
and U27925 (N_27925,N_27522,N_27111);
or U27926 (N_27926,N_27147,N_26536);
xnor U27927 (N_27927,N_27541,N_27358);
or U27928 (N_27928,N_27514,N_27053);
nand U27929 (N_27929,N_27203,N_27347);
nor U27930 (N_27930,N_26813,N_26411);
xnor U27931 (N_27931,N_26826,N_27475);
nor U27932 (N_27932,N_26967,N_26981);
nand U27933 (N_27933,N_27216,N_27474);
xnor U27934 (N_27934,N_27419,N_26921);
xnor U27935 (N_27935,N_26787,N_26678);
and U27936 (N_27936,N_27328,N_26990);
or U27937 (N_27937,N_27238,N_27398);
nand U27938 (N_27938,N_26462,N_27584);
xor U27939 (N_27939,N_26671,N_27266);
xor U27940 (N_27940,N_27102,N_26635);
and U27941 (N_27941,N_27277,N_26710);
or U27942 (N_27942,N_26510,N_26803);
and U27943 (N_27943,N_26553,N_27299);
nor U27944 (N_27944,N_26614,N_27058);
nand U27945 (N_27945,N_27245,N_27162);
nand U27946 (N_27946,N_27052,N_26582);
xor U27947 (N_27947,N_26734,N_27516);
nor U27948 (N_27948,N_27455,N_27019);
nor U27949 (N_27949,N_26733,N_26625);
xor U27950 (N_27950,N_27066,N_27059);
or U27951 (N_27951,N_27085,N_27457);
and U27952 (N_27952,N_26581,N_27291);
nand U27953 (N_27953,N_26896,N_27184);
nor U27954 (N_27954,N_27552,N_27364);
and U27955 (N_27955,N_27573,N_26685);
xnor U27956 (N_27956,N_26939,N_26732);
and U27957 (N_27957,N_26518,N_27135);
nor U27958 (N_27958,N_27463,N_26759);
xor U27959 (N_27959,N_26641,N_27385);
xnor U27960 (N_27960,N_26405,N_26424);
nor U27961 (N_27961,N_26786,N_26463);
and U27962 (N_27962,N_27548,N_27540);
xnor U27963 (N_27963,N_26459,N_26961);
xnor U27964 (N_27964,N_26700,N_26775);
nand U27965 (N_27965,N_26983,N_26630);
nand U27966 (N_27966,N_26972,N_26823);
or U27967 (N_27967,N_27335,N_27287);
nor U27968 (N_27968,N_26848,N_27340);
nor U27969 (N_27969,N_26622,N_27267);
or U27970 (N_27970,N_27345,N_27447);
nor U27971 (N_27971,N_27283,N_27511);
or U27972 (N_27972,N_27436,N_26796);
or U27973 (N_27973,N_27072,N_27282);
xor U27974 (N_27974,N_26724,N_26633);
nand U27975 (N_27975,N_26855,N_26979);
nor U27976 (N_27976,N_27089,N_26702);
nor U27977 (N_27977,N_27415,N_26766);
and U27978 (N_27978,N_27281,N_27009);
or U27979 (N_27979,N_27130,N_26688);
and U27980 (N_27980,N_26745,N_27586);
nand U27981 (N_27981,N_27125,N_27232);
xor U27982 (N_27982,N_26956,N_27166);
nor U27983 (N_27983,N_26431,N_27360);
or U27984 (N_27984,N_26933,N_27131);
xnor U27985 (N_27985,N_27175,N_26494);
or U27986 (N_27986,N_27538,N_26860);
or U27987 (N_27987,N_26406,N_26684);
and U27988 (N_27988,N_27376,N_27301);
or U27989 (N_27989,N_27309,N_27443);
nand U27990 (N_27990,N_26617,N_27262);
nor U27991 (N_27991,N_27018,N_27562);
or U27992 (N_27992,N_27582,N_27380);
xnor U27993 (N_27993,N_27167,N_26869);
and U27994 (N_27994,N_26818,N_26994);
or U27995 (N_27995,N_26640,N_26677);
nor U27996 (N_27996,N_27536,N_26806);
xor U27997 (N_27997,N_26579,N_26477);
nor U27998 (N_27998,N_27000,N_27339);
nor U27999 (N_27999,N_26455,N_26772);
xor U28000 (N_28000,N_27591,N_26697);
nand U28001 (N_28001,N_26770,N_26534);
xnor U28002 (N_28002,N_26509,N_26451);
xnor U28003 (N_28003,N_27179,N_26530);
xnor U28004 (N_28004,N_26955,N_26801);
or U28005 (N_28005,N_27397,N_26749);
nor U28006 (N_28006,N_26583,N_27316);
xor U28007 (N_28007,N_26941,N_26903);
and U28008 (N_28008,N_26658,N_27126);
and U28009 (N_28009,N_26916,N_26670);
or U28010 (N_28010,N_27479,N_27025);
nor U28011 (N_28011,N_27374,N_27483);
xnor U28012 (N_28012,N_27344,N_26709);
nor U28013 (N_28013,N_26422,N_27217);
nor U28014 (N_28014,N_26610,N_26615);
nor U28015 (N_28015,N_26507,N_26528);
xor U28016 (N_28016,N_26944,N_27576);
and U28017 (N_28017,N_27384,N_26958);
xnor U28018 (N_28018,N_26436,N_26777);
and U28019 (N_28019,N_26862,N_26551);
nor U28020 (N_28020,N_26727,N_26458);
xnor U28021 (N_28021,N_26410,N_27523);
nor U28022 (N_28022,N_26789,N_27515);
nor U28023 (N_28023,N_26975,N_27088);
or U28024 (N_28024,N_27590,N_27502);
or U28025 (N_28025,N_27334,N_27248);
nor U28026 (N_28026,N_26793,N_26989);
and U28027 (N_28027,N_26467,N_26816);
xnor U28028 (N_28028,N_26810,N_27564);
nor U28029 (N_28029,N_26465,N_27265);
nor U28030 (N_28030,N_27539,N_27598);
nor U28031 (N_28031,N_27431,N_27378);
xor U28032 (N_28032,N_26598,N_27307);
and U28033 (N_28033,N_26481,N_26883);
and U28034 (N_28034,N_27272,N_27406);
xnor U28035 (N_28035,N_26613,N_26698);
xor U28036 (N_28036,N_26492,N_26886);
nand U28037 (N_28037,N_27209,N_26792);
nand U28038 (N_28038,N_27302,N_26737);
nand U28039 (N_28039,N_27137,N_27592);
nor U28040 (N_28040,N_26741,N_26682);
xor U28041 (N_28041,N_27127,N_27106);
and U28042 (N_28042,N_26659,N_27213);
xor U28043 (N_28043,N_26662,N_27004);
and U28044 (N_28044,N_27223,N_26586);
and U28045 (N_28045,N_26704,N_26512);
nand U28046 (N_28046,N_26508,N_27362);
and U28047 (N_28047,N_27002,N_26456);
or U28048 (N_28048,N_26647,N_26604);
nor U28049 (N_28049,N_26506,N_26448);
xor U28050 (N_28050,N_27503,N_27553);
and U28051 (N_28051,N_26603,N_27532);
nor U28052 (N_28052,N_27251,N_27091);
nand U28053 (N_28053,N_26529,N_27433);
or U28054 (N_28054,N_26541,N_27439);
xor U28055 (N_28055,N_27230,N_26735);
xor U28056 (N_28056,N_27485,N_26623);
xor U28057 (N_28057,N_26667,N_26781);
and U28058 (N_28058,N_26547,N_27509);
xnor U28059 (N_28059,N_26968,N_27481);
and U28060 (N_28060,N_27161,N_27496);
and U28061 (N_28061,N_26637,N_26564);
or U28062 (N_28062,N_26690,N_27094);
xnor U28063 (N_28063,N_27190,N_27271);
or U28064 (N_28064,N_27249,N_26427);
and U28065 (N_28065,N_26831,N_27403);
or U28066 (N_28066,N_26627,N_26783);
nand U28067 (N_28067,N_26746,N_27551);
and U28068 (N_28068,N_27507,N_26444);
nor U28069 (N_28069,N_27418,N_27181);
or U28070 (N_28070,N_27163,N_27547);
or U28071 (N_28071,N_27202,N_27361);
nand U28072 (N_28072,N_27461,N_27186);
nand U28073 (N_28073,N_27191,N_26825);
nand U28074 (N_28074,N_26893,N_27211);
and U28075 (N_28075,N_27346,N_26784);
nor U28076 (N_28076,N_26538,N_27341);
or U28077 (N_28077,N_26540,N_27022);
nor U28078 (N_28078,N_27315,N_27256);
and U28079 (N_28079,N_26881,N_27535);
or U28080 (N_28080,N_27208,N_26584);
nand U28081 (N_28081,N_26864,N_26607);
and U28082 (N_28082,N_27142,N_27446);
xnor U28083 (N_28083,N_26703,N_27037);
and U28084 (N_28084,N_26445,N_26566);
nand U28085 (N_28085,N_26847,N_27227);
nand U28086 (N_28086,N_27075,N_27442);
nand U28087 (N_28087,N_27268,N_27143);
or U28088 (N_28088,N_27314,N_26491);
xor U28089 (N_28089,N_27326,N_27428);
nor U28090 (N_28090,N_26938,N_27451);
or U28091 (N_28091,N_27336,N_27574);
nand U28092 (N_28092,N_26895,N_26621);
and U28093 (N_28093,N_26998,N_27140);
xor U28094 (N_28094,N_27297,N_27580);
xnor U28095 (N_28095,N_26676,N_26595);
and U28096 (N_28096,N_26754,N_27010);
nor U28097 (N_28097,N_26572,N_27204);
and U28098 (N_28098,N_26695,N_27391);
nor U28099 (N_28099,N_27402,N_26503);
or U28100 (N_28100,N_27404,N_27546);
nand U28101 (N_28101,N_26984,N_26548);
xnor U28102 (N_28102,N_27048,N_27003);
or U28103 (N_28103,N_27557,N_26763);
nand U28104 (N_28104,N_26601,N_27395);
nand U28105 (N_28105,N_27555,N_26840);
nor U28106 (N_28106,N_26873,N_26824);
and U28107 (N_28107,N_26432,N_27124);
or U28108 (N_28108,N_26674,N_27067);
or U28109 (N_28109,N_26705,N_26785);
or U28110 (N_28110,N_27401,N_27366);
nor U28111 (N_28111,N_26409,N_27121);
xor U28112 (N_28112,N_26713,N_27015);
and U28113 (N_28113,N_26473,N_27132);
or U28114 (N_28114,N_27337,N_27423);
and U28115 (N_28115,N_27104,N_27006);
or U28116 (N_28116,N_27043,N_26537);
and U28117 (N_28117,N_27518,N_27399);
or U28118 (N_28118,N_27505,N_26931);
xor U28119 (N_28119,N_26602,N_27054);
nand U28120 (N_28120,N_27241,N_27530);
or U28121 (N_28121,N_27504,N_27275);
and U28122 (N_28122,N_26486,N_27556);
xor U28123 (N_28123,N_26736,N_27512);
xor U28124 (N_28124,N_27469,N_26997);
nor U28125 (N_28125,N_27445,N_26906);
xnor U28126 (N_28126,N_26948,N_27324);
xnor U28127 (N_28127,N_26863,N_26588);
and U28128 (N_28128,N_26693,N_27032);
xor U28129 (N_28129,N_27182,N_26681);
or U28130 (N_28130,N_26520,N_27064);
nand U28131 (N_28131,N_27049,N_27068);
xor U28132 (N_28132,N_27500,N_27174);
nand U28133 (N_28133,N_26845,N_26438);
nand U28134 (N_28134,N_27061,N_26856);
or U28135 (N_28135,N_26799,N_27045);
nand U28136 (N_28136,N_27118,N_26897);
or U28137 (N_28137,N_27040,N_26832);
xnor U28138 (N_28138,N_27138,N_26888);
and U28139 (N_28139,N_27544,N_26751);
and U28140 (N_28140,N_26841,N_27571);
nor U28141 (N_28141,N_27322,N_27149);
and U28142 (N_28142,N_27325,N_26472);
nand U28143 (N_28143,N_27098,N_27369);
nor U28144 (N_28144,N_26694,N_27062);
nand U28145 (N_28145,N_26711,N_26914);
nor U28146 (N_28146,N_26415,N_26400);
nand U28147 (N_28147,N_27298,N_26919);
and U28148 (N_28148,N_26805,N_27372);
or U28149 (N_28149,N_27097,N_27144);
or U28150 (N_28150,N_27425,N_26946);
nand U28151 (N_28151,N_27120,N_26765);
nor U28152 (N_28152,N_27460,N_27173);
nand U28153 (N_28153,N_26752,N_26974);
or U28154 (N_28154,N_26959,N_27083);
and U28155 (N_28155,N_27383,N_26814);
nor U28156 (N_28156,N_26585,N_26558);
or U28157 (N_28157,N_26740,N_27466);
nor U28158 (N_28158,N_27246,N_27195);
or U28159 (N_28159,N_26833,N_27185);
nor U28160 (N_28160,N_26649,N_26672);
nand U28161 (N_28161,N_27373,N_26757);
or U28162 (N_28162,N_27228,N_26493);
xnor U28163 (N_28163,N_26877,N_26743);
or U28164 (N_28164,N_27148,N_26523);
nand U28165 (N_28165,N_26439,N_27210);
xor U28166 (N_28166,N_27499,N_27311);
xnor U28167 (N_28167,N_27560,N_27342);
nor U28168 (N_28168,N_27160,N_26940);
or U28169 (N_28169,N_27234,N_27482);
nor U28170 (N_28170,N_27501,N_27099);
xnor U28171 (N_28171,N_26945,N_27452);
or U28172 (N_28172,N_27276,N_27396);
xor U28173 (N_28173,N_26926,N_27114);
xnor U28174 (N_28174,N_26626,N_26692);
nor U28175 (N_28175,N_27069,N_26879);
and U28176 (N_28176,N_26798,N_26466);
nor U28177 (N_28177,N_27016,N_27330);
or U28178 (N_28178,N_26661,N_26756);
nor U28179 (N_28179,N_27038,N_27593);
xnor U28180 (N_28180,N_26597,N_26457);
nand U28181 (N_28181,N_26804,N_26499);
and U28182 (N_28182,N_27533,N_27226);
and U28183 (N_28183,N_26552,N_27146);
xor U28184 (N_28184,N_27331,N_26865);
and U28185 (N_28185,N_27379,N_26590);
nor U28186 (N_28186,N_26565,N_26468);
and U28187 (N_28187,N_27274,N_27254);
nand U28188 (N_28188,N_26502,N_27529);
and U28189 (N_28189,N_26470,N_27599);
xnor U28190 (N_28190,N_26794,N_26576);
nor U28191 (N_28191,N_26991,N_26609);
nor U28192 (N_28192,N_26976,N_26571);
xnor U28193 (N_28193,N_27145,N_26773);
or U28194 (N_28194,N_27168,N_26882);
xnor U28195 (N_28195,N_27074,N_27047);
or U28196 (N_28196,N_26807,N_27531);
or U28197 (N_28197,N_26657,N_27490);
nand U28198 (N_28198,N_26768,N_27577);
or U28199 (N_28199,N_26779,N_26821);
and U28200 (N_28200,N_27396,N_26800);
nand U28201 (N_28201,N_26992,N_26790);
nand U28202 (N_28202,N_27167,N_27089);
and U28203 (N_28203,N_26984,N_27565);
or U28204 (N_28204,N_26486,N_27211);
nor U28205 (N_28205,N_26809,N_27409);
xor U28206 (N_28206,N_27298,N_27288);
and U28207 (N_28207,N_27341,N_27141);
xor U28208 (N_28208,N_27322,N_26876);
or U28209 (N_28209,N_26714,N_27099);
nand U28210 (N_28210,N_27076,N_26898);
or U28211 (N_28211,N_27269,N_27438);
nand U28212 (N_28212,N_26800,N_26428);
or U28213 (N_28213,N_26921,N_26687);
nor U28214 (N_28214,N_27274,N_26914);
and U28215 (N_28215,N_27334,N_26547);
nor U28216 (N_28216,N_27424,N_26442);
xor U28217 (N_28217,N_27014,N_26430);
or U28218 (N_28218,N_27317,N_26929);
xnor U28219 (N_28219,N_27287,N_27444);
nand U28220 (N_28220,N_26989,N_26922);
and U28221 (N_28221,N_26610,N_26865);
and U28222 (N_28222,N_26680,N_27323);
xor U28223 (N_28223,N_27480,N_27161);
xor U28224 (N_28224,N_26496,N_27392);
or U28225 (N_28225,N_27468,N_26605);
and U28226 (N_28226,N_27089,N_27325);
and U28227 (N_28227,N_27385,N_26618);
xnor U28228 (N_28228,N_27526,N_27451);
xor U28229 (N_28229,N_26453,N_27470);
xor U28230 (N_28230,N_27064,N_26770);
xnor U28231 (N_28231,N_27558,N_26959);
or U28232 (N_28232,N_27039,N_27222);
and U28233 (N_28233,N_26917,N_26949);
nor U28234 (N_28234,N_26803,N_27460);
nand U28235 (N_28235,N_27128,N_27079);
nor U28236 (N_28236,N_26907,N_26814);
xor U28237 (N_28237,N_26832,N_26520);
xor U28238 (N_28238,N_26508,N_27167);
or U28239 (N_28239,N_26494,N_26585);
xnor U28240 (N_28240,N_26483,N_27492);
xnor U28241 (N_28241,N_26678,N_26627);
or U28242 (N_28242,N_27119,N_27260);
and U28243 (N_28243,N_27268,N_26400);
or U28244 (N_28244,N_27129,N_26409);
nor U28245 (N_28245,N_26481,N_27426);
nor U28246 (N_28246,N_27200,N_26932);
nand U28247 (N_28247,N_27072,N_27138);
xor U28248 (N_28248,N_27339,N_26430);
nor U28249 (N_28249,N_27295,N_27404);
xor U28250 (N_28250,N_26946,N_27109);
xnor U28251 (N_28251,N_27046,N_27350);
or U28252 (N_28252,N_26491,N_27517);
xor U28253 (N_28253,N_27179,N_27334);
nand U28254 (N_28254,N_26938,N_27276);
nand U28255 (N_28255,N_27156,N_27531);
nand U28256 (N_28256,N_26864,N_26546);
or U28257 (N_28257,N_26961,N_26937);
and U28258 (N_28258,N_27556,N_26878);
and U28259 (N_28259,N_26901,N_27358);
and U28260 (N_28260,N_27586,N_26996);
nor U28261 (N_28261,N_26700,N_27249);
or U28262 (N_28262,N_27468,N_26760);
nand U28263 (N_28263,N_27520,N_27040);
and U28264 (N_28264,N_27540,N_27422);
and U28265 (N_28265,N_27116,N_27290);
and U28266 (N_28266,N_26975,N_27447);
nand U28267 (N_28267,N_27321,N_26549);
nand U28268 (N_28268,N_26459,N_27049);
or U28269 (N_28269,N_27312,N_26418);
nor U28270 (N_28270,N_26944,N_26493);
or U28271 (N_28271,N_26789,N_27130);
nand U28272 (N_28272,N_26498,N_27118);
nand U28273 (N_28273,N_26607,N_26636);
xnor U28274 (N_28274,N_26564,N_26945);
and U28275 (N_28275,N_27200,N_27587);
or U28276 (N_28276,N_27498,N_26418);
nand U28277 (N_28277,N_27205,N_26502);
nor U28278 (N_28278,N_26588,N_27229);
nand U28279 (N_28279,N_26477,N_27287);
nor U28280 (N_28280,N_26798,N_27139);
nand U28281 (N_28281,N_26435,N_26622);
nor U28282 (N_28282,N_27028,N_26522);
and U28283 (N_28283,N_26774,N_26464);
and U28284 (N_28284,N_26965,N_27161);
nor U28285 (N_28285,N_27012,N_27451);
xor U28286 (N_28286,N_26920,N_26704);
nor U28287 (N_28287,N_27028,N_27096);
xnor U28288 (N_28288,N_26532,N_26598);
or U28289 (N_28289,N_27441,N_27438);
and U28290 (N_28290,N_27216,N_26962);
nor U28291 (N_28291,N_26880,N_27030);
nand U28292 (N_28292,N_26454,N_26443);
nor U28293 (N_28293,N_27119,N_27471);
xor U28294 (N_28294,N_26437,N_26539);
nor U28295 (N_28295,N_27250,N_26604);
and U28296 (N_28296,N_26765,N_26846);
nor U28297 (N_28297,N_26595,N_26623);
or U28298 (N_28298,N_27452,N_26432);
nor U28299 (N_28299,N_26854,N_26899);
and U28300 (N_28300,N_27418,N_27090);
nor U28301 (N_28301,N_27125,N_26791);
nor U28302 (N_28302,N_27371,N_27195);
nor U28303 (N_28303,N_26754,N_26664);
or U28304 (N_28304,N_26886,N_27301);
or U28305 (N_28305,N_26561,N_26975);
nand U28306 (N_28306,N_27033,N_27275);
and U28307 (N_28307,N_27115,N_26908);
nor U28308 (N_28308,N_27138,N_27506);
and U28309 (N_28309,N_26558,N_26784);
xor U28310 (N_28310,N_26685,N_27068);
nor U28311 (N_28311,N_27308,N_27483);
xor U28312 (N_28312,N_27544,N_27551);
nor U28313 (N_28313,N_26512,N_27382);
nor U28314 (N_28314,N_27206,N_26585);
or U28315 (N_28315,N_27513,N_26600);
nand U28316 (N_28316,N_26817,N_27510);
xor U28317 (N_28317,N_26892,N_27426);
nand U28318 (N_28318,N_26462,N_26403);
xor U28319 (N_28319,N_27220,N_26962);
or U28320 (N_28320,N_27525,N_27230);
xor U28321 (N_28321,N_26611,N_26452);
or U28322 (N_28322,N_27313,N_26940);
nand U28323 (N_28323,N_26502,N_26628);
xor U28324 (N_28324,N_27533,N_26537);
nor U28325 (N_28325,N_26775,N_27169);
nand U28326 (N_28326,N_27295,N_26704);
and U28327 (N_28327,N_27382,N_26677);
nand U28328 (N_28328,N_26532,N_26509);
nand U28329 (N_28329,N_26578,N_27172);
nand U28330 (N_28330,N_27073,N_27224);
nor U28331 (N_28331,N_27123,N_27150);
nand U28332 (N_28332,N_26883,N_26841);
xor U28333 (N_28333,N_26751,N_26653);
xnor U28334 (N_28334,N_27137,N_27456);
xnor U28335 (N_28335,N_26762,N_26906);
or U28336 (N_28336,N_27566,N_27283);
xor U28337 (N_28337,N_27336,N_26868);
nor U28338 (N_28338,N_27428,N_26908);
or U28339 (N_28339,N_27304,N_27516);
xnor U28340 (N_28340,N_26985,N_27472);
and U28341 (N_28341,N_26755,N_27524);
and U28342 (N_28342,N_26580,N_27182);
xor U28343 (N_28343,N_27418,N_26966);
or U28344 (N_28344,N_27526,N_26413);
xnor U28345 (N_28345,N_26522,N_26807);
nor U28346 (N_28346,N_27599,N_27404);
or U28347 (N_28347,N_27377,N_26868);
nand U28348 (N_28348,N_26807,N_26844);
and U28349 (N_28349,N_27236,N_26913);
and U28350 (N_28350,N_27460,N_27340);
nand U28351 (N_28351,N_26854,N_26965);
or U28352 (N_28352,N_27048,N_26401);
xnor U28353 (N_28353,N_26916,N_26424);
and U28354 (N_28354,N_26756,N_27230);
and U28355 (N_28355,N_27336,N_27157);
nor U28356 (N_28356,N_26753,N_27442);
nand U28357 (N_28357,N_26745,N_27139);
nand U28358 (N_28358,N_27175,N_26518);
xnor U28359 (N_28359,N_26458,N_27532);
nor U28360 (N_28360,N_27470,N_27091);
nor U28361 (N_28361,N_27362,N_26441);
nand U28362 (N_28362,N_26419,N_26501);
nand U28363 (N_28363,N_27262,N_26473);
or U28364 (N_28364,N_27577,N_26698);
and U28365 (N_28365,N_26787,N_27382);
nor U28366 (N_28366,N_26594,N_26464);
xnor U28367 (N_28367,N_26505,N_27109);
nor U28368 (N_28368,N_27178,N_26478);
and U28369 (N_28369,N_27479,N_27569);
nand U28370 (N_28370,N_26525,N_27109);
xor U28371 (N_28371,N_27306,N_26426);
and U28372 (N_28372,N_26959,N_27578);
nor U28373 (N_28373,N_27201,N_26904);
nand U28374 (N_28374,N_27398,N_26434);
nor U28375 (N_28375,N_26459,N_26988);
nand U28376 (N_28376,N_26698,N_27302);
xnor U28377 (N_28377,N_27086,N_26935);
xnor U28378 (N_28378,N_27032,N_26754);
and U28379 (N_28379,N_27047,N_26419);
or U28380 (N_28380,N_26543,N_27094);
nand U28381 (N_28381,N_27484,N_26600);
nor U28382 (N_28382,N_27196,N_27026);
or U28383 (N_28383,N_26524,N_26643);
nand U28384 (N_28384,N_27099,N_27526);
nand U28385 (N_28385,N_26629,N_26762);
xnor U28386 (N_28386,N_27596,N_27142);
or U28387 (N_28387,N_27062,N_27224);
and U28388 (N_28388,N_27237,N_26774);
nand U28389 (N_28389,N_26626,N_26527);
xor U28390 (N_28390,N_26613,N_26792);
nor U28391 (N_28391,N_27506,N_27437);
nand U28392 (N_28392,N_26849,N_27381);
or U28393 (N_28393,N_26746,N_27444);
or U28394 (N_28394,N_26822,N_26418);
and U28395 (N_28395,N_26702,N_27222);
xnor U28396 (N_28396,N_27136,N_27463);
nor U28397 (N_28397,N_27189,N_27113);
xor U28398 (N_28398,N_26993,N_27188);
nor U28399 (N_28399,N_27340,N_26432);
or U28400 (N_28400,N_26530,N_27108);
or U28401 (N_28401,N_27379,N_26648);
nor U28402 (N_28402,N_26740,N_27034);
nand U28403 (N_28403,N_27594,N_26478);
or U28404 (N_28404,N_26998,N_26731);
xor U28405 (N_28405,N_27036,N_27087);
xnor U28406 (N_28406,N_26990,N_27368);
or U28407 (N_28407,N_26414,N_27393);
nor U28408 (N_28408,N_26413,N_26684);
and U28409 (N_28409,N_26466,N_27406);
or U28410 (N_28410,N_26833,N_27468);
or U28411 (N_28411,N_27314,N_27206);
nor U28412 (N_28412,N_26996,N_26794);
or U28413 (N_28413,N_27408,N_26951);
or U28414 (N_28414,N_27079,N_27221);
or U28415 (N_28415,N_27457,N_27137);
xnor U28416 (N_28416,N_26664,N_26904);
nand U28417 (N_28417,N_27392,N_27580);
nor U28418 (N_28418,N_26581,N_26572);
and U28419 (N_28419,N_26545,N_26799);
or U28420 (N_28420,N_27490,N_27034);
xor U28421 (N_28421,N_27198,N_27527);
nand U28422 (N_28422,N_27126,N_26405);
xnor U28423 (N_28423,N_27433,N_27219);
and U28424 (N_28424,N_27418,N_27127);
nand U28425 (N_28425,N_27448,N_26735);
and U28426 (N_28426,N_27034,N_27411);
or U28427 (N_28427,N_27155,N_26523);
nor U28428 (N_28428,N_27317,N_27136);
or U28429 (N_28429,N_26656,N_27147);
xor U28430 (N_28430,N_27511,N_26674);
or U28431 (N_28431,N_27485,N_26647);
nand U28432 (N_28432,N_26460,N_26918);
or U28433 (N_28433,N_27526,N_27274);
and U28434 (N_28434,N_27107,N_27080);
nand U28435 (N_28435,N_26621,N_27333);
and U28436 (N_28436,N_26511,N_26590);
and U28437 (N_28437,N_27037,N_27337);
nor U28438 (N_28438,N_27384,N_27473);
and U28439 (N_28439,N_26820,N_27594);
nand U28440 (N_28440,N_27428,N_26885);
and U28441 (N_28441,N_27496,N_27551);
or U28442 (N_28442,N_26641,N_26969);
and U28443 (N_28443,N_27350,N_26992);
or U28444 (N_28444,N_26529,N_26881);
xnor U28445 (N_28445,N_27400,N_26413);
nand U28446 (N_28446,N_27108,N_27306);
and U28447 (N_28447,N_27303,N_26704);
nor U28448 (N_28448,N_26457,N_26690);
and U28449 (N_28449,N_27136,N_26719);
xnor U28450 (N_28450,N_26555,N_27429);
nor U28451 (N_28451,N_27136,N_27520);
nor U28452 (N_28452,N_26850,N_27450);
or U28453 (N_28453,N_27597,N_26998);
nand U28454 (N_28454,N_26847,N_27581);
xor U28455 (N_28455,N_26775,N_27305);
and U28456 (N_28456,N_26649,N_27307);
and U28457 (N_28457,N_27168,N_27346);
nand U28458 (N_28458,N_27375,N_27162);
or U28459 (N_28459,N_26670,N_27353);
xor U28460 (N_28460,N_27258,N_27276);
xor U28461 (N_28461,N_26944,N_26584);
nor U28462 (N_28462,N_27444,N_26479);
nor U28463 (N_28463,N_26946,N_26427);
xnor U28464 (N_28464,N_27175,N_27052);
nor U28465 (N_28465,N_26980,N_26529);
xor U28466 (N_28466,N_27558,N_27250);
nor U28467 (N_28467,N_27290,N_27513);
or U28468 (N_28468,N_26946,N_27130);
and U28469 (N_28469,N_27416,N_27325);
xor U28470 (N_28470,N_26833,N_27429);
and U28471 (N_28471,N_26486,N_26412);
xnor U28472 (N_28472,N_26517,N_26881);
and U28473 (N_28473,N_27209,N_26786);
nor U28474 (N_28474,N_27058,N_27480);
nand U28475 (N_28475,N_27558,N_26770);
and U28476 (N_28476,N_27274,N_26507);
nand U28477 (N_28477,N_26650,N_27388);
and U28478 (N_28478,N_26518,N_27536);
and U28479 (N_28479,N_26783,N_27446);
nor U28480 (N_28480,N_26870,N_27364);
nor U28481 (N_28481,N_26737,N_26670);
xnor U28482 (N_28482,N_27130,N_27361);
and U28483 (N_28483,N_26836,N_26923);
nor U28484 (N_28484,N_27226,N_26425);
nand U28485 (N_28485,N_27056,N_26975);
xor U28486 (N_28486,N_27548,N_26505);
and U28487 (N_28487,N_27353,N_26462);
nand U28488 (N_28488,N_26481,N_27311);
nand U28489 (N_28489,N_26904,N_26510);
xor U28490 (N_28490,N_27088,N_27129);
nor U28491 (N_28491,N_26787,N_26420);
xnor U28492 (N_28492,N_26743,N_27454);
and U28493 (N_28493,N_27186,N_27084);
nand U28494 (N_28494,N_27495,N_27364);
nor U28495 (N_28495,N_27190,N_27578);
xor U28496 (N_28496,N_26705,N_27001);
and U28497 (N_28497,N_26797,N_26825);
xnor U28498 (N_28498,N_27403,N_26980);
or U28499 (N_28499,N_26782,N_27500);
nand U28500 (N_28500,N_27072,N_27229);
and U28501 (N_28501,N_26635,N_27344);
and U28502 (N_28502,N_27456,N_27008);
and U28503 (N_28503,N_27509,N_26872);
nor U28504 (N_28504,N_26839,N_26565);
nor U28505 (N_28505,N_27397,N_26549);
nor U28506 (N_28506,N_26660,N_27140);
nand U28507 (N_28507,N_27306,N_27201);
nor U28508 (N_28508,N_27305,N_26423);
nand U28509 (N_28509,N_27481,N_26996);
nand U28510 (N_28510,N_26661,N_26700);
or U28511 (N_28511,N_27440,N_27555);
xnor U28512 (N_28512,N_26796,N_27055);
xnor U28513 (N_28513,N_26523,N_27383);
or U28514 (N_28514,N_26681,N_27025);
xnor U28515 (N_28515,N_27346,N_26983);
or U28516 (N_28516,N_26720,N_26674);
and U28517 (N_28517,N_27039,N_26476);
nand U28518 (N_28518,N_27573,N_27437);
xnor U28519 (N_28519,N_27055,N_27587);
nand U28520 (N_28520,N_27164,N_27461);
nor U28521 (N_28521,N_26725,N_27483);
nor U28522 (N_28522,N_26997,N_27001);
and U28523 (N_28523,N_27102,N_27048);
nor U28524 (N_28524,N_27505,N_26509);
nand U28525 (N_28525,N_27239,N_26725);
xor U28526 (N_28526,N_26984,N_27007);
or U28527 (N_28527,N_26797,N_27592);
xnor U28528 (N_28528,N_26517,N_27521);
nor U28529 (N_28529,N_26736,N_26789);
or U28530 (N_28530,N_26575,N_26873);
nand U28531 (N_28531,N_27006,N_27441);
nand U28532 (N_28532,N_27168,N_27372);
xor U28533 (N_28533,N_27427,N_26826);
or U28534 (N_28534,N_27279,N_26663);
nor U28535 (N_28535,N_26524,N_26631);
nor U28536 (N_28536,N_27281,N_26624);
or U28537 (N_28537,N_27451,N_26889);
xnor U28538 (N_28538,N_27268,N_27002);
nand U28539 (N_28539,N_27058,N_26970);
and U28540 (N_28540,N_26980,N_27483);
nor U28541 (N_28541,N_26754,N_26750);
and U28542 (N_28542,N_27494,N_26750);
xor U28543 (N_28543,N_27434,N_27086);
xor U28544 (N_28544,N_27351,N_26826);
nand U28545 (N_28545,N_26832,N_26611);
or U28546 (N_28546,N_27544,N_27478);
nor U28547 (N_28547,N_26638,N_26592);
xor U28548 (N_28548,N_27480,N_26568);
or U28549 (N_28549,N_26494,N_27108);
and U28550 (N_28550,N_26869,N_27585);
nand U28551 (N_28551,N_26583,N_27209);
nor U28552 (N_28552,N_26774,N_26799);
or U28553 (N_28553,N_26974,N_26518);
nor U28554 (N_28554,N_27514,N_27070);
and U28555 (N_28555,N_27013,N_27143);
and U28556 (N_28556,N_26990,N_27303);
nor U28557 (N_28557,N_27590,N_27112);
or U28558 (N_28558,N_27035,N_27251);
nor U28559 (N_28559,N_27524,N_26757);
nand U28560 (N_28560,N_27222,N_26668);
or U28561 (N_28561,N_26834,N_26815);
xor U28562 (N_28562,N_26969,N_27482);
nand U28563 (N_28563,N_26943,N_27037);
xnor U28564 (N_28564,N_26813,N_26483);
nand U28565 (N_28565,N_27361,N_26585);
xnor U28566 (N_28566,N_26980,N_27555);
xnor U28567 (N_28567,N_26773,N_26822);
and U28568 (N_28568,N_27179,N_27363);
or U28569 (N_28569,N_27410,N_27430);
or U28570 (N_28570,N_26837,N_26426);
nor U28571 (N_28571,N_27334,N_26849);
or U28572 (N_28572,N_27495,N_26858);
nand U28573 (N_28573,N_26483,N_27317);
nand U28574 (N_28574,N_27594,N_26839);
or U28575 (N_28575,N_26901,N_26408);
or U28576 (N_28576,N_27374,N_27014);
nand U28577 (N_28577,N_26930,N_27292);
and U28578 (N_28578,N_27036,N_26760);
and U28579 (N_28579,N_26897,N_27026);
xnor U28580 (N_28580,N_27416,N_26869);
xor U28581 (N_28581,N_27129,N_26819);
nand U28582 (N_28582,N_26841,N_26877);
nor U28583 (N_28583,N_26690,N_26547);
xnor U28584 (N_28584,N_27125,N_27181);
and U28585 (N_28585,N_26447,N_26717);
nand U28586 (N_28586,N_26401,N_26783);
xnor U28587 (N_28587,N_27265,N_27425);
xor U28588 (N_28588,N_26497,N_27094);
xnor U28589 (N_28589,N_26454,N_27558);
nor U28590 (N_28590,N_26401,N_26695);
nor U28591 (N_28591,N_26411,N_26568);
nor U28592 (N_28592,N_26747,N_27158);
and U28593 (N_28593,N_27409,N_26476);
nor U28594 (N_28594,N_27247,N_26895);
nand U28595 (N_28595,N_27387,N_26753);
nand U28596 (N_28596,N_27592,N_27221);
or U28597 (N_28597,N_26917,N_27243);
nor U28598 (N_28598,N_27003,N_26625);
xor U28599 (N_28599,N_27545,N_26511);
or U28600 (N_28600,N_26425,N_27293);
nor U28601 (N_28601,N_27479,N_26904);
nor U28602 (N_28602,N_26443,N_27358);
nor U28603 (N_28603,N_27374,N_26613);
xor U28604 (N_28604,N_27535,N_27108);
nand U28605 (N_28605,N_26566,N_27501);
nor U28606 (N_28606,N_26782,N_26771);
nor U28607 (N_28607,N_27097,N_27122);
nand U28608 (N_28608,N_26766,N_27026);
xnor U28609 (N_28609,N_26538,N_26849);
xnor U28610 (N_28610,N_26669,N_27415);
nor U28611 (N_28611,N_27371,N_27338);
or U28612 (N_28612,N_26669,N_27043);
and U28613 (N_28613,N_26443,N_27490);
nand U28614 (N_28614,N_26736,N_26665);
and U28615 (N_28615,N_26983,N_26633);
nor U28616 (N_28616,N_27086,N_26490);
or U28617 (N_28617,N_26618,N_26970);
or U28618 (N_28618,N_26874,N_26606);
xor U28619 (N_28619,N_27201,N_27164);
and U28620 (N_28620,N_27032,N_27278);
or U28621 (N_28621,N_26714,N_26911);
and U28622 (N_28622,N_27494,N_27335);
and U28623 (N_28623,N_27122,N_27281);
or U28624 (N_28624,N_27381,N_27169);
xnor U28625 (N_28625,N_26773,N_26480);
nor U28626 (N_28626,N_26808,N_26833);
or U28627 (N_28627,N_26540,N_26495);
nand U28628 (N_28628,N_27085,N_27348);
nand U28629 (N_28629,N_26656,N_27353);
nor U28630 (N_28630,N_27396,N_27249);
nor U28631 (N_28631,N_26713,N_27082);
or U28632 (N_28632,N_27282,N_26897);
or U28633 (N_28633,N_26742,N_27141);
nand U28634 (N_28634,N_26505,N_26650);
nand U28635 (N_28635,N_27213,N_26631);
and U28636 (N_28636,N_26759,N_26987);
nor U28637 (N_28637,N_26893,N_26878);
nor U28638 (N_28638,N_27556,N_27510);
or U28639 (N_28639,N_26877,N_27498);
xnor U28640 (N_28640,N_27398,N_26724);
nand U28641 (N_28641,N_26580,N_27290);
or U28642 (N_28642,N_26547,N_27054);
xor U28643 (N_28643,N_27216,N_26660);
nand U28644 (N_28644,N_27378,N_27318);
or U28645 (N_28645,N_26529,N_26428);
nor U28646 (N_28646,N_26936,N_27002);
nor U28647 (N_28647,N_26936,N_27069);
or U28648 (N_28648,N_27567,N_26581);
nor U28649 (N_28649,N_27029,N_27118);
and U28650 (N_28650,N_26992,N_26510);
xor U28651 (N_28651,N_26547,N_27114);
xnor U28652 (N_28652,N_26732,N_27250);
and U28653 (N_28653,N_26785,N_27560);
or U28654 (N_28654,N_26627,N_27303);
or U28655 (N_28655,N_27257,N_27275);
nor U28656 (N_28656,N_27189,N_27408);
nor U28657 (N_28657,N_27137,N_26458);
nor U28658 (N_28658,N_27016,N_27060);
and U28659 (N_28659,N_27110,N_26807);
or U28660 (N_28660,N_27097,N_27437);
or U28661 (N_28661,N_26926,N_26643);
and U28662 (N_28662,N_27146,N_27229);
or U28663 (N_28663,N_27198,N_27108);
or U28664 (N_28664,N_27049,N_27148);
or U28665 (N_28665,N_26520,N_26777);
nor U28666 (N_28666,N_27074,N_26669);
nor U28667 (N_28667,N_27512,N_27530);
or U28668 (N_28668,N_26636,N_26421);
nand U28669 (N_28669,N_26539,N_27347);
nand U28670 (N_28670,N_26696,N_27314);
nand U28671 (N_28671,N_27292,N_27299);
and U28672 (N_28672,N_26637,N_26432);
and U28673 (N_28673,N_27277,N_27091);
nor U28674 (N_28674,N_27306,N_27480);
or U28675 (N_28675,N_27578,N_27373);
xnor U28676 (N_28676,N_26773,N_27452);
xnor U28677 (N_28677,N_26620,N_27059);
xor U28678 (N_28678,N_26834,N_27365);
and U28679 (N_28679,N_26531,N_26466);
nor U28680 (N_28680,N_27010,N_26592);
nand U28681 (N_28681,N_26832,N_26447);
or U28682 (N_28682,N_26893,N_26605);
and U28683 (N_28683,N_27189,N_27353);
nor U28684 (N_28684,N_26996,N_27230);
xor U28685 (N_28685,N_26730,N_26509);
and U28686 (N_28686,N_27293,N_26765);
and U28687 (N_28687,N_27380,N_26835);
xnor U28688 (N_28688,N_27062,N_26537);
and U28689 (N_28689,N_27348,N_26745);
or U28690 (N_28690,N_26436,N_27168);
nor U28691 (N_28691,N_26717,N_26601);
xnor U28692 (N_28692,N_27439,N_26527);
nand U28693 (N_28693,N_26958,N_27350);
or U28694 (N_28694,N_27197,N_26446);
nor U28695 (N_28695,N_26728,N_26464);
or U28696 (N_28696,N_26871,N_27223);
xnor U28697 (N_28697,N_26899,N_26758);
xor U28698 (N_28698,N_26825,N_27410);
nand U28699 (N_28699,N_27147,N_27538);
or U28700 (N_28700,N_27164,N_27468);
xnor U28701 (N_28701,N_26614,N_27593);
nor U28702 (N_28702,N_26871,N_26725);
or U28703 (N_28703,N_27428,N_27053);
nor U28704 (N_28704,N_26703,N_27472);
or U28705 (N_28705,N_26606,N_26722);
nor U28706 (N_28706,N_26428,N_27358);
and U28707 (N_28707,N_27441,N_27045);
xnor U28708 (N_28708,N_27496,N_26932);
nor U28709 (N_28709,N_26533,N_26556);
xor U28710 (N_28710,N_27556,N_26968);
nor U28711 (N_28711,N_27234,N_26604);
and U28712 (N_28712,N_27437,N_27084);
and U28713 (N_28713,N_27404,N_26814);
nand U28714 (N_28714,N_27109,N_27157);
nand U28715 (N_28715,N_27052,N_27117);
nand U28716 (N_28716,N_27511,N_27169);
and U28717 (N_28717,N_27143,N_27005);
nor U28718 (N_28718,N_26599,N_27018);
xnor U28719 (N_28719,N_26428,N_26950);
nand U28720 (N_28720,N_27273,N_26493);
xor U28721 (N_28721,N_26915,N_27283);
and U28722 (N_28722,N_26870,N_27489);
and U28723 (N_28723,N_27341,N_26539);
xnor U28724 (N_28724,N_26546,N_26473);
and U28725 (N_28725,N_27076,N_26410);
or U28726 (N_28726,N_26735,N_27588);
nor U28727 (N_28727,N_27336,N_26608);
or U28728 (N_28728,N_26687,N_26576);
nor U28729 (N_28729,N_27021,N_26705);
nor U28730 (N_28730,N_26677,N_27413);
nor U28731 (N_28731,N_27595,N_27475);
and U28732 (N_28732,N_26684,N_27163);
nand U28733 (N_28733,N_26983,N_27411);
or U28734 (N_28734,N_27106,N_26829);
nor U28735 (N_28735,N_26491,N_27495);
and U28736 (N_28736,N_27050,N_27390);
nor U28737 (N_28737,N_27497,N_27460);
and U28738 (N_28738,N_26900,N_26699);
and U28739 (N_28739,N_27002,N_26625);
and U28740 (N_28740,N_27469,N_26599);
nor U28741 (N_28741,N_27275,N_26673);
nand U28742 (N_28742,N_26791,N_27325);
and U28743 (N_28743,N_26973,N_26813);
xnor U28744 (N_28744,N_26543,N_27065);
nand U28745 (N_28745,N_27226,N_26606);
nand U28746 (N_28746,N_26737,N_26741);
nand U28747 (N_28747,N_26603,N_26517);
and U28748 (N_28748,N_27199,N_27407);
nand U28749 (N_28749,N_27111,N_26971);
and U28750 (N_28750,N_27378,N_27383);
nor U28751 (N_28751,N_27146,N_26653);
and U28752 (N_28752,N_26441,N_26656);
or U28753 (N_28753,N_26860,N_27000);
nand U28754 (N_28754,N_26584,N_27309);
xnor U28755 (N_28755,N_27229,N_26561);
xor U28756 (N_28756,N_27187,N_27482);
or U28757 (N_28757,N_26939,N_26599);
and U28758 (N_28758,N_27339,N_26980);
and U28759 (N_28759,N_27188,N_27230);
xnor U28760 (N_28760,N_27403,N_27529);
nor U28761 (N_28761,N_27376,N_26706);
xor U28762 (N_28762,N_27291,N_27178);
xor U28763 (N_28763,N_26434,N_26513);
xor U28764 (N_28764,N_27061,N_26665);
nand U28765 (N_28765,N_27522,N_26719);
or U28766 (N_28766,N_27113,N_26818);
or U28767 (N_28767,N_27314,N_26772);
nand U28768 (N_28768,N_27494,N_27015);
nand U28769 (N_28769,N_26982,N_26661);
nand U28770 (N_28770,N_27052,N_26564);
xor U28771 (N_28771,N_26545,N_26832);
nand U28772 (N_28772,N_26551,N_27105);
xnor U28773 (N_28773,N_27429,N_26592);
nand U28774 (N_28774,N_26956,N_27266);
and U28775 (N_28775,N_27286,N_27098);
xor U28776 (N_28776,N_27297,N_27154);
xnor U28777 (N_28777,N_27204,N_26753);
nor U28778 (N_28778,N_26588,N_26554);
nand U28779 (N_28779,N_26634,N_26847);
xnor U28780 (N_28780,N_27569,N_27414);
or U28781 (N_28781,N_26849,N_26564);
and U28782 (N_28782,N_27429,N_27426);
nor U28783 (N_28783,N_26675,N_27121);
xnor U28784 (N_28784,N_27524,N_27297);
or U28785 (N_28785,N_26744,N_26866);
and U28786 (N_28786,N_27439,N_27113);
xor U28787 (N_28787,N_27428,N_26946);
or U28788 (N_28788,N_27206,N_27250);
and U28789 (N_28789,N_26772,N_26988);
and U28790 (N_28790,N_26743,N_27576);
nand U28791 (N_28791,N_27415,N_26462);
and U28792 (N_28792,N_26893,N_27118);
nand U28793 (N_28793,N_27321,N_27277);
and U28794 (N_28794,N_27325,N_26401);
nand U28795 (N_28795,N_26470,N_26581);
nor U28796 (N_28796,N_26665,N_26487);
or U28797 (N_28797,N_27198,N_26837);
nand U28798 (N_28798,N_27532,N_26690);
or U28799 (N_28799,N_26457,N_26911);
nor U28800 (N_28800,N_28381,N_27702);
nor U28801 (N_28801,N_28171,N_28305);
and U28802 (N_28802,N_28391,N_28474);
xnor U28803 (N_28803,N_28257,N_28253);
or U28804 (N_28804,N_27777,N_27878);
nand U28805 (N_28805,N_27742,N_28691);
nor U28806 (N_28806,N_28520,N_28266);
xnor U28807 (N_28807,N_28028,N_28345);
or U28808 (N_28808,N_28692,N_28259);
nand U28809 (N_28809,N_28762,N_27866);
xor U28810 (N_28810,N_28160,N_27674);
nand U28811 (N_28811,N_28516,N_28733);
xor U28812 (N_28812,N_28047,N_27851);
xor U28813 (N_28813,N_28610,N_28006);
nor U28814 (N_28814,N_28270,N_28038);
xor U28815 (N_28815,N_28103,N_28225);
nor U28816 (N_28816,N_27741,N_27633);
and U28817 (N_28817,N_27672,N_28036);
or U28818 (N_28818,N_28050,N_28098);
or U28819 (N_28819,N_28764,N_28600);
nand U28820 (N_28820,N_28793,N_28153);
nor U28821 (N_28821,N_28644,N_28426);
nand U28822 (N_28822,N_28642,N_28236);
xor U28823 (N_28823,N_27649,N_28330);
nor U28824 (N_28824,N_28455,N_27669);
xor U28825 (N_28825,N_28732,N_28629);
nand U28826 (N_28826,N_27729,N_28687);
xor U28827 (N_28827,N_28163,N_28138);
nand U28828 (N_28828,N_27626,N_27725);
nor U28829 (N_28829,N_28658,N_27604);
nor U28830 (N_28830,N_28507,N_28382);
or U28831 (N_28831,N_28641,N_28140);
nand U28832 (N_28832,N_27969,N_27852);
nand U28833 (N_28833,N_28619,N_27648);
or U28834 (N_28834,N_28054,N_28191);
and U28835 (N_28835,N_27930,N_28473);
and U28836 (N_28836,N_28135,N_27752);
nor U28837 (N_28837,N_28745,N_28718);
or U28838 (N_28838,N_28194,N_28134);
xnor U28839 (N_28839,N_28375,N_27620);
nor U28840 (N_28840,N_28144,N_27917);
nand U28841 (N_28841,N_28433,N_28374);
nand U28842 (N_28842,N_28483,N_28504);
or U28843 (N_28843,N_27635,N_27801);
and U28844 (N_28844,N_28099,N_28190);
xor U28845 (N_28845,N_27877,N_28210);
and U28846 (N_28846,N_27952,N_27910);
xor U28847 (N_28847,N_27692,N_28187);
or U28848 (N_28848,N_28148,N_28450);
and U28849 (N_28849,N_28434,N_28274);
or U28850 (N_28850,N_28636,N_28445);
nor U28851 (N_28851,N_28268,N_28113);
nand U28852 (N_28852,N_27935,N_28120);
or U28853 (N_28853,N_28747,N_28016);
or U28854 (N_28854,N_27730,N_28765);
and U28855 (N_28855,N_28324,N_28627);
xor U28856 (N_28856,N_28093,N_28638);
xor U28857 (N_28857,N_28751,N_28515);
nor U28858 (N_28858,N_28682,N_28186);
xnor U28859 (N_28859,N_28218,N_27748);
and U28860 (N_28860,N_27639,N_28416);
or U28861 (N_28861,N_27815,N_28693);
nand U28862 (N_28862,N_28769,N_28238);
nand U28863 (N_28863,N_28774,N_28372);
xor U28864 (N_28864,N_27764,N_28609);
or U28865 (N_28865,N_28403,N_27734);
or U28866 (N_28866,N_28606,N_28326);
nor U28867 (N_28867,N_28396,N_28503);
or U28868 (N_28868,N_28311,N_28332);
nand U28869 (N_28869,N_28487,N_27846);
xnor U28870 (N_28870,N_28199,N_28249);
and U28871 (N_28871,N_27960,N_28552);
nor U28872 (N_28872,N_28481,N_28791);
or U28873 (N_28873,N_28536,N_27860);
and U28874 (N_28874,N_27782,N_28652);
nand U28875 (N_28875,N_27731,N_28735);
nor U28876 (N_28876,N_28502,N_27803);
or U28877 (N_28877,N_28369,N_27636);
nor U28878 (N_28878,N_28159,N_27873);
nand U28879 (N_28879,N_28079,N_27942);
xor U28880 (N_28880,N_27956,N_28157);
nand U28881 (N_28881,N_28308,N_28221);
or U28882 (N_28882,N_28757,N_27733);
nand U28883 (N_28883,N_28457,N_28530);
or U28884 (N_28884,N_28383,N_28040);
or U28885 (N_28885,N_28023,N_28674);
and U28886 (N_28886,N_27656,N_27971);
and U28887 (N_28887,N_27855,N_28621);
xnor U28888 (N_28888,N_28413,N_27607);
xnor U28889 (N_28889,N_27915,N_27948);
or U28890 (N_28890,N_28598,N_28165);
nand U28891 (N_28891,N_27710,N_27651);
or U28892 (N_28892,N_28067,N_27659);
or U28893 (N_28893,N_28032,N_28560);
nor U28894 (N_28894,N_28522,N_28243);
xor U28895 (N_28895,N_28068,N_28545);
and U28896 (N_28896,N_28725,N_28360);
or U28897 (N_28897,N_28525,N_28586);
xnor U28898 (N_28898,N_28130,N_27601);
or U28899 (N_28899,N_28405,N_28783);
nor U28900 (N_28900,N_28280,N_28364);
and U28901 (N_28901,N_28367,N_28297);
nand U28902 (N_28902,N_28690,N_27757);
and U28903 (N_28903,N_27695,N_28009);
nand U28904 (N_28904,N_28262,N_28740);
xor U28905 (N_28905,N_27914,N_28484);
and U28906 (N_28906,N_28203,N_27632);
and U28907 (N_28907,N_28538,N_28623);
or U28908 (N_28908,N_27883,N_28409);
or U28909 (N_28909,N_28271,N_27947);
xnor U28910 (N_28910,N_28737,N_28339);
and U28911 (N_28911,N_28529,N_28389);
xnor U28912 (N_28912,N_28703,N_28716);
xor U28913 (N_28913,N_28460,N_27617);
nor U28914 (N_28914,N_27940,N_28648);
or U28915 (N_28915,N_27623,N_27653);
and U28916 (N_28916,N_27970,N_28559);
or U28917 (N_28917,N_27839,N_28343);
xnor U28918 (N_28918,N_28787,N_27621);
nand U28919 (N_28919,N_28097,N_28561);
xnor U28920 (N_28920,N_28004,N_28059);
and U28921 (N_28921,N_28132,N_28233);
nand U28922 (N_28922,N_28161,N_27797);
nand U28923 (N_28923,N_27679,N_27629);
and U28924 (N_28924,N_27765,N_28741);
nand U28925 (N_28925,N_27658,N_28331);
nand U28926 (N_28926,N_27890,N_27637);
and U28927 (N_28927,N_27657,N_28288);
nand U28928 (N_28928,N_28125,N_28178);
xnor U28929 (N_28929,N_28301,N_27834);
nor U28930 (N_28930,N_28707,N_28075);
and U28931 (N_28931,N_28258,N_28250);
xor U28932 (N_28932,N_28334,N_27755);
or U28933 (N_28933,N_28353,N_28151);
xnor U28934 (N_28934,N_28645,N_28408);
and U28935 (N_28935,N_28709,N_28498);
xnor U28936 (N_28936,N_28406,N_27600);
and U28937 (N_28937,N_27724,N_28094);
and U28938 (N_28938,N_28282,N_27787);
and U28939 (N_28939,N_28518,N_27966);
or U28940 (N_28940,N_28084,N_27732);
xnor U28941 (N_28941,N_28688,N_28281);
nand U28942 (N_28942,N_27753,N_28251);
nor U28943 (N_28943,N_28149,N_28051);
xor U28944 (N_28944,N_28037,N_27831);
nor U28945 (N_28945,N_28117,N_27697);
xnor U28946 (N_28946,N_27962,N_28048);
nor U28947 (N_28947,N_28657,N_28625);
or U28948 (N_28948,N_27916,N_28778);
nand U28949 (N_28949,N_27677,N_27832);
xor U28950 (N_28950,N_27664,N_28476);
xor U28951 (N_28951,N_28168,N_28497);
xor U28952 (N_28952,N_28670,N_28611);
nor U28953 (N_28953,N_28749,N_28506);
nor U28954 (N_28954,N_28797,N_28284);
nor U28955 (N_28955,N_28392,N_28286);
xnor U28956 (N_28956,N_27631,N_27896);
xor U28957 (N_28957,N_28724,N_28323);
nor U28958 (N_28958,N_27663,N_28466);
nand U28959 (N_28959,N_28775,N_27811);
nand U28960 (N_28960,N_27728,N_28315);
nand U28961 (N_28961,N_28482,N_28567);
or U28962 (N_28962,N_28356,N_28034);
xor U28963 (N_28963,N_28422,N_28010);
nand U28964 (N_28964,N_27726,N_28240);
or U28965 (N_28965,N_28124,N_28541);
nor U28966 (N_28966,N_28340,N_28206);
nor U28967 (N_28967,N_28208,N_28336);
and U28968 (N_28968,N_27876,N_28526);
or U28969 (N_28969,N_28033,N_28255);
xor U28970 (N_28970,N_27938,N_27684);
and U28971 (N_28971,N_27903,N_27954);
and U28972 (N_28972,N_28485,N_27976);
or U28973 (N_28973,N_27762,N_28451);
and U28974 (N_28974,N_27837,N_28175);
or U28975 (N_28975,N_27880,N_28402);
nor U28976 (N_28976,N_28070,N_28316);
and U28977 (N_28977,N_28685,N_28746);
nor U28978 (N_28978,N_28260,N_28277);
nand U28979 (N_28979,N_28376,N_28302);
nor U28980 (N_28980,N_27776,N_28204);
or U28981 (N_28981,N_27875,N_28357);
nor U28982 (N_28982,N_27849,N_28349);
xor U28983 (N_28983,N_28794,N_27665);
nand U28984 (N_28984,N_28342,N_28509);
nand U28985 (N_28985,N_28112,N_28407);
nor U28986 (N_28986,N_28300,N_27967);
nand U28987 (N_28987,N_27871,N_28573);
or U28988 (N_28988,N_28201,N_28501);
nor U28989 (N_28989,N_28404,N_28579);
nor U28990 (N_28990,N_28779,N_27993);
nor U28991 (N_28991,N_28026,N_28440);
and U28992 (N_28992,N_28617,N_28314);
xnor U28993 (N_28993,N_27708,N_27820);
nand U28994 (N_28994,N_27887,N_28744);
nand U28995 (N_28995,N_28275,N_28361);
and U28996 (N_28996,N_28246,N_28133);
and U28997 (N_28997,N_28758,N_27608);
nor U28998 (N_28998,N_28431,N_27937);
or U28999 (N_28999,N_28058,N_27908);
and U29000 (N_29000,N_28592,N_27686);
and U29001 (N_29001,N_27721,N_28256);
or U29002 (N_29002,N_28563,N_28756);
or U29003 (N_29003,N_27783,N_27840);
nor U29004 (N_29004,N_28123,N_28524);
or U29005 (N_29005,N_28574,N_28283);
nand U29006 (N_29006,N_28790,N_27859);
and U29007 (N_29007,N_27619,N_28583);
nor U29008 (N_29008,N_28667,N_27602);
or U29009 (N_29009,N_28180,N_28550);
nand U29010 (N_29010,N_28072,N_28215);
xor U29011 (N_29011,N_27616,N_28773);
xor U29012 (N_29012,N_28569,N_27768);
or U29013 (N_29013,N_28661,N_27992);
xor U29014 (N_29014,N_28479,N_28193);
nand U29015 (N_29015,N_28777,N_28046);
or U29016 (N_29016,N_27805,N_28363);
and U29017 (N_29017,N_28115,N_28705);
xor U29018 (N_29018,N_27614,N_28102);
nor U29019 (N_29019,N_27893,N_28386);
xnor U29020 (N_29020,N_28615,N_27863);
nor U29021 (N_29021,N_28796,N_28772);
xor U29022 (N_29022,N_28664,N_28443);
nor U29023 (N_29023,N_28141,N_28517);
and U29024 (N_29024,N_27701,N_28385);
or U29025 (N_29025,N_28337,N_27668);
nand U29026 (N_29026,N_28241,N_28585);
nor U29027 (N_29027,N_27769,N_27738);
or U29028 (N_29028,N_28729,N_28365);
xor U29029 (N_29029,N_28448,N_28220);
or U29030 (N_29030,N_27899,N_28304);
nand U29031 (N_29031,N_27911,N_28587);
and U29032 (N_29032,N_28207,N_28454);
nand U29033 (N_29033,N_28211,N_27838);
and U29034 (N_29034,N_28182,N_28197);
and U29035 (N_29035,N_28090,N_28557);
and U29036 (N_29036,N_27913,N_28647);
xor U29037 (N_29037,N_27789,N_28303);
and U29038 (N_29038,N_28734,N_28662);
and U29039 (N_29039,N_28338,N_28209);
nor U29040 (N_29040,N_28083,N_27982);
nor U29041 (N_29041,N_28398,N_27628);
or U29042 (N_29042,N_28119,N_27881);
nand U29043 (N_29043,N_28717,N_27958);
xnor U29044 (N_29044,N_28095,N_28379);
and U29045 (N_29045,N_27988,N_28571);
nand U29046 (N_29046,N_28154,N_28435);
xor U29047 (N_29047,N_28462,N_28432);
nand U29048 (N_29048,N_28671,N_28137);
nor U29049 (N_29049,N_28789,N_28499);
nand U29050 (N_29050,N_27955,N_28291);
xnor U29051 (N_29051,N_27950,N_27968);
nand U29052 (N_29052,N_28798,N_28697);
xor U29053 (N_29053,N_27822,N_28387);
nor U29054 (N_29054,N_27879,N_27712);
xor U29055 (N_29055,N_27870,N_28676);
and U29056 (N_29056,N_28728,N_28767);
and U29057 (N_29057,N_28755,N_28085);
and U29058 (N_29058,N_27898,N_28738);
nand U29059 (N_29059,N_27704,N_27907);
xor U29060 (N_29060,N_28468,N_28665);
nor U29061 (N_29061,N_27977,N_27606);
and U29062 (N_29062,N_27722,N_27909);
nor U29063 (N_29063,N_28106,N_27858);
and U29064 (N_29064,N_28295,N_28643);
xnor U29065 (N_29065,N_28593,N_28198);
nor U29066 (N_29066,N_28071,N_28306);
and U29067 (N_29067,N_28227,N_27756);
and U29068 (N_29068,N_28702,N_27798);
nor U29069 (N_29069,N_27990,N_27941);
xnor U29070 (N_29070,N_28254,N_27716);
or U29071 (N_29071,N_27793,N_28490);
xor U29072 (N_29072,N_27747,N_27847);
nor U29073 (N_29073,N_28030,N_28176);
and U29074 (N_29074,N_28589,N_28022);
and U29075 (N_29075,N_27804,N_27646);
and U29076 (N_29076,N_27799,N_28213);
xor U29077 (N_29077,N_28118,N_28710);
and U29078 (N_29078,N_28390,N_28293);
nor U29079 (N_29079,N_28354,N_28017);
xnor U29080 (N_29080,N_27605,N_27854);
nor U29081 (N_29081,N_28588,N_27882);
and U29082 (N_29082,N_28465,N_28065);
or U29083 (N_29083,N_27688,N_28668);
nand U29084 (N_29084,N_27760,N_28761);
nor U29085 (N_29085,N_28640,N_28519);
and U29086 (N_29086,N_28469,N_28351);
nor U29087 (N_29087,N_28162,N_27671);
or U29088 (N_29088,N_27869,N_27933);
and U29089 (N_29089,N_27979,N_27819);
and U29090 (N_29090,N_27934,N_27660);
nor U29091 (N_29091,N_27786,N_27681);
nor U29092 (N_29092,N_27778,N_28189);
nand U29093 (N_29093,N_27735,N_27624);
xor U29094 (N_29094,N_27817,N_28726);
nand U29095 (N_29095,N_28045,N_27791);
or U29096 (N_29096,N_27745,N_28247);
xor U29097 (N_29097,N_28649,N_28318);
xor U29098 (N_29098,N_27699,N_27823);
nor U29099 (N_29099,N_27641,N_27864);
nor U29100 (N_29100,N_28183,N_27743);
nand U29101 (N_29101,N_28411,N_28566);
xor U29102 (N_29102,N_28591,N_27640);
or U29103 (N_29103,N_28155,N_28152);
and U29104 (N_29104,N_27773,N_28570);
xnor U29105 (N_29105,N_27685,N_27809);
xnor U29106 (N_29106,N_28373,N_27981);
and U29107 (N_29107,N_27812,N_27824);
and U29108 (N_29108,N_28540,N_28031);
nand U29109 (N_29109,N_28771,N_28131);
or U29110 (N_29110,N_27936,N_27759);
nand U29111 (N_29111,N_28470,N_27615);
nor U29112 (N_29112,N_28229,N_27690);
and U29113 (N_29113,N_28678,N_28350);
and U29114 (N_29114,N_28601,N_28174);
or U29115 (N_29115,N_28572,N_28005);
nor U29116 (N_29116,N_28442,N_28368);
or U29117 (N_29117,N_27985,N_28359);
and U29118 (N_29118,N_28265,N_28394);
and U29119 (N_29119,N_28366,N_28002);
xnor U29120 (N_29120,N_27642,N_28602);
xor U29121 (N_29121,N_28510,N_27918);
and U29122 (N_29122,N_27670,N_28521);
xor U29123 (N_29123,N_28272,N_27997);
or U29124 (N_29124,N_28177,N_28327);
nor U29125 (N_29125,N_28508,N_28267);
and U29126 (N_29126,N_28142,N_28035);
nand U29127 (N_29127,N_28087,N_28073);
nor U29128 (N_29128,N_28397,N_28720);
nand U29129 (N_29129,N_28289,N_28076);
and U29130 (N_29130,N_28414,N_28329);
xor U29131 (N_29131,N_28616,N_28788);
and U29132 (N_29132,N_28539,N_28384);
xnor U29133 (N_29133,N_28401,N_28495);
or U29134 (N_29134,N_27766,N_28185);
nand U29135 (N_29135,N_27949,N_28212);
nand U29136 (N_29136,N_28686,N_27932);
nor U29137 (N_29137,N_28321,N_28410);
or U29138 (N_29138,N_28493,N_28049);
or U29139 (N_29139,N_28715,N_28412);
and U29140 (N_29140,N_28459,N_28164);
and U29141 (N_29141,N_28666,N_28528);
or U29142 (N_29142,N_28237,N_28532);
nand U29143 (N_29143,N_27698,N_27696);
and U29144 (N_29144,N_27654,N_27775);
and U29145 (N_29145,N_28156,N_27939);
or U29146 (N_29146,N_27666,N_28264);
or U29147 (N_29147,N_28478,N_28776);
nand U29148 (N_29148,N_28158,N_28074);
nand U29149 (N_29149,N_28000,N_28276);
nand U29150 (N_29150,N_28415,N_28461);
nand U29151 (N_29151,N_28378,N_28108);
and U29152 (N_29152,N_28655,N_28309);
or U29153 (N_29153,N_28496,N_28603);
nand U29154 (N_29154,N_28143,N_27717);
nor U29155 (N_29155,N_27998,N_28217);
and U29156 (N_29156,N_28234,N_28001);
xor U29157 (N_29157,N_28173,N_28377);
and U29158 (N_29158,N_28296,N_27715);
xnor U29159 (N_29159,N_28192,N_28635);
nand U29160 (N_29160,N_28344,N_28167);
nor U29161 (N_29161,N_28231,N_28126);
xnor U29162 (N_29162,N_28428,N_28634);
and U29163 (N_29163,N_28620,N_28341);
xor U29164 (N_29164,N_27780,N_28328);
nand U29165 (N_29165,N_28505,N_28320);
nor U29166 (N_29166,N_27807,N_28604);
or U29167 (N_29167,N_28677,N_28044);
nand U29168 (N_29168,N_27630,N_28273);
or U29169 (N_29169,N_28252,N_28056);
xor U29170 (N_29170,N_28371,N_28799);
or U29171 (N_29171,N_28639,N_27996);
nand U29172 (N_29172,N_28053,N_28078);
nor U29173 (N_29173,N_28730,N_28553);
xnor U29174 (N_29174,N_27891,N_27779);
nand U29175 (N_29175,N_28294,N_27613);
or U29176 (N_29176,N_28568,N_27689);
and U29177 (N_29177,N_27650,N_28659);
or U29178 (N_29178,N_28088,N_28679);
nand U29179 (N_29179,N_27676,N_27951);
or U29180 (N_29180,N_27711,N_28420);
xor U29181 (N_29181,N_27965,N_28695);
nand U29182 (N_29182,N_28651,N_28564);
or U29183 (N_29183,N_27785,N_28100);
or U29184 (N_29184,N_28063,N_28723);
xor U29185 (N_29185,N_28166,N_28121);
or U29186 (N_29186,N_27627,N_28024);
or U29187 (N_29187,N_27895,N_28512);
and U29188 (N_29188,N_27751,N_28731);
xor U29189 (N_29189,N_27922,N_28551);
or U29190 (N_29190,N_28456,N_27770);
nand U29191 (N_29191,N_28195,N_28543);
and U29192 (N_29192,N_27758,N_28352);
and U29193 (N_29193,N_27693,N_27995);
nand U29194 (N_29194,N_27928,N_28395);
nand U29195 (N_29195,N_28597,N_28244);
or U29196 (N_29196,N_27923,N_28109);
or U29197 (N_29197,N_28607,N_27610);
nor U29198 (N_29198,N_28711,N_28007);
and U29199 (N_29199,N_28511,N_28575);
or U29200 (N_29200,N_28494,N_28043);
and U29201 (N_29201,N_28475,N_28436);
nor U29202 (N_29202,N_28419,N_27836);
and U29203 (N_29203,N_28580,N_28599);
xnor U29204 (N_29204,N_28472,N_28292);
or U29205 (N_29205,N_28488,N_28346);
nor U29206 (N_29206,N_27667,N_28089);
and U29207 (N_29207,N_28136,N_28013);
nor U29208 (N_29208,N_27609,N_28129);
and U29209 (N_29209,N_28224,N_28681);
or U29210 (N_29210,N_28449,N_28139);
xnor U29211 (N_29211,N_28750,N_27844);
nand U29212 (N_29212,N_27975,N_28279);
or U29213 (N_29213,N_27884,N_27808);
xnor U29214 (N_29214,N_28605,N_28298);
xnor U29215 (N_29215,N_28786,N_27814);
xor U29216 (N_29216,N_28523,N_28269);
or U29217 (N_29217,N_28169,N_28424);
or U29218 (N_29218,N_28624,N_28548);
xnor U29219 (N_29219,N_27784,N_28489);
or U29220 (N_29220,N_28285,N_28722);
nor U29221 (N_29221,N_28228,N_27718);
nor U29222 (N_29222,N_27953,N_27796);
nor U29223 (N_29223,N_27921,N_28719);
xor U29224 (N_29224,N_27788,N_28347);
xnor U29225 (N_29225,N_27912,N_28618);
xnor U29226 (N_29226,N_27983,N_27974);
and U29227 (N_29227,N_27926,N_28694);
or U29228 (N_29228,N_28708,N_28578);
or U29229 (N_29229,N_27813,N_27792);
xor U29230 (N_29230,N_28425,N_28188);
and U29231 (N_29231,N_28114,N_28721);
nor U29232 (N_29232,N_27700,N_28128);
nor U29233 (N_29233,N_28242,N_28052);
nor U29234 (N_29234,N_28400,N_28760);
xor U29235 (N_29235,N_28628,N_27739);
nor U29236 (N_29236,N_28577,N_28452);
xor U29237 (N_29237,N_27959,N_27603);
and U29238 (N_29238,N_27845,N_28261);
and U29239 (N_29239,N_27647,N_28216);
nor U29240 (N_29240,N_28091,N_28654);
nand U29241 (N_29241,N_28753,N_27680);
nand U29242 (N_29242,N_28514,N_28015);
or U29243 (N_29243,N_28307,N_28727);
and U29244 (N_29244,N_28675,N_27931);
xnor U29245 (N_29245,N_28355,N_28008);
and U29246 (N_29246,N_28042,N_27767);
nand U29247 (N_29247,N_28596,N_28196);
xor U29248 (N_29248,N_27991,N_27943);
xnor U29249 (N_29249,N_28226,N_27961);
and U29250 (N_29250,N_28742,N_28312);
nand U29251 (N_29251,N_27645,N_28780);
xnor U29252 (N_29252,N_28653,N_27946);
nor U29253 (N_29253,N_27694,N_27972);
xor U29254 (N_29254,N_27625,N_27920);
nand U29255 (N_29255,N_28019,N_28427);
nand U29256 (N_29256,N_28491,N_28235);
or U29257 (N_29257,N_28322,N_28792);
and U29258 (N_29258,N_27723,N_28626);
and U29259 (N_29259,N_27963,N_28680);
nand U29260 (N_29260,N_28055,N_27737);
nand U29261 (N_29261,N_28107,N_28446);
or U29262 (N_29262,N_28146,N_27790);
nand U29263 (N_29263,N_28684,N_27714);
nor U29264 (N_29264,N_28086,N_28399);
xnor U29265 (N_29265,N_27772,N_28358);
or U29266 (N_29266,N_27740,N_27853);
nor U29267 (N_29267,N_27622,N_28531);
xor U29268 (N_29268,N_28632,N_27841);
nor U29269 (N_29269,N_27828,N_28437);
xnor U29270 (N_29270,N_28689,N_28096);
nor U29271 (N_29271,N_28062,N_27889);
xor U29272 (N_29272,N_28430,N_27806);
nor U29273 (N_29273,N_28111,N_27618);
nor U29274 (N_29274,N_28181,N_28077);
nor U29275 (N_29275,N_27774,N_28700);
and U29276 (N_29276,N_28219,N_28417);
or U29277 (N_29277,N_27888,N_28441);
or U29278 (N_29278,N_27861,N_27794);
nor U29279 (N_29279,N_27829,N_28453);
nor U29280 (N_29280,N_28663,N_28713);
nand U29281 (N_29281,N_28631,N_27925);
xnor U29282 (N_29282,N_27919,N_28477);
and U29283 (N_29283,N_27874,N_27678);
and U29284 (N_29284,N_27736,N_27986);
xnor U29285 (N_29285,N_27944,N_28438);
or U29286 (N_29286,N_28061,N_27862);
nand U29287 (N_29287,N_28544,N_28423);
nor U29288 (N_29288,N_27810,N_28782);
nand U29289 (N_29289,N_27713,N_27652);
or U29290 (N_29290,N_28057,N_27687);
nor U29291 (N_29291,N_28712,N_27857);
nand U29292 (N_29292,N_28669,N_28633);
nor U29293 (N_29293,N_28781,N_27754);
nor U29294 (N_29294,N_27833,N_28766);
nor U29295 (N_29295,N_27761,N_28060);
xnor U29296 (N_29296,N_28535,N_28554);
xor U29297 (N_29297,N_27927,N_27612);
xor U29298 (N_29298,N_28683,N_27978);
and U29299 (N_29299,N_28202,N_27843);
xor U29300 (N_29300,N_28486,N_28590);
nand U29301 (N_29301,N_27825,N_27973);
or U29302 (N_29302,N_27826,N_27661);
nand U29303 (N_29303,N_28263,N_27818);
nand U29304 (N_29304,N_28122,N_27744);
nor U29305 (N_29305,N_28595,N_27750);
nand U29306 (N_29306,N_28230,N_28739);
and U29307 (N_29307,N_28025,N_28613);
and U29308 (N_29308,N_27706,N_28020);
and U29309 (N_29309,N_28582,N_28533);
or U29310 (N_29310,N_27901,N_28795);
nand U29311 (N_29311,N_28594,N_28527);
or U29312 (N_29312,N_28278,N_28471);
xnor U29313 (N_29313,N_28222,N_28101);
nor U29314 (N_29314,N_28064,N_28418);
nor U29315 (N_29315,N_27638,N_28232);
and U29316 (N_29316,N_28500,N_27673);
and U29317 (N_29317,N_27872,N_28105);
xor U29318 (N_29318,N_28576,N_28027);
and U29319 (N_29319,N_28388,N_27980);
xor U29320 (N_29320,N_28018,N_27842);
xor U29321 (N_29321,N_28170,N_28696);
nor U29322 (N_29322,N_28082,N_28754);
xor U29323 (N_29323,N_27703,N_28698);
or U29324 (N_29324,N_28147,N_28759);
nor U29325 (N_29325,N_28714,N_27865);
nand U29326 (N_29326,N_28069,N_28248);
or U29327 (N_29327,N_27800,N_27781);
xnor U29328 (N_29328,N_28637,N_27727);
xnor U29329 (N_29329,N_27897,N_28558);
nand U29330 (N_29330,N_28701,N_28299);
and U29331 (N_29331,N_28200,N_27763);
xor U29332 (N_29332,N_27655,N_27905);
or U29333 (N_29333,N_28421,N_28110);
nand U29334 (N_29334,N_28012,N_28172);
and U29335 (N_29335,N_28319,N_27634);
nor U29336 (N_29336,N_27989,N_28584);
and U29337 (N_29337,N_28039,N_27683);
xor U29338 (N_29338,N_28770,N_28370);
nor U29339 (N_29339,N_28630,N_27987);
or U29340 (N_29340,N_28784,N_27999);
xnor U29341 (N_29341,N_28014,N_27675);
nand U29342 (N_29342,N_27848,N_28287);
nand U29343 (N_29343,N_28214,N_28179);
and U29344 (N_29344,N_28537,N_28029);
nor U29345 (N_29345,N_27611,N_28480);
nand U29346 (N_29346,N_28660,N_28116);
nor U29347 (N_29347,N_27709,N_27827);
nor U29348 (N_29348,N_27906,N_28556);
nor U29349 (N_29349,N_28393,N_28748);
xor U29350 (N_29350,N_27984,N_28362);
nand U29351 (N_29351,N_28743,N_28614);
xnor U29352 (N_29352,N_27994,N_28463);
and U29353 (N_29353,N_28581,N_28290);
xnor U29354 (N_29354,N_27821,N_28699);
nor U29355 (N_29355,N_28313,N_28223);
and U29356 (N_29356,N_27720,N_28547);
and U29357 (N_29357,N_28546,N_28239);
and U29358 (N_29358,N_27644,N_27892);
or U29359 (N_29359,N_28380,N_27749);
xor U29360 (N_29360,N_27945,N_27830);
nand U29361 (N_29361,N_28534,N_28317);
or U29362 (N_29362,N_27816,N_28672);
nand U29363 (N_29363,N_28562,N_27707);
or U29364 (N_29364,N_28081,N_28447);
and U29365 (N_29365,N_27719,N_27662);
nor U29366 (N_29366,N_28763,N_28325);
and U29367 (N_29367,N_28565,N_28003);
xnor U29368 (N_29368,N_27886,N_27856);
nand U29369 (N_29369,N_28444,N_28145);
xnor U29370 (N_29370,N_28768,N_28092);
or U29371 (N_29371,N_28704,N_28184);
and U29372 (N_29372,N_27868,N_28333);
or U29373 (N_29373,N_28335,N_27682);
or U29374 (N_29374,N_28439,N_27867);
nand U29375 (N_29375,N_27894,N_27902);
or U29376 (N_29376,N_27705,N_28011);
nand U29377 (N_29377,N_27795,N_28612);
nand U29378 (N_29378,N_28785,N_28080);
nor U29379 (N_29379,N_28513,N_28752);
and U29380 (N_29380,N_27964,N_27771);
nand U29381 (N_29381,N_27850,N_28673);
xor U29382 (N_29382,N_28706,N_28646);
nand U29383 (N_29383,N_28656,N_28021);
xnor U29384 (N_29384,N_27904,N_28736);
and U29385 (N_29385,N_27835,N_27957);
nand U29386 (N_29386,N_28464,N_27885);
xor U29387 (N_29387,N_27929,N_27691);
xnor U29388 (N_29388,N_28492,N_28555);
nor U29389 (N_29389,N_28041,N_27802);
and U29390 (N_29390,N_28310,N_28608);
or U29391 (N_29391,N_28104,N_28429);
and U29392 (N_29392,N_28622,N_28650);
xor U29393 (N_29393,N_27643,N_28348);
and U29394 (N_29394,N_27746,N_28066);
xnor U29395 (N_29395,N_27924,N_28127);
and U29396 (N_29396,N_28245,N_28150);
and U29397 (N_29397,N_28549,N_28458);
or U29398 (N_29398,N_28205,N_28542);
or U29399 (N_29399,N_28467,N_27900);
nand U29400 (N_29400,N_27664,N_27903);
nor U29401 (N_29401,N_28338,N_27970);
nor U29402 (N_29402,N_28132,N_27690);
and U29403 (N_29403,N_28397,N_27711);
or U29404 (N_29404,N_27813,N_28622);
nor U29405 (N_29405,N_27834,N_28117);
and U29406 (N_29406,N_27994,N_28052);
xnor U29407 (N_29407,N_27991,N_27767);
nor U29408 (N_29408,N_28014,N_28207);
nor U29409 (N_29409,N_27959,N_27621);
or U29410 (N_29410,N_28488,N_28014);
xnor U29411 (N_29411,N_28131,N_28025);
nor U29412 (N_29412,N_28060,N_28608);
xor U29413 (N_29413,N_27811,N_28168);
or U29414 (N_29414,N_28192,N_28350);
nor U29415 (N_29415,N_27824,N_28451);
and U29416 (N_29416,N_27895,N_28345);
nor U29417 (N_29417,N_28114,N_27683);
or U29418 (N_29418,N_28232,N_27847);
or U29419 (N_29419,N_28498,N_28115);
or U29420 (N_29420,N_27693,N_28455);
nor U29421 (N_29421,N_28227,N_28648);
nand U29422 (N_29422,N_28722,N_27916);
nand U29423 (N_29423,N_28277,N_28160);
and U29424 (N_29424,N_28651,N_28583);
nand U29425 (N_29425,N_27644,N_28152);
or U29426 (N_29426,N_27874,N_28215);
or U29427 (N_29427,N_27917,N_27816);
xor U29428 (N_29428,N_28782,N_28526);
xnor U29429 (N_29429,N_28709,N_27885);
nor U29430 (N_29430,N_28379,N_28785);
nor U29431 (N_29431,N_28427,N_28649);
nor U29432 (N_29432,N_28483,N_27842);
and U29433 (N_29433,N_27764,N_28392);
nor U29434 (N_29434,N_28289,N_27822);
xor U29435 (N_29435,N_27824,N_28360);
nor U29436 (N_29436,N_27893,N_27817);
nor U29437 (N_29437,N_27971,N_28085);
and U29438 (N_29438,N_28096,N_28388);
nand U29439 (N_29439,N_27893,N_27874);
and U29440 (N_29440,N_28470,N_28474);
nor U29441 (N_29441,N_28378,N_28654);
nor U29442 (N_29442,N_28058,N_27701);
nor U29443 (N_29443,N_27998,N_28349);
or U29444 (N_29444,N_27954,N_27698);
nor U29445 (N_29445,N_28549,N_28445);
nand U29446 (N_29446,N_28340,N_28517);
nor U29447 (N_29447,N_28637,N_27864);
or U29448 (N_29448,N_27880,N_28515);
or U29449 (N_29449,N_28687,N_28552);
or U29450 (N_29450,N_28239,N_28321);
nand U29451 (N_29451,N_28066,N_28644);
and U29452 (N_29452,N_28435,N_28437);
nor U29453 (N_29453,N_28214,N_27938);
nand U29454 (N_29454,N_28189,N_28791);
xor U29455 (N_29455,N_27841,N_28489);
nor U29456 (N_29456,N_27958,N_27806);
nand U29457 (N_29457,N_27603,N_28518);
and U29458 (N_29458,N_28239,N_28694);
nand U29459 (N_29459,N_28564,N_28753);
xor U29460 (N_29460,N_27600,N_27837);
nor U29461 (N_29461,N_27659,N_27797);
xor U29462 (N_29462,N_28219,N_28571);
xor U29463 (N_29463,N_28317,N_27931);
nand U29464 (N_29464,N_28749,N_27857);
nand U29465 (N_29465,N_28749,N_28666);
and U29466 (N_29466,N_28150,N_28796);
nand U29467 (N_29467,N_28258,N_27627);
xnor U29468 (N_29468,N_28284,N_28376);
xnor U29469 (N_29469,N_28120,N_28337);
xor U29470 (N_29470,N_28132,N_28343);
xnor U29471 (N_29471,N_28373,N_27830);
nor U29472 (N_29472,N_28311,N_27860);
or U29473 (N_29473,N_27806,N_28319);
nor U29474 (N_29474,N_28633,N_28405);
xnor U29475 (N_29475,N_27924,N_28089);
or U29476 (N_29476,N_27603,N_28574);
xnor U29477 (N_29477,N_28022,N_28762);
nand U29478 (N_29478,N_28218,N_28783);
and U29479 (N_29479,N_28297,N_28788);
xor U29480 (N_29480,N_28540,N_28590);
nor U29481 (N_29481,N_28510,N_27789);
or U29482 (N_29482,N_28249,N_27860);
nand U29483 (N_29483,N_28131,N_28384);
or U29484 (N_29484,N_28184,N_28372);
or U29485 (N_29485,N_28575,N_28447);
nand U29486 (N_29486,N_28694,N_28121);
or U29487 (N_29487,N_27751,N_28070);
or U29488 (N_29488,N_27659,N_28043);
and U29489 (N_29489,N_28430,N_28635);
xor U29490 (N_29490,N_28686,N_27827);
xnor U29491 (N_29491,N_28528,N_27645);
and U29492 (N_29492,N_27725,N_28051);
nand U29493 (N_29493,N_28792,N_28552);
or U29494 (N_29494,N_28335,N_27673);
xnor U29495 (N_29495,N_27972,N_28321);
and U29496 (N_29496,N_28406,N_28157);
or U29497 (N_29497,N_28128,N_28616);
xor U29498 (N_29498,N_27687,N_28204);
nor U29499 (N_29499,N_28142,N_27675);
and U29500 (N_29500,N_28580,N_28796);
nor U29501 (N_29501,N_28286,N_28030);
and U29502 (N_29502,N_27865,N_28323);
xnor U29503 (N_29503,N_28008,N_27727);
xor U29504 (N_29504,N_27720,N_28673);
and U29505 (N_29505,N_28044,N_28421);
or U29506 (N_29506,N_28668,N_27619);
nor U29507 (N_29507,N_28590,N_28279);
and U29508 (N_29508,N_28541,N_27663);
xnor U29509 (N_29509,N_28021,N_28699);
and U29510 (N_29510,N_28575,N_27654);
nor U29511 (N_29511,N_28404,N_28784);
nor U29512 (N_29512,N_27600,N_28090);
nor U29513 (N_29513,N_28394,N_28589);
and U29514 (N_29514,N_28217,N_27702);
and U29515 (N_29515,N_28592,N_28698);
and U29516 (N_29516,N_28699,N_28301);
and U29517 (N_29517,N_28586,N_27674);
and U29518 (N_29518,N_28672,N_28654);
xor U29519 (N_29519,N_28192,N_28093);
xnor U29520 (N_29520,N_28527,N_28679);
nand U29521 (N_29521,N_28575,N_27874);
nor U29522 (N_29522,N_27958,N_28467);
and U29523 (N_29523,N_28416,N_28399);
and U29524 (N_29524,N_27863,N_27773);
nand U29525 (N_29525,N_28000,N_28365);
or U29526 (N_29526,N_28489,N_27655);
or U29527 (N_29527,N_27921,N_28021);
and U29528 (N_29528,N_28700,N_27923);
nand U29529 (N_29529,N_28118,N_27620);
xor U29530 (N_29530,N_28166,N_28242);
nand U29531 (N_29531,N_27909,N_27988);
or U29532 (N_29532,N_28251,N_28348);
nand U29533 (N_29533,N_27749,N_28136);
and U29534 (N_29534,N_28630,N_27874);
nand U29535 (N_29535,N_28556,N_27778);
xor U29536 (N_29536,N_27820,N_28107);
or U29537 (N_29537,N_27928,N_28526);
xor U29538 (N_29538,N_28772,N_27633);
or U29539 (N_29539,N_27848,N_27705);
nor U29540 (N_29540,N_27841,N_28309);
or U29541 (N_29541,N_27873,N_28208);
nor U29542 (N_29542,N_28128,N_28038);
nand U29543 (N_29543,N_28418,N_28225);
or U29544 (N_29544,N_28225,N_28271);
and U29545 (N_29545,N_27777,N_28207);
and U29546 (N_29546,N_28711,N_28610);
nand U29547 (N_29547,N_28120,N_27954);
or U29548 (N_29548,N_27986,N_27797);
nor U29549 (N_29549,N_28744,N_28707);
nand U29550 (N_29550,N_28644,N_28083);
xor U29551 (N_29551,N_28701,N_28565);
nand U29552 (N_29552,N_28646,N_28007);
or U29553 (N_29553,N_28546,N_28370);
nand U29554 (N_29554,N_28486,N_28548);
nand U29555 (N_29555,N_28563,N_28668);
xor U29556 (N_29556,N_27863,N_27618);
and U29557 (N_29557,N_28404,N_27866);
and U29558 (N_29558,N_28267,N_27986);
and U29559 (N_29559,N_27868,N_27779);
nor U29560 (N_29560,N_28244,N_27834);
or U29561 (N_29561,N_28356,N_28186);
or U29562 (N_29562,N_28142,N_28385);
nor U29563 (N_29563,N_28392,N_28353);
nor U29564 (N_29564,N_27665,N_27993);
nor U29565 (N_29565,N_28385,N_27867);
and U29566 (N_29566,N_27754,N_28666);
xor U29567 (N_29567,N_27652,N_28423);
nand U29568 (N_29568,N_28491,N_27634);
nor U29569 (N_29569,N_27701,N_27885);
or U29570 (N_29570,N_27660,N_28750);
and U29571 (N_29571,N_28447,N_28778);
nor U29572 (N_29572,N_27620,N_28363);
and U29573 (N_29573,N_28329,N_27953);
nor U29574 (N_29574,N_28326,N_27791);
and U29575 (N_29575,N_28289,N_28402);
xor U29576 (N_29576,N_27918,N_27654);
and U29577 (N_29577,N_28035,N_27836);
or U29578 (N_29578,N_28748,N_28147);
nor U29579 (N_29579,N_27678,N_28444);
or U29580 (N_29580,N_28527,N_28603);
or U29581 (N_29581,N_28664,N_28190);
and U29582 (N_29582,N_28472,N_28463);
and U29583 (N_29583,N_27887,N_28096);
nor U29584 (N_29584,N_28568,N_27983);
and U29585 (N_29585,N_27739,N_27627);
nand U29586 (N_29586,N_28322,N_27756);
xor U29587 (N_29587,N_27918,N_27695);
and U29588 (N_29588,N_28263,N_28646);
xor U29589 (N_29589,N_28673,N_28181);
or U29590 (N_29590,N_28405,N_28147);
or U29591 (N_29591,N_28089,N_28565);
or U29592 (N_29592,N_28150,N_27964);
xnor U29593 (N_29593,N_28710,N_28188);
nand U29594 (N_29594,N_28066,N_28491);
nor U29595 (N_29595,N_28676,N_28674);
xnor U29596 (N_29596,N_27724,N_28159);
and U29597 (N_29597,N_28404,N_28659);
or U29598 (N_29598,N_28232,N_28510);
xor U29599 (N_29599,N_27633,N_28783);
and U29600 (N_29600,N_28317,N_27701);
nand U29601 (N_29601,N_28275,N_27632);
nor U29602 (N_29602,N_28041,N_28437);
nor U29603 (N_29603,N_28318,N_28588);
or U29604 (N_29604,N_27913,N_28053);
xnor U29605 (N_29605,N_28505,N_27939);
nand U29606 (N_29606,N_27905,N_28714);
nor U29607 (N_29607,N_28225,N_28510);
nor U29608 (N_29608,N_28689,N_27927);
xnor U29609 (N_29609,N_28249,N_28132);
nor U29610 (N_29610,N_28362,N_28384);
or U29611 (N_29611,N_28265,N_28506);
and U29612 (N_29612,N_28429,N_27896);
or U29613 (N_29613,N_27689,N_27758);
nand U29614 (N_29614,N_28438,N_27868);
xor U29615 (N_29615,N_28433,N_28544);
nor U29616 (N_29616,N_28543,N_28428);
nor U29617 (N_29617,N_27969,N_28053);
xnor U29618 (N_29618,N_28336,N_28070);
nor U29619 (N_29619,N_27690,N_28540);
nor U29620 (N_29620,N_28637,N_28081);
xnor U29621 (N_29621,N_27826,N_28300);
xnor U29622 (N_29622,N_27789,N_27672);
nand U29623 (N_29623,N_28200,N_28351);
nor U29624 (N_29624,N_28152,N_27885);
or U29625 (N_29625,N_27701,N_27896);
and U29626 (N_29626,N_28647,N_28190);
xnor U29627 (N_29627,N_28184,N_28498);
or U29628 (N_29628,N_27722,N_27824);
and U29629 (N_29629,N_28100,N_28330);
and U29630 (N_29630,N_27950,N_28454);
nor U29631 (N_29631,N_28164,N_28662);
nand U29632 (N_29632,N_28777,N_27910);
and U29633 (N_29633,N_27861,N_27955);
nand U29634 (N_29634,N_28205,N_28350);
xnor U29635 (N_29635,N_27889,N_28109);
and U29636 (N_29636,N_28363,N_27884);
nor U29637 (N_29637,N_27956,N_27744);
nand U29638 (N_29638,N_28427,N_28426);
xor U29639 (N_29639,N_28285,N_28433);
nor U29640 (N_29640,N_27743,N_28591);
xnor U29641 (N_29641,N_28000,N_27815);
xor U29642 (N_29642,N_28549,N_28213);
nor U29643 (N_29643,N_28618,N_28666);
nor U29644 (N_29644,N_27643,N_28577);
and U29645 (N_29645,N_28144,N_28559);
and U29646 (N_29646,N_28502,N_28551);
xor U29647 (N_29647,N_28602,N_27963);
or U29648 (N_29648,N_28608,N_28666);
xor U29649 (N_29649,N_27954,N_28095);
xnor U29650 (N_29650,N_27824,N_28453);
xor U29651 (N_29651,N_27665,N_27916);
nor U29652 (N_29652,N_28014,N_28326);
nor U29653 (N_29653,N_28126,N_27726);
nor U29654 (N_29654,N_28779,N_28711);
nand U29655 (N_29655,N_27954,N_28065);
xnor U29656 (N_29656,N_28012,N_27854);
xnor U29657 (N_29657,N_27874,N_28657);
and U29658 (N_29658,N_27912,N_27856);
nor U29659 (N_29659,N_28562,N_28232);
and U29660 (N_29660,N_27780,N_27798);
nand U29661 (N_29661,N_27877,N_28001);
or U29662 (N_29662,N_27648,N_28356);
nor U29663 (N_29663,N_28423,N_28362);
nor U29664 (N_29664,N_28180,N_27804);
and U29665 (N_29665,N_27897,N_28412);
or U29666 (N_29666,N_28639,N_27686);
and U29667 (N_29667,N_28741,N_28716);
and U29668 (N_29668,N_28310,N_27681);
and U29669 (N_29669,N_28422,N_27926);
or U29670 (N_29670,N_28100,N_28704);
xor U29671 (N_29671,N_28531,N_27908);
xnor U29672 (N_29672,N_28535,N_27695);
and U29673 (N_29673,N_27751,N_28620);
or U29674 (N_29674,N_28325,N_28334);
nand U29675 (N_29675,N_28121,N_27667);
nor U29676 (N_29676,N_28747,N_28543);
and U29677 (N_29677,N_28226,N_27976);
nand U29678 (N_29678,N_28740,N_28434);
nor U29679 (N_29679,N_28008,N_28614);
or U29680 (N_29680,N_28504,N_28358);
xor U29681 (N_29681,N_28057,N_27847);
nand U29682 (N_29682,N_28576,N_27837);
nor U29683 (N_29683,N_28103,N_27713);
nor U29684 (N_29684,N_28610,N_28199);
xnor U29685 (N_29685,N_28435,N_28579);
or U29686 (N_29686,N_28541,N_28384);
and U29687 (N_29687,N_28730,N_28021);
nor U29688 (N_29688,N_27742,N_27664);
xor U29689 (N_29689,N_28102,N_27948);
or U29690 (N_29690,N_28588,N_28277);
nor U29691 (N_29691,N_28060,N_28729);
nor U29692 (N_29692,N_27713,N_28720);
nor U29693 (N_29693,N_28541,N_28583);
xnor U29694 (N_29694,N_28594,N_27883);
and U29695 (N_29695,N_27751,N_28211);
nand U29696 (N_29696,N_27970,N_27736);
and U29697 (N_29697,N_28073,N_27693);
or U29698 (N_29698,N_28709,N_28079);
and U29699 (N_29699,N_28213,N_28359);
xor U29700 (N_29700,N_27714,N_28412);
nand U29701 (N_29701,N_28110,N_28624);
xnor U29702 (N_29702,N_28604,N_27977);
or U29703 (N_29703,N_27603,N_28013);
xor U29704 (N_29704,N_28791,N_27892);
xor U29705 (N_29705,N_27923,N_28162);
or U29706 (N_29706,N_28426,N_28078);
nand U29707 (N_29707,N_28386,N_28521);
nor U29708 (N_29708,N_28234,N_28128);
and U29709 (N_29709,N_28053,N_27894);
nand U29710 (N_29710,N_27930,N_27612);
nand U29711 (N_29711,N_28218,N_27878);
or U29712 (N_29712,N_28742,N_28140);
nor U29713 (N_29713,N_27793,N_28555);
nand U29714 (N_29714,N_28718,N_27634);
xor U29715 (N_29715,N_27804,N_27744);
or U29716 (N_29716,N_28694,N_28579);
and U29717 (N_29717,N_27960,N_28228);
and U29718 (N_29718,N_28295,N_27637);
or U29719 (N_29719,N_28645,N_28541);
or U29720 (N_29720,N_27706,N_28652);
xor U29721 (N_29721,N_27724,N_28572);
nor U29722 (N_29722,N_27901,N_28225);
and U29723 (N_29723,N_27808,N_28397);
xor U29724 (N_29724,N_27835,N_27998);
xnor U29725 (N_29725,N_28273,N_27792);
nand U29726 (N_29726,N_28262,N_28180);
or U29727 (N_29727,N_28677,N_28249);
or U29728 (N_29728,N_28108,N_27953);
nor U29729 (N_29729,N_28655,N_27816);
nand U29730 (N_29730,N_27879,N_27873);
nand U29731 (N_29731,N_27786,N_28003);
and U29732 (N_29732,N_28422,N_27628);
nand U29733 (N_29733,N_28015,N_28281);
nor U29734 (N_29734,N_27952,N_28243);
nand U29735 (N_29735,N_27846,N_28777);
nor U29736 (N_29736,N_27697,N_27972);
or U29737 (N_29737,N_27947,N_28704);
nor U29738 (N_29738,N_27860,N_27655);
xor U29739 (N_29739,N_28065,N_27860);
or U29740 (N_29740,N_27749,N_27965);
or U29741 (N_29741,N_27849,N_27798);
and U29742 (N_29742,N_28228,N_28734);
nor U29743 (N_29743,N_27919,N_28573);
and U29744 (N_29744,N_28368,N_28555);
and U29745 (N_29745,N_27724,N_28362);
nand U29746 (N_29746,N_28097,N_27921);
and U29747 (N_29747,N_28445,N_27870);
xor U29748 (N_29748,N_27641,N_27948);
nand U29749 (N_29749,N_27695,N_28350);
xnor U29750 (N_29750,N_28711,N_28359);
xnor U29751 (N_29751,N_27892,N_28030);
nor U29752 (N_29752,N_28425,N_27795);
nand U29753 (N_29753,N_28097,N_27779);
nand U29754 (N_29754,N_27676,N_28715);
nand U29755 (N_29755,N_27869,N_28546);
or U29756 (N_29756,N_27667,N_28238);
nand U29757 (N_29757,N_27756,N_28299);
and U29758 (N_29758,N_27883,N_28210);
nor U29759 (N_29759,N_28110,N_28738);
and U29760 (N_29760,N_27651,N_27777);
nand U29761 (N_29761,N_28224,N_27751);
and U29762 (N_29762,N_27615,N_27998);
nand U29763 (N_29763,N_28353,N_28756);
and U29764 (N_29764,N_27703,N_28223);
xnor U29765 (N_29765,N_28488,N_27874);
nand U29766 (N_29766,N_28639,N_28431);
or U29767 (N_29767,N_27700,N_28327);
or U29768 (N_29768,N_27957,N_28578);
and U29769 (N_29769,N_28390,N_27908);
xor U29770 (N_29770,N_28664,N_28740);
nand U29771 (N_29771,N_27965,N_28782);
nand U29772 (N_29772,N_27910,N_27694);
nand U29773 (N_29773,N_28597,N_28207);
and U29774 (N_29774,N_27894,N_27702);
and U29775 (N_29775,N_28648,N_27636);
nand U29776 (N_29776,N_28272,N_28725);
nand U29777 (N_29777,N_28176,N_28209);
xnor U29778 (N_29778,N_28410,N_28123);
nor U29779 (N_29779,N_28400,N_27775);
nor U29780 (N_29780,N_28552,N_28455);
or U29781 (N_29781,N_28194,N_28652);
or U29782 (N_29782,N_28027,N_27902);
nor U29783 (N_29783,N_28184,N_27808);
or U29784 (N_29784,N_27851,N_28322);
and U29785 (N_29785,N_28567,N_28223);
xor U29786 (N_29786,N_28446,N_27946);
and U29787 (N_29787,N_28360,N_28333);
and U29788 (N_29788,N_27974,N_27697);
nand U29789 (N_29789,N_27891,N_28389);
and U29790 (N_29790,N_28612,N_27845);
nor U29791 (N_29791,N_28521,N_28448);
xor U29792 (N_29792,N_28193,N_28219);
or U29793 (N_29793,N_28545,N_28100);
or U29794 (N_29794,N_28131,N_28141);
nor U29795 (N_29795,N_28731,N_28458);
nor U29796 (N_29796,N_27985,N_27951);
and U29797 (N_29797,N_28708,N_28730);
nor U29798 (N_29798,N_28129,N_28143);
nor U29799 (N_29799,N_28227,N_28225);
xnor U29800 (N_29800,N_28632,N_28659);
nor U29801 (N_29801,N_28075,N_27815);
nand U29802 (N_29802,N_28291,N_27986);
xor U29803 (N_29803,N_27989,N_28017);
or U29804 (N_29804,N_28792,N_28627);
and U29805 (N_29805,N_27913,N_28131);
nor U29806 (N_29806,N_27641,N_27620);
nor U29807 (N_29807,N_28135,N_28282);
nand U29808 (N_29808,N_28469,N_28120);
and U29809 (N_29809,N_28144,N_28752);
nor U29810 (N_29810,N_28760,N_28398);
nor U29811 (N_29811,N_27927,N_27640);
xnor U29812 (N_29812,N_28042,N_28439);
and U29813 (N_29813,N_27679,N_28605);
xor U29814 (N_29814,N_28774,N_28191);
nor U29815 (N_29815,N_27653,N_28145);
xnor U29816 (N_29816,N_28027,N_27885);
nand U29817 (N_29817,N_28653,N_28619);
or U29818 (N_29818,N_28365,N_28502);
or U29819 (N_29819,N_27943,N_28399);
nor U29820 (N_29820,N_27916,N_27653);
nor U29821 (N_29821,N_28101,N_27963);
nor U29822 (N_29822,N_27936,N_28116);
and U29823 (N_29823,N_28218,N_28326);
or U29824 (N_29824,N_28398,N_27603);
or U29825 (N_29825,N_28459,N_28488);
xor U29826 (N_29826,N_28458,N_28176);
nand U29827 (N_29827,N_28220,N_28402);
nor U29828 (N_29828,N_28755,N_28726);
nand U29829 (N_29829,N_28370,N_28475);
nand U29830 (N_29830,N_28014,N_28227);
or U29831 (N_29831,N_28052,N_27906);
or U29832 (N_29832,N_28170,N_27942);
and U29833 (N_29833,N_28061,N_28575);
nand U29834 (N_29834,N_28348,N_28221);
and U29835 (N_29835,N_27789,N_28229);
or U29836 (N_29836,N_28256,N_27952);
xnor U29837 (N_29837,N_27697,N_27806);
or U29838 (N_29838,N_28177,N_28487);
or U29839 (N_29839,N_27996,N_28174);
nand U29840 (N_29840,N_28485,N_27726);
nand U29841 (N_29841,N_28137,N_27684);
nand U29842 (N_29842,N_28086,N_28209);
xor U29843 (N_29843,N_28194,N_27900);
nor U29844 (N_29844,N_27990,N_27877);
or U29845 (N_29845,N_27718,N_28291);
nor U29846 (N_29846,N_27701,N_28642);
and U29847 (N_29847,N_28338,N_28238);
xnor U29848 (N_29848,N_28463,N_28234);
and U29849 (N_29849,N_28401,N_27659);
or U29850 (N_29850,N_28021,N_27889);
nand U29851 (N_29851,N_27600,N_28041);
nor U29852 (N_29852,N_27638,N_28710);
nand U29853 (N_29853,N_27822,N_28214);
and U29854 (N_29854,N_27719,N_27645);
nor U29855 (N_29855,N_28371,N_28303);
nand U29856 (N_29856,N_28676,N_28619);
nand U29857 (N_29857,N_28761,N_28544);
or U29858 (N_29858,N_27908,N_28573);
nand U29859 (N_29859,N_28776,N_27908);
nand U29860 (N_29860,N_28036,N_28226);
and U29861 (N_29861,N_28246,N_28557);
nand U29862 (N_29862,N_28088,N_28412);
nor U29863 (N_29863,N_28360,N_28263);
nand U29864 (N_29864,N_28175,N_28451);
nor U29865 (N_29865,N_27967,N_27897);
and U29866 (N_29866,N_27846,N_28157);
or U29867 (N_29867,N_27823,N_27795);
and U29868 (N_29868,N_28656,N_28677);
nor U29869 (N_29869,N_27796,N_27716);
or U29870 (N_29870,N_28006,N_28138);
xor U29871 (N_29871,N_27650,N_27979);
nor U29872 (N_29872,N_28175,N_28273);
nand U29873 (N_29873,N_27887,N_28319);
nor U29874 (N_29874,N_27775,N_27819);
xor U29875 (N_29875,N_28336,N_27699);
nand U29876 (N_29876,N_27662,N_28785);
or U29877 (N_29877,N_28212,N_28509);
and U29878 (N_29878,N_28501,N_28051);
xnor U29879 (N_29879,N_28020,N_28699);
or U29880 (N_29880,N_27971,N_27898);
nor U29881 (N_29881,N_28094,N_28052);
nor U29882 (N_29882,N_28770,N_28019);
or U29883 (N_29883,N_27843,N_28654);
nor U29884 (N_29884,N_28142,N_28752);
and U29885 (N_29885,N_28598,N_28447);
or U29886 (N_29886,N_28461,N_28542);
xor U29887 (N_29887,N_28724,N_28334);
nor U29888 (N_29888,N_28011,N_27600);
xnor U29889 (N_29889,N_27766,N_28184);
and U29890 (N_29890,N_28042,N_27655);
and U29891 (N_29891,N_28721,N_28092);
and U29892 (N_29892,N_28258,N_27626);
and U29893 (N_29893,N_28708,N_28675);
or U29894 (N_29894,N_28789,N_27975);
nor U29895 (N_29895,N_28274,N_28047);
nor U29896 (N_29896,N_28148,N_28424);
nand U29897 (N_29897,N_27828,N_28079);
nor U29898 (N_29898,N_28278,N_28284);
and U29899 (N_29899,N_28044,N_28141);
xnor U29900 (N_29900,N_28360,N_27774);
nand U29901 (N_29901,N_28717,N_27938);
xor U29902 (N_29902,N_28028,N_27913);
nor U29903 (N_29903,N_28578,N_28224);
nor U29904 (N_29904,N_27611,N_28645);
and U29905 (N_29905,N_27654,N_28273);
nor U29906 (N_29906,N_28293,N_27867);
and U29907 (N_29907,N_27733,N_27928);
and U29908 (N_29908,N_27640,N_28147);
nand U29909 (N_29909,N_28664,N_27944);
nand U29910 (N_29910,N_27959,N_27629);
or U29911 (N_29911,N_28578,N_27906);
or U29912 (N_29912,N_27851,N_27793);
or U29913 (N_29913,N_28404,N_27711);
xor U29914 (N_29914,N_28381,N_27807);
or U29915 (N_29915,N_28129,N_27978);
nand U29916 (N_29916,N_27679,N_27911);
nand U29917 (N_29917,N_28625,N_27805);
xnor U29918 (N_29918,N_28776,N_27702);
nand U29919 (N_29919,N_28488,N_28174);
and U29920 (N_29920,N_28554,N_28510);
nor U29921 (N_29921,N_28738,N_27838);
xnor U29922 (N_29922,N_28495,N_28090);
or U29923 (N_29923,N_28699,N_27940);
xor U29924 (N_29924,N_28301,N_28032);
and U29925 (N_29925,N_28797,N_28310);
nand U29926 (N_29926,N_28015,N_27825);
and U29927 (N_29927,N_28716,N_28691);
nand U29928 (N_29928,N_28147,N_28117);
and U29929 (N_29929,N_28423,N_28675);
nand U29930 (N_29930,N_28591,N_28787);
nor U29931 (N_29931,N_28725,N_28762);
and U29932 (N_29932,N_28365,N_28113);
nor U29933 (N_29933,N_28632,N_28572);
nor U29934 (N_29934,N_28384,N_28202);
or U29935 (N_29935,N_28027,N_28193);
and U29936 (N_29936,N_28661,N_27728);
xnor U29937 (N_29937,N_27670,N_28418);
xor U29938 (N_29938,N_28158,N_27794);
and U29939 (N_29939,N_28578,N_27731);
nand U29940 (N_29940,N_28126,N_27830);
nor U29941 (N_29941,N_28660,N_28239);
nand U29942 (N_29942,N_28493,N_28379);
or U29943 (N_29943,N_28400,N_27747);
xor U29944 (N_29944,N_27770,N_27998);
nand U29945 (N_29945,N_28152,N_28617);
xor U29946 (N_29946,N_28075,N_28634);
or U29947 (N_29947,N_28367,N_27802);
and U29948 (N_29948,N_28722,N_28375);
xnor U29949 (N_29949,N_27896,N_28776);
nand U29950 (N_29950,N_28691,N_28578);
and U29951 (N_29951,N_28100,N_27752);
and U29952 (N_29952,N_28332,N_27771);
xnor U29953 (N_29953,N_27745,N_27663);
or U29954 (N_29954,N_27859,N_27849);
and U29955 (N_29955,N_28263,N_28072);
xnor U29956 (N_29956,N_27691,N_27865);
xnor U29957 (N_29957,N_28556,N_28720);
nor U29958 (N_29958,N_27813,N_28229);
nor U29959 (N_29959,N_27670,N_28620);
or U29960 (N_29960,N_28567,N_28594);
nand U29961 (N_29961,N_28716,N_28582);
nand U29962 (N_29962,N_28302,N_27640);
xor U29963 (N_29963,N_28649,N_27839);
nand U29964 (N_29964,N_27658,N_27790);
and U29965 (N_29965,N_27955,N_27826);
or U29966 (N_29966,N_27603,N_28194);
and U29967 (N_29967,N_27626,N_27905);
nor U29968 (N_29968,N_28056,N_27853);
xnor U29969 (N_29969,N_28481,N_27905);
nor U29970 (N_29970,N_28035,N_27917);
xnor U29971 (N_29971,N_27861,N_28466);
nand U29972 (N_29972,N_28600,N_28390);
nand U29973 (N_29973,N_28526,N_28422);
nor U29974 (N_29974,N_28269,N_27910);
nor U29975 (N_29975,N_28543,N_28387);
or U29976 (N_29976,N_28118,N_28593);
xor U29977 (N_29977,N_28079,N_28683);
and U29978 (N_29978,N_28168,N_28742);
or U29979 (N_29979,N_28478,N_28635);
nor U29980 (N_29980,N_28356,N_27654);
xnor U29981 (N_29981,N_27648,N_28049);
nand U29982 (N_29982,N_28273,N_28299);
nor U29983 (N_29983,N_28281,N_27820);
or U29984 (N_29984,N_28189,N_27906);
nand U29985 (N_29985,N_28327,N_28535);
and U29986 (N_29986,N_27916,N_27771);
xnor U29987 (N_29987,N_28446,N_28531);
or U29988 (N_29988,N_27696,N_27996);
or U29989 (N_29989,N_28783,N_28295);
and U29990 (N_29990,N_28653,N_27864);
and U29991 (N_29991,N_27820,N_28371);
nand U29992 (N_29992,N_27714,N_27762);
or U29993 (N_29993,N_27980,N_28110);
nor U29994 (N_29994,N_28673,N_27908);
xor U29995 (N_29995,N_27871,N_28477);
and U29996 (N_29996,N_28569,N_28009);
and U29997 (N_29997,N_28775,N_28716);
and U29998 (N_29998,N_28101,N_28762);
or U29999 (N_29999,N_27983,N_27766);
nand UO_0 (O_0,N_29525,N_29231);
or UO_1 (O_1,N_29340,N_28892);
xor UO_2 (O_2,N_29094,N_29297);
or UO_3 (O_3,N_29183,N_28979);
xnor UO_4 (O_4,N_29415,N_29011);
or UO_5 (O_5,N_29913,N_29866);
or UO_6 (O_6,N_29926,N_29928);
xnor UO_7 (O_7,N_29603,N_29571);
and UO_8 (O_8,N_28904,N_29002);
or UO_9 (O_9,N_29921,N_29604);
nand UO_10 (O_10,N_29001,N_29541);
or UO_11 (O_11,N_29022,N_29375);
nor UO_12 (O_12,N_29148,N_29523);
and UO_13 (O_13,N_29042,N_28984);
nand UO_14 (O_14,N_29071,N_29981);
nor UO_15 (O_15,N_29566,N_29968);
xor UO_16 (O_16,N_29796,N_29791);
xor UO_17 (O_17,N_29643,N_29450);
or UO_18 (O_18,N_29099,N_29170);
or UO_19 (O_19,N_29295,N_29033);
nand UO_20 (O_20,N_28983,N_29740);
nor UO_21 (O_21,N_29768,N_29987);
or UO_22 (O_22,N_29537,N_29114);
or UO_23 (O_23,N_29472,N_29721);
nor UO_24 (O_24,N_29091,N_28921);
nand UO_25 (O_25,N_28831,N_29140);
or UO_26 (O_26,N_28902,N_28895);
xnor UO_27 (O_27,N_29137,N_29786);
xnor UO_28 (O_28,N_29276,N_29451);
xor UO_29 (O_29,N_29467,N_29560);
or UO_30 (O_30,N_29751,N_28823);
xnor UO_31 (O_31,N_29304,N_28830);
nor UO_32 (O_32,N_29063,N_28941);
xnor UO_33 (O_33,N_29485,N_29238);
xor UO_34 (O_34,N_29186,N_29310);
or UO_35 (O_35,N_29182,N_29120);
and UO_36 (O_36,N_29346,N_28940);
and UO_37 (O_37,N_29809,N_29652);
and UO_38 (O_38,N_29426,N_28874);
nand UO_39 (O_39,N_29126,N_28840);
xor UO_40 (O_40,N_29464,N_29963);
and UO_41 (O_41,N_29247,N_29733);
nor UO_42 (O_42,N_29436,N_29175);
and UO_43 (O_43,N_29106,N_29399);
nor UO_44 (O_44,N_29108,N_29694);
and UO_45 (O_45,N_29365,N_28884);
nand UO_46 (O_46,N_29765,N_28910);
nand UO_47 (O_47,N_29258,N_29457);
or UO_48 (O_48,N_29670,N_29717);
nand UO_49 (O_49,N_29507,N_29452);
or UO_50 (O_50,N_29995,N_28943);
or UO_51 (O_51,N_29152,N_29318);
xnor UO_52 (O_52,N_29852,N_29727);
and UO_53 (O_53,N_28924,N_28836);
xnor UO_54 (O_54,N_29379,N_29089);
or UO_55 (O_55,N_28825,N_29028);
or UO_56 (O_56,N_29916,N_28938);
or UO_57 (O_57,N_28880,N_29435);
nand UO_58 (O_58,N_29096,N_28956);
or UO_59 (O_59,N_29520,N_29087);
nand UO_60 (O_60,N_29356,N_29532);
xor UO_61 (O_61,N_29893,N_29813);
xor UO_62 (O_62,N_29868,N_29688);
xor UO_63 (O_63,N_29699,N_29815);
and UO_64 (O_64,N_29376,N_29848);
xor UO_65 (O_65,N_29955,N_28817);
nor UO_66 (O_66,N_29103,N_29121);
nand UO_67 (O_67,N_29335,N_28872);
nor UO_68 (O_68,N_29040,N_29147);
nor UO_69 (O_69,N_29644,N_29219);
or UO_70 (O_70,N_29403,N_29506);
nand UO_71 (O_71,N_28826,N_28862);
and UO_72 (O_72,N_29931,N_28809);
nand UO_73 (O_73,N_29320,N_29620);
or UO_74 (O_74,N_29650,N_29187);
or UO_75 (O_75,N_29930,N_29691);
or UO_76 (O_76,N_29059,N_29783);
nor UO_77 (O_77,N_28970,N_29927);
nand UO_78 (O_78,N_28821,N_28978);
nand UO_79 (O_79,N_29263,N_28975);
and UO_80 (O_80,N_29818,N_29802);
nand UO_81 (O_81,N_29156,N_29385);
or UO_82 (O_82,N_29900,N_29766);
nor UO_83 (O_83,N_29296,N_29902);
nand UO_84 (O_84,N_29171,N_29594);
or UO_85 (O_85,N_29195,N_29224);
nor UO_86 (O_86,N_28959,N_29221);
xnor UO_87 (O_87,N_29865,N_29366);
nand UO_88 (O_88,N_28863,N_29706);
nand UO_89 (O_89,N_29045,N_29445);
nor UO_90 (O_90,N_29642,N_29159);
nor UO_91 (O_91,N_29012,N_29715);
and UO_92 (O_92,N_29653,N_28873);
nor UO_93 (O_93,N_29135,N_29861);
nand UO_94 (O_94,N_29651,N_29648);
and UO_95 (O_95,N_29085,N_29299);
nand UO_96 (O_96,N_29458,N_29855);
xnor UO_97 (O_97,N_28912,N_29634);
nand UO_98 (O_98,N_29947,N_29943);
xor UO_99 (O_99,N_29784,N_29845);
and UO_100 (O_100,N_29790,N_29701);
nand UO_101 (O_101,N_28991,N_29716);
nand UO_102 (O_102,N_29118,N_29991);
nor UO_103 (O_103,N_29847,N_29627);
and UO_104 (O_104,N_29919,N_29162);
nand UO_105 (O_105,N_29803,N_29607);
nor UO_106 (O_106,N_29361,N_29075);
nand UO_107 (O_107,N_29777,N_28837);
nand UO_108 (O_108,N_29495,N_29392);
nand UO_109 (O_109,N_29592,N_29516);
nand UO_110 (O_110,N_29542,N_29758);
and UO_111 (O_111,N_29239,N_29637);
xnor UO_112 (O_112,N_29241,N_29111);
nor UO_113 (O_113,N_29128,N_29117);
xnor UO_114 (O_114,N_29227,N_29885);
xor UO_115 (O_115,N_29508,N_29044);
and UO_116 (O_116,N_29273,N_29317);
nor UO_117 (O_117,N_29110,N_29976);
nand UO_118 (O_118,N_29799,N_29709);
nand UO_119 (O_119,N_29115,N_29867);
nor UO_120 (O_120,N_29671,N_28866);
nor UO_121 (O_121,N_29797,N_29951);
or UO_122 (O_122,N_29029,N_29685);
xnor UO_123 (O_123,N_29368,N_28923);
nor UO_124 (O_124,N_29084,N_29223);
or UO_125 (O_125,N_29271,N_28888);
nand UO_126 (O_126,N_29354,N_29226);
nand UO_127 (O_127,N_29357,N_29262);
xnor UO_128 (O_128,N_29817,N_29025);
nor UO_129 (O_129,N_29536,N_29582);
nand UO_130 (O_130,N_29477,N_29208);
nor UO_131 (O_131,N_29819,N_29104);
nand UO_132 (O_132,N_28833,N_29077);
xor UO_133 (O_133,N_29251,N_29401);
and UO_134 (O_134,N_29617,N_29568);
nand UO_135 (O_135,N_28914,N_29490);
nand UO_136 (O_136,N_29672,N_28887);
and UO_137 (O_137,N_28942,N_29336);
xor UO_138 (O_138,N_28977,N_29267);
nor UO_139 (O_139,N_29422,N_29377);
nor UO_140 (O_140,N_29447,N_28841);
and UO_141 (O_141,N_29906,N_29132);
or UO_142 (O_142,N_29362,N_29441);
or UO_143 (O_143,N_29048,N_29315);
and UO_144 (O_144,N_29475,N_29614);
nor UO_145 (O_145,N_29101,N_28818);
xor UO_146 (O_146,N_29693,N_29524);
xnor UO_147 (O_147,N_29641,N_29222);
xor UO_148 (O_148,N_29489,N_29351);
nand UO_149 (O_149,N_29405,N_29983);
xnor UO_150 (O_150,N_29034,N_29851);
and UO_151 (O_151,N_29204,N_28882);
or UO_152 (O_152,N_28964,N_28930);
xor UO_153 (O_153,N_29288,N_29246);
or UO_154 (O_154,N_29439,N_29367);
nand UO_155 (O_155,N_29774,N_29997);
or UO_156 (O_156,N_29655,N_29546);
and UO_157 (O_157,N_29825,N_29255);
or UO_158 (O_158,N_29697,N_29453);
or UO_159 (O_159,N_29824,N_29984);
xor UO_160 (O_160,N_29944,N_29862);
xnor UO_161 (O_161,N_29918,N_29789);
nor UO_162 (O_162,N_28919,N_29437);
nand UO_163 (O_163,N_29373,N_29563);
nor UO_164 (O_164,N_29260,N_29965);
and UO_165 (O_165,N_29561,N_29167);
and UO_166 (O_166,N_29726,N_29556);
nand UO_167 (O_167,N_29008,N_29319);
nor UO_168 (O_168,N_29282,N_28849);
and UO_169 (O_169,N_29083,N_29946);
and UO_170 (O_170,N_29213,N_28990);
xnor UO_171 (O_171,N_29780,N_29687);
nand UO_172 (O_172,N_28992,N_29901);
xor UO_173 (O_173,N_28987,N_29193);
xor UO_174 (O_174,N_29431,N_29513);
xnor UO_175 (O_175,N_28898,N_28929);
xor UO_176 (O_176,N_29631,N_29748);
nand UO_177 (O_177,N_29678,N_29611);
nand UO_178 (O_178,N_29492,N_29434);
or UO_179 (O_179,N_29081,N_29338);
nor UO_180 (O_180,N_29989,N_29657);
or UO_181 (O_181,N_29142,N_29707);
and UO_182 (O_182,N_29076,N_28814);
nand UO_183 (O_183,N_29181,N_29498);
nand UO_184 (O_184,N_29584,N_29949);
nand UO_185 (O_185,N_29762,N_29739);
nand UO_186 (O_186,N_29662,N_29849);
and UO_187 (O_187,N_29805,N_29579);
and UO_188 (O_188,N_29858,N_28935);
nand UO_189 (O_189,N_29889,N_29158);
xor UO_190 (O_190,N_28850,N_29214);
and UO_191 (O_191,N_29149,N_29487);
and UO_192 (O_192,N_28973,N_29062);
nor UO_193 (O_193,N_29754,N_29736);
xor UO_194 (O_194,N_28877,N_29290);
xor UO_195 (O_195,N_29912,N_28847);
xor UO_196 (O_196,N_29937,N_29681);
xnor UO_197 (O_197,N_29842,N_28952);
xnor UO_198 (O_198,N_29755,N_29261);
nor UO_199 (O_199,N_29808,N_29278);
nand UO_200 (O_200,N_29138,N_29703);
nand UO_201 (O_201,N_29713,N_29032);
and UO_202 (O_202,N_29667,N_29551);
or UO_203 (O_203,N_29811,N_29558);
or UO_204 (O_204,N_29610,N_29359);
nor UO_205 (O_205,N_28846,N_29207);
nand UO_206 (O_206,N_29067,N_29632);
or UO_207 (O_207,N_29831,N_28805);
nor UO_208 (O_208,N_29112,N_29006);
nor UO_209 (O_209,N_29689,N_29712);
or UO_210 (O_210,N_29035,N_28865);
or UO_211 (O_211,N_28807,N_29229);
nand UO_212 (O_212,N_29312,N_29872);
or UO_213 (O_213,N_29870,N_28999);
nand UO_214 (O_214,N_29234,N_29342);
or UO_215 (O_215,N_28864,N_29522);
xnor UO_216 (O_216,N_29027,N_28918);
or UO_217 (O_217,N_29601,N_28813);
xnor UO_218 (O_218,N_29932,N_29800);
nand UO_219 (O_219,N_29917,N_29185);
nand UO_220 (O_220,N_28913,N_29455);
or UO_221 (O_221,N_29599,N_29857);
and UO_222 (O_222,N_29844,N_28804);
xor UO_223 (O_223,N_29188,N_29178);
xnor UO_224 (O_224,N_29125,N_28982);
and UO_225 (O_225,N_29444,N_29009);
and UO_226 (O_226,N_28867,N_28876);
nand UO_227 (O_227,N_29016,N_29358);
nand UO_228 (O_228,N_29539,N_29624);
or UO_229 (O_229,N_29230,N_29243);
and UO_230 (O_230,N_29734,N_29216);
or UO_231 (O_231,N_29378,N_28907);
nor UO_232 (O_232,N_29722,N_28934);
nor UO_233 (O_233,N_29547,N_29846);
or UO_234 (O_234,N_29041,N_29690);
and UO_235 (O_235,N_29512,N_29854);
and UO_236 (O_236,N_29549,N_28875);
nand UO_237 (O_237,N_29890,N_29036);
xnor UO_238 (O_238,N_29019,N_29211);
or UO_239 (O_239,N_29286,N_29904);
xor UO_240 (O_240,N_29910,N_29837);
and UO_241 (O_241,N_29202,N_29285);
and UO_242 (O_242,N_29978,N_29788);
nor UO_243 (O_243,N_28967,N_29920);
and UO_244 (O_244,N_29324,N_29350);
or UO_245 (O_245,N_29771,N_29575);
xor UO_246 (O_246,N_29371,N_29822);
xor UO_247 (O_247,N_29272,N_29533);
nand UO_248 (O_248,N_28899,N_29414);
and UO_249 (O_249,N_29051,N_29596);
xor UO_250 (O_250,N_29958,N_29554);
and UO_251 (O_251,N_29275,N_29669);
or UO_252 (O_252,N_29654,N_29518);
xor UO_253 (O_253,N_29664,N_29370);
nor UO_254 (O_254,N_29388,N_29322);
nor UO_255 (O_255,N_29107,N_29668);
or UO_256 (O_256,N_29122,N_29155);
nand UO_257 (O_257,N_29218,N_29418);
or UO_258 (O_258,N_29374,N_28911);
xnor UO_259 (O_259,N_29645,N_29412);
or UO_260 (O_260,N_29612,N_29759);
and UO_261 (O_261,N_29079,N_29382);
nor UO_262 (O_262,N_29684,N_29938);
nor UO_263 (O_263,N_29109,N_29443);
nand UO_264 (O_264,N_29280,N_29303);
nor UO_265 (O_265,N_29469,N_29823);
or UO_266 (O_266,N_29479,N_29725);
and UO_267 (O_267,N_29665,N_28926);
nor UO_268 (O_268,N_29924,N_29225);
nand UO_269 (O_269,N_29764,N_28852);
xor UO_270 (O_270,N_29562,N_29004);
nor UO_271 (O_271,N_29602,N_28858);
nor UO_272 (O_272,N_29745,N_29360);
nand UO_273 (O_273,N_29066,N_29173);
nor UO_274 (O_274,N_28961,N_28922);
xor UO_275 (O_275,N_29491,N_29807);
nand UO_276 (O_276,N_29269,N_28933);
and UO_277 (O_277,N_29836,N_29994);
or UO_278 (O_278,N_29124,N_28932);
or UO_279 (O_279,N_29074,N_28960);
and UO_280 (O_280,N_29567,N_28829);
nor UO_281 (O_281,N_29500,N_28915);
and UO_282 (O_282,N_29199,N_28845);
nand UO_283 (O_283,N_29274,N_29738);
nor UO_284 (O_284,N_29907,N_29220);
and UO_285 (O_285,N_29527,N_29871);
nor UO_286 (O_286,N_29249,N_29496);
and UO_287 (O_287,N_29037,N_29018);
nand UO_288 (O_288,N_29086,N_29293);
and UO_289 (O_289,N_29640,N_28844);
or UO_290 (O_290,N_29502,N_29702);
and UO_291 (O_291,N_29100,N_29682);
nor UO_292 (O_292,N_29886,N_29078);
and UO_293 (O_293,N_29198,N_29157);
and UO_294 (O_294,N_29517,N_28883);
xnor UO_295 (O_295,N_29194,N_29795);
nand UO_296 (O_296,N_28801,N_29153);
nand UO_297 (O_297,N_29894,N_29898);
and UO_298 (O_298,N_29308,N_29459);
nor UO_299 (O_299,N_29565,N_29511);
xnor UO_300 (O_300,N_29573,N_28897);
xnor UO_301 (O_301,N_29971,N_29323);
xor UO_302 (O_302,N_29020,N_29497);
or UO_303 (O_303,N_29929,N_29268);
nand UO_304 (O_304,N_29164,N_29804);
xor UO_305 (O_305,N_28945,N_29301);
nand UO_306 (O_306,N_29600,N_29184);
or UO_307 (O_307,N_29394,N_29052);
nor UO_308 (O_308,N_28878,N_28954);
or UO_309 (O_309,N_29339,N_29948);
nor UO_310 (O_310,N_28997,N_29154);
xnor UO_311 (O_311,N_28966,N_29840);
xnor UO_312 (O_312,N_29772,N_29030);
or UO_313 (O_313,N_29460,N_29179);
xor UO_314 (O_314,N_29364,N_29410);
xnor UO_315 (O_315,N_29625,N_29345);
nand UO_316 (O_316,N_29630,N_29742);
xor UO_317 (O_317,N_29781,N_29191);
and UO_318 (O_318,N_29950,N_29408);
or UO_319 (O_319,N_29209,N_29972);
and UO_320 (O_320,N_29105,N_29675);
or UO_321 (O_321,N_28976,N_29623);
and UO_322 (O_322,N_29065,N_29986);
nand UO_323 (O_323,N_29925,N_29139);
nor UO_324 (O_324,N_29869,N_28860);
xnor UO_325 (O_325,N_29881,N_28803);
or UO_326 (O_326,N_29704,N_29746);
or UO_327 (O_327,N_29663,N_28812);
nand UO_328 (O_328,N_29245,N_29821);
and UO_329 (O_329,N_28900,N_29834);
or UO_330 (O_330,N_29420,N_29387);
or UO_331 (O_331,N_28920,N_29070);
and UO_332 (O_332,N_29311,N_29935);
xor UO_333 (O_333,N_29429,N_29550);
and UO_334 (O_334,N_29283,N_29969);
nor UO_335 (O_335,N_29060,N_28859);
xor UO_336 (O_336,N_29123,N_29966);
and UO_337 (O_337,N_29521,N_29705);
nand UO_338 (O_338,N_29143,N_29695);
xor UO_339 (O_339,N_29528,N_29021);
xor UO_340 (O_340,N_29874,N_29386);
nand UO_341 (O_341,N_28903,N_29134);
or UO_342 (O_342,N_29448,N_29967);
or UO_343 (O_343,N_29905,N_29656);
and UO_344 (O_344,N_29692,N_29775);
or UO_345 (O_345,N_29337,N_29720);
xor UO_346 (O_346,N_29875,N_29960);
nand UO_347 (O_347,N_29794,N_28917);
nor UO_348 (O_348,N_29015,N_29332);
and UO_349 (O_349,N_29144,N_29259);
nor UO_350 (O_350,N_29760,N_28916);
nor UO_351 (O_351,N_29635,N_28824);
and UO_352 (O_352,N_29622,N_29856);
or UO_353 (O_353,N_29348,N_29880);
nor UO_354 (O_354,N_29330,N_28981);
nand UO_355 (O_355,N_29253,N_29146);
or UO_356 (O_356,N_29406,N_29119);
and UO_357 (O_357,N_29676,N_29432);
nor UO_358 (O_358,N_29731,N_29572);
or UO_359 (O_359,N_29718,N_28905);
or UO_360 (O_360,N_28962,N_29787);
or UO_361 (O_361,N_29163,N_29628);
and UO_362 (O_362,N_29977,N_29024);
xnor UO_363 (O_363,N_29493,N_29534);
or UO_364 (O_364,N_29266,N_29683);
and UO_365 (O_365,N_29499,N_29992);
xnor UO_366 (O_366,N_29633,N_29730);
or UO_367 (O_367,N_29996,N_29569);
and UO_368 (O_368,N_29933,N_29402);
xor UO_369 (O_369,N_28946,N_29934);
nor UO_370 (O_370,N_28816,N_28851);
nor UO_371 (O_371,N_29480,N_29769);
xnor UO_372 (O_372,N_29820,N_29659);
and UO_373 (O_373,N_29284,N_29409);
nand UO_374 (O_374,N_28810,N_29999);
xnor UO_375 (O_375,N_29309,N_29250);
nor UO_376 (O_376,N_29017,N_29333);
nand UO_377 (O_377,N_29093,N_29470);
and UO_378 (O_378,N_29054,N_29626);
nand UO_379 (O_379,N_29723,N_29169);
and UO_380 (O_380,N_28819,N_28994);
xor UO_381 (O_381,N_29363,N_29419);
xor UO_382 (O_382,N_29454,N_28868);
and UO_383 (O_383,N_28906,N_29352);
nand UO_384 (O_384,N_29168,N_29215);
nand UO_385 (O_385,N_29150,N_29236);
xor UO_386 (O_386,N_29779,N_28842);
xnor UO_387 (O_387,N_29982,N_28835);
and UO_388 (O_388,N_28890,N_29830);
nand UO_389 (O_389,N_29585,N_29553);
and UO_390 (O_390,N_29843,N_29133);
nand UO_391 (O_391,N_29555,N_29744);
and UO_392 (O_392,N_29589,N_29233);
and UO_393 (O_393,N_28998,N_29763);
or UO_394 (O_394,N_29488,N_29090);
nor UO_395 (O_395,N_29072,N_29192);
nand UO_396 (O_396,N_29430,N_29714);
or UO_397 (O_397,N_29400,N_29292);
or UO_398 (O_398,N_29073,N_29265);
and UO_399 (O_399,N_29793,N_29031);
and UO_400 (O_400,N_29782,N_29026);
and UO_401 (O_401,N_29302,N_29095);
nor UO_402 (O_402,N_28953,N_29879);
and UO_403 (O_403,N_28908,N_29264);
nor UO_404 (O_404,N_29092,N_29621);
or UO_405 (O_405,N_29911,N_29334);
xor UO_406 (O_406,N_29428,N_29177);
xnor UO_407 (O_407,N_29055,N_29883);
xor UO_408 (O_408,N_29395,N_29313);
or UO_409 (O_409,N_29859,N_29270);
and UO_410 (O_410,N_29411,N_29636);
nand UO_411 (O_411,N_29914,N_29891);
or UO_412 (O_412,N_29985,N_29129);
or UO_413 (O_413,N_29413,N_28834);
nand UO_414 (O_414,N_29679,N_29038);
or UO_415 (O_415,N_28848,N_29344);
nor UO_416 (O_416,N_29398,N_28832);
xor UO_417 (O_417,N_29484,N_28891);
nor UO_418 (O_418,N_28869,N_29940);
nor UO_419 (O_419,N_29959,N_29732);
nor UO_420 (O_420,N_29529,N_29729);
or UO_421 (O_421,N_29853,N_28963);
or UO_422 (O_422,N_29466,N_29993);
or UO_423 (O_423,N_29331,N_29098);
nor UO_424 (O_424,N_29835,N_29962);
and UO_425 (O_425,N_29980,N_29446);
nand UO_426 (O_426,N_28937,N_29442);
and UO_427 (O_427,N_28993,N_28986);
nor UO_428 (O_428,N_28822,N_29242);
nor UO_429 (O_429,N_28969,N_29014);
and UO_430 (O_430,N_29580,N_29393);
and UO_431 (O_431,N_29544,N_29023);
or UO_432 (O_432,N_29974,N_29277);
nor UO_433 (O_433,N_28901,N_29828);
and UO_434 (O_434,N_28957,N_28985);
or UO_435 (O_435,N_29494,N_29510);
nand UO_436 (O_436,N_29396,N_28988);
xnor UO_437 (O_437,N_28854,N_28861);
nor UO_438 (O_438,N_29583,N_29449);
xor UO_439 (O_439,N_29903,N_29145);
nand UO_440 (O_440,N_28995,N_29899);
or UO_441 (O_441,N_29289,N_29240);
nand UO_442 (O_442,N_29761,N_29770);
xnor UO_443 (O_443,N_29741,N_29792);
nor UO_444 (O_444,N_29468,N_29053);
and UO_445 (O_445,N_29456,N_29203);
and UO_446 (O_446,N_28955,N_29535);
xnor UO_447 (O_447,N_29248,N_29039);
and UO_448 (O_448,N_29570,N_28968);
or UO_449 (O_449,N_29973,N_29578);
and UO_450 (O_450,N_29839,N_28808);
and UO_451 (O_451,N_29189,N_29609);
nand UO_452 (O_452,N_29281,N_29353);
xnor UO_453 (O_453,N_29082,N_28815);
or UO_454 (O_454,N_29674,N_29314);
xor UO_455 (O_455,N_29166,N_29708);
xor UO_456 (O_456,N_29404,N_29176);
and UO_457 (O_457,N_29327,N_29505);
and UO_458 (O_458,N_29827,N_29235);
nand UO_459 (O_459,N_29936,N_29658);
xnor UO_460 (O_460,N_29922,N_29049);
nor UO_461 (O_461,N_29069,N_29471);
xnor UO_462 (O_462,N_28948,N_29257);
nor UO_463 (O_463,N_29425,N_29397);
nor UO_464 (O_464,N_29212,N_29228);
or UO_465 (O_465,N_29616,N_29478);
xnor UO_466 (O_466,N_29097,N_28802);
xnor UO_467 (O_467,N_29957,N_29975);
xnor UO_468 (O_468,N_29673,N_29329);
xor UO_469 (O_469,N_29884,N_29618);
and UO_470 (O_470,N_29649,N_29606);
or UO_471 (O_471,N_28838,N_28811);
nand UO_472 (O_472,N_28843,N_28965);
nor UO_473 (O_473,N_29232,N_29990);
nand UO_474 (O_474,N_29619,N_29538);
nor UO_475 (O_475,N_29050,N_29961);
xnor UO_476 (O_476,N_29666,N_29829);
and UO_477 (O_477,N_29509,N_29998);
and UO_478 (O_478,N_29588,N_29279);
nor UO_479 (O_479,N_29530,N_29954);
xnor UO_480 (O_480,N_28853,N_29325);
xor UO_481 (O_481,N_29476,N_29964);
and UO_482 (O_482,N_29576,N_28896);
nor UO_483 (O_483,N_29131,N_29941);
and UO_484 (O_484,N_29841,N_29013);
nor UO_485 (O_485,N_29463,N_28856);
nor UO_486 (O_486,N_28839,N_29728);
nor UO_487 (O_487,N_29557,N_28980);
nand UO_488 (O_488,N_29380,N_29390);
xor UO_489 (O_489,N_29328,N_29056);
nor UO_490 (O_490,N_28927,N_29814);
nand UO_491 (O_491,N_29613,N_29136);
or UO_492 (O_492,N_29481,N_29165);
xnor UO_493 (O_493,N_29160,N_29088);
xor UO_494 (O_494,N_29172,N_29200);
and UO_495 (O_495,N_29660,N_29307);
xnor UO_496 (O_496,N_28871,N_28951);
or UO_497 (O_497,N_28996,N_29306);
or UO_498 (O_498,N_29838,N_29423);
nand UO_499 (O_499,N_29895,N_29559);
nor UO_500 (O_500,N_28909,N_28936);
or UO_501 (O_501,N_29347,N_29298);
or UO_502 (O_502,N_29064,N_29503);
nand UO_503 (O_503,N_29876,N_29174);
nor UO_504 (O_504,N_29190,N_29294);
nor UO_505 (O_505,N_28828,N_29942);
or UO_506 (O_506,N_29773,N_28870);
nor UO_507 (O_507,N_29438,N_29776);
nor UO_508 (O_508,N_29326,N_29724);
nand UO_509 (O_509,N_29465,N_29696);
nor UO_510 (O_510,N_29979,N_29711);
nor UO_511 (O_511,N_29750,N_29638);
and UO_512 (O_512,N_29564,N_29427);
or UO_513 (O_513,N_29287,N_29381);
nor UO_514 (O_514,N_29877,N_29545);
nand UO_515 (O_515,N_29826,N_29970);
nor UO_516 (O_516,N_29526,N_28879);
nand UO_517 (O_517,N_28800,N_29908);
nand UO_518 (O_518,N_29369,N_29882);
nand UO_519 (O_519,N_29595,N_29068);
xnor UO_520 (O_520,N_29543,N_29909);
xor UO_521 (O_521,N_29756,N_29719);
and UO_522 (O_522,N_28972,N_29433);
or UO_523 (O_523,N_29349,N_29749);
or UO_524 (O_524,N_29300,N_29531);
nor UO_525 (O_525,N_29141,N_29615);
xnor UO_526 (O_526,N_28971,N_29341);
nor UO_527 (O_527,N_29515,N_29680);
and UO_528 (O_528,N_29586,N_29597);
nor UO_529 (O_529,N_29254,N_29737);
nor UO_530 (O_530,N_29629,N_29196);
xor UO_531 (O_531,N_28893,N_29832);
xor UO_532 (O_532,N_28806,N_29519);
xor UO_533 (O_533,N_29355,N_29753);
xnor UO_534 (O_534,N_29806,N_29873);
xor UO_535 (O_535,N_28886,N_29608);
xor UO_536 (O_536,N_29474,N_29047);
nor UO_537 (O_537,N_29237,N_29197);
nand UO_538 (O_538,N_29514,N_29252);
or UO_539 (O_539,N_29540,N_29587);
nand UO_540 (O_540,N_29593,N_29113);
and UO_541 (O_541,N_29007,N_28950);
xnor UO_542 (O_542,N_29391,N_28855);
xnor UO_543 (O_543,N_28931,N_29833);
nand UO_544 (O_544,N_29161,N_29953);
xor UO_545 (O_545,N_29057,N_29205);
xnor UO_546 (O_546,N_29757,N_29860);
and UO_547 (O_547,N_29180,N_29710);
nand UO_548 (O_548,N_29752,N_29591);
xnor UO_549 (O_549,N_29735,N_29210);
and UO_550 (O_550,N_29343,N_29574);
nor UO_551 (O_551,N_29863,N_29256);
and UO_552 (O_552,N_29878,N_29798);
nand UO_553 (O_553,N_29372,N_28894);
nor UO_554 (O_554,N_28944,N_29058);
xor UO_555 (O_555,N_29217,N_29416);
nand UO_556 (O_556,N_29473,N_29700);
or UO_557 (O_557,N_29639,N_28939);
nand UO_558 (O_558,N_29801,N_29850);
nand UO_559 (O_559,N_29389,N_29005);
nand UO_560 (O_560,N_29061,N_29812);
xor UO_561 (O_561,N_29778,N_29440);
xor UO_562 (O_562,N_28827,N_29151);
xnor UO_563 (O_563,N_29043,N_29000);
nor UO_564 (O_564,N_28958,N_29605);
and UO_565 (O_565,N_29810,N_29010);
xnor UO_566 (O_566,N_29482,N_29767);
and UO_567 (O_567,N_29206,N_29407);
or UO_568 (O_568,N_29646,N_29698);
or UO_569 (O_569,N_29417,N_29945);
or UO_570 (O_570,N_29501,N_29483);
xnor UO_571 (O_571,N_29552,N_28949);
nand UO_572 (O_572,N_29102,N_29577);
nand UO_573 (O_573,N_29424,N_29915);
nand UO_574 (O_574,N_28889,N_29080);
nor UO_575 (O_575,N_29598,N_29923);
or UO_576 (O_576,N_29677,N_29462);
or UO_577 (O_577,N_29291,N_29661);
xor UO_578 (O_578,N_28928,N_29316);
and UO_579 (O_579,N_29816,N_29504);
and UO_580 (O_580,N_29686,N_29201);
nor UO_581 (O_581,N_29305,N_29003);
and UO_582 (O_582,N_28857,N_29747);
nor UO_583 (O_583,N_29321,N_29383);
nand UO_584 (O_584,N_29581,N_28974);
xor UO_585 (O_585,N_29956,N_29939);
xor UO_586 (O_586,N_29116,N_29988);
xor UO_587 (O_587,N_29590,N_28820);
nand UO_588 (O_588,N_28885,N_29548);
or UO_589 (O_589,N_29952,N_29888);
nor UO_590 (O_590,N_29743,N_28989);
xnor UO_591 (O_591,N_29130,N_29244);
nor UO_592 (O_592,N_29486,N_29461);
and UO_593 (O_593,N_28947,N_29647);
or UO_594 (O_594,N_29046,N_29892);
and UO_595 (O_595,N_29887,N_29127);
xnor UO_596 (O_596,N_28925,N_29785);
nor UO_597 (O_597,N_29897,N_29384);
nand UO_598 (O_598,N_29864,N_29896);
or UO_599 (O_599,N_29421,N_28881);
xnor UO_600 (O_600,N_29694,N_29313);
xor UO_601 (O_601,N_29024,N_28832);
nor UO_602 (O_602,N_29011,N_29970);
nor UO_603 (O_603,N_29419,N_29869);
xor UO_604 (O_604,N_29213,N_29464);
xor UO_605 (O_605,N_29176,N_28955);
or UO_606 (O_606,N_29555,N_29004);
or UO_607 (O_607,N_29462,N_29943);
or UO_608 (O_608,N_29895,N_29814);
xor UO_609 (O_609,N_28850,N_29001);
nand UO_610 (O_610,N_28991,N_29916);
or UO_611 (O_611,N_29971,N_29192);
and UO_612 (O_612,N_28800,N_29305);
or UO_613 (O_613,N_29934,N_29586);
and UO_614 (O_614,N_29517,N_29780);
xor UO_615 (O_615,N_28888,N_28905);
nand UO_616 (O_616,N_28856,N_29071);
xnor UO_617 (O_617,N_29402,N_29072);
nor UO_618 (O_618,N_29680,N_29930);
and UO_619 (O_619,N_29470,N_29412);
nor UO_620 (O_620,N_29583,N_29977);
nor UO_621 (O_621,N_29826,N_29827);
or UO_622 (O_622,N_29750,N_29924);
and UO_623 (O_623,N_29188,N_29291);
nor UO_624 (O_624,N_29982,N_29808);
or UO_625 (O_625,N_29165,N_29762);
xnor UO_626 (O_626,N_29050,N_29344);
nor UO_627 (O_627,N_29753,N_28896);
and UO_628 (O_628,N_29285,N_29400);
nor UO_629 (O_629,N_28893,N_29499);
and UO_630 (O_630,N_29174,N_28832);
and UO_631 (O_631,N_29073,N_29218);
nand UO_632 (O_632,N_29898,N_29643);
nor UO_633 (O_633,N_28977,N_28831);
nand UO_634 (O_634,N_29356,N_29963);
nor UO_635 (O_635,N_29585,N_29333);
xnor UO_636 (O_636,N_29067,N_29494);
xor UO_637 (O_637,N_29767,N_29643);
xnor UO_638 (O_638,N_29451,N_29886);
nand UO_639 (O_639,N_29825,N_29310);
nor UO_640 (O_640,N_28861,N_29752);
nand UO_641 (O_641,N_29557,N_29214);
or UO_642 (O_642,N_29934,N_29184);
and UO_643 (O_643,N_29133,N_29328);
nand UO_644 (O_644,N_29525,N_29386);
xnor UO_645 (O_645,N_29368,N_29940);
or UO_646 (O_646,N_29681,N_29911);
nand UO_647 (O_647,N_29042,N_28965);
and UO_648 (O_648,N_29878,N_29907);
or UO_649 (O_649,N_29219,N_29274);
or UO_650 (O_650,N_29217,N_29066);
nor UO_651 (O_651,N_29015,N_28914);
nand UO_652 (O_652,N_29290,N_29926);
nand UO_653 (O_653,N_29081,N_28905);
xnor UO_654 (O_654,N_29842,N_29602);
xor UO_655 (O_655,N_29698,N_29469);
xnor UO_656 (O_656,N_29855,N_29649);
nor UO_657 (O_657,N_29893,N_29517);
or UO_658 (O_658,N_29445,N_28890);
or UO_659 (O_659,N_29969,N_29938);
nand UO_660 (O_660,N_29007,N_28841);
or UO_661 (O_661,N_29974,N_29348);
nor UO_662 (O_662,N_28917,N_29901);
nand UO_663 (O_663,N_29466,N_29791);
nor UO_664 (O_664,N_29394,N_29346);
nor UO_665 (O_665,N_29374,N_29338);
and UO_666 (O_666,N_29513,N_29153);
nor UO_667 (O_667,N_29726,N_28978);
nand UO_668 (O_668,N_29268,N_29805);
nor UO_669 (O_669,N_29406,N_28868);
and UO_670 (O_670,N_29701,N_29349);
xor UO_671 (O_671,N_29236,N_29584);
and UO_672 (O_672,N_29362,N_29523);
and UO_673 (O_673,N_29566,N_29948);
and UO_674 (O_674,N_29834,N_29199);
nor UO_675 (O_675,N_28976,N_29776);
and UO_676 (O_676,N_28960,N_29271);
nand UO_677 (O_677,N_29454,N_29880);
xor UO_678 (O_678,N_29359,N_29059);
and UO_679 (O_679,N_29972,N_28861);
xor UO_680 (O_680,N_29357,N_29162);
nand UO_681 (O_681,N_28891,N_29256);
nor UO_682 (O_682,N_29772,N_29555);
or UO_683 (O_683,N_29687,N_29452);
or UO_684 (O_684,N_29016,N_29558);
nor UO_685 (O_685,N_28854,N_29151);
and UO_686 (O_686,N_29326,N_29458);
xor UO_687 (O_687,N_29311,N_29224);
nand UO_688 (O_688,N_29733,N_29105);
and UO_689 (O_689,N_29727,N_29731);
nor UO_690 (O_690,N_29429,N_29491);
and UO_691 (O_691,N_29172,N_29919);
and UO_692 (O_692,N_29143,N_28807);
xor UO_693 (O_693,N_29423,N_29196);
and UO_694 (O_694,N_29369,N_29136);
xor UO_695 (O_695,N_29522,N_29461);
nor UO_696 (O_696,N_29700,N_29662);
nor UO_697 (O_697,N_29261,N_29109);
or UO_698 (O_698,N_29524,N_29253);
or UO_699 (O_699,N_29186,N_29526);
or UO_700 (O_700,N_29712,N_29042);
xnor UO_701 (O_701,N_29596,N_29139);
nor UO_702 (O_702,N_29147,N_29455);
and UO_703 (O_703,N_29495,N_29699);
nand UO_704 (O_704,N_29900,N_29280);
and UO_705 (O_705,N_29449,N_28998);
nand UO_706 (O_706,N_29016,N_28879);
and UO_707 (O_707,N_29964,N_29294);
nand UO_708 (O_708,N_29591,N_29985);
nand UO_709 (O_709,N_29731,N_29379);
xor UO_710 (O_710,N_29253,N_29641);
or UO_711 (O_711,N_29064,N_29420);
nor UO_712 (O_712,N_28819,N_28888);
and UO_713 (O_713,N_29269,N_29523);
nand UO_714 (O_714,N_29685,N_28989);
or UO_715 (O_715,N_29167,N_29313);
xor UO_716 (O_716,N_29715,N_29539);
nor UO_717 (O_717,N_29915,N_29333);
nor UO_718 (O_718,N_28935,N_29555);
nor UO_719 (O_719,N_29427,N_29251);
and UO_720 (O_720,N_28870,N_28900);
nor UO_721 (O_721,N_29117,N_28810);
nand UO_722 (O_722,N_29942,N_29560);
nor UO_723 (O_723,N_29475,N_28996);
nor UO_724 (O_724,N_28895,N_29068);
nor UO_725 (O_725,N_29226,N_28847);
or UO_726 (O_726,N_29998,N_29348);
and UO_727 (O_727,N_28908,N_29670);
xnor UO_728 (O_728,N_29151,N_28915);
nand UO_729 (O_729,N_29392,N_28800);
nor UO_730 (O_730,N_29389,N_29061);
or UO_731 (O_731,N_29479,N_29086);
xnor UO_732 (O_732,N_28943,N_29938);
or UO_733 (O_733,N_29911,N_29321);
nand UO_734 (O_734,N_29293,N_29173);
and UO_735 (O_735,N_29882,N_29075);
nor UO_736 (O_736,N_29520,N_29950);
xnor UO_737 (O_737,N_28869,N_28816);
and UO_738 (O_738,N_28888,N_29854);
nor UO_739 (O_739,N_29183,N_28806);
nor UO_740 (O_740,N_29926,N_28939);
nand UO_741 (O_741,N_29661,N_28953);
nand UO_742 (O_742,N_29095,N_29897);
xnor UO_743 (O_743,N_29738,N_29122);
nand UO_744 (O_744,N_29139,N_29479);
or UO_745 (O_745,N_29471,N_29016);
and UO_746 (O_746,N_29965,N_29991);
and UO_747 (O_747,N_29879,N_29219);
and UO_748 (O_748,N_29784,N_29296);
nand UO_749 (O_749,N_29500,N_29816);
and UO_750 (O_750,N_29900,N_29012);
nor UO_751 (O_751,N_29123,N_29622);
or UO_752 (O_752,N_29207,N_28894);
nand UO_753 (O_753,N_29899,N_29822);
and UO_754 (O_754,N_29658,N_29577);
and UO_755 (O_755,N_29841,N_29905);
nand UO_756 (O_756,N_29644,N_29183);
and UO_757 (O_757,N_29761,N_28961);
nor UO_758 (O_758,N_29928,N_29739);
xor UO_759 (O_759,N_28895,N_29605);
and UO_760 (O_760,N_29854,N_29490);
or UO_761 (O_761,N_28974,N_29779);
nor UO_762 (O_762,N_29292,N_29316);
xor UO_763 (O_763,N_29658,N_29059);
nor UO_764 (O_764,N_29088,N_28945);
xor UO_765 (O_765,N_29768,N_29095);
or UO_766 (O_766,N_29519,N_29831);
xor UO_767 (O_767,N_29777,N_29900);
nand UO_768 (O_768,N_29908,N_29266);
or UO_769 (O_769,N_29349,N_29856);
or UO_770 (O_770,N_29324,N_29292);
nand UO_771 (O_771,N_29088,N_29124);
and UO_772 (O_772,N_29876,N_29300);
nand UO_773 (O_773,N_28970,N_29460);
nand UO_774 (O_774,N_28829,N_29968);
nor UO_775 (O_775,N_29503,N_29166);
xnor UO_776 (O_776,N_29090,N_29173);
or UO_777 (O_777,N_29688,N_29043);
xnor UO_778 (O_778,N_29488,N_29673);
xor UO_779 (O_779,N_28985,N_29861);
nand UO_780 (O_780,N_29787,N_29127);
or UO_781 (O_781,N_29117,N_28800);
or UO_782 (O_782,N_29677,N_29620);
and UO_783 (O_783,N_28915,N_29828);
or UO_784 (O_784,N_28993,N_29643);
and UO_785 (O_785,N_29354,N_29400);
or UO_786 (O_786,N_29495,N_29732);
xor UO_787 (O_787,N_29707,N_29961);
and UO_788 (O_788,N_29447,N_28962);
nor UO_789 (O_789,N_29658,N_29665);
or UO_790 (O_790,N_29851,N_29087);
xor UO_791 (O_791,N_29711,N_29443);
nor UO_792 (O_792,N_29999,N_28840);
nand UO_793 (O_793,N_29818,N_28966);
xor UO_794 (O_794,N_29534,N_29294);
nand UO_795 (O_795,N_29667,N_29052);
nand UO_796 (O_796,N_28999,N_29729);
or UO_797 (O_797,N_29855,N_29327);
nor UO_798 (O_798,N_29501,N_29745);
or UO_799 (O_799,N_29673,N_28926);
nor UO_800 (O_800,N_29374,N_29040);
xnor UO_801 (O_801,N_29683,N_29433);
or UO_802 (O_802,N_29137,N_29614);
xor UO_803 (O_803,N_28967,N_29579);
xnor UO_804 (O_804,N_29097,N_29275);
nor UO_805 (O_805,N_29590,N_29797);
nor UO_806 (O_806,N_29922,N_28895);
and UO_807 (O_807,N_29464,N_29797);
nor UO_808 (O_808,N_29788,N_29669);
nand UO_809 (O_809,N_29863,N_28840);
nor UO_810 (O_810,N_29012,N_29452);
or UO_811 (O_811,N_29684,N_29884);
and UO_812 (O_812,N_28944,N_29846);
nor UO_813 (O_813,N_29251,N_29192);
nor UO_814 (O_814,N_29447,N_29520);
nand UO_815 (O_815,N_29069,N_29615);
nand UO_816 (O_816,N_29958,N_29742);
or UO_817 (O_817,N_29645,N_29594);
nand UO_818 (O_818,N_29181,N_29527);
nor UO_819 (O_819,N_28888,N_29478);
nor UO_820 (O_820,N_29154,N_28903);
nor UO_821 (O_821,N_29397,N_29984);
and UO_822 (O_822,N_28888,N_29265);
and UO_823 (O_823,N_29630,N_29649);
xnor UO_824 (O_824,N_29319,N_29633);
xnor UO_825 (O_825,N_29016,N_28846);
nand UO_826 (O_826,N_29326,N_29494);
or UO_827 (O_827,N_29736,N_29497);
or UO_828 (O_828,N_29798,N_29952);
or UO_829 (O_829,N_29145,N_29987);
nor UO_830 (O_830,N_29974,N_29540);
and UO_831 (O_831,N_29824,N_29205);
nor UO_832 (O_832,N_29660,N_29231);
xnor UO_833 (O_833,N_29102,N_29839);
nand UO_834 (O_834,N_28961,N_28901);
or UO_835 (O_835,N_29397,N_29699);
nand UO_836 (O_836,N_29240,N_29161);
or UO_837 (O_837,N_29079,N_29727);
xor UO_838 (O_838,N_29576,N_29711);
xnor UO_839 (O_839,N_29996,N_29470);
and UO_840 (O_840,N_29140,N_29518);
or UO_841 (O_841,N_29389,N_29191);
nand UO_842 (O_842,N_29436,N_29588);
nor UO_843 (O_843,N_29119,N_29431);
nor UO_844 (O_844,N_29323,N_29070);
nor UO_845 (O_845,N_29002,N_29371);
nand UO_846 (O_846,N_29276,N_29094);
xnor UO_847 (O_847,N_28814,N_29861);
and UO_848 (O_848,N_29202,N_29633);
xnor UO_849 (O_849,N_28984,N_29785);
nor UO_850 (O_850,N_29851,N_29708);
xor UO_851 (O_851,N_29140,N_29993);
and UO_852 (O_852,N_29027,N_28873);
nand UO_853 (O_853,N_29849,N_29320);
nand UO_854 (O_854,N_29186,N_29169);
xor UO_855 (O_855,N_28877,N_29681);
nor UO_856 (O_856,N_29055,N_29622);
nand UO_857 (O_857,N_29849,N_29579);
or UO_858 (O_858,N_28808,N_29679);
nor UO_859 (O_859,N_29095,N_29637);
xor UO_860 (O_860,N_29643,N_29705);
xnor UO_861 (O_861,N_29299,N_29573);
nor UO_862 (O_862,N_29788,N_29455);
and UO_863 (O_863,N_29867,N_29833);
nand UO_864 (O_864,N_28962,N_29282);
and UO_865 (O_865,N_28984,N_29060);
nor UO_866 (O_866,N_29170,N_29175);
nand UO_867 (O_867,N_29020,N_29038);
nand UO_868 (O_868,N_29841,N_29545);
nand UO_869 (O_869,N_29318,N_29021);
and UO_870 (O_870,N_29428,N_29461);
and UO_871 (O_871,N_29757,N_29954);
xnor UO_872 (O_872,N_29882,N_29094);
and UO_873 (O_873,N_28901,N_28951);
and UO_874 (O_874,N_29713,N_29442);
nor UO_875 (O_875,N_29714,N_28920);
and UO_876 (O_876,N_29616,N_29189);
nor UO_877 (O_877,N_28882,N_29949);
xnor UO_878 (O_878,N_29706,N_29013);
or UO_879 (O_879,N_29359,N_29424);
and UO_880 (O_880,N_29344,N_29389);
nand UO_881 (O_881,N_29828,N_29260);
xnor UO_882 (O_882,N_29052,N_29189);
and UO_883 (O_883,N_29926,N_29081);
xor UO_884 (O_884,N_29580,N_28937);
and UO_885 (O_885,N_29132,N_29436);
nor UO_886 (O_886,N_29529,N_29688);
xor UO_887 (O_887,N_29039,N_29067);
xnor UO_888 (O_888,N_29810,N_28943);
xnor UO_889 (O_889,N_29137,N_29191);
and UO_890 (O_890,N_29894,N_29834);
nor UO_891 (O_891,N_29850,N_29660);
nand UO_892 (O_892,N_29455,N_29326);
nand UO_893 (O_893,N_28823,N_29235);
and UO_894 (O_894,N_29176,N_29615);
xnor UO_895 (O_895,N_29504,N_28992);
and UO_896 (O_896,N_29442,N_29962);
nor UO_897 (O_897,N_29885,N_29252);
xnor UO_898 (O_898,N_29503,N_28969);
and UO_899 (O_899,N_29185,N_29785);
nand UO_900 (O_900,N_28885,N_29976);
nand UO_901 (O_901,N_29227,N_29203);
nor UO_902 (O_902,N_29440,N_29057);
xnor UO_903 (O_903,N_29627,N_28876);
nor UO_904 (O_904,N_29617,N_29658);
nor UO_905 (O_905,N_29269,N_29440);
or UO_906 (O_906,N_29067,N_29565);
or UO_907 (O_907,N_29018,N_29027);
xnor UO_908 (O_908,N_29426,N_29979);
or UO_909 (O_909,N_28941,N_29282);
xnor UO_910 (O_910,N_29466,N_29523);
xnor UO_911 (O_911,N_29704,N_29201);
xor UO_912 (O_912,N_29210,N_29203);
xor UO_913 (O_913,N_29061,N_29143);
nand UO_914 (O_914,N_29251,N_29167);
and UO_915 (O_915,N_29987,N_29185);
or UO_916 (O_916,N_29734,N_29132);
or UO_917 (O_917,N_29587,N_29104);
or UO_918 (O_918,N_29765,N_29465);
or UO_919 (O_919,N_28977,N_29705);
nand UO_920 (O_920,N_29680,N_29154);
or UO_921 (O_921,N_29922,N_29486);
nor UO_922 (O_922,N_29754,N_29943);
nor UO_923 (O_923,N_28893,N_29676);
nand UO_924 (O_924,N_28977,N_29991);
or UO_925 (O_925,N_29620,N_29794);
and UO_926 (O_926,N_29829,N_29861);
xnor UO_927 (O_927,N_29769,N_28922);
and UO_928 (O_928,N_29395,N_29943);
nand UO_929 (O_929,N_29928,N_29072);
and UO_930 (O_930,N_29769,N_29560);
nand UO_931 (O_931,N_29078,N_28980);
or UO_932 (O_932,N_29587,N_29679);
or UO_933 (O_933,N_29900,N_29218);
and UO_934 (O_934,N_28995,N_29474);
nor UO_935 (O_935,N_29021,N_29559);
nor UO_936 (O_936,N_29080,N_29286);
and UO_937 (O_937,N_29537,N_28952);
or UO_938 (O_938,N_28948,N_29333);
and UO_939 (O_939,N_29091,N_29749);
or UO_940 (O_940,N_29809,N_29435);
and UO_941 (O_941,N_29911,N_29424);
nand UO_942 (O_942,N_29331,N_29404);
or UO_943 (O_943,N_28851,N_29518);
or UO_944 (O_944,N_29673,N_28901);
nor UO_945 (O_945,N_29974,N_29641);
xnor UO_946 (O_946,N_28807,N_29759);
or UO_947 (O_947,N_28826,N_29197);
xnor UO_948 (O_948,N_29083,N_28952);
or UO_949 (O_949,N_29511,N_29219);
nor UO_950 (O_950,N_29526,N_29041);
nor UO_951 (O_951,N_29211,N_29519);
and UO_952 (O_952,N_29691,N_29884);
nor UO_953 (O_953,N_29298,N_29602);
xnor UO_954 (O_954,N_29106,N_29741);
or UO_955 (O_955,N_29619,N_29048);
or UO_956 (O_956,N_29772,N_28906);
xnor UO_957 (O_957,N_29042,N_29684);
nor UO_958 (O_958,N_29742,N_29305);
nand UO_959 (O_959,N_29152,N_29241);
nor UO_960 (O_960,N_29524,N_29229);
and UO_961 (O_961,N_29329,N_29463);
nor UO_962 (O_962,N_29925,N_29309);
nand UO_963 (O_963,N_29194,N_29571);
xnor UO_964 (O_964,N_29418,N_29047);
or UO_965 (O_965,N_28978,N_29036);
or UO_966 (O_966,N_28958,N_29093);
xnor UO_967 (O_967,N_29759,N_29098);
or UO_968 (O_968,N_29787,N_28857);
and UO_969 (O_969,N_29573,N_29776);
or UO_970 (O_970,N_29483,N_28964);
nand UO_971 (O_971,N_28877,N_29180);
xnor UO_972 (O_972,N_29710,N_29901);
and UO_973 (O_973,N_29918,N_29535);
nand UO_974 (O_974,N_29653,N_29140);
and UO_975 (O_975,N_29383,N_29276);
xnor UO_976 (O_976,N_29893,N_29713);
nand UO_977 (O_977,N_29718,N_29016);
nor UO_978 (O_978,N_29608,N_28877);
or UO_979 (O_979,N_28806,N_28846);
nor UO_980 (O_980,N_29866,N_29470);
and UO_981 (O_981,N_29859,N_29893);
xor UO_982 (O_982,N_28865,N_28912);
and UO_983 (O_983,N_29957,N_29043);
and UO_984 (O_984,N_28850,N_29957);
nand UO_985 (O_985,N_29824,N_29915);
nand UO_986 (O_986,N_29751,N_29776);
or UO_987 (O_987,N_29317,N_29124);
xnor UO_988 (O_988,N_28841,N_29952);
nand UO_989 (O_989,N_29821,N_29112);
nand UO_990 (O_990,N_29502,N_29576);
and UO_991 (O_991,N_29425,N_29915);
nand UO_992 (O_992,N_29729,N_29875);
xor UO_993 (O_993,N_29241,N_29661);
nand UO_994 (O_994,N_29438,N_28968);
or UO_995 (O_995,N_29901,N_29319);
nor UO_996 (O_996,N_28989,N_28922);
nor UO_997 (O_997,N_29988,N_29081);
nor UO_998 (O_998,N_29974,N_29735);
and UO_999 (O_999,N_28931,N_29954);
nand UO_1000 (O_1000,N_28813,N_29574);
nor UO_1001 (O_1001,N_29802,N_29516);
or UO_1002 (O_1002,N_29955,N_29956);
nand UO_1003 (O_1003,N_28852,N_29890);
nand UO_1004 (O_1004,N_29164,N_29387);
nor UO_1005 (O_1005,N_29266,N_29054);
or UO_1006 (O_1006,N_29643,N_29911);
or UO_1007 (O_1007,N_28820,N_29527);
nor UO_1008 (O_1008,N_29224,N_29810);
or UO_1009 (O_1009,N_29925,N_29175);
and UO_1010 (O_1010,N_29165,N_29347);
nand UO_1011 (O_1011,N_29747,N_28955);
nand UO_1012 (O_1012,N_29206,N_29288);
xor UO_1013 (O_1013,N_28827,N_29082);
or UO_1014 (O_1014,N_29661,N_29986);
nand UO_1015 (O_1015,N_29047,N_29001);
xor UO_1016 (O_1016,N_29808,N_29230);
and UO_1017 (O_1017,N_29348,N_29931);
or UO_1018 (O_1018,N_29735,N_29902);
nand UO_1019 (O_1019,N_29920,N_29295);
and UO_1020 (O_1020,N_29061,N_28800);
and UO_1021 (O_1021,N_29847,N_29090);
and UO_1022 (O_1022,N_29473,N_29688);
or UO_1023 (O_1023,N_29222,N_28975);
nand UO_1024 (O_1024,N_28926,N_29714);
or UO_1025 (O_1025,N_29855,N_29544);
nand UO_1026 (O_1026,N_29588,N_29608);
or UO_1027 (O_1027,N_29710,N_29545);
nand UO_1028 (O_1028,N_29170,N_29411);
xor UO_1029 (O_1029,N_29095,N_29799);
and UO_1030 (O_1030,N_29918,N_29488);
nor UO_1031 (O_1031,N_29362,N_29359);
and UO_1032 (O_1032,N_29382,N_29274);
nor UO_1033 (O_1033,N_29425,N_29158);
xor UO_1034 (O_1034,N_29401,N_29818);
or UO_1035 (O_1035,N_29233,N_29845);
and UO_1036 (O_1036,N_29766,N_28805);
nor UO_1037 (O_1037,N_29462,N_29618);
and UO_1038 (O_1038,N_29079,N_29295);
and UO_1039 (O_1039,N_28884,N_28955);
or UO_1040 (O_1040,N_29126,N_29808);
nor UO_1041 (O_1041,N_29963,N_29887);
or UO_1042 (O_1042,N_29620,N_29461);
or UO_1043 (O_1043,N_28857,N_29474);
nor UO_1044 (O_1044,N_29774,N_29647);
and UO_1045 (O_1045,N_29592,N_29044);
nand UO_1046 (O_1046,N_29326,N_29692);
nand UO_1047 (O_1047,N_29079,N_29246);
and UO_1048 (O_1048,N_29741,N_29144);
xor UO_1049 (O_1049,N_29893,N_29954);
or UO_1050 (O_1050,N_29109,N_28993);
nand UO_1051 (O_1051,N_29701,N_28805);
xor UO_1052 (O_1052,N_29792,N_29453);
or UO_1053 (O_1053,N_28837,N_29112);
nand UO_1054 (O_1054,N_29674,N_29596);
nand UO_1055 (O_1055,N_28890,N_28954);
or UO_1056 (O_1056,N_29136,N_29981);
xor UO_1057 (O_1057,N_29719,N_28983);
xnor UO_1058 (O_1058,N_28852,N_29850);
xor UO_1059 (O_1059,N_29422,N_29068);
nand UO_1060 (O_1060,N_29086,N_29745);
or UO_1061 (O_1061,N_29586,N_28927);
nand UO_1062 (O_1062,N_29711,N_29804);
and UO_1063 (O_1063,N_29614,N_29529);
xor UO_1064 (O_1064,N_29122,N_28939);
nand UO_1065 (O_1065,N_28900,N_29141);
or UO_1066 (O_1066,N_29065,N_29359);
or UO_1067 (O_1067,N_29202,N_29724);
nand UO_1068 (O_1068,N_28884,N_29532);
nor UO_1069 (O_1069,N_29684,N_29844);
xnor UO_1070 (O_1070,N_29166,N_29225);
nand UO_1071 (O_1071,N_29601,N_29066);
xor UO_1072 (O_1072,N_29863,N_29810);
xor UO_1073 (O_1073,N_29980,N_29225);
and UO_1074 (O_1074,N_29690,N_29279);
and UO_1075 (O_1075,N_29499,N_29276);
nand UO_1076 (O_1076,N_28842,N_29768);
and UO_1077 (O_1077,N_29464,N_29544);
nor UO_1078 (O_1078,N_29632,N_29127);
nand UO_1079 (O_1079,N_29935,N_29918);
nand UO_1080 (O_1080,N_29556,N_28884);
nand UO_1081 (O_1081,N_29342,N_29910);
nand UO_1082 (O_1082,N_29865,N_29419);
or UO_1083 (O_1083,N_29013,N_29050);
or UO_1084 (O_1084,N_29371,N_28819);
xnor UO_1085 (O_1085,N_29983,N_29465);
nor UO_1086 (O_1086,N_28898,N_29204);
nand UO_1087 (O_1087,N_29107,N_28880);
xnor UO_1088 (O_1088,N_29877,N_29296);
xor UO_1089 (O_1089,N_29940,N_29555);
and UO_1090 (O_1090,N_28887,N_29331);
nand UO_1091 (O_1091,N_29016,N_28931);
nor UO_1092 (O_1092,N_29775,N_29752);
nand UO_1093 (O_1093,N_29828,N_28817);
and UO_1094 (O_1094,N_28855,N_29193);
nor UO_1095 (O_1095,N_29023,N_29993);
and UO_1096 (O_1096,N_29779,N_28978);
nor UO_1097 (O_1097,N_28885,N_29060);
nand UO_1098 (O_1098,N_29023,N_29101);
nand UO_1099 (O_1099,N_29494,N_28958);
or UO_1100 (O_1100,N_29260,N_28923);
nand UO_1101 (O_1101,N_29475,N_29085);
and UO_1102 (O_1102,N_28913,N_29084);
or UO_1103 (O_1103,N_29708,N_29839);
and UO_1104 (O_1104,N_29468,N_29048);
nand UO_1105 (O_1105,N_29621,N_28825);
or UO_1106 (O_1106,N_29673,N_29314);
nor UO_1107 (O_1107,N_29891,N_29536);
and UO_1108 (O_1108,N_29975,N_29077);
nand UO_1109 (O_1109,N_29645,N_29698);
nor UO_1110 (O_1110,N_28830,N_29909);
xor UO_1111 (O_1111,N_29073,N_29256);
xor UO_1112 (O_1112,N_29398,N_29459);
or UO_1113 (O_1113,N_28860,N_29694);
nor UO_1114 (O_1114,N_29442,N_29275);
nor UO_1115 (O_1115,N_29136,N_29694);
and UO_1116 (O_1116,N_29837,N_29719);
nor UO_1117 (O_1117,N_29742,N_29637);
nor UO_1118 (O_1118,N_28869,N_29634);
or UO_1119 (O_1119,N_28928,N_29733);
nand UO_1120 (O_1120,N_29952,N_29643);
xor UO_1121 (O_1121,N_29015,N_29727);
or UO_1122 (O_1122,N_29888,N_29625);
and UO_1123 (O_1123,N_29250,N_29648);
nand UO_1124 (O_1124,N_29892,N_29453);
xor UO_1125 (O_1125,N_29944,N_29868);
nand UO_1126 (O_1126,N_29904,N_29705);
nor UO_1127 (O_1127,N_29570,N_29528);
and UO_1128 (O_1128,N_29701,N_28953);
xor UO_1129 (O_1129,N_29824,N_29924);
xnor UO_1130 (O_1130,N_28990,N_29591);
and UO_1131 (O_1131,N_29381,N_28869);
xor UO_1132 (O_1132,N_29129,N_29533);
nor UO_1133 (O_1133,N_29291,N_29232);
and UO_1134 (O_1134,N_29694,N_29566);
nand UO_1135 (O_1135,N_29815,N_29269);
xnor UO_1136 (O_1136,N_29074,N_29382);
nor UO_1137 (O_1137,N_29604,N_29356);
xnor UO_1138 (O_1138,N_29908,N_29972);
xor UO_1139 (O_1139,N_29199,N_29539);
or UO_1140 (O_1140,N_29234,N_29411);
and UO_1141 (O_1141,N_28934,N_28926);
xnor UO_1142 (O_1142,N_28953,N_29078);
nor UO_1143 (O_1143,N_28979,N_28909);
and UO_1144 (O_1144,N_29117,N_28813);
and UO_1145 (O_1145,N_29128,N_29484);
or UO_1146 (O_1146,N_29238,N_29525);
nand UO_1147 (O_1147,N_29487,N_28918);
or UO_1148 (O_1148,N_29287,N_29849);
nor UO_1149 (O_1149,N_29697,N_29672);
nand UO_1150 (O_1150,N_29487,N_29266);
nand UO_1151 (O_1151,N_29736,N_29935);
nor UO_1152 (O_1152,N_29985,N_29360);
nor UO_1153 (O_1153,N_29343,N_29674);
and UO_1154 (O_1154,N_29837,N_29554);
xor UO_1155 (O_1155,N_29047,N_29378);
xor UO_1156 (O_1156,N_28941,N_29337);
and UO_1157 (O_1157,N_29306,N_29295);
nor UO_1158 (O_1158,N_29742,N_29183);
nand UO_1159 (O_1159,N_29906,N_29837);
nand UO_1160 (O_1160,N_28974,N_29020);
or UO_1161 (O_1161,N_29811,N_28998);
xor UO_1162 (O_1162,N_29495,N_29001);
nand UO_1163 (O_1163,N_29173,N_29291);
xnor UO_1164 (O_1164,N_29615,N_29837);
nand UO_1165 (O_1165,N_29738,N_29231);
nand UO_1166 (O_1166,N_29316,N_29980);
and UO_1167 (O_1167,N_28866,N_28820);
nand UO_1168 (O_1168,N_28804,N_29387);
and UO_1169 (O_1169,N_28879,N_29705);
nand UO_1170 (O_1170,N_28886,N_29620);
or UO_1171 (O_1171,N_29386,N_29505);
and UO_1172 (O_1172,N_28913,N_29138);
and UO_1173 (O_1173,N_28880,N_29016);
or UO_1174 (O_1174,N_29886,N_28822);
nand UO_1175 (O_1175,N_29210,N_29248);
nor UO_1176 (O_1176,N_29627,N_29928);
xor UO_1177 (O_1177,N_29258,N_29297);
nand UO_1178 (O_1178,N_29624,N_29090);
or UO_1179 (O_1179,N_29081,N_29293);
xnor UO_1180 (O_1180,N_29434,N_29402);
and UO_1181 (O_1181,N_28916,N_29083);
and UO_1182 (O_1182,N_29803,N_29173);
nand UO_1183 (O_1183,N_29574,N_29106);
nor UO_1184 (O_1184,N_28854,N_28964);
nor UO_1185 (O_1185,N_29232,N_29250);
nand UO_1186 (O_1186,N_29112,N_29766);
xor UO_1187 (O_1187,N_29101,N_29915);
or UO_1188 (O_1188,N_29482,N_29872);
and UO_1189 (O_1189,N_29102,N_29125);
xor UO_1190 (O_1190,N_28837,N_28879);
and UO_1191 (O_1191,N_29067,N_29583);
or UO_1192 (O_1192,N_29013,N_29436);
nand UO_1193 (O_1193,N_29577,N_29926);
nand UO_1194 (O_1194,N_29962,N_28818);
or UO_1195 (O_1195,N_29831,N_29399);
xor UO_1196 (O_1196,N_29946,N_28925);
and UO_1197 (O_1197,N_29519,N_29208);
or UO_1198 (O_1198,N_29732,N_29867);
and UO_1199 (O_1199,N_29909,N_29329);
xnor UO_1200 (O_1200,N_29995,N_29032);
nand UO_1201 (O_1201,N_29735,N_29615);
xor UO_1202 (O_1202,N_29206,N_29148);
nor UO_1203 (O_1203,N_29782,N_29201);
nand UO_1204 (O_1204,N_29726,N_29306);
and UO_1205 (O_1205,N_28950,N_29130);
nand UO_1206 (O_1206,N_29714,N_29671);
nor UO_1207 (O_1207,N_29371,N_28885);
nand UO_1208 (O_1208,N_29518,N_29288);
xor UO_1209 (O_1209,N_29492,N_29035);
or UO_1210 (O_1210,N_29627,N_28981);
nand UO_1211 (O_1211,N_29864,N_29078);
xor UO_1212 (O_1212,N_29802,N_29310);
nor UO_1213 (O_1213,N_29227,N_29811);
or UO_1214 (O_1214,N_29956,N_29133);
and UO_1215 (O_1215,N_29610,N_28972);
or UO_1216 (O_1216,N_28943,N_28979);
or UO_1217 (O_1217,N_29367,N_29651);
or UO_1218 (O_1218,N_29932,N_29047);
xnor UO_1219 (O_1219,N_28982,N_28828);
xor UO_1220 (O_1220,N_29826,N_29758);
nor UO_1221 (O_1221,N_29620,N_28988);
or UO_1222 (O_1222,N_29813,N_29256);
or UO_1223 (O_1223,N_29127,N_29259);
nor UO_1224 (O_1224,N_29213,N_29336);
and UO_1225 (O_1225,N_29593,N_29733);
xnor UO_1226 (O_1226,N_29280,N_29695);
and UO_1227 (O_1227,N_29286,N_29899);
xnor UO_1228 (O_1228,N_29216,N_29272);
nand UO_1229 (O_1229,N_29780,N_29865);
and UO_1230 (O_1230,N_28826,N_28943);
or UO_1231 (O_1231,N_29094,N_29413);
and UO_1232 (O_1232,N_28995,N_29798);
nor UO_1233 (O_1233,N_29876,N_29096);
nand UO_1234 (O_1234,N_29396,N_29469);
xor UO_1235 (O_1235,N_29294,N_29232);
nor UO_1236 (O_1236,N_28911,N_28956);
xnor UO_1237 (O_1237,N_29299,N_28941);
nor UO_1238 (O_1238,N_29072,N_29557);
nand UO_1239 (O_1239,N_29620,N_29305);
nand UO_1240 (O_1240,N_28915,N_28973);
or UO_1241 (O_1241,N_29307,N_29581);
nand UO_1242 (O_1242,N_28905,N_29179);
and UO_1243 (O_1243,N_29997,N_29093);
and UO_1244 (O_1244,N_28809,N_29464);
or UO_1245 (O_1245,N_29771,N_29980);
or UO_1246 (O_1246,N_29571,N_29169);
or UO_1247 (O_1247,N_29894,N_29627);
or UO_1248 (O_1248,N_28887,N_29239);
or UO_1249 (O_1249,N_29976,N_29848);
nor UO_1250 (O_1250,N_29638,N_29278);
or UO_1251 (O_1251,N_29736,N_29878);
nand UO_1252 (O_1252,N_28882,N_29916);
nor UO_1253 (O_1253,N_29607,N_28805);
nor UO_1254 (O_1254,N_29139,N_29287);
and UO_1255 (O_1255,N_29744,N_29311);
nand UO_1256 (O_1256,N_29193,N_28816);
or UO_1257 (O_1257,N_28851,N_28977);
nand UO_1258 (O_1258,N_29212,N_29792);
nand UO_1259 (O_1259,N_29997,N_29632);
nand UO_1260 (O_1260,N_29261,N_29292);
nand UO_1261 (O_1261,N_29076,N_29822);
nand UO_1262 (O_1262,N_28812,N_29779);
nor UO_1263 (O_1263,N_29588,N_29480);
or UO_1264 (O_1264,N_29820,N_29711);
nand UO_1265 (O_1265,N_28858,N_29124);
or UO_1266 (O_1266,N_29758,N_29559);
nor UO_1267 (O_1267,N_29449,N_29452);
nand UO_1268 (O_1268,N_29594,N_28845);
or UO_1269 (O_1269,N_29251,N_29155);
xnor UO_1270 (O_1270,N_29965,N_29546);
nor UO_1271 (O_1271,N_29002,N_29093);
nor UO_1272 (O_1272,N_29799,N_29318);
nor UO_1273 (O_1273,N_28911,N_29568);
nor UO_1274 (O_1274,N_28960,N_29050);
or UO_1275 (O_1275,N_29821,N_29288);
and UO_1276 (O_1276,N_29987,N_29542);
or UO_1277 (O_1277,N_29078,N_28938);
nor UO_1278 (O_1278,N_29836,N_29183);
nand UO_1279 (O_1279,N_29238,N_28910);
and UO_1280 (O_1280,N_29552,N_29727);
nor UO_1281 (O_1281,N_29380,N_29411);
nor UO_1282 (O_1282,N_29559,N_29038);
nand UO_1283 (O_1283,N_28919,N_29114);
or UO_1284 (O_1284,N_29483,N_29459);
and UO_1285 (O_1285,N_29599,N_29341);
or UO_1286 (O_1286,N_28996,N_29978);
or UO_1287 (O_1287,N_29318,N_28903);
nand UO_1288 (O_1288,N_29504,N_29150);
xnor UO_1289 (O_1289,N_29590,N_28904);
nor UO_1290 (O_1290,N_28965,N_29706);
or UO_1291 (O_1291,N_28947,N_29005);
nand UO_1292 (O_1292,N_29945,N_29725);
xnor UO_1293 (O_1293,N_29810,N_29914);
nor UO_1294 (O_1294,N_29220,N_29238);
or UO_1295 (O_1295,N_29766,N_29741);
xor UO_1296 (O_1296,N_28964,N_29136);
xor UO_1297 (O_1297,N_29774,N_29176);
nand UO_1298 (O_1298,N_29560,N_29588);
and UO_1299 (O_1299,N_29698,N_29630);
and UO_1300 (O_1300,N_29231,N_29858);
and UO_1301 (O_1301,N_28827,N_29858);
xor UO_1302 (O_1302,N_29469,N_28921);
or UO_1303 (O_1303,N_28823,N_28854);
and UO_1304 (O_1304,N_28893,N_29597);
nor UO_1305 (O_1305,N_29657,N_29978);
nor UO_1306 (O_1306,N_29852,N_29458);
nor UO_1307 (O_1307,N_29483,N_28921);
or UO_1308 (O_1308,N_29883,N_28818);
or UO_1309 (O_1309,N_29376,N_29604);
xnor UO_1310 (O_1310,N_29454,N_29808);
nand UO_1311 (O_1311,N_29242,N_29271);
xor UO_1312 (O_1312,N_28896,N_29581);
or UO_1313 (O_1313,N_29152,N_29008);
nor UO_1314 (O_1314,N_28895,N_29394);
nand UO_1315 (O_1315,N_29618,N_29746);
xnor UO_1316 (O_1316,N_29450,N_29503);
nor UO_1317 (O_1317,N_29672,N_29428);
xnor UO_1318 (O_1318,N_29810,N_29249);
nor UO_1319 (O_1319,N_29234,N_29586);
xor UO_1320 (O_1320,N_29262,N_29702);
nand UO_1321 (O_1321,N_29888,N_29005);
or UO_1322 (O_1322,N_29933,N_29374);
nor UO_1323 (O_1323,N_28957,N_29480);
xor UO_1324 (O_1324,N_29419,N_29925);
xor UO_1325 (O_1325,N_29769,N_29007);
nor UO_1326 (O_1326,N_29021,N_29812);
nand UO_1327 (O_1327,N_29377,N_29079);
nor UO_1328 (O_1328,N_29346,N_29354);
and UO_1329 (O_1329,N_29761,N_28870);
xor UO_1330 (O_1330,N_29451,N_29086);
or UO_1331 (O_1331,N_29294,N_29529);
nand UO_1332 (O_1332,N_29264,N_29546);
or UO_1333 (O_1333,N_28964,N_29282);
nand UO_1334 (O_1334,N_29497,N_29761);
nand UO_1335 (O_1335,N_29444,N_29076);
or UO_1336 (O_1336,N_28801,N_29641);
or UO_1337 (O_1337,N_28932,N_29632);
or UO_1338 (O_1338,N_29492,N_29585);
and UO_1339 (O_1339,N_29865,N_29685);
xor UO_1340 (O_1340,N_29856,N_29402);
nor UO_1341 (O_1341,N_29861,N_28990);
xnor UO_1342 (O_1342,N_29932,N_29292);
nor UO_1343 (O_1343,N_29689,N_29955);
nand UO_1344 (O_1344,N_28987,N_29158);
nor UO_1345 (O_1345,N_29223,N_29379);
or UO_1346 (O_1346,N_29184,N_29098);
nor UO_1347 (O_1347,N_29020,N_29985);
or UO_1348 (O_1348,N_29676,N_29946);
xor UO_1349 (O_1349,N_29163,N_29974);
and UO_1350 (O_1350,N_29456,N_29977);
nor UO_1351 (O_1351,N_28917,N_29734);
and UO_1352 (O_1352,N_29551,N_29198);
xnor UO_1353 (O_1353,N_29276,N_29515);
xor UO_1354 (O_1354,N_28933,N_29777);
nor UO_1355 (O_1355,N_29551,N_29579);
and UO_1356 (O_1356,N_29211,N_29804);
or UO_1357 (O_1357,N_29340,N_29819);
nand UO_1358 (O_1358,N_29990,N_29307);
xor UO_1359 (O_1359,N_29311,N_29486);
or UO_1360 (O_1360,N_28835,N_29731);
xor UO_1361 (O_1361,N_28805,N_29008);
nor UO_1362 (O_1362,N_29240,N_29754);
nor UO_1363 (O_1363,N_29500,N_29631);
xor UO_1364 (O_1364,N_29645,N_29695);
or UO_1365 (O_1365,N_29878,N_29777);
and UO_1366 (O_1366,N_29837,N_29420);
or UO_1367 (O_1367,N_29281,N_29819);
and UO_1368 (O_1368,N_29111,N_29457);
or UO_1369 (O_1369,N_29846,N_29646);
nor UO_1370 (O_1370,N_29864,N_29690);
xor UO_1371 (O_1371,N_29181,N_29032);
nand UO_1372 (O_1372,N_29283,N_29405);
and UO_1373 (O_1373,N_28890,N_29714);
xor UO_1374 (O_1374,N_29903,N_28949);
and UO_1375 (O_1375,N_29294,N_29982);
xnor UO_1376 (O_1376,N_29549,N_29653);
and UO_1377 (O_1377,N_29120,N_29599);
nor UO_1378 (O_1378,N_29173,N_28812);
xor UO_1379 (O_1379,N_28880,N_29695);
xor UO_1380 (O_1380,N_29311,N_29657);
nand UO_1381 (O_1381,N_29767,N_28870);
nand UO_1382 (O_1382,N_29433,N_29293);
xor UO_1383 (O_1383,N_29808,N_28967);
nor UO_1384 (O_1384,N_29637,N_29836);
or UO_1385 (O_1385,N_28874,N_29430);
xnor UO_1386 (O_1386,N_28996,N_29984);
and UO_1387 (O_1387,N_29435,N_29032);
nor UO_1388 (O_1388,N_28867,N_29081);
and UO_1389 (O_1389,N_29458,N_29910);
nand UO_1390 (O_1390,N_29598,N_29086);
nand UO_1391 (O_1391,N_29991,N_29271);
nand UO_1392 (O_1392,N_29490,N_29068);
or UO_1393 (O_1393,N_29603,N_28867);
nor UO_1394 (O_1394,N_29126,N_29498);
nor UO_1395 (O_1395,N_29620,N_29315);
xor UO_1396 (O_1396,N_28975,N_29954);
xor UO_1397 (O_1397,N_28900,N_29814);
xor UO_1398 (O_1398,N_29535,N_29480);
nand UO_1399 (O_1399,N_28837,N_29216);
and UO_1400 (O_1400,N_29727,N_29006);
nand UO_1401 (O_1401,N_29409,N_29724);
nor UO_1402 (O_1402,N_29832,N_29897);
nor UO_1403 (O_1403,N_28881,N_28826);
and UO_1404 (O_1404,N_28826,N_29681);
nor UO_1405 (O_1405,N_29790,N_29184);
xor UO_1406 (O_1406,N_29118,N_29748);
xor UO_1407 (O_1407,N_29753,N_29309);
or UO_1408 (O_1408,N_29622,N_29064);
or UO_1409 (O_1409,N_29683,N_29513);
xnor UO_1410 (O_1410,N_28927,N_29690);
nor UO_1411 (O_1411,N_29799,N_29229);
and UO_1412 (O_1412,N_29481,N_28806);
nor UO_1413 (O_1413,N_29677,N_29496);
or UO_1414 (O_1414,N_29109,N_29991);
and UO_1415 (O_1415,N_29230,N_29839);
nor UO_1416 (O_1416,N_29735,N_29422);
and UO_1417 (O_1417,N_29405,N_29837);
xor UO_1418 (O_1418,N_28988,N_29998);
or UO_1419 (O_1419,N_29406,N_29240);
nor UO_1420 (O_1420,N_29213,N_29196);
or UO_1421 (O_1421,N_29233,N_29612);
or UO_1422 (O_1422,N_29650,N_29250);
nand UO_1423 (O_1423,N_29215,N_29474);
nor UO_1424 (O_1424,N_28801,N_29124);
xor UO_1425 (O_1425,N_29257,N_29566);
xnor UO_1426 (O_1426,N_29887,N_29429);
or UO_1427 (O_1427,N_29829,N_29373);
and UO_1428 (O_1428,N_29467,N_29301);
nor UO_1429 (O_1429,N_29752,N_29980);
or UO_1430 (O_1430,N_29880,N_29489);
xor UO_1431 (O_1431,N_29894,N_29897);
nor UO_1432 (O_1432,N_28912,N_29050);
nand UO_1433 (O_1433,N_28920,N_29801);
or UO_1434 (O_1434,N_29557,N_29514);
or UO_1435 (O_1435,N_29068,N_29033);
and UO_1436 (O_1436,N_29792,N_29215);
xor UO_1437 (O_1437,N_28802,N_29133);
and UO_1438 (O_1438,N_29245,N_29943);
nand UO_1439 (O_1439,N_29347,N_29389);
nor UO_1440 (O_1440,N_29184,N_29885);
or UO_1441 (O_1441,N_29331,N_29921);
xor UO_1442 (O_1442,N_29372,N_29649);
nand UO_1443 (O_1443,N_29720,N_29188);
or UO_1444 (O_1444,N_29320,N_28840);
nand UO_1445 (O_1445,N_28983,N_29401);
or UO_1446 (O_1446,N_29586,N_29627);
or UO_1447 (O_1447,N_28902,N_29965);
nand UO_1448 (O_1448,N_29547,N_29207);
and UO_1449 (O_1449,N_29942,N_29727);
and UO_1450 (O_1450,N_28887,N_29448);
xnor UO_1451 (O_1451,N_29795,N_29632);
xor UO_1452 (O_1452,N_29276,N_28838);
nor UO_1453 (O_1453,N_29948,N_28848);
nor UO_1454 (O_1454,N_28995,N_29286);
and UO_1455 (O_1455,N_29587,N_29299);
nor UO_1456 (O_1456,N_29305,N_29232);
nand UO_1457 (O_1457,N_29100,N_29536);
nor UO_1458 (O_1458,N_29867,N_29541);
xor UO_1459 (O_1459,N_29548,N_29139);
and UO_1460 (O_1460,N_29012,N_28904);
nand UO_1461 (O_1461,N_28904,N_28860);
nand UO_1462 (O_1462,N_29973,N_29023);
and UO_1463 (O_1463,N_29784,N_29537);
or UO_1464 (O_1464,N_29355,N_29562);
xnor UO_1465 (O_1465,N_29760,N_28818);
nor UO_1466 (O_1466,N_29495,N_28824);
xnor UO_1467 (O_1467,N_29987,N_29274);
xor UO_1468 (O_1468,N_29003,N_29077);
nand UO_1469 (O_1469,N_28906,N_28878);
nor UO_1470 (O_1470,N_29828,N_29264);
or UO_1471 (O_1471,N_29261,N_29001);
nand UO_1472 (O_1472,N_29423,N_29107);
or UO_1473 (O_1473,N_28829,N_29203);
nand UO_1474 (O_1474,N_29007,N_29088);
and UO_1475 (O_1475,N_29073,N_29513);
or UO_1476 (O_1476,N_29168,N_28912);
nand UO_1477 (O_1477,N_29990,N_29223);
xor UO_1478 (O_1478,N_29211,N_29129);
nor UO_1479 (O_1479,N_29282,N_29302);
and UO_1480 (O_1480,N_29182,N_29088);
nand UO_1481 (O_1481,N_28812,N_29922);
nand UO_1482 (O_1482,N_29461,N_29032);
xor UO_1483 (O_1483,N_29850,N_29324);
xnor UO_1484 (O_1484,N_29999,N_29783);
xor UO_1485 (O_1485,N_29847,N_29422);
xnor UO_1486 (O_1486,N_29705,N_29645);
xor UO_1487 (O_1487,N_29664,N_28800);
xor UO_1488 (O_1488,N_29795,N_29809);
and UO_1489 (O_1489,N_29133,N_29209);
and UO_1490 (O_1490,N_28928,N_29352);
nor UO_1491 (O_1491,N_28947,N_28832);
and UO_1492 (O_1492,N_28900,N_28964);
xnor UO_1493 (O_1493,N_28815,N_29215);
and UO_1494 (O_1494,N_29866,N_28976);
or UO_1495 (O_1495,N_29723,N_28945);
and UO_1496 (O_1496,N_29426,N_29717);
nor UO_1497 (O_1497,N_29435,N_29795);
nor UO_1498 (O_1498,N_29970,N_29141);
nand UO_1499 (O_1499,N_29475,N_29590);
nor UO_1500 (O_1500,N_29523,N_29568);
nand UO_1501 (O_1501,N_28937,N_29777);
or UO_1502 (O_1502,N_29320,N_29244);
or UO_1503 (O_1503,N_28949,N_29097);
nor UO_1504 (O_1504,N_29369,N_29028);
nor UO_1505 (O_1505,N_29326,N_29763);
nor UO_1506 (O_1506,N_29910,N_29941);
or UO_1507 (O_1507,N_29760,N_28884);
nor UO_1508 (O_1508,N_29706,N_28856);
nand UO_1509 (O_1509,N_29587,N_28948);
and UO_1510 (O_1510,N_28966,N_29449);
nand UO_1511 (O_1511,N_29222,N_29793);
nor UO_1512 (O_1512,N_29259,N_28954);
nand UO_1513 (O_1513,N_29507,N_29127);
or UO_1514 (O_1514,N_29549,N_29979);
or UO_1515 (O_1515,N_29070,N_29706);
nor UO_1516 (O_1516,N_29639,N_29426);
or UO_1517 (O_1517,N_29286,N_29356);
or UO_1518 (O_1518,N_28803,N_29689);
xnor UO_1519 (O_1519,N_29739,N_29348);
nand UO_1520 (O_1520,N_29260,N_29081);
xnor UO_1521 (O_1521,N_29180,N_29291);
and UO_1522 (O_1522,N_29809,N_29974);
nand UO_1523 (O_1523,N_29370,N_29160);
nand UO_1524 (O_1524,N_29431,N_29892);
or UO_1525 (O_1525,N_29114,N_29887);
and UO_1526 (O_1526,N_29076,N_29700);
xnor UO_1527 (O_1527,N_28841,N_29094);
xor UO_1528 (O_1528,N_29760,N_29327);
nand UO_1529 (O_1529,N_29657,N_29804);
xor UO_1530 (O_1530,N_29191,N_29467);
nand UO_1531 (O_1531,N_29448,N_29797);
nand UO_1532 (O_1532,N_29374,N_29227);
nand UO_1533 (O_1533,N_29808,N_29569);
nand UO_1534 (O_1534,N_29703,N_29603);
and UO_1535 (O_1535,N_29686,N_29385);
and UO_1536 (O_1536,N_29732,N_29752);
or UO_1537 (O_1537,N_29255,N_29360);
and UO_1538 (O_1538,N_28916,N_29293);
and UO_1539 (O_1539,N_29927,N_29030);
and UO_1540 (O_1540,N_29227,N_29873);
nand UO_1541 (O_1541,N_29886,N_29625);
xnor UO_1542 (O_1542,N_29219,N_29186);
or UO_1543 (O_1543,N_29325,N_28927);
and UO_1544 (O_1544,N_29359,N_29622);
xor UO_1545 (O_1545,N_29883,N_29704);
xnor UO_1546 (O_1546,N_29924,N_29233);
nand UO_1547 (O_1547,N_29359,N_29245);
and UO_1548 (O_1548,N_29667,N_29750);
and UO_1549 (O_1549,N_29962,N_29727);
and UO_1550 (O_1550,N_29022,N_29944);
xnor UO_1551 (O_1551,N_29312,N_29132);
xnor UO_1552 (O_1552,N_29722,N_29606);
nor UO_1553 (O_1553,N_28924,N_29976);
and UO_1554 (O_1554,N_29711,N_29182);
xor UO_1555 (O_1555,N_29565,N_29606);
xor UO_1556 (O_1556,N_29190,N_29827);
nand UO_1557 (O_1557,N_29769,N_29813);
and UO_1558 (O_1558,N_29272,N_29819);
xor UO_1559 (O_1559,N_29878,N_29856);
or UO_1560 (O_1560,N_29723,N_29018);
or UO_1561 (O_1561,N_28956,N_29307);
nand UO_1562 (O_1562,N_29009,N_29651);
or UO_1563 (O_1563,N_29791,N_29106);
xnor UO_1564 (O_1564,N_29558,N_29611);
or UO_1565 (O_1565,N_29987,N_29896);
xor UO_1566 (O_1566,N_29151,N_29395);
nor UO_1567 (O_1567,N_29723,N_28946);
nand UO_1568 (O_1568,N_28863,N_29803);
nand UO_1569 (O_1569,N_28938,N_29998);
nand UO_1570 (O_1570,N_29253,N_29853);
or UO_1571 (O_1571,N_29604,N_29370);
nand UO_1572 (O_1572,N_28883,N_29919);
or UO_1573 (O_1573,N_29734,N_29591);
and UO_1574 (O_1574,N_29073,N_29999);
xnor UO_1575 (O_1575,N_29258,N_29004);
nor UO_1576 (O_1576,N_29209,N_28979);
and UO_1577 (O_1577,N_29374,N_29758);
xor UO_1578 (O_1578,N_29824,N_29808);
or UO_1579 (O_1579,N_29951,N_29137);
and UO_1580 (O_1580,N_29000,N_29651);
nand UO_1581 (O_1581,N_29543,N_29400);
nor UO_1582 (O_1582,N_29987,N_28837);
xnor UO_1583 (O_1583,N_29541,N_29990);
nor UO_1584 (O_1584,N_29158,N_28978);
nand UO_1585 (O_1585,N_28849,N_29724);
or UO_1586 (O_1586,N_29637,N_29046);
or UO_1587 (O_1587,N_29076,N_28810);
or UO_1588 (O_1588,N_29569,N_29247);
and UO_1589 (O_1589,N_29016,N_29835);
nand UO_1590 (O_1590,N_29628,N_29014);
nor UO_1591 (O_1591,N_29115,N_29517);
nand UO_1592 (O_1592,N_29733,N_29360);
nor UO_1593 (O_1593,N_29909,N_28972);
xor UO_1594 (O_1594,N_29335,N_29048);
and UO_1595 (O_1595,N_29463,N_29128);
or UO_1596 (O_1596,N_29780,N_29945);
xnor UO_1597 (O_1597,N_29414,N_29196);
xnor UO_1598 (O_1598,N_29222,N_29002);
or UO_1599 (O_1599,N_28956,N_29233);
or UO_1600 (O_1600,N_29304,N_29695);
or UO_1601 (O_1601,N_29655,N_28894);
nor UO_1602 (O_1602,N_29124,N_29628);
nand UO_1603 (O_1603,N_29499,N_28959);
xor UO_1604 (O_1604,N_29495,N_29623);
nand UO_1605 (O_1605,N_29816,N_29589);
or UO_1606 (O_1606,N_28933,N_28939);
xor UO_1607 (O_1607,N_29360,N_29032);
nor UO_1608 (O_1608,N_28957,N_29616);
xor UO_1609 (O_1609,N_29767,N_29850);
nand UO_1610 (O_1610,N_29155,N_29983);
and UO_1611 (O_1611,N_29334,N_29256);
xnor UO_1612 (O_1612,N_28965,N_29917);
or UO_1613 (O_1613,N_29676,N_28828);
nor UO_1614 (O_1614,N_29082,N_29663);
and UO_1615 (O_1615,N_29280,N_29346);
xnor UO_1616 (O_1616,N_29853,N_28953);
or UO_1617 (O_1617,N_28801,N_29530);
nand UO_1618 (O_1618,N_28838,N_29293);
or UO_1619 (O_1619,N_29379,N_29382);
nor UO_1620 (O_1620,N_29582,N_29424);
nor UO_1621 (O_1621,N_29290,N_29900);
nor UO_1622 (O_1622,N_29544,N_29222);
nand UO_1623 (O_1623,N_29215,N_29846);
nand UO_1624 (O_1624,N_29167,N_29852);
and UO_1625 (O_1625,N_29199,N_29712);
nand UO_1626 (O_1626,N_29527,N_29213);
xor UO_1627 (O_1627,N_29116,N_29823);
nand UO_1628 (O_1628,N_28922,N_29089);
xor UO_1629 (O_1629,N_29032,N_29363);
and UO_1630 (O_1630,N_29672,N_29787);
and UO_1631 (O_1631,N_29829,N_29362);
nor UO_1632 (O_1632,N_29214,N_29101);
nor UO_1633 (O_1633,N_29342,N_29780);
nor UO_1634 (O_1634,N_29343,N_29149);
xnor UO_1635 (O_1635,N_29125,N_29681);
nor UO_1636 (O_1636,N_29476,N_29343);
xnor UO_1637 (O_1637,N_28863,N_29979);
or UO_1638 (O_1638,N_29947,N_29675);
and UO_1639 (O_1639,N_29022,N_29680);
nor UO_1640 (O_1640,N_29121,N_28829);
xnor UO_1641 (O_1641,N_28949,N_29542);
nor UO_1642 (O_1642,N_29226,N_29065);
xor UO_1643 (O_1643,N_29513,N_29269);
nand UO_1644 (O_1644,N_29178,N_28947);
nor UO_1645 (O_1645,N_29994,N_29282);
nor UO_1646 (O_1646,N_29731,N_29284);
and UO_1647 (O_1647,N_29242,N_29875);
nor UO_1648 (O_1648,N_29732,N_29427);
xor UO_1649 (O_1649,N_29156,N_29402);
xor UO_1650 (O_1650,N_29072,N_29994);
nand UO_1651 (O_1651,N_29363,N_29742);
nand UO_1652 (O_1652,N_29862,N_29164);
or UO_1653 (O_1653,N_29257,N_29449);
and UO_1654 (O_1654,N_29741,N_29248);
nand UO_1655 (O_1655,N_29244,N_29377);
nor UO_1656 (O_1656,N_29699,N_29881);
nor UO_1657 (O_1657,N_29640,N_29665);
xor UO_1658 (O_1658,N_29572,N_29708);
or UO_1659 (O_1659,N_29540,N_29051);
nand UO_1660 (O_1660,N_29404,N_29022);
nor UO_1661 (O_1661,N_29974,N_29825);
nand UO_1662 (O_1662,N_29667,N_29610);
xnor UO_1663 (O_1663,N_28802,N_28963);
and UO_1664 (O_1664,N_29587,N_29255);
or UO_1665 (O_1665,N_29689,N_29642);
or UO_1666 (O_1666,N_29880,N_29616);
or UO_1667 (O_1667,N_29632,N_29882);
nor UO_1668 (O_1668,N_29348,N_29852);
xor UO_1669 (O_1669,N_29737,N_28945);
or UO_1670 (O_1670,N_29151,N_28919);
and UO_1671 (O_1671,N_28847,N_29326);
xnor UO_1672 (O_1672,N_29909,N_29527);
nand UO_1673 (O_1673,N_28852,N_29282);
xnor UO_1674 (O_1674,N_29724,N_29223);
nor UO_1675 (O_1675,N_29144,N_29198);
nand UO_1676 (O_1676,N_28833,N_29239);
nand UO_1677 (O_1677,N_29995,N_29085);
and UO_1678 (O_1678,N_29260,N_29319);
or UO_1679 (O_1679,N_29449,N_28894);
nand UO_1680 (O_1680,N_29859,N_29861);
and UO_1681 (O_1681,N_29433,N_29077);
nand UO_1682 (O_1682,N_29402,N_28932);
or UO_1683 (O_1683,N_28937,N_28987);
nand UO_1684 (O_1684,N_29313,N_29251);
and UO_1685 (O_1685,N_29104,N_29281);
or UO_1686 (O_1686,N_29389,N_28890);
and UO_1687 (O_1687,N_29072,N_28960);
and UO_1688 (O_1688,N_29626,N_29524);
and UO_1689 (O_1689,N_29346,N_29875);
xor UO_1690 (O_1690,N_29659,N_29663);
xnor UO_1691 (O_1691,N_29620,N_29706);
nand UO_1692 (O_1692,N_29806,N_29807);
or UO_1693 (O_1693,N_29165,N_28948);
nand UO_1694 (O_1694,N_29415,N_29359);
and UO_1695 (O_1695,N_29273,N_29516);
nor UO_1696 (O_1696,N_29523,N_29441);
or UO_1697 (O_1697,N_29565,N_29540);
nand UO_1698 (O_1698,N_28842,N_29984);
nor UO_1699 (O_1699,N_29895,N_29890);
and UO_1700 (O_1700,N_29159,N_29560);
and UO_1701 (O_1701,N_29651,N_29921);
nor UO_1702 (O_1702,N_29597,N_29939);
nand UO_1703 (O_1703,N_29989,N_29902);
or UO_1704 (O_1704,N_29136,N_28871);
and UO_1705 (O_1705,N_29868,N_29917);
and UO_1706 (O_1706,N_29004,N_29145);
and UO_1707 (O_1707,N_29144,N_28892);
nor UO_1708 (O_1708,N_28920,N_29716);
nor UO_1709 (O_1709,N_28852,N_28942);
nand UO_1710 (O_1710,N_29045,N_29318);
nor UO_1711 (O_1711,N_29855,N_29095);
and UO_1712 (O_1712,N_28841,N_29904);
nor UO_1713 (O_1713,N_29370,N_29195);
and UO_1714 (O_1714,N_28953,N_28848);
xnor UO_1715 (O_1715,N_29213,N_28849);
nor UO_1716 (O_1716,N_29342,N_29361);
and UO_1717 (O_1717,N_29268,N_28905);
nand UO_1718 (O_1718,N_29593,N_28833);
nand UO_1719 (O_1719,N_28838,N_29369);
xnor UO_1720 (O_1720,N_28893,N_29213);
and UO_1721 (O_1721,N_29733,N_28972);
nor UO_1722 (O_1722,N_29300,N_29241);
or UO_1723 (O_1723,N_29588,N_29896);
or UO_1724 (O_1724,N_29417,N_29344);
nor UO_1725 (O_1725,N_29723,N_29304);
xor UO_1726 (O_1726,N_29804,N_29232);
or UO_1727 (O_1727,N_29533,N_29358);
nand UO_1728 (O_1728,N_29478,N_28950);
or UO_1729 (O_1729,N_29581,N_29628);
xnor UO_1730 (O_1730,N_29199,N_29571);
and UO_1731 (O_1731,N_29018,N_29583);
and UO_1732 (O_1732,N_29159,N_29504);
and UO_1733 (O_1733,N_29052,N_29920);
or UO_1734 (O_1734,N_29021,N_29159);
xnor UO_1735 (O_1735,N_29568,N_28844);
nand UO_1736 (O_1736,N_29951,N_28959);
or UO_1737 (O_1737,N_29912,N_29204);
xnor UO_1738 (O_1738,N_29842,N_29553);
xnor UO_1739 (O_1739,N_29408,N_28894);
or UO_1740 (O_1740,N_29738,N_29233);
and UO_1741 (O_1741,N_29732,N_29895);
nand UO_1742 (O_1742,N_29613,N_29468);
xnor UO_1743 (O_1743,N_29688,N_29974);
or UO_1744 (O_1744,N_29222,N_29658);
xor UO_1745 (O_1745,N_28853,N_28866);
and UO_1746 (O_1746,N_29236,N_29251);
nand UO_1747 (O_1747,N_29559,N_29685);
and UO_1748 (O_1748,N_29844,N_29141);
xnor UO_1749 (O_1749,N_28999,N_29541);
or UO_1750 (O_1750,N_29624,N_29584);
xnor UO_1751 (O_1751,N_29334,N_29270);
nand UO_1752 (O_1752,N_29867,N_29205);
xor UO_1753 (O_1753,N_29913,N_29477);
and UO_1754 (O_1754,N_29441,N_29595);
or UO_1755 (O_1755,N_29156,N_29740);
nor UO_1756 (O_1756,N_29824,N_29502);
nor UO_1757 (O_1757,N_29580,N_29982);
xnor UO_1758 (O_1758,N_29936,N_29817);
or UO_1759 (O_1759,N_29807,N_28918);
or UO_1760 (O_1760,N_29114,N_29247);
or UO_1761 (O_1761,N_28976,N_29839);
and UO_1762 (O_1762,N_28862,N_29870);
nor UO_1763 (O_1763,N_29905,N_29664);
nor UO_1764 (O_1764,N_29605,N_29748);
and UO_1765 (O_1765,N_29690,N_29641);
and UO_1766 (O_1766,N_29204,N_29212);
nor UO_1767 (O_1767,N_29374,N_29663);
xnor UO_1768 (O_1768,N_28851,N_29988);
xor UO_1769 (O_1769,N_29732,N_28921);
nor UO_1770 (O_1770,N_29788,N_29890);
or UO_1771 (O_1771,N_29825,N_29677);
nor UO_1772 (O_1772,N_29619,N_29327);
xnor UO_1773 (O_1773,N_29504,N_29792);
and UO_1774 (O_1774,N_29196,N_29708);
nand UO_1775 (O_1775,N_28810,N_29041);
nand UO_1776 (O_1776,N_29652,N_28991);
and UO_1777 (O_1777,N_29246,N_29339);
nor UO_1778 (O_1778,N_29326,N_29688);
and UO_1779 (O_1779,N_29928,N_29106);
xor UO_1780 (O_1780,N_29991,N_29777);
nand UO_1781 (O_1781,N_29239,N_29648);
and UO_1782 (O_1782,N_29533,N_29334);
or UO_1783 (O_1783,N_29390,N_29520);
and UO_1784 (O_1784,N_29862,N_29276);
or UO_1785 (O_1785,N_29804,N_29670);
and UO_1786 (O_1786,N_29616,N_28868);
and UO_1787 (O_1787,N_28823,N_29644);
and UO_1788 (O_1788,N_29092,N_29601);
and UO_1789 (O_1789,N_29157,N_29918);
or UO_1790 (O_1790,N_29142,N_28882);
and UO_1791 (O_1791,N_29994,N_29294);
nand UO_1792 (O_1792,N_29541,N_29066);
and UO_1793 (O_1793,N_29196,N_29268);
or UO_1794 (O_1794,N_29932,N_29642);
xor UO_1795 (O_1795,N_29026,N_29917);
xnor UO_1796 (O_1796,N_29140,N_29339);
nand UO_1797 (O_1797,N_29302,N_29676);
and UO_1798 (O_1798,N_29759,N_29615);
nand UO_1799 (O_1799,N_29230,N_29302);
and UO_1800 (O_1800,N_28863,N_29778);
xor UO_1801 (O_1801,N_29256,N_29629);
nand UO_1802 (O_1802,N_29631,N_29958);
nor UO_1803 (O_1803,N_29615,N_28957);
nor UO_1804 (O_1804,N_29693,N_29574);
and UO_1805 (O_1805,N_29790,N_29119);
nor UO_1806 (O_1806,N_29599,N_29952);
and UO_1807 (O_1807,N_29937,N_29757);
xnor UO_1808 (O_1808,N_28862,N_29327);
nor UO_1809 (O_1809,N_29504,N_28851);
xor UO_1810 (O_1810,N_29862,N_29034);
or UO_1811 (O_1811,N_29103,N_28845);
nor UO_1812 (O_1812,N_29446,N_29917);
nand UO_1813 (O_1813,N_28834,N_29852);
or UO_1814 (O_1814,N_29142,N_29135);
or UO_1815 (O_1815,N_29750,N_29548);
nand UO_1816 (O_1816,N_28955,N_29682);
xnor UO_1817 (O_1817,N_28957,N_28870);
nor UO_1818 (O_1818,N_29996,N_29245);
or UO_1819 (O_1819,N_29467,N_29165);
or UO_1820 (O_1820,N_29512,N_28892);
nand UO_1821 (O_1821,N_28952,N_29273);
or UO_1822 (O_1822,N_29493,N_29624);
nand UO_1823 (O_1823,N_29694,N_29842);
nor UO_1824 (O_1824,N_29133,N_29932);
xor UO_1825 (O_1825,N_29972,N_29040);
or UO_1826 (O_1826,N_29600,N_29648);
and UO_1827 (O_1827,N_29707,N_29774);
nand UO_1828 (O_1828,N_29691,N_29137);
nor UO_1829 (O_1829,N_29189,N_28899);
nor UO_1830 (O_1830,N_29029,N_29192);
or UO_1831 (O_1831,N_28845,N_29020);
nand UO_1832 (O_1832,N_29172,N_29549);
or UO_1833 (O_1833,N_29810,N_28910);
nand UO_1834 (O_1834,N_28918,N_29197);
and UO_1835 (O_1835,N_29283,N_29202);
and UO_1836 (O_1836,N_29773,N_28981);
or UO_1837 (O_1837,N_29595,N_28956);
and UO_1838 (O_1838,N_29998,N_29088);
nand UO_1839 (O_1839,N_29039,N_29470);
nor UO_1840 (O_1840,N_29607,N_28881);
nor UO_1841 (O_1841,N_29155,N_29449);
nor UO_1842 (O_1842,N_29369,N_29006);
and UO_1843 (O_1843,N_29926,N_28813);
nor UO_1844 (O_1844,N_29975,N_29033);
and UO_1845 (O_1845,N_29909,N_29145);
and UO_1846 (O_1846,N_29982,N_29008);
and UO_1847 (O_1847,N_28945,N_29255);
nand UO_1848 (O_1848,N_29556,N_28978);
nor UO_1849 (O_1849,N_29334,N_29074);
nand UO_1850 (O_1850,N_29011,N_29535);
nand UO_1851 (O_1851,N_28952,N_29105);
nand UO_1852 (O_1852,N_29160,N_29383);
or UO_1853 (O_1853,N_29595,N_29816);
nand UO_1854 (O_1854,N_29947,N_29330);
nand UO_1855 (O_1855,N_29545,N_29057);
and UO_1856 (O_1856,N_29957,N_29034);
and UO_1857 (O_1857,N_29635,N_29811);
and UO_1858 (O_1858,N_29430,N_29202);
and UO_1859 (O_1859,N_29848,N_29657);
nand UO_1860 (O_1860,N_29927,N_29851);
and UO_1861 (O_1861,N_29773,N_29398);
nor UO_1862 (O_1862,N_29973,N_29563);
xor UO_1863 (O_1863,N_28905,N_29229);
and UO_1864 (O_1864,N_28849,N_29182);
xnor UO_1865 (O_1865,N_29173,N_29168);
or UO_1866 (O_1866,N_29939,N_29535);
xnor UO_1867 (O_1867,N_29481,N_29013);
and UO_1868 (O_1868,N_29788,N_29821);
or UO_1869 (O_1869,N_28945,N_29658);
nand UO_1870 (O_1870,N_29056,N_29800);
and UO_1871 (O_1871,N_29132,N_29243);
and UO_1872 (O_1872,N_29907,N_29291);
nand UO_1873 (O_1873,N_29215,N_28988);
or UO_1874 (O_1874,N_29839,N_29389);
xnor UO_1875 (O_1875,N_28829,N_29826);
xor UO_1876 (O_1876,N_29207,N_29050);
and UO_1877 (O_1877,N_29072,N_29151);
nor UO_1878 (O_1878,N_29370,N_29929);
nand UO_1879 (O_1879,N_29804,N_29664);
and UO_1880 (O_1880,N_29030,N_28863);
nand UO_1881 (O_1881,N_29116,N_29508);
nor UO_1882 (O_1882,N_28815,N_29025);
nand UO_1883 (O_1883,N_29034,N_29502);
nand UO_1884 (O_1884,N_29558,N_29826);
and UO_1885 (O_1885,N_29504,N_29723);
and UO_1886 (O_1886,N_29940,N_29345);
nand UO_1887 (O_1887,N_29179,N_29973);
or UO_1888 (O_1888,N_29858,N_28818);
and UO_1889 (O_1889,N_29810,N_29795);
xor UO_1890 (O_1890,N_29844,N_29962);
xor UO_1891 (O_1891,N_29429,N_29413);
nand UO_1892 (O_1892,N_28886,N_29887);
nor UO_1893 (O_1893,N_29427,N_29406);
nor UO_1894 (O_1894,N_28905,N_29405);
nor UO_1895 (O_1895,N_29616,N_28976);
and UO_1896 (O_1896,N_28908,N_29733);
or UO_1897 (O_1897,N_28887,N_29243);
nor UO_1898 (O_1898,N_29365,N_29221);
nor UO_1899 (O_1899,N_28897,N_29413);
nand UO_1900 (O_1900,N_29333,N_29316);
nor UO_1901 (O_1901,N_29592,N_29920);
xnor UO_1902 (O_1902,N_29547,N_29887);
xnor UO_1903 (O_1903,N_29261,N_29829);
xor UO_1904 (O_1904,N_29890,N_29892);
xor UO_1905 (O_1905,N_28995,N_28949);
and UO_1906 (O_1906,N_29519,N_29546);
nand UO_1907 (O_1907,N_29994,N_29186);
xor UO_1908 (O_1908,N_29521,N_29555);
nor UO_1909 (O_1909,N_29231,N_29427);
xnor UO_1910 (O_1910,N_29393,N_29070);
nor UO_1911 (O_1911,N_29031,N_29046);
or UO_1912 (O_1912,N_28882,N_28982);
or UO_1913 (O_1913,N_28938,N_29297);
or UO_1914 (O_1914,N_29124,N_28865);
nand UO_1915 (O_1915,N_29944,N_29179);
xor UO_1916 (O_1916,N_29627,N_29267);
nand UO_1917 (O_1917,N_29069,N_29731);
xor UO_1918 (O_1918,N_29078,N_29018);
or UO_1919 (O_1919,N_28903,N_29081);
nor UO_1920 (O_1920,N_29616,N_29356);
and UO_1921 (O_1921,N_29213,N_29888);
and UO_1922 (O_1922,N_28839,N_29987);
nand UO_1923 (O_1923,N_29436,N_29291);
nand UO_1924 (O_1924,N_29762,N_28900);
and UO_1925 (O_1925,N_29849,N_29385);
or UO_1926 (O_1926,N_28819,N_29327);
or UO_1927 (O_1927,N_28837,N_29083);
and UO_1928 (O_1928,N_29726,N_29245);
xor UO_1929 (O_1929,N_29500,N_29374);
and UO_1930 (O_1930,N_29544,N_29080);
xnor UO_1931 (O_1931,N_29155,N_29838);
or UO_1932 (O_1932,N_28862,N_29812);
and UO_1933 (O_1933,N_29895,N_29090);
xor UO_1934 (O_1934,N_29808,N_29053);
nor UO_1935 (O_1935,N_29550,N_29380);
and UO_1936 (O_1936,N_29555,N_29640);
or UO_1937 (O_1937,N_29862,N_29957);
nand UO_1938 (O_1938,N_29782,N_29951);
and UO_1939 (O_1939,N_28919,N_29655);
and UO_1940 (O_1940,N_29998,N_28929);
xor UO_1941 (O_1941,N_29090,N_28947);
nor UO_1942 (O_1942,N_29563,N_29511);
or UO_1943 (O_1943,N_29905,N_29278);
nand UO_1944 (O_1944,N_29486,N_28949);
nor UO_1945 (O_1945,N_29650,N_29691);
nor UO_1946 (O_1946,N_29769,N_29744);
nand UO_1947 (O_1947,N_29046,N_28846);
and UO_1948 (O_1948,N_29959,N_29645);
nand UO_1949 (O_1949,N_28848,N_29570);
nand UO_1950 (O_1950,N_29683,N_28931);
nand UO_1951 (O_1951,N_28814,N_29681);
xor UO_1952 (O_1952,N_29926,N_29961);
or UO_1953 (O_1953,N_28941,N_28976);
nor UO_1954 (O_1954,N_29711,N_29608);
nor UO_1955 (O_1955,N_29632,N_29706);
or UO_1956 (O_1956,N_29207,N_29710);
or UO_1957 (O_1957,N_29357,N_29510);
nand UO_1958 (O_1958,N_29513,N_29207);
nor UO_1959 (O_1959,N_29556,N_29633);
and UO_1960 (O_1960,N_29950,N_29265);
nor UO_1961 (O_1961,N_29557,N_29217);
or UO_1962 (O_1962,N_29974,N_29465);
nor UO_1963 (O_1963,N_29501,N_28982);
xor UO_1964 (O_1964,N_29827,N_29315);
nand UO_1965 (O_1965,N_29861,N_29549);
nand UO_1966 (O_1966,N_29335,N_29588);
and UO_1967 (O_1967,N_28827,N_29367);
xor UO_1968 (O_1968,N_29040,N_29341);
nand UO_1969 (O_1969,N_29201,N_29995);
and UO_1970 (O_1970,N_29573,N_29516);
nand UO_1971 (O_1971,N_29529,N_29509);
and UO_1972 (O_1972,N_29155,N_29974);
and UO_1973 (O_1973,N_29050,N_29134);
nor UO_1974 (O_1974,N_29041,N_29663);
and UO_1975 (O_1975,N_29205,N_28846);
or UO_1976 (O_1976,N_28819,N_29439);
nor UO_1977 (O_1977,N_29170,N_29676);
nor UO_1978 (O_1978,N_29284,N_29992);
xnor UO_1979 (O_1979,N_29841,N_29265);
xor UO_1980 (O_1980,N_29202,N_29835);
nand UO_1981 (O_1981,N_29738,N_29188);
nor UO_1982 (O_1982,N_29761,N_29210);
and UO_1983 (O_1983,N_29880,N_29358);
and UO_1984 (O_1984,N_29968,N_28905);
and UO_1985 (O_1985,N_28906,N_29845);
and UO_1986 (O_1986,N_29982,N_29441);
nand UO_1987 (O_1987,N_29839,N_29071);
or UO_1988 (O_1988,N_29756,N_29283);
xnor UO_1989 (O_1989,N_28922,N_29245);
nand UO_1990 (O_1990,N_29800,N_29700);
nor UO_1991 (O_1991,N_29156,N_29561);
xnor UO_1992 (O_1992,N_29357,N_29368);
xnor UO_1993 (O_1993,N_28968,N_29429);
or UO_1994 (O_1994,N_29325,N_29673);
nor UO_1995 (O_1995,N_29904,N_29745);
nand UO_1996 (O_1996,N_29095,N_29523);
and UO_1997 (O_1997,N_29469,N_28892);
nor UO_1998 (O_1998,N_29517,N_29508);
xnor UO_1999 (O_1999,N_29959,N_29791);
or UO_2000 (O_2000,N_29138,N_29169);
or UO_2001 (O_2001,N_28842,N_29102);
xor UO_2002 (O_2002,N_29180,N_29001);
nand UO_2003 (O_2003,N_29278,N_29043);
xor UO_2004 (O_2004,N_29928,N_29446);
xor UO_2005 (O_2005,N_29794,N_29326);
nor UO_2006 (O_2006,N_29907,N_29374);
nand UO_2007 (O_2007,N_29566,N_28947);
and UO_2008 (O_2008,N_28919,N_29790);
xnor UO_2009 (O_2009,N_29690,N_29803);
nor UO_2010 (O_2010,N_29820,N_29706);
nor UO_2011 (O_2011,N_29954,N_29835);
xnor UO_2012 (O_2012,N_28863,N_29219);
xnor UO_2013 (O_2013,N_29464,N_28815);
and UO_2014 (O_2014,N_29942,N_28918);
nor UO_2015 (O_2015,N_29012,N_29778);
nand UO_2016 (O_2016,N_29440,N_28857);
nand UO_2017 (O_2017,N_29231,N_29132);
nand UO_2018 (O_2018,N_29636,N_28830);
xor UO_2019 (O_2019,N_29346,N_28948);
or UO_2020 (O_2020,N_28945,N_28862);
nor UO_2021 (O_2021,N_29397,N_29383);
xnor UO_2022 (O_2022,N_29226,N_29905);
or UO_2023 (O_2023,N_29148,N_29806);
xor UO_2024 (O_2024,N_28998,N_28974);
and UO_2025 (O_2025,N_29683,N_28966);
or UO_2026 (O_2026,N_29853,N_29295);
and UO_2027 (O_2027,N_29776,N_29493);
xor UO_2028 (O_2028,N_29612,N_29697);
nand UO_2029 (O_2029,N_29513,N_29652);
xor UO_2030 (O_2030,N_29481,N_29105);
or UO_2031 (O_2031,N_29071,N_28824);
nand UO_2032 (O_2032,N_28911,N_29440);
xor UO_2033 (O_2033,N_28839,N_29313);
nor UO_2034 (O_2034,N_29892,N_29947);
nor UO_2035 (O_2035,N_29625,N_29001);
nand UO_2036 (O_2036,N_29789,N_28892);
or UO_2037 (O_2037,N_29859,N_28853);
and UO_2038 (O_2038,N_29810,N_29007);
and UO_2039 (O_2039,N_29834,N_29458);
nor UO_2040 (O_2040,N_29581,N_29553);
and UO_2041 (O_2041,N_28868,N_29511);
nor UO_2042 (O_2042,N_29587,N_29715);
xor UO_2043 (O_2043,N_29047,N_29832);
nor UO_2044 (O_2044,N_28998,N_29125);
or UO_2045 (O_2045,N_29354,N_29587);
nand UO_2046 (O_2046,N_29150,N_29042);
nand UO_2047 (O_2047,N_29892,N_29591);
nand UO_2048 (O_2048,N_29217,N_29756);
xor UO_2049 (O_2049,N_29400,N_29046);
nor UO_2050 (O_2050,N_29911,N_28859);
nand UO_2051 (O_2051,N_28996,N_29259);
nor UO_2052 (O_2052,N_29459,N_29079);
or UO_2053 (O_2053,N_29401,N_28814);
or UO_2054 (O_2054,N_29107,N_29854);
nand UO_2055 (O_2055,N_28973,N_29798);
xnor UO_2056 (O_2056,N_29471,N_28958);
or UO_2057 (O_2057,N_29462,N_28809);
or UO_2058 (O_2058,N_29651,N_29515);
nor UO_2059 (O_2059,N_29229,N_29130);
nand UO_2060 (O_2060,N_29214,N_29482);
nor UO_2061 (O_2061,N_29749,N_29214);
nand UO_2062 (O_2062,N_29972,N_28846);
nand UO_2063 (O_2063,N_29727,N_29320);
or UO_2064 (O_2064,N_29747,N_29339);
or UO_2065 (O_2065,N_29044,N_29281);
nand UO_2066 (O_2066,N_29727,N_29487);
nand UO_2067 (O_2067,N_28984,N_29938);
and UO_2068 (O_2068,N_29778,N_29319);
nand UO_2069 (O_2069,N_28986,N_29944);
or UO_2070 (O_2070,N_29358,N_29082);
nor UO_2071 (O_2071,N_29303,N_29335);
nand UO_2072 (O_2072,N_29899,N_29575);
and UO_2073 (O_2073,N_29568,N_29327);
nor UO_2074 (O_2074,N_29933,N_29673);
nand UO_2075 (O_2075,N_29545,N_29086);
and UO_2076 (O_2076,N_29673,N_29430);
nor UO_2077 (O_2077,N_28887,N_29858);
and UO_2078 (O_2078,N_29836,N_29127);
and UO_2079 (O_2079,N_29753,N_29248);
xor UO_2080 (O_2080,N_29480,N_29584);
xor UO_2081 (O_2081,N_29461,N_29105);
nor UO_2082 (O_2082,N_29057,N_29043);
or UO_2083 (O_2083,N_29456,N_29526);
or UO_2084 (O_2084,N_29062,N_29205);
nand UO_2085 (O_2085,N_29699,N_29341);
xnor UO_2086 (O_2086,N_29452,N_29057);
or UO_2087 (O_2087,N_29585,N_28844);
nor UO_2088 (O_2088,N_28875,N_29608);
nand UO_2089 (O_2089,N_29157,N_29757);
xnor UO_2090 (O_2090,N_28843,N_29737);
xor UO_2091 (O_2091,N_29449,N_29705);
or UO_2092 (O_2092,N_29146,N_28914);
and UO_2093 (O_2093,N_29250,N_29550);
and UO_2094 (O_2094,N_29227,N_29986);
or UO_2095 (O_2095,N_29190,N_29891);
nor UO_2096 (O_2096,N_29603,N_29188);
xor UO_2097 (O_2097,N_29035,N_28849);
nand UO_2098 (O_2098,N_29747,N_29336);
or UO_2099 (O_2099,N_29120,N_29882);
or UO_2100 (O_2100,N_29233,N_29757);
nor UO_2101 (O_2101,N_29210,N_29297);
nor UO_2102 (O_2102,N_29012,N_29420);
and UO_2103 (O_2103,N_29499,N_28864);
nand UO_2104 (O_2104,N_29154,N_29699);
xnor UO_2105 (O_2105,N_29619,N_28820);
nand UO_2106 (O_2106,N_28915,N_29484);
nand UO_2107 (O_2107,N_29213,N_29913);
nor UO_2108 (O_2108,N_29818,N_29036);
nand UO_2109 (O_2109,N_29428,N_29235);
or UO_2110 (O_2110,N_29968,N_29522);
and UO_2111 (O_2111,N_29601,N_28909);
nand UO_2112 (O_2112,N_29810,N_29046);
and UO_2113 (O_2113,N_29401,N_29094);
or UO_2114 (O_2114,N_29914,N_29277);
or UO_2115 (O_2115,N_29123,N_29508);
and UO_2116 (O_2116,N_29673,N_28821);
and UO_2117 (O_2117,N_29311,N_29814);
xnor UO_2118 (O_2118,N_29767,N_29091);
or UO_2119 (O_2119,N_29928,N_29516);
xor UO_2120 (O_2120,N_29645,N_29953);
and UO_2121 (O_2121,N_29179,N_29776);
nor UO_2122 (O_2122,N_29553,N_29172);
xnor UO_2123 (O_2123,N_29696,N_29954);
xor UO_2124 (O_2124,N_29216,N_28927);
xnor UO_2125 (O_2125,N_29563,N_29614);
or UO_2126 (O_2126,N_29600,N_29221);
or UO_2127 (O_2127,N_29282,N_29970);
or UO_2128 (O_2128,N_28966,N_29807);
nand UO_2129 (O_2129,N_29671,N_29939);
nand UO_2130 (O_2130,N_29875,N_29088);
and UO_2131 (O_2131,N_29033,N_28960);
nor UO_2132 (O_2132,N_29761,N_28948);
nor UO_2133 (O_2133,N_29521,N_29939);
or UO_2134 (O_2134,N_29090,N_29521);
or UO_2135 (O_2135,N_29358,N_29447);
or UO_2136 (O_2136,N_29675,N_29313);
or UO_2137 (O_2137,N_29960,N_29153);
nand UO_2138 (O_2138,N_28987,N_28928);
nand UO_2139 (O_2139,N_29312,N_28806);
and UO_2140 (O_2140,N_28847,N_29489);
xnor UO_2141 (O_2141,N_29102,N_29859);
or UO_2142 (O_2142,N_29650,N_29720);
or UO_2143 (O_2143,N_29604,N_29794);
and UO_2144 (O_2144,N_29299,N_29328);
and UO_2145 (O_2145,N_29526,N_29011);
or UO_2146 (O_2146,N_29650,N_28835);
or UO_2147 (O_2147,N_29468,N_29178);
nand UO_2148 (O_2148,N_29094,N_28855);
nor UO_2149 (O_2149,N_28919,N_29894);
xor UO_2150 (O_2150,N_29467,N_29833);
or UO_2151 (O_2151,N_29871,N_29620);
and UO_2152 (O_2152,N_29006,N_29928);
and UO_2153 (O_2153,N_29819,N_29323);
nor UO_2154 (O_2154,N_29825,N_29439);
and UO_2155 (O_2155,N_29496,N_29130);
or UO_2156 (O_2156,N_29337,N_29099);
nor UO_2157 (O_2157,N_29473,N_29845);
and UO_2158 (O_2158,N_29131,N_29146);
nand UO_2159 (O_2159,N_28937,N_29120);
and UO_2160 (O_2160,N_29300,N_28835);
nand UO_2161 (O_2161,N_29413,N_29674);
xnor UO_2162 (O_2162,N_29390,N_29822);
or UO_2163 (O_2163,N_28878,N_29258);
and UO_2164 (O_2164,N_28822,N_29701);
nor UO_2165 (O_2165,N_29456,N_29377);
xnor UO_2166 (O_2166,N_29116,N_29628);
or UO_2167 (O_2167,N_28862,N_29731);
or UO_2168 (O_2168,N_29908,N_29094);
nand UO_2169 (O_2169,N_29487,N_29729);
nor UO_2170 (O_2170,N_29060,N_29953);
nor UO_2171 (O_2171,N_29185,N_29359);
xnor UO_2172 (O_2172,N_29669,N_29990);
xor UO_2173 (O_2173,N_29613,N_29197);
or UO_2174 (O_2174,N_29467,N_29041);
nor UO_2175 (O_2175,N_29550,N_29194);
xor UO_2176 (O_2176,N_29097,N_29240);
and UO_2177 (O_2177,N_29690,N_29256);
and UO_2178 (O_2178,N_29968,N_29687);
xor UO_2179 (O_2179,N_29204,N_29973);
and UO_2180 (O_2180,N_29542,N_28975);
nand UO_2181 (O_2181,N_29383,N_29651);
nor UO_2182 (O_2182,N_29552,N_29246);
nor UO_2183 (O_2183,N_29999,N_29239);
xor UO_2184 (O_2184,N_29726,N_29585);
and UO_2185 (O_2185,N_28981,N_29977);
xnor UO_2186 (O_2186,N_29577,N_28915);
nand UO_2187 (O_2187,N_29473,N_28913);
nand UO_2188 (O_2188,N_29559,N_29310);
xnor UO_2189 (O_2189,N_29264,N_29299);
or UO_2190 (O_2190,N_28961,N_29412);
or UO_2191 (O_2191,N_29675,N_29057);
or UO_2192 (O_2192,N_29156,N_29019);
and UO_2193 (O_2193,N_29753,N_29760);
nand UO_2194 (O_2194,N_29527,N_28874);
nand UO_2195 (O_2195,N_29015,N_29435);
and UO_2196 (O_2196,N_28938,N_29391);
or UO_2197 (O_2197,N_29146,N_29020);
xor UO_2198 (O_2198,N_29867,N_29905);
and UO_2199 (O_2199,N_29994,N_29540);
or UO_2200 (O_2200,N_29321,N_29540);
xor UO_2201 (O_2201,N_28836,N_29622);
nor UO_2202 (O_2202,N_29235,N_29270);
xor UO_2203 (O_2203,N_29149,N_29184);
nor UO_2204 (O_2204,N_29371,N_29597);
and UO_2205 (O_2205,N_29356,N_29023);
and UO_2206 (O_2206,N_29419,N_28883);
nand UO_2207 (O_2207,N_29034,N_29307);
nand UO_2208 (O_2208,N_29042,N_29694);
xor UO_2209 (O_2209,N_29058,N_29287);
or UO_2210 (O_2210,N_29923,N_29560);
and UO_2211 (O_2211,N_29803,N_28811);
or UO_2212 (O_2212,N_29878,N_29376);
nor UO_2213 (O_2213,N_29017,N_29782);
xnor UO_2214 (O_2214,N_29631,N_29475);
nand UO_2215 (O_2215,N_28955,N_29466);
or UO_2216 (O_2216,N_29502,N_28978);
and UO_2217 (O_2217,N_29151,N_29769);
xor UO_2218 (O_2218,N_29049,N_29427);
and UO_2219 (O_2219,N_29183,N_29992);
xor UO_2220 (O_2220,N_29528,N_28872);
nand UO_2221 (O_2221,N_29615,N_29122);
and UO_2222 (O_2222,N_29461,N_29372);
nand UO_2223 (O_2223,N_29214,N_29127);
xnor UO_2224 (O_2224,N_29389,N_29640);
xnor UO_2225 (O_2225,N_29150,N_28987);
and UO_2226 (O_2226,N_28967,N_29623);
or UO_2227 (O_2227,N_29506,N_29641);
nand UO_2228 (O_2228,N_28923,N_29128);
nor UO_2229 (O_2229,N_29977,N_29852);
xor UO_2230 (O_2230,N_29926,N_29832);
xor UO_2231 (O_2231,N_29780,N_29379);
nor UO_2232 (O_2232,N_29198,N_29811);
and UO_2233 (O_2233,N_29713,N_29526);
and UO_2234 (O_2234,N_29026,N_28923);
nor UO_2235 (O_2235,N_29195,N_29620);
and UO_2236 (O_2236,N_29117,N_29800);
xor UO_2237 (O_2237,N_29169,N_29848);
xnor UO_2238 (O_2238,N_29590,N_29278);
nand UO_2239 (O_2239,N_28806,N_29796);
and UO_2240 (O_2240,N_29632,N_28896);
or UO_2241 (O_2241,N_29915,N_28970);
nor UO_2242 (O_2242,N_28931,N_29324);
nor UO_2243 (O_2243,N_29334,N_29993);
and UO_2244 (O_2244,N_29215,N_29534);
or UO_2245 (O_2245,N_29656,N_29814);
or UO_2246 (O_2246,N_28939,N_29402);
nor UO_2247 (O_2247,N_28930,N_29168);
nor UO_2248 (O_2248,N_29710,N_29863);
xor UO_2249 (O_2249,N_29849,N_28900);
or UO_2250 (O_2250,N_29312,N_29412);
or UO_2251 (O_2251,N_29185,N_29880);
or UO_2252 (O_2252,N_29546,N_29424);
nand UO_2253 (O_2253,N_29895,N_29342);
or UO_2254 (O_2254,N_29459,N_29957);
xor UO_2255 (O_2255,N_28978,N_29675);
nand UO_2256 (O_2256,N_28955,N_28833);
and UO_2257 (O_2257,N_29970,N_29915);
or UO_2258 (O_2258,N_29044,N_28943);
xnor UO_2259 (O_2259,N_29997,N_29953);
nor UO_2260 (O_2260,N_29018,N_29303);
xor UO_2261 (O_2261,N_29536,N_29485);
xor UO_2262 (O_2262,N_28968,N_29437);
nand UO_2263 (O_2263,N_28809,N_29518);
xnor UO_2264 (O_2264,N_29964,N_29149);
nand UO_2265 (O_2265,N_29759,N_29213);
nand UO_2266 (O_2266,N_29359,N_29811);
or UO_2267 (O_2267,N_29188,N_28877);
xnor UO_2268 (O_2268,N_29145,N_29073);
or UO_2269 (O_2269,N_28825,N_29690);
nand UO_2270 (O_2270,N_29757,N_29942);
xor UO_2271 (O_2271,N_29705,N_29992);
nand UO_2272 (O_2272,N_29425,N_29680);
xnor UO_2273 (O_2273,N_29055,N_29348);
xor UO_2274 (O_2274,N_29068,N_29477);
nor UO_2275 (O_2275,N_29067,N_29648);
nand UO_2276 (O_2276,N_28819,N_29275);
nand UO_2277 (O_2277,N_29792,N_29364);
xnor UO_2278 (O_2278,N_29688,N_29537);
and UO_2279 (O_2279,N_28964,N_29716);
nor UO_2280 (O_2280,N_29809,N_29821);
or UO_2281 (O_2281,N_29173,N_28900);
and UO_2282 (O_2282,N_29260,N_28808);
or UO_2283 (O_2283,N_29108,N_29234);
nor UO_2284 (O_2284,N_29271,N_29860);
nor UO_2285 (O_2285,N_29496,N_29342);
xor UO_2286 (O_2286,N_29124,N_29845);
xor UO_2287 (O_2287,N_29716,N_29003);
nand UO_2288 (O_2288,N_29532,N_29051);
nor UO_2289 (O_2289,N_29400,N_29077);
nand UO_2290 (O_2290,N_29024,N_28940);
nand UO_2291 (O_2291,N_29189,N_29403);
or UO_2292 (O_2292,N_29753,N_29588);
or UO_2293 (O_2293,N_29850,N_29735);
xnor UO_2294 (O_2294,N_29842,N_29104);
xnor UO_2295 (O_2295,N_29507,N_29451);
xnor UO_2296 (O_2296,N_29196,N_29887);
and UO_2297 (O_2297,N_29690,N_29443);
or UO_2298 (O_2298,N_28883,N_29847);
nand UO_2299 (O_2299,N_28973,N_29359);
or UO_2300 (O_2300,N_29196,N_28854);
and UO_2301 (O_2301,N_29403,N_29889);
or UO_2302 (O_2302,N_29692,N_29235);
nand UO_2303 (O_2303,N_29129,N_28803);
xor UO_2304 (O_2304,N_29871,N_29789);
nor UO_2305 (O_2305,N_28843,N_29298);
xnor UO_2306 (O_2306,N_29903,N_29940);
and UO_2307 (O_2307,N_29829,N_29055);
or UO_2308 (O_2308,N_29794,N_29552);
and UO_2309 (O_2309,N_28808,N_29569);
nor UO_2310 (O_2310,N_29152,N_29131);
and UO_2311 (O_2311,N_29714,N_29572);
and UO_2312 (O_2312,N_29679,N_28960);
nand UO_2313 (O_2313,N_29883,N_29098);
nor UO_2314 (O_2314,N_28930,N_29785);
and UO_2315 (O_2315,N_29988,N_28941);
nand UO_2316 (O_2316,N_29741,N_29504);
xor UO_2317 (O_2317,N_29654,N_29936);
or UO_2318 (O_2318,N_29634,N_29171);
nor UO_2319 (O_2319,N_29132,N_29404);
nor UO_2320 (O_2320,N_29053,N_29628);
and UO_2321 (O_2321,N_29537,N_29436);
xor UO_2322 (O_2322,N_29564,N_29409);
xor UO_2323 (O_2323,N_29128,N_29287);
nor UO_2324 (O_2324,N_29657,N_29247);
or UO_2325 (O_2325,N_29579,N_29031);
nand UO_2326 (O_2326,N_29455,N_29400);
nor UO_2327 (O_2327,N_29649,N_29331);
nor UO_2328 (O_2328,N_29568,N_29907);
nor UO_2329 (O_2329,N_29078,N_29639);
nand UO_2330 (O_2330,N_29871,N_29244);
or UO_2331 (O_2331,N_29748,N_29969);
or UO_2332 (O_2332,N_29679,N_29320);
or UO_2333 (O_2333,N_29736,N_28944);
or UO_2334 (O_2334,N_29141,N_29002);
and UO_2335 (O_2335,N_29807,N_29621);
and UO_2336 (O_2336,N_29864,N_29026);
xor UO_2337 (O_2337,N_29119,N_29698);
nor UO_2338 (O_2338,N_29300,N_29025);
or UO_2339 (O_2339,N_29960,N_29930);
xor UO_2340 (O_2340,N_29230,N_29882);
or UO_2341 (O_2341,N_29079,N_28954);
or UO_2342 (O_2342,N_29919,N_29173);
nand UO_2343 (O_2343,N_29266,N_29819);
and UO_2344 (O_2344,N_28994,N_28968);
or UO_2345 (O_2345,N_29349,N_28803);
or UO_2346 (O_2346,N_29940,N_29151);
xnor UO_2347 (O_2347,N_29157,N_29972);
nor UO_2348 (O_2348,N_29996,N_29266);
xnor UO_2349 (O_2349,N_28946,N_29380);
nor UO_2350 (O_2350,N_28917,N_29026);
nand UO_2351 (O_2351,N_29975,N_29639);
nor UO_2352 (O_2352,N_28899,N_29100);
xor UO_2353 (O_2353,N_29248,N_28822);
nor UO_2354 (O_2354,N_29580,N_29649);
or UO_2355 (O_2355,N_28906,N_29846);
xor UO_2356 (O_2356,N_29271,N_29357);
nand UO_2357 (O_2357,N_29872,N_28843);
or UO_2358 (O_2358,N_29203,N_29361);
nor UO_2359 (O_2359,N_29403,N_28849);
nand UO_2360 (O_2360,N_29833,N_29882);
and UO_2361 (O_2361,N_29591,N_29317);
or UO_2362 (O_2362,N_29456,N_29028);
nor UO_2363 (O_2363,N_29217,N_28887);
and UO_2364 (O_2364,N_29427,N_28834);
nand UO_2365 (O_2365,N_28901,N_29022);
or UO_2366 (O_2366,N_29668,N_29188);
nand UO_2367 (O_2367,N_29014,N_29799);
nand UO_2368 (O_2368,N_29343,N_29137);
xnor UO_2369 (O_2369,N_29081,N_29039);
xnor UO_2370 (O_2370,N_29411,N_28894);
xor UO_2371 (O_2371,N_29926,N_29788);
and UO_2372 (O_2372,N_29312,N_28884);
nand UO_2373 (O_2373,N_29366,N_29677);
nor UO_2374 (O_2374,N_29131,N_28807);
or UO_2375 (O_2375,N_29292,N_29103);
nand UO_2376 (O_2376,N_29252,N_29154);
and UO_2377 (O_2377,N_28801,N_29528);
nand UO_2378 (O_2378,N_29881,N_29678);
nor UO_2379 (O_2379,N_29070,N_29896);
and UO_2380 (O_2380,N_29784,N_29211);
nor UO_2381 (O_2381,N_29892,N_29597);
xor UO_2382 (O_2382,N_29133,N_29066);
nand UO_2383 (O_2383,N_29833,N_29924);
or UO_2384 (O_2384,N_29098,N_29894);
nand UO_2385 (O_2385,N_29942,N_29951);
nor UO_2386 (O_2386,N_29825,N_29268);
xnor UO_2387 (O_2387,N_29622,N_29723);
or UO_2388 (O_2388,N_28871,N_29397);
and UO_2389 (O_2389,N_29197,N_29478);
nand UO_2390 (O_2390,N_29827,N_29747);
nand UO_2391 (O_2391,N_29552,N_28891);
xor UO_2392 (O_2392,N_29576,N_28870);
xnor UO_2393 (O_2393,N_29441,N_29659);
xor UO_2394 (O_2394,N_29297,N_29412);
and UO_2395 (O_2395,N_29799,N_29234);
nor UO_2396 (O_2396,N_29581,N_29224);
nand UO_2397 (O_2397,N_29948,N_28809);
xnor UO_2398 (O_2398,N_29884,N_29744);
nor UO_2399 (O_2399,N_29130,N_29002);
xor UO_2400 (O_2400,N_29379,N_29926);
nor UO_2401 (O_2401,N_29126,N_29604);
xor UO_2402 (O_2402,N_29673,N_28930);
xor UO_2403 (O_2403,N_29630,N_29465);
or UO_2404 (O_2404,N_29116,N_29134);
and UO_2405 (O_2405,N_29303,N_29059);
xor UO_2406 (O_2406,N_29283,N_29400);
and UO_2407 (O_2407,N_28940,N_29955);
nand UO_2408 (O_2408,N_29766,N_28979);
nand UO_2409 (O_2409,N_29851,N_29923);
nand UO_2410 (O_2410,N_29860,N_29260);
xnor UO_2411 (O_2411,N_29856,N_29389);
xnor UO_2412 (O_2412,N_28939,N_29180);
xnor UO_2413 (O_2413,N_29744,N_29345);
xor UO_2414 (O_2414,N_29341,N_28851);
xnor UO_2415 (O_2415,N_29643,N_29682);
xnor UO_2416 (O_2416,N_29177,N_29131);
nor UO_2417 (O_2417,N_28987,N_29650);
and UO_2418 (O_2418,N_29954,N_29199);
or UO_2419 (O_2419,N_28955,N_29977);
xnor UO_2420 (O_2420,N_29454,N_29706);
nand UO_2421 (O_2421,N_29295,N_29818);
or UO_2422 (O_2422,N_29696,N_29935);
nor UO_2423 (O_2423,N_29581,N_29572);
or UO_2424 (O_2424,N_29385,N_28915);
nand UO_2425 (O_2425,N_29202,N_28968);
and UO_2426 (O_2426,N_29845,N_29431);
and UO_2427 (O_2427,N_29356,N_29975);
and UO_2428 (O_2428,N_29013,N_29344);
and UO_2429 (O_2429,N_29673,N_29180);
and UO_2430 (O_2430,N_29048,N_29995);
xnor UO_2431 (O_2431,N_28845,N_29090);
nand UO_2432 (O_2432,N_28919,N_29861);
or UO_2433 (O_2433,N_29966,N_29850);
nand UO_2434 (O_2434,N_29938,N_29637);
or UO_2435 (O_2435,N_29894,N_28917);
xnor UO_2436 (O_2436,N_29484,N_29668);
or UO_2437 (O_2437,N_29503,N_29354);
or UO_2438 (O_2438,N_29724,N_28946);
and UO_2439 (O_2439,N_29847,N_29320);
nor UO_2440 (O_2440,N_29184,N_29157);
and UO_2441 (O_2441,N_29438,N_28894);
and UO_2442 (O_2442,N_29733,N_29959);
and UO_2443 (O_2443,N_29638,N_29179);
xor UO_2444 (O_2444,N_28911,N_29743);
nor UO_2445 (O_2445,N_28854,N_29166);
xnor UO_2446 (O_2446,N_29733,N_29583);
or UO_2447 (O_2447,N_29540,N_29747);
or UO_2448 (O_2448,N_29344,N_29522);
nor UO_2449 (O_2449,N_29698,N_29783);
xor UO_2450 (O_2450,N_29347,N_29899);
and UO_2451 (O_2451,N_29261,N_29510);
xor UO_2452 (O_2452,N_29963,N_28817);
and UO_2453 (O_2453,N_29467,N_29232);
nand UO_2454 (O_2454,N_29771,N_29699);
and UO_2455 (O_2455,N_29032,N_28872);
or UO_2456 (O_2456,N_29876,N_29799);
xnor UO_2457 (O_2457,N_29207,N_28815);
or UO_2458 (O_2458,N_28967,N_28910);
xor UO_2459 (O_2459,N_28949,N_29107);
nand UO_2460 (O_2460,N_28857,N_29672);
and UO_2461 (O_2461,N_28851,N_28961);
or UO_2462 (O_2462,N_29542,N_29800);
nor UO_2463 (O_2463,N_28953,N_29475);
or UO_2464 (O_2464,N_29359,N_29279);
nand UO_2465 (O_2465,N_28808,N_28817);
nand UO_2466 (O_2466,N_29451,N_29963);
and UO_2467 (O_2467,N_29591,N_29420);
nand UO_2468 (O_2468,N_29385,N_29891);
nor UO_2469 (O_2469,N_29360,N_29642);
nor UO_2470 (O_2470,N_29743,N_29806);
and UO_2471 (O_2471,N_29772,N_28907);
xor UO_2472 (O_2472,N_29971,N_29535);
and UO_2473 (O_2473,N_29747,N_29638);
xor UO_2474 (O_2474,N_29301,N_29506);
and UO_2475 (O_2475,N_29032,N_29143);
or UO_2476 (O_2476,N_29899,N_29845);
nand UO_2477 (O_2477,N_29508,N_29879);
and UO_2478 (O_2478,N_29704,N_29419);
nor UO_2479 (O_2479,N_28920,N_29715);
nand UO_2480 (O_2480,N_29178,N_29304);
and UO_2481 (O_2481,N_29978,N_29283);
nand UO_2482 (O_2482,N_29920,N_29319);
and UO_2483 (O_2483,N_28826,N_29656);
and UO_2484 (O_2484,N_29290,N_29712);
or UO_2485 (O_2485,N_29583,N_29382);
nor UO_2486 (O_2486,N_29571,N_29681);
or UO_2487 (O_2487,N_28855,N_29385);
xnor UO_2488 (O_2488,N_29099,N_29477);
xnor UO_2489 (O_2489,N_29515,N_29738);
xor UO_2490 (O_2490,N_29555,N_29289);
xnor UO_2491 (O_2491,N_29792,N_29376);
and UO_2492 (O_2492,N_29444,N_29658);
xnor UO_2493 (O_2493,N_29294,N_29709);
nor UO_2494 (O_2494,N_29582,N_29196);
or UO_2495 (O_2495,N_29670,N_29878);
nand UO_2496 (O_2496,N_29848,N_29770);
nor UO_2497 (O_2497,N_29289,N_28818);
nor UO_2498 (O_2498,N_29989,N_29954);
nand UO_2499 (O_2499,N_29633,N_29505);
nand UO_2500 (O_2500,N_29469,N_28920);
xor UO_2501 (O_2501,N_29325,N_29428);
and UO_2502 (O_2502,N_29289,N_28858);
nor UO_2503 (O_2503,N_29995,N_28922);
and UO_2504 (O_2504,N_29805,N_29337);
nor UO_2505 (O_2505,N_29601,N_29174);
or UO_2506 (O_2506,N_29842,N_29636);
or UO_2507 (O_2507,N_29791,N_28940);
nand UO_2508 (O_2508,N_28954,N_29561);
or UO_2509 (O_2509,N_29497,N_29523);
nand UO_2510 (O_2510,N_29641,N_29812);
xnor UO_2511 (O_2511,N_28972,N_29107);
xnor UO_2512 (O_2512,N_29519,N_29285);
and UO_2513 (O_2513,N_29425,N_29704);
nor UO_2514 (O_2514,N_28872,N_29718);
or UO_2515 (O_2515,N_29387,N_29405);
nand UO_2516 (O_2516,N_28927,N_28969);
nand UO_2517 (O_2517,N_29654,N_28872);
and UO_2518 (O_2518,N_29795,N_29932);
and UO_2519 (O_2519,N_28811,N_29424);
and UO_2520 (O_2520,N_29180,N_29498);
and UO_2521 (O_2521,N_28880,N_29179);
or UO_2522 (O_2522,N_29893,N_28854);
nand UO_2523 (O_2523,N_29883,N_28852);
xnor UO_2524 (O_2524,N_29884,N_29041);
nor UO_2525 (O_2525,N_28834,N_29791);
or UO_2526 (O_2526,N_28943,N_29290);
xor UO_2527 (O_2527,N_29090,N_28889);
or UO_2528 (O_2528,N_29180,N_29500);
xnor UO_2529 (O_2529,N_29667,N_28916);
nand UO_2530 (O_2530,N_29630,N_28987);
xor UO_2531 (O_2531,N_29765,N_29193);
or UO_2532 (O_2532,N_29240,N_29456);
or UO_2533 (O_2533,N_29248,N_29778);
or UO_2534 (O_2534,N_29099,N_29154);
xor UO_2535 (O_2535,N_29289,N_28957);
or UO_2536 (O_2536,N_29561,N_28925);
nand UO_2537 (O_2537,N_29063,N_29353);
and UO_2538 (O_2538,N_29785,N_29040);
xor UO_2539 (O_2539,N_29290,N_29057);
and UO_2540 (O_2540,N_28954,N_29421);
and UO_2541 (O_2541,N_29481,N_29795);
nand UO_2542 (O_2542,N_29334,N_29988);
nand UO_2543 (O_2543,N_29803,N_29503);
and UO_2544 (O_2544,N_28942,N_28944);
xnor UO_2545 (O_2545,N_29611,N_29966);
or UO_2546 (O_2546,N_29267,N_28987);
and UO_2547 (O_2547,N_28901,N_28998);
xnor UO_2548 (O_2548,N_29258,N_29663);
and UO_2549 (O_2549,N_29084,N_28811);
and UO_2550 (O_2550,N_29098,N_29468);
and UO_2551 (O_2551,N_29795,N_29431);
and UO_2552 (O_2552,N_29157,N_29638);
nand UO_2553 (O_2553,N_29796,N_29325);
nor UO_2554 (O_2554,N_29067,N_29721);
xnor UO_2555 (O_2555,N_29106,N_29318);
or UO_2556 (O_2556,N_29063,N_29174);
nand UO_2557 (O_2557,N_29092,N_29132);
nor UO_2558 (O_2558,N_29464,N_29130);
nand UO_2559 (O_2559,N_29937,N_29380);
or UO_2560 (O_2560,N_28928,N_29582);
or UO_2561 (O_2561,N_29834,N_29606);
or UO_2562 (O_2562,N_29759,N_29851);
or UO_2563 (O_2563,N_29868,N_28948);
nand UO_2564 (O_2564,N_29775,N_29803);
nor UO_2565 (O_2565,N_29925,N_29526);
nor UO_2566 (O_2566,N_29157,N_29450);
or UO_2567 (O_2567,N_29175,N_29816);
xnor UO_2568 (O_2568,N_29519,N_29653);
nor UO_2569 (O_2569,N_29126,N_29349);
or UO_2570 (O_2570,N_29886,N_28961);
nand UO_2571 (O_2571,N_29813,N_29333);
or UO_2572 (O_2572,N_29914,N_29652);
nand UO_2573 (O_2573,N_29810,N_29993);
or UO_2574 (O_2574,N_29612,N_29406);
xor UO_2575 (O_2575,N_29796,N_29165);
xor UO_2576 (O_2576,N_29599,N_29361);
nand UO_2577 (O_2577,N_29101,N_29357);
or UO_2578 (O_2578,N_29547,N_29777);
xnor UO_2579 (O_2579,N_28839,N_29112);
nand UO_2580 (O_2580,N_28993,N_28879);
or UO_2581 (O_2581,N_28891,N_29789);
or UO_2582 (O_2582,N_29114,N_29110);
or UO_2583 (O_2583,N_29253,N_29772);
xnor UO_2584 (O_2584,N_28964,N_29200);
nand UO_2585 (O_2585,N_29365,N_28878);
nand UO_2586 (O_2586,N_29144,N_29028);
or UO_2587 (O_2587,N_29758,N_29120);
or UO_2588 (O_2588,N_29122,N_29843);
and UO_2589 (O_2589,N_29084,N_29022);
nor UO_2590 (O_2590,N_29133,N_29324);
nor UO_2591 (O_2591,N_29054,N_29929);
nand UO_2592 (O_2592,N_29766,N_28826);
or UO_2593 (O_2593,N_29909,N_28867);
xor UO_2594 (O_2594,N_29993,N_28952);
and UO_2595 (O_2595,N_29341,N_29614);
nand UO_2596 (O_2596,N_29918,N_29607);
nor UO_2597 (O_2597,N_29926,N_29678);
and UO_2598 (O_2598,N_29803,N_29275);
or UO_2599 (O_2599,N_29556,N_29511);
xor UO_2600 (O_2600,N_29233,N_28970);
nor UO_2601 (O_2601,N_28876,N_29105);
xnor UO_2602 (O_2602,N_28975,N_29242);
xor UO_2603 (O_2603,N_29534,N_29900);
and UO_2604 (O_2604,N_29443,N_29273);
and UO_2605 (O_2605,N_29368,N_29156);
or UO_2606 (O_2606,N_29405,N_29247);
nor UO_2607 (O_2607,N_29514,N_29771);
xor UO_2608 (O_2608,N_29414,N_29058);
or UO_2609 (O_2609,N_29412,N_29363);
or UO_2610 (O_2610,N_29788,N_29744);
nor UO_2611 (O_2611,N_29843,N_28819);
nand UO_2612 (O_2612,N_28914,N_28881);
and UO_2613 (O_2613,N_28995,N_29355);
nor UO_2614 (O_2614,N_29672,N_29135);
or UO_2615 (O_2615,N_29196,N_29264);
or UO_2616 (O_2616,N_28807,N_29664);
nand UO_2617 (O_2617,N_29368,N_29715);
nand UO_2618 (O_2618,N_29272,N_29468);
nand UO_2619 (O_2619,N_28808,N_29453);
or UO_2620 (O_2620,N_29707,N_29038);
nand UO_2621 (O_2621,N_29053,N_29781);
nand UO_2622 (O_2622,N_29690,N_29226);
nand UO_2623 (O_2623,N_29959,N_28902);
xor UO_2624 (O_2624,N_29920,N_29704);
and UO_2625 (O_2625,N_28983,N_28908);
or UO_2626 (O_2626,N_29253,N_29203);
xor UO_2627 (O_2627,N_29409,N_28882);
nor UO_2628 (O_2628,N_29894,N_29062);
and UO_2629 (O_2629,N_28827,N_29187);
nand UO_2630 (O_2630,N_29838,N_29259);
nor UO_2631 (O_2631,N_29230,N_29054);
nand UO_2632 (O_2632,N_29632,N_29588);
nand UO_2633 (O_2633,N_29335,N_29866);
nor UO_2634 (O_2634,N_29204,N_29558);
and UO_2635 (O_2635,N_29197,N_29670);
xnor UO_2636 (O_2636,N_29182,N_29981);
and UO_2637 (O_2637,N_29507,N_29455);
nand UO_2638 (O_2638,N_29947,N_29341);
nand UO_2639 (O_2639,N_29817,N_29925);
xnor UO_2640 (O_2640,N_29824,N_29788);
xnor UO_2641 (O_2641,N_29996,N_29707);
nor UO_2642 (O_2642,N_29850,N_29536);
or UO_2643 (O_2643,N_29976,N_29717);
xnor UO_2644 (O_2644,N_29129,N_29324);
xnor UO_2645 (O_2645,N_29323,N_29294);
and UO_2646 (O_2646,N_29657,N_28950);
or UO_2647 (O_2647,N_29092,N_28950);
nor UO_2648 (O_2648,N_29285,N_29069);
and UO_2649 (O_2649,N_29681,N_29988);
nor UO_2650 (O_2650,N_29767,N_29505);
and UO_2651 (O_2651,N_29298,N_29443);
or UO_2652 (O_2652,N_29413,N_29896);
nand UO_2653 (O_2653,N_29620,N_29841);
and UO_2654 (O_2654,N_29303,N_28854);
xnor UO_2655 (O_2655,N_29941,N_29863);
nand UO_2656 (O_2656,N_29122,N_29846);
nor UO_2657 (O_2657,N_28906,N_29012);
nor UO_2658 (O_2658,N_29270,N_29020);
nand UO_2659 (O_2659,N_29702,N_29936);
or UO_2660 (O_2660,N_29568,N_29388);
xnor UO_2661 (O_2661,N_29788,N_29695);
or UO_2662 (O_2662,N_29663,N_29520);
or UO_2663 (O_2663,N_29641,N_28937);
xnor UO_2664 (O_2664,N_29154,N_29155);
nor UO_2665 (O_2665,N_29546,N_28998);
or UO_2666 (O_2666,N_29359,N_29302);
or UO_2667 (O_2667,N_29298,N_29827);
and UO_2668 (O_2668,N_29171,N_29638);
nand UO_2669 (O_2669,N_29714,N_29366);
and UO_2670 (O_2670,N_29345,N_29444);
and UO_2671 (O_2671,N_28942,N_29501);
nor UO_2672 (O_2672,N_29773,N_29381);
nor UO_2673 (O_2673,N_29746,N_29438);
or UO_2674 (O_2674,N_28945,N_29715);
or UO_2675 (O_2675,N_29052,N_28987);
xor UO_2676 (O_2676,N_29821,N_29279);
or UO_2677 (O_2677,N_29073,N_29912);
nor UO_2678 (O_2678,N_29803,N_29215);
or UO_2679 (O_2679,N_29562,N_29632);
and UO_2680 (O_2680,N_29268,N_29123);
nand UO_2681 (O_2681,N_29669,N_29664);
nand UO_2682 (O_2682,N_29382,N_29812);
or UO_2683 (O_2683,N_29544,N_29155);
or UO_2684 (O_2684,N_29988,N_29307);
or UO_2685 (O_2685,N_29852,N_29319);
or UO_2686 (O_2686,N_29326,N_29509);
xor UO_2687 (O_2687,N_29669,N_29866);
nand UO_2688 (O_2688,N_29083,N_29444);
and UO_2689 (O_2689,N_28858,N_28980);
nand UO_2690 (O_2690,N_28968,N_29506);
nand UO_2691 (O_2691,N_29363,N_28916);
nor UO_2692 (O_2692,N_29568,N_29928);
xnor UO_2693 (O_2693,N_28899,N_29353);
nand UO_2694 (O_2694,N_29414,N_29782);
or UO_2695 (O_2695,N_29264,N_29674);
xnor UO_2696 (O_2696,N_29880,N_29135);
nand UO_2697 (O_2697,N_29799,N_29724);
and UO_2698 (O_2698,N_28827,N_29660);
or UO_2699 (O_2699,N_29297,N_29715);
nor UO_2700 (O_2700,N_29025,N_29376);
nor UO_2701 (O_2701,N_29524,N_29575);
nand UO_2702 (O_2702,N_29297,N_29429);
or UO_2703 (O_2703,N_29879,N_29399);
nand UO_2704 (O_2704,N_29123,N_29282);
nand UO_2705 (O_2705,N_29761,N_29642);
xor UO_2706 (O_2706,N_29102,N_28928);
xnor UO_2707 (O_2707,N_29325,N_29459);
and UO_2708 (O_2708,N_29288,N_29479);
or UO_2709 (O_2709,N_29075,N_29908);
nor UO_2710 (O_2710,N_29937,N_29377);
nand UO_2711 (O_2711,N_29523,N_29572);
or UO_2712 (O_2712,N_29839,N_29832);
xnor UO_2713 (O_2713,N_29385,N_29041);
and UO_2714 (O_2714,N_29182,N_29593);
nand UO_2715 (O_2715,N_29248,N_29089);
xor UO_2716 (O_2716,N_28927,N_29067);
nor UO_2717 (O_2717,N_29848,N_29988);
nor UO_2718 (O_2718,N_29065,N_29772);
nor UO_2719 (O_2719,N_28883,N_29638);
or UO_2720 (O_2720,N_29263,N_29104);
xnor UO_2721 (O_2721,N_28921,N_29919);
and UO_2722 (O_2722,N_29260,N_29818);
xor UO_2723 (O_2723,N_28828,N_29580);
or UO_2724 (O_2724,N_28963,N_29719);
nor UO_2725 (O_2725,N_29890,N_29247);
nor UO_2726 (O_2726,N_29174,N_29333);
nand UO_2727 (O_2727,N_29856,N_29514);
and UO_2728 (O_2728,N_29358,N_29184);
or UO_2729 (O_2729,N_29319,N_29027);
nor UO_2730 (O_2730,N_29287,N_29863);
or UO_2731 (O_2731,N_29830,N_29008);
nand UO_2732 (O_2732,N_29015,N_29561);
xnor UO_2733 (O_2733,N_29021,N_29435);
xor UO_2734 (O_2734,N_29653,N_28992);
nand UO_2735 (O_2735,N_28884,N_29012);
xnor UO_2736 (O_2736,N_29324,N_29436);
nand UO_2737 (O_2737,N_29493,N_29898);
or UO_2738 (O_2738,N_29030,N_29948);
xnor UO_2739 (O_2739,N_29203,N_29038);
nand UO_2740 (O_2740,N_28974,N_29547);
nand UO_2741 (O_2741,N_29825,N_29969);
and UO_2742 (O_2742,N_29873,N_29332);
xnor UO_2743 (O_2743,N_29347,N_29069);
nor UO_2744 (O_2744,N_29435,N_29445);
xor UO_2745 (O_2745,N_29326,N_29638);
xor UO_2746 (O_2746,N_29571,N_29950);
nand UO_2747 (O_2747,N_29952,N_29363);
and UO_2748 (O_2748,N_28835,N_29125);
nand UO_2749 (O_2749,N_29240,N_29604);
and UO_2750 (O_2750,N_29309,N_29292);
nand UO_2751 (O_2751,N_29332,N_29191);
or UO_2752 (O_2752,N_29538,N_29228);
nor UO_2753 (O_2753,N_29633,N_29880);
nor UO_2754 (O_2754,N_29223,N_29936);
and UO_2755 (O_2755,N_29100,N_29350);
nor UO_2756 (O_2756,N_29417,N_29946);
or UO_2757 (O_2757,N_29463,N_29931);
and UO_2758 (O_2758,N_29238,N_28816);
nor UO_2759 (O_2759,N_29689,N_29166);
xor UO_2760 (O_2760,N_29913,N_29041);
and UO_2761 (O_2761,N_29595,N_29514);
xnor UO_2762 (O_2762,N_29010,N_29096);
nor UO_2763 (O_2763,N_29940,N_29642);
and UO_2764 (O_2764,N_29430,N_29406);
nor UO_2765 (O_2765,N_28953,N_29729);
xor UO_2766 (O_2766,N_29217,N_29977);
xor UO_2767 (O_2767,N_29257,N_29896);
or UO_2768 (O_2768,N_29793,N_28812);
nand UO_2769 (O_2769,N_29168,N_29060);
or UO_2770 (O_2770,N_29892,N_29546);
or UO_2771 (O_2771,N_29554,N_29057);
xor UO_2772 (O_2772,N_29871,N_29684);
and UO_2773 (O_2773,N_29509,N_29524);
nor UO_2774 (O_2774,N_28842,N_29939);
or UO_2775 (O_2775,N_29089,N_29670);
xnor UO_2776 (O_2776,N_28908,N_28889);
nor UO_2777 (O_2777,N_29863,N_28839);
nor UO_2778 (O_2778,N_29855,N_28946);
nand UO_2779 (O_2779,N_29901,N_29396);
and UO_2780 (O_2780,N_29108,N_29904);
or UO_2781 (O_2781,N_29616,N_29437);
xnor UO_2782 (O_2782,N_29943,N_29945);
or UO_2783 (O_2783,N_28812,N_29431);
or UO_2784 (O_2784,N_29140,N_28816);
or UO_2785 (O_2785,N_29962,N_29015);
nor UO_2786 (O_2786,N_29151,N_29498);
xnor UO_2787 (O_2787,N_29328,N_29436);
or UO_2788 (O_2788,N_29130,N_29223);
or UO_2789 (O_2789,N_29123,N_29629);
nor UO_2790 (O_2790,N_29634,N_29595);
nand UO_2791 (O_2791,N_29629,N_28844);
and UO_2792 (O_2792,N_28968,N_29483);
xor UO_2793 (O_2793,N_29496,N_29040);
and UO_2794 (O_2794,N_29563,N_29487);
and UO_2795 (O_2795,N_29273,N_29682);
or UO_2796 (O_2796,N_29838,N_29192);
nor UO_2797 (O_2797,N_29370,N_29497);
nand UO_2798 (O_2798,N_29791,N_29580);
nor UO_2799 (O_2799,N_29835,N_29308);
nand UO_2800 (O_2800,N_29939,N_28974);
nor UO_2801 (O_2801,N_29984,N_29182);
nor UO_2802 (O_2802,N_29612,N_29302);
or UO_2803 (O_2803,N_29235,N_29494);
nor UO_2804 (O_2804,N_29212,N_29013);
and UO_2805 (O_2805,N_29787,N_29059);
or UO_2806 (O_2806,N_28800,N_29083);
and UO_2807 (O_2807,N_28833,N_29806);
nand UO_2808 (O_2808,N_29010,N_29387);
xnor UO_2809 (O_2809,N_28895,N_28958);
nor UO_2810 (O_2810,N_29875,N_29450);
nor UO_2811 (O_2811,N_29122,N_29744);
xnor UO_2812 (O_2812,N_29802,N_29735);
nor UO_2813 (O_2813,N_29708,N_28896);
nor UO_2814 (O_2814,N_29646,N_29176);
xor UO_2815 (O_2815,N_29653,N_28984);
nor UO_2816 (O_2816,N_28857,N_28870);
or UO_2817 (O_2817,N_28916,N_29541);
nand UO_2818 (O_2818,N_28860,N_29441);
or UO_2819 (O_2819,N_28932,N_29610);
and UO_2820 (O_2820,N_29304,N_28814);
and UO_2821 (O_2821,N_29470,N_29817);
nor UO_2822 (O_2822,N_29191,N_29051);
nand UO_2823 (O_2823,N_29626,N_29080);
nand UO_2824 (O_2824,N_28844,N_29227);
xnor UO_2825 (O_2825,N_29632,N_29122);
nor UO_2826 (O_2826,N_29673,N_29834);
or UO_2827 (O_2827,N_28867,N_28919);
nand UO_2828 (O_2828,N_29983,N_29394);
xor UO_2829 (O_2829,N_29267,N_29520);
nor UO_2830 (O_2830,N_29095,N_28879);
nand UO_2831 (O_2831,N_29640,N_29914);
or UO_2832 (O_2832,N_29679,N_29053);
xor UO_2833 (O_2833,N_29106,N_29848);
xor UO_2834 (O_2834,N_29394,N_29006);
nor UO_2835 (O_2835,N_28959,N_29014);
xnor UO_2836 (O_2836,N_29363,N_28986);
nor UO_2837 (O_2837,N_29606,N_28853);
and UO_2838 (O_2838,N_29590,N_29051);
xor UO_2839 (O_2839,N_29912,N_29392);
and UO_2840 (O_2840,N_29688,N_29081);
nand UO_2841 (O_2841,N_29722,N_29895);
and UO_2842 (O_2842,N_29295,N_29123);
and UO_2843 (O_2843,N_29565,N_29327);
nand UO_2844 (O_2844,N_29044,N_28828);
xor UO_2845 (O_2845,N_29139,N_29699);
xor UO_2846 (O_2846,N_29228,N_29199);
xor UO_2847 (O_2847,N_29231,N_29442);
nand UO_2848 (O_2848,N_29867,N_29246);
nand UO_2849 (O_2849,N_29943,N_29153);
nand UO_2850 (O_2850,N_29145,N_28957);
and UO_2851 (O_2851,N_29550,N_29985);
nor UO_2852 (O_2852,N_29577,N_29848);
xor UO_2853 (O_2853,N_29161,N_29237);
nor UO_2854 (O_2854,N_29231,N_28904);
nand UO_2855 (O_2855,N_29662,N_29139);
and UO_2856 (O_2856,N_29503,N_29035);
xor UO_2857 (O_2857,N_29230,N_29102);
and UO_2858 (O_2858,N_29692,N_29251);
xor UO_2859 (O_2859,N_29531,N_29655);
or UO_2860 (O_2860,N_29366,N_29711);
nand UO_2861 (O_2861,N_29134,N_29350);
and UO_2862 (O_2862,N_29204,N_29710);
and UO_2863 (O_2863,N_28870,N_29500);
or UO_2864 (O_2864,N_28855,N_29877);
nand UO_2865 (O_2865,N_29029,N_29451);
and UO_2866 (O_2866,N_29476,N_28811);
nor UO_2867 (O_2867,N_29935,N_29511);
nor UO_2868 (O_2868,N_29150,N_29624);
or UO_2869 (O_2869,N_28864,N_29597);
and UO_2870 (O_2870,N_29110,N_29320);
nand UO_2871 (O_2871,N_29010,N_29208);
or UO_2872 (O_2872,N_29828,N_29904);
nand UO_2873 (O_2873,N_29850,N_29316);
xnor UO_2874 (O_2874,N_29062,N_28802);
and UO_2875 (O_2875,N_29924,N_29126);
xor UO_2876 (O_2876,N_29722,N_29788);
nand UO_2877 (O_2877,N_29870,N_29157);
or UO_2878 (O_2878,N_29626,N_29625);
nand UO_2879 (O_2879,N_29458,N_29141);
nand UO_2880 (O_2880,N_29983,N_28836);
nand UO_2881 (O_2881,N_28826,N_28995);
xor UO_2882 (O_2882,N_29199,N_29129);
nand UO_2883 (O_2883,N_29138,N_29903);
nand UO_2884 (O_2884,N_29318,N_29641);
nor UO_2885 (O_2885,N_29209,N_28999);
nor UO_2886 (O_2886,N_29426,N_29852);
nor UO_2887 (O_2887,N_28845,N_29534);
nor UO_2888 (O_2888,N_29958,N_29009);
and UO_2889 (O_2889,N_28954,N_28872);
nor UO_2890 (O_2890,N_29756,N_29267);
xor UO_2891 (O_2891,N_29424,N_29287);
and UO_2892 (O_2892,N_29677,N_29331);
and UO_2893 (O_2893,N_29805,N_29474);
nor UO_2894 (O_2894,N_29666,N_29569);
xnor UO_2895 (O_2895,N_29271,N_29280);
nor UO_2896 (O_2896,N_29820,N_29995);
xnor UO_2897 (O_2897,N_29554,N_29636);
and UO_2898 (O_2898,N_28870,N_29717);
nand UO_2899 (O_2899,N_29233,N_28898);
nor UO_2900 (O_2900,N_28933,N_29772);
or UO_2901 (O_2901,N_29859,N_29642);
and UO_2902 (O_2902,N_29703,N_29954);
nand UO_2903 (O_2903,N_29014,N_28847);
or UO_2904 (O_2904,N_29642,N_29561);
nor UO_2905 (O_2905,N_29996,N_29960);
xnor UO_2906 (O_2906,N_28856,N_29270);
and UO_2907 (O_2907,N_29056,N_29116);
or UO_2908 (O_2908,N_29196,N_29199);
nand UO_2909 (O_2909,N_29472,N_29544);
nand UO_2910 (O_2910,N_28961,N_29262);
and UO_2911 (O_2911,N_29039,N_29790);
nand UO_2912 (O_2912,N_29681,N_28951);
xnor UO_2913 (O_2913,N_29557,N_29100);
or UO_2914 (O_2914,N_29641,N_29427);
xor UO_2915 (O_2915,N_29099,N_29718);
nor UO_2916 (O_2916,N_29655,N_29516);
and UO_2917 (O_2917,N_29224,N_29000);
and UO_2918 (O_2918,N_29814,N_29339);
nor UO_2919 (O_2919,N_29131,N_29487);
or UO_2920 (O_2920,N_29183,N_29206);
or UO_2921 (O_2921,N_29314,N_29488);
or UO_2922 (O_2922,N_29205,N_28866);
xor UO_2923 (O_2923,N_29247,N_28853);
and UO_2924 (O_2924,N_29695,N_29927);
or UO_2925 (O_2925,N_28952,N_29527);
xnor UO_2926 (O_2926,N_29919,N_29801);
xor UO_2927 (O_2927,N_29207,N_29958);
and UO_2928 (O_2928,N_29690,N_29336);
xnor UO_2929 (O_2929,N_29873,N_29534);
or UO_2930 (O_2930,N_29145,N_29592);
xnor UO_2931 (O_2931,N_28860,N_29728);
xor UO_2932 (O_2932,N_29721,N_29077);
and UO_2933 (O_2933,N_28949,N_29441);
nor UO_2934 (O_2934,N_29293,N_29471);
nand UO_2935 (O_2935,N_29527,N_29603);
nor UO_2936 (O_2936,N_29516,N_28820);
or UO_2937 (O_2937,N_29036,N_29675);
or UO_2938 (O_2938,N_29949,N_29591);
nand UO_2939 (O_2939,N_29557,N_29364);
or UO_2940 (O_2940,N_29656,N_28928);
and UO_2941 (O_2941,N_29314,N_29943);
nor UO_2942 (O_2942,N_29848,N_29138);
and UO_2943 (O_2943,N_29649,N_28891);
nor UO_2944 (O_2944,N_29397,N_28982);
or UO_2945 (O_2945,N_29734,N_29628);
and UO_2946 (O_2946,N_28985,N_29592);
nor UO_2947 (O_2947,N_28873,N_29165);
and UO_2948 (O_2948,N_29386,N_29776);
or UO_2949 (O_2949,N_29084,N_28830);
or UO_2950 (O_2950,N_29525,N_29107);
and UO_2951 (O_2951,N_29026,N_29180);
nand UO_2952 (O_2952,N_29477,N_29328);
xnor UO_2953 (O_2953,N_29178,N_29078);
and UO_2954 (O_2954,N_28926,N_29453);
or UO_2955 (O_2955,N_29556,N_29080);
nand UO_2956 (O_2956,N_29646,N_28888);
and UO_2957 (O_2957,N_29568,N_29070);
nor UO_2958 (O_2958,N_29548,N_28990);
nand UO_2959 (O_2959,N_29296,N_29789);
nor UO_2960 (O_2960,N_29002,N_29317);
xnor UO_2961 (O_2961,N_29202,N_28884);
xnor UO_2962 (O_2962,N_29806,N_29398);
xor UO_2963 (O_2963,N_29492,N_29888);
or UO_2964 (O_2964,N_29751,N_29967);
nand UO_2965 (O_2965,N_29306,N_29472);
nand UO_2966 (O_2966,N_29082,N_28849);
nor UO_2967 (O_2967,N_29763,N_29848);
nand UO_2968 (O_2968,N_29350,N_28975);
or UO_2969 (O_2969,N_29779,N_28891);
and UO_2970 (O_2970,N_29002,N_29549);
xor UO_2971 (O_2971,N_28969,N_29282);
xnor UO_2972 (O_2972,N_29312,N_29532);
and UO_2973 (O_2973,N_29499,N_29049);
or UO_2974 (O_2974,N_28811,N_29768);
xnor UO_2975 (O_2975,N_29930,N_29583);
nor UO_2976 (O_2976,N_29170,N_28852);
and UO_2977 (O_2977,N_29988,N_29168);
or UO_2978 (O_2978,N_29419,N_29946);
xor UO_2979 (O_2979,N_28922,N_29941);
or UO_2980 (O_2980,N_29149,N_29237);
and UO_2981 (O_2981,N_29936,N_29028);
and UO_2982 (O_2982,N_29712,N_28986);
or UO_2983 (O_2983,N_29123,N_29318);
nor UO_2984 (O_2984,N_29756,N_29645);
and UO_2985 (O_2985,N_29040,N_29495);
nor UO_2986 (O_2986,N_29934,N_29502);
nor UO_2987 (O_2987,N_29782,N_29338);
or UO_2988 (O_2988,N_28978,N_29532);
and UO_2989 (O_2989,N_29282,N_29849);
nand UO_2990 (O_2990,N_29858,N_28976);
nand UO_2991 (O_2991,N_29362,N_28893);
xor UO_2992 (O_2992,N_29182,N_29748);
nor UO_2993 (O_2993,N_29933,N_28953);
nor UO_2994 (O_2994,N_29249,N_29137);
xnor UO_2995 (O_2995,N_29701,N_29444);
or UO_2996 (O_2996,N_28840,N_29955);
nand UO_2997 (O_2997,N_29994,N_29833);
and UO_2998 (O_2998,N_29292,N_29506);
xor UO_2999 (O_2999,N_29191,N_29996);
nand UO_3000 (O_3000,N_29290,N_28990);
nor UO_3001 (O_3001,N_29768,N_29818);
xnor UO_3002 (O_3002,N_29828,N_29612);
nor UO_3003 (O_3003,N_29886,N_28908);
and UO_3004 (O_3004,N_29519,N_29621);
xnor UO_3005 (O_3005,N_29175,N_29321);
xor UO_3006 (O_3006,N_29512,N_29268);
or UO_3007 (O_3007,N_29634,N_28803);
xor UO_3008 (O_3008,N_29449,N_29218);
nor UO_3009 (O_3009,N_29745,N_29505);
xor UO_3010 (O_3010,N_29496,N_29080);
nor UO_3011 (O_3011,N_29948,N_29949);
nor UO_3012 (O_3012,N_29085,N_29304);
or UO_3013 (O_3013,N_29232,N_29730);
xor UO_3014 (O_3014,N_29509,N_29416);
or UO_3015 (O_3015,N_29960,N_29331);
and UO_3016 (O_3016,N_29389,N_29847);
nand UO_3017 (O_3017,N_29737,N_28916);
nor UO_3018 (O_3018,N_29397,N_29820);
and UO_3019 (O_3019,N_29248,N_28992);
nor UO_3020 (O_3020,N_29664,N_29511);
and UO_3021 (O_3021,N_29580,N_29610);
nand UO_3022 (O_3022,N_29163,N_29718);
xor UO_3023 (O_3023,N_29265,N_29928);
nand UO_3024 (O_3024,N_29794,N_29801);
or UO_3025 (O_3025,N_28896,N_29565);
nor UO_3026 (O_3026,N_29765,N_29322);
nand UO_3027 (O_3027,N_29776,N_28834);
nor UO_3028 (O_3028,N_29307,N_29478);
xor UO_3029 (O_3029,N_28962,N_29907);
and UO_3030 (O_3030,N_28835,N_28854);
nand UO_3031 (O_3031,N_29788,N_29076);
nor UO_3032 (O_3032,N_29918,N_29892);
xor UO_3033 (O_3033,N_29059,N_29988);
or UO_3034 (O_3034,N_29973,N_29715);
and UO_3035 (O_3035,N_29307,N_29162);
nor UO_3036 (O_3036,N_29570,N_28804);
and UO_3037 (O_3037,N_29183,N_29130);
nand UO_3038 (O_3038,N_29820,N_29597);
and UO_3039 (O_3039,N_29247,N_29215);
or UO_3040 (O_3040,N_28969,N_29039);
or UO_3041 (O_3041,N_29321,N_28921);
nand UO_3042 (O_3042,N_29785,N_29914);
and UO_3043 (O_3043,N_29883,N_29027);
xnor UO_3044 (O_3044,N_29528,N_29932);
xor UO_3045 (O_3045,N_29221,N_29704);
nand UO_3046 (O_3046,N_29617,N_29628);
xor UO_3047 (O_3047,N_29505,N_28856);
nand UO_3048 (O_3048,N_29822,N_29452);
nand UO_3049 (O_3049,N_29507,N_29286);
and UO_3050 (O_3050,N_29403,N_29536);
nor UO_3051 (O_3051,N_29285,N_29112);
xor UO_3052 (O_3052,N_29581,N_29604);
nand UO_3053 (O_3053,N_29361,N_29854);
nor UO_3054 (O_3054,N_29383,N_29772);
nand UO_3055 (O_3055,N_29222,N_28874);
nor UO_3056 (O_3056,N_29703,N_29693);
nand UO_3057 (O_3057,N_28928,N_29283);
and UO_3058 (O_3058,N_29568,N_29350);
nand UO_3059 (O_3059,N_29650,N_29624);
nand UO_3060 (O_3060,N_29652,N_29476);
or UO_3061 (O_3061,N_29473,N_29858);
xor UO_3062 (O_3062,N_29637,N_28830);
and UO_3063 (O_3063,N_29105,N_29070);
or UO_3064 (O_3064,N_28821,N_29439);
or UO_3065 (O_3065,N_29483,N_28809);
or UO_3066 (O_3066,N_29778,N_29877);
and UO_3067 (O_3067,N_29343,N_29959);
nand UO_3068 (O_3068,N_29691,N_29226);
or UO_3069 (O_3069,N_29472,N_29389);
and UO_3070 (O_3070,N_29940,N_29210);
nor UO_3071 (O_3071,N_29791,N_29067);
or UO_3072 (O_3072,N_29843,N_29810);
nor UO_3073 (O_3073,N_29298,N_28811);
nor UO_3074 (O_3074,N_29203,N_29084);
nand UO_3075 (O_3075,N_29226,N_29191);
nor UO_3076 (O_3076,N_29038,N_29752);
or UO_3077 (O_3077,N_29123,N_29437);
xor UO_3078 (O_3078,N_29618,N_29557);
or UO_3079 (O_3079,N_29975,N_29399);
or UO_3080 (O_3080,N_29207,N_29286);
or UO_3081 (O_3081,N_29378,N_29242);
xnor UO_3082 (O_3082,N_28893,N_28844);
nor UO_3083 (O_3083,N_29492,N_29780);
xnor UO_3084 (O_3084,N_29620,N_29768);
nand UO_3085 (O_3085,N_29647,N_29749);
nand UO_3086 (O_3086,N_28931,N_29195);
and UO_3087 (O_3087,N_29189,N_29322);
nor UO_3088 (O_3088,N_29449,N_29414);
and UO_3089 (O_3089,N_28888,N_29723);
and UO_3090 (O_3090,N_29050,N_29864);
nand UO_3091 (O_3091,N_29420,N_28994);
and UO_3092 (O_3092,N_29467,N_29755);
or UO_3093 (O_3093,N_29405,N_29563);
nor UO_3094 (O_3094,N_28923,N_29503);
nor UO_3095 (O_3095,N_29452,N_29933);
and UO_3096 (O_3096,N_29747,N_29881);
nand UO_3097 (O_3097,N_29654,N_29139);
and UO_3098 (O_3098,N_29941,N_29593);
nor UO_3099 (O_3099,N_29080,N_29485);
xor UO_3100 (O_3100,N_28811,N_29435);
xnor UO_3101 (O_3101,N_29944,N_28940);
nor UO_3102 (O_3102,N_28843,N_29662);
nand UO_3103 (O_3103,N_29071,N_29246);
xor UO_3104 (O_3104,N_29782,N_29801);
or UO_3105 (O_3105,N_29606,N_29830);
nand UO_3106 (O_3106,N_29296,N_29241);
or UO_3107 (O_3107,N_29174,N_29718);
nor UO_3108 (O_3108,N_29562,N_29980);
and UO_3109 (O_3109,N_29142,N_28915);
and UO_3110 (O_3110,N_29984,N_29093);
xor UO_3111 (O_3111,N_29753,N_29825);
or UO_3112 (O_3112,N_29187,N_29361);
nor UO_3113 (O_3113,N_29879,N_29786);
and UO_3114 (O_3114,N_29536,N_29138);
xor UO_3115 (O_3115,N_29687,N_29558);
and UO_3116 (O_3116,N_29152,N_28983);
nand UO_3117 (O_3117,N_29472,N_28801);
and UO_3118 (O_3118,N_29887,N_29956);
or UO_3119 (O_3119,N_28917,N_29757);
nand UO_3120 (O_3120,N_29521,N_29304);
nor UO_3121 (O_3121,N_28850,N_29080);
and UO_3122 (O_3122,N_29594,N_29585);
nand UO_3123 (O_3123,N_29459,N_29424);
nand UO_3124 (O_3124,N_29042,N_29471);
xnor UO_3125 (O_3125,N_29524,N_29889);
nand UO_3126 (O_3126,N_29697,N_28813);
xnor UO_3127 (O_3127,N_29369,N_29800);
nand UO_3128 (O_3128,N_29738,N_28911);
nand UO_3129 (O_3129,N_29953,N_29028);
and UO_3130 (O_3130,N_28984,N_29029);
xnor UO_3131 (O_3131,N_29799,N_28841);
xnor UO_3132 (O_3132,N_29139,N_29757);
and UO_3133 (O_3133,N_29083,N_29524);
or UO_3134 (O_3134,N_29667,N_28964);
or UO_3135 (O_3135,N_28964,N_29837);
nand UO_3136 (O_3136,N_29671,N_29646);
nor UO_3137 (O_3137,N_28863,N_29368);
nor UO_3138 (O_3138,N_29513,N_29184);
nor UO_3139 (O_3139,N_29664,N_29047);
nor UO_3140 (O_3140,N_29529,N_29937);
nand UO_3141 (O_3141,N_29618,N_29120);
and UO_3142 (O_3142,N_29405,N_29054);
xor UO_3143 (O_3143,N_29246,N_29742);
xnor UO_3144 (O_3144,N_29225,N_29647);
xnor UO_3145 (O_3145,N_29428,N_29998);
nand UO_3146 (O_3146,N_28804,N_29748);
or UO_3147 (O_3147,N_29067,N_29146);
and UO_3148 (O_3148,N_29860,N_29694);
nor UO_3149 (O_3149,N_28849,N_28839);
nor UO_3150 (O_3150,N_29830,N_29512);
xnor UO_3151 (O_3151,N_29578,N_29018);
or UO_3152 (O_3152,N_29772,N_29238);
nor UO_3153 (O_3153,N_29997,N_29609);
or UO_3154 (O_3154,N_28918,N_28941);
and UO_3155 (O_3155,N_29952,N_29587);
and UO_3156 (O_3156,N_29335,N_29569);
nor UO_3157 (O_3157,N_29294,N_29462);
nand UO_3158 (O_3158,N_29169,N_29767);
or UO_3159 (O_3159,N_29302,N_29666);
and UO_3160 (O_3160,N_29250,N_28875);
xnor UO_3161 (O_3161,N_29516,N_29410);
nand UO_3162 (O_3162,N_29859,N_29198);
nor UO_3163 (O_3163,N_29968,N_29672);
nand UO_3164 (O_3164,N_28993,N_29635);
or UO_3165 (O_3165,N_28915,N_29846);
and UO_3166 (O_3166,N_28910,N_29808);
or UO_3167 (O_3167,N_28823,N_29025);
xnor UO_3168 (O_3168,N_29161,N_29589);
nand UO_3169 (O_3169,N_29401,N_29286);
or UO_3170 (O_3170,N_29247,N_29939);
nand UO_3171 (O_3171,N_29950,N_29366);
nand UO_3172 (O_3172,N_29221,N_29624);
xor UO_3173 (O_3173,N_29607,N_29717);
nand UO_3174 (O_3174,N_29683,N_28977);
nor UO_3175 (O_3175,N_29148,N_29462);
xor UO_3176 (O_3176,N_29872,N_29076);
nor UO_3177 (O_3177,N_29967,N_29434);
xnor UO_3178 (O_3178,N_29572,N_29700);
and UO_3179 (O_3179,N_29940,N_28824);
nand UO_3180 (O_3180,N_29687,N_29091);
or UO_3181 (O_3181,N_29374,N_28901);
nand UO_3182 (O_3182,N_28813,N_28984);
or UO_3183 (O_3183,N_29175,N_28901);
xor UO_3184 (O_3184,N_28865,N_29468);
nand UO_3185 (O_3185,N_29111,N_29251);
xnor UO_3186 (O_3186,N_29744,N_29938);
nor UO_3187 (O_3187,N_29608,N_29431);
nand UO_3188 (O_3188,N_29711,N_29750);
or UO_3189 (O_3189,N_29849,N_29948);
nand UO_3190 (O_3190,N_29244,N_29040);
and UO_3191 (O_3191,N_29054,N_29866);
and UO_3192 (O_3192,N_29399,N_29501);
and UO_3193 (O_3193,N_28907,N_28949);
or UO_3194 (O_3194,N_29696,N_29752);
and UO_3195 (O_3195,N_29178,N_29736);
or UO_3196 (O_3196,N_29928,N_29331);
nand UO_3197 (O_3197,N_29019,N_29914);
and UO_3198 (O_3198,N_29868,N_29468);
or UO_3199 (O_3199,N_29317,N_29444);
nand UO_3200 (O_3200,N_29737,N_29589);
nand UO_3201 (O_3201,N_28805,N_29876);
nor UO_3202 (O_3202,N_29866,N_29942);
nand UO_3203 (O_3203,N_28958,N_29290);
nor UO_3204 (O_3204,N_29035,N_29939);
xnor UO_3205 (O_3205,N_28930,N_29403);
xnor UO_3206 (O_3206,N_29490,N_29843);
xnor UO_3207 (O_3207,N_29352,N_29450);
nand UO_3208 (O_3208,N_28997,N_29728);
nand UO_3209 (O_3209,N_29436,N_29380);
xnor UO_3210 (O_3210,N_29713,N_29689);
and UO_3211 (O_3211,N_29119,N_29859);
and UO_3212 (O_3212,N_29728,N_29246);
or UO_3213 (O_3213,N_29923,N_29772);
or UO_3214 (O_3214,N_29263,N_29865);
nor UO_3215 (O_3215,N_29292,N_29959);
xor UO_3216 (O_3216,N_28895,N_29443);
nor UO_3217 (O_3217,N_29706,N_29345);
and UO_3218 (O_3218,N_28906,N_29638);
or UO_3219 (O_3219,N_29589,N_28820);
nand UO_3220 (O_3220,N_29494,N_29960);
and UO_3221 (O_3221,N_29337,N_29346);
and UO_3222 (O_3222,N_29784,N_29422);
or UO_3223 (O_3223,N_29212,N_29135);
or UO_3224 (O_3224,N_29592,N_28865);
or UO_3225 (O_3225,N_29857,N_29446);
and UO_3226 (O_3226,N_29915,N_29350);
or UO_3227 (O_3227,N_29395,N_28802);
or UO_3228 (O_3228,N_28988,N_29116);
or UO_3229 (O_3229,N_29228,N_28950);
xor UO_3230 (O_3230,N_29458,N_29095);
nand UO_3231 (O_3231,N_29910,N_29885);
and UO_3232 (O_3232,N_29752,N_28850);
or UO_3233 (O_3233,N_29528,N_28820);
nand UO_3234 (O_3234,N_28856,N_28981);
nor UO_3235 (O_3235,N_28927,N_29333);
xnor UO_3236 (O_3236,N_28920,N_29597);
nor UO_3237 (O_3237,N_28941,N_29938);
and UO_3238 (O_3238,N_29969,N_28976);
nor UO_3239 (O_3239,N_29457,N_29640);
or UO_3240 (O_3240,N_29838,N_29404);
nand UO_3241 (O_3241,N_29513,N_29496);
xnor UO_3242 (O_3242,N_29892,N_29545);
nand UO_3243 (O_3243,N_29272,N_29190);
nor UO_3244 (O_3244,N_29729,N_29586);
nand UO_3245 (O_3245,N_28850,N_29166);
nand UO_3246 (O_3246,N_29053,N_29313);
nor UO_3247 (O_3247,N_29673,N_29859);
and UO_3248 (O_3248,N_29945,N_29336);
or UO_3249 (O_3249,N_29959,N_29198);
and UO_3250 (O_3250,N_29459,N_29636);
nand UO_3251 (O_3251,N_28840,N_28835);
xor UO_3252 (O_3252,N_29313,N_29213);
or UO_3253 (O_3253,N_29794,N_29322);
nor UO_3254 (O_3254,N_29468,N_29682);
and UO_3255 (O_3255,N_29818,N_29774);
nand UO_3256 (O_3256,N_29192,N_29155);
xnor UO_3257 (O_3257,N_29495,N_28888);
xnor UO_3258 (O_3258,N_29898,N_29697);
and UO_3259 (O_3259,N_28821,N_29074);
and UO_3260 (O_3260,N_29463,N_29604);
nor UO_3261 (O_3261,N_29276,N_29774);
and UO_3262 (O_3262,N_29191,N_29422);
or UO_3263 (O_3263,N_29903,N_29633);
nand UO_3264 (O_3264,N_29207,N_29851);
or UO_3265 (O_3265,N_28843,N_28859);
xor UO_3266 (O_3266,N_29247,N_29923);
and UO_3267 (O_3267,N_29511,N_29480);
nor UO_3268 (O_3268,N_29055,N_28881);
nor UO_3269 (O_3269,N_29864,N_29526);
xor UO_3270 (O_3270,N_29926,N_29014);
nand UO_3271 (O_3271,N_29602,N_29730);
nand UO_3272 (O_3272,N_29682,N_29689);
xnor UO_3273 (O_3273,N_29860,N_29091);
xor UO_3274 (O_3274,N_29812,N_29351);
xor UO_3275 (O_3275,N_29053,N_29928);
or UO_3276 (O_3276,N_29322,N_29153);
and UO_3277 (O_3277,N_29260,N_29550);
nand UO_3278 (O_3278,N_28809,N_29728);
and UO_3279 (O_3279,N_28972,N_29677);
and UO_3280 (O_3280,N_28819,N_29667);
and UO_3281 (O_3281,N_29550,N_29119);
nand UO_3282 (O_3282,N_29874,N_29776);
and UO_3283 (O_3283,N_29203,N_29712);
and UO_3284 (O_3284,N_29653,N_29405);
and UO_3285 (O_3285,N_29051,N_29069);
or UO_3286 (O_3286,N_29777,N_29923);
or UO_3287 (O_3287,N_28949,N_28872);
nand UO_3288 (O_3288,N_29066,N_29398);
nand UO_3289 (O_3289,N_29349,N_29130);
nor UO_3290 (O_3290,N_29101,N_29440);
xor UO_3291 (O_3291,N_29683,N_29451);
nor UO_3292 (O_3292,N_29809,N_29748);
nor UO_3293 (O_3293,N_29797,N_29855);
xnor UO_3294 (O_3294,N_29574,N_29724);
xnor UO_3295 (O_3295,N_29690,N_29120);
nand UO_3296 (O_3296,N_29465,N_29451);
and UO_3297 (O_3297,N_29825,N_28864);
or UO_3298 (O_3298,N_29041,N_29582);
nand UO_3299 (O_3299,N_29249,N_28895);
and UO_3300 (O_3300,N_29882,N_29201);
or UO_3301 (O_3301,N_29946,N_28981);
xor UO_3302 (O_3302,N_29408,N_28884);
nor UO_3303 (O_3303,N_29073,N_29040);
and UO_3304 (O_3304,N_29649,N_29449);
nand UO_3305 (O_3305,N_29104,N_29442);
nand UO_3306 (O_3306,N_29979,N_29894);
nand UO_3307 (O_3307,N_29263,N_28804);
and UO_3308 (O_3308,N_29011,N_29761);
or UO_3309 (O_3309,N_28920,N_29382);
or UO_3310 (O_3310,N_29263,N_29246);
xor UO_3311 (O_3311,N_29619,N_29139);
nand UO_3312 (O_3312,N_29740,N_29604);
or UO_3313 (O_3313,N_29744,N_28893);
and UO_3314 (O_3314,N_29889,N_29922);
nand UO_3315 (O_3315,N_28934,N_29387);
or UO_3316 (O_3316,N_29458,N_29034);
xor UO_3317 (O_3317,N_29706,N_29923);
nor UO_3318 (O_3318,N_29457,N_29536);
or UO_3319 (O_3319,N_29640,N_29125);
xor UO_3320 (O_3320,N_29025,N_29664);
and UO_3321 (O_3321,N_28877,N_28803);
nand UO_3322 (O_3322,N_29678,N_28887);
and UO_3323 (O_3323,N_28879,N_29889);
nand UO_3324 (O_3324,N_29853,N_28913);
nand UO_3325 (O_3325,N_29252,N_29176);
nor UO_3326 (O_3326,N_29762,N_29795);
nor UO_3327 (O_3327,N_29383,N_29602);
xnor UO_3328 (O_3328,N_28945,N_29491);
nor UO_3329 (O_3329,N_29122,N_29314);
xnor UO_3330 (O_3330,N_29675,N_29055);
nor UO_3331 (O_3331,N_28803,N_29215);
nor UO_3332 (O_3332,N_29152,N_29541);
nand UO_3333 (O_3333,N_29294,N_29702);
xor UO_3334 (O_3334,N_29039,N_29562);
or UO_3335 (O_3335,N_29313,N_29312);
and UO_3336 (O_3336,N_28938,N_29693);
xor UO_3337 (O_3337,N_29285,N_29078);
xnor UO_3338 (O_3338,N_28929,N_29457);
and UO_3339 (O_3339,N_28981,N_29442);
nor UO_3340 (O_3340,N_29278,N_29073);
or UO_3341 (O_3341,N_29839,N_29881);
or UO_3342 (O_3342,N_29286,N_28832);
nor UO_3343 (O_3343,N_29415,N_29686);
xnor UO_3344 (O_3344,N_28840,N_29470);
nand UO_3345 (O_3345,N_29723,N_29882);
nor UO_3346 (O_3346,N_29315,N_29836);
nor UO_3347 (O_3347,N_29255,N_29444);
nor UO_3348 (O_3348,N_29040,N_29823);
nand UO_3349 (O_3349,N_29592,N_29060);
or UO_3350 (O_3350,N_29547,N_29149);
and UO_3351 (O_3351,N_29861,N_29541);
or UO_3352 (O_3352,N_29872,N_29078);
nand UO_3353 (O_3353,N_28883,N_28953);
nor UO_3354 (O_3354,N_29658,N_29549);
and UO_3355 (O_3355,N_29106,N_29589);
and UO_3356 (O_3356,N_29407,N_29826);
and UO_3357 (O_3357,N_29625,N_29568);
and UO_3358 (O_3358,N_28823,N_29747);
xor UO_3359 (O_3359,N_29168,N_29679);
xnor UO_3360 (O_3360,N_29773,N_29159);
or UO_3361 (O_3361,N_29883,N_29599);
nor UO_3362 (O_3362,N_29757,N_29745);
or UO_3363 (O_3363,N_29501,N_29865);
nand UO_3364 (O_3364,N_29550,N_28846);
or UO_3365 (O_3365,N_29387,N_29484);
xor UO_3366 (O_3366,N_29329,N_29409);
nor UO_3367 (O_3367,N_29364,N_29008);
or UO_3368 (O_3368,N_29660,N_29817);
nor UO_3369 (O_3369,N_29831,N_29630);
xor UO_3370 (O_3370,N_28828,N_29772);
nor UO_3371 (O_3371,N_29518,N_29947);
and UO_3372 (O_3372,N_29155,N_29612);
and UO_3373 (O_3373,N_28849,N_29299);
nor UO_3374 (O_3374,N_29779,N_28846);
nor UO_3375 (O_3375,N_29453,N_29983);
xor UO_3376 (O_3376,N_29537,N_29139);
or UO_3377 (O_3377,N_28875,N_29315);
nand UO_3378 (O_3378,N_29350,N_29708);
and UO_3379 (O_3379,N_29866,N_29376);
nor UO_3380 (O_3380,N_29227,N_29459);
nand UO_3381 (O_3381,N_29286,N_29869);
or UO_3382 (O_3382,N_29388,N_29417);
and UO_3383 (O_3383,N_28804,N_29573);
nand UO_3384 (O_3384,N_29523,N_29262);
or UO_3385 (O_3385,N_28954,N_29214);
or UO_3386 (O_3386,N_29771,N_29418);
and UO_3387 (O_3387,N_29400,N_29704);
nor UO_3388 (O_3388,N_28854,N_29771);
or UO_3389 (O_3389,N_29985,N_29737);
and UO_3390 (O_3390,N_28860,N_29759);
nand UO_3391 (O_3391,N_29015,N_29980);
nor UO_3392 (O_3392,N_29254,N_29642);
nand UO_3393 (O_3393,N_29762,N_29502);
xnor UO_3394 (O_3394,N_28899,N_29524);
nor UO_3395 (O_3395,N_29494,N_29034);
nand UO_3396 (O_3396,N_29113,N_29114);
nor UO_3397 (O_3397,N_29045,N_29223);
or UO_3398 (O_3398,N_29289,N_29534);
and UO_3399 (O_3399,N_29213,N_29089);
xnor UO_3400 (O_3400,N_29397,N_29136);
nor UO_3401 (O_3401,N_29097,N_29449);
and UO_3402 (O_3402,N_29882,N_29532);
or UO_3403 (O_3403,N_28965,N_29620);
nand UO_3404 (O_3404,N_29100,N_29113);
or UO_3405 (O_3405,N_28849,N_29800);
xor UO_3406 (O_3406,N_28814,N_29813);
nand UO_3407 (O_3407,N_29910,N_29115);
nand UO_3408 (O_3408,N_28943,N_29294);
nor UO_3409 (O_3409,N_28892,N_29271);
or UO_3410 (O_3410,N_29551,N_29090);
or UO_3411 (O_3411,N_29177,N_29797);
nand UO_3412 (O_3412,N_29660,N_29393);
or UO_3413 (O_3413,N_29307,N_29073);
and UO_3414 (O_3414,N_28976,N_28862);
nand UO_3415 (O_3415,N_29864,N_29591);
nor UO_3416 (O_3416,N_29707,N_29358);
nand UO_3417 (O_3417,N_29187,N_28880);
nor UO_3418 (O_3418,N_29352,N_29809);
xor UO_3419 (O_3419,N_29261,N_29509);
or UO_3420 (O_3420,N_29109,N_29273);
nor UO_3421 (O_3421,N_29569,N_29526);
and UO_3422 (O_3422,N_29109,N_29635);
nand UO_3423 (O_3423,N_29205,N_29336);
or UO_3424 (O_3424,N_29445,N_28875);
nand UO_3425 (O_3425,N_29323,N_29415);
nor UO_3426 (O_3426,N_29017,N_29844);
nor UO_3427 (O_3427,N_29153,N_29495);
and UO_3428 (O_3428,N_29335,N_29668);
and UO_3429 (O_3429,N_29312,N_29099);
and UO_3430 (O_3430,N_29955,N_29352);
nand UO_3431 (O_3431,N_29678,N_29548);
nor UO_3432 (O_3432,N_29883,N_28979);
or UO_3433 (O_3433,N_29064,N_29445);
xor UO_3434 (O_3434,N_29573,N_28824);
nor UO_3435 (O_3435,N_29764,N_29356);
nand UO_3436 (O_3436,N_28889,N_29124);
and UO_3437 (O_3437,N_29453,N_29395);
nor UO_3438 (O_3438,N_29783,N_29041);
nand UO_3439 (O_3439,N_28912,N_29714);
nor UO_3440 (O_3440,N_29277,N_29214);
nand UO_3441 (O_3441,N_29549,N_29983);
or UO_3442 (O_3442,N_29053,N_29237);
or UO_3443 (O_3443,N_29921,N_29156);
and UO_3444 (O_3444,N_29776,N_29116);
nand UO_3445 (O_3445,N_29038,N_28818);
xnor UO_3446 (O_3446,N_29746,N_29309);
nand UO_3447 (O_3447,N_29595,N_29932);
or UO_3448 (O_3448,N_29031,N_29037);
xnor UO_3449 (O_3449,N_29779,N_29883);
or UO_3450 (O_3450,N_28955,N_28891);
and UO_3451 (O_3451,N_29193,N_29270);
xnor UO_3452 (O_3452,N_29017,N_29178);
and UO_3453 (O_3453,N_29359,N_29106);
and UO_3454 (O_3454,N_29658,N_28968);
and UO_3455 (O_3455,N_28918,N_29886);
xor UO_3456 (O_3456,N_28805,N_29287);
nand UO_3457 (O_3457,N_29528,N_29443);
xor UO_3458 (O_3458,N_29903,N_29935);
xor UO_3459 (O_3459,N_29486,N_28819);
nor UO_3460 (O_3460,N_28934,N_28921);
nand UO_3461 (O_3461,N_28860,N_29156);
xor UO_3462 (O_3462,N_29973,N_29003);
nor UO_3463 (O_3463,N_29746,N_29883);
xor UO_3464 (O_3464,N_29437,N_29768);
nor UO_3465 (O_3465,N_29230,N_29564);
and UO_3466 (O_3466,N_29914,N_29311);
xor UO_3467 (O_3467,N_29766,N_29194);
and UO_3468 (O_3468,N_29444,N_29795);
xor UO_3469 (O_3469,N_29018,N_29280);
and UO_3470 (O_3470,N_28808,N_29702);
nor UO_3471 (O_3471,N_29710,N_29470);
xor UO_3472 (O_3472,N_29220,N_29573);
nand UO_3473 (O_3473,N_29984,N_28905);
and UO_3474 (O_3474,N_29692,N_29748);
nand UO_3475 (O_3475,N_28855,N_29382);
xor UO_3476 (O_3476,N_28894,N_29315);
and UO_3477 (O_3477,N_29026,N_28822);
nand UO_3478 (O_3478,N_29212,N_29285);
and UO_3479 (O_3479,N_29676,N_29362);
xnor UO_3480 (O_3480,N_29230,N_29656);
and UO_3481 (O_3481,N_28937,N_29670);
xnor UO_3482 (O_3482,N_29087,N_29017);
or UO_3483 (O_3483,N_29078,N_29624);
and UO_3484 (O_3484,N_29403,N_29389);
nand UO_3485 (O_3485,N_29935,N_29398);
and UO_3486 (O_3486,N_29079,N_29141);
or UO_3487 (O_3487,N_29599,N_29944);
xor UO_3488 (O_3488,N_29105,N_29055);
nor UO_3489 (O_3489,N_29602,N_29099);
and UO_3490 (O_3490,N_28976,N_29299);
or UO_3491 (O_3491,N_29064,N_29245);
and UO_3492 (O_3492,N_29148,N_29683);
xnor UO_3493 (O_3493,N_28884,N_29484);
and UO_3494 (O_3494,N_29487,N_29385);
xor UO_3495 (O_3495,N_29810,N_29491);
xnor UO_3496 (O_3496,N_29574,N_29301);
nor UO_3497 (O_3497,N_29960,N_28935);
nand UO_3498 (O_3498,N_29135,N_29140);
xnor UO_3499 (O_3499,N_28840,N_29818);
endmodule