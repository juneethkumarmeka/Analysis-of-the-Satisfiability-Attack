module basic_1500_15000_2000_60_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_425,In_960);
nor U1 (N_1,In_850,In_1260);
xnor U2 (N_2,In_1246,In_1374);
nand U3 (N_3,In_1438,In_940);
or U4 (N_4,In_456,In_1497);
nand U5 (N_5,In_1489,In_1253);
xnor U6 (N_6,In_621,In_1069);
nor U7 (N_7,In_970,In_293);
nand U8 (N_8,In_570,In_1272);
and U9 (N_9,In_827,In_934);
nor U10 (N_10,In_734,In_202);
xor U11 (N_11,In_890,In_330);
nor U12 (N_12,In_180,In_463);
nand U13 (N_13,In_925,In_1393);
xnor U14 (N_14,In_525,In_259);
nand U15 (N_15,In_1238,In_955);
or U16 (N_16,In_709,In_279);
or U17 (N_17,In_181,In_365);
nor U18 (N_18,In_312,In_167);
and U19 (N_19,In_37,In_1402);
xnor U20 (N_20,In_27,In_1234);
xor U21 (N_21,In_383,In_521);
nor U22 (N_22,In_922,In_1405);
xor U23 (N_23,In_134,In_944);
and U24 (N_24,In_1353,In_711);
xnor U25 (N_25,In_1040,In_904);
or U26 (N_26,In_154,In_580);
or U27 (N_27,In_208,In_1248);
xor U28 (N_28,In_842,In_986);
nand U29 (N_29,In_227,In_978);
or U30 (N_30,In_856,In_1134);
and U31 (N_31,In_691,In_1109);
xnor U32 (N_32,In_651,In_880);
or U33 (N_33,In_1154,In_1148);
or U34 (N_34,In_913,In_1233);
nand U35 (N_35,In_561,In_921);
nor U36 (N_36,In_1344,In_398);
nand U37 (N_37,In_1059,In_1219);
and U38 (N_38,In_417,In_1472);
nand U39 (N_39,In_1217,In_1301);
and U40 (N_40,In_1195,In_286);
or U41 (N_41,In_1048,In_531);
xor U42 (N_42,In_1007,In_733);
and U43 (N_43,In_83,In_229);
nor U44 (N_44,In_1172,In_67);
xnor U45 (N_45,In_624,In_1485);
xnor U46 (N_46,In_1076,In_53);
and U47 (N_47,In_1243,In_1196);
nor U48 (N_48,In_581,In_720);
nor U49 (N_49,In_1403,In_794);
or U50 (N_50,In_716,In_341);
xor U51 (N_51,In_451,In_24);
and U52 (N_52,In_269,In_1444);
and U53 (N_53,In_32,In_697);
nand U54 (N_54,In_9,In_297);
xnor U55 (N_55,In_798,In_1292);
nor U56 (N_56,In_681,In_834);
and U57 (N_57,In_1269,In_975);
xor U58 (N_58,In_1095,In_482);
nand U59 (N_59,In_657,In_1187);
nor U60 (N_60,In_433,In_757);
nor U61 (N_61,In_26,In_888);
and U62 (N_62,In_1481,In_548);
and U63 (N_63,In_1035,In_1430);
nor U64 (N_64,In_828,In_635);
xor U65 (N_65,In_427,In_443);
or U66 (N_66,In_864,In_614);
nand U67 (N_67,In_1005,In_1369);
nand U68 (N_68,In_675,In_424);
nand U69 (N_69,In_1370,In_1279);
xor U70 (N_70,In_680,In_568);
or U71 (N_71,In_644,In_1070);
or U72 (N_72,In_305,In_186);
and U73 (N_73,In_722,In_1491);
or U74 (N_74,In_349,In_141);
xnor U75 (N_75,In_194,In_846);
or U76 (N_76,In_240,In_615);
or U77 (N_77,In_1063,In_72);
nor U78 (N_78,In_15,In_1051);
nor U79 (N_79,In_235,In_324);
or U80 (N_80,In_679,In_800);
or U81 (N_81,In_1214,In_52);
nor U82 (N_82,In_549,In_1469);
nor U83 (N_83,In_1262,In_873);
or U84 (N_84,In_225,In_566);
xnor U85 (N_85,In_164,In_489);
and U86 (N_86,In_105,In_737);
xor U87 (N_87,In_589,In_1323);
xnor U88 (N_88,In_968,In_152);
and U89 (N_89,In_1457,In_303);
nand U90 (N_90,In_1064,In_830);
or U91 (N_91,In_162,In_402);
nand U92 (N_92,In_1437,In_376);
nor U93 (N_93,In_1170,In_380);
and U94 (N_94,In_518,In_1387);
and U95 (N_95,In_1454,In_1399);
or U96 (N_96,In_1021,In_599);
or U97 (N_97,In_719,In_177);
nor U98 (N_98,In_881,In_811);
nor U99 (N_99,In_564,In_163);
nor U100 (N_100,In_511,In_1442);
or U101 (N_101,In_223,In_682);
or U102 (N_102,In_192,In_1098);
xnor U103 (N_103,In_1421,In_853);
and U104 (N_104,In_677,In_209);
nor U105 (N_105,In_1322,In_1382);
or U106 (N_106,In_928,In_1299);
nand U107 (N_107,In_203,In_1346);
nand U108 (N_108,In_434,In_1014);
and U109 (N_109,In_779,In_702);
or U110 (N_110,In_470,In_40);
or U111 (N_111,In_284,In_438);
xor U112 (N_112,In_301,In_870);
xor U113 (N_113,In_1397,In_497);
xnor U114 (N_114,In_686,In_997);
nor U115 (N_115,In_260,In_810);
nand U116 (N_116,In_1389,In_360);
xnor U117 (N_117,In_546,In_507);
or U118 (N_118,In_732,In_1441);
or U119 (N_119,In_748,In_1097);
nor U120 (N_120,In_887,In_1255);
or U121 (N_121,In_1153,In_288);
nor U122 (N_122,In_385,In_1293);
or U123 (N_123,In_619,In_275);
nor U124 (N_124,In_900,In_941);
or U125 (N_125,In_325,In_1462);
nor U126 (N_126,In_761,In_1202);
nand U127 (N_127,In_854,In_1254);
xor U128 (N_128,In_819,In_661);
and U129 (N_129,In_1045,In_1455);
or U130 (N_130,In_1194,In_1203);
and U131 (N_131,In_1288,In_1065);
nor U132 (N_132,In_444,In_122);
nor U133 (N_133,In_161,In_1365);
and U134 (N_134,In_419,In_65);
xor U135 (N_135,In_1416,In_442);
or U136 (N_136,In_769,In_1006);
xnor U137 (N_137,In_1345,In_465);
or U138 (N_138,In_658,In_204);
nand U139 (N_139,In_622,In_406);
and U140 (N_140,In_504,In_1114);
and U141 (N_141,In_829,In_704);
nand U142 (N_142,In_191,In_1314);
nand U143 (N_143,In_572,In_958);
xnor U144 (N_144,In_1074,In_573);
nor U145 (N_145,In_613,In_195);
nand U146 (N_146,In_266,In_347);
nand U147 (N_147,In_458,In_950);
or U148 (N_148,In_1499,In_375);
and U149 (N_149,In_1230,In_1132);
nor U150 (N_150,In_539,In_1049);
and U151 (N_151,In_1282,In_440);
nand U152 (N_152,In_1464,In_1424);
nand U153 (N_153,In_1380,In_176);
nor U154 (N_154,In_1107,In_1036);
or U155 (N_155,In_633,In_281);
or U156 (N_156,In_236,In_781);
or U157 (N_157,In_0,In_481);
nand U158 (N_158,In_1024,In_931);
and U159 (N_159,In_653,In_963);
nand U160 (N_160,In_1081,In_588);
xor U161 (N_161,In_961,In_821);
xor U162 (N_162,In_1037,In_1259);
and U163 (N_163,In_724,In_608);
or U164 (N_164,In_58,In_1326);
nand U165 (N_165,In_807,In_607);
nor U166 (N_166,In_108,In_1027);
nor U167 (N_167,In_714,In_538);
nor U168 (N_168,In_1088,In_35);
nand U169 (N_169,In_1354,In_1155);
and U170 (N_170,In_517,In_1392);
nor U171 (N_171,In_390,In_144);
nand U172 (N_172,In_584,In_774);
nand U173 (N_173,In_1117,In_678);
xor U174 (N_174,In_824,In_315);
or U175 (N_175,In_796,In_468);
or U176 (N_176,In_1276,In_1342);
and U177 (N_177,In_61,In_535);
nand U178 (N_178,In_418,In_50);
and U179 (N_179,In_252,In_1480);
or U180 (N_180,In_1284,In_377);
nand U181 (N_181,In_715,In_1164);
nand U182 (N_182,In_946,In_78);
and U183 (N_183,In_731,In_1015);
xnor U184 (N_184,In_578,In_1016);
nor U185 (N_185,In_201,In_693);
nand U186 (N_186,In_413,In_338);
nand U187 (N_187,In_1283,In_415);
nand U188 (N_188,In_778,In_519);
or U189 (N_189,In_1332,In_363);
nand U190 (N_190,In_687,In_471);
or U191 (N_191,In_1307,In_759);
or U192 (N_192,In_1275,In_554);
nand U193 (N_193,In_562,In_802);
nor U194 (N_194,In_373,In_1029);
or U195 (N_195,In_66,In_983);
and U196 (N_196,In_1384,In_1433);
nand U197 (N_197,In_903,In_649);
nand U198 (N_198,In_927,In_1108);
nand U199 (N_199,In_212,In_1092);
or U200 (N_200,In_909,In_250);
nor U201 (N_201,In_871,In_908);
nand U202 (N_202,In_22,In_896);
and U203 (N_203,In_689,In_220);
and U204 (N_204,In_1483,In_1038);
nor U205 (N_205,In_60,In_547);
nand U206 (N_206,In_1308,In_454);
nor U207 (N_207,In_117,In_1476);
or U208 (N_208,In_912,In_910);
nor U209 (N_209,In_1319,In_1366);
nand U210 (N_210,In_938,In_1042);
xnor U211 (N_211,In_1337,In_1305);
nor U212 (N_212,In_1482,In_1136);
nor U213 (N_213,In_175,In_787);
nor U214 (N_214,In_1010,In_645);
nor U215 (N_215,In_763,In_891);
nor U216 (N_216,In_487,In_1329);
and U217 (N_217,In_740,In_82);
or U218 (N_218,In_1463,In_104);
and U219 (N_219,In_48,In_1343);
or U220 (N_220,In_1071,In_858);
xnor U221 (N_221,In_47,In_309);
nand U222 (N_222,In_876,In_1102);
and U223 (N_223,In_118,In_728);
xor U224 (N_224,In_1199,In_1213);
or U225 (N_225,In_845,In_94);
nand U226 (N_226,In_437,In_1075);
or U227 (N_227,In_636,In_1356);
xnor U228 (N_228,In_1298,In_472);
or U229 (N_229,In_1300,In_508);
and U230 (N_230,In_46,In_1443);
and U231 (N_231,In_1394,In_1122);
nor U232 (N_232,In_905,In_157);
and U233 (N_233,In_762,In_1495);
nor U234 (N_234,In_1285,In_1104);
nand U235 (N_235,In_294,In_848);
or U236 (N_236,In_966,In_1336);
nor U237 (N_237,In_491,In_626);
and U238 (N_238,In_972,In_337);
and U239 (N_239,In_857,In_295);
and U240 (N_240,In_1414,In_182);
and U241 (N_241,In_1296,In_1079);
nand U242 (N_242,In_127,In_285);
xor U243 (N_243,In_883,In_701);
nor U244 (N_244,In_129,In_92);
or U245 (N_245,In_1101,In_1486);
nand U246 (N_246,In_973,In_628);
nor U247 (N_247,In_964,In_348);
nor U248 (N_248,In_1177,In_289);
nor U249 (N_249,In_34,In_838);
or U250 (N_250,In_115,In_1189);
xor U251 (N_251,In_727,In_1140);
or U252 (N_252,In_782,In_673);
or U253 (N_253,In_300,In_1341);
and U254 (N_254,In_710,In_461);
or U255 (N_255,In_1182,In_149);
nand U256 (N_256,In_261,In_110);
xor U257 (N_257,In_1458,In_1431);
nor U258 (N_258,In_1426,In_1432);
nand U259 (N_259,In_1496,N_121);
nand U260 (N_260,In_1244,N_21);
nor U261 (N_261,N_130,In_1468);
and U262 (N_262,N_117,In_351);
and U263 (N_263,In_1317,In_918);
and U264 (N_264,In_336,In_290);
and U265 (N_265,In_5,In_13);
or U266 (N_266,N_138,In_1440);
and U267 (N_267,In_216,N_186);
nand U268 (N_268,In_1335,In_1224);
and U269 (N_269,In_768,In_1161);
and U270 (N_270,In_1204,N_29);
nand U271 (N_271,N_239,In_917);
nand U272 (N_272,N_248,In_576);
nor U273 (N_273,In_754,In_746);
nor U274 (N_274,N_32,In_184);
nor U275 (N_275,N_197,N_207);
nor U276 (N_276,In_587,In_1127);
and U277 (N_277,In_685,In_831);
xor U278 (N_278,In_313,In_672);
and U279 (N_279,In_906,In_843);
nand U280 (N_280,In_543,In_902);
nor U281 (N_281,N_61,In_863);
xnor U282 (N_282,In_441,In_1084);
and U283 (N_283,N_70,In_630);
xor U284 (N_284,In_1473,N_203);
xnor U285 (N_285,N_8,In_924);
nor U286 (N_286,In_77,In_473);
or U287 (N_287,In_490,In_89);
nand U288 (N_288,In_382,In_1266);
nor U289 (N_289,In_962,In_1350);
and U290 (N_290,In_1340,N_242);
xnor U291 (N_291,In_793,N_182);
nand U292 (N_292,In_1361,In_460);
nor U293 (N_293,N_38,In_878);
or U294 (N_294,In_1325,In_703);
nor U295 (N_295,N_99,In_999);
and U296 (N_296,In_1239,In_664);
xnor U297 (N_297,In_484,N_216);
or U298 (N_298,In_408,In_151);
or U299 (N_299,N_77,In_23);
xor U300 (N_300,In_291,In_799);
or U301 (N_301,In_91,In_1235);
and U302 (N_302,In_1498,In_270);
nand U303 (N_303,In_190,In_55);
nand U304 (N_304,In_453,N_218);
nor U305 (N_305,In_741,In_1359);
nor U306 (N_306,In_159,In_867);
nand U307 (N_307,In_555,In_1256);
nand U308 (N_308,In_29,N_211);
nand U309 (N_309,In_841,In_1082);
or U310 (N_310,In_1193,In_1228);
xnor U311 (N_311,N_157,N_245);
nand U312 (N_312,In_171,In_1025);
xnor U313 (N_313,In_30,N_233);
nor U314 (N_314,In_1297,In_391);
nor U315 (N_315,In_648,In_17);
nand U316 (N_316,In_1470,In_329);
or U317 (N_317,N_146,In_262);
nand U318 (N_318,N_215,N_148);
xnor U319 (N_319,In_62,In_183);
xor U320 (N_320,In_1068,In_1475);
nor U321 (N_321,In_676,In_1210);
or U322 (N_322,N_9,N_168);
or U323 (N_323,In_659,In_951);
nor U324 (N_324,In_355,In_1218);
nor U325 (N_325,N_170,In_567);
or U326 (N_326,In_31,In_606);
nand U327 (N_327,In_1131,In_1383);
and U328 (N_328,N_178,In_1032);
nand U329 (N_329,In_196,N_217);
xnor U330 (N_330,In_1372,N_22);
nand U331 (N_331,In_529,In_367);
or U332 (N_332,In_977,In_459);
nor U333 (N_333,In_146,In_1115);
nor U334 (N_334,N_185,In_331);
and U335 (N_335,In_920,N_43);
nor U336 (N_336,In_556,In_412);
or U337 (N_337,N_154,In_718);
nand U338 (N_338,In_147,In_1100);
nand U339 (N_339,In_14,In_1080);
xor U340 (N_340,In_1143,In_243);
nand U341 (N_341,In_872,In_911);
or U342 (N_342,In_1197,N_188);
or U343 (N_343,In_985,In_68);
nor U344 (N_344,In_752,In_170);
xor U345 (N_345,N_89,In_852);
xnor U346 (N_346,In_1306,In_1371);
nor U347 (N_347,In_156,In_494);
nor U348 (N_348,In_1106,In_394);
xor U349 (N_349,In_1395,In_590);
and U350 (N_350,N_241,In_945);
or U351 (N_351,In_666,In_447);
xor U352 (N_352,In_1471,In_435);
nor U353 (N_353,In_1287,In_403);
or U354 (N_354,In_323,In_368);
nand U355 (N_355,N_176,In_1004);
nand U356 (N_356,In_839,N_111);
nand U357 (N_357,In_185,In_51);
or U358 (N_358,In_534,In_894);
nand U359 (N_359,In_404,In_276);
and U360 (N_360,In_1000,N_179);
nor U361 (N_361,In_136,N_73);
xnor U362 (N_362,In_421,In_932);
or U363 (N_363,In_1429,In_428);
xnor U364 (N_364,In_1390,N_88);
xor U365 (N_365,In_1240,In_755);
or U366 (N_366,N_166,In_197);
xor U367 (N_367,In_474,N_150);
nor U368 (N_368,In_647,In_875);
nand U369 (N_369,In_1191,N_140);
xor U370 (N_370,In_1033,N_128);
and U371 (N_371,N_230,N_91);
and U372 (N_372,In_1236,In_230);
nor U373 (N_373,In_749,N_172);
xor U374 (N_374,In_935,In_822);
xor U375 (N_375,In_585,In_73);
nor U376 (N_376,In_1111,In_1339);
xnor U377 (N_377,In_967,In_971);
or U378 (N_378,In_102,In_550);
xor U379 (N_379,N_180,In_981);
nand U380 (N_380,In_995,N_87);
or U381 (N_381,In_210,In_885);
nand U382 (N_382,In_1215,In_1351);
xor U383 (N_383,In_751,In_145);
and U384 (N_384,N_227,In_953);
xnor U385 (N_385,N_129,In_825);
nor U386 (N_386,N_11,In_745);
or U387 (N_387,In_1162,In_155);
xnor U388 (N_388,In_299,In_976);
nor U389 (N_389,In_116,N_201);
and U390 (N_390,N_59,In_516);
nor U391 (N_391,In_583,In_1459);
nand U392 (N_392,In_874,In_1252);
xnor U393 (N_393,N_114,In_542);
and U394 (N_394,In_1175,In_1427);
or U395 (N_395,In_1087,N_85);
and U396 (N_396,In_226,In_1205);
nand U397 (N_397,In_231,In_42);
or U398 (N_398,In_892,In_844);
and U399 (N_399,N_127,In_777);
nor U400 (N_400,In_1160,In_321);
xnor U401 (N_401,In_292,In_1188);
xor U402 (N_402,In_334,In_1363);
nand U403 (N_403,In_429,In_1355);
xor U404 (N_404,In_1461,In_274);
or U405 (N_405,In_1302,In_241);
and U406 (N_406,In_221,N_221);
and U407 (N_407,N_28,In_1137);
nand U408 (N_408,In_1099,In_1241);
and U409 (N_409,In_298,In_69);
nor U410 (N_410,N_184,In_948);
nor U411 (N_411,In_609,In_916);
xor U412 (N_412,In_698,N_149);
nand U413 (N_413,In_639,N_205);
or U414 (N_414,In_736,In_610);
nor U415 (N_415,In_860,In_199);
and U416 (N_416,N_57,N_106);
xnor U417 (N_417,In_952,In_586);
xor U418 (N_418,In_837,In_278);
or U419 (N_419,In_1460,In_533);
nand U420 (N_420,In_96,In_646);
xor U421 (N_421,In_1334,In_263);
or U422 (N_422,In_814,In_813);
xnor U423 (N_423,In_1490,In_106);
nand U424 (N_424,In_708,In_317);
nand U425 (N_425,In_123,In_344);
nor U426 (N_426,In_1375,N_229);
xor U427 (N_427,In_253,In_1159);
nor U428 (N_428,In_54,In_283);
nand U429 (N_429,In_1413,In_287);
xor U430 (N_430,N_90,N_35);
or U431 (N_431,In_1477,In_242);
nor U432 (N_432,In_1493,In_114);
nor U433 (N_433,N_18,In_1112);
nand U434 (N_434,In_479,In_462);
xnor U435 (N_435,In_173,In_1453);
and U436 (N_436,In_617,In_717);
nor U437 (N_437,In_3,In_695);
and U438 (N_438,In_322,In_327);
nor U439 (N_439,N_56,In_700);
nand U440 (N_440,In_1220,In_634);
nand U441 (N_441,N_159,N_7);
nor U442 (N_442,In_407,In_816);
and U443 (N_443,In_1123,In_1083);
nand U444 (N_444,In_643,In_574);
xnor U445 (N_445,N_60,N_153);
xor U446 (N_446,In_11,In_744);
and U447 (N_447,In_485,In_7);
xnor U448 (N_448,In_90,In_1022);
nand U449 (N_449,In_805,In_396);
xor U450 (N_450,In_354,In_1373);
and U451 (N_451,N_58,In_1312);
xnor U452 (N_452,In_1418,In_1227);
or U453 (N_453,In_943,In_865);
and U454 (N_454,N_69,N_13);
nor U455 (N_455,In_255,In_801);
and U456 (N_456,N_108,In_1318);
or U457 (N_457,N_173,In_1056);
nand U458 (N_458,In_211,In_1019);
nor U459 (N_459,In_120,N_0);
and U460 (N_460,In_352,In_1352);
nand U461 (N_461,In_1103,In_527);
and U462 (N_462,In_1105,In_809);
or U463 (N_463,N_199,N_143);
nand U464 (N_464,In_1121,N_96);
xnor U465 (N_465,N_19,In_826);
nand U466 (N_466,In_1381,In_445);
or U467 (N_467,In_430,N_17);
nand U468 (N_468,In_353,In_510);
nand U469 (N_469,In_342,In_38);
and U470 (N_470,In_130,In_750);
nand U471 (N_471,In_132,In_773);
nor U472 (N_472,N_16,In_994);
xor U473 (N_473,N_125,In_356);
xnor U474 (N_474,In_742,In_148);
and U475 (N_475,In_565,In_379);
and U476 (N_476,In_1479,In_206);
xnor U477 (N_477,In_650,In_1396);
or U478 (N_478,In_1448,In_1200);
nand U479 (N_479,In_1118,In_1090);
or U480 (N_480,In_81,In_655);
nand U481 (N_481,N_116,In_272);
and U482 (N_482,In_1150,In_1167);
and U483 (N_483,In_6,In_907);
xor U484 (N_484,In_764,In_44);
xnor U485 (N_485,In_99,In_25);
nand U486 (N_486,In_1410,N_231);
nor U487 (N_487,In_1128,In_128);
nor U488 (N_488,In_502,In_1125);
and U489 (N_489,N_47,In_244);
nand U490 (N_490,In_919,N_147);
nand U491 (N_491,In_1133,N_223);
or U492 (N_492,In_1327,In_1261);
nor U493 (N_493,In_256,In_1206);
and U494 (N_494,N_134,In_1057);
xnor U495 (N_495,In_528,In_1169);
or U496 (N_496,N_177,In_1052);
and U497 (N_497,N_26,In_707);
nand U498 (N_498,In_620,In_1411);
or U499 (N_499,In_1278,In_1047);
nand U500 (N_500,In_36,In_862);
and U501 (N_501,N_405,In_604);
nor U502 (N_502,N_175,In_215);
nand U503 (N_503,In_654,N_34);
and U504 (N_504,In_1020,In_12);
xor U505 (N_505,N_246,In_1176);
or U506 (N_506,In_780,In_45);
nand U507 (N_507,N_132,N_66);
nor U508 (N_508,In_254,N_353);
nor U509 (N_509,In_1349,In_739);
and U510 (N_510,In_1331,In_1277);
and U511 (N_511,In_420,N_452);
or U512 (N_512,In_1089,In_205);
nor U513 (N_513,In_815,N_382);
xnor U514 (N_514,In_1321,N_484);
nor U515 (N_515,N_164,N_156);
and U516 (N_516,In_1183,N_6);
or U517 (N_517,N_213,In_467);
or U518 (N_518,In_627,In_1385);
and U519 (N_519,In_868,In_786);
or U520 (N_520,In_135,N_464);
nand U521 (N_521,N_299,N_302);
xnor U522 (N_522,In_597,N_288);
and U523 (N_523,In_452,In_1474);
or U524 (N_524,N_466,In_670);
xor U525 (N_525,N_374,In_178);
or U526 (N_526,In_668,N_133);
xnor U527 (N_527,N_171,N_25);
xor U528 (N_528,In_1237,N_212);
xnor U529 (N_529,In_1046,N_446);
nand U530 (N_530,In_665,In_20);
or U531 (N_531,In_143,In_339);
and U532 (N_532,In_1412,N_453);
xnor U533 (N_533,In_1011,In_267);
or U534 (N_534,In_1434,N_498);
and U535 (N_535,In_696,N_39);
nand U536 (N_536,In_792,In_1401);
nor U537 (N_537,N_447,N_273);
xor U538 (N_538,N_316,In_1494);
nor U539 (N_539,In_457,In_683);
and U540 (N_540,N_45,In_431);
xor U541 (N_541,N_460,N_397);
or U542 (N_542,In_772,In_63);
xnor U543 (N_543,N_458,In_1232);
xor U544 (N_544,N_433,In_137);
xor U545 (N_545,In_168,N_475);
nor U546 (N_546,N_407,In_866);
nor U547 (N_547,N_376,In_1289);
and U548 (N_548,In_605,In_1043);
nand U549 (N_549,In_1073,In_1222);
nand U550 (N_550,N_20,In_832);
nand U551 (N_551,In_747,In_409);
nand U552 (N_552,N_489,In_930);
nand U553 (N_553,N_341,N_436);
nor U554 (N_554,N_102,In_381);
nor U555 (N_555,In_1138,In_611);
nor U556 (N_556,In_111,In_766);
nor U557 (N_557,In_1400,N_361);
xor U558 (N_558,In_1280,N_434);
and U559 (N_559,N_478,In_316);
and U560 (N_560,In_1119,In_897);
and U561 (N_561,N_337,N_240);
xor U562 (N_562,N_105,N_49);
xnor U563 (N_563,N_75,In_308);
or U564 (N_564,In_100,N_206);
nand U565 (N_565,N_281,N_74);
xnor U566 (N_566,N_232,N_444);
and U567 (N_567,In_788,In_790);
nand U568 (N_568,In_399,In_222);
xor U569 (N_569,In_1467,In_499);
or U570 (N_570,N_459,In_125);
or U571 (N_571,In_569,In_1165);
and U572 (N_572,N_409,N_368);
xnor U573 (N_573,In_1466,In_656);
nor U574 (N_574,In_1062,N_420);
or U575 (N_575,N_386,In_1286);
xnor U576 (N_576,In_836,In_84);
xor U577 (N_577,N_303,N_442);
nor U578 (N_578,N_435,In_165);
and U579 (N_579,In_1192,In_193);
or U580 (N_580,In_993,In_302);
or U581 (N_581,In_663,In_817);
nor U582 (N_582,N_399,N_383);
or U583 (N_583,N_499,N_276);
nand U584 (N_584,N_333,N_236);
or U585 (N_585,N_272,N_210);
xor U586 (N_586,In_93,N_224);
and U587 (N_587,In_1139,N_37);
and U588 (N_588,In_638,In_10);
or U589 (N_589,In_1408,In_362);
nor U590 (N_590,In_642,N_95);
and U591 (N_591,N_160,In_729);
and U592 (N_592,N_120,In_450);
or U593 (N_593,In_392,In_280);
and U594 (N_594,In_849,N_490);
or U595 (N_595,In_296,N_167);
xnor U596 (N_596,N_243,In_1181);
or U597 (N_597,In_56,In_372);
and U598 (N_598,In_213,In_738);
and U599 (N_599,N_362,In_1420);
or U600 (N_600,N_113,In_1124);
nor U601 (N_601,In_160,In_735);
nand U602 (N_602,In_1247,In_1303);
nor U603 (N_603,In_1171,In_343);
nor U604 (N_604,In_332,In_1377);
and U605 (N_605,In_969,N_183);
and U606 (N_606,N_124,In_469);
and U607 (N_607,N_439,N_63);
or U608 (N_608,N_401,In_75);
nand U609 (N_609,In_1017,In_384);
xnor U610 (N_610,In_306,N_331);
and U611 (N_611,In_1379,In_901);
and U612 (N_612,N_352,In_74);
and U613 (N_613,In_706,In_884);
and U614 (N_614,In_820,In_1428);
nand U615 (N_615,N_93,In_1264);
nor U616 (N_616,In_1357,In_480);
xnor U617 (N_617,N_450,In_1044);
and U618 (N_618,In_1221,In_307);
or U619 (N_619,N_15,In_1360);
nand U620 (N_620,N_366,N_101);
nor U621 (N_621,In_448,N_338);
xnor U622 (N_622,In_1050,N_340);
xor U623 (N_623,In_616,In_1409);
or U624 (N_624,N_289,In_540);
or U625 (N_625,N_145,In_947);
or U626 (N_626,N_417,N_322);
and U627 (N_627,In_956,In_1184);
nor U628 (N_628,In_623,N_247);
xnor U629 (N_629,N_292,N_78);
nor U630 (N_630,In_632,In_688);
or U631 (N_631,In_1226,In_95);
nor U632 (N_632,In_219,N_271);
xnor U633 (N_633,In_803,In_414);
and U634 (N_634,In_358,N_165);
and U635 (N_635,In_965,In_949);
or U636 (N_636,N_158,In_1149);
nand U637 (N_637,In_797,N_310);
nor U638 (N_638,In_1066,In_563);
or U639 (N_639,In_466,N_394);
nor U640 (N_640,N_492,N_364);
or U641 (N_641,In_488,N_295);
or U642 (N_642,In_723,In_4);
or U643 (N_643,In_629,In_486);
xnor U644 (N_644,N_115,N_200);
nand U645 (N_645,In_1211,N_424);
nand U646 (N_646,In_1129,In_915);
xnor U647 (N_647,In_400,N_67);
nor U648 (N_648,In_699,N_268);
nand U649 (N_649,N_208,In_113);
or U650 (N_650,N_318,N_136);
nor U651 (N_651,N_326,In_771);
nor U652 (N_652,N_220,N_327);
nand U653 (N_653,N_485,N_419);
or U654 (N_654,N_457,N_423);
and U655 (N_655,N_467,In_88);
nand U656 (N_656,N_191,N_12);
nand U657 (N_657,N_430,In_1002);
nand U658 (N_658,In_1417,In_39);
or U659 (N_659,N_235,In_1251);
and U660 (N_660,In_1488,In_1185);
nand U661 (N_661,In_1257,N_455);
xor U662 (N_662,In_600,In_1116);
nor U663 (N_663,N_249,N_42);
or U664 (N_664,In_189,In_557);
and U665 (N_665,In_401,N_471);
xnor U666 (N_666,N_193,In_505);
nand U667 (N_667,N_315,In_449);
or U668 (N_668,N_219,In_1291);
or U669 (N_669,N_252,N_319);
nor U670 (N_670,N_228,In_851);
xnor U671 (N_671,In_1358,In_602);
or U672 (N_672,In_512,N_107);
or U673 (N_673,N_278,In_509);
nand U674 (N_674,In_1451,In_1313);
nand U675 (N_675,In_1190,N_152);
or U676 (N_676,In_1041,In_1093);
or U677 (N_677,In_593,In_1311);
nor U678 (N_678,In_265,In_1367);
xor U679 (N_679,In_397,In_544);
or U680 (N_680,In_808,N_472);
nand U681 (N_681,In_455,N_122);
nor U682 (N_682,In_725,N_413);
nand U683 (N_683,In_933,N_448);
nor U684 (N_684,N_301,In_577);
nand U685 (N_685,In_612,In_174);
nand U686 (N_686,In_246,N_62);
or U687 (N_687,In_974,In_598);
and U688 (N_688,N_400,N_262);
or U689 (N_689,In_526,In_1146);
xnor U690 (N_690,In_1086,In_319);
nand U691 (N_691,In_551,In_33);
nand U692 (N_692,N_494,In_361);
xor U693 (N_693,In_345,In_1406);
or U694 (N_694,In_140,N_30);
nand U695 (N_695,N_282,In_340);
or U696 (N_696,In_405,In_1078);
or U697 (N_697,In_1446,In_553);
or U698 (N_698,In_652,N_189);
and U699 (N_699,In_422,In_1315);
nor U700 (N_700,N_488,N_266);
xnor U701 (N_701,In_237,N_422);
nor U702 (N_702,In_158,In_1072);
nor U703 (N_703,In_1364,N_328);
nand U704 (N_704,In_328,N_40);
nor U705 (N_705,N_142,N_126);
nand U706 (N_706,N_118,In_1144);
and U707 (N_707,In_895,In_49);
or U708 (N_708,In_1186,N_98);
or U709 (N_709,In_503,In_705);
xnor U710 (N_710,N_131,N_402);
or U711 (N_711,In_1415,In_169);
and U712 (N_712,In_478,N_311);
nor U713 (N_713,N_64,In_214);
and U714 (N_714,N_244,In_514);
xnor U715 (N_715,N_144,N_100);
nor U716 (N_716,N_162,In_595);
or U717 (N_717,In_1135,In_959);
nor U718 (N_718,N_370,In_1094);
and U719 (N_719,In_1271,In_1058);
or U720 (N_720,In_1452,In_1198);
xnor U721 (N_721,N_396,N_151);
xor U722 (N_722,In_1039,N_41);
xor U723 (N_723,In_251,In_257);
nor U724 (N_724,In_1445,In_936);
xnor U725 (N_725,In_1120,In_1096);
nor U726 (N_726,In_603,In_1001);
and U727 (N_727,In_1265,In_524);
nand U728 (N_728,In_674,In_426);
or U729 (N_729,N_418,In_684);
nand U730 (N_730,In_501,N_349);
and U731 (N_731,N_440,In_395);
or U732 (N_732,In_1249,In_1449);
nor U733 (N_733,In_942,N_330);
xor U734 (N_734,In_374,In_492);
or U735 (N_735,In_1330,N_141);
and U736 (N_736,In_1013,N_251);
nor U737 (N_737,N_392,N_234);
and U738 (N_738,In_1295,In_264);
or U739 (N_739,In_726,In_789);
and U740 (N_740,N_44,N_325);
nand U741 (N_741,N_1,In_277);
or U742 (N_742,In_767,In_1130);
xnor U743 (N_743,In_436,In_101);
and U744 (N_744,In_500,In_594);
or U745 (N_745,In_247,N_51);
xor U746 (N_746,In_992,In_1231);
nand U747 (N_747,N_385,In_98);
xnor U748 (N_748,N_380,In_79);
and U749 (N_749,In_97,In_483);
nor U750 (N_750,In_775,N_591);
and U751 (N_751,N_648,In_393);
or U752 (N_752,In_1166,N_537);
nor U753 (N_753,N_715,N_94);
nor U754 (N_754,N_543,N_495);
nor U755 (N_755,N_280,In_350);
and U756 (N_756,N_483,In_1225);
nor U757 (N_757,N_110,N_660);
or U758 (N_758,N_226,N_555);
and U759 (N_759,N_545,In_318);
or U760 (N_760,N_553,N_746);
nor U761 (N_761,N_526,N_258);
nand U762 (N_762,In_1207,N_3);
or U763 (N_763,In_984,In_1012);
xor U764 (N_764,In_818,N_733);
nand U765 (N_765,In_1003,N_414);
xor U766 (N_766,N_384,In_804);
or U767 (N_767,In_552,N_293);
and U768 (N_768,In_1268,N_679);
nor U769 (N_769,N_540,N_372);
nand U770 (N_770,In_495,In_1023);
nor U771 (N_771,N_55,In_41);
nand U772 (N_772,In_756,N_441);
or U773 (N_773,N_72,In_558);
and U774 (N_774,In_1145,N_542);
nor U775 (N_775,N_119,N_557);
nand U776 (N_776,N_619,In_1309);
xor U777 (N_777,In_1009,In_1263);
nor U778 (N_778,N_190,N_476);
xor U779 (N_779,N_238,N_354);
and U780 (N_780,N_516,In_886);
nor U781 (N_781,N_639,In_207);
and U782 (N_782,In_346,In_238);
nand U783 (N_783,N_744,N_336);
nor U784 (N_784,N_260,N_556);
nor U785 (N_785,N_718,N_31);
nand U786 (N_786,In_138,In_446);
nor U787 (N_787,In_228,In_758);
or U788 (N_788,In_743,In_1267);
or U789 (N_789,In_1245,N_602);
nor U790 (N_790,N_86,N_194);
nor U791 (N_791,N_48,N_607);
and U792 (N_792,In_1436,In_1294);
nand U793 (N_793,In_59,N_699);
and U794 (N_794,In_172,In_1376);
nor U795 (N_795,N_702,N_332);
nand U796 (N_796,N_515,N_691);
nand U797 (N_797,In_8,In_667);
nand U798 (N_798,N_720,N_672);
xnor U799 (N_799,In_991,In_166);
xnor U800 (N_800,In_692,N_673);
nor U801 (N_801,In_188,N_698);
nor U802 (N_802,In_596,N_406);
or U803 (N_803,N_462,N_692);
xor U804 (N_804,In_1398,N_474);
and U805 (N_805,N_527,N_558);
nor U806 (N_806,In_791,N_645);
xnor U807 (N_807,In_579,In_224);
nand U808 (N_808,In_1158,In_150);
and U809 (N_809,N_456,N_668);
or U810 (N_810,In_753,In_1091);
nor U811 (N_811,N_163,N_508);
nand U812 (N_812,N_371,N_631);
nor U813 (N_813,N_519,N_747);
nand U814 (N_814,In_730,N_487);
or U815 (N_815,N_618,In_1055);
or U816 (N_816,In_571,In_1258);
nor U817 (N_817,In_1422,N_644);
and U818 (N_818,In_1067,N_534);
xnor U819 (N_819,In_198,In_1028);
nand U820 (N_820,N_547,N_308);
or U821 (N_821,N_613,In_1447);
or U822 (N_822,N_703,N_343);
xnor U823 (N_823,In_1163,N_279);
nor U824 (N_824,N_307,N_187);
nand U825 (N_825,N_623,N_321);
or U826 (N_826,In_582,In_1034);
xnor U827 (N_827,In_765,N_657);
nand U828 (N_828,N_314,N_14);
nor U829 (N_829,N_290,N_538);
nand U830 (N_830,In_1290,N_261);
xnor U831 (N_831,N_569,In_87);
nor U832 (N_832,N_530,In_1333);
or U833 (N_833,N_646,In_1273);
or U834 (N_834,In_660,N_632);
xnor U835 (N_835,N_209,In_637);
or U836 (N_836,N_287,N_730);
and U837 (N_837,N_255,N_465);
xnor U838 (N_838,N_347,In_939);
nor U839 (N_839,N_544,In_1368);
xnor U840 (N_840,N_377,N_638);
and U841 (N_841,N_570,In_1274);
nor U842 (N_842,N_614,N_112);
xor U843 (N_843,In_1388,In_893);
nor U844 (N_844,In_239,N_137);
nor U845 (N_845,In_536,N_381);
nor U846 (N_846,In_520,N_653);
nand U847 (N_847,In_823,In_1391);
nand U848 (N_848,In_923,In_1492);
xnor U849 (N_849,N_363,In_43);
nor U850 (N_850,In_1250,N_597);
xor U851 (N_851,N_346,N_53);
and U852 (N_852,In_541,N_317);
xor U853 (N_853,In_1242,N_554);
xnor U854 (N_854,N_393,N_658);
nor U855 (N_855,N_606,N_250);
nor U856 (N_856,N_659,N_46);
nor U857 (N_857,In_19,In_112);
nor U858 (N_858,N_344,N_549);
nor U859 (N_859,N_503,N_582);
xor U860 (N_860,In_694,In_861);
xor U861 (N_861,N_65,N_562);
nor U862 (N_862,N_706,N_520);
nor U863 (N_863,In_304,N_196);
nand U864 (N_864,N_689,In_1324);
and U865 (N_865,In_785,N_550);
nand U866 (N_866,N_621,N_561);
and U867 (N_867,In_545,In_770);
nor U868 (N_868,N_576,In_1407);
or U869 (N_869,N_735,N_714);
and U870 (N_870,N_551,N_506);
and U871 (N_871,N_54,In_1465);
or U872 (N_872,N_2,N_583);
or U873 (N_873,N_500,In_1310);
xnor U874 (N_874,In_1223,N_663);
xor U875 (N_875,N_740,N_36);
or U876 (N_876,N_438,In_859);
nor U877 (N_877,In_1,N_560);
and U878 (N_878,N_701,N_517);
nand U879 (N_879,In_310,N_548);
nor U880 (N_880,N_711,N_599);
nand U881 (N_881,N_681,N_622);
and U882 (N_882,N_509,In_1157);
nand U883 (N_883,N_655,N_265);
or U884 (N_884,In_1425,N_378);
nor U885 (N_885,N_5,N_202);
or U886 (N_886,N_566,N_611);
nand U887 (N_887,In_371,In_899);
or U888 (N_888,In_591,N_357);
nor U889 (N_889,N_214,In_1212);
or U890 (N_890,In_314,In_640);
or U891 (N_891,N_710,N_313);
and U892 (N_892,N_688,N_443);
nor U893 (N_893,N_571,In_795);
nand U894 (N_894,In_1209,In_957);
xor U895 (N_895,N_567,N_595);
nor U896 (N_896,N_27,In_179);
nand U897 (N_897,In_1126,In_1142);
xnor U898 (N_898,N_505,N_486);
nor U899 (N_899,N_429,In_107);
or U900 (N_900,N_33,N_700);
and U901 (N_901,In_879,N_723);
nor U902 (N_902,N_590,N_712);
or U903 (N_903,N_76,N_709);
nor U904 (N_904,In_1031,N_539);
or U905 (N_905,In_233,In_669);
xor U906 (N_906,N_389,In_245);
or U907 (N_907,N_451,In_631);
nor U908 (N_908,N_79,N_320);
nand U909 (N_909,N_298,N_470);
nor U910 (N_910,In_1147,N_4);
nor U911 (N_911,N_552,N_588);
nand U912 (N_912,N_573,In_249);
or U913 (N_913,In_1061,N_408);
nor U914 (N_914,N_670,In_432);
and U915 (N_915,N_225,N_264);
and U916 (N_916,In_439,In_1439);
nor U917 (N_917,N_529,In_989);
or U918 (N_918,N_192,In_124);
xor U919 (N_919,N_564,N_736);
nand U920 (N_920,N_651,In_1419);
nor U921 (N_921,N_513,N_690);
xnor U922 (N_922,In_833,N_727);
or U923 (N_923,N_274,N_512);
nand U924 (N_924,In_1304,N_481);
or U925 (N_925,N_390,N_643);
nand U926 (N_926,N_578,In_515);
nand U927 (N_927,N_630,In_464);
xnor U928 (N_928,N_334,In_71);
nand U929 (N_929,N_463,N_627);
and U930 (N_930,N_367,N_518);
nor U931 (N_931,N_312,In_475);
nor U932 (N_932,N_491,N_696);
or U933 (N_933,N_335,N_257);
xor U934 (N_934,N_395,N_559);
and U935 (N_935,N_375,N_82);
nor U936 (N_936,In_783,In_1054);
nand U937 (N_937,In_273,In_1178);
and U938 (N_938,In_70,In_889);
or U939 (N_939,N_624,N_535);
nand U940 (N_940,In_1168,N_398);
xnor U941 (N_941,In_76,In_530);
nand U942 (N_942,N_687,In_423);
or U943 (N_943,N_104,N_726);
or U944 (N_944,N_286,N_356);
and U945 (N_945,In_378,In_1316);
nor U946 (N_946,N_532,N_647);
xnor U947 (N_947,In_806,In_1484);
or U948 (N_948,In_86,N_521);
or U949 (N_949,N_350,N_195);
nor U950 (N_950,N_739,In_357);
nor U951 (N_951,In_139,N_572);
xnor U952 (N_952,N_596,N_198);
xnor U953 (N_953,N_628,In_812);
or U954 (N_954,N_323,N_204);
xnor U955 (N_955,N_620,N_348);
or U956 (N_956,N_437,N_748);
or U957 (N_957,N_721,N_345);
xor U958 (N_958,In_232,N_605);
xor U959 (N_959,In_200,N_640);
and U960 (N_960,In_1423,N_359);
and U961 (N_961,N_269,N_577);
or U962 (N_962,N_412,In_979);
nor U963 (N_963,In_366,N_52);
and U964 (N_964,In_1077,In_28);
or U965 (N_965,In_234,N_294);
and U966 (N_966,In_16,In_1338);
xnor U967 (N_967,In_869,In_410);
nand U968 (N_968,N_161,N_479);
and U969 (N_969,In_271,N_635);
or U970 (N_970,In_1362,In_133);
or U971 (N_971,N_324,In_333);
or U972 (N_972,In_560,N_734);
and U973 (N_973,N_253,N_729);
nand U974 (N_974,In_1018,In_625);
nor U975 (N_975,In_1060,N_502);
xor U976 (N_976,N_237,N_285);
and U977 (N_977,N_270,N_680);
xor U978 (N_978,N_473,In_1113);
nand U979 (N_979,N_80,In_57);
nor U980 (N_980,In_389,In_1156);
and U981 (N_981,In_1110,N_575);
nor U982 (N_982,N_636,N_387);
and U983 (N_983,N_427,N_677);
or U984 (N_984,N_421,In_121);
and U985 (N_985,N_501,In_760);
nor U986 (N_986,In_996,N_482);
nand U987 (N_987,N_722,N_522);
xor U988 (N_988,In_187,N_694);
and U989 (N_989,In_523,N_665);
and U990 (N_990,N_10,N_480);
nand U991 (N_991,In_1347,N_68);
nand U992 (N_992,N_174,In_506);
or U993 (N_993,N_445,N_342);
or U994 (N_994,In_217,N_682);
nand U995 (N_995,N_256,N_275);
and U996 (N_996,N_634,N_431);
and U997 (N_997,In_914,In_370);
nor U998 (N_998,N_425,In_80);
nand U999 (N_999,In_1053,N_97);
xnor U1000 (N_1000,N_765,N_784);
or U1001 (N_1001,N_750,N_806);
xnor U1002 (N_1002,N_832,In_721);
and U1003 (N_1003,N_824,N_911);
nor U1004 (N_1004,N_525,N_969);
nand U1005 (N_1005,In_690,N_937);
nor U1006 (N_1006,N_675,N_531);
xnor U1007 (N_1007,N_351,N_895);
or U1008 (N_1008,N_819,N_985);
nor U1009 (N_1009,N_123,N_762);
and U1010 (N_1010,N_857,N_865);
xnor U1011 (N_1011,N_683,In_126);
or U1012 (N_1012,N_981,N_885);
and U1013 (N_1013,In_1450,N_523);
or U1014 (N_1014,In_1348,N_626);
nand U1015 (N_1015,In_847,N_305);
and U1016 (N_1016,N_608,N_910);
or U1017 (N_1017,N_892,N_379);
and U1018 (N_1018,N_589,N_813);
xor U1019 (N_1019,N_872,In_1030);
or U1020 (N_1020,N_934,N_943);
and U1021 (N_1021,N_755,N_254);
and U1022 (N_1022,N_907,N_81);
nor U1023 (N_1023,N_609,In_1173);
nor U1024 (N_1024,N_772,N_925);
or U1025 (N_1025,N_822,N_841);
and U1026 (N_1026,N_831,N_881);
or U1027 (N_1027,N_477,N_979);
and U1028 (N_1028,N_996,N_805);
or U1029 (N_1029,N_695,N_994);
or U1030 (N_1030,N_92,N_791);
and U1031 (N_1031,In_575,N_284);
and U1032 (N_1032,N_846,In_496);
or U1033 (N_1033,In_21,N_884);
or U1034 (N_1034,N_373,N_964);
nand U1035 (N_1035,N_941,In_416);
or U1036 (N_1036,N_972,In_248);
xor U1037 (N_1037,In_513,N_829);
and U1038 (N_1038,N_998,In_712);
and U1039 (N_1039,In_1456,N_834);
nand U1040 (N_1040,In_855,N_939);
or U1041 (N_1041,N_811,N_789);
and U1042 (N_1042,N_633,N_957);
nand U1043 (N_1043,N_860,N_708);
nor U1044 (N_1044,N_904,In_592);
nor U1045 (N_1045,In_618,In_840);
nand U1046 (N_1046,N_838,N_732);
xnor U1047 (N_1047,N_365,N_641);
nor U1048 (N_1048,In_982,N_103);
nand U1049 (N_1049,N_890,N_867);
and U1050 (N_1050,N_912,N_771);
xor U1051 (N_1051,N_906,N_942);
nor U1052 (N_1052,N_612,N_752);
nor U1053 (N_1053,N_585,N_891);
nand U1054 (N_1054,N_879,N_587);
nor U1055 (N_1055,N_358,N_411);
nand U1056 (N_1056,In_537,N_992);
xnor U1057 (N_1057,N_932,N_454);
and U1058 (N_1058,In_18,N_642);
and U1059 (N_1059,N_923,N_960);
nand U1060 (N_1060,N_581,N_827);
or U1061 (N_1061,N_795,N_705);
nand U1062 (N_1062,N_963,N_987);
nor U1063 (N_1063,N_83,N_666);
or U1064 (N_1064,N_514,N_432);
xor U1065 (N_1065,N_461,N_958);
or U1066 (N_1066,N_724,N_654);
and U1067 (N_1067,N_404,N_637);
or U1068 (N_1068,N_825,N_304);
xor U1069 (N_1069,In_387,N_719);
nand U1070 (N_1070,N_50,N_751);
or U1071 (N_1071,N_135,In_320);
nand U1072 (N_1072,N_962,N_836);
nor U1073 (N_1073,N_528,In_980);
nor U1074 (N_1074,N_913,N_497);
or U1075 (N_1075,N_649,N_593);
nand U1076 (N_1076,N_603,N_953);
or U1077 (N_1077,N_844,N_667);
xnor U1078 (N_1078,In_1152,N_770);
nor U1079 (N_1079,N_259,N_277);
or U1080 (N_1080,N_355,N_469);
xor U1081 (N_1081,N_815,N_754);
nand U1082 (N_1082,N_742,N_927);
nand U1083 (N_1083,N_650,N_741);
and U1084 (N_1084,In_1435,N_970);
or U1085 (N_1085,N_847,N_896);
or U1086 (N_1086,N_533,N_760);
nand U1087 (N_1087,N_671,N_139);
nand U1088 (N_1088,N_948,N_971);
xor U1089 (N_1089,N_861,N_916);
and U1090 (N_1090,N_968,N_601);
nand U1091 (N_1091,N_656,In_1229);
nand U1092 (N_1092,N_862,N_661);
nand U1093 (N_1093,N_803,N_774);
or U1094 (N_1094,N_835,N_917);
and U1095 (N_1095,N_574,N_792);
nor U1096 (N_1096,N_616,In_2);
nor U1097 (N_1097,N_798,N_933);
and U1098 (N_1098,N_84,N_919);
and U1099 (N_1099,N_339,N_169);
nand U1100 (N_1100,N_615,N_808);
xnor U1101 (N_1101,N_848,N_753);
or U1102 (N_1102,N_403,N_967);
nand U1103 (N_1103,N_511,N_851);
or U1104 (N_1104,N_617,N_875);
or U1105 (N_1105,In_369,N_928);
or U1106 (N_1106,N_973,N_924);
and U1107 (N_1107,In_218,N_850);
xnor U1108 (N_1108,In_119,N_830);
or U1109 (N_1109,N_579,In_1320);
nor U1110 (N_1110,In_1208,N_871);
nand U1111 (N_1111,N_763,N_889);
and U1112 (N_1112,In_282,N_893);
xor U1113 (N_1113,N_563,In_1478);
nand U1114 (N_1114,N_71,N_24);
nor U1115 (N_1115,N_759,N_949);
and U1116 (N_1116,In_998,N_837);
or U1117 (N_1117,N_713,In_1085);
nand U1118 (N_1118,N_776,N_761);
or U1119 (N_1119,N_586,N_267);
or U1120 (N_1120,N_329,N_902);
nor U1121 (N_1121,N_845,N_728);
and U1122 (N_1122,N_507,N_23);
nand U1123 (N_1123,N_984,N_369);
or U1124 (N_1124,N_783,In_662);
xnor U1125 (N_1125,N_817,N_877);
xnor U1126 (N_1126,In_671,N_787);
nand U1127 (N_1127,N_812,N_669);
and U1128 (N_1128,N_864,N_743);
xor U1129 (N_1129,N_674,N_956);
nand U1130 (N_1130,N_678,N_809);
or U1131 (N_1131,In_364,N_955);
and U1132 (N_1132,In_1487,N_797);
and U1133 (N_1133,N_600,N_360);
nor U1134 (N_1134,In_601,In_359);
and U1135 (N_1135,N_415,N_391);
nand U1136 (N_1136,In_532,N_991);
or U1137 (N_1137,In_522,In_131);
nand U1138 (N_1138,N_777,In_268);
nand U1139 (N_1139,N_863,N_428);
and U1140 (N_1140,In_926,N_820);
or U1141 (N_1141,In_311,N_109);
and U1142 (N_1142,N_717,N_779);
and U1143 (N_1143,N_766,N_878);
or U1144 (N_1144,N_565,In_109);
nand U1145 (N_1145,N_737,In_1216);
nor U1146 (N_1146,N_938,N_801);
and U1147 (N_1147,N_704,N_897);
nand U1148 (N_1148,N_914,In_987);
and U1149 (N_1149,N_297,N_888);
or U1150 (N_1150,N_945,N_995);
and U1151 (N_1151,N_977,N_662);
nand U1152 (N_1152,N_947,N_767);
and U1153 (N_1153,N_905,N_946);
nand U1154 (N_1154,N_951,N_676);
and U1155 (N_1155,N_782,N_388);
xnor U1156 (N_1156,N_707,N_839);
or U1157 (N_1157,In_103,N_826);
or U1158 (N_1158,N_944,N_909);
and U1159 (N_1159,N_524,N_980);
nand U1160 (N_1160,N_738,N_222);
or U1161 (N_1161,N_745,In_1404);
and U1162 (N_1162,In_1201,N_853);
nor U1163 (N_1163,N_954,In_713);
or U1164 (N_1164,N_920,In_335);
and U1165 (N_1165,N_799,N_493);
xor U1166 (N_1166,N_887,N_965);
nand U1167 (N_1167,N_309,In_326);
nor U1168 (N_1168,N_868,N_693);
nand U1169 (N_1169,N_291,N_870);
or U1170 (N_1170,N_988,In_1386);
xor U1171 (N_1171,N_686,N_952);
or U1172 (N_1172,N_684,N_921);
nand U1173 (N_1173,N_800,N_592);
nand U1174 (N_1174,In_386,N_899);
nand U1175 (N_1175,In_877,N_449);
and U1176 (N_1176,N_793,N_629);
nand U1177 (N_1177,In_954,N_580);
nand U1178 (N_1178,N_785,N_931);
or U1179 (N_1179,N_731,N_416);
nand U1180 (N_1180,N_898,In_1008);
or U1181 (N_1181,N_858,In_476);
and U1182 (N_1182,N_873,N_426);
nand U1183 (N_1183,N_604,N_978);
xnor U1184 (N_1184,N_903,N_966);
and U1185 (N_1185,N_306,In_937);
nor U1186 (N_1186,In_1378,In_1328);
nor U1187 (N_1187,N_536,N_697);
and U1188 (N_1188,In_784,N_410);
nand U1189 (N_1189,N_816,In_1141);
nand U1190 (N_1190,N_950,N_807);
and U1191 (N_1191,In_85,N_883);
and U1192 (N_1192,N_900,N_852);
nor U1193 (N_1193,In_1180,N_997);
and U1194 (N_1194,N_866,N_959);
or U1195 (N_1195,In_1281,In_835);
or U1196 (N_1196,In_411,N_725);
nand U1197 (N_1197,In_929,N_598);
xor U1198 (N_1198,N_842,N_869);
xnor U1199 (N_1199,N_918,N_769);
or U1200 (N_1200,In_1026,N_986);
nand U1201 (N_1201,N_989,N_802);
nand U1202 (N_1202,N_940,N_843);
nand U1203 (N_1203,In_153,N_961);
or U1204 (N_1204,N_468,N_155);
and U1205 (N_1205,N_790,In_493);
and U1206 (N_1206,In_641,N_856);
nand U1207 (N_1207,N_773,N_300);
and U1208 (N_1208,In_258,N_756);
xnor U1209 (N_1209,N_828,N_936);
nand U1210 (N_1210,N_610,N_685);
and U1211 (N_1211,N_778,N_993);
nor U1212 (N_1212,N_786,N_775);
nand U1213 (N_1213,N_894,N_546);
and U1214 (N_1214,N_758,In_1179);
nor U1215 (N_1215,N_283,N_584);
and U1216 (N_1216,N_859,N_922);
or U1217 (N_1217,In_776,N_664);
or U1218 (N_1218,N_541,N_780);
or U1219 (N_1219,N_882,N_796);
or U1220 (N_1220,N_263,N_886);
nor U1221 (N_1221,N_880,N_990);
nand U1222 (N_1222,N_804,In_882);
nand U1223 (N_1223,N_840,N_821);
or U1224 (N_1224,N_935,N_757);
or U1225 (N_1225,In_142,In_559);
nor U1226 (N_1226,N_908,N_749);
nand U1227 (N_1227,N_181,N_849);
or U1228 (N_1228,In_1174,N_982);
xnor U1229 (N_1229,N_568,N_915);
or U1230 (N_1230,In_898,N_999);
and U1231 (N_1231,N_930,N_974);
nand U1232 (N_1232,N_983,In_388);
xnor U1233 (N_1233,N_975,N_496);
and U1234 (N_1234,In_1270,In_64);
xor U1235 (N_1235,N_781,N_876);
and U1236 (N_1236,N_788,N_874);
and U1237 (N_1237,In_477,N_652);
or U1238 (N_1238,N_764,N_976);
nor U1239 (N_1239,N_854,N_625);
nand U1240 (N_1240,In_988,N_818);
xor U1241 (N_1241,N_901,N_926);
nand U1242 (N_1242,N_504,In_498);
and U1243 (N_1243,N_823,N_855);
nand U1244 (N_1244,N_510,In_990);
and U1245 (N_1245,N_814,N_296);
and U1246 (N_1246,N_716,N_833);
nand U1247 (N_1247,N_768,N_810);
xnor U1248 (N_1248,In_1151,N_794);
nand U1249 (N_1249,N_594,N_929);
xnor U1250 (N_1250,N_1180,N_1067);
nand U1251 (N_1251,N_1043,N_1226);
and U1252 (N_1252,N_1104,N_1166);
and U1253 (N_1253,N_1079,N_1145);
or U1254 (N_1254,N_1186,N_1101);
xor U1255 (N_1255,N_1209,N_1005);
nor U1256 (N_1256,N_1222,N_1068);
nor U1257 (N_1257,N_1134,N_1162);
nand U1258 (N_1258,N_1143,N_1224);
xnor U1259 (N_1259,N_1212,N_1002);
nand U1260 (N_1260,N_1049,N_1015);
or U1261 (N_1261,N_1130,N_1246);
nand U1262 (N_1262,N_1105,N_1241);
nand U1263 (N_1263,N_1201,N_1062);
and U1264 (N_1264,N_1009,N_1050);
nor U1265 (N_1265,N_1030,N_1014);
nor U1266 (N_1266,N_1233,N_1026);
or U1267 (N_1267,N_1041,N_1058);
or U1268 (N_1268,N_1210,N_1206);
nor U1269 (N_1269,N_1012,N_1046);
xnor U1270 (N_1270,N_1150,N_1095);
and U1271 (N_1271,N_1115,N_1245);
xnor U1272 (N_1272,N_1223,N_1184);
nor U1273 (N_1273,N_1194,N_1084);
or U1274 (N_1274,N_1240,N_1003);
or U1275 (N_1275,N_1199,N_1220);
nand U1276 (N_1276,N_1195,N_1020);
and U1277 (N_1277,N_1120,N_1070);
xnor U1278 (N_1278,N_1013,N_1103);
xor U1279 (N_1279,N_1089,N_1042);
or U1280 (N_1280,N_1074,N_1168);
and U1281 (N_1281,N_1221,N_1249);
xor U1282 (N_1282,N_1200,N_1248);
nand U1283 (N_1283,N_1085,N_1019);
and U1284 (N_1284,N_1000,N_1188);
nand U1285 (N_1285,N_1029,N_1088);
and U1286 (N_1286,N_1154,N_1011);
xor U1287 (N_1287,N_1114,N_1169);
and U1288 (N_1288,N_1236,N_1056);
or U1289 (N_1289,N_1028,N_1183);
nand U1290 (N_1290,N_1110,N_1148);
nand U1291 (N_1291,N_1064,N_1207);
and U1292 (N_1292,N_1108,N_1112);
and U1293 (N_1293,N_1087,N_1179);
or U1294 (N_1294,N_1048,N_1229);
nand U1295 (N_1295,N_1117,N_1116);
nor U1296 (N_1296,N_1149,N_1205);
nor U1297 (N_1297,N_1204,N_1165);
xor U1298 (N_1298,N_1021,N_1025);
and U1299 (N_1299,N_1091,N_1096);
nand U1300 (N_1300,N_1007,N_1203);
xor U1301 (N_1301,N_1036,N_1172);
nand U1302 (N_1302,N_1023,N_1109);
xnor U1303 (N_1303,N_1140,N_1044);
nand U1304 (N_1304,N_1001,N_1057);
xnor U1305 (N_1305,N_1202,N_1093);
nor U1306 (N_1306,N_1004,N_1128);
or U1307 (N_1307,N_1040,N_1190);
and U1308 (N_1308,N_1139,N_1059);
xor U1309 (N_1309,N_1135,N_1008);
or U1310 (N_1310,N_1032,N_1211);
and U1311 (N_1311,N_1192,N_1047);
or U1312 (N_1312,N_1144,N_1034);
or U1313 (N_1313,N_1238,N_1124);
or U1314 (N_1314,N_1156,N_1107);
xnor U1315 (N_1315,N_1177,N_1118);
xor U1316 (N_1316,N_1141,N_1176);
or U1317 (N_1317,N_1151,N_1182);
or U1318 (N_1318,N_1173,N_1022);
or U1319 (N_1319,N_1242,N_1217);
nor U1320 (N_1320,N_1076,N_1185);
nand U1321 (N_1321,N_1227,N_1137);
and U1322 (N_1322,N_1051,N_1158);
and U1323 (N_1323,N_1138,N_1247);
or U1324 (N_1324,N_1171,N_1039);
xor U1325 (N_1325,N_1147,N_1216);
and U1326 (N_1326,N_1066,N_1102);
nand U1327 (N_1327,N_1045,N_1098);
nand U1328 (N_1328,N_1146,N_1174);
or U1329 (N_1329,N_1086,N_1031);
or U1330 (N_1330,N_1094,N_1065);
and U1331 (N_1331,N_1080,N_1125);
nor U1332 (N_1332,N_1129,N_1081);
and U1333 (N_1333,N_1092,N_1234);
nand U1334 (N_1334,N_1214,N_1123);
and U1335 (N_1335,N_1127,N_1152);
nand U1336 (N_1336,N_1244,N_1063);
and U1337 (N_1337,N_1213,N_1054);
nor U1338 (N_1338,N_1197,N_1132);
and U1339 (N_1339,N_1016,N_1073);
or U1340 (N_1340,N_1161,N_1061);
or U1341 (N_1341,N_1006,N_1010);
nor U1342 (N_1342,N_1159,N_1090);
xnor U1343 (N_1343,N_1239,N_1133);
or U1344 (N_1344,N_1155,N_1196);
or U1345 (N_1345,N_1017,N_1142);
nor U1346 (N_1346,N_1232,N_1078);
xnor U1347 (N_1347,N_1037,N_1187);
or U1348 (N_1348,N_1157,N_1121);
nor U1349 (N_1349,N_1225,N_1033);
or U1350 (N_1350,N_1122,N_1231);
xnor U1351 (N_1351,N_1027,N_1071);
and U1352 (N_1352,N_1131,N_1055);
xor U1353 (N_1353,N_1136,N_1208);
or U1354 (N_1354,N_1060,N_1072);
nand U1355 (N_1355,N_1193,N_1113);
xor U1356 (N_1356,N_1035,N_1218);
xor U1357 (N_1357,N_1069,N_1215);
or U1358 (N_1358,N_1191,N_1082);
nand U1359 (N_1359,N_1189,N_1100);
nor U1360 (N_1360,N_1243,N_1175);
nand U1361 (N_1361,N_1153,N_1160);
nor U1362 (N_1362,N_1198,N_1024);
nor U1363 (N_1363,N_1038,N_1181);
nand U1364 (N_1364,N_1106,N_1119);
nand U1365 (N_1365,N_1235,N_1167);
and U1366 (N_1366,N_1097,N_1111);
xor U1367 (N_1367,N_1075,N_1018);
nor U1368 (N_1368,N_1219,N_1178);
xor U1369 (N_1369,N_1170,N_1230);
nor U1370 (N_1370,N_1052,N_1126);
xor U1371 (N_1371,N_1077,N_1083);
nor U1372 (N_1372,N_1164,N_1099);
and U1373 (N_1373,N_1237,N_1163);
xnor U1374 (N_1374,N_1053,N_1228);
nand U1375 (N_1375,N_1057,N_1053);
nor U1376 (N_1376,N_1232,N_1249);
or U1377 (N_1377,N_1123,N_1048);
nor U1378 (N_1378,N_1204,N_1076);
nor U1379 (N_1379,N_1085,N_1020);
nand U1380 (N_1380,N_1082,N_1237);
nand U1381 (N_1381,N_1053,N_1060);
nor U1382 (N_1382,N_1162,N_1052);
xor U1383 (N_1383,N_1131,N_1141);
or U1384 (N_1384,N_1170,N_1179);
xnor U1385 (N_1385,N_1069,N_1156);
and U1386 (N_1386,N_1222,N_1143);
xnor U1387 (N_1387,N_1041,N_1188);
nor U1388 (N_1388,N_1013,N_1241);
nand U1389 (N_1389,N_1077,N_1059);
xnor U1390 (N_1390,N_1194,N_1207);
xnor U1391 (N_1391,N_1098,N_1096);
nor U1392 (N_1392,N_1214,N_1121);
and U1393 (N_1393,N_1070,N_1033);
nor U1394 (N_1394,N_1086,N_1027);
nand U1395 (N_1395,N_1091,N_1221);
xor U1396 (N_1396,N_1195,N_1134);
and U1397 (N_1397,N_1196,N_1124);
nand U1398 (N_1398,N_1139,N_1001);
nor U1399 (N_1399,N_1048,N_1016);
nand U1400 (N_1400,N_1066,N_1013);
and U1401 (N_1401,N_1124,N_1208);
or U1402 (N_1402,N_1210,N_1155);
nand U1403 (N_1403,N_1167,N_1138);
nor U1404 (N_1404,N_1094,N_1126);
xor U1405 (N_1405,N_1115,N_1194);
or U1406 (N_1406,N_1039,N_1239);
and U1407 (N_1407,N_1236,N_1034);
and U1408 (N_1408,N_1244,N_1202);
and U1409 (N_1409,N_1182,N_1027);
xnor U1410 (N_1410,N_1053,N_1058);
xor U1411 (N_1411,N_1090,N_1170);
or U1412 (N_1412,N_1166,N_1209);
nor U1413 (N_1413,N_1153,N_1243);
nor U1414 (N_1414,N_1084,N_1090);
xor U1415 (N_1415,N_1218,N_1102);
xor U1416 (N_1416,N_1180,N_1087);
xnor U1417 (N_1417,N_1157,N_1084);
or U1418 (N_1418,N_1075,N_1081);
nand U1419 (N_1419,N_1032,N_1091);
nand U1420 (N_1420,N_1222,N_1247);
nand U1421 (N_1421,N_1245,N_1205);
and U1422 (N_1422,N_1173,N_1044);
nor U1423 (N_1423,N_1236,N_1134);
nand U1424 (N_1424,N_1065,N_1142);
nor U1425 (N_1425,N_1192,N_1118);
xor U1426 (N_1426,N_1031,N_1013);
nor U1427 (N_1427,N_1163,N_1199);
and U1428 (N_1428,N_1067,N_1003);
nand U1429 (N_1429,N_1024,N_1188);
and U1430 (N_1430,N_1069,N_1101);
nor U1431 (N_1431,N_1165,N_1125);
nor U1432 (N_1432,N_1052,N_1063);
xnor U1433 (N_1433,N_1004,N_1209);
nor U1434 (N_1434,N_1235,N_1029);
xnor U1435 (N_1435,N_1032,N_1114);
and U1436 (N_1436,N_1197,N_1136);
or U1437 (N_1437,N_1123,N_1200);
and U1438 (N_1438,N_1112,N_1101);
xor U1439 (N_1439,N_1149,N_1085);
or U1440 (N_1440,N_1078,N_1143);
and U1441 (N_1441,N_1211,N_1044);
nand U1442 (N_1442,N_1244,N_1227);
xnor U1443 (N_1443,N_1206,N_1058);
nor U1444 (N_1444,N_1095,N_1078);
xor U1445 (N_1445,N_1157,N_1166);
and U1446 (N_1446,N_1174,N_1018);
nor U1447 (N_1447,N_1126,N_1020);
and U1448 (N_1448,N_1034,N_1194);
xnor U1449 (N_1449,N_1059,N_1097);
and U1450 (N_1450,N_1113,N_1030);
and U1451 (N_1451,N_1217,N_1188);
and U1452 (N_1452,N_1016,N_1122);
or U1453 (N_1453,N_1160,N_1046);
and U1454 (N_1454,N_1030,N_1007);
or U1455 (N_1455,N_1202,N_1171);
and U1456 (N_1456,N_1096,N_1099);
and U1457 (N_1457,N_1103,N_1206);
nor U1458 (N_1458,N_1124,N_1194);
and U1459 (N_1459,N_1044,N_1075);
nor U1460 (N_1460,N_1213,N_1002);
and U1461 (N_1461,N_1011,N_1028);
and U1462 (N_1462,N_1246,N_1174);
nand U1463 (N_1463,N_1138,N_1073);
xor U1464 (N_1464,N_1249,N_1137);
and U1465 (N_1465,N_1073,N_1002);
nand U1466 (N_1466,N_1210,N_1147);
and U1467 (N_1467,N_1024,N_1155);
or U1468 (N_1468,N_1246,N_1186);
nor U1469 (N_1469,N_1039,N_1104);
or U1470 (N_1470,N_1183,N_1080);
and U1471 (N_1471,N_1240,N_1202);
and U1472 (N_1472,N_1103,N_1204);
and U1473 (N_1473,N_1116,N_1175);
nand U1474 (N_1474,N_1208,N_1031);
or U1475 (N_1475,N_1236,N_1138);
nor U1476 (N_1476,N_1232,N_1153);
and U1477 (N_1477,N_1193,N_1050);
or U1478 (N_1478,N_1009,N_1243);
nor U1479 (N_1479,N_1133,N_1195);
xnor U1480 (N_1480,N_1045,N_1068);
xnor U1481 (N_1481,N_1067,N_1100);
and U1482 (N_1482,N_1206,N_1234);
and U1483 (N_1483,N_1093,N_1221);
and U1484 (N_1484,N_1066,N_1110);
or U1485 (N_1485,N_1151,N_1244);
xor U1486 (N_1486,N_1210,N_1094);
or U1487 (N_1487,N_1105,N_1217);
nor U1488 (N_1488,N_1133,N_1080);
nor U1489 (N_1489,N_1216,N_1166);
xor U1490 (N_1490,N_1237,N_1060);
nand U1491 (N_1491,N_1140,N_1092);
xor U1492 (N_1492,N_1181,N_1119);
and U1493 (N_1493,N_1125,N_1137);
nor U1494 (N_1494,N_1039,N_1228);
and U1495 (N_1495,N_1164,N_1200);
and U1496 (N_1496,N_1144,N_1163);
xor U1497 (N_1497,N_1076,N_1231);
xor U1498 (N_1498,N_1003,N_1013);
and U1499 (N_1499,N_1068,N_1149);
and U1500 (N_1500,N_1490,N_1411);
nand U1501 (N_1501,N_1251,N_1334);
and U1502 (N_1502,N_1297,N_1273);
nor U1503 (N_1503,N_1495,N_1401);
nor U1504 (N_1504,N_1397,N_1396);
nor U1505 (N_1505,N_1498,N_1314);
nor U1506 (N_1506,N_1461,N_1329);
and U1507 (N_1507,N_1446,N_1370);
nand U1508 (N_1508,N_1294,N_1373);
nand U1509 (N_1509,N_1315,N_1316);
nand U1510 (N_1510,N_1386,N_1318);
nand U1511 (N_1511,N_1345,N_1288);
xor U1512 (N_1512,N_1346,N_1476);
and U1513 (N_1513,N_1387,N_1298);
or U1514 (N_1514,N_1257,N_1264);
or U1515 (N_1515,N_1357,N_1431);
nor U1516 (N_1516,N_1354,N_1458);
nand U1517 (N_1517,N_1343,N_1259);
and U1518 (N_1518,N_1389,N_1465);
or U1519 (N_1519,N_1301,N_1252);
or U1520 (N_1520,N_1390,N_1300);
nand U1521 (N_1521,N_1361,N_1489);
nand U1522 (N_1522,N_1494,N_1413);
and U1523 (N_1523,N_1444,N_1284);
xnor U1524 (N_1524,N_1393,N_1380);
or U1525 (N_1525,N_1378,N_1462);
nand U1526 (N_1526,N_1466,N_1423);
nand U1527 (N_1527,N_1291,N_1254);
nor U1528 (N_1528,N_1414,N_1341);
and U1529 (N_1529,N_1456,N_1270);
and U1530 (N_1530,N_1473,N_1302);
or U1531 (N_1531,N_1303,N_1325);
and U1532 (N_1532,N_1438,N_1313);
nor U1533 (N_1533,N_1289,N_1364);
nor U1534 (N_1534,N_1372,N_1321);
and U1535 (N_1535,N_1497,N_1385);
and U1536 (N_1536,N_1355,N_1381);
xor U1537 (N_1537,N_1406,N_1488);
nor U1538 (N_1538,N_1342,N_1290);
nor U1539 (N_1539,N_1317,N_1368);
and U1540 (N_1540,N_1356,N_1307);
and U1541 (N_1541,N_1336,N_1293);
nor U1542 (N_1542,N_1344,N_1425);
nor U1543 (N_1543,N_1402,N_1337);
and U1544 (N_1544,N_1482,N_1319);
nand U1545 (N_1545,N_1295,N_1268);
nor U1546 (N_1546,N_1282,N_1353);
nand U1547 (N_1547,N_1398,N_1256);
and U1548 (N_1548,N_1374,N_1296);
and U1549 (N_1549,N_1471,N_1440);
or U1550 (N_1550,N_1258,N_1312);
and U1551 (N_1551,N_1333,N_1349);
nor U1552 (N_1552,N_1475,N_1347);
or U1553 (N_1553,N_1299,N_1340);
nand U1554 (N_1554,N_1272,N_1308);
and U1555 (N_1555,N_1429,N_1277);
nand U1556 (N_1556,N_1285,N_1279);
xor U1557 (N_1557,N_1365,N_1304);
or U1558 (N_1558,N_1427,N_1492);
and U1559 (N_1559,N_1455,N_1428);
or U1560 (N_1560,N_1348,N_1384);
and U1561 (N_1561,N_1460,N_1306);
nand U1562 (N_1562,N_1405,N_1369);
or U1563 (N_1563,N_1328,N_1474);
xnor U1564 (N_1564,N_1468,N_1453);
and U1565 (N_1565,N_1448,N_1278);
xnor U1566 (N_1566,N_1292,N_1382);
xor U1567 (N_1567,N_1375,N_1480);
xor U1568 (N_1568,N_1266,N_1358);
nand U1569 (N_1569,N_1371,N_1260);
nor U1570 (N_1570,N_1323,N_1324);
nor U1571 (N_1571,N_1379,N_1250);
or U1572 (N_1572,N_1267,N_1280);
nor U1573 (N_1573,N_1470,N_1437);
nor U1574 (N_1574,N_1441,N_1286);
xnor U1575 (N_1575,N_1322,N_1335);
or U1576 (N_1576,N_1399,N_1477);
nor U1577 (N_1577,N_1434,N_1499);
or U1578 (N_1578,N_1276,N_1443);
or U1579 (N_1579,N_1362,N_1388);
nand U1580 (N_1580,N_1392,N_1281);
nor U1581 (N_1581,N_1309,N_1450);
and U1582 (N_1582,N_1481,N_1404);
nand U1583 (N_1583,N_1261,N_1487);
or U1584 (N_1584,N_1424,N_1452);
or U1585 (N_1585,N_1436,N_1269);
nor U1586 (N_1586,N_1496,N_1383);
nor U1587 (N_1587,N_1472,N_1491);
nand U1588 (N_1588,N_1310,N_1320);
and U1589 (N_1589,N_1447,N_1339);
or U1590 (N_1590,N_1463,N_1366);
and U1591 (N_1591,N_1422,N_1426);
and U1592 (N_1592,N_1479,N_1412);
and U1593 (N_1593,N_1400,N_1262);
or U1594 (N_1594,N_1360,N_1271);
and U1595 (N_1595,N_1416,N_1459);
or U1596 (N_1596,N_1338,N_1408);
nand U1597 (N_1597,N_1421,N_1255);
or U1598 (N_1598,N_1351,N_1352);
or U1599 (N_1599,N_1377,N_1457);
and U1600 (N_1600,N_1432,N_1430);
or U1601 (N_1601,N_1449,N_1311);
xnor U1602 (N_1602,N_1410,N_1403);
xnor U1603 (N_1603,N_1332,N_1417);
or U1604 (N_1604,N_1305,N_1420);
and U1605 (N_1605,N_1326,N_1376);
xnor U1606 (N_1606,N_1435,N_1274);
nor U1607 (N_1607,N_1469,N_1439);
nand U1608 (N_1608,N_1483,N_1415);
and U1609 (N_1609,N_1451,N_1485);
and U1610 (N_1610,N_1265,N_1283);
and U1611 (N_1611,N_1331,N_1493);
or U1612 (N_1612,N_1433,N_1367);
xor U1613 (N_1613,N_1442,N_1486);
nor U1614 (N_1614,N_1407,N_1467);
and U1615 (N_1615,N_1454,N_1395);
xnor U1616 (N_1616,N_1478,N_1287);
and U1617 (N_1617,N_1391,N_1253);
nor U1618 (N_1618,N_1327,N_1418);
nand U1619 (N_1619,N_1363,N_1394);
nor U1620 (N_1620,N_1330,N_1484);
or U1621 (N_1621,N_1359,N_1263);
xor U1622 (N_1622,N_1464,N_1350);
xnor U1623 (N_1623,N_1445,N_1275);
or U1624 (N_1624,N_1419,N_1409);
nand U1625 (N_1625,N_1477,N_1255);
nand U1626 (N_1626,N_1258,N_1417);
xnor U1627 (N_1627,N_1334,N_1365);
or U1628 (N_1628,N_1400,N_1380);
nand U1629 (N_1629,N_1331,N_1358);
or U1630 (N_1630,N_1349,N_1486);
and U1631 (N_1631,N_1433,N_1464);
xnor U1632 (N_1632,N_1265,N_1391);
xnor U1633 (N_1633,N_1259,N_1460);
nand U1634 (N_1634,N_1405,N_1282);
and U1635 (N_1635,N_1428,N_1389);
or U1636 (N_1636,N_1269,N_1273);
or U1637 (N_1637,N_1327,N_1473);
and U1638 (N_1638,N_1371,N_1366);
and U1639 (N_1639,N_1433,N_1310);
or U1640 (N_1640,N_1488,N_1318);
or U1641 (N_1641,N_1351,N_1416);
nand U1642 (N_1642,N_1374,N_1329);
and U1643 (N_1643,N_1467,N_1489);
nor U1644 (N_1644,N_1347,N_1352);
xnor U1645 (N_1645,N_1314,N_1335);
or U1646 (N_1646,N_1312,N_1346);
nor U1647 (N_1647,N_1329,N_1457);
xor U1648 (N_1648,N_1390,N_1326);
nand U1649 (N_1649,N_1360,N_1384);
and U1650 (N_1650,N_1398,N_1254);
xnor U1651 (N_1651,N_1326,N_1488);
or U1652 (N_1652,N_1441,N_1321);
nor U1653 (N_1653,N_1393,N_1367);
nor U1654 (N_1654,N_1307,N_1300);
nand U1655 (N_1655,N_1457,N_1282);
or U1656 (N_1656,N_1267,N_1458);
xnor U1657 (N_1657,N_1291,N_1487);
nor U1658 (N_1658,N_1421,N_1479);
xnor U1659 (N_1659,N_1402,N_1414);
and U1660 (N_1660,N_1365,N_1448);
or U1661 (N_1661,N_1309,N_1289);
nor U1662 (N_1662,N_1342,N_1409);
nor U1663 (N_1663,N_1312,N_1482);
and U1664 (N_1664,N_1422,N_1270);
and U1665 (N_1665,N_1269,N_1381);
nand U1666 (N_1666,N_1485,N_1491);
and U1667 (N_1667,N_1492,N_1384);
and U1668 (N_1668,N_1252,N_1397);
xor U1669 (N_1669,N_1499,N_1257);
nor U1670 (N_1670,N_1338,N_1491);
nor U1671 (N_1671,N_1488,N_1301);
nor U1672 (N_1672,N_1303,N_1472);
or U1673 (N_1673,N_1434,N_1323);
nand U1674 (N_1674,N_1276,N_1369);
and U1675 (N_1675,N_1341,N_1450);
or U1676 (N_1676,N_1460,N_1365);
and U1677 (N_1677,N_1422,N_1370);
nor U1678 (N_1678,N_1399,N_1384);
nand U1679 (N_1679,N_1290,N_1478);
or U1680 (N_1680,N_1280,N_1401);
xnor U1681 (N_1681,N_1292,N_1327);
and U1682 (N_1682,N_1337,N_1341);
xor U1683 (N_1683,N_1260,N_1404);
and U1684 (N_1684,N_1366,N_1294);
nand U1685 (N_1685,N_1274,N_1437);
and U1686 (N_1686,N_1442,N_1401);
nand U1687 (N_1687,N_1358,N_1318);
and U1688 (N_1688,N_1497,N_1419);
nand U1689 (N_1689,N_1316,N_1417);
nand U1690 (N_1690,N_1384,N_1300);
or U1691 (N_1691,N_1371,N_1421);
nand U1692 (N_1692,N_1487,N_1256);
nor U1693 (N_1693,N_1277,N_1439);
nand U1694 (N_1694,N_1307,N_1442);
or U1695 (N_1695,N_1426,N_1450);
or U1696 (N_1696,N_1267,N_1290);
nand U1697 (N_1697,N_1362,N_1376);
nand U1698 (N_1698,N_1388,N_1307);
nor U1699 (N_1699,N_1378,N_1353);
nand U1700 (N_1700,N_1261,N_1269);
nand U1701 (N_1701,N_1333,N_1411);
or U1702 (N_1702,N_1426,N_1307);
nand U1703 (N_1703,N_1464,N_1254);
nor U1704 (N_1704,N_1382,N_1475);
nor U1705 (N_1705,N_1412,N_1387);
or U1706 (N_1706,N_1435,N_1411);
xor U1707 (N_1707,N_1474,N_1400);
and U1708 (N_1708,N_1299,N_1313);
nor U1709 (N_1709,N_1250,N_1494);
nor U1710 (N_1710,N_1474,N_1457);
or U1711 (N_1711,N_1466,N_1346);
nand U1712 (N_1712,N_1425,N_1481);
nand U1713 (N_1713,N_1478,N_1304);
nand U1714 (N_1714,N_1484,N_1388);
or U1715 (N_1715,N_1340,N_1254);
nand U1716 (N_1716,N_1360,N_1399);
or U1717 (N_1717,N_1285,N_1405);
xnor U1718 (N_1718,N_1407,N_1481);
and U1719 (N_1719,N_1279,N_1491);
or U1720 (N_1720,N_1280,N_1494);
or U1721 (N_1721,N_1311,N_1358);
xor U1722 (N_1722,N_1405,N_1375);
or U1723 (N_1723,N_1398,N_1267);
nor U1724 (N_1724,N_1329,N_1273);
xor U1725 (N_1725,N_1344,N_1412);
or U1726 (N_1726,N_1299,N_1413);
and U1727 (N_1727,N_1275,N_1456);
nand U1728 (N_1728,N_1417,N_1263);
nor U1729 (N_1729,N_1493,N_1475);
or U1730 (N_1730,N_1325,N_1343);
nand U1731 (N_1731,N_1396,N_1366);
nand U1732 (N_1732,N_1450,N_1313);
nand U1733 (N_1733,N_1412,N_1410);
xnor U1734 (N_1734,N_1356,N_1278);
xor U1735 (N_1735,N_1469,N_1255);
or U1736 (N_1736,N_1491,N_1460);
xnor U1737 (N_1737,N_1362,N_1451);
or U1738 (N_1738,N_1369,N_1385);
or U1739 (N_1739,N_1374,N_1262);
or U1740 (N_1740,N_1387,N_1325);
and U1741 (N_1741,N_1494,N_1256);
nand U1742 (N_1742,N_1452,N_1363);
nor U1743 (N_1743,N_1438,N_1306);
nand U1744 (N_1744,N_1280,N_1333);
or U1745 (N_1745,N_1453,N_1267);
or U1746 (N_1746,N_1412,N_1458);
or U1747 (N_1747,N_1490,N_1413);
and U1748 (N_1748,N_1497,N_1302);
nor U1749 (N_1749,N_1385,N_1303);
nand U1750 (N_1750,N_1581,N_1536);
or U1751 (N_1751,N_1597,N_1671);
or U1752 (N_1752,N_1534,N_1670);
nor U1753 (N_1753,N_1619,N_1524);
or U1754 (N_1754,N_1562,N_1656);
nor U1755 (N_1755,N_1724,N_1566);
nand U1756 (N_1756,N_1526,N_1653);
nor U1757 (N_1757,N_1690,N_1647);
nor U1758 (N_1758,N_1626,N_1677);
nor U1759 (N_1759,N_1665,N_1510);
nand U1760 (N_1760,N_1684,N_1732);
and U1761 (N_1761,N_1564,N_1598);
nand U1762 (N_1762,N_1682,N_1596);
or U1763 (N_1763,N_1603,N_1655);
xor U1764 (N_1764,N_1539,N_1700);
or U1765 (N_1765,N_1629,N_1585);
nor U1766 (N_1766,N_1680,N_1576);
xnor U1767 (N_1767,N_1645,N_1636);
or U1768 (N_1768,N_1569,N_1711);
and U1769 (N_1769,N_1516,N_1698);
nand U1770 (N_1770,N_1742,N_1702);
nand U1771 (N_1771,N_1533,N_1587);
or U1772 (N_1772,N_1568,N_1554);
and U1773 (N_1773,N_1578,N_1520);
nor U1774 (N_1774,N_1641,N_1550);
nor U1775 (N_1775,N_1588,N_1628);
xnor U1776 (N_1776,N_1639,N_1509);
xnor U1777 (N_1777,N_1584,N_1730);
nor U1778 (N_1778,N_1624,N_1693);
nand U1779 (N_1779,N_1747,N_1609);
xnor U1780 (N_1780,N_1685,N_1560);
or U1781 (N_1781,N_1540,N_1630);
xor U1782 (N_1782,N_1608,N_1625);
nor U1783 (N_1783,N_1664,N_1661);
nor U1784 (N_1784,N_1638,N_1692);
nand U1785 (N_1785,N_1527,N_1604);
nand U1786 (N_1786,N_1716,N_1743);
or U1787 (N_1787,N_1521,N_1707);
nor U1788 (N_1788,N_1574,N_1513);
nand U1789 (N_1789,N_1740,N_1676);
or U1790 (N_1790,N_1531,N_1659);
or U1791 (N_1791,N_1544,N_1662);
or U1792 (N_1792,N_1719,N_1508);
xnor U1793 (N_1793,N_1652,N_1731);
nor U1794 (N_1794,N_1723,N_1557);
nor U1795 (N_1795,N_1642,N_1696);
and U1796 (N_1796,N_1709,N_1612);
or U1797 (N_1797,N_1607,N_1591);
nand U1798 (N_1798,N_1669,N_1646);
or U1799 (N_1799,N_1571,N_1699);
nor U1800 (N_1800,N_1737,N_1717);
xor U1801 (N_1801,N_1749,N_1725);
and U1802 (N_1802,N_1617,N_1522);
nor U1803 (N_1803,N_1722,N_1697);
nor U1804 (N_1804,N_1673,N_1552);
xnor U1805 (N_1805,N_1570,N_1573);
or U1806 (N_1806,N_1691,N_1715);
or U1807 (N_1807,N_1729,N_1643);
and U1808 (N_1808,N_1586,N_1710);
nor U1809 (N_1809,N_1601,N_1728);
nand U1810 (N_1810,N_1721,N_1736);
nor U1811 (N_1811,N_1618,N_1713);
nor U1812 (N_1812,N_1518,N_1529);
or U1813 (N_1813,N_1541,N_1735);
xor U1814 (N_1814,N_1590,N_1651);
or U1815 (N_1815,N_1551,N_1650);
nand U1816 (N_1816,N_1741,N_1592);
xor U1817 (N_1817,N_1549,N_1720);
or U1818 (N_1818,N_1565,N_1575);
nor U1819 (N_1819,N_1595,N_1616);
nand U1820 (N_1820,N_1632,N_1627);
xor U1821 (N_1821,N_1678,N_1610);
or U1822 (N_1822,N_1503,N_1558);
and U1823 (N_1823,N_1714,N_1640);
and U1824 (N_1824,N_1660,N_1688);
or U1825 (N_1825,N_1648,N_1532);
and U1826 (N_1826,N_1745,N_1502);
or U1827 (N_1827,N_1704,N_1599);
nand U1828 (N_1828,N_1602,N_1613);
or U1829 (N_1829,N_1580,N_1667);
nand U1830 (N_1830,N_1583,N_1695);
nor U1831 (N_1831,N_1621,N_1579);
xnor U1832 (N_1832,N_1738,N_1548);
xnor U1833 (N_1833,N_1706,N_1528);
nor U1834 (N_1834,N_1572,N_1589);
or U1835 (N_1835,N_1537,N_1663);
nor U1836 (N_1836,N_1683,N_1734);
nand U1837 (N_1837,N_1681,N_1654);
nor U1838 (N_1838,N_1644,N_1594);
and U1839 (N_1839,N_1559,N_1507);
nand U1840 (N_1840,N_1567,N_1600);
or U1841 (N_1841,N_1582,N_1556);
or U1842 (N_1842,N_1686,N_1744);
or U1843 (N_1843,N_1514,N_1666);
nor U1844 (N_1844,N_1615,N_1674);
and U1845 (N_1845,N_1623,N_1675);
nor U1846 (N_1846,N_1635,N_1525);
or U1847 (N_1847,N_1542,N_1733);
xor U1848 (N_1848,N_1506,N_1689);
nor U1849 (N_1849,N_1593,N_1555);
and U1850 (N_1850,N_1546,N_1519);
or U1851 (N_1851,N_1672,N_1748);
or U1852 (N_1852,N_1511,N_1605);
nor U1853 (N_1853,N_1543,N_1614);
xor U1854 (N_1854,N_1739,N_1708);
or U1855 (N_1855,N_1703,N_1535);
nand U1856 (N_1856,N_1658,N_1545);
or U1857 (N_1857,N_1718,N_1668);
and U1858 (N_1858,N_1712,N_1727);
or U1859 (N_1859,N_1634,N_1746);
or U1860 (N_1860,N_1501,N_1606);
or U1861 (N_1861,N_1517,N_1553);
xor U1862 (N_1862,N_1500,N_1657);
nand U1863 (N_1863,N_1530,N_1547);
xnor U1864 (N_1864,N_1633,N_1512);
xor U1865 (N_1865,N_1561,N_1705);
or U1866 (N_1866,N_1701,N_1563);
nor U1867 (N_1867,N_1622,N_1649);
xnor U1868 (N_1868,N_1505,N_1687);
or U1869 (N_1869,N_1694,N_1523);
or U1870 (N_1870,N_1538,N_1726);
and U1871 (N_1871,N_1577,N_1637);
or U1872 (N_1872,N_1679,N_1620);
nand U1873 (N_1873,N_1515,N_1631);
nand U1874 (N_1874,N_1611,N_1504);
nand U1875 (N_1875,N_1625,N_1585);
and U1876 (N_1876,N_1607,N_1730);
xor U1877 (N_1877,N_1648,N_1604);
nand U1878 (N_1878,N_1623,N_1641);
nor U1879 (N_1879,N_1716,N_1631);
or U1880 (N_1880,N_1722,N_1666);
nand U1881 (N_1881,N_1573,N_1563);
and U1882 (N_1882,N_1676,N_1725);
nand U1883 (N_1883,N_1627,N_1607);
nand U1884 (N_1884,N_1575,N_1554);
nand U1885 (N_1885,N_1690,N_1619);
nor U1886 (N_1886,N_1697,N_1745);
or U1887 (N_1887,N_1721,N_1567);
xnor U1888 (N_1888,N_1568,N_1524);
xor U1889 (N_1889,N_1630,N_1533);
nor U1890 (N_1890,N_1614,N_1620);
or U1891 (N_1891,N_1558,N_1746);
nand U1892 (N_1892,N_1710,N_1726);
and U1893 (N_1893,N_1535,N_1534);
nand U1894 (N_1894,N_1747,N_1690);
nor U1895 (N_1895,N_1562,N_1569);
xnor U1896 (N_1896,N_1658,N_1690);
xor U1897 (N_1897,N_1539,N_1651);
nand U1898 (N_1898,N_1502,N_1533);
or U1899 (N_1899,N_1678,N_1530);
and U1900 (N_1900,N_1512,N_1698);
or U1901 (N_1901,N_1525,N_1706);
or U1902 (N_1902,N_1704,N_1542);
nand U1903 (N_1903,N_1582,N_1735);
and U1904 (N_1904,N_1632,N_1503);
nand U1905 (N_1905,N_1611,N_1712);
or U1906 (N_1906,N_1508,N_1749);
nor U1907 (N_1907,N_1711,N_1578);
nor U1908 (N_1908,N_1521,N_1645);
nor U1909 (N_1909,N_1723,N_1541);
and U1910 (N_1910,N_1734,N_1568);
and U1911 (N_1911,N_1616,N_1606);
and U1912 (N_1912,N_1698,N_1660);
or U1913 (N_1913,N_1723,N_1602);
or U1914 (N_1914,N_1733,N_1617);
nor U1915 (N_1915,N_1546,N_1659);
nand U1916 (N_1916,N_1501,N_1621);
nor U1917 (N_1917,N_1543,N_1719);
xor U1918 (N_1918,N_1741,N_1609);
or U1919 (N_1919,N_1532,N_1674);
nand U1920 (N_1920,N_1707,N_1604);
and U1921 (N_1921,N_1657,N_1565);
and U1922 (N_1922,N_1591,N_1718);
nor U1923 (N_1923,N_1585,N_1690);
nand U1924 (N_1924,N_1708,N_1730);
nand U1925 (N_1925,N_1693,N_1626);
nand U1926 (N_1926,N_1590,N_1707);
and U1927 (N_1927,N_1744,N_1674);
and U1928 (N_1928,N_1555,N_1724);
nand U1929 (N_1929,N_1734,N_1710);
nand U1930 (N_1930,N_1560,N_1606);
xor U1931 (N_1931,N_1713,N_1679);
or U1932 (N_1932,N_1609,N_1589);
xor U1933 (N_1933,N_1549,N_1676);
nor U1934 (N_1934,N_1609,N_1626);
or U1935 (N_1935,N_1507,N_1632);
or U1936 (N_1936,N_1519,N_1670);
and U1937 (N_1937,N_1634,N_1726);
nor U1938 (N_1938,N_1735,N_1574);
and U1939 (N_1939,N_1605,N_1607);
nand U1940 (N_1940,N_1739,N_1631);
xor U1941 (N_1941,N_1585,N_1511);
xor U1942 (N_1942,N_1721,N_1554);
or U1943 (N_1943,N_1568,N_1669);
nand U1944 (N_1944,N_1725,N_1572);
xor U1945 (N_1945,N_1646,N_1502);
nor U1946 (N_1946,N_1518,N_1641);
and U1947 (N_1947,N_1542,N_1656);
and U1948 (N_1948,N_1551,N_1547);
nor U1949 (N_1949,N_1660,N_1663);
nand U1950 (N_1950,N_1702,N_1684);
nor U1951 (N_1951,N_1746,N_1544);
or U1952 (N_1952,N_1575,N_1727);
nor U1953 (N_1953,N_1589,N_1583);
and U1954 (N_1954,N_1500,N_1542);
or U1955 (N_1955,N_1608,N_1586);
nor U1956 (N_1956,N_1530,N_1622);
or U1957 (N_1957,N_1660,N_1608);
nor U1958 (N_1958,N_1702,N_1671);
and U1959 (N_1959,N_1542,N_1560);
and U1960 (N_1960,N_1732,N_1585);
xnor U1961 (N_1961,N_1642,N_1511);
nand U1962 (N_1962,N_1744,N_1709);
or U1963 (N_1963,N_1638,N_1599);
xnor U1964 (N_1964,N_1576,N_1503);
xor U1965 (N_1965,N_1612,N_1613);
xor U1966 (N_1966,N_1693,N_1602);
xor U1967 (N_1967,N_1529,N_1710);
nor U1968 (N_1968,N_1568,N_1732);
nor U1969 (N_1969,N_1630,N_1605);
nor U1970 (N_1970,N_1607,N_1524);
or U1971 (N_1971,N_1667,N_1724);
nor U1972 (N_1972,N_1626,N_1509);
or U1973 (N_1973,N_1604,N_1724);
and U1974 (N_1974,N_1720,N_1647);
xor U1975 (N_1975,N_1627,N_1521);
and U1976 (N_1976,N_1617,N_1749);
nand U1977 (N_1977,N_1613,N_1533);
and U1978 (N_1978,N_1512,N_1654);
nor U1979 (N_1979,N_1534,N_1548);
xnor U1980 (N_1980,N_1575,N_1690);
xor U1981 (N_1981,N_1526,N_1588);
xor U1982 (N_1982,N_1694,N_1576);
nand U1983 (N_1983,N_1657,N_1530);
xnor U1984 (N_1984,N_1548,N_1551);
xnor U1985 (N_1985,N_1588,N_1738);
or U1986 (N_1986,N_1542,N_1623);
xor U1987 (N_1987,N_1608,N_1641);
and U1988 (N_1988,N_1545,N_1503);
and U1989 (N_1989,N_1601,N_1707);
nand U1990 (N_1990,N_1614,N_1687);
and U1991 (N_1991,N_1643,N_1672);
and U1992 (N_1992,N_1613,N_1521);
or U1993 (N_1993,N_1738,N_1733);
nor U1994 (N_1994,N_1700,N_1699);
or U1995 (N_1995,N_1522,N_1710);
nor U1996 (N_1996,N_1720,N_1718);
nor U1997 (N_1997,N_1724,N_1616);
nand U1998 (N_1998,N_1636,N_1623);
and U1999 (N_1999,N_1709,N_1697);
nor U2000 (N_2000,N_1927,N_1771);
xor U2001 (N_2001,N_1946,N_1956);
or U2002 (N_2002,N_1859,N_1849);
xnor U2003 (N_2003,N_1963,N_1841);
and U2004 (N_2004,N_1881,N_1842);
nand U2005 (N_2005,N_1924,N_1777);
nand U2006 (N_2006,N_1900,N_1853);
and U2007 (N_2007,N_1840,N_1988);
nand U2008 (N_2008,N_1913,N_1949);
nand U2009 (N_2009,N_1957,N_1827);
xor U2010 (N_2010,N_1871,N_1984);
and U2011 (N_2011,N_1939,N_1756);
xnor U2012 (N_2012,N_1981,N_1903);
or U2013 (N_2013,N_1834,N_1790);
and U2014 (N_2014,N_1891,N_1921);
xor U2015 (N_2015,N_1966,N_1964);
and U2016 (N_2016,N_1815,N_1996);
nand U2017 (N_2017,N_1839,N_1794);
and U2018 (N_2018,N_1967,N_1935);
or U2019 (N_2019,N_1951,N_1819);
xnor U2020 (N_2020,N_1847,N_1772);
xnor U2021 (N_2021,N_1888,N_1800);
nor U2022 (N_2022,N_1923,N_1974);
and U2023 (N_2023,N_1803,N_1764);
nor U2024 (N_2024,N_1979,N_1797);
and U2025 (N_2025,N_1953,N_1767);
nand U2026 (N_2026,N_1813,N_1829);
nand U2027 (N_2027,N_1962,N_1879);
xnor U2028 (N_2028,N_1992,N_1798);
and U2029 (N_2029,N_1865,N_1959);
nand U2030 (N_2030,N_1808,N_1750);
and U2031 (N_2031,N_1997,N_1761);
nor U2032 (N_2032,N_1751,N_1862);
xor U2033 (N_2033,N_1778,N_1878);
and U2034 (N_2034,N_1788,N_1826);
nor U2035 (N_2035,N_1940,N_1932);
nor U2036 (N_2036,N_1978,N_1844);
nor U2037 (N_2037,N_1854,N_1817);
xnor U2038 (N_2038,N_1783,N_1898);
and U2039 (N_2039,N_1763,N_1926);
xnor U2040 (N_2040,N_1933,N_1948);
nand U2041 (N_2041,N_1848,N_1782);
xor U2042 (N_2042,N_1781,N_1931);
and U2043 (N_2043,N_1902,N_1983);
nor U2044 (N_2044,N_1875,N_1780);
nand U2045 (N_2045,N_1768,N_1961);
xnor U2046 (N_2046,N_1912,N_1954);
and U2047 (N_2047,N_1887,N_1754);
and U2048 (N_2048,N_1928,N_1773);
xor U2049 (N_2049,N_1874,N_1977);
and U2050 (N_2050,N_1972,N_1904);
and U2051 (N_2051,N_1799,N_1910);
and U2052 (N_2052,N_1989,N_1938);
or U2053 (N_2053,N_1925,N_1828);
nand U2054 (N_2054,N_1918,N_1911);
xnor U2055 (N_2055,N_1762,N_1973);
or U2056 (N_2056,N_1994,N_1876);
nand U2057 (N_2057,N_1870,N_1811);
and U2058 (N_2058,N_1917,N_1814);
xnor U2059 (N_2059,N_1864,N_1915);
nor U2060 (N_2060,N_1892,N_1944);
and U2061 (N_2061,N_1982,N_1929);
nand U2062 (N_2062,N_1970,N_1796);
and U2063 (N_2063,N_1775,N_1872);
nand U2064 (N_2064,N_1909,N_1823);
and U2065 (N_2065,N_1943,N_1965);
xor U2066 (N_2066,N_1784,N_1896);
nor U2067 (N_2067,N_1866,N_1846);
and U2068 (N_2068,N_1884,N_1863);
and U2069 (N_2069,N_1786,N_1753);
nand U2070 (N_2070,N_1986,N_1882);
nand U2071 (N_2071,N_1975,N_1789);
nand U2072 (N_2072,N_1894,N_1920);
or U2073 (N_2073,N_1976,N_1890);
nand U2074 (N_2074,N_1779,N_1820);
and U2075 (N_2075,N_1895,N_1873);
or U2076 (N_2076,N_1934,N_1883);
xor U2077 (N_2077,N_1969,N_1889);
nor U2078 (N_2078,N_1804,N_1760);
xor U2079 (N_2079,N_1893,N_1980);
nor U2080 (N_2080,N_1810,N_1812);
nand U2081 (N_2081,N_1809,N_1987);
nand U2082 (N_2082,N_1958,N_1845);
xnor U2083 (N_2083,N_1880,N_1752);
nand U2084 (N_2084,N_1985,N_1999);
xor U2085 (N_2085,N_1919,N_1825);
and U2086 (N_2086,N_1792,N_1776);
nand U2087 (N_2087,N_1937,N_1858);
and U2088 (N_2088,N_1830,N_1869);
nor U2089 (N_2089,N_1795,N_1836);
xnor U2090 (N_2090,N_1991,N_1816);
nor U2091 (N_2091,N_1765,N_1856);
or U2092 (N_2092,N_1766,N_1906);
nor U2093 (N_2093,N_1899,N_1821);
or U2094 (N_2094,N_1916,N_1952);
xor U2095 (N_2095,N_1855,N_1838);
nand U2096 (N_2096,N_1907,N_1843);
and U2097 (N_2097,N_1950,N_1990);
nor U2098 (N_2098,N_1785,N_1914);
nor U2099 (N_2099,N_1835,N_1831);
and U2100 (N_2100,N_1801,N_1908);
nor U2101 (N_2101,N_1755,N_1852);
nor U2102 (N_2102,N_1930,N_1757);
nand U2103 (N_2103,N_1861,N_1837);
nand U2104 (N_2104,N_1787,N_1806);
or U2105 (N_2105,N_1922,N_1868);
nor U2106 (N_2106,N_1960,N_1968);
or U2107 (N_2107,N_1941,N_1758);
xor U2108 (N_2108,N_1993,N_1769);
or U2109 (N_2109,N_1877,N_1885);
or U2110 (N_2110,N_1905,N_1774);
nor U2111 (N_2111,N_1793,N_1998);
xor U2112 (N_2112,N_1971,N_1942);
nor U2113 (N_2113,N_1995,N_1802);
nand U2114 (N_2114,N_1833,N_1897);
nand U2115 (N_2115,N_1857,N_1886);
nand U2116 (N_2116,N_1818,N_1860);
and U2117 (N_2117,N_1770,N_1955);
nor U2118 (N_2118,N_1945,N_1759);
and U2119 (N_2119,N_1867,N_1851);
nor U2120 (N_2120,N_1901,N_1807);
nor U2121 (N_2121,N_1832,N_1805);
or U2122 (N_2122,N_1822,N_1791);
nor U2123 (N_2123,N_1936,N_1947);
and U2124 (N_2124,N_1850,N_1824);
nand U2125 (N_2125,N_1790,N_1914);
nor U2126 (N_2126,N_1983,N_1800);
or U2127 (N_2127,N_1819,N_1987);
xnor U2128 (N_2128,N_1813,N_1844);
or U2129 (N_2129,N_1890,N_1965);
xnor U2130 (N_2130,N_1802,N_1814);
and U2131 (N_2131,N_1845,N_1957);
xor U2132 (N_2132,N_1983,N_1961);
nor U2133 (N_2133,N_1882,N_1874);
and U2134 (N_2134,N_1772,N_1812);
and U2135 (N_2135,N_1968,N_1819);
nor U2136 (N_2136,N_1775,N_1773);
xnor U2137 (N_2137,N_1986,N_1793);
nor U2138 (N_2138,N_1992,N_1909);
xor U2139 (N_2139,N_1941,N_1781);
xor U2140 (N_2140,N_1891,N_1925);
and U2141 (N_2141,N_1897,N_1805);
nor U2142 (N_2142,N_1923,N_1926);
nand U2143 (N_2143,N_1802,N_1896);
and U2144 (N_2144,N_1796,N_1985);
xnor U2145 (N_2145,N_1978,N_1754);
and U2146 (N_2146,N_1981,N_1797);
and U2147 (N_2147,N_1980,N_1750);
or U2148 (N_2148,N_1948,N_1776);
xor U2149 (N_2149,N_1772,N_1750);
and U2150 (N_2150,N_1961,N_1904);
xnor U2151 (N_2151,N_1865,N_1784);
or U2152 (N_2152,N_1878,N_1812);
nand U2153 (N_2153,N_1754,N_1944);
nand U2154 (N_2154,N_1765,N_1919);
or U2155 (N_2155,N_1756,N_1835);
xnor U2156 (N_2156,N_1990,N_1954);
nand U2157 (N_2157,N_1871,N_1924);
or U2158 (N_2158,N_1811,N_1925);
or U2159 (N_2159,N_1879,N_1813);
nand U2160 (N_2160,N_1891,N_1923);
nor U2161 (N_2161,N_1937,N_1864);
xnor U2162 (N_2162,N_1931,N_1939);
nand U2163 (N_2163,N_1823,N_1965);
and U2164 (N_2164,N_1785,N_1918);
nand U2165 (N_2165,N_1770,N_1779);
nand U2166 (N_2166,N_1926,N_1773);
xnor U2167 (N_2167,N_1779,N_1867);
nor U2168 (N_2168,N_1778,N_1829);
or U2169 (N_2169,N_1958,N_1860);
nor U2170 (N_2170,N_1853,N_1862);
nor U2171 (N_2171,N_1926,N_1976);
xor U2172 (N_2172,N_1949,N_1826);
nor U2173 (N_2173,N_1988,N_1851);
nand U2174 (N_2174,N_1929,N_1768);
or U2175 (N_2175,N_1755,N_1861);
or U2176 (N_2176,N_1764,N_1853);
or U2177 (N_2177,N_1916,N_1902);
xnor U2178 (N_2178,N_1902,N_1860);
or U2179 (N_2179,N_1956,N_1988);
nand U2180 (N_2180,N_1851,N_1968);
nand U2181 (N_2181,N_1954,N_1757);
nor U2182 (N_2182,N_1987,N_1900);
and U2183 (N_2183,N_1984,N_1935);
xor U2184 (N_2184,N_1917,N_1971);
and U2185 (N_2185,N_1922,N_1998);
or U2186 (N_2186,N_1911,N_1874);
nor U2187 (N_2187,N_1837,N_1820);
xnor U2188 (N_2188,N_1782,N_1780);
nand U2189 (N_2189,N_1770,N_1962);
and U2190 (N_2190,N_1829,N_1816);
nor U2191 (N_2191,N_1974,N_1794);
nor U2192 (N_2192,N_1833,N_1892);
nor U2193 (N_2193,N_1994,N_1920);
nand U2194 (N_2194,N_1883,N_1943);
nand U2195 (N_2195,N_1794,N_1768);
or U2196 (N_2196,N_1999,N_1815);
nor U2197 (N_2197,N_1946,N_1771);
nand U2198 (N_2198,N_1912,N_1990);
nand U2199 (N_2199,N_1877,N_1860);
xnor U2200 (N_2200,N_1910,N_1962);
or U2201 (N_2201,N_1983,N_1761);
xnor U2202 (N_2202,N_1812,N_1807);
nand U2203 (N_2203,N_1794,N_1808);
nand U2204 (N_2204,N_1956,N_1872);
or U2205 (N_2205,N_1998,N_1941);
nand U2206 (N_2206,N_1960,N_1893);
xor U2207 (N_2207,N_1782,N_1974);
or U2208 (N_2208,N_1954,N_1892);
nor U2209 (N_2209,N_1756,N_1777);
nor U2210 (N_2210,N_1784,N_1979);
xor U2211 (N_2211,N_1797,N_1774);
and U2212 (N_2212,N_1881,N_1800);
or U2213 (N_2213,N_1774,N_1870);
nand U2214 (N_2214,N_1824,N_1763);
xnor U2215 (N_2215,N_1954,N_1827);
xor U2216 (N_2216,N_1998,N_1988);
xor U2217 (N_2217,N_1898,N_1880);
nor U2218 (N_2218,N_1849,N_1862);
xnor U2219 (N_2219,N_1964,N_1757);
nor U2220 (N_2220,N_1836,N_1967);
or U2221 (N_2221,N_1957,N_1911);
and U2222 (N_2222,N_1885,N_1858);
or U2223 (N_2223,N_1814,N_1924);
nor U2224 (N_2224,N_1902,N_1828);
nand U2225 (N_2225,N_1905,N_1895);
and U2226 (N_2226,N_1894,N_1907);
xnor U2227 (N_2227,N_1817,N_1970);
xnor U2228 (N_2228,N_1983,N_1988);
nor U2229 (N_2229,N_1980,N_1787);
or U2230 (N_2230,N_1885,N_1750);
nand U2231 (N_2231,N_1846,N_1892);
xnor U2232 (N_2232,N_1837,N_1939);
or U2233 (N_2233,N_1797,N_1883);
xnor U2234 (N_2234,N_1983,N_1990);
nor U2235 (N_2235,N_1935,N_1986);
and U2236 (N_2236,N_1961,N_1943);
or U2237 (N_2237,N_1892,N_1802);
nand U2238 (N_2238,N_1896,N_1844);
and U2239 (N_2239,N_1918,N_1967);
nand U2240 (N_2240,N_1878,N_1886);
or U2241 (N_2241,N_1866,N_1901);
or U2242 (N_2242,N_1978,N_1800);
and U2243 (N_2243,N_1778,N_1837);
or U2244 (N_2244,N_1990,N_1782);
nor U2245 (N_2245,N_1881,N_1942);
or U2246 (N_2246,N_1784,N_1807);
nor U2247 (N_2247,N_1982,N_1899);
nor U2248 (N_2248,N_1840,N_1902);
or U2249 (N_2249,N_1793,N_1925);
nand U2250 (N_2250,N_2102,N_2055);
or U2251 (N_2251,N_2037,N_2026);
and U2252 (N_2252,N_2160,N_2205);
and U2253 (N_2253,N_2113,N_2098);
and U2254 (N_2254,N_2210,N_2175);
and U2255 (N_2255,N_2245,N_2018);
or U2256 (N_2256,N_2233,N_2215);
or U2257 (N_2257,N_2019,N_2216);
and U2258 (N_2258,N_2114,N_2115);
xor U2259 (N_2259,N_2053,N_2099);
nor U2260 (N_2260,N_2234,N_2035);
or U2261 (N_2261,N_2156,N_2198);
xnor U2262 (N_2262,N_2145,N_2066);
xnor U2263 (N_2263,N_2000,N_2208);
nor U2264 (N_2264,N_2191,N_2069);
and U2265 (N_2265,N_2087,N_2050);
nand U2266 (N_2266,N_2101,N_2075);
nand U2267 (N_2267,N_2025,N_2039);
and U2268 (N_2268,N_2243,N_2119);
nor U2269 (N_2269,N_2047,N_2034);
xor U2270 (N_2270,N_2057,N_2015);
or U2271 (N_2271,N_2096,N_2189);
and U2272 (N_2272,N_2067,N_2150);
xor U2273 (N_2273,N_2173,N_2029);
or U2274 (N_2274,N_2152,N_2120);
nand U2275 (N_2275,N_2185,N_2202);
nand U2276 (N_2276,N_2190,N_2092);
or U2277 (N_2277,N_2011,N_2169);
nor U2278 (N_2278,N_2227,N_2064);
or U2279 (N_2279,N_2084,N_2036);
nor U2280 (N_2280,N_2006,N_2248);
nand U2281 (N_2281,N_2164,N_2027);
xor U2282 (N_2282,N_2007,N_2103);
nand U2283 (N_2283,N_2242,N_2163);
and U2284 (N_2284,N_2123,N_2199);
nand U2285 (N_2285,N_2105,N_2144);
and U2286 (N_2286,N_2182,N_2054);
and U2287 (N_2287,N_2080,N_2060);
or U2288 (N_2288,N_2091,N_2238);
and U2289 (N_2289,N_2082,N_2168);
nand U2290 (N_2290,N_2237,N_2016);
nor U2291 (N_2291,N_2009,N_2194);
nand U2292 (N_2292,N_2157,N_2042);
nand U2293 (N_2293,N_2112,N_2241);
xor U2294 (N_2294,N_2229,N_2062);
nor U2295 (N_2295,N_2024,N_2228);
and U2296 (N_2296,N_2162,N_2124);
nand U2297 (N_2297,N_2158,N_2240);
or U2298 (N_2298,N_2170,N_2032);
and U2299 (N_2299,N_2030,N_2065);
xnor U2300 (N_2300,N_2209,N_2140);
or U2301 (N_2301,N_2131,N_2121);
nand U2302 (N_2302,N_2077,N_2108);
nand U2303 (N_2303,N_2063,N_2188);
nor U2304 (N_2304,N_2212,N_2038);
and U2305 (N_2305,N_2197,N_2088);
xnor U2306 (N_2306,N_2225,N_2154);
and U2307 (N_2307,N_2127,N_2122);
and U2308 (N_2308,N_2213,N_2167);
xnor U2309 (N_2309,N_2236,N_2166);
nand U2310 (N_2310,N_2085,N_2222);
and U2311 (N_2311,N_2071,N_2200);
nand U2312 (N_2312,N_2070,N_2044);
nor U2313 (N_2313,N_2218,N_2141);
xor U2314 (N_2314,N_2181,N_2004);
and U2315 (N_2315,N_2072,N_2220);
or U2316 (N_2316,N_2049,N_2184);
nor U2317 (N_2317,N_2183,N_2224);
and U2318 (N_2318,N_2109,N_2143);
nor U2319 (N_2319,N_2142,N_2023);
and U2320 (N_2320,N_2043,N_2132);
nor U2321 (N_2321,N_2155,N_2020);
and U2322 (N_2322,N_2244,N_2217);
nor U2323 (N_2323,N_2081,N_2079);
or U2324 (N_2324,N_2097,N_2001);
or U2325 (N_2325,N_2161,N_2178);
nand U2326 (N_2326,N_2171,N_2147);
xnor U2327 (N_2327,N_2211,N_2110);
nand U2328 (N_2328,N_2136,N_2028);
xor U2329 (N_2329,N_2204,N_2090);
nor U2330 (N_2330,N_2022,N_2203);
nor U2331 (N_2331,N_2104,N_2179);
nor U2332 (N_2332,N_2031,N_2247);
xnor U2333 (N_2333,N_2040,N_2125);
nand U2334 (N_2334,N_2058,N_2094);
nand U2335 (N_2335,N_2153,N_2187);
and U2336 (N_2336,N_2186,N_2116);
and U2337 (N_2337,N_2008,N_2107);
xnor U2338 (N_2338,N_2100,N_2207);
nor U2339 (N_2339,N_2195,N_2012);
xnor U2340 (N_2340,N_2048,N_2073);
and U2341 (N_2341,N_2021,N_2014);
or U2342 (N_2342,N_2126,N_2149);
nand U2343 (N_2343,N_2111,N_2095);
nor U2344 (N_2344,N_2106,N_2045);
or U2345 (N_2345,N_2135,N_2076);
and U2346 (N_2346,N_2172,N_2059);
nand U2347 (N_2347,N_2176,N_2231);
or U2348 (N_2348,N_2010,N_2005);
xor U2349 (N_2349,N_2083,N_2138);
xnor U2350 (N_2350,N_2133,N_2130);
xnor U2351 (N_2351,N_2128,N_2051);
nand U2352 (N_2352,N_2196,N_2017);
xor U2353 (N_2353,N_2239,N_2118);
xor U2354 (N_2354,N_2129,N_2219);
and U2355 (N_2355,N_2221,N_2052);
or U2356 (N_2356,N_2201,N_2232);
and U2357 (N_2357,N_2061,N_2013);
or U2358 (N_2358,N_2246,N_2074);
and U2359 (N_2359,N_2180,N_2146);
nand U2360 (N_2360,N_2177,N_2159);
and U2361 (N_2361,N_2117,N_2093);
or U2362 (N_2362,N_2046,N_2235);
and U2363 (N_2363,N_2206,N_2056);
xnor U2364 (N_2364,N_2068,N_2003);
nand U2365 (N_2365,N_2002,N_2193);
xor U2366 (N_2366,N_2151,N_2230);
or U2367 (N_2367,N_2134,N_2086);
nor U2368 (N_2368,N_2192,N_2137);
and U2369 (N_2369,N_2078,N_2165);
xor U2370 (N_2370,N_2226,N_2033);
xnor U2371 (N_2371,N_2223,N_2249);
or U2372 (N_2372,N_2148,N_2174);
and U2373 (N_2373,N_2214,N_2139);
or U2374 (N_2374,N_2089,N_2041);
nand U2375 (N_2375,N_2238,N_2069);
or U2376 (N_2376,N_2051,N_2240);
nor U2377 (N_2377,N_2227,N_2079);
nor U2378 (N_2378,N_2041,N_2101);
and U2379 (N_2379,N_2195,N_2190);
or U2380 (N_2380,N_2052,N_2228);
and U2381 (N_2381,N_2175,N_2123);
xnor U2382 (N_2382,N_2015,N_2002);
xor U2383 (N_2383,N_2228,N_2021);
nand U2384 (N_2384,N_2201,N_2106);
and U2385 (N_2385,N_2085,N_2130);
nand U2386 (N_2386,N_2217,N_2049);
nor U2387 (N_2387,N_2166,N_2161);
nor U2388 (N_2388,N_2234,N_2235);
and U2389 (N_2389,N_2062,N_2244);
and U2390 (N_2390,N_2240,N_2003);
nand U2391 (N_2391,N_2248,N_2206);
nor U2392 (N_2392,N_2001,N_2020);
xor U2393 (N_2393,N_2115,N_2168);
nor U2394 (N_2394,N_2087,N_2145);
or U2395 (N_2395,N_2225,N_2244);
xnor U2396 (N_2396,N_2128,N_2191);
nor U2397 (N_2397,N_2133,N_2111);
or U2398 (N_2398,N_2154,N_2089);
or U2399 (N_2399,N_2127,N_2031);
and U2400 (N_2400,N_2220,N_2209);
nor U2401 (N_2401,N_2130,N_2201);
nand U2402 (N_2402,N_2098,N_2176);
nor U2403 (N_2403,N_2028,N_2080);
or U2404 (N_2404,N_2047,N_2024);
and U2405 (N_2405,N_2011,N_2120);
and U2406 (N_2406,N_2183,N_2083);
or U2407 (N_2407,N_2013,N_2129);
nor U2408 (N_2408,N_2090,N_2190);
or U2409 (N_2409,N_2114,N_2128);
and U2410 (N_2410,N_2067,N_2245);
nand U2411 (N_2411,N_2055,N_2091);
or U2412 (N_2412,N_2232,N_2249);
or U2413 (N_2413,N_2213,N_2097);
nor U2414 (N_2414,N_2150,N_2164);
nand U2415 (N_2415,N_2004,N_2213);
or U2416 (N_2416,N_2061,N_2174);
or U2417 (N_2417,N_2119,N_2125);
and U2418 (N_2418,N_2133,N_2061);
xnor U2419 (N_2419,N_2013,N_2041);
or U2420 (N_2420,N_2146,N_2044);
xnor U2421 (N_2421,N_2110,N_2238);
or U2422 (N_2422,N_2008,N_2087);
nand U2423 (N_2423,N_2185,N_2156);
xor U2424 (N_2424,N_2070,N_2073);
nand U2425 (N_2425,N_2032,N_2169);
nand U2426 (N_2426,N_2065,N_2221);
or U2427 (N_2427,N_2162,N_2050);
or U2428 (N_2428,N_2232,N_2008);
and U2429 (N_2429,N_2082,N_2088);
nand U2430 (N_2430,N_2191,N_2176);
xor U2431 (N_2431,N_2094,N_2019);
xor U2432 (N_2432,N_2219,N_2082);
xnor U2433 (N_2433,N_2119,N_2246);
nor U2434 (N_2434,N_2149,N_2144);
or U2435 (N_2435,N_2136,N_2115);
nand U2436 (N_2436,N_2006,N_2152);
xor U2437 (N_2437,N_2143,N_2160);
xnor U2438 (N_2438,N_2130,N_2015);
xor U2439 (N_2439,N_2155,N_2024);
xor U2440 (N_2440,N_2041,N_2120);
xnor U2441 (N_2441,N_2208,N_2165);
or U2442 (N_2442,N_2181,N_2186);
xnor U2443 (N_2443,N_2155,N_2236);
nor U2444 (N_2444,N_2110,N_2127);
xnor U2445 (N_2445,N_2233,N_2244);
and U2446 (N_2446,N_2205,N_2085);
nor U2447 (N_2447,N_2100,N_2173);
xnor U2448 (N_2448,N_2149,N_2140);
nand U2449 (N_2449,N_2078,N_2105);
xor U2450 (N_2450,N_2024,N_2082);
and U2451 (N_2451,N_2052,N_2188);
xor U2452 (N_2452,N_2133,N_2217);
nor U2453 (N_2453,N_2155,N_2209);
xor U2454 (N_2454,N_2156,N_2060);
nor U2455 (N_2455,N_2048,N_2090);
nand U2456 (N_2456,N_2203,N_2023);
nor U2457 (N_2457,N_2014,N_2195);
nor U2458 (N_2458,N_2204,N_2149);
and U2459 (N_2459,N_2041,N_2057);
xor U2460 (N_2460,N_2127,N_2114);
nand U2461 (N_2461,N_2129,N_2241);
nand U2462 (N_2462,N_2236,N_2200);
xor U2463 (N_2463,N_2057,N_2161);
and U2464 (N_2464,N_2058,N_2161);
or U2465 (N_2465,N_2047,N_2079);
and U2466 (N_2466,N_2151,N_2114);
nand U2467 (N_2467,N_2032,N_2016);
xor U2468 (N_2468,N_2248,N_2181);
nor U2469 (N_2469,N_2017,N_2149);
or U2470 (N_2470,N_2074,N_2079);
xnor U2471 (N_2471,N_2080,N_2003);
xor U2472 (N_2472,N_2224,N_2246);
or U2473 (N_2473,N_2150,N_2023);
and U2474 (N_2474,N_2187,N_2069);
and U2475 (N_2475,N_2184,N_2236);
and U2476 (N_2476,N_2037,N_2001);
nor U2477 (N_2477,N_2233,N_2127);
nand U2478 (N_2478,N_2084,N_2089);
nor U2479 (N_2479,N_2241,N_2237);
or U2480 (N_2480,N_2170,N_2212);
nor U2481 (N_2481,N_2106,N_2196);
nand U2482 (N_2482,N_2203,N_2216);
nor U2483 (N_2483,N_2193,N_2237);
and U2484 (N_2484,N_2021,N_2130);
or U2485 (N_2485,N_2112,N_2098);
and U2486 (N_2486,N_2071,N_2080);
xor U2487 (N_2487,N_2123,N_2133);
nand U2488 (N_2488,N_2116,N_2069);
xor U2489 (N_2489,N_2125,N_2204);
nand U2490 (N_2490,N_2241,N_2206);
and U2491 (N_2491,N_2248,N_2237);
and U2492 (N_2492,N_2040,N_2020);
nor U2493 (N_2493,N_2004,N_2088);
and U2494 (N_2494,N_2222,N_2083);
or U2495 (N_2495,N_2186,N_2151);
nand U2496 (N_2496,N_2228,N_2179);
and U2497 (N_2497,N_2165,N_2194);
and U2498 (N_2498,N_2021,N_2042);
and U2499 (N_2499,N_2243,N_2081);
xor U2500 (N_2500,N_2440,N_2327);
xor U2501 (N_2501,N_2449,N_2454);
or U2502 (N_2502,N_2334,N_2391);
or U2503 (N_2503,N_2411,N_2419);
or U2504 (N_2504,N_2258,N_2371);
nand U2505 (N_2505,N_2387,N_2310);
nand U2506 (N_2506,N_2279,N_2294);
and U2507 (N_2507,N_2403,N_2357);
and U2508 (N_2508,N_2393,N_2392);
or U2509 (N_2509,N_2376,N_2490);
xnor U2510 (N_2510,N_2486,N_2434);
xnor U2511 (N_2511,N_2460,N_2343);
or U2512 (N_2512,N_2308,N_2420);
and U2513 (N_2513,N_2396,N_2283);
nor U2514 (N_2514,N_2312,N_2274);
or U2515 (N_2515,N_2452,N_2468);
and U2516 (N_2516,N_2293,N_2325);
nand U2517 (N_2517,N_2394,N_2342);
nor U2518 (N_2518,N_2444,N_2455);
or U2519 (N_2519,N_2286,N_2443);
and U2520 (N_2520,N_2442,N_2317);
and U2521 (N_2521,N_2470,N_2353);
nor U2522 (N_2522,N_2412,N_2356);
and U2523 (N_2523,N_2451,N_2472);
nor U2524 (N_2524,N_2354,N_2474);
nor U2525 (N_2525,N_2370,N_2290);
xor U2526 (N_2526,N_2263,N_2288);
or U2527 (N_2527,N_2358,N_2402);
or U2528 (N_2528,N_2422,N_2269);
nor U2529 (N_2529,N_2477,N_2453);
nand U2530 (N_2530,N_2259,N_2368);
or U2531 (N_2531,N_2298,N_2331);
and U2532 (N_2532,N_2446,N_2311);
and U2533 (N_2533,N_2377,N_2268);
or U2534 (N_2534,N_2487,N_2302);
nand U2535 (N_2535,N_2417,N_2359);
xnor U2536 (N_2536,N_2266,N_2438);
or U2537 (N_2537,N_2471,N_2345);
nand U2538 (N_2538,N_2480,N_2355);
or U2539 (N_2539,N_2265,N_2448);
xnor U2540 (N_2540,N_2260,N_2459);
and U2541 (N_2541,N_2369,N_2306);
xnor U2542 (N_2542,N_2257,N_2352);
nor U2543 (N_2543,N_2299,N_2300);
and U2544 (N_2544,N_2284,N_2305);
and U2545 (N_2545,N_2322,N_2333);
or U2546 (N_2546,N_2496,N_2366);
xnor U2547 (N_2547,N_2278,N_2253);
and U2548 (N_2548,N_2330,N_2479);
or U2549 (N_2549,N_2489,N_2292);
nand U2550 (N_2550,N_2273,N_2491);
nand U2551 (N_2551,N_2493,N_2383);
xor U2552 (N_2552,N_2349,N_2484);
and U2553 (N_2553,N_2347,N_2436);
and U2554 (N_2554,N_2262,N_2335);
nor U2555 (N_2555,N_2375,N_2339);
nor U2556 (N_2556,N_2428,N_2314);
or U2557 (N_2557,N_2432,N_2447);
xor U2558 (N_2558,N_2388,N_2464);
or U2559 (N_2559,N_2285,N_2457);
and U2560 (N_2560,N_2261,N_2476);
xnor U2561 (N_2561,N_2337,N_2297);
or U2562 (N_2562,N_2316,N_2418);
nor U2563 (N_2563,N_2341,N_2367);
or U2564 (N_2564,N_2344,N_2276);
nand U2565 (N_2565,N_2326,N_2431);
nor U2566 (N_2566,N_2473,N_2414);
or U2567 (N_2567,N_2360,N_2365);
and U2568 (N_2568,N_2324,N_2483);
and U2569 (N_2569,N_2421,N_2475);
nand U2570 (N_2570,N_2406,N_2423);
nand U2571 (N_2571,N_2320,N_2361);
and U2572 (N_2572,N_2433,N_2315);
or U2573 (N_2573,N_2296,N_2427);
xnor U2574 (N_2574,N_2374,N_2463);
xor U2575 (N_2575,N_2372,N_2363);
nor U2576 (N_2576,N_2348,N_2362);
or U2577 (N_2577,N_2267,N_2282);
or U2578 (N_2578,N_2413,N_2478);
nand U2579 (N_2579,N_2287,N_2424);
nor U2580 (N_2580,N_2425,N_2405);
xnor U2581 (N_2581,N_2398,N_2323);
xor U2582 (N_2582,N_2439,N_2329);
xnor U2583 (N_2583,N_2498,N_2488);
or U2584 (N_2584,N_2461,N_2381);
nor U2585 (N_2585,N_2379,N_2401);
and U2586 (N_2586,N_2280,N_2408);
nand U2587 (N_2587,N_2373,N_2271);
nand U2588 (N_2588,N_2307,N_2437);
or U2589 (N_2589,N_2336,N_2499);
nand U2590 (N_2590,N_2426,N_2275);
or U2591 (N_2591,N_2321,N_2364);
nor U2592 (N_2592,N_2482,N_2458);
nor U2593 (N_2593,N_2252,N_2407);
nand U2594 (N_2594,N_2304,N_2469);
xnor U2595 (N_2595,N_2497,N_2466);
nor U2596 (N_2596,N_2389,N_2303);
or U2597 (N_2597,N_2465,N_2462);
and U2598 (N_2598,N_2380,N_2390);
nand U2599 (N_2599,N_2378,N_2250);
or U2600 (N_2600,N_2386,N_2485);
nand U2601 (N_2601,N_2289,N_2251);
and U2602 (N_2602,N_2399,N_2291);
nor U2603 (N_2603,N_2467,N_2346);
or U2604 (N_2604,N_2456,N_2301);
or U2605 (N_2605,N_2309,N_2350);
or U2606 (N_2606,N_2332,N_2319);
xor U2607 (N_2607,N_2494,N_2277);
or U2608 (N_2608,N_2264,N_2318);
and U2609 (N_2609,N_2410,N_2481);
nor U2610 (N_2610,N_2435,N_2256);
xor U2611 (N_2611,N_2430,N_2404);
and U2612 (N_2612,N_2382,N_2272);
or U2613 (N_2613,N_2328,N_2397);
or U2614 (N_2614,N_2400,N_2313);
nand U2615 (N_2615,N_2385,N_2384);
or U2616 (N_2616,N_2495,N_2295);
xor U2617 (N_2617,N_2270,N_2450);
xor U2618 (N_2618,N_2255,N_2429);
nor U2619 (N_2619,N_2416,N_2492);
nand U2620 (N_2620,N_2409,N_2254);
nor U2621 (N_2621,N_2441,N_2445);
xor U2622 (N_2622,N_2351,N_2338);
or U2623 (N_2623,N_2340,N_2281);
nor U2624 (N_2624,N_2395,N_2415);
nand U2625 (N_2625,N_2273,N_2254);
and U2626 (N_2626,N_2408,N_2423);
nand U2627 (N_2627,N_2495,N_2339);
nand U2628 (N_2628,N_2368,N_2283);
xnor U2629 (N_2629,N_2266,N_2358);
nor U2630 (N_2630,N_2307,N_2294);
xor U2631 (N_2631,N_2319,N_2398);
nor U2632 (N_2632,N_2427,N_2408);
nor U2633 (N_2633,N_2307,N_2322);
nand U2634 (N_2634,N_2498,N_2338);
or U2635 (N_2635,N_2495,N_2328);
nor U2636 (N_2636,N_2371,N_2387);
or U2637 (N_2637,N_2492,N_2413);
or U2638 (N_2638,N_2446,N_2498);
xnor U2639 (N_2639,N_2450,N_2339);
nand U2640 (N_2640,N_2337,N_2315);
or U2641 (N_2641,N_2361,N_2260);
or U2642 (N_2642,N_2332,N_2468);
nand U2643 (N_2643,N_2313,N_2377);
and U2644 (N_2644,N_2432,N_2301);
nor U2645 (N_2645,N_2280,N_2393);
or U2646 (N_2646,N_2458,N_2495);
nand U2647 (N_2647,N_2385,N_2263);
and U2648 (N_2648,N_2369,N_2400);
or U2649 (N_2649,N_2258,N_2269);
and U2650 (N_2650,N_2333,N_2313);
nor U2651 (N_2651,N_2448,N_2487);
nand U2652 (N_2652,N_2276,N_2269);
xnor U2653 (N_2653,N_2381,N_2490);
nor U2654 (N_2654,N_2366,N_2255);
xnor U2655 (N_2655,N_2324,N_2419);
or U2656 (N_2656,N_2420,N_2488);
xnor U2657 (N_2657,N_2432,N_2366);
xnor U2658 (N_2658,N_2421,N_2258);
nor U2659 (N_2659,N_2327,N_2466);
nor U2660 (N_2660,N_2347,N_2304);
xor U2661 (N_2661,N_2479,N_2387);
nand U2662 (N_2662,N_2382,N_2485);
nand U2663 (N_2663,N_2298,N_2296);
or U2664 (N_2664,N_2278,N_2341);
nand U2665 (N_2665,N_2427,N_2433);
or U2666 (N_2666,N_2292,N_2403);
and U2667 (N_2667,N_2408,N_2312);
xor U2668 (N_2668,N_2289,N_2487);
or U2669 (N_2669,N_2434,N_2443);
nor U2670 (N_2670,N_2496,N_2419);
nand U2671 (N_2671,N_2252,N_2493);
and U2672 (N_2672,N_2469,N_2402);
nor U2673 (N_2673,N_2255,N_2445);
xor U2674 (N_2674,N_2493,N_2256);
or U2675 (N_2675,N_2490,N_2306);
xnor U2676 (N_2676,N_2432,N_2460);
and U2677 (N_2677,N_2470,N_2250);
or U2678 (N_2678,N_2352,N_2264);
xnor U2679 (N_2679,N_2466,N_2282);
xnor U2680 (N_2680,N_2480,N_2415);
and U2681 (N_2681,N_2353,N_2327);
nor U2682 (N_2682,N_2325,N_2468);
or U2683 (N_2683,N_2439,N_2438);
nor U2684 (N_2684,N_2427,N_2338);
and U2685 (N_2685,N_2462,N_2458);
or U2686 (N_2686,N_2449,N_2426);
and U2687 (N_2687,N_2383,N_2359);
or U2688 (N_2688,N_2424,N_2341);
nor U2689 (N_2689,N_2394,N_2387);
and U2690 (N_2690,N_2434,N_2499);
xnor U2691 (N_2691,N_2393,N_2493);
and U2692 (N_2692,N_2391,N_2381);
xor U2693 (N_2693,N_2498,N_2360);
xnor U2694 (N_2694,N_2343,N_2489);
nand U2695 (N_2695,N_2357,N_2309);
and U2696 (N_2696,N_2359,N_2275);
nor U2697 (N_2697,N_2335,N_2476);
nor U2698 (N_2698,N_2348,N_2361);
nand U2699 (N_2699,N_2474,N_2388);
nand U2700 (N_2700,N_2483,N_2264);
xor U2701 (N_2701,N_2314,N_2398);
or U2702 (N_2702,N_2353,N_2430);
nand U2703 (N_2703,N_2371,N_2289);
xor U2704 (N_2704,N_2349,N_2489);
nand U2705 (N_2705,N_2298,N_2278);
and U2706 (N_2706,N_2422,N_2291);
nand U2707 (N_2707,N_2300,N_2425);
and U2708 (N_2708,N_2376,N_2345);
nor U2709 (N_2709,N_2352,N_2266);
nor U2710 (N_2710,N_2477,N_2480);
nor U2711 (N_2711,N_2451,N_2431);
or U2712 (N_2712,N_2278,N_2375);
and U2713 (N_2713,N_2497,N_2332);
nand U2714 (N_2714,N_2470,N_2404);
and U2715 (N_2715,N_2490,N_2408);
or U2716 (N_2716,N_2374,N_2402);
nor U2717 (N_2717,N_2353,N_2260);
nor U2718 (N_2718,N_2299,N_2347);
nand U2719 (N_2719,N_2449,N_2262);
xor U2720 (N_2720,N_2254,N_2460);
nand U2721 (N_2721,N_2382,N_2412);
nand U2722 (N_2722,N_2338,N_2487);
and U2723 (N_2723,N_2461,N_2398);
xnor U2724 (N_2724,N_2455,N_2317);
xor U2725 (N_2725,N_2451,N_2310);
xnor U2726 (N_2726,N_2488,N_2433);
nand U2727 (N_2727,N_2428,N_2288);
nor U2728 (N_2728,N_2397,N_2418);
or U2729 (N_2729,N_2470,N_2491);
nand U2730 (N_2730,N_2296,N_2461);
xor U2731 (N_2731,N_2490,N_2255);
and U2732 (N_2732,N_2412,N_2399);
nand U2733 (N_2733,N_2428,N_2418);
and U2734 (N_2734,N_2479,N_2287);
and U2735 (N_2735,N_2414,N_2360);
nor U2736 (N_2736,N_2365,N_2410);
or U2737 (N_2737,N_2291,N_2391);
nand U2738 (N_2738,N_2414,N_2295);
and U2739 (N_2739,N_2469,N_2458);
nor U2740 (N_2740,N_2396,N_2422);
or U2741 (N_2741,N_2278,N_2371);
xnor U2742 (N_2742,N_2306,N_2266);
and U2743 (N_2743,N_2290,N_2344);
nand U2744 (N_2744,N_2317,N_2394);
and U2745 (N_2745,N_2481,N_2264);
nand U2746 (N_2746,N_2496,N_2386);
xnor U2747 (N_2747,N_2288,N_2411);
nor U2748 (N_2748,N_2259,N_2455);
nor U2749 (N_2749,N_2495,N_2342);
nor U2750 (N_2750,N_2516,N_2614);
nor U2751 (N_2751,N_2569,N_2581);
and U2752 (N_2752,N_2660,N_2565);
nand U2753 (N_2753,N_2582,N_2633);
or U2754 (N_2754,N_2539,N_2719);
or U2755 (N_2755,N_2650,N_2747);
and U2756 (N_2756,N_2667,N_2654);
and U2757 (N_2757,N_2697,N_2518);
xnor U2758 (N_2758,N_2597,N_2585);
nand U2759 (N_2759,N_2668,N_2725);
and U2760 (N_2760,N_2560,N_2662);
nand U2761 (N_2761,N_2503,N_2551);
or U2762 (N_2762,N_2591,N_2708);
nand U2763 (N_2763,N_2600,N_2621);
or U2764 (N_2764,N_2521,N_2746);
nand U2765 (N_2765,N_2717,N_2615);
nand U2766 (N_2766,N_2564,N_2679);
nand U2767 (N_2767,N_2715,N_2527);
nor U2768 (N_2768,N_2693,N_2661);
or U2769 (N_2769,N_2744,N_2557);
nand U2770 (N_2770,N_2622,N_2664);
nand U2771 (N_2771,N_2563,N_2721);
or U2772 (N_2772,N_2674,N_2580);
xor U2773 (N_2773,N_2528,N_2710);
or U2774 (N_2774,N_2540,N_2500);
or U2775 (N_2775,N_2685,N_2530);
nor U2776 (N_2776,N_2683,N_2651);
and U2777 (N_2777,N_2570,N_2656);
or U2778 (N_2778,N_2595,N_2678);
and U2779 (N_2779,N_2634,N_2712);
xor U2780 (N_2780,N_2576,N_2554);
nand U2781 (N_2781,N_2548,N_2684);
xor U2782 (N_2782,N_2562,N_2502);
or U2783 (N_2783,N_2749,N_2698);
or U2784 (N_2784,N_2707,N_2639);
and U2785 (N_2785,N_2645,N_2726);
or U2786 (N_2786,N_2687,N_2533);
xor U2787 (N_2787,N_2640,N_2529);
and U2788 (N_2788,N_2523,N_2543);
or U2789 (N_2789,N_2709,N_2511);
nand U2790 (N_2790,N_2583,N_2561);
and U2791 (N_2791,N_2524,N_2696);
or U2792 (N_2792,N_2512,N_2659);
nand U2793 (N_2793,N_2720,N_2627);
nor U2794 (N_2794,N_2691,N_2599);
nand U2795 (N_2795,N_2596,N_2532);
xnor U2796 (N_2796,N_2745,N_2743);
xor U2797 (N_2797,N_2713,N_2740);
nand U2798 (N_2798,N_2559,N_2604);
or U2799 (N_2799,N_2728,N_2623);
or U2800 (N_2800,N_2578,N_2724);
xnor U2801 (N_2801,N_2537,N_2670);
and U2802 (N_2802,N_2702,N_2658);
nor U2803 (N_2803,N_2647,N_2626);
nand U2804 (N_2804,N_2606,N_2619);
or U2805 (N_2805,N_2699,N_2526);
nor U2806 (N_2806,N_2663,N_2677);
xnor U2807 (N_2807,N_2598,N_2630);
nor U2808 (N_2808,N_2686,N_2558);
or U2809 (N_2809,N_2680,N_2690);
xnor U2810 (N_2810,N_2592,N_2566);
xnor U2811 (N_2811,N_2586,N_2733);
xor U2812 (N_2812,N_2673,N_2737);
xnor U2813 (N_2813,N_2642,N_2588);
or U2814 (N_2814,N_2629,N_2544);
and U2815 (N_2815,N_2652,N_2522);
or U2816 (N_2816,N_2590,N_2504);
nand U2817 (N_2817,N_2631,N_2605);
or U2818 (N_2818,N_2714,N_2546);
nand U2819 (N_2819,N_2550,N_2517);
nor U2820 (N_2820,N_2632,N_2635);
nand U2821 (N_2821,N_2716,N_2701);
nor U2822 (N_2822,N_2587,N_2536);
and U2823 (N_2823,N_2613,N_2735);
nand U2824 (N_2824,N_2601,N_2602);
nor U2825 (N_2825,N_2547,N_2695);
nand U2826 (N_2826,N_2669,N_2739);
xnor U2827 (N_2827,N_2542,N_2637);
nor U2828 (N_2828,N_2625,N_2531);
xor U2829 (N_2829,N_2589,N_2567);
nand U2830 (N_2830,N_2723,N_2603);
xnor U2831 (N_2831,N_2722,N_2549);
xor U2832 (N_2832,N_2552,N_2538);
xor U2833 (N_2833,N_2742,N_2649);
xnor U2834 (N_2834,N_2688,N_2545);
and U2835 (N_2835,N_2655,N_2718);
nor U2836 (N_2836,N_2577,N_2700);
or U2837 (N_2837,N_2643,N_2572);
and U2838 (N_2838,N_2553,N_2617);
nor U2839 (N_2839,N_2506,N_2675);
xnor U2840 (N_2840,N_2519,N_2568);
or U2841 (N_2841,N_2556,N_2736);
nand U2842 (N_2842,N_2584,N_2731);
or U2843 (N_2843,N_2681,N_2738);
nor U2844 (N_2844,N_2513,N_2648);
and U2845 (N_2845,N_2579,N_2611);
nand U2846 (N_2846,N_2732,N_2628);
and U2847 (N_2847,N_2594,N_2657);
nor U2848 (N_2848,N_2555,N_2620);
xor U2849 (N_2849,N_2509,N_2727);
xnor U2850 (N_2850,N_2535,N_2571);
nand U2851 (N_2851,N_2741,N_2734);
or U2852 (N_2852,N_2609,N_2520);
nor U2853 (N_2853,N_2618,N_2607);
and U2854 (N_2854,N_2671,N_2510);
nor U2855 (N_2855,N_2730,N_2705);
or U2856 (N_2856,N_2624,N_2676);
nand U2857 (N_2857,N_2636,N_2508);
and U2858 (N_2858,N_2505,N_2610);
nor U2859 (N_2859,N_2672,N_2748);
nand U2860 (N_2860,N_2689,N_2501);
or U2861 (N_2861,N_2682,N_2612);
nand U2862 (N_2862,N_2575,N_2616);
nand U2863 (N_2863,N_2541,N_2534);
xor U2864 (N_2864,N_2666,N_2706);
or U2865 (N_2865,N_2646,N_2573);
nand U2866 (N_2866,N_2704,N_2515);
nand U2867 (N_2867,N_2665,N_2641);
nor U2868 (N_2868,N_2711,N_2692);
xor U2869 (N_2869,N_2608,N_2694);
and U2870 (N_2870,N_2729,N_2525);
or U2871 (N_2871,N_2644,N_2514);
nor U2872 (N_2872,N_2653,N_2574);
and U2873 (N_2873,N_2638,N_2593);
or U2874 (N_2874,N_2507,N_2703);
nor U2875 (N_2875,N_2593,N_2708);
nor U2876 (N_2876,N_2708,N_2706);
xnor U2877 (N_2877,N_2601,N_2703);
nand U2878 (N_2878,N_2530,N_2666);
and U2879 (N_2879,N_2534,N_2727);
nor U2880 (N_2880,N_2569,N_2644);
and U2881 (N_2881,N_2682,N_2625);
nor U2882 (N_2882,N_2591,N_2656);
nand U2883 (N_2883,N_2517,N_2711);
and U2884 (N_2884,N_2594,N_2625);
nand U2885 (N_2885,N_2573,N_2664);
xor U2886 (N_2886,N_2609,N_2558);
nand U2887 (N_2887,N_2608,N_2553);
xor U2888 (N_2888,N_2595,N_2630);
xor U2889 (N_2889,N_2706,N_2574);
and U2890 (N_2890,N_2556,N_2523);
nand U2891 (N_2891,N_2560,N_2611);
nand U2892 (N_2892,N_2529,N_2571);
nor U2893 (N_2893,N_2575,N_2619);
nand U2894 (N_2894,N_2686,N_2631);
nor U2895 (N_2895,N_2718,N_2700);
nand U2896 (N_2896,N_2722,N_2690);
xor U2897 (N_2897,N_2613,N_2576);
nand U2898 (N_2898,N_2512,N_2723);
xor U2899 (N_2899,N_2589,N_2602);
nand U2900 (N_2900,N_2611,N_2594);
xor U2901 (N_2901,N_2656,N_2518);
or U2902 (N_2902,N_2584,N_2631);
or U2903 (N_2903,N_2597,N_2728);
or U2904 (N_2904,N_2738,N_2515);
xor U2905 (N_2905,N_2643,N_2539);
xor U2906 (N_2906,N_2633,N_2521);
nand U2907 (N_2907,N_2514,N_2602);
and U2908 (N_2908,N_2589,N_2508);
nor U2909 (N_2909,N_2679,N_2734);
or U2910 (N_2910,N_2557,N_2708);
nand U2911 (N_2911,N_2701,N_2690);
nor U2912 (N_2912,N_2653,N_2576);
xor U2913 (N_2913,N_2633,N_2595);
nor U2914 (N_2914,N_2656,N_2546);
xnor U2915 (N_2915,N_2708,N_2570);
and U2916 (N_2916,N_2576,N_2517);
nand U2917 (N_2917,N_2656,N_2627);
and U2918 (N_2918,N_2546,N_2697);
nand U2919 (N_2919,N_2530,N_2697);
or U2920 (N_2920,N_2591,N_2654);
or U2921 (N_2921,N_2600,N_2669);
or U2922 (N_2922,N_2566,N_2631);
or U2923 (N_2923,N_2550,N_2573);
nor U2924 (N_2924,N_2544,N_2628);
xor U2925 (N_2925,N_2507,N_2546);
xnor U2926 (N_2926,N_2669,N_2534);
or U2927 (N_2927,N_2708,N_2515);
xnor U2928 (N_2928,N_2680,N_2567);
nor U2929 (N_2929,N_2612,N_2607);
nor U2930 (N_2930,N_2580,N_2558);
nand U2931 (N_2931,N_2534,N_2744);
nor U2932 (N_2932,N_2698,N_2735);
nor U2933 (N_2933,N_2574,N_2697);
or U2934 (N_2934,N_2614,N_2552);
and U2935 (N_2935,N_2533,N_2624);
xor U2936 (N_2936,N_2670,N_2602);
or U2937 (N_2937,N_2708,N_2673);
xor U2938 (N_2938,N_2637,N_2569);
nand U2939 (N_2939,N_2576,N_2601);
xnor U2940 (N_2940,N_2603,N_2707);
or U2941 (N_2941,N_2568,N_2586);
nor U2942 (N_2942,N_2550,N_2530);
or U2943 (N_2943,N_2503,N_2706);
xor U2944 (N_2944,N_2606,N_2528);
or U2945 (N_2945,N_2715,N_2623);
or U2946 (N_2946,N_2599,N_2564);
nand U2947 (N_2947,N_2663,N_2506);
or U2948 (N_2948,N_2593,N_2744);
nand U2949 (N_2949,N_2680,N_2607);
xor U2950 (N_2950,N_2601,N_2733);
xor U2951 (N_2951,N_2634,N_2519);
nand U2952 (N_2952,N_2548,N_2718);
or U2953 (N_2953,N_2501,N_2699);
xnor U2954 (N_2954,N_2683,N_2518);
and U2955 (N_2955,N_2720,N_2715);
nand U2956 (N_2956,N_2749,N_2662);
and U2957 (N_2957,N_2636,N_2569);
nor U2958 (N_2958,N_2534,N_2501);
nand U2959 (N_2959,N_2601,N_2647);
and U2960 (N_2960,N_2710,N_2713);
xnor U2961 (N_2961,N_2651,N_2627);
xnor U2962 (N_2962,N_2624,N_2520);
and U2963 (N_2963,N_2662,N_2668);
nand U2964 (N_2964,N_2606,N_2684);
xnor U2965 (N_2965,N_2594,N_2613);
nor U2966 (N_2966,N_2508,N_2714);
xnor U2967 (N_2967,N_2716,N_2671);
and U2968 (N_2968,N_2501,N_2585);
and U2969 (N_2969,N_2693,N_2660);
and U2970 (N_2970,N_2728,N_2524);
or U2971 (N_2971,N_2694,N_2689);
nand U2972 (N_2972,N_2511,N_2612);
xnor U2973 (N_2973,N_2702,N_2707);
xnor U2974 (N_2974,N_2546,N_2570);
and U2975 (N_2975,N_2518,N_2695);
nor U2976 (N_2976,N_2549,N_2631);
nand U2977 (N_2977,N_2505,N_2676);
nor U2978 (N_2978,N_2539,N_2512);
xnor U2979 (N_2979,N_2748,N_2726);
nor U2980 (N_2980,N_2649,N_2612);
xnor U2981 (N_2981,N_2707,N_2503);
nor U2982 (N_2982,N_2519,N_2541);
nand U2983 (N_2983,N_2722,N_2726);
or U2984 (N_2984,N_2591,N_2746);
and U2985 (N_2985,N_2678,N_2532);
xor U2986 (N_2986,N_2611,N_2719);
or U2987 (N_2987,N_2571,N_2580);
or U2988 (N_2988,N_2651,N_2613);
nand U2989 (N_2989,N_2510,N_2630);
nand U2990 (N_2990,N_2626,N_2639);
and U2991 (N_2991,N_2654,N_2693);
xor U2992 (N_2992,N_2500,N_2693);
nand U2993 (N_2993,N_2527,N_2746);
and U2994 (N_2994,N_2729,N_2614);
and U2995 (N_2995,N_2700,N_2544);
and U2996 (N_2996,N_2669,N_2504);
xnor U2997 (N_2997,N_2543,N_2733);
or U2998 (N_2998,N_2643,N_2653);
and U2999 (N_2999,N_2507,N_2516);
or U3000 (N_3000,N_2776,N_2782);
nor U3001 (N_3001,N_2941,N_2821);
or U3002 (N_3002,N_2789,N_2867);
xnor U3003 (N_3003,N_2940,N_2804);
nand U3004 (N_3004,N_2755,N_2797);
or U3005 (N_3005,N_2953,N_2920);
xnor U3006 (N_3006,N_2904,N_2838);
nand U3007 (N_3007,N_2849,N_2769);
nor U3008 (N_3008,N_2894,N_2842);
and U3009 (N_3009,N_2937,N_2784);
nor U3010 (N_3010,N_2989,N_2929);
or U3011 (N_3011,N_2936,N_2913);
nor U3012 (N_3012,N_2990,N_2974);
and U3013 (N_3013,N_2970,N_2877);
xor U3014 (N_3014,N_2779,N_2865);
xor U3015 (N_3015,N_2973,N_2983);
and U3016 (N_3016,N_2787,N_2984);
xor U3017 (N_3017,N_2793,N_2889);
nor U3018 (N_3018,N_2902,N_2852);
or U3019 (N_3019,N_2949,N_2854);
nor U3020 (N_3020,N_2806,N_2764);
nor U3021 (N_3021,N_2795,N_2843);
xnor U3022 (N_3022,N_2810,N_2977);
or U3023 (N_3023,N_2911,N_2816);
xnor U3024 (N_3024,N_2813,N_2909);
nor U3025 (N_3025,N_2905,N_2908);
xor U3026 (N_3026,N_2979,N_2995);
or U3027 (N_3027,N_2982,N_2765);
nand U3028 (N_3028,N_2863,N_2963);
xnor U3029 (N_3029,N_2895,N_2762);
nor U3030 (N_3030,N_2956,N_2967);
or U3031 (N_3031,N_2899,N_2759);
or U3032 (N_3032,N_2955,N_2850);
or U3033 (N_3033,N_2896,N_2772);
xor U3034 (N_3034,N_2845,N_2825);
and U3035 (N_3035,N_2968,N_2777);
or U3036 (N_3036,N_2976,N_2946);
nor U3037 (N_3037,N_2785,N_2800);
and U3038 (N_3038,N_2954,N_2809);
nand U3039 (N_3039,N_2752,N_2786);
nor U3040 (N_3040,N_2917,N_2866);
and U3041 (N_3041,N_2798,N_2882);
xnor U3042 (N_3042,N_2751,N_2872);
nor U3043 (N_3043,N_2829,N_2888);
xnor U3044 (N_3044,N_2932,N_2774);
nor U3045 (N_3045,N_2808,N_2942);
or U3046 (N_3046,N_2883,N_2818);
or U3047 (N_3047,N_2966,N_2837);
and U3048 (N_3048,N_2969,N_2910);
xor U3049 (N_3049,N_2851,N_2830);
or U3050 (N_3050,N_2938,N_2887);
nand U3051 (N_3051,N_2961,N_2934);
nand U3052 (N_3052,N_2931,N_2870);
nand U3053 (N_3053,N_2900,N_2750);
nor U3054 (N_3054,N_2815,N_2844);
nor U3055 (N_3055,N_2812,N_2988);
nor U3056 (N_3056,N_2763,N_2986);
and U3057 (N_3057,N_2848,N_2879);
nor U3058 (N_3058,N_2791,N_2880);
xnor U3059 (N_3059,N_2805,N_2835);
nand U3060 (N_3060,N_2897,N_2760);
xor U3061 (N_3061,N_2853,N_2871);
and U3062 (N_3062,N_2839,N_2939);
and U3063 (N_3063,N_2757,N_2881);
or U3064 (N_3064,N_2778,N_2901);
nand U3065 (N_3065,N_2891,N_2826);
or U3066 (N_3066,N_2788,N_2962);
nand U3067 (N_3067,N_2773,N_2916);
nand U3068 (N_3068,N_2822,N_2978);
nor U3069 (N_3069,N_2952,N_2903);
nand U3070 (N_3070,N_2907,N_2921);
nand U3071 (N_3071,N_2975,N_2998);
nor U3072 (N_3072,N_2875,N_2861);
and U3073 (N_3073,N_2958,N_2964);
nor U3074 (N_3074,N_2832,N_2768);
and U3075 (N_3075,N_2796,N_2912);
nand U3076 (N_3076,N_2981,N_2925);
xnor U3077 (N_3077,N_2802,N_2756);
nand U3078 (N_3078,N_2948,N_2935);
and U3079 (N_3079,N_2886,N_2824);
and U3080 (N_3080,N_2766,N_2943);
nor U3081 (N_3081,N_2801,N_2928);
and U3082 (N_3082,N_2933,N_2914);
nand U3083 (N_3083,N_2987,N_2930);
and U3084 (N_3084,N_2820,N_2873);
and U3085 (N_3085,N_2792,N_2924);
and U3086 (N_3086,N_2775,N_2951);
nand U3087 (N_3087,N_2959,N_2864);
xor U3088 (N_3088,N_2817,N_2996);
xnor U3089 (N_3089,N_2836,N_2999);
and U3090 (N_3090,N_2980,N_2950);
nand U3091 (N_3091,N_2831,N_2770);
and U3092 (N_3092,N_2834,N_2868);
nor U3093 (N_3093,N_2927,N_2919);
xnor U3094 (N_3094,N_2926,N_2827);
xor U3095 (N_3095,N_2858,N_2790);
and U3096 (N_3096,N_2960,N_2957);
and U3097 (N_3097,N_2833,N_2819);
xor U3098 (N_3098,N_2754,N_2890);
and U3099 (N_3099,N_2965,N_2893);
or U3100 (N_3100,N_2811,N_2856);
xnor U3101 (N_3101,N_2898,N_2972);
and U3102 (N_3102,N_2753,N_2918);
or U3103 (N_3103,N_2885,N_2876);
xor U3104 (N_3104,N_2767,N_2771);
and U3105 (N_3105,N_2761,N_2857);
nand U3106 (N_3106,N_2922,N_2781);
or U3107 (N_3107,N_2993,N_2780);
and U3108 (N_3108,N_2991,N_2859);
nand U3109 (N_3109,N_2803,N_2915);
nand U3110 (N_3110,N_2814,N_2846);
nor U3111 (N_3111,N_2874,N_2878);
nor U3112 (N_3112,N_2799,N_2841);
and U3113 (N_3113,N_2862,N_2992);
xnor U3114 (N_3114,N_2860,N_2947);
xor U3115 (N_3115,N_2906,N_2994);
or U3116 (N_3116,N_2823,N_2945);
nand U3117 (N_3117,N_2985,N_2997);
or U3118 (N_3118,N_2892,N_2944);
nand U3119 (N_3119,N_2847,N_2783);
nor U3120 (N_3120,N_2840,N_2794);
nor U3121 (N_3121,N_2807,N_2869);
or U3122 (N_3122,N_2828,N_2923);
xor U3123 (N_3123,N_2884,N_2855);
and U3124 (N_3124,N_2971,N_2758);
xnor U3125 (N_3125,N_2916,N_2866);
xnor U3126 (N_3126,N_2872,N_2860);
xor U3127 (N_3127,N_2974,N_2889);
and U3128 (N_3128,N_2860,N_2950);
nand U3129 (N_3129,N_2868,N_2826);
and U3130 (N_3130,N_2963,N_2764);
nor U3131 (N_3131,N_2951,N_2780);
nand U3132 (N_3132,N_2770,N_2892);
or U3133 (N_3133,N_2886,N_2942);
or U3134 (N_3134,N_2878,N_2796);
or U3135 (N_3135,N_2884,N_2987);
and U3136 (N_3136,N_2864,N_2991);
nand U3137 (N_3137,N_2876,N_2943);
or U3138 (N_3138,N_2788,N_2777);
and U3139 (N_3139,N_2830,N_2814);
and U3140 (N_3140,N_2988,N_2756);
and U3141 (N_3141,N_2834,N_2821);
or U3142 (N_3142,N_2919,N_2798);
nor U3143 (N_3143,N_2859,N_2834);
xor U3144 (N_3144,N_2777,N_2913);
nand U3145 (N_3145,N_2907,N_2898);
or U3146 (N_3146,N_2895,N_2951);
xor U3147 (N_3147,N_2907,N_2771);
and U3148 (N_3148,N_2938,N_2772);
nor U3149 (N_3149,N_2950,N_2890);
or U3150 (N_3150,N_2923,N_2907);
nand U3151 (N_3151,N_2776,N_2778);
nand U3152 (N_3152,N_2796,N_2964);
nand U3153 (N_3153,N_2946,N_2926);
and U3154 (N_3154,N_2997,N_2828);
xor U3155 (N_3155,N_2938,N_2940);
xnor U3156 (N_3156,N_2998,N_2799);
and U3157 (N_3157,N_2861,N_2824);
or U3158 (N_3158,N_2755,N_2851);
nor U3159 (N_3159,N_2811,N_2760);
nand U3160 (N_3160,N_2836,N_2879);
nor U3161 (N_3161,N_2767,N_2990);
nor U3162 (N_3162,N_2909,N_2828);
nand U3163 (N_3163,N_2832,N_2756);
nor U3164 (N_3164,N_2869,N_2808);
nor U3165 (N_3165,N_2795,N_2915);
nor U3166 (N_3166,N_2792,N_2877);
nor U3167 (N_3167,N_2933,N_2957);
xnor U3168 (N_3168,N_2953,N_2971);
or U3169 (N_3169,N_2979,N_2976);
nor U3170 (N_3170,N_2771,N_2896);
nor U3171 (N_3171,N_2762,N_2850);
nand U3172 (N_3172,N_2818,N_2896);
xnor U3173 (N_3173,N_2769,N_2842);
nor U3174 (N_3174,N_2947,N_2991);
or U3175 (N_3175,N_2765,N_2890);
or U3176 (N_3176,N_2854,N_2819);
and U3177 (N_3177,N_2754,N_2826);
and U3178 (N_3178,N_2952,N_2823);
xnor U3179 (N_3179,N_2931,N_2855);
and U3180 (N_3180,N_2911,N_2781);
xor U3181 (N_3181,N_2820,N_2969);
or U3182 (N_3182,N_2921,N_2965);
nor U3183 (N_3183,N_2954,N_2915);
nor U3184 (N_3184,N_2897,N_2774);
nand U3185 (N_3185,N_2935,N_2846);
xor U3186 (N_3186,N_2751,N_2939);
xor U3187 (N_3187,N_2902,N_2890);
and U3188 (N_3188,N_2857,N_2841);
nand U3189 (N_3189,N_2906,N_2892);
nor U3190 (N_3190,N_2772,N_2793);
nor U3191 (N_3191,N_2897,N_2971);
nor U3192 (N_3192,N_2934,N_2999);
and U3193 (N_3193,N_2760,N_2981);
and U3194 (N_3194,N_2964,N_2869);
nor U3195 (N_3195,N_2784,N_2761);
xor U3196 (N_3196,N_2822,N_2910);
nand U3197 (N_3197,N_2842,N_2945);
xor U3198 (N_3198,N_2994,N_2887);
nand U3199 (N_3199,N_2893,N_2868);
xor U3200 (N_3200,N_2842,N_2752);
xor U3201 (N_3201,N_2769,N_2827);
or U3202 (N_3202,N_2826,N_2854);
and U3203 (N_3203,N_2985,N_2861);
or U3204 (N_3204,N_2758,N_2986);
xnor U3205 (N_3205,N_2877,N_2957);
or U3206 (N_3206,N_2805,N_2826);
and U3207 (N_3207,N_2776,N_2770);
xor U3208 (N_3208,N_2953,N_2840);
nor U3209 (N_3209,N_2978,N_2998);
xnor U3210 (N_3210,N_2880,N_2773);
and U3211 (N_3211,N_2827,N_2750);
or U3212 (N_3212,N_2987,N_2803);
nor U3213 (N_3213,N_2859,N_2908);
or U3214 (N_3214,N_2911,N_2904);
and U3215 (N_3215,N_2760,N_2932);
nor U3216 (N_3216,N_2900,N_2975);
and U3217 (N_3217,N_2936,N_2854);
xor U3218 (N_3218,N_2769,N_2992);
xor U3219 (N_3219,N_2976,N_2770);
nor U3220 (N_3220,N_2984,N_2821);
nand U3221 (N_3221,N_2757,N_2954);
nor U3222 (N_3222,N_2960,N_2986);
nor U3223 (N_3223,N_2774,N_2838);
nand U3224 (N_3224,N_2957,N_2981);
nor U3225 (N_3225,N_2850,N_2892);
or U3226 (N_3226,N_2849,N_2937);
nor U3227 (N_3227,N_2885,N_2889);
nand U3228 (N_3228,N_2763,N_2985);
or U3229 (N_3229,N_2883,N_2946);
or U3230 (N_3230,N_2948,N_2884);
nor U3231 (N_3231,N_2833,N_2826);
nor U3232 (N_3232,N_2997,N_2755);
xnor U3233 (N_3233,N_2854,N_2802);
nand U3234 (N_3234,N_2802,N_2811);
nand U3235 (N_3235,N_2821,N_2850);
nor U3236 (N_3236,N_2965,N_2941);
nor U3237 (N_3237,N_2848,N_2897);
nand U3238 (N_3238,N_2989,N_2846);
and U3239 (N_3239,N_2949,N_2947);
nand U3240 (N_3240,N_2858,N_2929);
or U3241 (N_3241,N_2823,N_2915);
and U3242 (N_3242,N_2966,N_2996);
nor U3243 (N_3243,N_2842,N_2879);
or U3244 (N_3244,N_2945,N_2953);
xnor U3245 (N_3245,N_2963,N_2935);
nor U3246 (N_3246,N_2939,N_2830);
or U3247 (N_3247,N_2773,N_2986);
or U3248 (N_3248,N_2967,N_2878);
nand U3249 (N_3249,N_2859,N_2857);
nand U3250 (N_3250,N_3105,N_3101);
nor U3251 (N_3251,N_3085,N_3029);
nand U3252 (N_3252,N_3248,N_3220);
or U3253 (N_3253,N_3201,N_3135);
nand U3254 (N_3254,N_3046,N_3145);
and U3255 (N_3255,N_3073,N_3215);
nor U3256 (N_3256,N_3140,N_3212);
and U3257 (N_3257,N_3130,N_3244);
and U3258 (N_3258,N_3142,N_3243);
nand U3259 (N_3259,N_3185,N_3177);
nand U3260 (N_3260,N_3088,N_3053);
or U3261 (N_3261,N_3058,N_3182);
nand U3262 (N_3262,N_3242,N_3178);
xor U3263 (N_3263,N_3056,N_3028);
and U3264 (N_3264,N_3200,N_3080);
and U3265 (N_3265,N_3231,N_3246);
and U3266 (N_3266,N_3203,N_3186);
xnor U3267 (N_3267,N_3143,N_3147);
nor U3268 (N_3268,N_3019,N_3159);
and U3269 (N_3269,N_3137,N_3075);
xnor U3270 (N_3270,N_3086,N_3059);
nor U3271 (N_3271,N_3035,N_3038);
nor U3272 (N_3272,N_3079,N_3025);
and U3273 (N_3273,N_3037,N_3115);
nor U3274 (N_3274,N_3221,N_3217);
and U3275 (N_3275,N_3240,N_3114);
and U3276 (N_3276,N_3012,N_3005);
and U3277 (N_3277,N_3117,N_3168);
nand U3278 (N_3278,N_3112,N_3009);
nor U3279 (N_3279,N_3083,N_3184);
xor U3280 (N_3280,N_3237,N_3131);
nand U3281 (N_3281,N_3069,N_3097);
xnor U3282 (N_3282,N_3156,N_3162);
and U3283 (N_3283,N_3107,N_3011);
nor U3284 (N_3284,N_3123,N_3074);
nand U3285 (N_3285,N_3048,N_3062);
nand U3286 (N_3286,N_3093,N_3090);
xnor U3287 (N_3287,N_3022,N_3064);
or U3288 (N_3288,N_3042,N_3146);
and U3289 (N_3289,N_3081,N_3227);
xor U3290 (N_3290,N_3078,N_3113);
or U3291 (N_3291,N_3096,N_3171);
nand U3292 (N_3292,N_3045,N_3180);
or U3293 (N_3293,N_3154,N_3136);
and U3294 (N_3294,N_3160,N_3172);
nand U3295 (N_3295,N_3132,N_3066);
xnor U3296 (N_3296,N_3014,N_3095);
and U3297 (N_3297,N_3148,N_3077);
xnor U3298 (N_3298,N_3104,N_3108);
and U3299 (N_3299,N_3099,N_3170);
or U3300 (N_3300,N_3175,N_3229);
nand U3301 (N_3301,N_3213,N_3034);
nand U3302 (N_3302,N_3234,N_3166);
xor U3303 (N_3303,N_3210,N_3043);
or U3304 (N_3304,N_3106,N_3249);
xor U3305 (N_3305,N_3188,N_3094);
xnor U3306 (N_3306,N_3223,N_3233);
nand U3307 (N_3307,N_3225,N_3070);
xnor U3308 (N_3308,N_3015,N_3026);
and U3309 (N_3309,N_3129,N_3193);
nand U3310 (N_3310,N_3087,N_3236);
xnor U3311 (N_3311,N_3205,N_3039);
nor U3312 (N_3312,N_3003,N_3209);
xor U3313 (N_3313,N_3001,N_3006);
and U3314 (N_3314,N_3152,N_3157);
xor U3315 (N_3315,N_3084,N_3247);
or U3316 (N_3316,N_3102,N_3000);
and U3317 (N_3317,N_3007,N_3052);
or U3318 (N_3318,N_3181,N_3230);
nand U3319 (N_3319,N_3120,N_3133);
nand U3320 (N_3320,N_3050,N_3226);
xor U3321 (N_3321,N_3020,N_3055);
xor U3322 (N_3322,N_3161,N_3224);
xnor U3323 (N_3323,N_3118,N_3030);
xnor U3324 (N_3324,N_3071,N_3004);
and U3325 (N_3325,N_3091,N_3061);
nor U3326 (N_3326,N_3206,N_3036);
nand U3327 (N_3327,N_3040,N_3109);
and U3328 (N_3328,N_3169,N_3195);
and U3329 (N_3329,N_3235,N_3128);
xor U3330 (N_3330,N_3150,N_3239);
or U3331 (N_3331,N_3187,N_3089);
nand U3332 (N_3332,N_3174,N_3183);
nor U3333 (N_3333,N_3044,N_3057);
or U3334 (N_3334,N_3241,N_3228);
xnor U3335 (N_3335,N_3010,N_3158);
and U3336 (N_3336,N_3119,N_3153);
and U3337 (N_3337,N_3068,N_3138);
nand U3338 (N_3338,N_3067,N_3196);
and U3339 (N_3339,N_3127,N_3031);
nor U3340 (N_3340,N_3121,N_3060);
xor U3341 (N_3341,N_3033,N_3222);
nor U3342 (N_3342,N_3092,N_3013);
or U3343 (N_3343,N_3041,N_3023);
and U3344 (N_3344,N_3167,N_3173);
or U3345 (N_3345,N_3054,N_3207);
nand U3346 (N_3346,N_3192,N_3144);
xor U3347 (N_3347,N_3149,N_3021);
nor U3348 (N_3348,N_3076,N_3111);
nor U3349 (N_3349,N_3082,N_3163);
xor U3350 (N_3350,N_3072,N_3194);
or U3351 (N_3351,N_3063,N_3126);
xor U3352 (N_3352,N_3199,N_3134);
and U3353 (N_3353,N_3179,N_3103);
nor U3354 (N_3354,N_3110,N_3202);
xnor U3355 (N_3355,N_3245,N_3139);
or U3356 (N_3356,N_3219,N_3155);
or U3357 (N_3357,N_3027,N_3100);
nor U3358 (N_3358,N_3165,N_3098);
and U3359 (N_3359,N_3032,N_3214);
xnor U3360 (N_3360,N_3008,N_3191);
and U3361 (N_3361,N_3116,N_3208);
nor U3362 (N_3362,N_3216,N_3218);
and U3363 (N_3363,N_3232,N_3002);
or U3364 (N_3364,N_3238,N_3151);
nor U3365 (N_3365,N_3122,N_3164);
nor U3366 (N_3366,N_3024,N_3017);
xnor U3367 (N_3367,N_3211,N_3016);
nor U3368 (N_3368,N_3176,N_3049);
xor U3369 (N_3369,N_3190,N_3189);
nor U3370 (N_3370,N_3197,N_3047);
nor U3371 (N_3371,N_3141,N_3198);
xnor U3372 (N_3372,N_3018,N_3051);
nand U3373 (N_3373,N_3125,N_3065);
xnor U3374 (N_3374,N_3204,N_3124);
or U3375 (N_3375,N_3009,N_3201);
nor U3376 (N_3376,N_3173,N_3044);
or U3377 (N_3377,N_3228,N_3081);
nand U3378 (N_3378,N_3027,N_3046);
xnor U3379 (N_3379,N_3027,N_3105);
nand U3380 (N_3380,N_3222,N_3098);
nand U3381 (N_3381,N_3119,N_3053);
nand U3382 (N_3382,N_3019,N_3171);
nor U3383 (N_3383,N_3184,N_3024);
or U3384 (N_3384,N_3079,N_3122);
xor U3385 (N_3385,N_3147,N_3197);
xor U3386 (N_3386,N_3156,N_3247);
nor U3387 (N_3387,N_3122,N_3058);
xnor U3388 (N_3388,N_3139,N_3134);
and U3389 (N_3389,N_3238,N_3179);
or U3390 (N_3390,N_3023,N_3002);
nor U3391 (N_3391,N_3039,N_3237);
nor U3392 (N_3392,N_3248,N_3039);
xnor U3393 (N_3393,N_3091,N_3050);
nor U3394 (N_3394,N_3132,N_3125);
xnor U3395 (N_3395,N_3244,N_3246);
or U3396 (N_3396,N_3200,N_3030);
or U3397 (N_3397,N_3029,N_3230);
or U3398 (N_3398,N_3173,N_3156);
xor U3399 (N_3399,N_3095,N_3185);
xnor U3400 (N_3400,N_3155,N_3209);
and U3401 (N_3401,N_3161,N_3088);
or U3402 (N_3402,N_3033,N_3208);
nand U3403 (N_3403,N_3071,N_3158);
and U3404 (N_3404,N_3065,N_3053);
nand U3405 (N_3405,N_3000,N_3025);
or U3406 (N_3406,N_3204,N_3077);
and U3407 (N_3407,N_3007,N_3203);
nand U3408 (N_3408,N_3187,N_3003);
nand U3409 (N_3409,N_3130,N_3036);
xor U3410 (N_3410,N_3227,N_3113);
and U3411 (N_3411,N_3215,N_3099);
and U3412 (N_3412,N_3163,N_3032);
or U3413 (N_3413,N_3049,N_3226);
xnor U3414 (N_3414,N_3217,N_3104);
nor U3415 (N_3415,N_3052,N_3030);
nor U3416 (N_3416,N_3064,N_3068);
or U3417 (N_3417,N_3234,N_3248);
xor U3418 (N_3418,N_3245,N_3068);
and U3419 (N_3419,N_3153,N_3126);
nand U3420 (N_3420,N_3115,N_3007);
or U3421 (N_3421,N_3087,N_3066);
and U3422 (N_3422,N_3073,N_3040);
nand U3423 (N_3423,N_3081,N_3226);
xnor U3424 (N_3424,N_3167,N_3103);
nand U3425 (N_3425,N_3115,N_3190);
nand U3426 (N_3426,N_3139,N_3086);
nand U3427 (N_3427,N_3020,N_3163);
and U3428 (N_3428,N_3141,N_3124);
nor U3429 (N_3429,N_3044,N_3149);
xnor U3430 (N_3430,N_3226,N_3036);
or U3431 (N_3431,N_3148,N_3249);
xnor U3432 (N_3432,N_3081,N_3066);
or U3433 (N_3433,N_3086,N_3035);
and U3434 (N_3434,N_3118,N_3082);
xor U3435 (N_3435,N_3013,N_3224);
xor U3436 (N_3436,N_3151,N_3230);
or U3437 (N_3437,N_3004,N_3024);
nor U3438 (N_3438,N_3044,N_3130);
and U3439 (N_3439,N_3013,N_3117);
and U3440 (N_3440,N_3203,N_3012);
nand U3441 (N_3441,N_3142,N_3151);
xor U3442 (N_3442,N_3150,N_3005);
and U3443 (N_3443,N_3180,N_3155);
xnor U3444 (N_3444,N_3240,N_3076);
and U3445 (N_3445,N_3073,N_3194);
nor U3446 (N_3446,N_3156,N_3042);
nor U3447 (N_3447,N_3220,N_3097);
nand U3448 (N_3448,N_3219,N_3066);
xnor U3449 (N_3449,N_3209,N_3158);
or U3450 (N_3450,N_3234,N_3159);
nor U3451 (N_3451,N_3214,N_3076);
nor U3452 (N_3452,N_3234,N_3170);
xor U3453 (N_3453,N_3027,N_3132);
nand U3454 (N_3454,N_3247,N_3244);
nand U3455 (N_3455,N_3187,N_3137);
xnor U3456 (N_3456,N_3192,N_3170);
and U3457 (N_3457,N_3032,N_3079);
or U3458 (N_3458,N_3161,N_3059);
or U3459 (N_3459,N_3123,N_3138);
xor U3460 (N_3460,N_3073,N_3014);
nor U3461 (N_3461,N_3124,N_3069);
xnor U3462 (N_3462,N_3089,N_3247);
or U3463 (N_3463,N_3128,N_3046);
or U3464 (N_3464,N_3061,N_3206);
and U3465 (N_3465,N_3210,N_3162);
nor U3466 (N_3466,N_3236,N_3186);
or U3467 (N_3467,N_3241,N_3204);
xnor U3468 (N_3468,N_3145,N_3042);
nor U3469 (N_3469,N_3158,N_3077);
xor U3470 (N_3470,N_3245,N_3046);
and U3471 (N_3471,N_3245,N_3175);
xor U3472 (N_3472,N_3121,N_3125);
xor U3473 (N_3473,N_3227,N_3245);
nand U3474 (N_3474,N_3014,N_3002);
and U3475 (N_3475,N_3209,N_3038);
and U3476 (N_3476,N_3014,N_3048);
nand U3477 (N_3477,N_3046,N_3097);
nand U3478 (N_3478,N_3232,N_3045);
and U3479 (N_3479,N_3115,N_3095);
xor U3480 (N_3480,N_3037,N_3139);
nor U3481 (N_3481,N_3173,N_3175);
nor U3482 (N_3482,N_3183,N_3085);
nor U3483 (N_3483,N_3247,N_3192);
and U3484 (N_3484,N_3054,N_3151);
nor U3485 (N_3485,N_3038,N_3181);
xnor U3486 (N_3486,N_3134,N_3193);
nor U3487 (N_3487,N_3006,N_3161);
xnor U3488 (N_3488,N_3134,N_3155);
and U3489 (N_3489,N_3183,N_3186);
and U3490 (N_3490,N_3174,N_3161);
nor U3491 (N_3491,N_3182,N_3108);
nor U3492 (N_3492,N_3186,N_3188);
and U3493 (N_3493,N_3089,N_3212);
or U3494 (N_3494,N_3140,N_3191);
or U3495 (N_3495,N_3152,N_3171);
nor U3496 (N_3496,N_3017,N_3191);
nand U3497 (N_3497,N_3103,N_3133);
xnor U3498 (N_3498,N_3129,N_3060);
and U3499 (N_3499,N_3058,N_3044);
xor U3500 (N_3500,N_3409,N_3395);
nor U3501 (N_3501,N_3451,N_3349);
or U3502 (N_3502,N_3412,N_3354);
and U3503 (N_3503,N_3391,N_3317);
and U3504 (N_3504,N_3393,N_3490);
nand U3505 (N_3505,N_3357,N_3254);
nand U3506 (N_3506,N_3484,N_3432);
nand U3507 (N_3507,N_3454,N_3491);
nor U3508 (N_3508,N_3399,N_3346);
xnor U3509 (N_3509,N_3355,N_3440);
nand U3510 (N_3510,N_3333,N_3278);
and U3511 (N_3511,N_3318,N_3381);
and U3512 (N_3512,N_3398,N_3289);
and U3513 (N_3513,N_3387,N_3266);
and U3514 (N_3514,N_3340,N_3385);
or U3515 (N_3515,N_3353,N_3262);
nor U3516 (N_3516,N_3389,N_3356);
and U3517 (N_3517,N_3388,N_3281);
and U3518 (N_3518,N_3433,N_3265);
nor U3519 (N_3519,N_3304,N_3319);
nor U3520 (N_3520,N_3397,N_3366);
nand U3521 (N_3521,N_3337,N_3445);
nand U3522 (N_3522,N_3450,N_3497);
or U3523 (N_3523,N_3256,N_3344);
or U3524 (N_3524,N_3459,N_3358);
nand U3525 (N_3525,N_3284,N_3373);
nand U3526 (N_3526,N_3331,N_3418);
xnor U3527 (N_3527,N_3296,N_3255);
nor U3528 (N_3528,N_3253,N_3477);
xor U3529 (N_3529,N_3458,N_3407);
xnor U3530 (N_3530,N_3309,N_3400);
or U3531 (N_3531,N_3292,N_3476);
or U3532 (N_3532,N_3367,N_3314);
nor U3533 (N_3533,N_3290,N_3430);
nand U3534 (N_3534,N_3257,N_3493);
and U3535 (N_3535,N_3321,N_3371);
xor U3536 (N_3536,N_3287,N_3428);
and U3537 (N_3537,N_3457,N_3377);
xnor U3538 (N_3538,N_3364,N_3359);
nand U3539 (N_3539,N_3335,N_3487);
and U3540 (N_3540,N_3456,N_3495);
or U3541 (N_3541,N_3452,N_3351);
nor U3542 (N_3542,N_3423,N_3376);
or U3543 (N_3543,N_3481,N_3414);
and U3544 (N_3544,N_3406,N_3302);
or U3545 (N_3545,N_3444,N_3369);
nor U3546 (N_3546,N_3384,N_3269);
xnor U3547 (N_3547,N_3489,N_3442);
nand U3548 (N_3548,N_3390,N_3485);
and U3549 (N_3549,N_3310,N_3473);
nor U3550 (N_3550,N_3275,N_3350);
nand U3551 (N_3551,N_3267,N_3261);
or U3552 (N_3552,N_3436,N_3362);
xor U3553 (N_3553,N_3453,N_3424);
and U3554 (N_3554,N_3330,N_3264);
nor U3555 (N_3555,N_3435,N_3498);
nor U3556 (N_3556,N_3401,N_3348);
xor U3557 (N_3557,N_3417,N_3271);
nand U3558 (N_3558,N_3250,N_3339);
and U3559 (N_3559,N_3404,N_3494);
xnor U3560 (N_3560,N_3394,N_3375);
nor U3561 (N_3561,N_3480,N_3336);
or U3562 (N_3562,N_3322,N_3426);
or U3563 (N_3563,N_3251,N_3268);
nor U3564 (N_3564,N_3293,N_3294);
or U3565 (N_3565,N_3386,N_3374);
and U3566 (N_3566,N_3334,N_3478);
or U3567 (N_3567,N_3380,N_3338);
nor U3568 (N_3568,N_3298,N_3365);
or U3569 (N_3569,N_3291,N_3259);
nand U3570 (N_3570,N_3443,N_3438);
or U3571 (N_3571,N_3474,N_3370);
nand U3572 (N_3572,N_3465,N_3499);
xor U3573 (N_3573,N_3408,N_3420);
or U3574 (N_3574,N_3496,N_3263);
nor U3575 (N_3575,N_3448,N_3411);
and U3576 (N_3576,N_3295,N_3475);
nand U3577 (N_3577,N_3460,N_3311);
nor U3578 (N_3578,N_3469,N_3361);
or U3579 (N_3579,N_3482,N_3382);
nor U3580 (N_3580,N_3461,N_3320);
and U3581 (N_3581,N_3383,N_3329);
nand U3582 (N_3582,N_3270,N_3441);
nor U3583 (N_3583,N_3300,N_3286);
and U3584 (N_3584,N_3328,N_3486);
or U3585 (N_3585,N_3280,N_3468);
xor U3586 (N_3586,N_3363,N_3277);
nand U3587 (N_3587,N_3252,N_3429);
and U3588 (N_3588,N_3396,N_3313);
or U3589 (N_3589,N_3431,N_3274);
xnor U3590 (N_3590,N_3368,N_3297);
nor U3591 (N_3591,N_3422,N_3416);
xnor U3592 (N_3592,N_3288,N_3343);
xnor U3593 (N_3593,N_3312,N_3392);
and U3594 (N_3594,N_3299,N_3303);
and U3595 (N_3595,N_3325,N_3427);
nand U3596 (N_3596,N_3455,N_3446);
nand U3597 (N_3597,N_3347,N_3282);
xor U3598 (N_3598,N_3324,N_3372);
nor U3599 (N_3599,N_3352,N_3308);
or U3600 (N_3600,N_3447,N_3316);
xnor U3601 (N_3601,N_3379,N_3327);
and U3602 (N_3602,N_3403,N_3273);
or U3603 (N_3603,N_3276,N_3315);
and U3604 (N_3604,N_3345,N_3402);
xnor U3605 (N_3605,N_3260,N_3466);
or U3606 (N_3606,N_3305,N_3439);
nor U3607 (N_3607,N_3470,N_3483);
nand U3608 (N_3608,N_3463,N_3479);
xor U3609 (N_3609,N_3421,N_3471);
xnor U3610 (N_3610,N_3413,N_3415);
nor U3611 (N_3611,N_3462,N_3492);
nor U3612 (N_3612,N_3467,N_3434);
or U3613 (N_3613,N_3488,N_3341);
nand U3614 (N_3614,N_3285,N_3464);
and U3615 (N_3615,N_3405,N_3258);
xnor U3616 (N_3616,N_3332,N_3301);
xor U3617 (N_3617,N_3360,N_3283);
or U3618 (N_3618,N_3279,N_3306);
or U3619 (N_3619,N_3410,N_3449);
xor U3620 (N_3620,N_3419,N_3425);
and U3621 (N_3621,N_3472,N_3378);
nor U3622 (N_3622,N_3326,N_3437);
nor U3623 (N_3623,N_3272,N_3323);
and U3624 (N_3624,N_3342,N_3307);
or U3625 (N_3625,N_3343,N_3348);
nand U3626 (N_3626,N_3417,N_3299);
nor U3627 (N_3627,N_3496,N_3477);
xnor U3628 (N_3628,N_3426,N_3449);
xor U3629 (N_3629,N_3356,N_3374);
and U3630 (N_3630,N_3404,N_3320);
nor U3631 (N_3631,N_3267,N_3402);
nand U3632 (N_3632,N_3433,N_3405);
nand U3633 (N_3633,N_3319,N_3267);
xor U3634 (N_3634,N_3271,N_3312);
xor U3635 (N_3635,N_3334,N_3401);
xor U3636 (N_3636,N_3337,N_3385);
xnor U3637 (N_3637,N_3486,N_3309);
nand U3638 (N_3638,N_3381,N_3346);
and U3639 (N_3639,N_3404,N_3379);
nand U3640 (N_3640,N_3475,N_3300);
or U3641 (N_3641,N_3268,N_3390);
nand U3642 (N_3642,N_3387,N_3485);
or U3643 (N_3643,N_3360,N_3386);
nand U3644 (N_3644,N_3394,N_3417);
or U3645 (N_3645,N_3389,N_3375);
nor U3646 (N_3646,N_3350,N_3491);
nand U3647 (N_3647,N_3325,N_3254);
or U3648 (N_3648,N_3481,N_3385);
and U3649 (N_3649,N_3486,N_3277);
and U3650 (N_3650,N_3443,N_3345);
nand U3651 (N_3651,N_3272,N_3463);
xnor U3652 (N_3652,N_3498,N_3374);
and U3653 (N_3653,N_3338,N_3458);
or U3654 (N_3654,N_3486,N_3410);
xor U3655 (N_3655,N_3444,N_3425);
xnor U3656 (N_3656,N_3411,N_3490);
and U3657 (N_3657,N_3357,N_3497);
or U3658 (N_3658,N_3344,N_3265);
nor U3659 (N_3659,N_3444,N_3279);
and U3660 (N_3660,N_3430,N_3454);
xnor U3661 (N_3661,N_3442,N_3388);
or U3662 (N_3662,N_3494,N_3361);
nand U3663 (N_3663,N_3455,N_3252);
nand U3664 (N_3664,N_3385,N_3496);
nand U3665 (N_3665,N_3310,N_3366);
nand U3666 (N_3666,N_3385,N_3270);
or U3667 (N_3667,N_3479,N_3493);
xnor U3668 (N_3668,N_3250,N_3309);
or U3669 (N_3669,N_3367,N_3419);
nand U3670 (N_3670,N_3492,N_3321);
xor U3671 (N_3671,N_3427,N_3397);
nand U3672 (N_3672,N_3337,N_3487);
or U3673 (N_3673,N_3470,N_3313);
nand U3674 (N_3674,N_3334,N_3279);
xor U3675 (N_3675,N_3392,N_3385);
or U3676 (N_3676,N_3301,N_3380);
or U3677 (N_3677,N_3284,N_3254);
nand U3678 (N_3678,N_3266,N_3306);
xor U3679 (N_3679,N_3353,N_3256);
and U3680 (N_3680,N_3361,N_3369);
nand U3681 (N_3681,N_3368,N_3434);
nor U3682 (N_3682,N_3396,N_3348);
xor U3683 (N_3683,N_3286,N_3394);
and U3684 (N_3684,N_3483,N_3265);
xnor U3685 (N_3685,N_3395,N_3287);
nand U3686 (N_3686,N_3411,N_3470);
nand U3687 (N_3687,N_3301,N_3309);
nand U3688 (N_3688,N_3396,N_3468);
xnor U3689 (N_3689,N_3386,N_3421);
xor U3690 (N_3690,N_3368,N_3488);
and U3691 (N_3691,N_3282,N_3463);
and U3692 (N_3692,N_3251,N_3309);
and U3693 (N_3693,N_3352,N_3294);
or U3694 (N_3694,N_3358,N_3386);
xnor U3695 (N_3695,N_3351,N_3461);
nor U3696 (N_3696,N_3313,N_3304);
xor U3697 (N_3697,N_3449,N_3458);
or U3698 (N_3698,N_3315,N_3474);
nand U3699 (N_3699,N_3334,N_3455);
and U3700 (N_3700,N_3300,N_3379);
xnor U3701 (N_3701,N_3287,N_3415);
nor U3702 (N_3702,N_3428,N_3430);
nor U3703 (N_3703,N_3327,N_3302);
xnor U3704 (N_3704,N_3465,N_3291);
and U3705 (N_3705,N_3290,N_3391);
nand U3706 (N_3706,N_3348,N_3282);
or U3707 (N_3707,N_3292,N_3444);
xor U3708 (N_3708,N_3341,N_3330);
nand U3709 (N_3709,N_3327,N_3400);
nor U3710 (N_3710,N_3324,N_3452);
or U3711 (N_3711,N_3275,N_3341);
and U3712 (N_3712,N_3388,N_3419);
xor U3713 (N_3713,N_3298,N_3393);
or U3714 (N_3714,N_3262,N_3336);
and U3715 (N_3715,N_3418,N_3338);
nor U3716 (N_3716,N_3427,N_3333);
nand U3717 (N_3717,N_3466,N_3411);
nand U3718 (N_3718,N_3392,N_3408);
and U3719 (N_3719,N_3395,N_3387);
nor U3720 (N_3720,N_3480,N_3473);
and U3721 (N_3721,N_3476,N_3491);
and U3722 (N_3722,N_3289,N_3435);
or U3723 (N_3723,N_3399,N_3435);
or U3724 (N_3724,N_3341,N_3308);
nand U3725 (N_3725,N_3338,N_3294);
nand U3726 (N_3726,N_3437,N_3460);
nand U3727 (N_3727,N_3329,N_3349);
and U3728 (N_3728,N_3358,N_3319);
nor U3729 (N_3729,N_3327,N_3278);
and U3730 (N_3730,N_3460,N_3338);
and U3731 (N_3731,N_3294,N_3407);
nor U3732 (N_3732,N_3466,N_3461);
nor U3733 (N_3733,N_3473,N_3273);
nor U3734 (N_3734,N_3425,N_3327);
nor U3735 (N_3735,N_3388,N_3396);
or U3736 (N_3736,N_3291,N_3429);
or U3737 (N_3737,N_3424,N_3498);
nand U3738 (N_3738,N_3393,N_3465);
nand U3739 (N_3739,N_3467,N_3390);
nor U3740 (N_3740,N_3409,N_3294);
and U3741 (N_3741,N_3348,N_3267);
and U3742 (N_3742,N_3312,N_3282);
xor U3743 (N_3743,N_3484,N_3414);
xor U3744 (N_3744,N_3324,N_3395);
nor U3745 (N_3745,N_3400,N_3295);
nand U3746 (N_3746,N_3437,N_3425);
nor U3747 (N_3747,N_3322,N_3476);
nand U3748 (N_3748,N_3250,N_3451);
nand U3749 (N_3749,N_3440,N_3272);
nand U3750 (N_3750,N_3726,N_3699);
xnor U3751 (N_3751,N_3654,N_3707);
nand U3752 (N_3752,N_3580,N_3607);
nand U3753 (N_3753,N_3565,N_3746);
nor U3754 (N_3754,N_3708,N_3720);
or U3755 (N_3755,N_3537,N_3506);
or U3756 (N_3756,N_3509,N_3552);
nand U3757 (N_3757,N_3557,N_3732);
xnor U3758 (N_3758,N_3717,N_3605);
or U3759 (N_3759,N_3630,N_3655);
nand U3760 (N_3760,N_3501,N_3675);
nor U3761 (N_3761,N_3520,N_3684);
or U3762 (N_3762,N_3550,N_3576);
xor U3763 (N_3763,N_3508,N_3636);
or U3764 (N_3764,N_3730,N_3621);
xnor U3765 (N_3765,N_3519,N_3690);
and U3766 (N_3766,N_3635,N_3725);
nand U3767 (N_3767,N_3568,N_3595);
nor U3768 (N_3768,N_3588,N_3504);
nand U3769 (N_3769,N_3613,N_3715);
and U3770 (N_3770,N_3656,N_3676);
and U3771 (N_3771,N_3632,N_3586);
nor U3772 (N_3772,N_3521,N_3529);
or U3773 (N_3773,N_3741,N_3693);
nor U3774 (N_3774,N_3539,N_3703);
xnor U3775 (N_3775,N_3591,N_3689);
nor U3776 (N_3776,N_3556,N_3533);
or U3777 (N_3777,N_3624,N_3625);
xnor U3778 (N_3778,N_3728,N_3634);
nor U3779 (N_3779,N_3640,N_3679);
or U3780 (N_3780,N_3695,N_3709);
and U3781 (N_3781,N_3513,N_3734);
nor U3782 (N_3782,N_3582,N_3604);
and U3783 (N_3783,N_3573,N_3677);
nand U3784 (N_3784,N_3596,N_3545);
xnor U3785 (N_3785,N_3618,N_3633);
nor U3786 (N_3786,N_3691,N_3548);
xor U3787 (N_3787,N_3516,N_3648);
nand U3788 (N_3788,N_3608,N_3590);
nand U3789 (N_3789,N_3645,N_3569);
xor U3790 (N_3790,N_3716,N_3531);
nor U3791 (N_3791,N_3571,N_3731);
nor U3792 (N_3792,N_3665,N_3502);
and U3793 (N_3793,N_3577,N_3535);
nand U3794 (N_3794,N_3579,N_3515);
or U3795 (N_3795,N_3745,N_3652);
nor U3796 (N_3796,N_3628,N_3532);
xor U3797 (N_3797,N_3638,N_3574);
xnor U3798 (N_3798,N_3536,N_3743);
nor U3799 (N_3799,N_3629,N_3542);
xnor U3800 (N_3800,N_3721,N_3659);
xor U3801 (N_3801,N_3662,N_3678);
nor U3802 (N_3802,N_3553,N_3555);
nand U3803 (N_3803,N_3742,N_3503);
nor U3804 (N_3804,N_3664,N_3609);
nand U3805 (N_3805,N_3694,N_3657);
or U3806 (N_3806,N_3524,N_3674);
and U3807 (N_3807,N_3615,N_3650);
nand U3808 (N_3808,N_3583,N_3688);
or U3809 (N_3809,N_3578,N_3510);
xnor U3810 (N_3810,N_3698,N_3612);
or U3811 (N_3811,N_3701,N_3600);
nor U3812 (N_3812,N_3599,N_3670);
and U3813 (N_3813,N_3626,N_3567);
nand U3814 (N_3814,N_3623,N_3598);
nor U3815 (N_3815,N_3671,N_3666);
or U3816 (N_3816,N_3696,N_3680);
xnor U3817 (N_3817,N_3507,N_3530);
and U3818 (N_3818,N_3643,N_3668);
and U3819 (N_3819,N_3641,N_3697);
nand U3820 (N_3820,N_3683,N_3558);
and U3821 (N_3821,N_3649,N_3749);
nor U3822 (N_3822,N_3512,N_3528);
or U3823 (N_3823,N_3692,N_3594);
or U3824 (N_3824,N_3637,N_3748);
xor U3825 (N_3825,N_3733,N_3735);
xnor U3826 (N_3826,N_3744,N_3587);
and U3827 (N_3827,N_3619,N_3672);
and U3828 (N_3828,N_3718,N_3700);
xnor U3829 (N_3829,N_3727,N_3661);
or U3830 (N_3830,N_3660,N_3712);
nor U3831 (N_3831,N_3686,N_3544);
or U3832 (N_3832,N_3602,N_3517);
nor U3833 (N_3833,N_3669,N_3658);
xor U3834 (N_3834,N_3592,N_3525);
nand U3835 (N_3835,N_3570,N_3547);
and U3836 (N_3836,N_3646,N_3549);
nor U3837 (N_3837,N_3647,N_3723);
and U3838 (N_3838,N_3546,N_3706);
nor U3839 (N_3839,N_3719,N_3740);
or U3840 (N_3840,N_3747,N_3681);
and U3841 (N_3841,N_3561,N_3739);
xor U3842 (N_3842,N_3551,N_3617);
or U3843 (N_3843,N_3702,N_3610);
nor U3844 (N_3844,N_3560,N_3682);
nor U3845 (N_3845,N_3616,N_3685);
xor U3846 (N_3846,N_3713,N_3514);
or U3847 (N_3847,N_3534,N_3584);
or U3848 (N_3848,N_3663,N_3518);
nor U3849 (N_3849,N_3597,N_3620);
nor U3850 (N_3850,N_3710,N_3603);
and U3851 (N_3851,N_3614,N_3540);
xor U3852 (N_3852,N_3572,N_3736);
xor U3853 (N_3853,N_3714,N_3575);
or U3854 (N_3854,N_3500,N_3593);
nor U3855 (N_3855,N_3705,N_3639);
xnor U3856 (N_3856,N_3631,N_3704);
xnor U3857 (N_3857,N_3687,N_3563);
nand U3858 (N_3858,N_3667,N_3738);
and U3859 (N_3859,N_3722,N_3511);
nand U3860 (N_3860,N_3554,N_3526);
or U3861 (N_3861,N_3644,N_3606);
nand U3862 (N_3862,N_3562,N_3627);
nand U3863 (N_3863,N_3622,N_3653);
nand U3864 (N_3864,N_3711,N_3585);
nand U3865 (N_3865,N_3729,N_3589);
or U3866 (N_3866,N_3564,N_3523);
nor U3867 (N_3867,N_3611,N_3651);
and U3868 (N_3868,N_3541,N_3522);
and U3869 (N_3869,N_3538,N_3642);
or U3870 (N_3870,N_3543,N_3559);
nand U3871 (N_3871,N_3505,N_3601);
xnor U3872 (N_3872,N_3527,N_3737);
nand U3873 (N_3873,N_3724,N_3566);
and U3874 (N_3874,N_3673,N_3581);
xor U3875 (N_3875,N_3735,N_3506);
or U3876 (N_3876,N_3521,N_3624);
xnor U3877 (N_3877,N_3655,N_3503);
nand U3878 (N_3878,N_3538,N_3658);
xor U3879 (N_3879,N_3672,N_3528);
and U3880 (N_3880,N_3610,N_3679);
xnor U3881 (N_3881,N_3527,N_3641);
or U3882 (N_3882,N_3694,N_3696);
xor U3883 (N_3883,N_3553,N_3676);
and U3884 (N_3884,N_3524,N_3603);
or U3885 (N_3885,N_3636,N_3662);
nand U3886 (N_3886,N_3611,N_3671);
nand U3887 (N_3887,N_3502,N_3510);
or U3888 (N_3888,N_3685,N_3552);
nand U3889 (N_3889,N_3663,N_3569);
nor U3890 (N_3890,N_3590,N_3655);
xnor U3891 (N_3891,N_3585,N_3734);
nor U3892 (N_3892,N_3747,N_3603);
nand U3893 (N_3893,N_3543,N_3641);
nor U3894 (N_3894,N_3618,N_3710);
or U3895 (N_3895,N_3543,N_3735);
nand U3896 (N_3896,N_3744,N_3570);
nand U3897 (N_3897,N_3508,N_3637);
nor U3898 (N_3898,N_3736,N_3609);
xor U3899 (N_3899,N_3625,N_3537);
or U3900 (N_3900,N_3502,N_3501);
xor U3901 (N_3901,N_3739,N_3748);
xnor U3902 (N_3902,N_3588,N_3613);
xor U3903 (N_3903,N_3505,N_3648);
xor U3904 (N_3904,N_3547,N_3599);
nand U3905 (N_3905,N_3601,N_3519);
nor U3906 (N_3906,N_3650,N_3603);
nand U3907 (N_3907,N_3662,N_3531);
nand U3908 (N_3908,N_3611,N_3681);
and U3909 (N_3909,N_3655,N_3618);
xor U3910 (N_3910,N_3659,N_3562);
xnor U3911 (N_3911,N_3645,N_3748);
or U3912 (N_3912,N_3574,N_3612);
and U3913 (N_3913,N_3644,N_3540);
and U3914 (N_3914,N_3680,N_3502);
or U3915 (N_3915,N_3672,N_3720);
or U3916 (N_3916,N_3600,N_3521);
xor U3917 (N_3917,N_3677,N_3528);
or U3918 (N_3918,N_3518,N_3656);
and U3919 (N_3919,N_3630,N_3722);
or U3920 (N_3920,N_3663,N_3652);
or U3921 (N_3921,N_3598,N_3565);
nand U3922 (N_3922,N_3634,N_3556);
or U3923 (N_3923,N_3657,N_3537);
xor U3924 (N_3924,N_3625,N_3676);
nor U3925 (N_3925,N_3710,N_3718);
nor U3926 (N_3926,N_3717,N_3705);
and U3927 (N_3927,N_3669,N_3554);
xor U3928 (N_3928,N_3568,N_3507);
or U3929 (N_3929,N_3610,N_3557);
nand U3930 (N_3930,N_3610,N_3589);
xor U3931 (N_3931,N_3600,N_3573);
or U3932 (N_3932,N_3537,N_3571);
and U3933 (N_3933,N_3634,N_3570);
nor U3934 (N_3934,N_3581,N_3617);
nor U3935 (N_3935,N_3538,N_3510);
or U3936 (N_3936,N_3616,N_3596);
nor U3937 (N_3937,N_3679,N_3646);
nor U3938 (N_3938,N_3609,N_3619);
and U3939 (N_3939,N_3602,N_3723);
or U3940 (N_3940,N_3647,N_3597);
or U3941 (N_3941,N_3724,N_3690);
nand U3942 (N_3942,N_3635,N_3558);
nand U3943 (N_3943,N_3635,N_3723);
or U3944 (N_3944,N_3640,N_3523);
nand U3945 (N_3945,N_3618,N_3667);
xnor U3946 (N_3946,N_3668,N_3525);
nand U3947 (N_3947,N_3707,N_3520);
nand U3948 (N_3948,N_3619,N_3657);
or U3949 (N_3949,N_3619,N_3508);
nand U3950 (N_3950,N_3687,N_3568);
xnor U3951 (N_3951,N_3641,N_3583);
nor U3952 (N_3952,N_3525,N_3519);
or U3953 (N_3953,N_3597,N_3618);
nand U3954 (N_3954,N_3593,N_3739);
and U3955 (N_3955,N_3646,N_3537);
or U3956 (N_3956,N_3672,N_3740);
nand U3957 (N_3957,N_3672,N_3727);
nand U3958 (N_3958,N_3530,N_3561);
or U3959 (N_3959,N_3738,N_3687);
xnor U3960 (N_3960,N_3716,N_3622);
or U3961 (N_3961,N_3665,N_3704);
or U3962 (N_3962,N_3574,N_3544);
or U3963 (N_3963,N_3521,N_3565);
xor U3964 (N_3964,N_3505,N_3684);
nor U3965 (N_3965,N_3718,N_3555);
nand U3966 (N_3966,N_3508,N_3694);
nand U3967 (N_3967,N_3566,N_3708);
nand U3968 (N_3968,N_3633,N_3689);
and U3969 (N_3969,N_3575,N_3731);
xnor U3970 (N_3970,N_3547,N_3745);
and U3971 (N_3971,N_3577,N_3656);
nand U3972 (N_3972,N_3558,N_3711);
xnor U3973 (N_3973,N_3581,N_3513);
nor U3974 (N_3974,N_3601,N_3717);
nand U3975 (N_3975,N_3595,N_3594);
nand U3976 (N_3976,N_3522,N_3667);
and U3977 (N_3977,N_3601,N_3596);
nand U3978 (N_3978,N_3556,N_3640);
and U3979 (N_3979,N_3744,N_3527);
and U3980 (N_3980,N_3575,N_3532);
or U3981 (N_3981,N_3651,N_3518);
nand U3982 (N_3982,N_3581,N_3536);
nand U3983 (N_3983,N_3548,N_3684);
or U3984 (N_3984,N_3575,N_3683);
nor U3985 (N_3985,N_3574,N_3543);
or U3986 (N_3986,N_3626,N_3670);
nor U3987 (N_3987,N_3648,N_3512);
nor U3988 (N_3988,N_3629,N_3732);
nor U3989 (N_3989,N_3609,N_3737);
or U3990 (N_3990,N_3663,N_3702);
and U3991 (N_3991,N_3514,N_3553);
nand U3992 (N_3992,N_3527,N_3502);
and U3993 (N_3993,N_3551,N_3588);
or U3994 (N_3994,N_3715,N_3559);
nand U3995 (N_3995,N_3719,N_3577);
and U3996 (N_3996,N_3618,N_3590);
xnor U3997 (N_3997,N_3558,N_3503);
nand U3998 (N_3998,N_3699,N_3601);
or U3999 (N_3999,N_3738,N_3593);
or U4000 (N_4000,N_3938,N_3921);
nor U4001 (N_4001,N_3988,N_3818);
nand U4002 (N_4002,N_3815,N_3924);
or U4003 (N_4003,N_3892,N_3998);
nand U4004 (N_4004,N_3826,N_3769);
nor U4005 (N_4005,N_3939,N_3775);
xor U4006 (N_4006,N_3880,N_3985);
or U4007 (N_4007,N_3822,N_3945);
and U4008 (N_4008,N_3819,N_3872);
xor U4009 (N_4009,N_3852,N_3786);
and U4010 (N_4010,N_3866,N_3838);
nor U4011 (N_4011,N_3936,N_3759);
xnor U4012 (N_4012,N_3929,N_3993);
nor U4013 (N_4013,N_3952,N_3991);
nand U4014 (N_4014,N_3834,N_3969);
xnor U4015 (N_4015,N_3802,N_3837);
xnor U4016 (N_4016,N_3867,N_3783);
nand U4017 (N_4017,N_3789,N_3946);
nand U4018 (N_4018,N_3996,N_3785);
nor U4019 (N_4019,N_3904,N_3974);
and U4020 (N_4020,N_3806,N_3784);
or U4021 (N_4021,N_3887,N_3888);
nand U4022 (N_4022,N_3782,N_3849);
xnor U4023 (N_4023,N_3925,N_3916);
or U4024 (N_4024,N_3937,N_3980);
nor U4025 (N_4025,N_3790,N_3752);
and U4026 (N_4026,N_3861,N_3879);
and U4027 (N_4027,N_3987,N_3828);
xnor U4028 (N_4028,N_3931,N_3793);
nor U4029 (N_4029,N_3915,N_3941);
nand U4030 (N_4030,N_3981,N_3885);
nor U4031 (N_4031,N_3859,N_3779);
and U4032 (N_4032,N_3889,N_3798);
nor U4033 (N_4033,N_3792,N_3964);
or U4034 (N_4034,N_3754,N_3796);
nand U4035 (N_4035,N_3997,N_3940);
xnor U4036 (N_4036,N_3927,N_3965);
and U4037 (N_4037,N_3928,N_3949);
and U4038 (N_4038,N_3830,N_3777);
and U4039 (N_4039,N_3829,N_3912);
or U4040 (N_4040,N_3771,N_3765);
and U4041 (N_4041,N_3918,N_3820);
nor U4042 (N_4042,N_3760,N_3907);
or U4043 (N_4043,N_3773,N_3770);
and U4044 (N_4044,N_3891,N_3906);
nand U4045 (N_4045,N_3886,N_3840);
xnor U4046 (N_4046,N_3972,N_3768);
and U4047 (N_4047,N_3901,N_3932);
xor U4048 (N_4048,N_3862,N_3767);
nand U4049 (N_4049,N_3951,N_3905);
or U4050 (N_4050,N_3816,N_3989);
or U4051 (N_4051,N_3761,N_3922);
and U4052 (N_4052,N_3902,N_3944);
xor U4053 (N_4053,N_3978,N_3763);
and U4054 (N_4054,N_3864,N_3957);
xor U4055 (N_4055,N_3883,N_3908);
and U4056 (N_4056,N_3968,N_3855);
xnor U4057 (N_4057,N_3999,N_3757);
and U4058 (N_4058,N_3825,N_3774);
xor U4059 (N_4059,N_3933,N_3800);
xor U4060 (N_4060,N_3841,N_3971);
nor U4061 (N_4061,N_3961,N_3958);
or U4062 (N_4062,N_3909,N_3853);
and U4063 (N_4063,N_3871,N_3984);
nor U4064 (N_4064,N_3856,N_3995);
nor U4065 (N_4065,N_3935,N_3835);
nand U4066 (N_4066,N_3801,N_3821);
xnor U4067 (N_4067,N_3882,N_3874);
nor U4068 (N_4068,N_3923,N_3954);
xnor U4069 (N_4069,N_3890,N_3794);
nor U4070 (N_4070,N_3810,N_3776);
and U4071 (N_4071,N_3750,N_3863);
xnor U4072 (N_4072,N_3884,N_3960);
xor U4073 (N_4073,N_3911,N_3808);
nor U4074 (N_4074,N_3824,N_3832);
xnor U4075 (N_4075,N_3898,N_3780);
nor U4076 (N_4076,N_3850,N_3955);
and U4077 (N_4077,N_3860,N_3982);
xnor U4078 (N_4078,N_3803,N_3772);
xnor U4079 (N_4079,N_3868,N_3787);
xor U4080 (N_4080,N_3751,N_3873);
nand U4081 (N_4081,N_3817,N_3833);
nor U4082 (N_4082,N_3878,N_3854);
nor U4083 (N_4083,N_3919,N_3762);
nand U4084 (N_4084,N_3836,N_3865);
xnor U4085 (N_4085,N_3877,N_3809);
or U4086 (N_4086,N_3869,N_3788);
nand U4087 (N_4087,N_3917,N_3842);
or U4088 (N_4088,N_3897,N_3839);
nor U4089 (N_4089,N_3983,N_3813);
and U4090 (N_4090,N_3797,N_3962);
and U4091 (N_4091,N_3875,N_3956);
nor U4092 (N_4092,N_3844,N_3910);
xor U4093 (N_4093,N_3992,N_3950);
nand U4094 (N_4094,N_3758,N_3942);
nor U4095 (N_4095,N_3870,N_3948);
and U4096 (N_4096,N_3827,N_3976);
xnor U4097 (N_4097,N_3990,N_3900);
nor U4098 (N_4098,N_3795,N_3764);
nor U4099 (N_4099,N_3994,N_3913);
and U4100 (N_4100,N_3814,N_3807);
or U4101 (N_4101,N_3920,N_3799);
and U4102 (N_4102,N_3778,N_3753);
nand U4103 (N_4103,N_3903,N_3896);
nor U4104 (N_4104,N_3953,N_3847);
xnor U4105 (N_4105,N_3755,N_3926);
nor U4106 (N_4106,N_3805,N_3977);
or U4107 (N_4107,N_3848,N_3899);
or U4108 (N_4108,N_3966,N_3756);
and U4109 (N_4109,N_3858,N_3831);
nand U4110 (N_4110,N_3881,N_3973);
nor U4111 (N_4111,N_3843,N_3979);
and U4112 (N_4112,N_3970,N_3967);
and U4113 (N_4113,N_3947,N_3766);
and U4114 (N_4114,N_3930,N_3963);
and U4115 (N_4115,N_3876,N_3851);
nand U4116 (N_4116,N_3986,N_3914);
nand U4117 (N_4117,N_3812,N_3846);
xnor U4118 (N_4118,N_3893,N_3823);
nand U4119 (N_4119,N_3894,N_3895);
or U4120 (N_4120,N_3804,N_3975);
nor U4121 (N_4121,N_3791,N_3845);
or U4122 (N_4122,N_3781,N_3934);
nand U4123 (N_4123,N_3857,N_3943);
nand U4124 (N_4124,N_3811,N_3959);
nor U4125 (N_4125,N_3914,N_3936);
nor U4126 (N_4126,N_3919,N_3776);
nor U4127 (N_4127,N_3956,N_3975);
nor U4128 (N_4128,N_3879,N_3781);
nor U4129 (N_4129,N_3908,N_3993);
nand U4130 (N_4130,N_3879,N_3892);
or U4131 (N_4131,N_3928,N_3769);
or U4132 (N_4132,N_3990,N_3908);
nand U4133 (N_4133,N_3814,N_3998);
nand U4134 (N_4134,N_3802,N_3750);
or U4135 (N_4135,N_3834,N_3753);
nor U4136 (N_4136,N_3952,N_3769);
or U4137 (N_4137,N_3788,N_3882);
nand U4138 (N_4138,N_3995,N_3848);
nand U4139 (N_4139,N_3959,N_3867);
and U4140 (N_4140,N_3753,N_3922);
nand U4141 (N_4141,N_3872,N_3964);
nand U4142 (N_4142,N_3863,N_3841);
and U4143 (N_4143,N_3758,N_3930);
and U4144 (N_4144,N_3947,N_3820);
xnor U4145 (N_4145,N_3874,N_3978);
xor U4146 (N_4146,N_3999,N_3989);
and U4147 (N_4147,N_3869,N_3764);
and U4148 (N_4148,N_3762,N_3789);
xor U4149 (N_4149,N_3796,N_3862);
xor U4150 (N_4150,N_3913,N_3991);
nand U4151 (N_4151,N_3885,N_3965);
and U4152 (N_4152,N_3849,N_3880);
xnor U4153 (N_4153,N_3978,N_3977);
nor U4154 (N_4154,N_3963,N_3774);
nand U4155 (N_4155,N_3985,N_3890);
xor U4156 (N_4156,N_3765,N_3769);
nor U4157 (N_4157,N_3775,N_3869);
and U4158 (N_4158,N_3785,N_3934);
nor U4159 (N_4159,N_3753,N_3818);
xnor U4160 (N_4160,N_3771,N_3889);
and U4161 (N_4161,N_3860,N_3769);
xor U4162 (N_4162,N_3751,N_3830);
or U4163 (N_4163,N_3802,N_3770);
nor U4164 (N_4164,N_3933,N_3868);
xnor U4165 (N_4165,N_3769,N_3855);
and U4166 (N_4166,N_3841,N_3848);
xor U4167 (N_4167,N_3961,N_3911);
and U4168 (N_4168,N_3776,N_3964);
xor U4169 (N_4169,N_3897,N_3970);
or U4170 (N_4170,N_3784,N_3916);
and U4171 (N_4171,N_3751,N_3823);
or U4172 (N_4172,N_3897,N_3795);
nor U4173 (N_4173,N_3801,N_3950);
xnor U4174 (N_4174,N_3772,N_3759);
nor U4175 (N_4175,N_3811,N_3981);
and U4176 (N_4176,N_3938,N_3891);
nand U4177 (N_4177,N_3833,N_3992);
nor U4178 (N_4178,N_3948,N_3942);
and U4179 (N_4179,N_3899,N_3780);
xor U4180 (N_4180,N_3834,N_3750);
xnor U4181 (N_4181,N_3793,N_3962);
and U4182 (N_4182,N_3824,N_3904);
nand U4183 (N_4183,N_3937,N_3772);
nand U4184 (N_4184,N_3914,N_3956);
nor U4185 (N_4185,N_3887,N_3780);
or U4186 (N_4186,N_3992,N_3953);
or U4187 (N_4187,N_3912,N_3901);
or U4188 (N_4188,N_3766,N_3974);
nand U4189 (N_4189,N_3935,N_3822);
xnor U4190 (N_4190,N_3833,N_3784);
nand U4191 (N_4191,N_3941,N_3956);
and U4192 (N_4192,N_3799,N_3987);
nor U4193 (N_4193,N_3796,N_3960);
nor U4194 (N_4194,N_3851,N_3826);
nor U4195 (N_4195,N_3939,N_3851);
or U4196 (N_4196,N_3823,N_3861);
and U4197 (N_4197,N_3791,N_3934);
and U4198 (N_4198,N_3831,N_3963);
and U4199 (N_4199,N_3750,N_3839);
nor U4200 (N_4200,N_3911,N_3805);
nand U4201 (N_4201,N_3937,N_3840);
nor U4202 (N_4202,N_3913,N_3813);
xor U4203 (N_4203,N_3821,N_3879);
xor U4204 (N_4204,N_3784,N_3774);
nand U4205 (N_4205,N_3845,N_3860);
xor U4206 (N_4206,N_3833,N_3977);
or U4207 (N_4207,N_3806,N_3870);
xor U4208 (N_4208,N_3840,N_3790);
and U4209 (N_4209,N_3762,N_3864);
nor U4210 (N_4210,N_3835,N_3954);
or U4211 (N_4211,N_3830,N_3860);
nand U4212 (N_4212,N_3835,N_3758);
or U4213 (N_4213,N_3851,N_3906);
xnor U4214 (N_4214,N_3831,N_3952);
or U4215 (N_4215,N_3844,N_3981);
nor U4216 (N_4216,N_3896,N_3872);
and U4217 (N_4217,N_3844,N_3804);
nand U4218 (N_4218,N_3846,N_3915);
or U4219 (N_4219,N_3760,N_3820);
and U4220 (N_4220,N_3969,N_3948);
nand U4221 (N_4221,N_3936,N_3840);
xnor U4222 (N_4222,N_3879,N_3770);
nor U4223 (N_4223,N_3759,N_3895);
or U4224 (N_4224,N_3757,N_3907);
and U4225 (N_4225,N_3910,N_3846);
and U4226 (N_4226,N_3871,N_3750);
xor U4227 (N_4227,N_3927,N_3855);
nand U4228 (N_4228,N_3868,N_3817);
nand U4229 (N_4229,N_3793,N_3935);
xor U4230 (N_4230,N_3927,N_3785);
xnor U4231 (N_4231,N_3964,N_3974);
xor U4232 (N_4232,N_3814,N_3995);
nor U4233 (N_4233,N_3954,N_3929);
and U4234 (N_4234,N_3843,N_3799);
and U4235 (N_4235,N_3944,N_3966);
nand U4236 (N_4236,N_3851,N_3967);
nand U4237 (N_4237,N_3910,N_3829);
and U4238 (N_4238,N_3990,N_3901);
or U4239 (N_4239,N_3925,N_3841);
or U4240 (N_4240,N_3880,N_3752);
or U4241 (N_4241,N_3924,N_3778);
or U4242 (N_4242,N_3790,N_3998);
nand U4243 (N_4243,N_3992,N_3971);
nor U4244 (N_4244,N_3884,N_3946);
or U4245 (N_4245,N_3802,N_3889);
xnor U4246 (N_4246,N_3807,N_3768);
or U4247 (N_4247,N_3950,N_3957);
nor U4248 (N_4248,N_3864,N_3844);
nor U4249 (N_4249,N_3986,N_3810);
xnor U4250 (N_4250,N_4053,N_4036);
nor U4251 (N_4251,N_4106,N_4044);
nand U4252 (N_4252,N_4197,N_4172);
nor U4253 (N_4253,N_4232,N_4098);
xor U4254 (N_4254,N_4242,N_4164);
nand U4255 (N_4255,N_4108,N_4227);
xor U4256 (N_4256,N_4169,N_4024);
xor U4257 (N_4257,N_4084,N_4145);
xnor U4258 (N_4258,N_4120,N_4231);
xnor U4259 (N_4259,N_4074,N_4161);
and U4260 (N_4260,N_4209,N_4059);
nor U4261 (N_4261,N_4207,N_4092);
or U4262 (N_4262,N_4191,N_4135);
nor U4263 (N_4263,N_4114,N_4151);
and U4264 (N_4264,N_4090,N_4236);
and U4265 (N_4265,N_4241,N_4221);
xnor U4266 (N_4266,N_4125,N_4113);
or U4267 (N_4267,N_4055,N_4035);
nand U4268 (N_4268,N_4111,N_4046);
nand U4269 (N_4269,N_4173,N_4229);
and U4270 (N_4270,N_4131,N_4147);
and U4271 (N_4271,N_4187,N_4204);
and U4272 (N_4272,N_4089,N_4050);
nor U4273 (N_4273,N_4008,N_4006);
or U4274 (N_4274,N_4034,N_4222);
and U4275 (N_4275,N_4015,N_4142);
or U4276 (N_4276,N_4117,N_4109);
or U4277 (N_4277,N_4121,N_4011);
and U4278 (N_4278,N_4212,N_4080);
xor U4279 (N_4279,N_4192,N_4021);
and U4280 (N_4280,N_4193,N_4026);
and U4281 (N_4281,N_4058,N_4130);
and U4282 (N_4282,N_4025,N_4051);
and U4283 (N_4283,N_4143,N_4223);
nand U4284 (N_4284,N_4004,N_4082);
or U4285 (N_4285,N_4023,N_4219);
or U4286 (N_4286,N_4183,N_4218);
nand U4287 (N_4287,N_4107,N_4194);
nand U4288 (N_4288,N_4163,N_4073);
nor U4289 (N_4289,N_4030,N_4152);
nor U4290 (N_4290,N_4160,N_4102);
and U4291 (N_4291,N_4019,N_4245);
xor U4292 (N_4292,N_4122,N_4129);
nand U4293 (N_4293,N_4017,N_4198);
or U4294 (N_4294,N_4119,N_4140);
xor U4295 (N_4295,N_4065,N_4237);
nand U4296 (N_4296,N_4244,N_4216);
nor U4297 (N_4297,N_4190,N_4031);
nand U4298 (N_4298,N_4047,N_4134);
nor U4299 (N_4299,N_4064,N_4180);
and U4300 (N_4300,N_4206,N_4081);
or U4301 (N_4301,N_4101,N_4174);
nor U4302 (N_4302,N_4040,N_4176);
nor U4303 (N_4303,N_4038,N_4203);
and U4304 (N_4304,N_4137,N_4002);
or U4305 (N_4305,N_4014,N_4226);
nor U4306 (N_4306,N_4105,N_4138);
and U4307 (N_4307,N_4115,N_4096);
or U4308 (N_4308,N_4007,N_4132);
nor U4309 (N_4309,N_4022,N_4230);
nand U4310 (N_4310,N_4016,N_4133);
nand U4311 (N_4311,N_4093,N_4063);
and U4312 (N_4312,N_4072,N_4099);
and U4313 (N_4313,N_4153,N_4154);
or U4314 (N_4314,N_4067,N_4078);
nand U4315 (N_4315,N_4139,N_4233);
nand U4316 (N_4316,N_4196,N_4056);
nor U4317 (N_4317,N_4200,N_4116);
xor U4318 (N_4318,N_4086,N_4248);
or U4319 (N_4319,N_4186,N_4042);
nor U4320 (N_4320,N_4094,N_4039);
nor U4321 (N_4321,N_4238,N_4032);
nor U4322 (N_4322,N_4168,N_4175);
nand U4323 (N_4323,N_4027,N_4087);
xor U4324 (N_4324,N_4217,N_4155);
xor U4325 (N_4325,N_4118,N_4201);
nand U4326 (N_4326,N_4210,N_4061);
and U4327 (N_4327,N_4185,N_4178);
and U4328 (N_4328,N_4124,N_4184);
nor U4329 (N_4329,N_4123,N_4127);
and U4330 (N_4330,N_4028,N_4071);
or U4331 (N_4331,N_4104,N_4158);
nand U4332 (N_4332,N_4213,N_4097);
or U4333 (N_4333,N_4181,N_4202);
nor U4334 (N_4334,N_4225,N_4239);
and U4335 (N_4335,N_4013,N_4220);
nand U4336 (N_4336,N_4159,N_4179);
and U4337 (N_4337,N_4020,N_4005);
nand U4338 (N_4338,N_4240,N_4085);
nor U4339 (N_4339,N_4057,N_4167);
or U4340 (N_4340,N_4045,N_4243);
xor U4341 (N_4341,N_4009,N_4049);
nand U4342 (N_4342,N_4228,N_4037);
nor U4343 (N_4343,N_4001,N_4141);
xor U4344 (N_4344,N_4208,N_4211);
or U4345 (N_4345,N_4079,N_4062);
nor U4346 (N_4346,N_4171,N_4060);
nor U4347 (N_4347,N_4249,N_4043);
and U4348 (N_4348,N_4166,N_4162);
nor U4349 (N_4349,N_4144,N_4170);
nor U4350 (N_4350,N_4157,N_4136);
or U4351 (N_4351,N_4215,N_4100);
or U4352 (N_4352,N_4018,N_4126);
nand U4353 (N_4353,N_4205,N_4091);
xnor U4354 (N_4354,N_4246,N_4095);
nor U4355 (N_4355,N_4112,N_4128);
or U4356 (N_4356,N_4066,N_4199);
xnor U4357 (N_4357,N_4214,N_4165);
and U4358 (N_4358,N_4003,N_4182);
nor U4359 (N_4359,N_4033,N_4076);
xnor U4360 (N_4360,N_4012,N_4156);
xnor U4361 (N_4361,N_4068,N_4150);
nor U4362 (N_4362,N_4148,N_4010);
xnor U4363 (N_4363,N_4075,N_4146);
nand U4364 (N_4364,N_4195,N_4048);
xor U4365 (N_4365,N_4077,N_4070);
nor U4366 (N_4366,N_4069,N_4224);
or U4367 (N_4367,N_4149,N_4247);
nor U4368 (N_4368,N_4234,N_4052);
or U4369 (N_4369,N_4041,N_4000);
nor U4370 (N_4370,N_4054,N_4103);
xnor U4371 (N_4371,N_4088,N_4235);
xnor U4372 (N_4372,N_4083,N_4110);
nand U4373 (N_4373,N_4177,N_4029);
xor U4374 (N_4374,N_4189,N_4188);
or U4375 (N_4375,N_4180,N_4192);
and U4376 (N_4376,N_4238,N_4107);
or U4377 (N_4377,N_4223,N_4085);
nand U4378 (N_4378,N_4114,N_4112);
nand U4379 (N_4379,N_4072,N_4150);
or U4380 (N_4380,N_4044,N_4200);
xnor U4381 (N_4381,N_4185,N_4119);
xor U4382 (N_4382,N_4150,N_4077);
nand U4383 (N_4383,N_4142,N_4124);
and U4384 (N_4384,N_4032,N_4055);
xnor U4385 (N_4385,N_4188,N_4077);
nand U4386 (N_4386,N_4171,N_4244);
nor U4387 (N_4387,N_4007,N_4017);
or U4388 (N_4388,N_4057,N_4123);
and U4389 (N_4389,N_4242,N_4175);
or U4390 (N_4390,N_4141,N_4075);
nand U4391 (N_4391,N_4010,N_4020);
nor U4392 (N_4392,N_4207,N_4133);
xor U4393 (N_4393,N_4126,N_4013);
nor U4394 (N_4394,N_4091,N_4114);
or U4395 (N_4395,N_4120,N_4168);
xor U4396 (N_4396,N_4194,N_4009);
xnor U4397 (N_4397,N_4078,N_4011);
or U4398 (N_4398,N_4216,N_4033);
xor U4399 (N_4399,N_4086,N_4209);
xor U4400 (N_4400,N_4027,N_4075);
or U4401 (N_4401,N_4208,N_4063);
nor U4402 (N_4402,N_4046,N_4049);
xor U4403 (N_4403,N_4004,N_4191);
nor U4404 (N_4404,N_4160,N_4172);
and U4405 (N_4405,N_4193,N_4221);
nand U4406 (N_4406,N_4033,N_4010);
xnor U4407 (N_4407,N_4229,N_4120);
or U4408 (N_4408,N_4143,N_4210);
and U4409 (N_4409,N_4031,N_4154);
xnor U4410 (N_4410,N_4031,N_4011);
and U4411 (N_4411,N_4073,N_4016);
xor U4412 (N_4412,N_4122,N_4133);
and U4413 (N_4413,N_4135,N_4034);
nand U4414 (N_4414,N_4107,N_4097);
xnor U4415 (N_4415,N_4191,N_4249);
nand U4416 (N_4416,N_4161,N_4198);
nand U4417 (N_4417,N_4023,N_4188);
nor U4418 (N_4418,N_4199,N_4032);
or U4419 (N_4419,N_4076,N_4151);
xnor U4420 (N_4420,N_4041,N_4086);
nand U4421 (N_4421,N_4080,N_4166);
or U4422 (N_4422,N_4175,N_4185);
and U4423 (N_4423,N_4067,N_4002);
nand U4424 (N_4424,N_4178,N_4069);
xnor U4425 (N_4425,N_4087,N_4167);
nor U4426 (N_4426,N_4072,N_4128);
and U4427 (N_4427,N_4033,N_4128);
and U4428 (N_4428,N_4118,N_4223);
or U4429 (N_4429,N_4023,N_4181);
nor U4430 (N_4430,N_4011,N_4199);
nand U4431 (N_4431,N_4000,N_4057);
xor U4432 (N_4432,N_4108,N_4193);
and U4433 (N_4433,N_4142,N_4102);
and U4434 (N_4434,N_4111,N_4129);
nor U4435 (N_4435,N_4089,N_4122);
and U4436 (N_4436,N_4221,N_4106);
xor U4437 (N_4437,N_4101,N_4249);
or U4438 (N_4438,N_4131,N_4015);
nand U4439 (N_4439,N_4077,N_4050);
and U4440 (N_4440,N_4120,N_4122);
and U4441 (N_4441,N_4072,N_4027);
nand U4442 (N_4442,N_4237,N_4021);
nor U4443 (N_4443,N_4081,N_4048);
or U4444 (N_4444,N_4030,N_4170);
nand U4445 (N_4445,N_4082,N_4065);
xnor U4446 (N_4446,N_4115,N_4109);
and U4447 (N_4447,N_4165,N_4115);
xor U4448 (N_4448,N_4082,N_4023);
nor U4449 (N_4449,N_4198,N_4041);
nand U4450 (N_4450,N_4009,N_4176);
nand U4451 (N_4451,N_4096,N_4038);
nor U4452 (N_4452,N_4185,N_4215);
nand U4453 (N_4453,N_4035,N_4088);
nand U4454 (N_4454,N_4097,N_4059);
and U4455 (N_4455,N_4239,N_4248);
or U4456 (N_4456,N_4219,N_4058);
or U4457 (N_4457,N_4161,N_4156);
nor U4458 (N_4458,N_4034,N_4131);
nor U4459 (N_4459,N_4004,N_4114);
xor U4460 (N_4460,N_4016,N_4104);
nor U4461 (N_4461,N_4165,N_4125);
nor U4462 (N_4462,N_4012,N_4128);
or U4463 (N_4463,N_4020,N_4078);
or U4464 (N_4464,N_4001,N_4038);
and U4465 (N_4465,N_4241,N_4085);
xnor U4466 (N_4466,N_4162,N_4146);
or U4467 (N_4467,N_4139,N_4099);
and U4468 (N_4468,N_4040,N_4017);
xor U4469 (N_4469,N_4186,N_4128);
nand U4470 (N_4470,N_4030,N_4208);
or U4471 (N_4471,N_4010,N_4131);
or U4472 (N_4472,N_4187,N_4099);
and U4473 (N_4473,N_4062,N_4100);
or U4474 (N_4474,N_4103,N_4139);
nand U4475 (N_4475,N_4047,N_4159);
nor U4476 (N_4476,N_4036,N_4101);
and U4477 (N_4477,N_4030,N_4064);
xnor U4478 (N_4478,N_4233,N_4002);
or U4479 (N_4479,N_4083,N_4068);
xor U4480 (N_4480,N_4170,N_4091);
xor U4481 (N_4481,N_4082,N_4204);
nor U4482 (N_4482,N_4213,N_4212);
nor U4483 (N_4483,N_4164,N_4226);
nor U4484 (N_4484,N_4145,N_4049);
nor U4485 (N_4485,N_4183,N_4160);
nor U4486 (N_4486,N_4067,N_4136);
or U4487 (N_4487,N_4091,N_4070);
nor U4488 (N_4488,N_4232,N_4124);
nor U4489 (N_4489,N_4236,N_4087);
and U4490 (N_4490,N_4239,N_4058);
or U4491 (N_4491,N_4158,N_4235);
and U4492 (N_4492,N_4055,N_4105);
and U4493 (N_4493,N_4036,N_4059);
nor U4494 (N_4494,N_4012,N_4124);
or U4495 (N_4495,N_4153,N_4246);
or U4496 (N_4496,N_4002,N_4143);
and U4497 (N_4497,N_4057,N_4194);
nand U4498 (N_4498,N_4210,N_4128);
nand U4499 (N_4499,N_4152,N_4057);
nor U4500 (N_4500,N_4441,N_4314);
nor U4501 (N_4501,N_4376,N_4440);
and U4502 (N_4502,N_4436,N_4364);
xnor U4503 (N_4503,N_4311,N_4448);
or U4504 (N_4504,N_4462,N_4359);
nand U4505 (N_4505,N_4250,N_4413);
nor U4506 (N_4506,N_4377,N_4253);
nand U4507 (N_4507,N_4469,N_4295);
xnor U4508 (N_4508,N_4452,N_4433);
nor U4509 (N_4509,N_4287,N_4453);
xor U4510 (N_4510,N_4428,N_4327);
or U4511 (N_4511,N_4497,N_4350);
nor U4512 (N_4512,N_4389,N_4284);
nand U4513 (N_4513,N_4361,N_4269);
and U4514 (N_4514,N_4353,N_4483);
or U4515 (N_4515,N_4496,N_4379);
or U4516 (N_4516,N_4339,N_4352);
xnor U4517 (N_4517,N_4255,N_4263);
nand U4518 (N_4518,N_4267,N_4400);
or U4519 (N_4519,N_4490,N_4477);
nor U4520 (N_4520,N_4378,N_4320);
xnor U4521 (N_4521,N_4473,N_4435);
or U4522 (N_4522,N_4439,N_4485);
or U4523 (N_4523,N_4310,N_4375);
nor U4524 (N_4524,N_4398,N_4272);
or U4525 (N_4525,N_4261,N_4312);
xnor U4526 (N_4526,N_4289,N_4293);
and U4527 (N_4527,N_4368,N_4494);
or U4528 (N_4528,N_4424,N_4273);
and U4529 (N_4529,N_4489,N_4437);
xnor U4530 (N_4530,N_4406,N_4427);
nor U4531 (N_4531,N_4450,N_4369);
or U4532 (N_4532,N_4401,N_4347);
or U4533 (N_4533,N_4421,N_4288);
nor U4534 (N_4534,N_4384,N_4499);
xor U4535 (N_4535,N_4296,N_4317);
and U4536 (N_4536,N_4336,N_4266);
or U4537 (N_4537,N_4372,N_4467);
and U4538 (N_4538,N_4345,N_4493);
or U4539 (N_4539,N_4470,N_4324);
xnor U4540 (N_4540,N_4438,N_4454);
or U4541 (N_4541,N_4323,N_4290);
nor U4542 (N_4542,N_4260,N_4471);
and U4543 (N_4543,N_4309,N_4276);
and U4544 (N_4544,N_4355,N_4264);
or U4545 (N_4545,N_4262,N_4465);
or U4546 (N_4546,N_4299,N_4358);
xnor U4547 (N_4547,N_4300,N_4283);
or U4548 (N_4548,N_4399,N_4380);
or U4549 (N_4549,N_4430,N_4444);
or U4550 (N_4550,N_4418,N_4387);
and U4551 (N_4551,N_4419,N_4486);
nor U4552 (N_4552,N_4363,N_4275);
nand U4553 (N_4553,N_4495,N_4366);
and U4554 (N_4554,N_4409,N_4482);
nand U4555 (N_4555,N_4270,N_4447);
nor U4556 (N_4556,N_4412,N_4395);
nor U4557 (N_4557,N_4331,N_4292);
nand U4558 (N_4558,N_4472,N_4252);
nor U4559 (N_4559,N_4426,N_4442);
or U4560 (N_4560,N_4476,N_4307);
and U4561 (N_4561,N_4414,N_4280);
xnor U4562 (N_4562,N_4468,N_4356);
xor U4563 (N_4563,N_4456,N_4431);
or U4564 (N_4564,N_4291,N_4333);
nor U4565 (N_4565,N_4349,N_4302);
or U4566 (N_4566,N_4411,N_4481);
nand U4567 (N_4567,N_4268,N_4383);
and U4568 (N_4568,N_4475,N_4397);
and U4569 (N_4569,N_4479,N_4308);
xnor U4570 (N_4570,N_4271,N_4251);
nor U4571 (N_4571,N_4342,N_4434);
nor U4572 (N_4572,N_4304,N_4254);
and U4573 (N_4573,N_4371,N_4257);
xnor U4574 (N_4574,N_4385,N_4321);
nor U4575 (N_4575,N_4391,N_4474);
nand U4576 (N_4576,N_4373,N_4492);
nor U4577 (N_4577,N_4281,N_4341);
xnor U4578 (N_4578,N_4423,N_4484);
or U4579 (N_4579,N_4298,N_4390);
or U4580 (N_4580,N_4370,N_4374);
and U4581 (N_4581,N_4330,N_4420);
nor U4582 (N_4582,N_4403,N_4357);
and U4583 (N_4583,N_4392,N_4259);
and U4584 (N_4584,N_4408,N_4449);
nor U4585 (N_4585,N_4458,N_4265);
nor U4586 (N_4586,N_4491,N_4416);
nor U4587 (N_4587,N_4394,N_4360);
nand U4588 (N_4588,N_4343,N_4301);
or U4589 (N_4589,N_4460,N_4381);
xor U4590 (N_4590,N_4354,N_4297);
nand U4591 (N_4591,N_4348,N_4480);
nand U4592 (N_4592,N_4386,N_4282);
xor U4593 (N_4593,N_4279,N_4325);
xnor U4594 (N_4594,N_4388,N_4415);
or U4595 (N_4595,N_4274,N_4329);
and U4596 (N_4596,N_4322,N_4258);
nand U4597 (N_4597,N_4455,N_4382);
xnor U4598 (N_4598,N_4396,N_4443);
nor U4599 (N_4599,N_4319,N_4464);
or U4600 (N_4600,N_4393,N_4316);
nand U4601 (N_4601,N_4285,N_4429);
nor U4602 (N_4602,N_4305,N_4362);
nand U4603 (N_4603,N_4417,N_4466);
nand U4604 (N_4604,N_4326,N_4256);
or U4605 (N_4605,N_4286,N_4328);
nand U4606 (N_4606,N_4459,N_4410);
xnor U4607 (N_4607,N_4478,N_4313);
nand U4608 (N_4608,N_4365,N_4346);
xnor U4609 (N_4609,N_4451,N_4498);
xor U4610 (N_4610,N_4335,N_4334);
nor U4611 (N_4611,N_4404,N_4432);
and U4612 (N_4612,N_4306,N_4337);
and U4613 (N_4613,N_4344,N_4367);
and U4614 (N_4614,N_4422,N_4278);
nand U4615 (N_4615,N_4445,N_4457);
or U4616 (N_4616,N_4338,N_4461);
and U4617 (N_4617,N_4332,N_4487);
and U4618 (N_4618,N_4405,N_4294);
nor U4619 (N_4619,N_4402,N_4277);
and U4620 (N_4620,N_4488,N_4446);
xor U4621 (N_4621,N_4315,N_4463);
xnor U4622 (N_4622,N_4340,N_4407);
xnor U4623 (N_4623,N_4425,N_4303);
nor U4624 (N_4624,N_4318,N_4351);
xor U4625 (N_4625,N_4285,N_4396);
and U4626 (N_4626,N_4360,N_4441);
nor U4627 (N_4627,N_4490,N_4357);
or U4628 (N_4628,N_4454,N_4371);
nor U4629 (N_4629,N_4262,N_4466);
and U4630 (N_4630,N_4438,N_4462);
or U4631 (N_4631,N_4471,N_4292);
and U4632 (N_4632,N_4305,N_4426);
xnor U4633 (N_4633,N_4306,N_4445);
nor U4634 (N_4634,N_4278,N_4480);
nor U4635 (N_4635,N_4416,N_4271);
xnor U4636 (N_4636,N_4321,N_4294);
nand U4637 (N_4637,N_4354,N_4376);
or U4638 (N_4638,N_4362,N_4351);
nor U4639 (N_4639,N_4483,N_4455);
nand U4640 (N_4640,N_4479,N_4417);
nand U4641 (N_4641,N_4477,N_4396);
xor U4642 (N_4642,N_4332,N_4465);
nand U4643 (N_4643,N_4273,N_4447);
and U4644 (N_4644,N_4355,N_4301);
and U4645 (N_4645,N_4394,N_4496);
nand U4646 (N_4646,N_4401,N_4308);
nor U4647 (N_4647,N_4449,N_4471);
or U4648 (N_4648,N_4489,N_4370);
and U4649 (N_4649,N_4458,N_4414);
xor U4650 (N_4650,N_4261,N_4480);
xor U4651 (N_4651,N_4341,N_4357);
and U4652 (N_4652,N_4271,N_4496);
and U4653 (N_4653,N_4288,N_4256);
and U4654 (N_4654,N_4259,N_4264);
or U4655 (N_4655,N_4318,N_4313);
nor U4656 (N_4656,N_4405,N_4456);
nor U4657 (N_4657,N_4296,N_4294);
and U4658 (N_4658,N_4305,N_4364);
or U4659 (N_4659,N_4332,N_4350);
xnor U4660 (N_4660,N_4358,N_4301);
or U4661 (N_4661,N_4278,N_4334);
and U4662 (N_4662,N_4269,N_4327);
nand U4663 (N_4663,N_4466,N_4313);
and U4664 (N_4664,N_4276,N_4302);
nand U4665 (N_4665,N_4316,N_4492);
or U4666 (N_4666,N_4415,N_4424);
nand U4667 (N_4667,N_4290,N_4277);
or U4668 (N_4668,N_4369,N_4454);
xnor U4669 (N_4669,N_4416,N_4351);
xor U4670 (N_4670,N_4434,N_4441);
or U4671 (N_4671,N_4477,N_4466);
and U4672 (N_4672,N_4336,N_4472);
xnor U4673 (N_4673,N_4440,N_4384);
nand U4674 (N_4674,N_4379,N_4269);
nor U4675 (N_4675,N_4422,N_4317);
xnor U4676 (N_4676,N_4356,N_4257);
and U4677 (N_4677,N_4420,N_4362);
xnor U4678 (N_4678,N_4350,N_4498);
nor U4679 (N_4679,N_4324,N_4269);
xor U4680 (N_4680,N_4363,N_4274);
and U4681 (N_4681,N_4456,N_4286);
xor U4682 (N_4682,N_4469,N_4256);
and U4683 (N_4683,N_4390,N_4451);
nor U4684 (N_4684,N_4270,N_4431);
nand U4685 (N_4685,N_4307,N_4469);
nor U4686 (N_4686,N_4358,N_4332);
nand U4687 (N_4687,N_4412,N_4462);
xor U4688 (N_4688,N_4455,N_4413);
xnor U4689 (N_4689,N_4467,N_4263);
and U4690 (N_4690,N_4261,N_4496);
or U4691 (N_4691,N_4380,N_4486);
xnor U4692 (N_4692,N_4461,N_4497);
xnor U4693 (N_4693,N_4267,N_4452);
nand U4694 (N_4694,N_4463,N_4340);
and U4695 (N_4695,N_4448,N_4336);
nor U4696 (N_4696,N_4310,N_4414);
nand U4697 (N_4697,N_4278,N_4312);
xnor U4698 (N_4698,N_4413,N_4433);
xor U4699 (N_4699,N_4399,N_4488);
nor U4700 (N_4700,N_4274,N_4482);
or U4701 (N_4701,N_4271,N_4405);
nor U4702 (N_4702,N_4291,N_4271);
or U4703 (N_4703,N_4462,N_4379);
nor U4704 (N_4704,N_4414,N_4271);
and U4705 (N_4705,N_4453,N_4299);
nand U4706 (N_4706,N_4289,N_4492);
and U4707 (N_4707,N_4492,N_4460);
xnor U4708 (N_4708,N_4325,N_4481);
nand U4709 (N_4709,N_4463,N_4382);
and U4710 (N_4710,N_4291,N_4374);
or U4711 (N_4711,N_4320,N_4395);
xor U4712 (N_4712,N_4254,N_4335);
nand U4713 (N_4713,N_4326,N_4323);
xor U4714 (N_4714,N_4289,N_4305);
nor U4715 (N_4715,N_4289,N_4388);
nand U4716 (N_4716,N_4385,N_4399);
nand U4717 (N_4717,N_4370,N_4253);
or U4718 (N_4718,N_4472,N_4311);
or U4719 (N_4719,N_4309,N_4302);
nor U4720 (N_4720,N_4283,N_4423);
and U4721 (N_4721,N_4298,N_4393);
or U4722 (N_4722,N_4453,N_4446);
nand U4723 (N_4723,N_4250,N_4330);
xnor U4724 (N_4724,N_4459,N_4341);
nand U4725 (N_4725,N_4499,N_4325);
xor U4726 (N_4726,N_4270,N_4422);
or U4727 (N_4727,N_4496,N_4357);
or U4728 (N_4728,N_4406,N_4301);
nand U4729 (N_4729,N_4480,N_4366);
xor U4730 (N_4730,N_4265,N_4253);
nand U4731 (N_4731,N_4452,N_4268);
nand U4732 (N_4732,N_4280,N_4468);
xnor U4733 (N_4733,N_4461,N_4372);
nand U4734 (N_4734,N_4334,N_4484);
and U4735 (N_4735,N_4287,N_4352);
xnor U4736 (N_4736,N_4283,N_4390);
xnor U4737 (N_4737,N_4306,N_4382);
nor U4738 (N_4738,N_4258,N_4426);
nor U4739 (N_4739,N_4434,N_4377);
and U4740 (N_4740,N_4321,N_4461);
or U4741 (N_4741,N_4325,N_4253);
xor U4742 (N_4742,N_4468,N_4359);
nand U4743 (N_4743,N_4269,N_4335);
nor U4744 (N_4744,N_4464,N_4337);
nor U4745 (N_4745,N_4398,N_4277);
nor U4746 (N_4746,N_4434,N_4492);
and U4747 (N_4747,N_4333,N_4373);
nor U4748 (N_4748,N_4318,N_4407);
and U4749 (N_4749,N_4394,N_4303);
nor U4750 (N_4750,N_4570,N_4748);
nor U4751 (N_4751,N_4680,N_4609);
or U4752 (N_4752,N_4623,N_4504);
or U4753 (N_4753,N_4659,N_4643);
or U4754 (N_4754,N_4638,N_4719);
xor U4755 (N_4755,N_4654,N_4528);
xnor U4756 (N_4756,N_4551,N_4517);
and U4757 (N_4757,N_4622,N_4565);
nand U4758 (N_4758,N_4685,N_4503);
xnor U4759 (N_4759,N_4629,N_4745);
nor U4760 (N_4760,N_4652,N_4675);
xnor U4761 (N_4761,N_4729,N_4558);
nand U4762 (N_4762,N_4522,N_4548);
nand U4763 (N_4763,N_4670,N_4605);
or U4764 (N_4764,N_4684,N_4710);
xnor U4765 (N_4765,N_4718,N_4656);
and U4766 (N_4766,N_4508,N_4529);
nor U4767 (N_4767,N_4704,N_4667);
xor U4768 (N_4768,N_4627,N_4635);
nor U4769 (N_4769,N_4688,N_4614);
nand U4770 (N_4770,N_4516,N_4573);
or U4771 (N_4771,N_4723,N_4537);
or U4772 (N_4772,N_4692,N_4519);
or U4773 (N_4773,N_4730,N_4501);
xnor U4774 (N_4774,N_4637,N_4713);
or U4775 (N_4775,N_4582,N_4703);
or U4776 (N_4776,N_4624,N_4673);
and U4777 (N_4777,N_4598,N_4708);
and U4778 (N_4778,N_4649,N_4615);
or U4779 (N_4779,N_4502,N_4647);
or U4780 (N_4780,N_4572,N_4523);
or U4781 (N_4781,N_4617,N_4698);
nand U4782 (N_4782,N_4541,N_4722);
nand U4783 (N_4783,N_4648,N_4734);
and U4784 (N_4784,N_4592,N_4535);
nor U4785 (N_4785,N_4613,N_4591);
nand U4786 (N_4786,N_4521,N_4612);
xor U4787 (N_4787,N_4737,N_4744);
or U4788 (N_4788,N_4539,N_4579);
or U4789 (N_4789,N_4662,N_4630);
and U4790 (N_4790,N_4634,N_4714);
and U4791 (N_4791,N_4686,N_4527);
or U4792 (N_4792,N_4542,N_4590);
and U4793 (N_4793,N_4661,N_4653);
or U4794 (N_4794,N_4561,N_4511);
and U4795 (N_4795,N_4538,N_4640);
and U4796 (N_4796,N_4666,N_4721);
xor U4797 (N_4797,N_4696,N_4520);
and U4798 (N_4798,N_4544,N_4694);
nor U4799 (N_4799,N_4687,N_4738);
or U4800 (N_4800,N_4583,N_4672);
nor U4801 (N_4801,N_4602,N_4608);
or U4802 (N_4802,N_4510,N_4611);
nand U4803 (N_4803,N_4540,N_4628);
nor U4804 (N_4804,N_4682,N_4702);
xor U4805 (N_4805,N_4607,N_4564);
xor U4806 (N_4806,N_4536,N_4644);
nand U4807 (N_4807,N_4724,N_4717);
nand U4808 (N_4808,N_4651,N_4525);
and U4809 (N_4809,N_4679,N_4709);
nand U4810 (N_4810,N_4557,N_4707);
nand U4811 (N_4811,N_4690,N_4509);
xnor U4812 (N_4812,N_4728,N_4683);
nor U4813 (N_4813,N_4545,N_4568);
xor U4814 (N_4814,N_4747,N_4681);
nor U4815 (N_4815,N_4618,N_4736);
xnor U4816 (N_4816,N_4720,N_4712);
nor U4817 (N_4817,N_4619,N_4515);
nor U4818 (N_4818,N_4631,N_4514);
xor U4819 (N_4819,N_4588,N_4610);
or U4820 (N_4820,N_4584,N_4726);
or U4821 (N_4821,N_4505,N_4559);
nor U4822 (N_4822,N_4576,N_4567);
xnor U4823 (N_4823,N_4616,N_4566);
nand U4824 (N_4824,N_4674,N_4595);
or U4825 (N_4825,N_4549,N_4636);
nand U4826 (N_4826,N_4639,N_4524);
nor U4827 (N_4827,N_4735,N_4668);
nand U4828 (N_4828,N_4660,N_4620);
and U4829 (N_4829,N_4589,N_4664);
nor U4830 (N_4830,N_4533,N_4531);
nor U4831 (N_4831,N_4518,N_4700);
and U4832 (N_4832,N_4739,N_4731);
xor U4833 (N_4833,N_4601,N_4733);
xnor U4834 (N_4834,N_4597,N_4701);
nand U4835 (N_4835,N_4574,N_4526);
or U4836 (N_4836,N_4578,N_4553);
xor U4837 (N_4837,N_4532,N_4550);
xor U4838 (N_4838,N_4650,N_4727);
nor U4839 (N_4839,N_4633,N_4569);
xor U4840 (N_4840,N_4586,N_4507);
nand U4841 (N_4841,N_4740,N_4506);
nor U4842 (N_4842,N_4706,N_4658);
and U4843 (N_4843,N_4715,N_4530);
or U4844 (N_4844,N_4562,N_4543);
or U4845 (N_4845,N_4749,N_4534);
and U4846 (N_4846,N_4594,N_4716);
xor U4847 (N_4847,N_4547,N_4604);
nand U4848 (N_4848,N_4599,N_4575);
or U4849 (N_4849,N_4626,N_4646);
nand U4850 (N_4850,N_4596,N_4711);
nand U4851 (N_4851,N_4600,N_4693);
xnor U4852 (N_4852,N_4705,N_4645);
nor U4853 (N_4853,N_4741,N_4677);
or U4854 (N_4854,N_4512,N_4742);
nor U4855 (N_4855,N_4746,N_4743);
and U4856 (N_4856,N_4689,N_4669);
and U4857 (N_4857,N_4671,N_4606);
and U4858 (N_4858,N_4732,N_4581);
nor U4859 (N_4859,N_4641,N_4546);
nand U4860 (N_4860,N_4655,N_4571);
and U4861 (N_4861,N_4603,N_4663);
and U4862 (N_4862,N_4621,N_4657);
and U4863 (N_4863,N_4555,N_4554);
nand U4864 (N_4864,N_4552,N_4560);
nor U4865 (N_4865,N_4676,N_4625);
and U4866 (N_4866,N_4678,N_4563);
xnor U4867 (N_4867,N_4513,N_4593);
nor U4868 (N_4868,N_4665,N_4556);
or U4869 (N_4869,N_4500,N_4699);
or U4870 (N_4870,N_4697,N_4695);
xor U4871 (N_4871,N_4642,N_4632);
nor U4872 (N_4872,N_4580,N_4585);
nor U4873 (N_4873,N_4691,N_4725);
and U4874 (N_4874,N_4587,N_4577);
or U4875 (N_4875,N_4630,N_4627);
or U4876 (N_4876,N_4674,N_4701);
or U4877 (N_4877,N_4730,N_4524);
or U4878 (N_4878,N_4509,N_4607);
nand U4879 (N_4879,N_4645,N_4729);
and U4880 (N_4880,N_4614,N_4545);
xnor U4881 (N_4881,N_4723,N_4584);
and U4882 (N_4882,N_4544,N_4542);
nand U4883 (N_4883,N_4577,N_4627);
xnor U4884 (N_4884,N_4604,N_4636);
nor U4885 (N_4885,N_4505,N_4648);
and U4886 (N_4886,N_4592,N_4695);
nand U4887 (N_4887,N_4520,N_4730);
nand U4888 (N_4888,N_4532,N_4596);
nand U4889 (N_4889,N_4609,N_4518);
nor U4890 (N_4890,N_4666,N_4537);
nand U4891 (N_4891,N_4698,N_4545);
nand U4892 (N_4892,N_4539,N_4707);
nand U4893 (N_4893,N_4666,N_4500);
and U4894 (N_4894,N_4658,N_4728);
and U4895 (N_4895,N_4558,N_4738);
nor U4896 (N_4896,N_4657,N_4710);
nand U4897 (N_4897,N_4743,N_4729);
nand U4898 (N_4898,N_4673,N_4507);
or U4899 (N_4899,N_4625,N_4666);
nor U4900 (N_4900,N_4559,N_4730);
or U4901 (N_4901,N_4669,N_4591);
xor U4902 (N_4902,N_4579,N_4553);
nor U4903 (N_4903,N_4542,N_4713);
and U4904 (N_4904,N_4709,N_4627);
xor U4905 (N_4905,N_4500,N_4615);
nor U4906 (N_4906,N_4589,N_4660);
or U4907 (N_4907,N_4588,N_4653);
xnor U4908 (N_4908,N_4525,N_4678);
or U4909 (N_4909,N_4674,N_4525);
or U4910 (N_4910,N_4663,N_4512);
or U4911 (N_4911,N_4541,N_4584);
xor U4912 (N_4912,N_4652,N_4534);
xor U4913 (N_4913,N_4573,N_4734);
nand U4914 (N_4914,N_4663,N_4671);
nand U4915 (N_4915,N_4746,N_4557);
xnor U4916 (N_4916,N_4739,N_4570);
or U4917 (N_4917,N_4538,N_4572);
and U4918 (N_4918,N_4646,N_4716);
or U4919 (N_4919,N_4731,N_4658);
or U4920 (N_4920,N_4651,N_4741);
xor U4921 (N_4921,N_4635,N_4651);
or U4922 (N_4922,N_4547,N_4741);
nand U4923 (N_4923,N_4691,N_4666);
nor U4924 (N_4924,N_4725,N_4635);
or U4925 (N_4925,N_4655,N_4698);
or U4926 (N_4926,N_4614,N_4608);
xnor U4927 (N_4927,N_4543,N_4622);
and U4928 (N_4928,N_4609,N_4521);
and U4929 (N_4929,N_4664,N_4554);
or U4930 (N_4930,N_4559,N_4703);
nor U4931 (N_4931,N_4600,N_4664);
and U4932 (N_4932,N_4638,N_4725);
xnor U4933 (N_4933,N_4546,N_4746);
nand U4934 (N_4934,N_4595,N_4649);
and U4935 (N_4935,N_4565,N_4657);
nor U4936 (N_4936,N_4548,N_4693);
or U4937 (N_4937,N_4671,N_4613);
or U4938 (N_4938,N_4607,N_4687);
nor U4939 (N_4939,N_4607,N_4694);
xor U4940 (N_4940,N_4518,N_4598);
and U4941 (N_4941,N_4650,N_4555);
or U4942 (N_4942,N_4688,N_4711);
and U4943 (N_4943,N_4712,N_4629);
xnor U4944 (N_4944,N_4740,N_4722);
or U4945 (N_4945,N_4531,N_4616);
nand U4946 (N_4946,N_4678,N_4688);
xnor U4947 (N_4947,N_4556,N_4599);
nor U4948 (N_4948,N_4733,N_4627);
xor U4949 (N_4949,N_4532,N_4681);
nor U4950 (N_4950,N_4506,N_4617);
nand U4951 (N_4951,N_4723,N_4687);
or U4952 (N_4952,N_4513,N_4743);
nand U4953 (N_4953,N_4501,N_4513);
and U4954 (N_4954,N_4672,N_4642);
nand U4955 (N_4955,N_4625,N_4506);
or U4956 (N_4956,N_4551,N_4570);
and U4957 (N_4957,N_4568,N_4539);
nand U4958 (N_4958,N_4684,N_4619);
or U4959 (N_4959,N_4549,N_4577);
xor U4960 (N_4960,N_4654,N_4587);
and U4961 (N_4961,N_4525,N_4526);
and U4962 (N_4962,N_4645,N_4603);
nand U4963 (N_4963,N_4588,N_4737);
nand U4964 (N_4964,N_4674,N_4627);
xor U4965 (N_4965,N_4638,N_4571);
nand U4966 (N_4966,N_4518,N_4528);
nand U4967 (N_4967,N_4727,N_4522);
nand U4968 (N_4968,N_4514,N_4533);
nor U4969 (N_4969,N_4698,N_4694);
or U4970 (N_4970,N_4676,N_4532);
xnor U4971 (N_4971,N_4584,N_4571);
nand U4972 (N_4972,N_4601,N_4734);
nor U4973 (N_4973,N_4641,N_4675);
or U4974 (N_4974,N_4686,N_4500);
nand U4975 (N_4975,N_4734,N_4506);
nor U4976 (N_4976,N_4666,N_4563);
and U4977 (N_4977,N_4542,N_4553);
xnor U4978 (N_4978,N_4717,N_4676);
and U4979 (N_4979,N_4544,N_4511);
nor U4980 (N_4980,N_4536,N_4689);
nand U4981 (N_4981,N_4650,N_4527);
and U4982 (N_4982,N_4618,N_4514);
nor U4983 (N_4983,N_4709,N_4729);
xor U4984 (N_4984,N_4733,N_4680);
nor U4985 (N_4985,N_4611,N_4596);
nand U4986 (N_4986,N_4522,N_4648);
and U4987 (N_4987,N_4621,N_4526);
nor U4988 (N_4988,N_4732,N_4634);
and U4989 (N_4989,N_4747,N_4597);
nand U4990 (N_4990,N_4725,N_4643);
and U4991 (N_4991,N_4706,N_4607);
nor U4992 (N_4992,N_4566,N_4645);
nand U4993 (N_4993,N_4642,N_4725);
nand U4994 (N_4994,N_4513,N_4599);
or U4995 (N_4995,N_4684,N_4587);
nor U4996 (N_4996,N_4710,N_4531);
nor U4997 (N_4997,N_4510,N_4581);
and U4998 (N_4998,N_4524,N_4679);
and U4999 (N_4999,N_4633,N_4500);
xor U5000 (N_5000,N_4937,N_4957);
xor U5001 (N_5001,N_4921,N_4782);
and U5002 (N_5002,N_4852,N_4929);
or U5003 (N_5003,N_4996,N_4877);
and U5004 (N_5004,N_4901,N_4864);
xor U5005 (N_5005,N_4862,N_4753);
and U5006 (N_5006,N_4941,N_4761);
xor U5007 (N_5007,N_4773,N_4850);
or U5008 (N_5008,N_4875,N_4785);
or U5009 (N_5009,N_4824,N_4907);
nand U5010 (N_5010,N_4943,N_4906);
nor U5011 (N_5011,N_4873,N_4940);
xnor U5012 (N_5012,N_4965,N_4895);
nand U5013 (N_5013,N_4944,N_4926);
xnor U5014 (N_5014,N_4964,N_4777);
xnor U5015 (N_5015,N_4841,N_4843);
nor U5016 (N_5016,N_4898,N_4893);
nor U5017 (N_5017,N_4867,N_4967);
or U5018 (N_5018,N_4978,N_4903);
or U5019 (N_5019,N_4869,N_4987);
nor U5020 (N_5020,N_4958,N_4879);
nand U5021 (N_5021,N_4771,N_4812);
or U5022 (N_5022,N_4952,N_4985);
nand U5023 (N_5023,N_4870,N_4857);
xnor U5024 (N_5024,N_4800,N_4991);
xnor U5025 (N_5025,N_4999,N_4979);
xnor U5026 (N_5026,N_4768,N_4874);
nor U5027 (N_5027,N_4751,N_4989);
nand U5028 (N_5028,N_4792,N_4805);
nor U5029 (N_5029,N_4886,N_4894);
xor U5030 (N_5030,N_4835,N_4838);
and U5031 (N_5031,N_4885,N_4814);
nor U5032 (N_5032,N_4819,N_4826);
or U5033 (N_5033,N_4930,N_4960);
or U5034 (N_5034,N_4863,N_4971);
and U5035 (N_5035,N_4808,N_4902);
nor U5036 (N_5036,N_4828,N_4849);
or U5037 (N_5037,N_4832,N_4917);
nor U5038 (N_5038,N_4914,N_4823);
or U5039 (N_5039,N_4966,N_4983);
xor U5040 (N_5040,N_4918,N_4837);
xor U5041 (N_5041,N_4781,N_4866);
xor U5042 (N_5042,N_4922,N_4846);
nand U5043 (N_5043,N_4775,N_4779);
or U5044 (N_5044,N_4975,N_4897);
or U5045 (N_5045,N_4816,N_4924);
or U5046 (N_5046,N_4908,N_4767);
and U5047 (N_5047,N_4853,N_4970);
nand U5048 (N_5048,N_4935,N_4892);
and U5049 (N_5049,N_4912,N_4807);
nor U5050 (N_5050,N_4859,N_4790);
nand U5051 (N_5051,N_4946,N_4931);
and U5052 (N_5052,N_4860,N_4797);
and U5053 (N_5053,N_4923,N_4774);
nand U5054 (N_5054,N_4968,N_4963);
or U5055 (N_5055,N_4995,N_4789);
nor U5056 (N_5056,N_4772,N_4802);
xor U5057 (N_5057,N_4762,N_4791);
or U5058 (N_5058,N_4810,N_4955);
and U5059 (N_5059,N_4990,N_4798);
nand U5060 (N_5060,N_4969,N_4988);
nand U5061 (N_5061,N_4899,N_4954);
or U5062 (N_5062,N_4851,N_4848);
xor U5063 (N_5063,N_4769,N_4801);
or U5064 (N_5064,N_4856,N_4915);
xor U5065 (N_5065,N_4951,N_4932);
or U5066 (N_5066,N_4878,N_4758);
and U5067 (N_5067,N_4759,N_4977);
xor U5068 (N_5068,N_4760,N_4845);
and U5069 (N_5069,N_4766,N_4981);
xnor U5070 (N_5070,N_4793,N_4905);
and U5071 (N_5071,N_4834,N_4858);
nor U5072 (N_5072,N_4750,N_4854);
nor U5073 (N_5073,N_4765,N_4953);
nor U5074 (N_5074,N_4982,N_4821);
or U5075 (N_5075,N_4804,N_4962);
and U5076 (N_5076,N_4919,N_4884);
or U5077 (N_5077,N_4936,N_4881);
nor U5078 (N_5078,N_4786,N_4910);
nand U5079 (N_5079,N_4795,N_4882);
or U5080 (N_5080,N_4840,N_4974);
nor U5081 (N_5081,N_4756,N_4815);
or U5082 (N_5082,N_4872,N_4799);
nand U5083 (N_5083,N_4865,N_4980);
or U5084 (N_5084,N_4757,N_4788);
or U5085 (N_5085,N_4992,N_4984);
nand U5086 (N_5086,N_4998,N_4778);
nor U5087 (N_5087,N_4945,N_4820);
xor U5088 (N_5088,N_4787,N_4920);
or U5089 (N_5089,N_4887,N_4770);
nand U5090 (N_5090,N_4831,N_4783);
or U5091 (N_5091,N_4818,N_4780);
nor U5092 (N_5092,N_4889,N_4947);
xor U5093 (N_5093,N_4871,N_4861);
nand U5094 (N_5094,N_4833,N_4827);
nand U5095 (N_5095,N_4809,N_4976);
or U5096 (N_5096,N_4855,N_4900);
nor U5097 (N_5097,N_4803,N_4916);
nand U5098 (N_5098,N_4993,N_4948);
or U5099 (N_5099,N_4847,N_4997);
xor U5100 (N_5100,N_4752,N_4825);
and U5101 (N_5101,N_4763,N_4776);
xor U5102 (N_5102,N_4868,N_4961);
xor U5103 (N_5103,N_4959,N_4813);
xor U5104 (N_5104,N_4891,N_4754);
xor U5105 (N_5105,N_4927,N_4876);
or U5106 (N_5106,N_4956,N_4806);
nor U5107 (N_5107,N_4896,N_4794);
nor U5108 (N_5108,N_4764,N_4839);
or U5109 (N_5109,N_4934,N_4817);
and U5110 (N_5110,N_4994,N_4830);
nor U5111 (N_5111,N_4890,N_4938);
and U5112 (N_5112,N_4755,N_4949);
nor U5113 (N_5113,N_4842,N_4911);
xnor U5114 (N_5114,N_4972,N_4909);
nor U5115 (N_5115,N_4939,N_4904);
xnor U5116 (N_5116,N_4973,N_4784);
or U5117 (N_5117,N_4836,N_4986);
nor U5118 (N_5118,N_4933,N_4883);
nand U5119 (N_5119,N_4811,N_4913);
nand U5120 (N_5120,N_4880,N_4822);
and U5121 (N_5121,N_4829,N_4925);
nand U5122 (N_5122,N_4928,N_4888);
and U5123 (N_5123,N_4950,N_4942);
nand U5124 (N_5124,N_4844,N_4796);
xor U5125 (N_5125,N_4784,N_4830);
or U5126 (N_5126,N_4983,N_4957);
or U5127 (N_5127,N_4972,N_4979);
and U5128 (N_5128,N_4803,N_4982);
and U5129 (N_5129,N_4920,N_4781);
nand U5130 (N_5130,N_4980,N_4872);
nand U5131 (N_5131,N_4825,N_4942);
nor U5132 (N_5132,N_4898,N_4926);
nor U5133 (N_5133,N_4847,N_4870);
or U5134 (N_5134,N_4950,N_4828);
or U5135 (N_5135,N_4891,N_4843);
xor U5136 (N_5136,N_4849,N_4843);
or U5137 (N_5137,N_4918,N_4805);
and U5138 (N_5138,N_4916,N_4815);
or U5139 (N_5139,N_4793,N_4940);
xor U5140 (N_5140,N_4988,N_4914);
and U5141 (N_5141,N_4975,N_4806);
or U5142 (N_5142,N_4773,N_4762);
or U5143 (N_5143,N_4989,N_4968);
nor U5144 (N_5144,N_4915,N_4818);
and U5145 (N_5145,N_4928,N_4807);
nor U5146 (N_5146,N_4995,N_4997);
and U5147 (N_5147,N_4919,N_4760);
xor U5148 (N_5148,N_4911,N_4848);
or U5149 (N_5149,N_4883,N_4814);
nor U5150 (N_5150,N_4809,N_4855);
or U5151 (N_5151,N_4982,N_4871);
nand U5152 (N_5152,N_4817,N_4854);
xor U5153 (N_5153,N_4953,N_4757);
or U5154 (N_5154,N_4836,N_4788);
or U5155 (N_5155,N_4958,N_4951);
xnor U5156 (N_5156,N_4856,N_4823);
nor U5157 (N_5157,N_4864,N_4829);
and U5158 (N_5158,N_4952,N_4821);
or U5159 (N_5159,N_4921,N_4917);
or U5160 (N_5160,N_4934,N_4919);
xor U5161 (N_5161,N_4998,N_4894);
and U5162 (N_5162,N_4812,N_4968);
or U5163 (N_5163,N_4847,N_4890);
and U5164 (N_5164,N_4843,N_4831);
or U5165 (N_5165,N_4895,N_4789);
nand U5166 (N_5166,N_4947,N_4822);
nor U5167 (N_5167,N_4962,N_4909);
nor U5168 (N_5168,N_4836,N_4881);
xor U5169 (N_5169,N_4832,N_4964);
or U5170 (N_5170,N_4845,N_4831);
nand U5171 (N_5171,N_4980,N_4944);
xnor U5172 (N_5172,N_4869,N_4948);
nand U5173 (N_5173,N_4846,N_4794);
or U5174 (N_5174,N_4812,N_4935);
or U5175 (N_5175,N_4852,N_4812);
nand U5176 (N_5176,N_4792,N_4975);
nor U5177 (N_5177,N_4807,N_4892);
nor U5178 (N_5178,N_4960,N_4779);
xnor U5179 (N_5179,N_4927,N_4804);
xor U5180 (N_5180,N_4889,N_4828);
and U5181 (N_5181,N_4764,N_4994);
or U5182 (N_5182,N_4809,N_4972);
nand U5183 (N_5183,N_4756,N_4941);
and U5184 (N_5184,N_4955,N_4820);
nor U5185 (N_5185,N_4855,N_4974);
xor U5186 (N_5186,N_4939,N_4949);
nor U5187 (N_5187,N_4758,N_4831);
nor U5188 (N_5188,N_4900,N_4819);
or U5189 (N_5189,N_4914,N_4880);
or U5190 (N_5190,N_4757,N_4992);
nand U5191 (N_5191,N_4888,N_4773);
or U5192 (N_5192,N_4819,N_4803);
nor U5193 (N_5193,N_4950,N_4785);
nand U5194 (N_5194,N_4985,N_4928);
nor U5195 (N_5195,N_4867,N_4962);
nor U5196 (N_5196,N_4835,N_4982);
nand U5197 (N_5197,N_4886,N_4972);
nor U5198 (N_5198,N_4924,N_4762);
or U5199 (N_5199,N_4968,N_4877);
and U5200 (N_5200,N_4937,N_4935);
xor U5201 (N_5201,N_4895,N_4999);
and U5202 (N_5202,N_4920,N_4865);
or U5203 (N_5203,N_4822,N_4960);
nand U5204 (N_5204,N_4750,N_4824);
nand U5205 (N_5205,N_4930,N_4757);
or U5206 (N_5206,N_4978,N_4930);
nand U5207 (N_5207,N_4860,N_4877);
and U5208 (N_5208,N_4770,N_4854);
xnor U5209 (N_5209,N_4877,N_4981);
nor U5210 (N_5210,N_4781,N_4958);
or U5211 (N_5211,N_4781,N_4878);
xor U5212 (N_5212,N_4781,N_4999);
or U5213 (N_5213,N_4875,N_4940);
nor U5214 (N_5214,N_4768,N_4818);
or U5215 (N_5215,N_4781,N_4970);
xor U5216 (N_5216,N_4805,N_4789);
xor U5217 (N_5217,N_4762,N_4942);
or U5218 (N_5218,N_4753,N_4965);
or U5219 (N_5219,N_4949,N_4828);
and U5220 (N_5220,N_4956,N_4775);
nand U5221 (N_5221,N_4823,N_4938);
xor U5222 (N_5222,N_4905,N_4917);
and U5223 (N_5223,N_4843,N_4778);
and U5224 (N_5224,N_4994,N_4850);
xor U5225 (N_5225,N_4950,N_4906);
nand U5226 (N_5226,N_4906,N_4764);
nor U5227 (N_5227,N_4813,N_4983);
and U5228 (N_5228,N_4802,N_4902);
nor U5229 (N_5229,N_4791,N_4913);
nor U5230 (N_5230,N_4752,N_4850);
or U5231 (N_5231,N_4829,N_4975);
nor U5232 (N_5232,N_4792,N_4873);
nor U5233 (N_5233,N_4981,N_4888);
nand U5234 (N_5234,N_4935,N_4817);
nor U5235 (N_5235,N_4945,N_4987);
nor U5236 (N_5236,N_4794,N_4980);
or U5237 (N_5237,N_4877,N_4755);
nor U5238 (N_5238,N_4768,N_4845);
xor U5239 (N_5239,N_4773,N_4764);
and U5240 (N_5240,N_4966,N_4860);
nor U5241 (N_5241,N_4806,N_4935);
and U5242 (N_5242,N_4937,N_4896);
nor U5243 (N_5243,N_4850,N_4824);
or U5244 (N_5244,N_4968,N_4802);
nor U5245 (N_5245,N_4892,N_4893);
nand U5246 (N_5246,N_4827,N_4797);
nand U5247 (N_5247,N_4973,N_4889);
xor U5248 (N_5248,N_4888,N_4921);
nand U5249 (N_5249,N_4933,N_4785);
nor U5250 (N_5250,N_5199,N_5053);
nand U5251 (N_5251,N_5056,N_5145);
or U5252 (N_5252,N_5197,N_5228);
nand U5253 (N_5253,N_5013,N_5128);
nor U5254 (N_5254,N_5046,N_5232);
nand U5255 (N_5255,N_5047,N_5104);
xnor U5256 (N_5256,N_5155,N_5102);
nor U5257 (N_5257,N_5168,N_5236);
xnor U5258 (N_5258,N_5138,N_5066);
nand U5259 (N_5259,N_5044,N_5022);
or U5260 (N_5260,N_5078,N_5057);
nand U5261 (N_5261,N_5100,N_5045);
nor U5262 (N_5262,N_5216,N_5152);
or U5263 (N_5263,N_5079,N_5051);
or U5264 (N_5264,N_5076,N_5121);
and U5265 (N_5265,N_5245,N_5021);
nand U5266 (N_5266,N_5159,N_5088);
nand U5267 (N_5267,N_5202,N_5136);
xnor U5268 (N_5268,N_5081,N_5017);
xnor U5269 (N_5269,N_5118,N_5038);
or U5270 (N_5270,N_5032,N_5134);
or U5271 (N_5271,N_5082,N_5224);
nor U5272 (N_5272,N_5211,N_5083);
or U5273 (N_5273,N_5068,N_5043);
nand U5274 (N_5274,N_5109,N_5111);
nor U5275 (N_5275,N_5133,N_5163);
nor U5276 (N_5276,N_5037,N_5174);
xnor U5277 (N_5277,N_5167,N_5049);
nand U5278 (N_5278,N_5143,N_5129);
xor U5279 (N_5279,N_5119,N_5234);
and U5280 (N_5280,N_5220,N_5214);
nor U5281 (N_5281,N_5203,N_5001);
xor U5282 (N_5282,N_5026,N_5008);
xor U5283 (N_5283,N_5069,N_5120);
xor U5284 (N_5284,N_5229,N_5186);
xor U5285 (N_5285,N_5025,N_5180);
or U5286 (N_5286,N_5108,N_5183);
or U5287 (N_5287,N_5029,N_5091);
and U5288 (N_5288,N_5188,N_5060);
nor U5289 (N_5289,N_5178,N_5139);
or U5290 (N_5290,N_5052,N_5135);
and U5291 (N_5291,N_5089,N_5077);
or U5292 (N_5292,N_5141,N_5223);
nand U5293 (N_5293,N_5010,N_5005);
nor U5294 (N_5294,N_5248,N_5124);
nor U5295 (N_5295,N_5182,N_5030);
or U5296 (N_5296,N_5226,N_5099);
and U5297 (N_5297,N_5191,N_5189);
or U5298 (N_5298,N_5249,N_5115);
nor U5299 (N_5299,N_5222,N_5170);
and U5300 (N_5300,N_5192,N_5006);
nor U5301 (N_5301,N_5116,N_5075);
nand U5302 (N_5302,N_5065,N_5096);
and U5303 (N_5303,N_5034,N_5073);
or U5304 (N_5304,N_5090,N_5080);
xor U5305 (N_5305,N_5055,N_5208);
xor U5306 (N_5306,N_5114,N_5110);
or U5307 (N_5307,N_5103,N_5117);
and U5308 (N_5308,N_5185,N_5207);
or U5309 (N_5309,N_5106,N_5156);
nor U5310 (N_5310,N_5243,N_5169);
nand U5311 (N_5311,N_5071,N_5002);
nand U5312 (N_5312,N_5242,N_5126);
and U5313 (N_5313,N_5086,N_5209);
and U5314 (N_5314,N_5087,N_5070);
xnor U5315 (N_5315,N_5003,N_5140);
and U5316 (N_5316,N_5132,N_5101);
nand U5317 (N_5317,N_5042,N_5112);
or U5318 (N_5318,N_5195,N_5206);
and U5319 (N_5319,N_5107,N_5059);
and U5320 (N_5320,N_5122,N_5048);
or U5321 (N_5321,N_5062,N_5241);
and U5322 (N_5322,N_5011,N_5205);
nand U5323 (N_5323,N_5092,N_5004);
or U5324 (N_5324,N_5028,N_5039);
nand U5325 (N_5325,N_5105,N_5148);
xnor U5326 (N_5326,N_5181,N_5033);
and U5327 (N_5327,N_5130,N_5084);
xor U5328 (N_5328,N_5210,N_5215);
xor U5329 (N_5329,N_5064,N_5007);
xnor U5330 (N_5330,N_5160,N_5161);
nor U5331 (N_5331,N_5023,N_5217);
or U5332 (N_5332,N_5173,N_5157);
nor U5333 (N_5333,N_5014,N_5175);
or U5334 (N_5334,N_5000,N_5098);
and U5335 (N_5335,N_5018,N_5200);
or U5336 (N_5336,N_5050,N_5054);
or U5337 (N_5337,N_5012,N_5162);
nand U5338 (N_5338,N_5193,N_5176);
and U5339 (N_5339,N_5019,N_5063);
and U5340 (N_5340,N_5027,N_5237);
or U5341 (N_5341,N_5154,N_5230);
nand U5342 (N_5342,N_5238,N_5219);
and U5343 (N_5343,N_5009,N_5153);
nor U5344 (N_5344,N_5212,N_5198);
nand U5345 (N_5345,N_5016,N_5072);
nand U5346 (N_5346,N_5231,N_5172);
nor U5347 (N_5347,N_5179,N_5142);
nor U5348 (N_5348,N_5097,N_5094);
nor U5349 (N_5349,N_5225,N_5024);
nor U5350 (N_5350,N_5147,N_5235);
nor U5351 (N_5351,N_5213,N_5244);
xor U5352 (N_5352,N_5151,N_5158);
nor U5353 (N_5353,N_5058,N_5137);
nand U5354 (N_5354,N_5095,N_5093);
nand U5355 (N_5355,N_5127,N_5246);
or U5356 (N_5356,N_5146,N_5190);
nor U5357 (N_5357,N_5194,N_5196);
or U5358 (N_5358,N_5218,N_5036);
or U5359 (N_5359,N_5247,N_5085);
nand U5360 (N_5360,N_5125,N_5239);
nor U5361 (N_5361,N_5201,N_5204);
or U5362 (N_5362,N_5240,N_5020);
nand U5363 (N_5363,N_5074,N_5131);
or U5364 (N_5364,N_5171,N_5233);
nor U5365 (N_5365,N_5164,N_5015);
nand U5366 (N_5366,N_5123,N_5187);
xor U5367 (N_5367,N_5040,N_5227);
or U5368 (N_5368,N_5035,N_5165);
nand U5369 (N_5369,N_5150,N_5184);
and U5370 (N_5370,N_5113,N_5221);
and U5371 (N_5371,N_5067,N_5041);
and U5372 (N_5372,N_5166,N_5061);
nor U5373 (N_5373,N_5144,N_5031);
or U5374 (N_5374,N_5177,N_5149);
or U5375 (N_5375,N_5028,N_5149);
xor U5376 (N_5376,N_5066,N_5234);
or U5377 (N_5377,N_5048,N_5075);
nand U5378 (N_5378,N_5009,N_5225);
nand U5379 (N_5379,N_5063,N_5091);
nand U5380 (N_5380,N_5126,N_5173);
or U5381 (N_5381,N_5100,N_5099);
nor U5382 (N_5382,N_5185,N_5151);
and U5383 (N_5383,N_5113,N_5231);
or U5384 (N_5384,N_5183,N_5224);
and U5385 (N_5385,N_5040,N_5212);
and U5386 (N_5386,N_5227,N_5243);
or U5387 (N_5387,N_5078,N_5183);
xnor U5388 (N_5388,N_5168,N_5165);
nand U5389 (N_5389,N_5046,N_5098);
nand U5390 (N_5390,N_5104,N_5242);
xor U5391 (N_5391,N_5028,N_5089);
xor U5392 (N_5392,N_5245,N_5036);
and U5393 (N_5393,N_5158,N_5019);
nand U5394 (N_5394,N_5057,N_5196);
xnor U5395 (N_5395,N_5086,N_5072);
or U5396 (N_5396,N_5173,N_5187);
xnor U5397 (N_5397,N_5015,N_5199);
or U5398 (N_5398,N_5011,N_5221);
xor U5399 (N_5399,N_5015,N_5012);
and U5400 (N_5400,N_5040,N_5091);
and U5401 (N_5401,N_5167,N_5202);
nor U5402 (N_5402,N_5124,N_5058);
or U5403 (N_5403,N_5187,N_5071);
nand U5404 (N_5404,N_5049,N_5039);
nand U5405 (N_5405,N_5188,N_5185);
nand U5406 (N_5406,N_5025,N_5016);
nand U5407 (N_5407,N_5008,N_5058);
or U5408 (N_5408,N_5088,N_5009);
xor U5409 (N_5409,N_5184,N_5219);
xnor U5410 (N_5410,N_5067,N_5130);
nor U5411 (N_5411,N_5026,N_5087);
xnor U5412 (N_5412,N_5171,N_5226);
and U5413 (N_5413,N_5173,N_5067);
nor U5414 (N_5414,N_5169,N_5192);
and U5415 (N_5415,N_5040,N_5121);
or U5416 (N_5416,N_5008,N_5002);
or U5417 (N_5417,N_5247,N_5165);
xnor U5418 (N_5418,N_5057,N_5212);
nand U5419 (N_5419,N_5009,N_5087);
or U5420 (N_5420,N_5168,N_5077);
xnor U5421 (N_5421,N_5025,N_5134);
and U5422 (N_5422,N_5151,N_5239);
nor U5423 (N_5423,N_5234,N_5061);
and U5424 (N_5424,N_5047,N_5170);
and U5425 (N_5425,N_5214,N_5013);
and U5426 (N_5426,N_5067,N_5024);
and U5427 (N_5427,N_5127,N_5228);
nand U5428 (N_5428,N_5168,N_5152);
or U5429 (N_5429,N_5054,N_5097);
xor U5430 (N_5430,N_5007,N_5000);
or U5431 (N_5431,N_5172,N_5071);
and U5432 (N_5432,N_5032,N_5047);
and U5433 (N_5433,N_5034,N_5046);
or U5434 (N_5434,N_5065,N_5176);
and U5435 (N_5435,N_5152,N_5102);
and U5436 (N_5436,N_5194,N_5060);
or U5437 (N_5437,N_5249,N_5225);
xnor U5438 (N_5438,N_5137,N_5089);
xor U5439 (N_5439,N_5090,N_5095);
nand U5440 (N_5440,N_5042,N_5241);
xnor U5441 (N_5441,N_5159,N_5008);
nor U5442 (N_5442,N_5006,N_5074);
nand U5443 (N_5443,N_5158,N_5093);
and U5444 (N_5444,N_5025,N_5171);
and U5445 (N_5445,N_5067,N_5194);
and U5446 (N_5446,N_5073,N_5052);
nor U5447 (N_5447,N_5180,N_5192);
and U5448 (N_5448,N_5114,N_5028);
nand U5449 (N_5449,N_5059,N_5147);
xnor U5450 (N_5450,N_5153,N_5239);
and U5451 (N_5451,N_5148,N_5207);
and U5452 (N_5452,N_5045,N_5166);
and U5453 (N_5453,N_5105,N_5249);
or U5454 (N_5454,N_5067,N_5119);
and U5455 (N_5455,N_5184,N_5119);
nor U5456 (N_5456,N_5119,N_5037);
or U5457 (N_5457,N_5104,N_5194);
nor U5458 (N_5458,N_5198,N_5174);
xor U5459 (N_5459,N_5219,N_5053);
nand U5460 (N_5460,N_5035,N_5107);
and U5461 (N_5461,N_5240,N_5218);
and U5462 (N_5462,N_5123,N_5063);
or U5463 (N_5463,N_5029,N_5093);
or U5464 (N_5464,N_5208,N_5051);
or U5465 (N_5465,N_5217,N_5163);
xnor U5466 (N_5466,N_5115,N_5084);
and U5467 (N_5467,N_5071,N_5086);
or U5468 (N_5468,N_5130,N_5173);
and U5469 (N_5469,N_5174,N_5184);
nand U5470 (N_5470,N_5148,N_5126);
xor U5471 (N_5471,N_5009,N_5135);
nand U5472 (N_5472,N_5190,N_5115);
nand U5473 (N_5473,N_5104,N_5051);
nand U5474 (N_5474,N_5145,N_5047);
nand U5475 (N_5475,N_5235,N_5035);
xnor U5476 (N_5476,N_5138,N_5081);
nor U5477 (N_5477,N_5103,N_5182);
or U5478 (N_5478,N_5074,N_5227);
and U5479 (N_5479,N_5215,N_5092);
nand U5480 (N_5480,N_5231,N_5018);
or U5481 (N_5481,N_5202,N_5091);
xor U5482 (N_5482,N_5058,N_5077);
and U5483 (N_5483,N_5054,N_5149);
nand U5484 (N_5484,N_5135,N_5067);
or U5485 (N_5485,N_5011,N_5207);
and U5486 (N_5486,N_5169,N_5234);
xnor U5487 (N_5487,N_5099,N_5182);
xnor U5488 (N_5488,N_5000,N_5179);
and U5489 (N_5489,N_5082,N_5181);
xor U5490 (N_5490,N_5010,N_5071);
xnor U5491 (N_5491,N_5004,N_5082);
or U5492 (N_5492,N_5028,N_5178);
and U5493 (N_5493,N_5139,N_5200);
nand U5494 (N_5494,N_5188,N_5206);
nor U5495 (N_5495,N_5154,N_5059);
or U5496 (N_5496,N_5225,N_5020);
nor U5497 (N_5497,N_5161,N_5026);
nand U5498 (N_5498,N_5060,N_5079);
and U5499 (N_5499,N_5218,N_5091);
or U5500 (N_5500,N_5396,N_5308);
nor U5501 (N_5501,N_5393,N_5430);
xor U5502 (N_5502,N_5484,N_5400);
nand U5503 (N_5503,N_5419,N_5341);
nor U5504 (N_5504,N_5276,N_5386);
nor U5505 (N_5505,N_5280,N_5435);
and U5506 (N_5506,N_5267,N_5262);
nand U5507 (N_5507,N_5487,N_5494);
nor U5508 (N_5508,N_5277,N_5436);
or U5509 (N_5509,N_5472,N_5254);
and U5510 (N_5510,N_5368,N_5265);
xnor U5511 (N_5511,N_5356,N_5363);
nor U5512 (N_5512,N_5495,N_5404);
and U5513 (N_5513,N_5295,N_5311);
xor U5514 (N_5514,N_5474,N_5314);
xnor U5515 (N_5515,N_5471,N_5409);
or U5516 (N_5516,N_5446,N_5447);
or U5517 (N_5517,N_5458,N_5370);
xor U5518 (N_5518,N_5469,N_5310);
xnor U5519 (N_5519,N_5366,N_5344);
or U5520 (N_5520,N_5457,N_5492);
xnor U5521 (N_5521,N_5470,N_5428);
xnor U5522 (N_5522,N_5454,N_5362);
nor U5523 (N_5523,N_5281,N_5408);
nand U5524 (N_5524,N_5353,N_5395);
nor U5525 (N_5525,N_5388,N_5326);
nor U5526 (N_5526,N_5486,N_5445);
nand U5527 (N_5527,N_5429,N_5389);
nand U5528 (N_5528,N_5422,N_5273);
nand U5529 (N_5529,N_5288,N_5424);
nand U5530 (N_5530,N_5357,N_5320);
nor U5531 (N_5531,N_5421,N_5251);
xor U5532 (N_5532,N_5384,N_5338);
or U5533 (N_5533,N_5387,N_5425);
and U5534 (N_5534,N_5437,N_5323);
nand U5535 (N_5535,N_5352,N_5431);
nor U5536 (N_5536,N_5279,N_5383);
nand U5537 (N_5537,N_5259,N_5291);
or U5538 (N_5538,N_5371,N_5364);
nor U5539 (N_5539,N_5444,N_5334);
xnor U5540 (N_5540,N_5345,N_5432);
nor U5541 (N_5541,N_5459,N_5333);
and U5542 (N_5542,N_5415,N_5328);
and U5543 (N_5543,N_5339,N_5252);
xor U5544 (N_5544,N_5467,N_5305);
or U5545 (N_5545,N_5303,N_5282);
xor U5546 (N_5546,N_5453,N_5478);
nand U5547 (N_5547,N_5378,N_5496);
and U5548 (N_5548,N_5448,N_5325);
nand U5549 (N_5549,N_5296,N_5312);
and U5550 (N_5550,N_5485,N_5391);
or U5551 (N_5551,N_5330,N_5309);
and U5552 (N_5552,N_5442,N_5473);
or U5553 (N_5553,N_5475,N_5464);
nand U5554 (N_5554,N_5385,N_5406);
or U5555 (N_5555,N_5250,N_5272);
xnor U5556 (N_5556,N_5373,N_5275);
or U5557 (N_5557,N_5412,N_5441);
nor U5558 (N_5558,N_5375,N_5318);
nand U5559 (N_5559,N_5351,N_5263);
or U5560 (N_5560,N_5499,N_5337);
nor U5561 (N_5561,N_5369,N_5255);
nand U5562 (N_5562,N_5253,N_5315);
xor U5563 (N_5563,N_5423,N_5298);
xnor U5564 (N_5564,N_5460,N_5350);
and U5565 (N_5565,N_5342,N_5294);
or U5566 (N_5566,N_5331,N_5416);
or U5567 (N_5567,N_5477,N_5414);
and U5568 (N_5568,N_5482,N_5292);
nand U5569 (N_5569,N_5407,N_5376);
xor U5570 (N_5570,N_5380,N_5420);
nor U5571 (N_5571,N_5270,N_5443);
and U5572 (N_5572,N_5397,N_5427);
nor U5573 (N_5573,N_5271,N_5258);
xnor U5574 (N_5574,N_5299,N_5256);
nand U5575 (N_5575,N_5274,N_5257);
xnor U5576 (N_5576,N_5480,N_5285);
xnor U5577 (N_5577,N_5463,N_5367);
xor U5578 (N_5578,N_5372,N_5476);
nor U5579 (N_5579,N_5426,N_5462);
xor U5580 (N_5580,N_5481,N_5358);
xor U5581 (N_5581,N_5321,N_5402);
nand U5582 (N_5582,N_5479,N_5269);
nor U5583 (N_5583,N_5336,N_5266);
nor U5584 (N_5584,N_5403,N_5306);
nand U5585 (N_5585,N_5466,N_5483);
or U5586 (N_5586,N_5264,N_5491);
or U5587 (N_5587,N_5349,N_5451);
or U5588 (N_5588,N_5399,N_5489);
nand U5589 (N_5589,N_5390,N_5346);
nor U5590 (N_5590,N_5417,N_5410);
or U5591 (N_5591,N_5398,N_5348);
or U5592 (N_5592,N_5456,N_5335);
or U5593 (N_5593,N_5418,N_5405);
nor U5594 (N_5594,N_5332,N_5327);
nand U5595 (N_5595,N_5283,N_5359);
nand U5596 (N_5596,N_5468,N_5382);
nand U5597 (N_5597,N_5439,N_5284);
nor U5598 (N_5598,N_5455,N_5304);
nor U5599 (N_5599,N_5343,N_5278);
nand U5600 (N_5600,N_5461,N_5301);
nand U5601 (N_5601,N_5324,N_5261);
or U5602 (N_5602,N_5493,N_5497);
xor U5603 (N_5603,N_5360,N_5490);
nand U5604 (N_5604,N_5293,N_5379);
xor U5605 (N_5605,N_5329,N_5411);
and U5606 (N_5606,N_5268,N_5381);
or U5607 (N_5607,N_5319,N_5313);
nor U5608 (N_5608,N_5377,N_5354);
and U5609 (N_5609,N_5286,N_5465);
nor U5610 (N_5610,N_5450,N_5488);
xnor U5611 (N_5611,N_5433,N_5316);
and U5612 (N_5612,N_5413,N_5452);
xor U5613 (N_5613,N_5361,N_5498);
xnor U5614 (N_5614,N_5365,N_5302);
nand U5615 (N_5615,N_5322,N_5297);
xnor U5616 (N_5616,N_5394,N_5374);
nand U5617 (N_5617,N_5440,N_5340);
nor U5618 (N_5618,N_5289,N_5260);
and U5619 (N_5619,N_5347,N_5287);
xor U5620 (N_5620,N_5392,N_5290);
xor U5621 (N_5621,N_5438,N_5355);
nand U5622 (N_5622,N_5307,N_5434);
or U5623 (N_5623,N_5401,N_5317);
or U5624 (N_5624,N_5300,N_5449);
xor U5625 (N_5625,N_5340,N_5406);
nand U5626 (N_5626,N_5367,N_5402);
nor U5627 (N_5627,N_5417,N_5356);
or U5628 (N_5628,N_5464,N_5496);
or U5629 (N_5629,N_5424,N_5384);
or U5630 (N_5630,N_5331,N_5397);
or U5631 (N_5631,N_5433,N_5461);
nor U5632 (N_5632,N_5432,N_5435);
or U5633 (N_5633,N_5261,N_5417);
nand U5634 (N_5634,N_5406,N_5497);
xor U5635 (N_5635,N_5483,N_5481);
nand U5636 (N_5636,N_5304,N_5361);
xor U5637 (N_5637,N_5285,N_5366);
nor U5638 (N_5638,N_5312,N_5266);
and U5639 (N_5639,N_5381,N_5475);
or U5640 (N_5640,N_5295,N_5274);
nor U5641 (N_5641,N_5269,N_5371);
nand U5642 (N_5642,N_5388,N_5497);
xnor U5643 (N_5643,N_5284,N_5369);
and U5644 (N_5644,N_5259,N_5456);
nor U5645 (N_5645,N_5264,N_5300);
and U5646 (N_5646,N_5408,N_5367);
xnor U5647 (N_5647,N_5352,N_5300);
xor U5648 (N_5648,N_5483,N_5317);
or U5649 (N_5649,N_5387,N_5339);
or U5650 (N_5650,N_5460,N_5412);
or U5651 (N_5651,N_5413,N_5311);
nor U5652 (N_5652,N_5276,N_5361);
and U5653 (N_5653,N_5354,N_5420);
nand U5654 (N_5654,N_5318,N_5276);
and U5655 (N_5655,N_5378,N_5320);
or U5656 (N_5656,N_5499,N_5462);
nor U5657 (N_5657,N_5259,N_5258);
nand U5658 (N_5658,N_5462,N_5431);
or U5659 (N_5659,N_5495,N_5258);
and U5660 (N_5660,N_5337,N_5353);
xor U5661 (N_5661,N_5492,N_5405);
and U5662 (N_5662,N_5388,N_5279);
nand U5663 (N_5663,N_5412,N_5458);
and U5664 (N_5664,N_5417,N_5338);
and U5665 (N_5665,N_5347,N_5495);
and U5666 (N_5666,N_5442,N_5422);
nand U5667 (N_5667,N_5274,N_5459);
nor U5668 (N_5668,N_5258,N_5342);
or U5669 (N_5669,N_5274,N_5423);
nor U5670 (N_5670,N_5304,N_5394);
xnor U5671 (N_5671,N_5441,N_5353);
nand U5672 (N_5672,N_5370,N_5389);
or U5673 (N_5673,N_5380,N_5479);
nand U5674 (N_5674,N_5314,N_5367);
nand U5675 (N_5675,N_5378,N_5387);
nand U5676 (N_5676,N_5378,N_5278);
and U5677 (N_5677,N_5495,N_5497);
or U5678 (N_5678,N_5314,N_5483);
nand U5679 (N_5679,N_5487,N_5331);
nand U5680 (N_5680,N_5462,N_5312);
xnor U5681 (N_5681,N_5327,N_5252);
and U5682 (N_5682,N_5342,N_5315);
xnor U5683 (N_5683,N_5321,N_5455);
xnor U5684 (N_5684,N_5430,N_5391);
nand U5685 (N_5685,N_5347,N_5300);
nand U5686 (N_5686,N_5379,N_5448);
and U5687 (N_5687,N_5384,N_5317);
nor U5688 (N_5688,N_5312,N_5471);
nand U5689 (N_5689,N_5345,N_5332);
and U5690 (N_5690,N_5323,N_5341);
nand U5691 (N_5691,N_5357,N_5358);
nand U5692 (N_5692,N_5317,N_5430);
or U5693 (N_5693,N_5451,N_5467);
xor U5694 (N_5694,N_5369,N_5278);
xnor U5695 (N_5695,N_5443,N_5305);
nor U5696 (N_5696,N_5265,N_5277);
and U5697 (N_5697,N_5289,N_5466);
and U5698 (N_5698,N_5299,N_5435);
or U5699 (N_5699,N_5429,N_5397);
nor U5700 (N_5700,N_5456,N_5262);
xor U5701 (N_5701,N_5260,N_5471);
and U5702 (N_5702,N_5335,N_5492);
or U5703 (N_5703,N_5275,N_5452);
or U5704 (N_5704,N_5426,N_5253);
and U5705 (N_5705,N_5460,N_5440);
nand U5706 (N_5706,N_5377,N_5489);
and U5707 (N_5707,N_5376,N_5338);
nor U5708 (N_5708,N_5460,N_5262);
nand U5709 (N_5709,N_5281,N_5392);
xor U5710 (N_5710,N_5370,N_5351);
and U5711 (N_5711,N_5269,N_5398);
nand U5712 (N_5712,N_5411,N_5363);
and U5713 (N_5713,N_5393,N_5498);
nor U5714 (N_5714,N_5335,N_5327);
or U5715 (N_5715,N_5426,N_5403);
nor U5716 (N_5716,N_5452,N_5433);
nor U5717 (N_5717,N_5490,N_5486);
or U5718 (N_5718,N_5496,N_5473);
nand U5719 (N_5719,N_5466,N_5416);
xor U5720 (N_5720,N_5431,N_5331);
xnor U5721 (N_5721,N_5496,N_5321);
xor U5722 (N_5722,N_5315,N_5291);
and U5723 (N_5723,N_5480,N_5406);
nand U5724 (N_5724,N_5492,N_5401);
xor U5725 (N_5725,N_5493,N_5491);
or U5726 (N_5726,N_5434,N_5284);
nor U5727 (N_5727,N_5306,N_5451);
or U5728 (N_5728,N_5286,N_5336);
and U5729 (N_5729,N_5486,N_5431);
and U5730 (N_5730,N_5344,N_5424);
nor U5731 (N_5731,N_5360,N_5324);
or U5732 (N_5732,N_5332,N_5385);
or U5733 (N_5733,N_5299,N_5395);
nand U5734 (N_5734,N_5336,N_5351);
nand U5735 (N_5735,N_5332,N_5438);
nand U5736 (N_5736,N_5475,N_5307);
nor U5737 (N_5737,N_5308,N_5309);
and U5738 (N_5738,N_5322,N_5370);
and U5739 (N_5739,N_5422,N_5458);
nand U5740 (N_5740,N_5289,N_5453);
and U5741 (N_5741,N_5467,N_5402);
xnor U5742 (N_5742,N_5450,N_5469);
nand U5743 (N_5743,N_5392,N_5451);
and U5744 (N_5744,N_5385,N_5307);
xnor U5745 (N_5745,N_5437,N_5335);
nor U5746 (N_5746,N_5291,N_5281);
nor U5747 (N_5747,N_5436,N_5266);
xnor U5748 (N_5748,N_5453,N_5485);
nor U5749 (N_5749,N_5397,N_5483);
xnor U5750 (N_5750,N_5709,N_5581);
or U5751 (N_5751,N_5745,N_5699);
and U5752 (N_5752,N_5598,N_5654);
and U5753 (N_5753,N_5541,N_5509);
xnor U5754 (N_5754,N_5623,N_5528);
and U5755 (N_5755,N_5634,N_5588);
and U5756 (N_5756,N_5723,N_5696);
and U5757 (N_5757,N_5516,N_5635);
and U5758 (N_5758,N_5662,N_5626);
nand U5759 (N_5759,N_5684,N_5667);
nand U5760 (N_5760,N_5731,N_5584);
nand U5761 (N_5761,N_5737,N_5694);
nor U5762 (N_5762,N_5739,N_5610);
nor U5763 (N_5763,N_5736,N_5665);
or U5764 (N_5764,N_5695,N_5670);
xor U5765 (N_5765,N_5741,N_5674);
and U5766 (N_5766,N_5642,N_5513);
nand U5767 (N_5767,N_5624,N_5562);
xor U5768 (N_5768,N_5644,N_5543);
nor U5769 (N_5769,N_5548,N_5605);
nand U5770 (N_5770,N_5532,N_5568);
nor U5771 (N_5771,N_5565,N_5703);
and U5772 (N_5772,N_5726,N_5648);
and U5773 (N_5773,N_5746,N_5554);
nand U5774 (N_5774,N_5603,N_5666);
nand U5775 (N_5775,N_5614,N_5658);
and U5776 (N_5776,N_5560,N_5545);
nand U5777 (N_5777,N_5711,N_5531);
or U5778 (N_5778,N_5638,N_5551);
xnor U5779 (N_5779,N_5738,N_5563);
nor U5780 (N_5780,N_5688,N_5578);
and U5781 (N_5781,N_5725,N_5650);
and U5782 (N_5782,N_5673,N_5606);
and U5783 (N_5783,N_5587,N_5530);
nor U5784 (N_5784,N_5552,N_5722);
nand U5785 (N_5785,N_5525,N_5629);
or U5786 (N_5786,N_5529,N_5715);
nor U5787 (N_5787,N_5633,N_5660);
or U5788 (N_5788,N_5728,N_5564);
xor U5789 (N_5789,N_5717,N_5518);
and U5790 (N_5790,N_5628,N_5546);
nor U5791 (N_5791,N_5567,N_5727);
nand U5792 (N_5792,N_5502,N_5625);
xnor U5793 (N_5793,N_5539,N_5708);
and U5794 (N_5794,N_5580,N_5720);
xnor U5795 (N_5795,N_5514,N_5679);
or U5796 (N_5796,N_5713,N_5749);
xor U5797 (N_5797,N_5595,N_5575);
xor U5798 (N_5798,N_5542,N_5616);
or U5799 (N_5799,N_5707,N_5718);
or U5800 (N_5800,N_5651,N_5706);
nand U5801 (N_5801,N_5517,N_5577);
nor U5802 (N_5802,N_5590,N_5505);
nand U5803 (N_5803,N_5682,N_5724);
xor U5804 (N_5804,N_5639,N_5500);
nand U5805 (N_5805,N_5599,N_5557);
xor U5806 (N_5806,N_5604,N_5740);
or U5807 (N_5807,N_5680,N_5523);
nand U5808 (N_5808,N_5643,N_5600);
nor U5809 (N_5809,N_5574,N_5663);
nor U5810 (N_5810,N_5591,N_5632);
nor U5811 (N_5811,N_5555,N_5618);
nand U5812 (N_5812,N_5705,N_5671);
or U5813 (N_5813,N_5647,N_5748);
xor U5814 (N_5814,N_5556,N_5747);
nand U5815 (N_5815,N_5649,N_5710);
nor U5816 (N_5816,N_5550,N_5637);
nor U5817 (N_5817,N_5526,N_5571);
nor U5818 (N_5818,N_5656,N_5608);
nor U5819 (N_5819,N_5645,N_5596);
or U5820 (N_5820,N_5612,N_5655);
or U5821 (N_5821,N_5508,N_5646);
and U5822 (N_5822,N_5689,N_5735);
nand U5823 (N_5823,N_5686,N_5510);
xor U5824 (N_5824,N_5672,N_5621);
xnor U5825 (N_5825,N_5700,N_5630);
nor U5826 (N_5826,N_5619,N_5657);
nor U5827 (N_5827,N_5640,N_5573);
nand U5828 (N_5828,N_5566,N_5627);
xnor U5829 (N_5829,N_5693,N_5675);
and U5830 (N_5830,N_5572,N_5583);
and U5831 (N_5831,N_5631,N_5561);
xor U5832 (N_5832,N_5602,N_5714);
nor U5833 (N_5833,N_5538,N_5734);
or U5834 (N_5834,N_5540,N_5512);
and U5835 (N_5835,N_5636,N_5537);
nand U5836 (N_5836,N_5527,N_5582);
nor U5837 (N_5837,N_5730,N_5558);
or U5838 (N_5838,N_5594,N_5729);
and U5839 (N_5839,N_5524,N_5579);
nand U5840 (N_5840,N_5742,N_5677);
xor U5841 (N_5841,N_5501,N_5697);
xnor U5842 (N_5842,N_5585,N_5601);
and U5843 (N_5843,N_5534,N_5661);
nand U5844 (N_5844,N_5553,N_5622);
or U5845 (N_5845,N_5570,N_5664);
or U5846 (N_5846,N_5586,N_5690);
and U5847 (N_5847,N_5569,N_5533);
nor U5848 (N_5848,N_5615,N_5521);
or U5849 (N_5849,N_5597,N_5536);
nor U5850 (N_5850,N_5733,N_5712);
nand U5851 (N_5851,N_5511,N_5668);
or U5852 (N_5852,N_5609,N_5743);
or U5853 (N_5853,N_5692,N_5515);
nor U5854 (N_5854,N_5506,N_5698);
xor U5855 (N_5855,N_5589,N_5611);
xnor U5856 (N_5856,N_5520,N_5702);
nand U5857 (N_5857,N_5522,N_5613);
or U5858 (N_5858,N_5592,N_5691);
and U5859 (N_5859,N_5676,N_5685);
or U5860 (N_5860,N_5744,N_5659);
and U5861 (N_5861,N_5519,N_5701);
and U5862 (N_5862,N_5716,N_5678);
xnor U5863 (N_5863,N_5683,N_5732);
nor U5864 (N_5864,N_5503,N_5544);
or U5865 (N_5865,N_5576,N_5504);
or U5866 (N_5866,N_5507,N_5687);
nor U5867 (N_5867,N_5641,N_5607);
or U5868 (N_5868,N_5617,N_5669);
nor U5869 (N_5869,N_5653,N_5535);
nand U5870 (N_5870,N_5681,N_5704);
nor U5871 (N_5871,N_5719,N_5652);
nand U5872 (N_5872,N_5620,N_5721);
xnor U5873 (N_5873,N_5593,N_5549);
nor U5874 (N_5874,N_5547,N_5559);
nand U5875 (N_5875,N_5624,N_5505);
xnor U5876 (N_5876,N_5672,N_5704);
or U5877 (N_5877,N_5610,N_5646);
xnor U5878 (N_5878,N_5564,N_5603);
or U5879 (N_5879,N_5666,N_5618);
xnor U5880 (N_5880,N_5737,N_5558);
and U5881 (N_5881,N_5658,N_5727);
or U5882 (N_5882,N_5588,N_5601);
or U5883 (N_5883,N_5652,N_5698);
xor U5884 (N_5884,N_5663,N_5660);
or U5885 (N_5885,N_5548,N_5541);
xnor U5886 (N_5886,N_5684,N_5530);
or U5887 (N_5887,N_5703,N_5628);
and U5888 (N_5888,N_5597,N_5723);
nand U5889 (N_5889,N_5507,N_5512);
nand U5890 (N_5890,N_5682,N_5568);
and U5891 (N_5891,N_5630,N_5690);
nor U5892 (N_5892,N_5653,N_5564);
nor U5893 (N_5893,N_5724,N_5586);
or U5894 (N_5894,N_5552,N_5632);
and U5895 (N_5895,N_5561,N_5539);
nand U5896 (N_5896,N_5552,N_5652);
nand U5897 (N_5897,N_5526,N_5695);
nand U5898 (N_5898,N_5627,N_5548);
nand U5899 (N_5899,N_5586,N_5536);
and U5900 (N_5900,N_5585,N_5573);
xor U5901 (N_5901,N_5518,N_5529);
nand U5902 (N_5902,N_5607,N_5736);
nand U5903 (N_5903,N_5563,N_5648);
or U5904 (N_5904,N_5631,N_5605);
nand U5905 (N_5905,N_5572,N_5500);
and U5906 (N_5906,N_5543,N_5564);
or U5907 (N_5907,N_5714,N_5715);
nor U5908 (N_5908,N_5720,N_5730);
nor U5909 (N_5909,N_5696,N_5518);
nand U5910 (N_5910,N_5662,N_5693);
nor U5911 (N_5911,N_5559,N_5689);
nand U5912 (N_5912,N_5638,N_5518);
and U5913 (N_5913,N_5691,N_5658);
xor U5914 (N_5914,N_5539,N_5597);
xnor U5915 (N_5915,N_5664,N_5597);
nor U5916 (N_5916,N_5713,N_5536);
or U5917 (N_5917,N_5514,N_5555);
nand U5918 (N_5918,N_5651,N_5742);
and U5919 (N_5919,N_5650,N_5593);
and U5920 (N_5920,N_5529,N_5627);
and U5921 (N_5921,N_5667,N_5716);
xnor U5922 (N_5922,N_5503,N_5658);
or U5923 (N_5923,N_5517,N_5520);
and U5924 (N_5924,N_5716,N_5573);
nor U5925 (N_5925,N_5698,N_5573);
or U5926 (N_5926,N_5567,N_5549);
nor U5927 (N_5927,N_5566,N_5554);
nand U5928 (N_5928,N_5603,N_5706);
nor U5929 (N_5929,N_5685,N_5684);
nor U5930 (N_5930,N_5749,N_5688);
nor U5931 (N_5931,N_5676,N_5624);
nand U5932 (N_5932,N_5537,N_5746);
and U5933 (N_5933,N_5646,N_5637);
or U5934 (N_5934,N_5564,N_5546);
or U5935 (N_5935,N_5502,N_5559);
xnor U5936 (N_5936,N_5550,N_5560);
and U5937 (N_5937,N_5673,N_5727);
and U5938 (N_5938,N_5619,N_5501);
or U5939 (N_5939,N_5733,N_5666);
or U5940 (N_5940,N_5513,N_5715);
nor U5941 (N_5941,N_5652,N_5691);
nand U5942 (N_5942,N_5605,N_5575);
or U5943 (N_5943,N_5590,N_5528);
and U5944 (N_5944,N_5529,N_5517);
nand U5945 (N_5945,N_5558,N_5597);
xnor U5946 (N_5946,N_5526,N_5531);
or U5947 (N_5947,N_5658,N_5700);
nand U5948 (N_5948,N_5520,N_5710);
xor U5949 (N_5949,N_5639,N_5721);
nor U5950 (N_5950,N_5651,N_5620);
nor U5951 (N_5951,N_5614,N_5664);
xor U5952 (N_5952,N_5590,N_5622);
nor U5953 (N_5953,N_5674,N_5634);
and U5954 (N_5954,N_5657,N_5578);
and U5955 (N_5955,N_5635,N_5503);
nand U5956 (N_5956,N_5700,N_5684);
nor U5957 (N_5957,N_5657,N_5736);
nor U5958 (N_5958,N_5591,N_5526);
nand U5959 (N_5959,N_5732,N_5687);
xor U5960 (N_5960,N_5719,N_5686);
xor U5961 (N_5961,N_5611,N_5677);
and U5962 (N_5962,N_5746,N_5705);
nand U5963 (N_5963,N_5664,N_5533);
nand U5964 (N_5964,N_5657,N_5535);
and U5965 (N_5965,N_5514,N_5662);
xnor U5966 (N_5966,N_5731,N_5505);
nand U5967 (N_5967,N_5508,N_5737);
xor U5968 (N_5968,N_5639,N_5584);
xor U5969 (N_5969,N_5730,N_5572);
or U5970 (N_5970,N_5541,N_5511);
and U5971 (N_5971,N_5509,N_5530);
xor U5972 (N_5972,N_5691,N_5711);
and U5973 (N_5973,N_5588,N_5737);
or U5974 (N_5974,N_5501,N_5730);
and U5975 (N_5975,N_5589,N_5692);
nor U5976 (N_5976,N_5744,N_5598);
xnor U5977 (N_5977,N_5667,N_5717);
and U5978 (N_5978,N_5507,N_5611);
nor U5979 (N_5979,N_5607,N_5553);
and U5980 (N_5980,N_5718,N_5665);
or U5981 (N_5981,N_5502,N_5618);
and U5982 (N_5982,N_5564,N_5716);
and U5983 (N_5983,N_5647,N_5598);
xnor U5984 (N_5984,N_5609,N_5683);
or U5985 (N_5985,N_5545,N_5513);
nor U5986 (N_5986,N_5625,N_5561);
xnor U5987 (N_5987,N_5571,N_5649);
or U5988 (N_5988,N_5547,N_5736);
and U5989 (N_5989,N_5639,N_5619);
xnor U5990 (N_5990,N_5668,N_5728);
nor U5991 (N_5991,N_5741,N_5573);
nand U5992 (N_5992,N_5558,N_5561);
and U5993 (N_5993,N_5587,N_5715);
nand U5994 (N_5994,N_5670,N_5684);
xnor U5995 (N_5995,N_5734,N_5596);
nor U5996 (N_5996,N_5687,N_5551);
or U5997 (N_5997,N_5560,N_5747);
xor U5998 (N_5998,N_5584,N_5553);
and U5999 (N_5999,N_5680,N_5667);
and U6000 (N_6000,N_5950,N_5895);
xor U6001 (N_6001,N_5798,N_5915);
and U6002 (N_6002,N_5960,N_5826);
nand U6003 (N_6003,N_5780,N_5973);
and U6004 (N_6004,N_5977,N_5864);
or U6005 (N_6005,N_5843,N_5754);
and U6006 (N_6006,N_5876,N_5980);
and U6007 (N_6007,N_5800,N_5900);
nor U6008 (N_6008,N_5778,N_5933);
xor U6009 (N_6009,N_5914,N_5878);
or U6010 (N_6010,N_5954,N_5777);
and U6011 (N_6011,N_5956,N_5987);
nor U6012 (N_6012,N_5814,N_5852);
nor U6013 (N_6013,N_5926,N_5896);
xor U6014 (N_6014,N_5993,N_5775);
nor U6015 (N_6015,N_5982,N_5804);
nand U6016 (N_6016,N_5851,N_5967);
nor U6017 (N_6017,N_5953,N_5809);
and U6018 (N_6018,N_5847,N_5881);
and U6019 (N_6019,N_5856,N_5840);
nor U6020 (N_6020,N_5825,N_5751);
nor U6021 (N_6021,N_5867,N_5998);
or U6022 (N_6022,N_5885,N_5916);
nand U6023 (N_6023,N_5909,N_5970);
and U6024 (N_6024,N_5795,N_5952);
or U6025 (N_6025,N_5925,N_5874);
and U6026 (N_6026,N_5964,N_5822);
xnor U6027 (N_6027,N_5877,N_5893);
xnor U6028 (N_6028,N_5784,N_5765);
or U6029 (N_6029,N_5943,N_5860);
nand U6030 (N_6030,N_5978,N_5756);
xor U6031 (N_6031,N_5892,N_5966);
or U6032 (N_6032,N_5946,N_5894);
xnor U6033 (N_6033,N_5997,N_5919);
and U6034 (N_6034,N_5924,N_5979);
or U6035 (N_6035,N_5813,N_5757);
xor U6036 (N_6036,N_5759,N_5986);
nor U6037 (N_6037,N_5853,N_5969);
nand U6038 (N_6038,N_5808,N_5988);
nor U6039 (N_6039,N_5769,N_5974);
nand U6040 (N_6040,N_5831,N_5790);
and U6041 (N_6041,N_5955,N_5806);
nand U6042 (N_6042,N_5761,N_5959);
nor U6043 (N_6043,N_5810,N_5930);
xor U6044 (N_6044,N_5802,N_5752);
nand U6045 (N_6045,N_5935,N_5891);
and U6046 (N_6046,N_5844,N_5971);
nor U6047 (N_6047,N_5842,N_5990);
and U6048 (N_6048,N_5942,N_5797);
or U6049 (N_6049,N_5849,N_5927);
or U6050 (N_6050,N_5995,N_5920);
nor U6051 (N_6051,N_5898,N_5968);
xnor U6052 (N_6052,N_5932,N_5815);
nor U6053 (N_6053,N_5833,N_5755);
or U6054 (N_6054,N_5817,N_5934);
nand U6055 (N_6055,N_5962,N_5903);
nor U6056 (N_6056,N_5855,N_5766);
and U6057 (N_6057,N_5904,N_5828);
nor U6058 (N_6058,N_5873,N_5886);
xnor U6059 (N_6059,N_5949,N_5807);
or U6060 (N_6060,N_5910,N_5936);
nand U6061 (N_6061,N_5792,N_5911);
and U6062 (N_6062,N_5989,N_5791);
or U6063 (N_6063,N_5803,N_5999);
nor U6064 (N_6064,N_5923,N_5753);
nand U6065 (N_6065,N_5846,N_5981);
or U6066 (N_6066,N_5805,N_5768);
and U6067 (N_6067,N_5829,N_5848);
nand U6068 (N_6068,N_5912,N_5882);
or U6069 (N_6069,N_5845,N_5870);
nor U6070 (N_6070,N_5830,N_5782);
xnor U6071 (N_6071,N_5996,N_5901);
nand U6072 (N_6072,N_5890,N_5834);
and U6073 (N_6073,N_5972,N_5868);
and U6074 (N_6074,N_5963,N_5992);
nand U6075 (N_6075,N_5779,N_5794);
nor U6076 (N_6076,N_5947,N_5839);
xnor U6077 (N_6077,N_5859,N_5783);
nor U6078 (N_6078,N_5945,N_5760);
nor U6079 (N_6079,N_5850,N_5832);
or U6080 (N_6080,N_5793,N_5965);
nor U6081 (N_6081,N_5957,N_5799);
and U6082 (N_6082,N_5824,N_5863);
xor U6083 (N_6083,N_5875,N_5883);
nor U6084 (N_6084,N_5884,N_5788);
and U6085 (N_6085,N_5819,N_5994);
xor U6086 (N_6086,N_5944,N_5958);
nand U6087 (N_6087,N_5871,N_5812);
and U6088 (N_6088,N_5938,N_5917);
nor U6089 (N_6089,N_5820,N_5771);
nand U6090 (N_6090,N_5776,N_5928);
and U6091 (N_6091,N_5816,N_5789);
xor U6092 (N_6092,N_5907,N_5818);
or U6093 (N_6093,N_5902,N_5836);
and U6094 (N_6094,N_5906,N_5931);
and U6095 (N_6095,N_5975,N_5905);
nor U6096 (N_6096,N_5835,N_5869);
nand U6097 (N_6097,N_5889,N_5948);
nand U6098 (N_6098,N_5858,N_5991);
or U6099 (N_6099,N_5880,N_5862);
or U6100 (N_6100,N_5940,N_5921);
xor U6101 (N_6101,N_5888,N_5861);
and U6102 (N_6102,N_5764,N_5854);
or U6103 (N_6103,N_5937,N_5796);
nand U6104 (N_6104,N_5801,N_5774);
nand U6105 (N_6105,N_5929,N_5786);
or U6106 (N_6106,N_5951,N_5787);
or U6107 (N_6107,N_5821,N_5785);
and U6108 (N_6108,N_5837,N_5976);
or U6109 (N_6109,N_5899,N_5872);
or U6110 (N_6110,N_5913,N_5823);
nor U6111 (N_6111,N_5879,N_5918);
or U6112 (N_6112,N_5781,N_5983);
nor U6113 (N_6113,N_5841,N_5985);
nand U6114 (N_6114,N_5811,N_5770);
xnor U6115 (N_6115,N_5887,N_5941);
and U6116 (N_6116,N_5857,N_5772);
xor U6117 (N_6117,N_5838,N_5922);
nor U6118 (N_6118,N_5758,N_5767);
and U6119 (N_6119,N_5908,N_5897);
xnor U6120 (N_6120,N_5865,N_5763);
and U6121 (N_6121,N_5773,N_5939);
nor U6122 (N_6122,N_5762,N_5750);
nor U6123 (N_6123,N_5827,N_5866);
or U6124 (N_6124,N_5961,N_5984);
nor U6125 (N_6125,N_5885,N_5810);
nand U6126 (N_6126,N_5857,N_5798);
nor U6127 (N_6127,N_5907,N_5813);
and U6128 (N_6128,N_5892,N_5846);
nor U6129 (N_6129,N_5902,N_5948);
nor U6130 (N_6130,N_5870,N_5916);
nand U6131 (N_6131,N_5848,N_5841);
and U6132 (N_6132,N_5773,N_5814);
or U6133 (N_6133,N_5994,N_5959);
xor U6134 (N_6134,N_5913,N_5923);
nand U6135 (N_6135,N_5819,N_5826);
nor U6136 (N_6136,N_5822,N_5771);
and U6137 (N_6137,N_5872,N_5969);
or U6138 (N_6138,N_5931,N_5878);
nor U6139 (N_6139,N_5919,N_5813);
or U6140 (N_6140,N_5954,N_5896);
nand U6141 (N_6141,N_5921,N_5891);
and U6142 (N_6142,N_5775,N_5969);
xor U6143 (N_6143,N_5975,N_5993);
nand U6144 (N_6144,N_5815,N_5942);
xnor U6145 (N_6145,N_5818,N_5967);
nand U6146 (N_6146,N_5782,N_5863);
xnor U6147 (N_6147,N_5925,N_5967);
xor U6148 (N_6148,N_5771,N_5762);
nor U6149 (N_6149,N_5962,N_5980);
nor U6150 (N_6150,N_5942,N_5847);
nor U6151 (N_6151,N_5835,N_5756);
nor U6152 (N_6152,N_5801,N_5809);
nand U6153 (N_6153,N_5880,N_5990);
nand U6154 (N_6154,N_5843,N_5830);
and U6155 (N_6155,N_5800,N_5964);
or U6156 (N_6156,N_5901,N_5952);
or U6157 (N_6157,N_5838,N_5900);
and U6158 (N_6158,N_5865,N_5833);
nor U6159 (N_6159,N_5973,N_5841);
or U6160 (N_6160,N_5899,N_5849);
nand U6161 (N_6161,N_5913,N_5863);
or U6162 (N_6162,N_5919,N_5856);
and U6163 (N_6163,N_5832,N_5929);
xnor U6164 (N_6164,N_5904,N_5917);
and U6165 (N_6165,N_5958,N_5968);
xor U6166 (N_6166,N_5841,N_5824);
or U6167 (N_6167,N_5850,N_5971);
nand U6168 (N_6168,N_5974,N_5835);
or U6169 (N_6169,N_5776,N_5874);
or U6170 (N_6170,N_5969,N_5783);
nor U6171 (N_6171,N_5786,N_5956);
xnor U6172 (N_6172,N_5954,N_5907);
or U6173 (N_6173,N_5823,N_5779);
or U6174 (N_6174,N_5794,N_5944);
or U6175 (N_6175,N_5823,N_5958);
nand U6176 (N_6176,N_5877,N_5853);
nor U6177 (N_6177,N_5767,N_5751);
nand U6178 (N_6178,N_5809,N_5891);
or U6179 (N_6179,N_5826,N_5779);
nand U6180 (N_6180,N_5819,N_5871);
nor U6181 (N_6181,N_5910,N_5773);
or U6182 (N_6182,N_5750,N_5967);
nand U6183 (N_6183,N_5778,N_5961);
xor U6184 (N_6184,N_5919,N_5911);
nand U6185 (N_6185,N_5887,N_5969);
or U6186 (N_6186,N_5876,N_5767);
or U6187 (N_6187,N_5892,N_5878);
nand U6188 (N_6188,N_5758,N_5859);
nor U6189 (N_6189,N_5758,N_5787);
xor U6190 (N_6190,N_5853,N_5933);
or U6191 (N_6191,N_5993,N_5904);
nor U6192 (N_6192,N_5891,N_5944);
nand U6193 (N_6193,N_5781,N_5795);
or U6194 (N_6194,N_5810,N_5902);
and U6195 (N_6195,N_5832,N_5827);
nor U6196 (N_6196,N_5756,N_5825);
or U6197 (N_6197,N_5808,N_5921);
nand U6198 (N_6198,N_5827,N_5999);
nand U6199 (N_6199,N_5899,N_5901);
nand U6200 (N_6200,N_5877,N_5902);
and U6201 (N_6201,N_5858,N_5813);
nor U6202 (N_6202,N_5901,N_5909);
or U6203 (N_6203,N_5966,N_5960);
nor U6204 (N_6204,N_5917,N_5973);
nand U6205 (N_6205,N_5798,N_5926);
and U6206 (N_6206,N_5899,N_5827);
nor U6207 (N_6207,N_5845,N_5981);
nor U6208 (N_6208,N_5991,N_5949);
or U6209 (N_6209,N_5836,N_5752);
nor U6210 (N_6210,N_5965,N_5845);
and U6211 (N_6211,N_5769,N_5767);
nand U6212 (N_6212,N_5885,N_5943);
or U6213 (N_6213,N_5781,N_5873);
and U6214 (N_6214,N_5940,N_5795);
and U6215 (N_6215,N_5798,N_5906);
nand U6216 (N_6216,N_5856,N_5774);
or U6217 (N_6217,N_5891,N_5772);
and U6218 (N_6218,N_5871,N_5833);
and U6219 (N_6219,N_5796,N_5891);
nor U6220 (N_6220,N_5797,N_5909);
nand U6221 (N_6221,N_5968,N_5996);
nand U6222 (N_6222,N_5927,N_5864);
nand U6223 (N_6223,N_5834,N_5753);
or U6224 (N_6224,N_5989,N_5773);
and U6225 (N_6225,N_5897,N_5947);
xor U6226 (N_6226,N_5906,N_5846);
and U6227 (N_6227,N_5850,N_5997);
xor U6228 (N_6228,N_5788,N_5752);
nand U6229 (N_6229,N_5873,N_5955);
nor U6230 (N_6230,N_5930,N_5962);
nor U6231 (N_6231,N_5973,N_5912);
nor U6232 (N_6232,N_5887,N_5899);
and U6233 (N_6233,N_5773,N_5962);
nor U6234 (N_6234,N_5984,N_5822);
nand U6235 (N_6235,N_5789,N_5911);
nor U6236 (N_6236,N_5876,N_5935);
nor U6237 (N_6237,N_5973,N_5750);
and U6238 (N_6238,N_5923,N_5938);
nand U6239 (N_6239,N_5829,N_5801);
and U6240 (N_6240,N_5776,N_5956);
and U6241 (N_6241,N_5917,N_5944);
or U6242 (N_6242,N_5773,N_5835);
nand U6243 (N_6243,N_5946,N_5978);
xnor U6244 (N_6244,N_5802,N_5898);
and U6245 (N_6245,N_5823,N_5775);
nor U6246 (N_6246,N_5830,N_5818);
or U6247 (N_6247,N_5780,N_5971);
xor U6248 (N_6248,N_5932,N_5907);
or U6249 (N_6249,N_5928,N_5930);
nor U6250 (N_6250,N_6218,N_6017);
or U6251 (N_6251,N_6075,N_6027);
nand U6252 (N_6252,N_6214,N_6106);
xor U6253 (N_6253,N_6217,N_6015);
nor U6254 (N_6254,N_6215,N_6105);
nor U6255 (N_6255,N_6048,N_6042);
nor U6256 (N_6256,N_6120,N_6131);
nand U6257 (N_6257,N_6158,N_6138);
nor U6258 (N_6258,N_6237,N_6087);
and U6259 (N_6259,N_6177,N_6242);
and U6260 (N_6260,N_6078,N_6047);
nand U6261 (N_6261,N_6189,N_6225);
nor U6262 (N_6262,N_6073,N_6179);
nand U6263 (N_6263,N_6039,N_6141);
or U6264 (N_6264,N_6228,N_6056);
or U6265 (N_6265,N_6031,N_6003);
nand U6266 (N_6266,N_6132,N_6170);
xor U6267 (N_6267,N_6098,N_6109);
nor U6268 (N_6268,N_6139,N_6057);
nor U6269 (N_6269,N_6033,N_6050);
or U6270 (N_6270,N_6197,N_6148);
and U6271 (N_6271,N_6239,N_6174);
or U6272 (N_6272,N_6081,N_6146);
and U6273 (N_6273,N_6240,N_6021);
xnor U6274 (N_6274,N_6200,N_6084);
and U6275 (N_6275,N_6180,N_6101);
xor U6276 (N_6276,N_6032,N_6066);
nor U6277 (N_6277,N_6199,N_6088);
and U6278 (N_6278,N_6072,N_6061);
nor U6279 (N_6279,N_6187,N_6007);
nor U6280 (N_6280,N_6096,N_6128);
nor U6281 (N_6281,N_6082,N_6207);
xnor U6282 (N_6282,N_6247,N_6059);
and U6283 (N_6283,N_6165,N_6183);
or U6284 (N_6284,N_6012,N_6150);
nor U6285 (N_6285,N_6094,N_6034);
xor U6286 (N_6286,N_6010,N_6029);
xor U6287 (N_6287,N_6112,N_6164);
or U6288 (N_6288,N_6091,N_6244);
and U6289 (N_6289,N_6016,N_6086);
or U6290 (N_6290,N_6245,N_6137);
nor U6291 (N_6291,N_6172,N_6142);
xor U6292 (N_6292,N_6102,N_6014);
and U6293 (N_6293,N_6219,N_6206);
and U6294 (N_6294,N_6001,N_6005);
or U6295 (N_6295,N_6117,N_6157);
nand U6296 (N_6296,N_6114,N_6103);
and U6297 (N_6297,N_6224,N_6230);
xnor U6298 (N_6298,N_6008,N_6093);
and U6299 (N_6299,N_6169,N_6104);
nand U6300 (N_6300,N_6036,N_6037);
or U6301 (N_6301,N_6249,N_6045);
or U6302 (N_6302,N_6205,N_6004);
nor U6303 (N_6303,N_6220,N_6231);
nand U6304 (N_6304,N_6153,N_6018);
xnor U6305 (N_6305,N_6130,N_6019);
xor U6306 (N_6306,N_6175,N_6182);
nand U6307 (N_6307,N_6166,N_6108);
nor U6308 (N_6308,N_6176,N_6089);
or U6309 (N_6309,N_6127,N_6213);
nor U6310 (N_6310,N_6063,N_6122);
and U6311 (N_6311,N_6229,N_6188);
nor U6312 (N_6312,N_6079,N_6196);
nor U6313 (N_6313,N_6080,N_6178);
and U6314 (N_6314,N_6092,N_6136);
nand U6315 (N_6315,N_6192,N_6025);
and U6316 (N_6316,N_6099,N_6083);
nor U6317 (N_6317,N_6155,N_6216);
or U6318 (N_6318,N_6134,N_6168);
xor U6319 (N_6319,N_6152,N_6121);
nor U6320 (N_6320,N_6062,N_6248);
nand U6321 (N_6321,N_6065,N_6233);
and U6322 (N_6322,N_6210,N_6203);
and U6323 (N_6323,N_6043,N_6013);
or U6324 (N_6324,N_6100,N_6191);
nor U6325 (N_6325,N_6069,N_6195);
nand U6326 (N_6326,N_6038,N_6173);
or U6327 (N_6327,N_6185,N_6208);
and U6328 (N_6328,N_6115,N_6044);
or U6329 (N_6329,N_6000,N_6041);
nand U6330 (N_6330,N_6133,N_6171);
or U6331 (N_6331,N_6194,N_6006);
nand U6332 (N_6332,N_6211,N_6028);
or U6333 (N_6333,N_6024,N_6160);
or U6334 (N_6334,N_6223,N_6035);
xnor U6335 (N_6335,N_6124,N_6147);
and U6336 (N_6336,N_6054,N_6209);
nor U6337 (N_6337,N_6140,N_6159);
and U6338 (N_6338,N_6184,N_6161);
nand U6339 (N_6339,N_6118,N_6090);
nor U6340 (N_6340,N_6111,N_6064);
nand U6341 (N_6341,N_6167,N_6151);
or U6342 (N_6342,N_6156,N_6235);
nand U6343 (N_6343,N_6107,N_6058);
or U6344 (N_6344,N_6222,N_6110);
nand U6345 (N_6345,N_6046,N_6049);
or U6346 (N_6346,N_6246,N_6076);
or U6347 (N_6347,N_6129,N_6011);
nand U6348 (N_6348,N_6113,N_6162);
or U6349 (N_6349,N_6055,N_6067);
nand U6350 (N_6350,N_6238,N_6026);
nand U6351 (N_6351,N_6085,N_6212);
or U6352 (N_6352,N_6236,N_6241);
nor U6353 (N_6353,N_6154,N_6202);
xor U6354 (N_6354,N_6125,N_6074);
nand U6355 (N_6355,N_6071,N_6226);
and U6356 (N_6356,N_6040,N_6190);
and U6357 (N_6357,N_6002,N_6135);
nor U6358 (N_6358,N_6051,N_6095);
nand U6359 (N_6359,N_6022,N_6116);
or U6360 (N_6360,N_6009,N_6204);
nand U6361 (N_6361,N_6232,N_6186);
or U6362 (N_6362,N_6181,N_6119);
nand U6363 (N_6363,N_6053,N_6227);
xnor U6364 (N_6364,N_6144,N_6052);
xor U6365 (N_6365,N_6149,N_6234);
nor U6366 (N_6366,N_6193,N_6163);
nor U6367 (N_6367,N_6077,N_6097);
nor U6368 (N_6368,N_6030,N_6070);
and U6369 (N_6369,N_6198,N_6143);
and U6370 (N_6370,N_6243,N_6060);
nand U6371 (N_6371,N_6221,N_6145);
or U6372 (N_6372,N_6201,N_6123);
and U6373 (N_6373,N_6126,N_6068);
nor U6374 (N_6374,N_6023,N_6020);
and U6375 (N_6375,N_6045,N_6221);
nand U6376 (N_6376,N_6015,N_6070);
xor U6377 (N_6377,N_6093,N_6127);
nand U6378 (N_6378,N_6181,N_6061);
nand U6379 (N_6379,N_6043,N_6128);
nor U6380 (N_6380,N_6153,N_6182);
and U6381 (N_6381,N_6019,N_6028);
nor U6382 (N_6382,N_6056,N_6226);
xor U6383 (N_6383,N_6152,N_6123);
xnor U6384 (N_6384,N_6205,N_6131);
xor U6385 (N_6385,N_6213,N_6192);
xor U6386 (N_6386,N_6101,N_6131);
xnor U6387 (N_6387,N_6068,N_6237);
or U6388 (N_6388,N_6228,N_6207);
nor U6389 (N_6389,N_6203,N_6145);
or U6390 (N_6390,N_6153,N_6207);
and U6391 (N_6391,N_6149,N_6207);
and U6392 (N_6392,N_6065,N_6026);
nor U6393 (N_6393,N_6072,N_6080);
nand U6394 (N_6394,N_6090,N_6233);
nand U6395 (N_6395,N_6236,N_6152);
nor U6396 (N_6396,N_6222,N_6183);
nor U6397 (N_6397,N_6049,N_6148);
or U6398 (N_6398,N_6199,N_6231);
nor U6399 (N_6399,N_6093,N_6156);
xnor U6400 (N_6400,N_6236,N_6100);
xor U6401 (N_6401,N_6015,N_6249);
nand U6402 (N_6402,N_6142,N_6204);
and U6403 (N_6403,N_6171,N_6192);
xor U6404 (N_6404,N_6084,N_6071);
nor U6405 (N_6405,N_6225,N_6230);
nand U6406 (N_6406,N_6032,N_6246);
xor U6407 (N_6407,N_6194,N_6138);
and U6408 (N_6408,N_6221,N_6014);
nor U6409 (N_6409,N_6087,N_6120);
nor U6410 (N_6410,N_6120,N_6221);
nand U6411 (N_6411,N_6082,N_6196);
nor U6412 (N_6412,N_6157,N_6095);
and U6413 (N_6413,N_6038,N_6001);
nand U6414 (N_6414,N_6019,N_6142);
or U6415 (N_6415,N_6138,N_6043);
nand U6416 (N_6416,N_6220,N_6139);
xnor U6417 (N_6417,N_6076,N_6127);
nor U6418 (N_6418,N_6032,N_6000);
xor U6419 (N_6419,N_6025,N_6007);
nor U6420 (N_6420,N_6216,N_6123);
or U6421 (N_6421,N_6216,N_6050);
nor U6422 (N_6422,N_6135,N_6147);
or U6423 (N_6423,N_6052,N_6188);
xor U6424 (N_6424,N_6129,N_6222);
nor U6425 (N_6425,N_6038,N_6009);
and U6426 (N_6426,N_6084,N_6166);
or U6427 (N_6427,N_6221,N_6205);
and U6428 (N_6428,N_6179,N_6219);
and U6429 (N_6429,N_6227,N_6100);
nand U6430 (N_6430,N_6127,N_6141);
nor U6431 (N_6431,N_6130,N_6077);
and U6432 (N_6432,N_6215,N_6012);
nand U6433 (N_6433,N_6063,N_6147);
or U6434 (N_6434,N_6103,N_6087);
or U6435 (N_6435,N_6055,N_6144);
nand U6436 (N_6436,N_6038,N_6114);
xor U6437 (N_6437,N_6047,N_6186);
or U6438 (N_6438,N_6232,N_6181);
and U6439 (N_6439,N_6063,N_6016);
or U6440 (N_6440,N_6158,N_6204);
or U6441 (N_6441,N_6199,N_6185);
xnor U6442 (N_6442,N_6051,N_6016);
xor U6443 (N_6443,N_6180,N_6041);
xnor U6444 (N_6444,N_6020,N_6042);
or U6445 (N_6445,N_6175,N_6174);
or U6446 (N_6446,N_6105,N_6082);
xnor U6447 (N_6447,N_6050,N_6226);
or U6448 (N_6448,N_6180,N_6017);
nor U6449 (N_6449,N_6036,N_6054);
and U6450 (N_6450,N_6237,N_6194);
nor U6451 (N_6451,N_6190,N_6011);
nor U6452 (N_6452,N_6018,N_6164);
or U6453 (N_6453,N_6034,N_6134);
or U6454 (N_6454,N_6028,N_6089);
or U6455 (N_6455,N_6080,N_6043);
xnor U6456 (N_6456,N_6178,N_6110);
or U6457 (N_6457,N_6146,N_6174);
or U6458 (N_6458,N_6149,N_6191);
and U6459 (N_6459,N_6245,N_6108);
xor U6460 (N_6460,N_6095,N_6000);
nor U6461 (N_6461,N_6020,N_6207);
nor U6462 (N_6462,N_6048,N_6007);
and U6463 (N_6463,N_6093,N_6155);
or U6464 (N_6464,N_6113,N_6140);
and U6465 (N_6465,N_6222,N_6219);
xnor U6466 (N_6466,N_6100,N_6169);
nor U6467 (N_6467,N_6191,N_6129);
nor U6468 (N_6468,N_6009,N_6008);
nor U6469 (N_6469,N_6074,N_6045);
and U6470 (N_6470,N_6121,N_6019);
and U6471 (N_6471,N_6196,N_6210);
nand U6472 (N_6472,N_6162,N_6182);
nor U6473 (N_6473,N_6151,N_6157);
or U6474 (N_6474,N_6237,N_6203);
nor U6475 (N_6475,N_6183,N_6085);
and U6476 (N_6476,N_6030,N_6049);
and U6477 (N_6477,N_6087,N_6168);
xor U6478 (N_6478,N_6099,N_6179);
nand U6479 (N_6479,N_6088,N_6041);
xor U6480 (N_6480,N_6079,N_6040);
or U6481 (N_6481,N_6225,N_6001);
or U6482 (N_6482,N_6010,N_6034);
xor U6483 (N_6483,N_6231,N_6172);
xor U6484 (N_6484,N_6230,N_6237);
and U6485 (N_6485,N_6162,N_6065);
xnor U6486 (N_6486,N_6225,N_6142);
nand U6487 (N_6487,N_6143,N_6216);
or U6488 (N_6488,N_6242,N_6028);
nand U6489 (N_6489,N_6026,N_6060);
and U6490 (N_6490,N_6108,N_6199);
and U6491 (N_6491,N_6117,N_6201);
nor U6492 (N_6492,N_6024,N_6220);
nand U6493 (N_6493,N_6106,N_6229);
nor U6494 (N_6494,N_6187,N_6053);
nand U6495 (N_6495,N_6167,N_6099);
and U6496 (N_6496,N_6179,N_6223);
nor U6497 (N_6497,N_6058,N_6193);
or U6498 (N_6498,N_6110,N_6022);
or U6499 (N_6499,N_6229,N_6192);
or U6500 (N_6500,N_6377,N_6338);
xnor U6501 (N_6501,N_6478,N_6407);
nand U6502 (N_6502,N_6266,N_6302);
nand U6503 (N_6503,N_6430,N_6410);
nor U6504 (N_6504,N_6461,N_6265);
xor U6505 (N_6505,N_6402,N_6450);
xnor U6506 (N_6506,N_6281,N_6417);
nand U6507 (N_6507,N_6457,N_6463);
nand U6508 (N_6508,N_6304,N_6484);
and U6509 (N_6509,N_6438,N_6373);
nor U6510 (N_6510,N_6258,N_6378);
nand U6511 (N_6511,N_6260,N_6291);
or U6512 (N_6512,N_6497,N_6372);
or U6513 (N_6513,N_6471,N_6375);
nand U6514 (N_6514,N_6350,N_6413);
and U6515 (N_6515,N_6252,N_6363);
xnor U6516 (N_6516,N_6351,N_6365);
and U6517 (N_6517,N_6434,N_6370);
nor U6518 (N_6518,N_6411,N_6381);
nor U6519 (N_6519,N_6468,N_6397);
nor U6520 (N_6520,N_6421,N_6432);
or U6521 (N_6521,N_6455,N_6286);
nand U6522 (N_6522,N_6420,N_6482);
or U6523 (N_6523,N_6383,N_6283);
xor U6524 (N_6524,N_6349,N_6337);
and U6525 (N_6525,N_6481,N_6262);
and U6526 (N_6526,N_6451,N_6334);
or U6527 (N_6527,N_6414,N_6314);
or U6528 (N_6528,N_6320,N_6400);
and U6529 (N_6529,N_6493,N_6435);
nor U6530 (N_6530,N_6394,N_6441);
nor U6531 (N_6531,N_6296,N_6331);
nor U6532 (N_6532,N_6469,N_6270);
xor U6533 (N_6533,N_6464,N_6251);
xnor U6534 (N_6534,N_6317,N_6426);
nand U6535 (N_6535,N_6292,N_6303);
xnor U6536 (N_6536,N_6366,N_6389);
xnor U6537 (N_6537,N_6295,N_6340);
xor U6538 (N_6538,N_6476,N_6391);
nor U6539 (N_6539,N_6385,N_6440);
and U6540 (N_6540,N_6294,N_6261);
nand U6541 (N_6541,N_6399,N_6355);
xor U6542 (N_6542,N_6442,N_6290);
nor U6543 (N_6543,N_6277,N_6353);
nor U6544 (N_6544,N_6475,N_6382);
or U6545 (N_6545,N_6452,N_6328);
or U6546 (N_6546,N_6395,N_6424);
and U6547 (N_6547,N_6288,N_6390);
or U6548 (N_6548,N_6406,N_6278);
xor U6549 (N_6549,N_6319,N_6496);
nand U6550 (N_6550,N_6490,N_6289);
xor U6551 (N_6551,N_6330,N_6322);
nand U6552 (N_6552,N_6362,N_6250);
and U6553 (N_6553,N_6306,N_6368);
nand U6554 (N_6554,N_6271,N_6364);
nand U6555 (N_6555,N_6479,N_6449);
nor U6556 (N_6556,N_6268,N_6473);
nand U6557 (N_6557,N_6300,N_6285);
and U6558 (N_6558,N_6333,N_6371);
nor U6559 (N_6559,N_6332,N_6398);
nor U6560 (N_6560,N_6428,N_6275);
nand U6561 (N_6561,N_6477,N_6418);
nand U6562 (N_6562,N_6256,N_6324);
and U6563 (N_6563,N_6307,N_6458);
nor U6564 (N_6564,N_6273,N_6339);
nor U6565 (N_6565,N_6485,N_6467);
nor U6566 (N_6566,N_6462,N_6433);
nor U6567 (N_6567,N_6466,N_6269);
xor U6568 (N_6568,N_6409,N_6257);
or U6569 (N_6569,N_6498,N_6264);
or U6570 (N_6570,N_6310,N_6446);
nand U6571 (N_6571,N_6315,N_6499);
xnor U6572 (N_6572,N_6343,N_6408);
or U6573 (N_6573,N_6361,N_6447);
or U6574 (N_6574,N_6436,N_6259);
nor U6575 (N_6575,N_6483,N_6369);
or U6576 (N_6576,N_6313,N_6341);
or U6577 (N_6577,N_6494,N_6492);
and U6578 (N_6578,N_6444,N_6405);
xor U6579 (N_6579,N_6293,N_6380);
nand U6580 (N_6580,N_6419,N_6445);
nand U6581 (N_6581,N_6354,N_6386);
xnor U6582 (N_6582,N_6393,N_6454);
and U6583 (N_6583,N_6352,N_6415);
or U6584 (N_6584,N_6325,N_6376);
and U6585 (N_6585,N_6460,N_6305);
or U6586 (N_6586,N_6412,N_6309);
xor U6587 (N_6587,N_6280,N_6427);
nor U6588 (N_6588,N_6486,N_6308);
nand U6589 (N_6589,N_6274,N_6298);
or U6590 (N_6590,N_6459,N_6416);
nor U6591 (N_6591,N_6299,N_6284);
nand U6592 (N_6592,N_6384,N_6392);
and U6593 (N_6593,N_6318,N_6495);
nand U6594 (N_6594,N_6347,N_6360);
nand U6595 (N_6595,N_6387,N_6344);
nand U6596 (N_6596,N_6253,N_6401);
or U6597 (N_6597,N_6379,N_6316);
nand U6598 (N_6598,N_6488,N_6431);
nor U6599 (N_6599,N_6472,N_6448);
xnor U6600 (N_6600,N_6396,N_6276);
and U6601 (N_6601,N_6388,N_6474);
and U6602 (N_6602,N_6358,N_6359);
nor U6603 (N_6603,N_6348,N_6403);
nand U6604 (N_6604,N_6423,N_6254);
nor U6605 (N_6605,N_6480,N_6312);
or U6606 (N_6606,N_6404,N_6487);
and U6607 (N_6607,N_6453,N_6342);
xor U6608 (N_6608,N_6267,N_6437);
nor U6609 (N_6609,N_6465,N_6272);
nor U6610 (N_6610,N_6323,N_6439);
xnor U6611 (N_6611,N_6336,N_6263);
or U6612 (N_6612,N_6345,N_6470);
nor U6613 (N_6613,N_6326,N_6301);
xor U6614 (N_6614,N_6327,N_6335);
nand U6615 (N_6615,N_6329,N_6311);
nand U6616 (N_6616,N_6346,N_6367);
xnor U6617 (N_6617,N_6422,N_6356);
or U6618 (N_6618,N_6425,N_6255);
nor U6619 (N_6619,N_6456,N_6491);
and U6620 (N_6620,N_6443,N_6374);
and U6621 (N_6621,N_6489,N_6279);
xor U6622 (N_6622,N_6429,N_6321);
nor U6623 (N_6623,N_6287,N_6297);
nor U6624 (N_6624,N_6357,N_6282);
and U6625 (N_6625,N_6484,N_6469);
xnor U6626 (N_6626,N_6457,N_6398);
nand U6627 (N_6627,N_6488,N_6300);
xnor U6628 (N_6628,N_6372,N_6379);
nor U6629 (N_6629,N_6488,N_6250);
xor U6630 (N_6630,N_6430,N_6424);
xnor U6631 (N_6631,N_6467,N_6338);
nor U6632 (N_6632,N_6467,N_6339);
or U6633 (N_6633,N_6302,N_6496);
nand U6634 (N_6634,N_6438,N_6468);
or U6635 (N_6635,N_6408,N_6354);
or U6636 (N_6636,N_6343,N_6353);
and U6637 (N_6637,N_6356,N_6481);
nand U6638 (N_6638,N_6379,N_6478);
nand U6639 (N_6639,N_6470,N_6341);
nand U6640 (N_6640,N_6488,N_6498);
and U6641 (N_6641,N_6492,N_6322);
or U6642 (N_6642,N_6447,N_6413);
or U6643 (N_6643,N_6268,N_6346);
xor U6644 (N_6644,N_6450,N_6473);
nand U6645 (N_6645,N_6435,N_6453);
or U6646 (N_6646,N_6333,N_6459);
nor U6647 (N_6647,N_6277,N_6432);
nand U6648 (N_6648,N_6253,N_6384);
xnor U6649 (N_6649,N_6254,N_6306);
nand U6650 (N_6650,N_6325,N_6455);
nor U6651 (N_6651,N_6358,N_6329);
nor U6652 (N_6652,N_6400,N_6460);
nor U6653 (N_6653,N_6256,N_6326);
xor U6654 (N_6654,N_6250,N_6305);
and U6655 (N_6655,N_6469,N_6324);
xnor U6656 (N_6656,N_6289,N_6487);
or U6657 (N_6657,N_6307,N_6482);
xnor U6658 (N_6658,N_6431,N_6391);
or U6659 (N_6659,N_6261,N_6337);
and U6660 (N_6660,N_6254,N_6413);
nand U6661 (N_6661,N_6319,N_6261);
nand U6662 (N_6662,N_6449,N_6290);
and U6663 (N_6663,N_6252,N_6407);
or U6664 (N_6664,N_6362,N_6308);
and U6665 (N_6665,N_6334,N_6327);
xor U6666 (N_6666,N_6252,N_6306);
and U6667 (N_6667,N_6405,N_6265);
or U6668 (N_6668,N_6318,N_6283);
nand U6669 (N_6669,N_6393,N_6361);
nor U6670 (N_6670,N_6273,N_6326);
and U6671 (N_6671,N_6254,N_6279);
nor U6672 (N_6672,N_6359,N_6250);
nor U6673 (N_6673,N_6448,N_6373);
and U6674 (N_6674,N_6271,N_6283);
xnor U6675 (N_6675,N_6289,N_6410);
and U6676 (N_6676,N_6310,N_6303);
xnor U6677 (N_6677,N_6378,N_6362);
nand U6678 (N_6678,N_6394,N_6299);
nor U6679 (N_6679,N_6354,N_6352);
and U6680 (N_6680,N_6485,N_6394);
nand U6681 (N_6681,N_6322,N_6419);
nand U6682 (N_6682,N_6435,N_6387);
nand U6683 (N_6683,N_6444,N_6322);
or U6684 (N_6684,N_6369,N_6347);
or U6685 (N_6685,N_6310,N_6487);
nor U6686 (N_6686,N_6381,N_6265);
and U6687 (N_6687,N_6336,N_6407);
nor U6688 (N_6688,N_6392,N_6253);
nand U6689 (N_6689,N_6435,N_6339);
and U6690 (N_6690,N_6314,N_6439);
nand U6691 (N_6691,N_6308,N_6316);
nand U6692 (N_6692,N_6392,N_6291);
and U6693 (N_6693,N_6439,N_6356);
nand U6694 (N_6694,N_6391,N_6308);
nor U6695 (N_6695,N_6284,N_6476);
and U6696 (N_6696,N_6422,N_6481);
nor U6697 (N_6697,N_6270,N_6298);
and U6698 (N_6698,N_6340,N_6488);
or U6699 (N_6699,N_6426,N_6394);
and U6700 (N_6700,N_6407,N_6278);
nor U6701 (N_6701,N_6366,N_6272);
or U6702 (N_6702,N_6298,N_6493);
xor U6703 (N_6703,N_6286,N_6374);
nand U6704 (N_6704,N_6271,N_6417);
or U6705 (N_6705,N_6280,N_6491);
nor U6706 (N_6706,N_6484,N_6451);
and U6707 (N_6707,N_6443,N_6332);
nor U6708 (N_6708,N_6358,N_6454);
nand U6709 (N_6709,N_6393,N_6336);
and U6710 (N_6710,N_6448,N_6446);
xor U6711 (N_6711,N_6341,N_6442);
or U6712 (N_6712,N_6434,N_6288);
and U6713 (N_6713,N_6291,N_6400);
and U6714 (N_6714,N_6497,N_6444);
or U6715 (N_6715,N_6336,N_6421);
nand U6716 (N_6716,N_6275,N_6422);
nand U6717 (N_6717,N_6393,N_6451);
nand U6718 (N_6718,N_6298,N_6395);
nand U6719 (N_6719,N_6355,N_6366);
and U6720 (N_6720,N_6253,N_6321);
nand U6721 (N_6721,N_6265,N_6404);
nand U6722 (N_6722,N_6359,N_6472);
and U6723 (N_6723,N_6283,N_6450);
nor U6724 (N_6724,N_6485,N_6325);
nor U6725 (N_6725,N_6417,N_6259);
or U6726 (N_6726,N_6326,N_6395);
xnor U6727 (N_6727,N_6398,N_6477);
nand U6728 (N_6728,N_6395,N_6252);
and U6729 (N_6729,N_6393,N_6392);
or U6730 (N_6730,N_6358,N_6372);
xor U6731 (N_6731,N_6383,N_6456);
and U6732 (N_6732,N_6306,N_6403);
xnor U6733 (N_6733,N_6368,N_6417);
and U6734 (N_6734,N_6320,N_6487);
nand U6735 (N_6735,N_6314,N_6491);
or U6736 (N_6736,N_6346,N_6448);
or U6737 (N_6737,N_6379,N_6345);
and U6738 (N_6738,N_6347,N_6412);
or U6739 (N_6739,N_6379,N_6482);
xnor U6740 (N_6740,N_6496,N_6335);
or U6741 (N_6741,N_6454,N_6349);
nor U6742 (N_6742,N_6284,N_6273);
or U6743 (N_6743,N_6344,N_6300);
nand U6744 (N_6744,N_6348,N_6388);
xnor U6745 (N_6745,N_6313,N_6422);
nand U6746 (N_6746,N_6327,N_6491);
or U6747 (N_6747,N_6488,N_6422);
and U6748 (N_6748,N_6394,N_6481);
nand U6749 (N_6749,N_6301,N_6270);
xor U6750 (N_6750,N_6503,N_6728);
xnor U6751 (N_6751,N_6606,N_6698);
and U6752 (N_6752,N_6710,N_6738);
nor U6753 (N_6753,N_6562,N_6625);
xor U6754 (N_6754,N_6556,N_6702);
or U6755 (N_6755,N_6590,N_6555);
nand U6756 (N_6756,N_6701,N_6723);
nor U6757 (N_6757,N_6641,N_6565);
nor U6758 (N_6758,N_6637,N_6713);
nor U6759 (N_6759,N_6682,N_6697);
and U6760 (N_6760,N_6517,N_6552);
xor U6761 (N_6761,N_6524,N_6621);
nand U6762 (N_6762,N_6733,N_6533);
nand U6763 (N_6763,N_6677,N_6523);
xnor U6764 (N_6764,N_6528,N_6674);
or U6765 (N_6765,N_6699,N_6632);
or U6766 (N_6766,N_6651,N_6539);
nor U6767 (N_6767,N_6530,N_6655);
nor U6768 (N_6768,N_6595,N_6649);
or U6769 (N_6769,N_6605,N_6719);
or U6770 (N_6770,N_6507,N_6737);
and U6771 (N_6771,N_6689,N_6564);
and U6772 (N_6772,N_6624,N_6508);
nand U6773 (N_6773,N_6616,N_6591);
or U6774 (N_6774,N_6665,N_6557);
nor U6775 (N_6775,N_6506,N_6505);
or U6776 (N_6776,N_6521,N_6714);
or U6777 (N_6777,N_6717,N_6549);
xor U6778 (N_6778,N_6726,N_6739);
xnor U6779 (N_6779,N_6500,N_6633);
xor U6780 (N_6780,N_6581,N_6703);
nor U6781 (N_6781,N_6585,N_6575);
or U6782 (N_6782,N_6631,N_6709);
nor U6783 (N_6783,N_6715,N_6529);
nor U6784 (N_6784,N_6598,N_6652);
nor U6785 (N_6785,N_6660,N_6614);
and U6786 (N_6786,N_6670,N_6687);
or U6787 (N_6787,N_6623,N_6573);
nor U6788 (N_6788,N_6619,N_6603);
or U6789 (N_6789,N_6695,N_6700);
and U6790 (N_6790,N_6519,N_6601);
nand U6791 (N_6791,N_6579,N_6622);
nand U6792 (N_6792,N_6536,N_6514);
and U6793 (N_6793,N_6730,N_6712);
xor U6794 (N_6794,N_6648,N_6629);
and U6795 (N_6795,N_6686,N_6742);
and U6796 (N_6796,N_6724,N_6567);
nor U6797 (N_6797,N_6735,N_6743);
nand U6798 (N_6798,N_6675,N_6676);
and U6799 (N_6799,N_6545,N_6662);
nand U6800 (N_6800,N_6571,N_6666);
xnor U6801 (N_6801,N_6515,N_6696);
nor U6802 (N_6802,N_6681,N_6547);
nand U6803 (N_6803,N_6646,N_6620);
nor U6804 (N_6804,N_6647,N_6520);
nor U6805 (N_6805,N_6596,N_6534);
and U6806 (N_6806,N_6580,N_6543);
nor U6807 (N_6807,N_6707,N_6576);
nor U6808 (N_6808,N_6740,N_6650);
xor U6809 (N_6809,N_6643,N_6570);
nor U6810 (N_6810,N_6692,N_6511);
nor U6811 (N_6811,N_6642,N_6691);
or U6812 (N_6812,N_6518,N_6747);
or U6813 (N_6813,N_6532,N_6512);
or U6814 (N_6814,N_6731,N_6634);
nor U6815 (N_6815,N_6716,N_6656);
nand U6816 (N_6816,N_6718,N_6548);
or U6817 (N_6817,N_6609,N_6531);
xnor U6818 (N_6818,N_6626,N_6617);
nand U6819 (N_6819,N_6741,N_6610);
nor U6820 (N_6820,N_6654,N_6586);
nand U6821 (N_6821,N_6568,N_6553);
xnor U6822 (N_6822,N_6736,N_6516);
nor U6823 (N_6823,N_6653,N_6688);
xnor U6824 (N_6824,N_6559,N_6535);
xor U6825 (N_6825,N_6540,N_6663);
xor U6826 (N_6826,N_6563,N_6639);
nand U6827 (N_6827,N_6588,N_6721);
xnor U6828 (N_6828,N_6748,N_6589);
and U6829 (N_6829,N_6658,N_6683);
and U6830 (N_6830,N_6611,N_6618);
nor U6831 (N_6831,N_6704,N_6566);
and U6832 (N_6832,N_6592,N_6636);
or U6833 (N_6833,N_6615,N_6664);
nor U6834 (N_6834,N_6685,N_6745);
xnor U6835 (N_6835,N_6510,N_6706);
xnor U6836 (N_6836,N_6657,N_6720);
xnor U6837 (N_6837,N_6577,N_6569);
or U6838 (N_6838,N_6732,N_6608);
or U6839 (N_6839,N_6599,N_6554);
and U6840 (N_6840,N_6638,N_6630);
nor U6841 (N_6841,N_6509,N_6644);
or U6842 (N_6842,N_6694,N_6705);
nand U6843 (N_6843,N_6561,N_6640);
nand U6844 (N_6844,N_6672,N_6584);
or U6845 (N_6845,N_6541,N_6746);
xor U6846 (N_6846,N_6645,N_6578);
xnor U6847 (N_6847,N_6725,N_6635);
nand U6848 (N_6848,N_6594,N_6607);
xor U6849 (N_6849,N_6708,N_6604);
nand U6850 (N_6850,N_6627,N_6722);
xor U6851 (N_6851,N_6600,N_6659);
and U6852 (N_6852,N_6558,N_6542);
xor U6853 (N_6853,N_6504,N_6693);
and U6854 (N_6854,N_6679,N_6669);
nand U6855 (N_6855,N_6550,N_6628);
xnor U6856 (N_6856,N_6734,N_6572);
nand U6857 (N_6857,N_6537,N_6690);
or U6858 (N_6858,N_6668,N_6661);
nor U6859 (N_6859,N_6671,N_6678);
or U6860 (N_6860,N_6501,N_6583);
and U6861 (N_6861,N_6502,N_6527);
xor U6862 (N_6862,N_6587,N_6582);
nor U6863 (N_6863,N_6538,N_6546);
or U6864 (N_6864,N_6684,N_6612);
xor U6865 (N_6865,N_6593,N_6574);
nor U6866 (N_6866,N_6526,N_6551);
nor U6867 (N_6867,N_6513,N_6544);
xnor U6868 (N_6868,N_6613,N_6744);
nor U6869 (N_6869,N_6711,N_6680);
nand U6870 (N_6870,N_6729,N_6525);
and U6871 (N_6871,N_6522,N_6602);
or U6872 (N_6872,N_6597,N_6560);
xnor U6873 (N_6873,N_6667,N_6673);
nand U6874 (N_6874,N_6727,N_6749);
nor U6875 (N_6875,N_6665,N_6502);
xor U6876 (N_6876,N_6702,N_6697);
or U6877 (N_6877,N_6627,N_6593);
xor U6878 (N_6878,N_6591,N_6650);
nand U6879 (N_6879,N_6619,N_6644);
nand U6880 (N_6880,N_6573,N_6670);
and U6881 (N_6881,N_6725,N_6696);
xnor U6882 (N_6882,N_6621,N_6656);
nor U6883 (N_6883,N_6734,N_6629);
or U6884 (N_6884,N_6692,N_6674);
xor U6885 (N_6885,N_6647,N_6713);
or U6886 (N_6886,N_6508,N_6730);
nor U6887 (N_6887,N_6607,N_6727);
nor U6888 (N_6888,N_6515,N_6672);
or U6889 (N_6889,N_6749,N_6660);
nand U6890 (N_6890,N_6582,N_6599);
and U6891 (N_6891,N_6743,N_6737);
nor U6892 (N_6892,N_6603,N_6731);
nor U6893 (N_6893,N_6519,N_6697);
and U6894 (N_6894,N_6549,N_6553);
nand U6895 (N_6895,N_6588,N_6713);
or U6896 (N_6896,N_6609,N_6575);
nand U6897 (N_6897,N_6610,N_6686);
xor U6898 (N_6898,N_6547,N_6593);
nand U6899 (N_6899,N_6611,N_6664);
xor U6900 (N_6900,N_6730,N_6541);
nand U6901 (N_6901,N_6684,N_6597);
and U6902 (N_6902,N_6595,N_6561);
or U6903 (N_6903,N_6684,N_6655);
nor U6904 (N_6904,N_6660,N_6578);
nand U6905 (N_6905,N_6624,N_6563);
xnor U6906 (N_6906,N_6588,N_6661);
nor U6907 (N_6907,N_6625,N_6536);
nor U6908 (N_6908,N_6735,N_6666);
xor U6909 (N_6909,N_6691,N_6564);
xnor U6910 (N_6910,N_6587,N_6586);
nor U6911 (N_6911,N_6540,N_6720);
nand U6912 (N_6912,N_6635,N_6677);
or U6913 (N_6913,N_6643,N_6739);
or U6914 (N_6914,N_6566,N_6633);
nand U6915 (N_6915,N_6526,N_6501);
and U6916 (N_6916,N_6653,N_6618);
nand U6917 (N_6917,N_6612,N_6545);
nand U6918 (N_6918,N_6670,N_6521);
nor U6919 (N_6919,N_6730,N_6635);
and U6920 (N_6920,N_6654,N_6564);
and U6921 (N_6921,N_6572,N_6739);
nand U6922 (N_6922,N_6737,N_6601);
or U6923 (N_6923,N_6618,N_6734);
xor U6924 (N_6924,N_6660,N_6650);
nor U6925 (N_6925,N_6649,N_6534);
nand U6926 (N_6926,N_6658,N_6556);
nor U6927 (N_6927,N_6540,N_6544);
xnor U6928 (N_6928,N_6741,N_6550);
and U6929 (N_6929,N_6735,N_6637);
or U6930 (N_6930,N_6736,N_6678);
xnor U6931 (N_6931,N_6609,N_6555);
xnor U6932 (N_6932,N_6659,N_6630);
nand U6933 (N_6933,N_6630,N_6735);
nor U6934 (N_6934,N_6520,N_6578);
or U6935 (N_6935,N_6645,N_6648);
nand U6936 (N_6936,N_6612,N_6591);
or U6937 (N_6937,N_6681,N_6517);
nand U6938 (N_6938,N_6748,N_6666);
nor U6939 (N_6939,N_6653,N_6693);
xnor U6940 (N_6940,N_6516,N_6562);
and U6941 (N_6941,N_6709,N_6610);
or U6942 (N_6942,N_6533,N_6556);
xnor U6943 (N_6943,N_6671,N_6522);
xor U6944 (N_6944,N_6534,N_6658);
xnor U6945 (N_6945,N_6644,N_6621);
nor U6946 (N_6946,N_6515,N_6659);
nor U6947 (N_6947,N_6534,N_6682);
and U6948 (N_6948,N_6551,N_6514);
xor U6949 (N_6949,N_6505,N_6747);
nand U6950 (N_6950,N_6628,N_6543);
nand U6951 (N_6951,N_6562,N_6645);
nand U6952 (N_6952,N_6730,N_6535);
nand U6953 (N_6953,N_6653,N_6720);
xor U6954 (N_6954,N_6591,N_6590);
nand U6955 (N_6955,N_6559,N_6695);
xor U6956 (N_6956,N_6637,N_6623);
and U6957 (N_6957,N_6635,N_6690);
nand U6958 (N_6958,N_6617,N_6543);
xor U6959 (N_6959,N_6543,N_6635);
and U6960 (N_6960,N_6529,N_6567);
nand U6961 (N_6961,N_6600,N_6622);
or U6962 (N_6962,N_6557,N_6566);
nand U6963 (N_6963,N_6642,N_6675);
nand U6964 (N_6964,N_6595,N_6593);
or U6965 (N_6965,N_6600,N_6510);
and U6966 (N_6966,N_6670,N_6728);
or U6967 (N_6967,N_6749,N_6530);
xnor U6968 (N_6968,N_6613,N_6677);
xor U6969 (N_6969,N_6540,N_6519);
nand U6970 (N_6970,N_6741,N_6678);
nor U6971 (N_6971,N_6659,N_6665);
nor U6972 (N_6972,N_6748,N_6617);
nor U6973 (N_6973,N_6561,N_6729);
nand U6974 (N_6974,N_6565,N_6553);
nand U6975 (N_6975,N_6577,N_6553);
xnor U6976 (N_6976,N_6583,N_6714);
or U6977 (N_6977,N_6702,N_6526);
xor U6978 (N_6978,N_6677,N_6597);
and U6979 (N_6979,N_6731,N_6722);
or U6980 (N_6980,N_6591,N_6523);
xnor U6981 (N_6981,N_6592,N_6522);
nand U6982 (N_6982,N_6710,N_6575);
nand U6983 (N_6983,N_6588,N_6512);
nand U6984 (N_6984,N_6594,N_6555);
or U6985 (N_6985,N_6595,N_6739);
xor U6986 (N_6986,N_6620,N_6550);
nand U6987 (N_6987,N_6712,N_6682);
or U6988 (N_6988,N_6525,N_6563);
nor U6989 (N_6989,N_6718,N_6653);
xor U6990 (N_6990,N_6681,N_6511);
nand U6991 (N_6991,N_6648,N_6683);
nand U6992 (N_6992,N_6509,N_6636);
or U6993 (N_6993,N_6503,N_6679);
and U6994 (N_6994,N_6611,N_6699);
and U6995 (N_6995,N_6740,N_6546);
and U6996 (N_6996,N_6650,N_6596);
xor U6997 (N_6997,N_6625,N_6635);
nand U6998 (N_6998,N_6708,N_6501);
or U6999 (N_6999,N_6583,N_6612);
nor U7000 (N_7000,N_6820,N_6939);
xnor U7001 (N_7001,N_6918,N_6792);
nand U7002 (N_7002,N_6825,N_6941);
nand U7003 (N_7003,N_6930,N_6983);
nor U7004 (N_7004,N_6947,N_6925);
nor U7005 (N_7005,N_6758,N_6862);
nand U7006 (N_7006,N_6754,N_6986);
or U7007 (N_7007,N_6966,N_6999);
or U7008 (N_7008,N_6830,N_6842);
xnor U7009 (N_7009,N_6819,N_6950);
xnor U7010 (N_7010,N_6837,N_6777);
nor U7011 (N_7011,N_6804,N_6946);
nand U7012 (N_7012,N_6884,N_6880);
nand U7013 (N_7013,N_6912,N_6943);
xnor U7014 (N_7014,N_6993,N_6960);
nor U7015 (N_7015,N_6883,N_6903);
nand U7016 (N_7016,N_6759,N_6970);
xor U7017 (N_7017,N_6803,N_6923);
nand U7018 (N_7018,N_6776,N_6834);
or U7019 (N_7019,N_6957,N_6847);
and U7020 (N_7020,N_6853,N_6784);
or U7021 (N_7021,N_6874,N_6865);
or U7022 (N_7022,N_6887,N_6761);
nand U7023 (N_7023,N_6952,N_6890);
and U7024 (N_7024,N_6882,N_6828);
nand U7025 (N_7025,N_6850,N_6873);
or U7026 (N_7026,N_6821,N_6789);
or U7027 (N_7027,N_6889,N_6813);
and U7028 (N_7028,N_6827,N_6801);
xor U7029 (N_7029,N_6948,N_6785);
nand U7030 (N_7030,N_6894,N_6797);
and U7031 (N_7031,N_6851,N_6756);
xnor U7032 (N_7032,N_6805,N_6843);
nor U7033 (N_7033,N_6823,N_6911);
nand U7034 (N_7034,N_6872,N_6814);
nor U7035 (N_7035,N_6877,N_6794);
xor U7036 (N_7036,N_6871,N_6864);
and U7037 (N_7037,N_6857,N_6974);
nand U7038 (N_7038,N_6962,N_6992);
or U7039 (N_7039,N_6881,N_6854);
xnor U7040 (N_7040,N_6831,N_6969);
nor U7041 (N_7041,N_6787,N_6815);
and U7042 (N_7042,N_6796,N_6888);
or U7043 (N_7043,N_6855,N_6818);
nor U7044 (N_7044,N_6762,N_6798);
and U7045 (N_7045,N_6755,N_6919);
xor U7046 (N_7046,N_6958,N_6771);
or U7047 (N_7047,N_6886,N_6878);
xnor U7048 (N_7048,N_6836,N_6915);
and U7049 (N_7049,N_6858,N_6965);
xnor U7050 (N_7050,N_6994,N_6932);
xor U7051 (N_7051,N_6942,N_6904);
xnor U7052 (N_7052,N_6793,N_6868);
nand U7053 (N_7053,N_6961,N_6775);
nand U7054 (N_7054,N_6891,N_6920);
nor U7055 (N_7055,N_6826,N_6786);
or U7056 (N_7056,N_6964,N_6895);
or U7057 (N_7057,N_6900,N_6806);
or U7058 (N_7058,N_6922,N_6938);
or U7059 (N_7059,N_6859,N_6959);
nand U7060 (N_7060,N_6833,N_6899);
xor U7061 (N_7061,N_6824,N_6972);
nor U7062 (N_7062,N_6778,N_6971);
or U7063 (N_7063,N_6991,N_6980);
and U7064 (N_7064,N_6954,N_6963);
nor U7065 (N_7065,N_6848,N_6779);
and U7066 (N_7066,N_6870,N_6844);
nor U7067 (N_7067,N_6816,N_6782);
and U7068 (N_7068,N_6808,N_6998);
nor U7069 (N_7069,N_6879,N_6913);
nand U7070 (N_7070,N_6973,N_6812);
xnor U7071 (N_7071,N_6800,N_6982);
nor U7072 (N_7072,N_6846,N_6917);
xor U7073 (N_7073,N_6910,N_6981);
and U7074 (N_7074,N_6997,N_6901);
and U7075 (N_7075,N_6835,N_6769);
and U7076 (N_7076,N_6945,N_6940);
xnor U7077 (N_7077,N_6929,N_6856);
nor U7078 (N_7078,N_6921,N_6896);
and U7079 (N_7079,N_6907,N_6953);
nand U7080 (N_7080,N_6924,N_6867);
and U7081 (N_7081,N_6984,N_6951);
xor U7082 (N_7082,N_6838,N_6841);
and U7083 (N_7083,N_6928,N_6773);
nand U7084 (N_7084,N_6995,N_6750);
and U7085 (N_7085,N_6916,N_6892);
and U7086 (N_7086,N_6977,N_6934);
xnor U7087 (N_7087,N_6944,N_6955);
or U7088 (N_7088,N_6988,N_6845);
nand U7089 (N_7089,N_6968,N_6768);
or U7090 (N_7090,N_6897,N_6757);
nand U7091 (N_7091,N_6764,N_6839);
nand U7092 (N_7092,N_6875,N_6906);
nand U7093 (N_7093,N_6937,N_6849);
nand U7094 (N_7094,N_6752,N_6876);
nor U7095 (N_7095,N_6765,N_6790);
and U7096 (N_7096,N_6753,N_6898);
or U7097 (N_7097,N_6772,N_6926);
nand U7098 (N_7098,N_6908,N_6817);
or U7099 (N_7099,N_6767,N_6989);
nor U7100 (N_7100,N_6780,N_6807);
nor U7101 (N_7101,N_6949,N_6976);
nor U7102 (N_7102,N_6852,N_6795);
and U7103 (N_7103,N_6933,N_6996);
and U7104 (N_7104,N_6979,N_6809);
and U7105 (N_7105,N_6902,N_6770);
xor U7106 (N_7106,N_6791,N_6935);
nor U7107 (N_7107,N_6802,N_6967);
and U7108 (N_7108,N_6810,N_6840);
xor U7109 (N_7109,N_6760,N_6766);
and U7110 (N_7110,N_6863,N_6799);
xnor U7111 (N_7111,N_6931,N_6861);
nor U7112 (N_7112,N_6832,N_6781);
xnor U7113 (N_7113,N_6860,N_6990);
and U7114 (N_7114,N_6751,N_6829);
nand U7115 (N_7115,N_6987,N_6893);
and U7116 (N_7116,N_6869,N_6788);
xor U7117 (N_7117,N_6885,N_6783);
and U7118 (N_7118,N_6975,N_6866);
nand U7119 (N_7119,N_6763,N_6822);
nor U7120 (N_7120,N_6985,N_6936);
or U7121 (N_7121,N_6905,N_6909);
or U7122 (N_7122,N_6811,N_6914);
or U7123 (N_7123,N_6956,N_6774);
and U7124 (N_7124,N_6927,N_6978);
or U7125 (N_7125,N_6953,N_6945);
nor U7126 (N_7126,N_6840,N_6750);
nand U7127 (N_7127,N_6980,N_6917);
nand U7128 (N_7128,N_6895,N_6974);
and U7129 (N_7129,N_6805,N_6755);
nor U7130 (N_7130,N_6855,N_6901);
xnor U7131 (N_7131,N_6792,N_6875);
xor U7132 (N_7132,N_6909,N_6973);
xor U7133 (N_7133,N_6964,N_6899);
and U7134 (N_7134,N_6985,N_6793);
xor U7135 (N_7135,N_6981,N_6899);
and U7136 (N_7136,N_6898,N_6915);
and U7137 (N_7137,N_6914,N_6822);
nor U7138 (N_7138,N_6987,N_6969);
or U7139 (N_7139,N_6750,N_6939);
and U7140 (N_7140,N_6823,N_6785);
nand U7141 (N_7141,N_6968,N_6866);
xnor U7142 (N_7142,N_6970,N_6843);
or U7143 (N_7143,N_6811,N_6880);
nor U7144 (N_7144,N_6833,N_6966);
nor U7145 (N_7145,N_6839,N_6900);
xnor U7146 (N_7146,N_6798,N_6896);
nand U7147 (N_7147,N_6882,N_6835);
or U7148 (N_7148,N_6776,N_6932);
or U7149 (N_7149,N_6811,N_6778);
and U7150 (N_7150,N_6930,N_6797);
or U7151 (N_7151,N_6936,N_6975);
or U7152 (N_7152,N_6968,N_6973);
and U7153 (N_7153,N_6851,N_6980);
xnor U7154 (N_7154,N_6988,N_6960);
nor U7155 (N_7155,N_6877,N_6974);
nor U7156 (N_7156,N_6916,N_6816);
nand U7157 (N_7157,N_6962,N_6996);
and U7158 (N_7158,N_6887,N_6831);
and U7159 (N_7159,N_6762,N_6917);
and U7160 (N_7160,N_6913,N_6865);
and U7161 (N_7161,N_6757,N_6934);
and U7162 (N_7162,N_6950,N_6796);
nand U7163 (N_7163,N_6811,N_6910);
nor U7164 (N_7164,N_6992,N_6955);
nand U7165 (N_7165,N_6955,N_6993);
xor U7166 (N_7166,N_6754,N_6834);
xor U7167 (N_7167,N_6898,N_6894);
xnor U7168 (N_7168,N_6912,N_6930);
nor U7169 (N_7169,N_6881,N_6985);
nand U7170 (N_7170,N_6881,N_6981);
or U7171 (N_7171,N_6825,N_6753);
nand U7172 (N_7172,N_6900,N_6788);
nor U7173 (N_7173,N_6768,N_6822);
xor U7174 (N_7174,N_6995,N_6794);
nand U7175 (N_7175,N_6945,N_6763);
nor U7176 (N_7176,N_6847,N_6927);
xnor U7177 (N_7177,N_6928,N_6878);
or U7178 (N_7178,N_6992,N_6917);
nor U7179 (N_7179,N_6868,N_6906);
xor U7180 (N_7180,N_6996,N_6894);
nor U7181 (N_7181,N_6857,N_6959);
or U7182 (N_7182,N_6835,N_6980);
and U7183 (N_7183,N_6968,N_6996);
or U7184 (N_7184,N_6973,N_6959);
or U7185 (N_7185,N_6878,N_6856);
nor U7186 (N_7186,N_6939,N_6763);
xnor U7187 (N_7187,N_6873,N_6753);
nor U7188 (N_7188,N_6993,N_6852);
nor U7189 (N_7189,N_6876,N_6970);
xnor U7190 (N_7190,N_6782,N_6844);
nand U7191 (N_7191,N_6963,N_6848);
or U7192 (N_7192,N_6780,N_6826);
xnor U7193 (N_7193,N_6808,N_6927);
and U7194 (N_7194,N_6859,N_6917);
nor U7195 (N_7195,N_6919,N_6962);
or U7196 (N_7196,N_6875,N_6899);
nor U7197 (N_7197,N_6753,N_6869);
nor U7198 (N_7198,N_6791,N_6918);
xnor U7199 (N_7199,N_6980,N_6815);
nand U7200 (N_7200,N_6993,N_6933);
or U7201 (N_7201,N_6929,N_6795);
or U7202 (N_7202,N_6892,N_6757);
or U7203 (N_7203,N_6818,N_6899);
nor U7204 (N_7204,N_6778,N_6903);
or U7205 (N_7205,N_6808,N_6987);
nand U7206 (N_7206,N_6948,N_6819);
nor U7207 (N_7207,N_6943,N_6882);
nor U7208 (N_7208,N_6766,N_6790);
nand U7209 (N_7209,N_6975,N_6766);
or U7210 (N_7210,N_6774,N_6813);
xor U7211 (N_7211,N_6895,N_6912);
and U7212 (N_7212,N_6835,N_6958);
or U7213 (N_7213,N_6987,N_6783);
or U7214 (N_7214,N_6780,N_6754);
nand U7215 (N_7215,N_6872,N_6910);
nand U7216 (N_7216,N_6889,N_6753);
xnor U7217 (N_7217,N_6848,N_6874);
xnor U7218 (N_7218,N_6994,N_6930);
or U7219 (N_7219,N_6822,N_6868);
nand U7220 (N_7220,N_6840,N_6757);
xnor U7221 (N_7221,N_6757,N_6810);
xnor U7222 (N_7222,N_6828,N_6830);
nor U7223 (N_7223,N_6803,N_6857);
xor U7224 (N_7224,N_6796,N_6869);
and U7225 (N_7225,N_6788,N_6805);
or U7226 (N_7226,N_6988,N_6856);
and U7227 (N_7227,N_6890,N_6857);
nand U7228 (N_7228,N_6879,N_6996);
nor U7229 (N_7229,N_6811,N_6755);
nand U7230 (N_7230,N_6776,N_6849);
xnor U7231 (N_7231,N_6812,N_6946);
xor U7232 (N_7232,N_6936,N_6849);
xnor U7233 (N_7233,N_6773,N_6809);
nand U7234 (N_7234,N_6884,N_6924);
or U7235 (N_7235,N_6920,N_6814);
nand U7236 (N_7236,N_6831,N_6886);
and U7237 (N_7237,N_6984,N_6845);
or U7238 (N_7238,N_6769,N_6973);
and U7239 (N_7239,N_6766,N_6917);
xor U7240 (N_7240,N_6891,N_6873);
xnor U7241 (N_7241,N_6933,N_6787);
nor U7242 (N_7242,N_6758,N_6796);
or U7243 (N_7243,N_6951,N_6831);
xor U7244 (N_7244,N_6870,N_6891);
nor U7245 (N_7245,N_6950,N_6771);
and U7246 (N_7246,N_6943,N_6951);
nor U7247 (N_7247,N_6905,N_6982);
xor U7248 (N_7248,N_6794,N_6930);
or U7249 (N_7249,N_6756,N_6838);
xnor U7250 (N_7250,N_7188,N_7221);
xor U7251 (N_7251,N_7134,N_7168);
and U7252 (N_7252,N_7101,N_7147);
or U7253 (N_7253,N_7138,N_7214);
nor U7254 (N_7254,N_7031,N_7226);
nand U7255 (N_7255,N_7099,N_7186);
nor U7256 (N_7256,N_7011,N_7128);
or U7257 (N_7257,N_7081,N_7193);
or U7258 (N_7258,N_7204,N_7001);
or U7259 (N_7259,N_7088,N_7240);
nor U7260 (N_7260,N_7005,N_7068);
and U7261 (N_7261,N_7104,N_7019);
or U7262 (N_7262,N_7034,N_7073);
nor U7263 (N_7263,N_7030,N_7151);
xnor U7264 (N_7264,N_7094,N_7141);
or U7265 (N_7265,N_7035,N_7085);
xor U7266 (N_7266,N_7126,N_7009);
and U7267 (N_7267,N_7122,N_7242);
and U7268 (N_7268,N_7023,N_7146);
nor U7269 (N_7269,N_7061,N_7022);
nor U7270 (N_7270,N_7143,N_7201);
nor U7271 (N_7271,N_7060,N_7096);
nor U7272 (N_7272,N_7131,N_7194);
nand U7273 (N_7273,N_7248,N_7236);
xor U7274 (N_7274,N_7004,N_7223);
nand U7275 (N_7275,N_7243,N_7070);
nor U7276 (N_7276,N_7229,N_7054);
or U7277 (N_7277,N_7212,N_7015);
nor U7278 (N_7278,N_7117,N_7189);
nand U7279 (N_7279,N_7167,N_7093);
and U7280 (N_7280,N_7207,N_7056);
nand U7281 (N_7281,N_7179,N_7007);
and U7282 (N_7282,N_7231,N_7109);
and U7283 (N_7283,N_7067,N_7198);
or U7284 (N_7284,N_7121,N_7043);
nor U7285 (N_7285,N_7006,N_7050);
and U7286 (N_7286,N_7148,N_7245);
or U7287 (N_7287,N_7244,N_7100);
nor U7288 (N_7288,N_7082,N_7132);
or U7289 (N_7289,N_7124,N_7063);
or U7290 (N_7290,N_7069,N_7213);
and U7291 (N_7291,N_7125,N_7097);
nand U7292 (N_7292,N_7028,N_7202);
xor U7293 (N_7293,N_7098,N_7080);
and U7294 (N_7294,N_7018,N_7105);
and U7295 (N_7295,N_7185,N_7029);
xor U7296 (N_7296,N_7205,N_7027);
xnor U7297 (N_7297,N_7181,N_7234);
xnor U7298 (N_7298,N_7110,N_7053);
nor U7299 (N_7299,N_7012,N_7076);
nor U7300 (N_7300,N_7045,N_7040);
nand U7301 (N_7301,N_7103,N_7108);
or U7302 (N_7302,N_7052,N_7142);
and U7303 (N_7303,N_7048,N_7075);
and U7304 (N_7304,N_7078,N_7164);
nor U7305 (N_7305,N_7171,N_7017);
nand U7306 (N_7306,N_7196,N_7175);
and U7307 (N_7307,N_7120,N_7086);
or U7308 (N_7308,N_7135,N_7008);
nor U7309 (N_7309,N_7062,N_7046);
or U7310 (N_7310,N_7089,N_7241);
nand U7311 (N_7311,N_7140,N_7118);
xnor U7312 (N_7312,N_7169,N_7042);
nor U7313 (N_7313,N_7037,N_7187);
and U7314 (N_7314,N_7021,N_7219);
xnor U7315 (N_7315,N_7064,N_7172);
or U7316 (N_7316,N_7049,N_7173);
or U7317 (N_7317,N_7183,N_7091);
xor U7318 (N_7318,N_7247,N_7136);
or U7319 (N_7319,N_7084,N_7210);
nor U7320 (N_7320,N_7209,N_7158);
and U7321 (N_7321,N_7227,N_7002);
xnor U7322 (N_7322,N_7051,N_7041);
nor U7323 (N_7323,N_7190,N_7203);
and U7324 (N_7324,N_7153,N_7127);
xnor U7325 (N_7325,N_7166,N_7032);
nand U7326 (N_7326,N_7152,N_7176);
and U7327 (N_7327,N_7154,N_7195);
xor U7328 (N_7328,N_7092,N_7079);
xor U7329 (N_7329,N_7129,N_7003);
nand U7330 (N_7330,N_7178,N_7139);
and U7331 (N_7331,N_7216,N_7016);
nand U7332 (N_7332,N_7233,N_7137);
nand U7333 (N_7333,N_7239,N_7013);
or U7334 (N_7334,N_7112,N_7115);
and U7335 (N_7335,N_7159,N_7000);
nor U7336 (N_7336,N_7058,N_7083);
or U7337 (N_7337,N_7206,N_7033);
nand U7338 (N_7338,N_7218,N_7200);
xnor U7339 (N_7339,N_7072,N_7235);
or U7340 (N_7340,N_7165,N_7025);
nand U7341 (N_7341,N_7228,N_7220);
or U7342 (N_7342,N_7149,N_7111);
xor U7343 (N_7343,N_7133,N_7066);
xor U7344 (N_7344,N_7059,N_7215);
and U7345 (N_7345,N_7238,N_7157);
nor U7346 (N_7346,N_7163,N_7071);
xor U7347 (N_7347,N_7182,N_7177);
nand U7348 (N_7348,N_7222,N_7156);
or U7349 (N_7349,N_7020,N_7047);
xnor U7350 (N_7350,N_7160,N_7184);
nor U7351 (N_7351,N_7044,N_7225);
xnor U7352 (N_7352,N_7217,N_7024);
or U7353 (N_7353,N_7211,N_7161);
xor U7354 (N_7354,N_7174,N_7114);
or U7355 (N_7355,N_7123,N_7116);
nand U7356 (N_7356,N_7026,N_7246);
nor U7357 (N_7357,N_7145,N_7119);
xnor U7358 (N_7358,N_7144,N_7150);
xnor U7359 (N_7359,N_7230,N_7102);
nor U7360 (N_7360,N_7074,N_7192);
nor U7361 (N_7361,N_7010,N_7162);
xor U7362 (N_7362,N_7224,N_7057);
and U7363 (N_7363,N_7090,N_7087);
and U7364 (N_7364,N_7170,N_7077);
nor U7365 (N_7365,N_7014,N_7106);
or U7366 (N_7366,N_7036,N_7197);
or U7367 (N_7367,N_7055,N_7232);
or U7368 (N_7368,N_7208,N_7237);
nand U7369 (N_7369,N_7095,N_7180);
or U7370 (N_7370,N_7065,N_7130);
xor U7371 (N_7371,N_7107,N_7155);
and U7372 (N_7372,N_7113,N_7039);
nand U7373 (N_7373,N_7191,N_7249);
and U7374 (N_7374,N_7038,N_7199);
and U7375 (N_7375,N_7158,N_7130);
xnor U7376 (N_7376,N_7193,N_7226);
and U7377 (N_7377,N_7092,N_7084);
nor U7378 (N_7378,N_7098,N_7249);
or U7379 (N_7379,N_7084,N_7115);
nor U7380 (N_7380,N_7130,N_7017);
and U7381 (N_7381,N_7106,N_7221);
nor U7382 (N_7382,N_7120,N_7142);
nand U7383 (N_7383,N_7081,N_7131);
xnor U7384 (N_7384,N_7136,N_7048);
or U7385 (N_7385,N_7066,N_7065);
or U7386 (N_7386,N_7100,N_7010);
and U7387 (N_7387,N_7025,N_7022);
or U7388 (N_7388,N_7204,N_7163);
and U7389 (N_7389,N_7042,N_7178);
and U7390 (N_7390,N_7067,N_7069);
or U7391 (N_7391,N_7011,N_7191);
xor U7392 (N_7392,N_7174,N_7056);
or U7393 (N_7393,N_7022,N_7134);
nor U7394 (N_7394,N_7123,N_7163);
or U7395 (N_7395,N_7171,N_7172);
and U7396 (N_7396,N_7033,N_7236);
or U7397 (N_7397,N_7043,N_7204);
and U7398 (N_7398,N_7191,N_7145);
xor U7399 (N_7399,N_7138,N_7190);
xor U7400 (N_7400,N_7137,N_7101);
or U7401 (N_7401,N_7006,N_7095);
xnor U7402 (N_7402,N_7087,N_7070);
xnor U7403 (N_7403,N_7084,N_7048);
or U7404 (N_7404,N_7034,N_7193);
and U7405 (N_7405,N_7239,N_7008);
nor U7406 (N_7406,N_7159,N_7238);
xnor U7407 (N_7407,N_7234,N_7140);
or U7408 (N_7408,N_7190,N_7015);
xnor U7409 (N_7409,N_7232,N_7196);
or U7410 (N_7410,N_7236,N_7193);
xor U7411 (N_7411,N_7188,N_7151);
or U7412 (N_7412,N_7015,N_7163);
and U7413 (N_7413,N_7227,N_7025);
nand U7414 (N_7414,N_7245,N_7174);
nor U7415 (N_7415,N_7189,N_7235);
and U7416 (N_7416,N_7106,N_7122);
nand U7417 (N_7417,N_7236,N_7006);
nand U7418 (N_7418,N_7185,N_7132);
nand U7419 (N_7419,N_7045,N_7099);
nand U7420 (N_7420,N_7098,N_7195);
and U7421 (N_7421,N_7119,N_7008);
and U7422 (N_7422,N_7228,N_7197);
nor U7423 (N_7423,N_7048,N_7013);
nand U7424 (N_7424,N_7206,N_7241);
nor U7425 (N_7425,N_7182,N_7118);
nor U7426 (N_7426,N_7007,N_7200);
and U7427 (N_7427,N_7203,N_7111);
nor U7428 (N_7428,N_7245,N_7080);
nor U7429 (N_7429,N_7124,N_7108);
or U7430 (N_7430,N_7032,N_7048);
and U7431 (N_7431,N_7248,N_7249);
nor U7432 (N_7432,N_7011,N_7189);
xor U7433 (N_7433,N_7216,N_7163);
and U7434 (N_7434,N_7052,N_7121);
and U7435 (N_7435,N_7221,N_7048);
and U7436 (N_7436,N_7104,N_7020);
nor U7437 (N_7437,N_7112,N_7023);
and U7438 (N_7438,N_7030,N_7172);
nor U7439 (N_7439,N_7040,N_7097);
nand U7440 (N_7440,N_7058,N_7178);
nor U7441 (N_7441,N_7230,N_7023);
xor U7442 (N_7442,N_7041,N_7137);
xnor U7443 (N_7443,N_7050,N_7014);
nor U7444 (N_7444,N_7047,N_7083);
xor U7445 (N_7445,N_7200,N_7044);
nand U7446 (N_7446,N_7074,N_7187);
or U7447 (N_7447,N_7181,N_7143);
nand U7448 (N_7448,N_7114,N_7201);
or U7449 (N_7449,N_7136,N_7000);
nand U7450 (N_7450,N_7160,N_7139);
or U7451 (N_7451,N_7158,N_7120);
and U7452 (N_7452,N_7068,N_7088);
or U7453 (N_7453,N_7229,N_7163);
nand U7454 (N_7454,N_7190,N_7213);
xnor U7455 (N_7455,N_7096,N_7190);
nand U7456 (N_7456,N_7093,N_7013);
and U7457 (N_7457,N_7071,N_7179);
xor U7458 (N_7458,N_7036,N_7051);
or U7459 (N_7459,N_7162,N_7042);
xor U7460 (N_7460,N_7101,N_7232);
nand U7461 (N_7461,N_7017,N_7221);
and U7462 (N_7462,N_7093,N_7230);
xnor U7463 (N_7463,N_7037,N_7097);
xnor U7464 (N_7464,N_7133,N_7222);
xnor U7465 (N_7465,N_7162,N_7080);
nor U7466 (N_7466,N_7004,N_7207);
or U7467 (N_7467,N_7081,N_7102);
nor U7468 (N_7468,N_7247,N_7193);
xnor U7469 (N_7469,N_7229,N_7198);
or U7470 (N_7470,N_7047,N_7194);
xor U7471 (N_7471,N_7146,N_7061);
or U7472 (N_7472,N_7144,N_7057);
xor U7473 (N_7473,N_7238,N_7219);
or U7474 (N_7474,N_7166,N_7094);
and U7475 (N_7475,N_7081,N_7187);
nor U7476 (N_7476,N_7018,N_7029);
nor U7477 (N_7477,N_7037,N_7157);
xnor U7478 (N_7478,N_7225,N_7058);
xnor U7479 (N_7479,N_7244,N_7081);
xnor U7480 (N_7480,N_7057,N_7246);
and U7481 (N_7481,N_7100,N_7063);
nor U7482 (N_7482,N_7119,N_7005);
or U7483 (N_7483,N_7245,N_7134);
nand U7484 (N_7484,N_7069,N_7161);
or U7485 (N_7485,N_7009,N_7246);
xor U7486 (N_7486,N_7081,N_7113);
xnor U7487 (N_7487,N_7083,N_7076);
xor U7488 (N_7488,N_7160,N_7170);
xnor U7489 (N_7489,N_7073,N_7208);
nor U7490 (N_7490,N_7115,N_7067);
nand U7491 (N_7491,N_7203,N_7033);
or U7492 (N_7492,N_7017,N_7164);
or U7493 (N_7493,N_7056,N_7012);
nor U7494 (N_7494,N_7139,N_7206);
nor U7495 (N_7495,N_7013,N_7143);
and U7496 (N_7496,N_7152,N_7087);
nor U7497 (N_7497,N_7039,N_7073);
xor U7498 (N_7498,N_7188,N_7035);
and U7499 (N_7499,N_7185,N_7085);
nand U7500 (N_7500,N_7457,N_7402);
nand U7501 (N_7501,N_7333,N_7290);
nand U7502 (N_7502,N_7267,N_7453);
and U7503 (N_7503,N_7259,N_7260);
xor U7504 (N_7504,N_7489,N_7344);
nand U7505 (N_7505,N_7346,N_7297);
and U7506 (N_7506,N_7268,N_7450);
nand U7507 (N_7507,N_7264,N_7354);
or U7508 (N_7508,N_7287,N_7488);
or U7509 (N_7509,N_7274,N_7451);
or U7510 (N_7510,N_7419,N_7433);
nor U7511 (N_7511,N_7360,N_7376);
or U7512 (N_7512,N_7455,N_7498);
nand U7513 (N_7513,N_7304,N_7439);
nand U7514 (N_7514,N_7397,N_7461);
or U7515 (N_7515,N_7383,N_7330);
xor U7516 (N_7516,N_7472,N_7255);
nand U7517 (N_7517,N_7432,N_7481);
or U7518 (N_7518,N_7312,N_7411);
nand U7519 (N_7519,N_7286,N_7308);
xnor U7520 (N_7520,N_7302,N_7283);
and U7521 (N_7521,N_7306,N_7284);
and U7522 (N_7522,N_7467,N_7493);
and U7523 (N_7523,N_7313,N_7321);
nor U7524 (N_7524,N_7323,N_7315);
or U7525 (N_7525,N_7320,N_7416);
nand U7526 (N_7526,N_7431,N_7311);
nor U7527 (N_7527,N_7483,N_7337);
and U7528 (N_7528,N_7299,N_7292);
and U7529 (N_7529,N_7462,N_7331);
nor U7530 (N_7530,N_7422,N_7296);
xor U7531 (N_7531,N_7480,N_7407);
nand U7532 (N_7532,N_7420,N_7396);
nor U7533 (N_7533,N_7497,N_7293);
xor U7534 (N_7534,N_7368,N_7252);
xnor U7535 (N_7535,N_7487,N_7348);
xnor U7536 (N_7536,N_7482,N_7262);
xor U7537 (N_7537,N_7265,N_7380);
xor U7538 (N_7538,N_7278,N_7374);
xnor U7539 (N_7539,N_7266,N_7400);
nand U7540 (N_7540,N_7458,N_7336);
nor U7541 (N_7541,N_7391,N_7414);
nand U7542 (N_7542,N_7327,N_7285);
and U7543 (N_7543,N_7486,N_7310);
xnor U7544 (N_7544,N_7393,N_7349);
xor U7545 (N_7545,N_7452,N_7258);
and U7546 (N_7546,N_7355,N_7466);
and U7547 (N_7547,N_7359,N_7317);
or U7548 (N_7548,N_7473,N_7273);
nor U7549 (N_7549,N_7443,N_7417);
and U7550 (N_7550,N_7386,N_7390);
and U7551 (N_7551,N_7424,N_7324);
and U7552 (N_7552,N_7362,N_7447);
nand U7553 (N_7553,N_7499,N_7387);
nor U7554 (N_7554,N_7428,N_7491);
xor U7555 (N_7555,N_7418,N_7394);
and U7556 (N_7556,N_7479,N_7470);
xnor U7557 (N_7557,N_7289,N_7395);
nor U7558 (N_7558,N_7485,N_7305);
nand U7559 (N_7559,N_7250,N_7465);
nand U7560 (N_7560,N_7280,N_7369);
xor U7561 (N_7561,N_7254,N_7353);
nand U7562 (N_7562,N_7270,N_7322);
and U7563 (N_7563,N_7375,N_7401);
nand U7564 (N_7564,N_7282,N_7410);
nor U7565 (N_7565,N_7316,N_7358);
and U7566 (N_7566,N_7378,N_7406);
and U7567 (N_7567,N_7345,N_7365);
nand U7568 (N_7568,N_7340,N_7468);
xnor U7569 (N_7569,N_7343,N_7440);
and U7570 (N_7570,N_7277,N_7469);
nand U7571 (N_7571,N_7446,N_7478);
or U7572 (N_7572,N_7399,N_7405);
and U7573 (N_7573,N_7474,N_7471);
xnor U7574 (N_7574,N_7435,N_7415);
and U7575 (N_7575,N_7373,N_7445);
nor U7576 (N_7576,N_7367,N_7256);
or U7577 (N_7577,N_7263,N_7303);
xor U7578 (N_7578,N_7456,N_7425);
or U7579 (N_7579,N_7364,N_7409);
nor U7580 (N_7580,N_7495,N_7436);
xor U7581 (N_7581,N_7492,N_7384);
xnor U7582 (N_7582,N_7326,N_7427);
nor U7583 (N_7583,N_7379,N_7261);
xor U7584 (N_7584,N_7423,N_7475);
and U7585 (N_7585,N_7490,N_7253);
xnor U7586 (N_7586,N_7463,N_7314);
or U7587 (N_7587,N_7476,N_7421);
and U7588 (N_7588,N_7385,N_7309);
nor U7589 (N_7589,N_7269,N_7350);
nand U7590 (N_7590,N_7442,N_7412);
or U7591 (N_7591,N_7363,N_7298);
xnor U7592 (N_7592,N_7430,N_7372);
nand U7593 (N_7593,N_7477,N_7413);
and U7594 (N_7594,N_7257,N_7325);
or U7595 (N_7595,N_7398,N_7295);
xnor U7596 (N_7596,N_7338,N_7279);
and U7597 (N_7597,N_7335,N_7341);
xnor U7598 (N_7598,N_7454,N_7272);
xnor U7599 (N_7599,N_7356,N_7449);
nor U7600 (N_7600,N_7370,N_7448);
xnor U7601 (N_7601,N_7464,N_7300);
xnor U7602 (N_7602,N_7351,N_7484);
nand U7603 (N_7603,N_7328,N_7392);
nand U7604 (N_7604,N_7307,N_7352);
or U7605 (N_7605,N_7294,N_7377);
xor U7606 (N_7606,N_7319,N_7403);
and U7607 (N_7607,N_7494,N_7438);
xnor U7608 (N_7608,N_7301,N_7444);
or U7609 (N_7609,N_7347,N_7426);
nor U7610 (N_7610,N_7366,N_7332);
or U7611 (N_7611,N_7388,N_7389);
nand U7612 (N_7612,N_7459,N_7329);
and U7613 (N_7613,N_7276,N_7318);
nor U7614 (N_7614,N_7361,N_7357);
and U7615 (N_7615,N_7371,N_7251);
xor U7616 (N_7616,N_7441,N_7408);
nor U7617 (N_7617,N_7381,N_7281);
or U7618 (N_7618,N_7334,N_7342);
and U7619 (N_7619,N_7382,N_7437);
nor U7620 (N_7620,N_7496,N_7404);
nand U7621 (N_7621,N_7339,N_7429);
nor U7622 (N_7622,N_7460,N_7291);
or U7623 (N_7623,N_7434,N_7275);
xor U7624 (N_7624,N_7288,N_7271);
or U7625 (N_7625,N_7293,N_7456);
or U7626 (N_7626,N_7408,N_7473);
xor U7627 (N_7627,N_7370,N_7421);
or U7628 (N_7628,N_7413,N_7340);
and U7629 (N_7629,N_7403,N_7387);
and U7630 (N_7630,N_7416,N_7358);
nand U7631 (N_7631,N_7292,N_7439);
or U7632 (N_7632,N_7258,N_7422);
and U7633 (N_7633,N_7369,N_7415);
nor U7634 (N_7634,N_7288,N_7448);
nand U7635 (N_7635,N_7355,N_7331);
xnor U7636 (N_7636,N_7437,N_7465);
xnor U7637 (N_7637,N_7338,N_7281);
and U7638 (N_7638,N_7264,N_7380);
and U7639 (N_7639,N_7491,N_7356);
xnor U7640 (N_7640,N_7403,N_7368);
xnor U7641 (N_7641,N_7327,N_7314);
nor U7642 (N_7642,N_7282,N_7358);
xnor U7643 (N_7643,N_7326,N_7301);
nor U7644 (N_7644,N_7411,N_7283);
and U7645 (N_7645,N_7338,N_7358);
nor U7646 (N_7646,N_7390,N_7470);
nor U7647 (N_7647,N_7324,N_7395);
nand U7648 (N_7648,N_7306,N_7436);
nand U7649 (N_7649,N_7296,N_7443);
and U7650 (N_7650,N_7418,N_7440);
xor U7651 (N_7651,N_7445,N_7388);
nand U7652 (N_7652,N_7489,N_7335);
nor U7653 (N_7653,N_7412,N_7353);
nand U7654 (N_7654,N_7378,N_7295);
nor U7655 (N_7655,N_7291,N_7479);
xor U7656 (N_7656,N_7328,N_7288);
and U7657 (N_7657,N_7382,N_7317);
nand U7658 (N_7658,N_7312,N_7449);
or U7659 (N_7659,N_7420,N_7251);
nand U7660 (N_7660,N_7372,N_7456);
or U7661 (N_7661,N_7287,N_7361);
and U7662 (N_7662,N_7461,N_7465);
xnor U7663 (N_7663,N_7479,N_7471);
or U7664 (N_7664,N_7414,N_7257);
or U7665 (N_7665,N_7490,N_7457);
nand U7666 (N_7666,N_7305,N_7371);
nand U7667 (N_7667,N_7422,N_7484);
nand U7668 (N_7668,N_7270,N_7404);
and U7669 (N_7669,N_7305,N_7250);
or U7670 (N_7670,N_7425,N_7359);
nand U7671 (N_7671,N_7489,N_7414);
and U7672 (N_7672,N_7379,N_7284);
nor U7673 (N_7673,N_7475,N_7305);
and U7674 (N_7674,N_7267,N_7326);
nor U7675 (N_7675,N_7313,N_7359);
or U7676 (N_7676,N_7416,N_7306);
nand U7677 (N_7677,N_7308,N_7293);
nand U7678 (N_7678,N_7251,N_7374);
xnor U7679 (N_7679,N_7459,N_7333);
and U7680 (N_7680,N_7261,N_7259);
xor U7681 (N_7681,N_7425,N_7271);
xnor U7682 (N_7682,N_7363,N_7401);
and U7683 (N_7683,N_7462,N_7295);
nand U7684 (N_7684,N_7327,N_7269);
nor U7685 (N_7685,N_7489,N_7375);
and U7686 (N_7686,N_7452,N_7368);
nand U7687 (N_7687,N_7316,N_7433);
nor U7688 (N_7688,N_7317,N_7284);
xor U7689 (N_7689,N_7320,N_7358);
and U7690 (N_7690,N_7295,N_7321);
xor U7691 (N_7691,N_7495,N_7499);
and U7692 (N_7692,N_7265,N_7385);
or U7693 (N_7693,N_7387,N_7413);
nand U7694 (N_7694,N_7308,N_7488);
nand U7695 (N_7695,N_7355,N_7413);
xor U7696 (N_7696,N_7418,N_7484);
nand U7697 (N_7697,N_7465,N_7264);
nor U7698 (N_7698,N_7298,N_7493);
and U7699 (N_7699,N_7477,N_7410);
nand U7700 (N_7700,N_7260,N_7370);
or U7701 (N_7701,N_7394,N_7434);
and U7702 (N_7702,N_7498,N_7365);
nor U7703 (N_7703,N_7436,N_7373);
xor U7704 (N_7704,N_7455,N_7295);
nand U7705 (N_7705,N_7436,N_7267);
or U7706 (N_7706,N_7385,N_7391);
or U7707 (N_7707,N_7307,N_7434);
nand U7708 (N_7708,N_7335,N_7268);
and U7709 (N_7709,N_7377,N_7258);
xor U7710 (N_7710,N_7343,N_7349);
nand U7711 (N_7711,N_7448,N_7386);
xnor U7712 (N_7712,N_7399,N_7442);
xor U7713 (N_7713,N_7414,N_7405);
nor U7714 (N_7714,N_7465,N_7496);
nor U7715 (N_7715,N_7345,N_7312);
xnor U7716 (N_7716,N_7310,N_7316);
nand U7717 (N_7717,N_7282,N_7294);
nand U7718 (N_7718,N_7414,N_7323);
nor U7719 (N_7719,N_7257,N_7342);
xor U7720 (N_7720,N_7482,N_7361);
nor U7721 (N_7721,N_7472,N_7381);
or U7722 (N_7722,N_7473,N_7269);
nor U7723 (N_7723,N_7341,N_7475);
xor U7724 (N_7724,N_7298,N_7256);
nand U7725 (N_7725,N_7388,N_7367);
and U7726 (N_7726,N_7450,N_7314);
or U7727 (N_7727,N_7314,N_7393);
nor U7728 (N_7728,N_7479,N_7397);
xnor U7729 (N_7729,N_7340,N_7380);
xnor U7730 (N_7730,N_7320,N_7496);
xnor U7731 (N_7731,N_7488,N_7431);
xnor U7732 (N_7732,N_7340,N_7293);
or U7733 (N_7733,N_7386,N_7417);
xor U7734 (N_7734,N_7499,N_7293);
or U7735 (N_7735,N_7414,N_7487);
nand U7736 (N_7736,N_7474,N_7363);
and U7737 (N_7737,N_7495,N_7463);
nand U7738 (N_7738,N_7342,N_7434);
or U7739 (N_7739,N_7416,N_7497);
nand U7740 (N_7740,N_7479,N_7461);
nor U7741 (N_7741,N_7279,N_7478);
nand U7742 (N_7742,N_7361,N_7487);
nor U7743 (N_7743,N_7435,N_7420);
and U7744 (N_7744,N_7253,N_7470);
xnor U7745 (N_7745,N_7402,N_7399);
nand U7746 (N_7746,N_7363,N_7325);
or U7747 (N_7747,N_7345,N_7373);
nand U7748 (N_7748,N_7475,N_7468);
or U7749 (N_7749,N_7371,N_7383);
or U7750 (N_7750,N_7533,N_7737);
nor U7751 (N_7751,N_7578,N_7671);
nor U7752 (N_7752,N_7733,N_7560);
and U7753 (N_7753,N_7701,N_7728);
or U7754 (N_7754,N_7515,N_7504);
xor U7755 (N_7755,N_7539,N_7691);
xnor U7756 (N_7756,N_7653,N_7627);
and U7757 (N_7757,N_7554,N_7657);
xnor U7758 (N_7758,N_7517,N_7615);
and U7759 (N_7759,N_7553,N_7664);
xor U7760 (N_7760,N_7534,N_7744);
or U7761 (N_7761,N_7655,N_7642);
xnor U7762 (N_7762,N_7654,N_7593);
nor U7763 (N_7763,N_7687,N_7723);
xor U7764 (N_7764,N_7632,N_7567);
and U7765 (N_7765,N_7693,N_7641);
nand U7766 (N_7766,N_7512,N_7611);
nand U7767 (N_7767,N_7636,N_7531);
nor U7768 (N_7768,N_7638,N_7573);
nand U7769 (N_7769,N_7536,N_7588);
nor U7770 (N_7770,N_7652,N_7633);
xnor U7771 (N_7771,N_7678,N_7511);
xor U7772 (N_7772,N_7543,N_7571);
nor U7773 (N_7773,N_7689,N_7587);
nand U7774 (N_7774,N_7563,N_7676);
or U7775 (N_7775,N_7736,N_7711);
nand U7776 (N_7776,N_7530,N_7518);
nor U7777 (N_7777,N_7668,N_7629);
xor U7778 (N_7778,N_7625,N_7637);
nor U7779 (N_7779,N_7730,N_7697);
and U7780 (N_7780,N_7714,N_7523);
or U7781 (N_7781,N_7510,N_7501);
nor U7782 (N_7782,N_7516,N_7525);
xnor U7783 (N_7783,N_7545,N_7538);
xnor U7784 (N_7784,N_7575,N_7639);
xnor U7785 (N_7785,N_7547,N_7577);
nor U7786 (N_7786,N_7631,N_7662);
or U7787 (N_7787,N_7708,N_7665);
nor U7788 (N_7788,N_7595,N_7734);
nor U7789 (N_7789,N_7596,N_7648);
xnor U7790 (N_7790,N_7601,N_7572);
or U7791 (N_7791,N_7581,N_7696);
nand U7792 (N_7792,N_7600,N_7570);
or U7793 (N_7793,N_7508,N_7589);
and U7794 (N_7794,N_7568,N_7540);
xnor U7795 (N_7795,N_7550,N_7594);
nand U7796 (N_7796,N_7695,N_7684);
xor U7797 (N_7797,N_7564,N_7729);
and U7798 (N_7798,N_7738,N_7565);
nand U7799 (N_7799,N_7619,N_7746);
nor U7800 (N_7800,N_7704,N_7592);
xor U7801 (N_7801,N_7614,N_7609);
nand U7802 (N_7802,N_7707,N_7732);
or U7803 (N_7803,N_7507,N_7505);
nor U7804 (N_7804,N_7698,N_7712);
nor U7805 (N_7805,N_7608,N_7556);
nor U7806 (N_7806,N_7586,N_7569);
xnor U7807 (N_7807,N_7705,N_7605);
xnor U7808 (N_7808,N_7502,N_7725);
or U7809 (N_7809,N_7672,N_7719);
nand U7810 (N_7810,N_7503,N_7535);
nor U7811 (N_7811,N_7727,N_7529);
nand U7812 (N_7812,N_7717,N_7514);
xnor U7813 (N_7813,N_7557,N_7667);
xor U7814 (N_7814,N_7740,N_7661);
nand U7815 (N_7815,N_7663,N_7674);
xnor U7816 (N_7816,N_7585,N_7643);
nor U7817 (N_7817,N_7690,N_7724);
or U7818 (N_7818,N_7673,N_7716);
xnor U7819 (N_7819,N_7542,N_7656);
xor U7820 (N_7820,N_7602,N_7669);
nor U7821 (N_7821,N_7660,N_7618);
nand U7822 (N_7822,N_7699,N_7620);
nor U7823 (N_7823,N_7709,N_7621);
nor U7824 (N_7824,N_7509,N_7552);
xnor U7825 (N_7825,N_7616,N_7541);
or U7826 (N_7826,N_7623,N_7537);
or U7827 (N_7827,N_7628,N_7650);
nand U7828 (N_7828,N_7692,N_7703);
nand U7829 (N_7829,N_7558,N_7574);
xnor U7830 (N_7830,N_7610,N_7549);
nor U7831 (N_7831,N_7670,N_7635);
and U7832 (N_7832,N_7688,N_7706);
nor U7833 (N_7833,N_7520,N_7582);
and U7834 (N_7834,N_7526,N_7584);
nor U7835 (N_7835,N_7710,N_7513);
or U7836 (N_7836,N_7713,N_7718);
nor U7837 (N_7837,N_7651,N_7722);
or U7838 (N_7838,N_7561,N_7735);
xor U7839 (N_7839,N_7646,N_7626);
nor U7840 (N_7840,N_7521,N_7527);
nor U7841 (N_7841,N_7745,N_7683);
and U7842 (N_7842,N_7694,N_7607);
nand U7843 (N_7843,N_7548,N_7721);
and U7844 (N_7844,N_7528,N_7658);
and U7845 (N_7845,N_7685,N_7603);
or U7846 (N_7846,N_7583,N_7686);
nand U7847 (N_7847,N_7680,N_7524);
nor U7848 (N_7848,N_7580,N_7742);
and U7849 (N_7849,N_7640,N_7579);
and U7850 (N_7850,N_7598,N_7562);
or U7851 (N_7851,N_7624,N_7613);
or U7852 (N_7852,N_7597,N_7715);
or U7853 (N_7853,N_7634,N_7647);
or U7854 (N_7854,N_7681,N_7576);
xor U7855 (N_7855,N_7612,N_7500);
nand U7856 (N_7856,N_7649,N_7559);
and U7857 (N_7857,N_7555,N_7743);
and U7858 (N_7858,N_7566,N_7700);
nor U7859 (N_7859,N_7677,N_7544);
nor U7860 (N_7860,N_7679,N_7739);
or U7861 (N_7861,N_7702,N_7604);
xnor U7862 (N_7862,N_7630,N_7659);
and U7863 (N_7863,N_7522,N_7726);
and U7864 (N_7864,N_7644,N_7519);
or U7865 (N_7865,N_7532,N_7675);
nor U7866 (N_7866,N_7617,N_7741);
or U7867 (N_7867,N_7590,N_7682);
and U7868 (N_7868,N_7606,N_7622);
xnor U7869 (N_7869,N_7546,N_7749);
and U7870 (N_7870,N_7720,N_7645);
or U7871 (N_7871,N_7591,N_7666);
nor U7872 (N_7872,N_7747,N_7599);
nor U7873 (N_7873,N_7748,N_7551);
nor U7874 (N_7874,N_7731,N_7506);
nor U7875 (N_7875,N_7735,N_7703);
xnor U7876 (N_7876,N_7623,N_7709);
nand U7877 (N_7877,N_7614,N_7601);
nand U7878 (N_7878,N_7507,N_7708);
or U7879 (N_7879,N_7551,N_7565);
nand U7880 (N_7880,N_7650,N_7609);
xnor U7881 (N_7881,N_7646,N_7648);
or U7882 (N_7882,N_7645,N_7603);
nand U7883 (N_7883,N_7666,N_7583);
xor U7884 (N_7884,N_7539,N_7676);
xor U7885 (N_7885,N_7724,N_7610);
nand U7886 (N_7886,N_7705,N_7741);
and U7887 (N_7887,N_7669,N_7719);
and U7888 (N_7888,N_7729,N_7698);
and U7889 (N_7889,N_7545,N_7602);
or U7890 (N_7890,N_7659,N_7555);
nand U7891 (N_7891,N_7588,N_7619);
nand U7892 (N_7892,N_7512,N_7749);
nor U7893 (N_7893,N_7595,N_7533);
nand U7894 (N_7894,N_7703,N_7670);
nand U7895 (N_7895,N_7643,N_7587);
and U7896 (N_7896,N_7656,N_7625);
nor U7897 (N_7897,N_7732,N_7728);
and U7898 (N_7898,N_7736,N_7634);
nand U7899 (N_7899,N_7549,N_7670);
xor U7900 (N_7900,N_7581,N_7569);
xor U7901 (N_7901,N_7673,N_7629);
or U7902 (N_7902,N_7664,N_7527);
nand U7903 (N_7903,N_7604,N_7669);
or U7904 (N_7904,N_7682,N_7586);
xnor U7905 (N_7905,N_7515,N_7506);
or U7906 (N_7906,N_7736,N_7632);
nor U7907 (N_7907,N_7545,N_7565);
and U7908 (N_7908,N_7519,N_7526);
and U7909 (N_7909,N_7542,N_7705);
nor U7910 (N_7910,N_7582,N_7618);
xor U7911 (N_7911,N_7693,N_7741);
nor U7912 (N_7912,N_7711,N_7703);
xor U7913 (N_7913,N_7722,N_7503);
xor U7914 (N_7914,N_7551,N_7704);
or U7915 (N_7915,N_7578,N_7567);
nand U7916 (N_7916,N_7545,N_7573);
nand U7917 (N_7917,N_7664,N_7638);
nand U7918 (N_7918,N_7560,N_7727);
nand U7919 (N_7919,N_7741,N_7528);
xor U7920 (N_7920,N_7741,N_7655);
and U7921 (N_7921,N_7515,N_7678);
xnor U7922 (N_7922,N_7734,N_7730);
or U7923 (N_7923,N_7527,N_7684);
and U7924 (N_7924,N_7573,N_7746);
xor U7925 (N_7925,N_7551,N_7712);
xnor U7926 (N_7926,N_7665,N_7650);
or U7927 (N_7927,N_7632,N_7652);
nand U7928 (N_7928,N_7690,N_7607);
or U7929 (N_7929,N_7543,N_7627);
and U7930 (N_7930,N_7739,N_7569);
or U7931 (N_7931,N_7740,N_7571);
and U7932 (N_7932,N_7611,N_7550);
nor U7933 (N_7933,N_7625,N_7546);
or U7934 (N_7934,N_7668,N_7525);
or U7935 (N_7935,N_7719,N_7566);
nand U7936 (N_7936,N_7739,N_7640);
xor U7937 (N_7937,N_7608,N_7599);
and U7938 (N_7938,N_7516,N_7633);
nand U7939 (N_7939,N_7583,N_7722);
or U7940 (N_7940,N_7696,N_7667);
or U7941 (N_7941,N_7619,N_7550);
xnor U7942 (N_7942,N_7603,N_7712);
nand U7943 (N_7943,N_7586,N_7729);
or U7944 (N_7944,N_7747,N_7524);
nand U7945 (N_7945,N_7600,N_7526);
nor U7946 (N_7946,N_7702,N_7628);
or U7947 (N_7947,N_7620,N_7548);
nor U7948 (N_7948,N_7514,N_7584);
xnor U7949 (N_7949,N_7647,N_7664);
or U7950 (N_7950,N_7524,N_7513);
or U7951 (N_7951,N_7573,N_7535);
or U7952 (N_7952,N_7594,N_7507);
and U7953 (N_7953,N_7647,N_7512);
nand U7954 (N_7954,N_7619,N_7508);
xnor U7955 (N_7955,N_7744,N_7573);
nand U7956 (N_7956,N_7570,N_7506);
xor U7957 (N_7957,N_7614,N_7690);
nor U7958 (N_7958,N_7655,N_7625);
xnor U7959 (N_7959,N_7541,N_7524);
and U7960 (N_7960,N_7603,N_7734);
and U7961 (N_7961,N_7616,N_7522);
and U7962 (N_7962,N_7621,N_7708);
nor U7963 (N_7963,N_7669,N_7737);
and U7964 (N_7964,N_7563,N_7642);
or U7965 (N_7965,N_7510,N_7515);
nand U7966 (N_7966,N_7540,N_7738);
nor U7967 (N_7967,N_7691,N_7572);
nand U7968 (N_7968,N_7567,N_7639);
xnor U7969 (N_7969,N_7701,N_7583);
or U7970 (N_7970,N_7624,N_7638);
or U7971 (N_7971,N_7589,N_7510);
nand U7972 (N_7972,N_7719,N_7583);
nand U7973 (N_7973,N_7664,N_7509);
xor U7974 (N_7974,N_7618,N_7540);
nand U7975 (N_7975,N_7624,N_7730);
nand U7976 (N_7976,N_7553,N_7732);
nor U7977 (N_7977,N_7529,N_7592);
xor U7978 (N_7978,N_7575,N_7603);
and U7979 (N_7979,N_7721,N_7515);
xnor U7980 (N_7980,N_7747,N_7563);
nor U7981 (N_7981,N_7613,N_7681);
and U7982 (N_7982,N_7705,N_7522);
xor U7983 (N_7983,N_7664,N_7539);
xor U7984 (N_7984,N_7686,N_7508);
and U7985 (N_7985,N_7578,N_7510);
or U7986 (N_7986,N_7651,N_7535);
nor U7987 (N_7987,N_7711,N_7714);
nand U7988 (N_7988,N_7600,N_7573);
or U7989 (N_7989,N_7528,N_7623);
xor U7990 (N_7990,N_7609,N_7705);
xor U7991 (N_7991,N_7641,N_7553);
nand U7992 (N_7992,N_7639,N_7633);
xor U7993 (N_7993,N_7715,N_7635);
and U7994 (N_7994,N_7615,N_7692);
or U7995 (N_7995,N_7598,N_7611);
nand U7996 (N_7996,N_7697,N_7577);
nor U7997 (N_7997,N_7705,N_7631);
and U7998 (N_7998,N_7551,N_7745);
or U7999 (N_7999,N_7552,N_7569);
nor U8000 (N_8000,N_7859,N_7997);
xor U8001 (N_8001,N_7967,N_7889);
nand U8002 (N_8002,N_7767,N_7879);
and U8003 (N_8003,N_7944,N_7939);
nor U8004 (N_8004,N_7918,N_7917);
and U8005 (N_8005,N_7894,N_7846);
or U8006 (N_8006,N_7972,N_7799);
xnor U8007 (N_8007,N_7842,N_7924);
nand U8008 (N_8008,N_7773,N_7772);
nor U8009 (N_8009,N_7943,N_7810);
and U8010 (N_8010,N_7996,N_7985);
nor U8011 (N_8011,N_7788,N_7835);
or U8012 (N_8012,N_7770,N_7963);
xor U8013 (N_8013,N_7969,N_7813);
nor U8014 (N_8014,N_7957,N_7960);
nor U8015 (N_8015,N_7932,N_7885);
and U8016 (N_8016,N_7954,N_7838);
nor U8017 (N_8017,N_7948,N_7914);
nor U8018 (N_8018,N_7911,N_7760);
nand U8019 (N_8019,N_7941,N_7916);
nand U8020 (N_8020,N_7905,N_7961);
or U8021 (N_8021,N_7909,N_7789);
or U8022 (N_8022,N_7869,N_7796);
or U8023 (N_8023,N_7982,N_7968);
and U8024 (N_8024,N_7890,N_7833);
or U8025 (N_8025,N_7784,N_7983);
nand U8026 (N_8026,N_7975,N_7834);
nor U8027 (N_8027,N_7930,N_7964);
and U8028 (N_8028,N_7949,N_7830);
nor U8029 (N_8029,N_7761,N_7962);
xnor U8030 (N_8030,N_7792,N_7808);
and U8031 (N_8031,N_7823,N_7915);
and U8032 (N_8032,N_7886,N_7920);
or U8033 (N_8033,N_7922,N_7874);
and U8034 (N_8034,N_7936,N_7990);
and U8035 (N_8035,N_7801,N_7805);
nor U8036 (N_8036,N_7933,N_7853);
xnor U8037 (N_8037,N_7979,N_7892);
nand U8038 (N_8038,N_7844,N_7898);
xor U8039 (N_8039,N_7751,N_7921);
or U8040 (N_8040,N_7955,N_7947);
xor U8041 (N_8041,N_7896,N_7871);
nor U8042 (N_8042,N_7926,N_7821);
nor U8043 (N_8043,N_7815,N_7897);
or U8044 (N_8044,N_7803,N_7895);
nand U8045 (N_8045,N_7904,N_7925);
or U8046 (N_8046,N_7816,N_7980);
xor U8047 (N_8047,N_7752,N_7976);
nor U8048 (N_8048,N_7776,N_7951);
and U8049 (N_8049,N_7876,N_7857);
nor U8050 (N_8050,N_7848,N_7882);
or U8051 (N_8051,N_7800,N_7927);
nand U8052 (N_8052,N_7817,N_7880);
nor U8053 (N_8053,N_7866,N_7902);
xor U8054 (N_8054,N_7900,N_7849);
nand U8055 (N_8055,N_7858,N_7820);
or U8056 (N_8056,N_7868,N_7974);
xor U8057 (N_8057,N_7806,N_7850);
nand U8058 (N_8058,N_7824,N_7756);
xnor U8059 (N_8059,N_7856,N_7901);
and U8060 (N_8060,N_7797,N_7910);
and U8061 (N_8061,N_7795,N_7931);
and U8062 (N_8062,N_7989,N_7769);
or U8063 (N_8063,N_7771,N_7995);
or U8064 (N_8064,N_7865,N_7785);
xnor U8065 (N_8065,N_7836,N_7781);
xor U8066 (N_8066,N_7791,N_7863);
or U8067 (N_8067,N_7998,N_7854);
xor U8068 (N_8068,N_7987,N_7811);
or U8069 (N_8069,N_7753,N_7822);
nor U8070 (N_8070,N_7937,N_7966);
xor U8071 (N_8071,N_7994,N_7837);
xnor U8072 (N_8072,N_7958,N_7766);
nor U8073 (N_8073,N_7794,N_7971);
or U8074 (N_8074,N_7888,N_7764);
nor U8075 (N_8075,N_7919,N_7775);
or U8076 (N_8076,N_7754,N_7790);
nand U8077 (N_8077,N_7814,N_7873);
nor U8078 (N_8078,N_7782,N_7950);
or U8079 (N_8079,N_7765,N_7906);
nand U8080 (N_8080,N_7829,N_7907);
and U8081 (N_8081,N_7929,N_7992);
xnor U8082 (N_8082,N_7956,N_7774);
nor U8083 (N_8083,N_7913,N_7807);
and U8084 (N_8084,N_7938,N_7988);
nor U8085 (N_8085,N_7851,N_7779);
xnor U8086 (N_8086,N_7965,N_7783);
and U8087 (N_8087,N_7942,N_7841);
nand U8088 (N_8088,N_7946,N_7828);
nand U8089 (N_8089,N_7993,N_7777);
and U8090 (N_8090,N_7970,N_7867);
or U8091 (N_8091,N_7780,N_7945);
nor U8092 (N_8092,N_7755,N_7818);
xnor U8093 (N_8093,N_7875,N_7881);
nand U8094 (N_8094,N_7861,N_7750);
xor U8095 (N_8095,N_7877,N_7884);
nand U8096 (N_8096,N_7862,N_7798);
nor U8097 (N_8097,N_7762,N_7845);
and U8098 (N_8098,N_7959,N_7986);
xor U8099 (N_8099,N_7809,N_7860);
xor U8100 (N_8100,N_7840,N_7903);
or U8101 (N_8101,N_7826,N_7847);
or U8102 (N_8102,N_7977,N_7758);
or U8103 (N_8103,N_7832,N_7893);
or U8104 (N_8104,N_7827,N_7831);
nand U8105 (N_8105,N_7883,N_7940);
and U8106 (N_8106,N_7991,N_7887);
nor U8107 (N_8107,N_7935,N_7899);
xor U8108 (N_8108,N_7934,N_7973);
nand U8109 (N_8109,N_7778,N_7757);
or U8110 (N_8110,N_7759,N_7864);
or U8111 (N_8111,N_7852,N_7786);
or U8112 (N_8112,N_7981,N_7928);
xor U8113 (N_8113,N_7908,N_7804);
nor U8114 (N_8114,N_7802,N_7839);
nand U8115 (N_8115,N_7870,N_7768);
xnor U8116 (N_8116,N_7999,N_7912);
xnor U8117 (N_8117,N_7763,N_7978);
and U8118 (N_8118,N_7843,N_7952);
or U8119 (N_8119,N_7872,N_7787);
nor U8120 (N_8120,N_7825,N_7878);
nor U8121 (N_8121,N_7984,N_7953);
nor U8122 (N_8122,N_7891,N_7819);
nor U8123 (N_8123,N_7855,N_7812);
nand U8124 (N_8124,N_7793,N_7923);
nor U8125 (N_8125,N_7983,N_7981);
nor U8126 (N_8126,N_7827,N_7987);
nor U8127 (N_8127,N_7930,N_7941);
nor U8128 (N_8128,N_7826,N_7827);
and U8129 (N_8129,N_7897,N_7932);
nor U8130 (N_8130,N_7801,N_7887);
or U8131 (N_8131,N_7986,N_7818);
xor U8132 (N_8132,N_7853,N_7979);
and U8133 (N_8133,N_7910,N_7879);
xnor U8134 (N_8134,N_7762,N_7759);
and U8135 (N_8135,N_7987,N_7995);
or U8136 (N_8136,N_7908,N_7774);
xnor U8137 (N_8137,N_7951,N_7807);
nor U8138 (N_8138,N_7964,N_7771);
or U8139 (N_8139,N_7975,N_7985);
and U8140 (N_8140,N_7804,N_7771);
and U8141 (N_8141,N_7929,N_7941);
nor U8142 (N_8142,N_7841,N_7816);
and U8143 (N_8143,N_7980,N_7859);
and U8144 (N_8144,N_7805,N_7971);
or U8145 (N_8145,N_7781,N_7753);
nor U8146 (N_8146,N_7823,N_7761);
nor U8147 (N_8147,N_7968,N_7804);
xnor U8148 (N_8148,N_7961,N_7867);
or U8149 (N_8149,N_7765,N_7778);
nand U8150 (N_8150,N_7875,N_7977);
xor U8151 (N_8151,N_7854,N_7992);
xnor U8152 (N_8152,N_7875,N_7781);
nand U8153 (N_8153,N_7897,N_7936);
or U8154 (N_8154,N_7792,N_7995);
and U8155 (N_8155,N_7953,N_7819);
xnor U8156 (N_8156,N_7823,N_7868);
nor U8157 (N_8157,N_7854,N_7966);
and U8158 (N_8158,N_7873,N_7962);
or U8159 (N_8159,N_7979,N_7859);
nand U8160 (N_8160,N_7942,N_7950);
or U8161 (N_8161,N_7906,N_7756);
or U8162 (N_8162,N_7759,N_7786);
and U8163 (N_8163,N_7827,N_7767);
nand U8164 (N_8164,N_7825,N_7912);
nor U8165 (N_8165,N_7938,N_7874);
and U8166 (N_8166,N_7895,N_7816);
or U8167 (N_8167,N_7929,N_7827);
and U8168 (N_8168,N_7857,N_7928);
and U8169 (N_8169,N_7897,N_7768);
and U8170 (N_8170,N_7862,N_7817);
nor U8171 (N_8171,N_7858,N_7753);
nand U8172 (N_8172,N_7860,N_7972);
and U8173 (N_8173,N_7768,N_7908);
nand U8174 (N_8174,N_7910,N_7911);
nand U8175 (N_8175,N_7869,N_7892);
xor U8176 (N_8176,N_7941,N_7765);
and U8177 (N_8177,N_7878,N_7833);
nor U8178 (N_8178,N_7883,N_7992);
nor U8179 (N_8179,N_7993,N_7836);
xor U8180 (N_8180,N_7775,N_7933);
and U8181 (N_8181,N_7919,N_7865);
nand U8182 (N_8182,N_7896,N_7876);
or U8183 (N_8183,N_7888,N_7913);
or U8184 (N_8184,N_7896,N_7964);
or U8185 (N_8185,N_7824,N_7753);
nand U8186 (N_8186,N_7872,N_7944);
nor U8187 (N_8187,N_7999,N_7887);
nor U8188 (N_8188,N_7835,N_7840);
nor U8189 (N_8189,N_7924,N_7887);
and U8190 (N_8190,N_7853,N_7942);
nand U8191 (N_8191,N_7804,N_7843);
and U8192 (N_8192,N_7835,N_7851);
or U8193 (N_8193,N_7867,N_7892);
xnor U8194 (N_8194,N_7816,N_7924);
nand U8195 (N_8195,N_7792,N_7890);
and U8196 (N_8196,N_7935,N_7794);
or U8197 (N_8197,N_7882,N_7993);
and U8198 (N_8198,N_7995,N_7824);
xnor U8199 (N_8199,N_7925,N_7795);
nor U8200 (N_8200,N_7857,N_7886);
nand U8201 (N_8201,N_7879,N_7941);
nand U8202 (N_8202,N_7835,N_7798);
and U8203 (N_8203,N_7947,N_7998);
or U8204 (N_8204,N_7917,N_7977);
or U8205 (N_8205,N_7770,N_7763);
and U8206 (N_8206,N_7959,N_7857);
xnor U8207 (N_8207,N_7859,N_7951);
nand U8208 (N_8208,N_7948,N_7966);
or U8209 (N_8209,N_7892,N_7995);
nand U8210 (N_8210,N_7851,N_7793);
or U8211 (N_8211,N_7866,N_7969);
or U8212 (N_8212,N_7827,N_7762);
and U8213 (N_8213,N_7883,N_7902);
xnor U8214 (N_8214,N_7766,N_7912);
and U8215 (N_8215,N_7960,N_7913);
or U8216 (N_8216,N_7952,N_7827);
xnor U8217 (N_8217,N_7921,N_7778);
nor U8218 (N_8218,N_7905,N_7940);
or U8219 (N_8219,N_7908,N_7910);
xnor U8220 (N_8220,N_7830,N_7924);
and U8221 (N_8221,N_7894,N_7779);
nand U8222 (N_8222,N_7906,N_7939);
xnor U8223 (N_8223,N_7824,N_7809);
or U8224 (N_8224,N_7992,N_7978);
xnor U8225 (N_8225,N_7879,N_7929);
nor U8226 (N_8226,N_7799,N_7759);
nor U8227 (N_8227,N_7959,N_7759);
and U8228 (N_8228,N_7968,N_7781);
and U8229 (N_8229,N_7828,N_7861);
or U8230 (N_8230,N_7795,N_7982);
xnor U8231 (N_8231,N_7819,N_7790);
or U8232 (N_8232,N_7834,N_7777);
nor U8233 (N_8233,N_7771,N_7810);
xor U8234 (N_8234,N_7942,N_7756);
nand U8235 (N_8235,N_7874,N_7843);
nand U8236 (N_8236,N_7775,N_7906);
and U8237 (N_8237,N_7964,N_7973);
or U8238 (N_8238,N_7809,N_7898);
nor U8239 (N_8239,N_7912,N_7838);
nand U8240 (N_8240,N_7778,N_7815);
nand U8241 (N_8241,N_7944,N_7992);
nand U8242 (N_8242,N_7752,N_7848);
or U8243 (N_8243,N_7977,N_7877);
and U8244 (N_8244,N_7766,N_7828);
xnor U8245 (N_8245,N_7934,N_7897);
and U8246 (N_8246,N_7758,N_7993);
or U8247 (N_8247,N_7752,N_7771);
nand U8248 (N_8248,N_7939,N_7910);
nand U8249 (N_8249,N_7857,N_7867);
xnor U8250 (N_8250,N_8016,N_8113);
xnor U8251 (N_8251,N_8082,N_8164);
and U8252 (N_8252,N_8070,N_8209);
nand U8253 (N_8253,N_8065,N_8168);
and U8254 (N_8254,N_8110,N_8138);
nor U8255 (N_8255,N_8066,N_8229);
xor U8256 (N_8256,N_8118,N_8081);
xnor U8257 (N_8257,N_8100,N_8183);
or U8258 (N_8258,N_8121,N_8028);
or U8259 (N_8259,N_8238,N_8015);
xor U8260 (N_8260,N_8205,N_8031);
and U8261 (N_8261,N_8071,N_8079);
nor U8262 (N_8262,N_8034,N_8068);
xnor U8263 (N_8263,N_8024,N_8010);
or U8264 (N_8264,N_8094,N_8074);
nor U8265 (N_8265,N_8241,N_8086);
nor U8266 (N_8266,N_8102,N_8053);
xor U8267 (N_8267,N_8109,N_8046);
nor U8268 (N_8268,N_8043,N_8129);
or U8269 (N_8269,N_8146,N_8096);
or U8270 (N_8270,N_8078,N_8222);
xnor U8271 (N_8271,N_8063,N_8149);
or U8272 (N_8272,N_8088,N_8181);
nor U8273 (N_8273,N_8214,N_8220);
xor U8274 (N_8274,N_8187,N_8002);
nor U8275 (N_8275,N_8178,N_8166);
and U8276 (N_8276,N_8120,N_8007);
and U8277 (N_8277,N_8006,N_8038);
or U8278 (N_8278,N_8116,N_8199);
nor U8279 (N_8279,N_8162,N_8221);
xnor U8280 (N_8280,N_8215,N_8223);
nor U8281 (N_8281,N_8182,N_8021);
nand U8282 (N_8282,N_8210,N_8026);
nand U8283 (N_8283,N_8114,N_8119);
xor U8284 (N_8284,N_8135,N_8005);
nor U8285 (N_8285,N_8092,N_8128);
nor U8286 (N_8286,N_8151,N_8226);
nor U8287 (N_8287,N_8051,N_8143);
nand U8288 (N_8288,N_8103,N_8052);
nand U8289 (N_8289,N_8018,N_8206);
nor U8290 (N_8290,N_8228,N_8011);
nand U8291 (N_8291,N_8249,N_8171);
or U8292 (N_8292,N_8035,N_8244);
nor U8293 (N_8293,N_8224,N_8083);
or U8294 (N_8294,N_8230,N_8247);
and U8295 (N_8295,N_8219,N_8055);
nor U8296 (N_8296,N_8087,N_8044);
nand U8297 (N_8297,N_8003,N_8159);
nor U8298 (N_8298,N_8165,N_8172);
and U8299 (N_8299,N_8148,N_8157);
nand U8300 (N_8300,N_8216,N_8132);
nand U8301 (N_8301,N_8158,N_8144);
and U8302 (N_8302,N_8195,N_8036);
nand U8303 (N_8303,N_8008,N_8170);
nand U8304 (N_8304,N_8064,N_8204);
nor U8305 (N_8305,N_8101,N_8232);
and U8306 (N_8306,N_8147,N_8192);
nand U8307 (N_8307,N_8042,N_8115);
xnor U8308 (N_8308,N_8059,N_8175);
xnor U8309 (N_8309,N_8145,N_8123);
or U8310 (N_8310,N_8106,N_8240);
nor U8311 (N_8311,N_8075,N_8033);
nor U8312 (N_8312,N_8095,N_8067);
nor U8313 (N_8313,N_8242,N_8212);
nand U8314 (N_8314,N_8069,N_8248);
xor U8315 (N_8315,N_8200,N_8030);
xnor U8316 (N_8316,N_8025,N_8104);
or U8317 (N_8317,N_8174,N_8217);
or U8318 (N_8318,N_8213,N_8133);
nor U8319 (N_8319,N_8156,N_8137);
nor U8320 (N_8320,N_8169,N_8084);
nand U8321 (N_8321,N_8239,N_8191);
nand U8322 (N_8322,N_8227,N_8093);
nand U8323 (N_8323,N_8009,N_8020);
nand U8324 (N_8324,N_8014,N_8139);
nand U8325 (N_8325,N_8180,N_8176);
nand U8326 (N_8326,N_8040,N_8189);
or U8327 (N_8327,N_8202,N_8184);
or U8328 (N_8328,N_8140,N_8203);
and U8329 (N_8329,N_8054,N_8000);
nand U8330 (N_8330,N_8207,N_8185);
xnor U8331 (N_8331,N_8237,N_8029);
and U8332 (N_8332,N_8173,N_8022);
and U8333 (N_8333,N_8134,N_8197);
xor U8334 (N_8334,N_8233,N_8124);
nor U8335 (N_8335,N_8179,N_8056);
xor U8336 (N_8336,N_8152,N_8057);
and U8337 (N_8337,N_8154,N_8194);
xnor U8338 (N_8338,N_8039,N_8050);
or U8339 (N_8339,N_8019,N_8072);
nor U8340 (N_8340,N_8231,N_8125);
nand U8341 (N_8341,N_8001,N_8193);
nor U8342 (N_8342,N_8190,N_8186);
nor U8343 (N_8343,N_8073,N_8004);
or U8344 (N_8344,N_8126,N_8023);
or U8345 (N_8345,N_8127,N_8198);
or U8346 (N_8346,N_8098,N_8012);
nor U8347 (N_8347,N_8047,N_8099);
or U8348 (N_8348,N_8243,N_8142);
nand U8349 (N_8349,N_8060,N_8234);
and U8350 (N_8350,N_8136,N_8013);
nand U8351 (N_8351,N_8153,N_8048);
and U8352 (N_8352,N_8049,N_8235);
nor U8353 (N_8353,N_8076,N_8117);
nand U8354 (N_8354,N_8211,N_8150);
xor U8355 (N_8355,N_8027,N_8045);
or U8356 (N_8356,N_8111,N_8077);
nand U8357 (N_8357,N_8061,N_8208);
xor U8358 (N_8358,N_8160,N_8091);
and U8359 (N_8359,N_8167,N_8163);
xor U8360 (N_8360,N_8085,N_8218);
xnor U8361 (N_8361,N_8130,N_8058);
or U8362 (N_8362,N_8236,N_8017);
or U8363 (N_8363,N_8161,N_8177);
or U8364 (N_8364,N_8141,N_8041);
xnor U8365 (N_8365,N_8196,N_8131);
and U8366 (N_8366,N_8080,N_8062);
nand U8367 (N_8367,N_8105,N_8188);
or U8368 (N_8368,N_8037,N_8032);
xnor U8369 (N_8369,N_8225,N_8089);
or U8370 (N_8370,N_8097,N_8201);
or U8371 (N_8371,N_8245,N_8107);
xor U8372 (N_8372,N_8246,N_8090);
or U8373 (N_8373,N_8112,N_8122);
nor U8374 (N_8374,N_8108,N_8155);
or U8375 (N_8375,N_8171,N_8240);
or U8376 (N_8376,N_8164,N_8115);
or U8377 (N_8377,N_8109,N_8029);
and U8378 (N_8378,N_8221,N_8006);
nand U8379 (N_8379,N_8191,N_8016);
xnor U8380 (N_8380,N_8236,N_8089);
and U8381 (N_8381,N_8106,N_8185);
or U8382 (N_8382,N_8228,N_8146);
and U8383 (N_8383,N_8019,N_8009);
and U8384 (N_8384,N_8191,N_8117);
xor U8385 (N_8385,N_8175,N_8026);
nor U8386 (N_8386,N_8244,N_8246);
xor U8387 (N_8387,N_8155,N_8185);
or U8388 (N_8388,N_8141,N_8124);
nor U8389 (N_8389,N_8077,N_8177);
nor U8390 (N_8390,N_8197,N_8086);
or U8391 (N_8391,N_8157,N_8172);
nor U8392 (N_8392,N_8218,N_8174);
nand U8393 (N_8393,N_8000,N_8049);
nand U8394 (N_8394,N_8223,N_8141);
nor U8395 (N_8395,N_8029,N_8034);
xnor U8396 (N_8396,N_8171,N_8197);
xnor U8397 (N_8397,N_8013,N_8218);
or U8398 (N_8398,N_8114,N_8198);
nor U8399 (N_8399,N_8166,N_8054);
xnor U8400 (N_8400,N_8193,N_8223);
nor U8401 (N_8401,N_8240,N_8000);
or U8402 (N_8402,N_8038,N_8198);
or U8403 (N_8403,N_8197,N_8209);
xor U8404 (N_8404,N_8045,N_8103);
xnor U8405 (N_8405,N_8154,N_8079);
xor U8406 (N_8406,N_8172,N_8227);
or U8407 (N_8407,N_8021,N_8080);
nor U8408 (N_8408,N_8186,N_8157);
nor U8409 (N_8409,N_8061,N_8239);
nand U8410 (N_8410,N_8195,N_8118);
nor U8411 (N_8411,N_8014,N_8053);
or U8412 (N_8412,N_8097,N_8214);
and U8413 (N_8413,N_8103,N_8047);
or U8414 (N_8414,N_8116,N_8070);
nand U8415 (N_8415,N_8087,N_8056);
nand U8416 (N_8416,N_8142,N_8219);
nor U8417 (N_8417,N_8032,N_8049);
xnor U8418 (N_8418,N_8180,N_8101);
nor U8419 (N_8419,N_8027,N_8125);
nand U8420 (N_8420,N_8060,N_8248);
nor U8421 (N_8421,N_8127,N_8212);
nor U8422 (N_8422,N_8233,N_8185);
nor U8423 (N_8423,N_8054,N_8245);
xnor U8424 (N_8424,N_8072,N_8238);
xor U8425 (N_8425,N_8023,N_8163);
xnor U8426 (N_8426,N_8163,N_8077);
nand U8427 (N_8427,N_8170,N_8009);
nand U8428 (N_8428,N_8010,N_8090);
xor U8429 (N_8429,N_8127,N_8037);
and U8430 (N_8430,N_8184,N_8232);
xnor U8431 (N_8431,N_8191,N_8088);
nand U8432 (N_8432,N_8006,N_8166);
xor U8433 (N_8433,N_8235,N_8172);
and U8434 (N_8434,N_8119,N_8103);
or U8435 (N_8435,N_8134,N_8000);
nor U8436 (N_8436,N_8185,N_8107);
or U8437 (N_8437,N_8236,N_8079);
or U8438 (N_8438,N_8243,N_8014);
nor U8439 (N_8439,N_8035,N_8130);
nor U8440 (N_8440,N_8032,N_8022);
xnor U8441 (N_8441,N_8071,N_8166);
xnor U8442 (N_8442,N_8149,N_8074);
xor U8443 (N_8443,N_8145,N_8019);
nand U8444 (N_8444,N_8030,N_8190);
xnor U8445 (N_8445,N_8227,N_8108);
or U8446 (N_8446,N_8175,N_8007);
nor U8447 (N_8447,N_8078,N_8119);
and U8448 (N_8448,N_8122,N_8061);
or U8449 (N_8449,N_8035,N_8090);
nand U8450 (N_8450,N_8131,N_8021);
xnor U8451 (N_8451,N_8225,N_8135);
nand U8452 (N_8452,N_8061,N_8242);
nor U8453 (N_8453,N_8067,N_8068);
nor U8454 (N_8454,N_8172,N_8174);
xor U8455 (N_8455,N_8199,N_8201);
xor U8456 (N_8456,N_8089,N_8151);
nand U8457 (N_8457,N_8171,N_8222);
and U8458 (N_8458,N_8033,N_8165);
nand U8459 (N_8459,N_8174,N_8127);
xnor U8460 (N_8460,N_8192,N_8228);
and U8461 (N_8461,N_8011,N_8217);
or U8462 (N_8462,N_8048,N_8178);
and U8463 (N_8463,N_8239,N_8067);
nand U8464 (N_8464,N_8240,N_8184);
nor U8465 (N_8465,N_8184,N_8233);
xnor U8466 (N_8466,N_8216,N_8240);
or U8467 (N_8467,N_8015,N_8118);
or U8468 (N_8468,N_8113,N_8081);
and U8469 (N_8469,N_8079,N_8102);
nor U8470 (N_8470,N_8000,N_8141);
nand U8471 (N_8471,N_8240,N_8183);
and U8472 (N_8472,N_8043,N_8079);
xnor U8473 (N_8473,N_8151,N_8162);
nor U8474 (N_8474,N_8097,N_8095);
and U8475 (N_8475,N_8126,N_8219);
or U8476 (N_8476,N_8169,N_8115);
or U8477 (N_8477,N_8102,N_8239);
or U8478 (N_8478,N_8082,N_8071);
and U8479 (N_8479,N_8155,N_8064);
nor U8480 (N_8480,N_8221,N_8192);
xor U8481 (N_8481,N_8109,N_8045);
nand U8482 (N_8482,N_8131,N_8002);
and U8483 (N_8483,N_8011,N_8234);
nand U8484 (N_8484,N_8001,N_8004);
and U8485 (N_8485,N_8243,N_8192);
nand U8486 (N_8486,N_8054,N_8072);
and U8487 (N_8487,N_8219,N_8220);
or U8488 (N_8488,N_8131,N_8152);
nand U8489 (N_8489,N_8102,N_8213);
xor U8490 (N_8490,N_8070,N_8042);
and U8491 (N_8491,N_8039,N_8059);
nand U8492 (N_8492,N_8172,N_8073);
xnor U8493 (N_8493,N_8159,N_8021);
and U8494 (N_8494,N_8035,N_8072);
or U8495 (N_8495,N_8226,N_8153);
xor U8496 (N_8496,N_8047,N_8244);
nor U8497 (N_8497,N_8143,N_8139);
nand U8498 (N_8498,N_8141,N_8053);
nand U8499 (N_8499,N_8221,N_8208);
and U8500 (N_8500,N_8440,N_8494);
and U8501 (N_8501,N_8490,N_8273);
xnor U8502 (N_8502,N_8389,N_8392);
nand U8503 (N_8503,N_8493,N_8486);
xor U8504 (N_8504,N_8498,N_8446);
and U8505 (N_8505,N_8300,N_8449);
nand U8506 (N_8506,N_8483,N_8384);
xnor U8507 (N_8507,N_8285,N_8321);
and U8508 (N_8508,N_8381,N_8308);
or U8509 (N_8509,N_8290,N_8478);
or U8510 (N_8510,N_8485,N_8419);
and U8511 (N_8511,N_8338,N_8350);
and U8512 (N_8512,N_8418,N_8356);
and U8513 (N_8513,N_8432,N_8332);
nand U8514 (N_8514,N_8293,N_8266);
xor U8515 (N_8515,N_8376,N_8408);
xnor U8516 (N_8516,N_8452,N_8475);
xnor U8517 (N_8517,N_8254,N_8344);
or U8518 (N_8518,N_8468,N_8302);
or U8519 (N_8519,N_8352,N_8465);
and U8520 (N_8520,N_8433,N_8366);
nor U8521 (N_8521,N_8345,N_8393);
nand U8522 (N_8522,N_8396,N_8289);
nand U8523 (N_8523,N_8430,N_8441);
nand U8524 (N_8524,N_8445,N_8412);
and U8525 (N_8525,N_8457,N_8434);
nor U8526 (N_8526,N_8322,N_8459);
xnor U8527 (N_8527,N_8354,N_8489);
or U8528 (N_8528,N_8400,N_8280);
xnor U8529 (N_8529,N_8399,N_8355);
or U8530 (N_8530,N_8391,N_8335);
nand U8531 (N_8531,N_8436,N_8279);
nor U8532 (N_8532,N_8385,N_8390);
or U8533 (N_8533,N_8477,N_8427);
nor U8534 (N_8534,N_8346,N_8472);
nor U8535 (N_8535,N_8460,N_8402);
nand U8536 (N_8536,N_8453,N_8450);
or U8537 (N_8537,N_8303,N_8313);
nor U8538 (N_8538,N_8275,N_8469);
and U8539 (N_8539,N_8361,N_8406);
nor U8540 (N_8540,N_8455,N_8420);
or U8541 (N_8541,N_8444,N_8301);
xnor U8542 (N_8542,N_8331,N_8263);
and U8543 (N_8543,N_8487,N_8251);
nand U8544 (N_8544,N_8421,N_8476);
and U8545 (N_8545,N_8340,N_8414);
xnor U8546 (N_8546,N_8380,N_8341);
xnor U8547 (N_8547,N_8461,N_8491);
or U8548 (N_8548,N_8343,N_8497);
xor U8549 (N_8549,N_8337,N_8394);
nor U8550 (N_8550,N_8309,N_8359);
and U8551 (N_8551,N_8353,N_8388);
nor U8552 (N_8552,N_8334,N_8492);
xnor U8553 (N_8553,N_8255,N_8287);
nand U8554 (N_8554,N_8422,N_8312);
nand U8555 (N_8555,N_8306,N_8443);
or U8556 (N_8556,N_8425,N_8297);
nand U8557 (N_8557,N_8462,N_8351);
nor U8558 (N_8558,N_8265,N_8362);
nor U8559 (N_8559,N_8277,N_8458);
nor U8560 (N_8560,N_8260,N_8466);
nor U8561 (N_8561,N_8358,N_8481);
xor U8562 (N_8562,N_8496,N_8268);
nand U8563 (N_8563,N_8271,N_8298);
nand U8564 (N_8564,N_8317,N_8375);
nand U8565 (N_8565,N_8272,N_8377);
or U8566 (N_8566,N_8426,N_8473);
nand U8567 (N_8567,N_8474,N_8292);
and U8568 (N_8568,N_8274,N_8259);
xnor U8569 (N_8569,N_8296,N_8336);
nand U8570 (N_8570,N_8363,N_8314);
and U8571 (N_8571,N_8428,N_8411);
nor U8572 (N_8572,N_8387,N_8278);
and U8573 (N_8573,N_8405,N_8311);
or U8574 (N_8574,N_8294,N_8282);
nor U8575 (N_8575,N_8423,N_8398);
xnor U8576 (N_8576,N_8401,N_8382);
nor U8577 (N_8577,N_8367,N_8373);
nand U8578 (N_8578,N_8464,N_8403);
or U8579 (N_8579,N_8328,N_8495);
or U8580 (N_8580,N_8320,N_8447);
nand U8581 (N_8581,N_8325,N_8261);
and U8582 (N_8582,N_8288,N_8439);
and U8583 (N_8583,N_8295,N_8397);
or U8584 (N_8584,N_8409,N_8438);
and U8585 (N_8585,N_8270,N_8480);
and U8586 (N_8586,N_8448,N_8437);
and U8587 (N_8587,N_8404,N_8413);
xor U8588 (N_8588,N_8451,N_8499);
and U8589 (N_8589,N_8454,N_8330);
xnor U8590 (N_8590,N_8372,N_8250);
nor U8591 (N_8591,N_8281,N_8347);
and U8592 (N_8592,N_8286,N_8386);
xnor U8593 (N_8593,N_8284,N_8371);
and U8594 (N_8594,N_8417,N_8258);
and U8595 (N_8595,N_8467,N_8407);
nand U8596 (N_8596,N_8442,N_8326);
and U8597 (N_8597,N_8318,N_8379);
nor U8598 (N_8598,N_8429,N_8315);
nand U8599 (N_8599,N_8365,N_8378);
xor U8600 (N_8600,N_8267,N_8252);
nand U8601 (N_8601,N_8374,N_8276);
and U8602 (N_8602,N_8316,N_8291);
nor U8603 (N_8603,N_8435,N_8319);
or U8604 (N_8604,N_8360,N_8415);
nor U8605 (N_8605,N_8364,N_8431);
nand U8606 (N_8606,N_8348,N_8304);
nand U8607 (N_8607,N_8323,N_8256);
nand U8608 (N_8608,N_8327,N_8484);
and U8609 (N_8609,N_8324,N_8357);
and U8610 (N_8610,N_8482,N_8333);
or U8611 (N_8611,N_8463,N_8369);
xnor U8612 (N_8612,N_8349,N_8299);
or U8613 (N_8613,N_8368,N_8253);
or U8614 (N_8614,N_8310,N_8410);
xor U8615 (N_8615,N_8339,N_8305);
xor U8616 (N_8616,N_8383,N_8471);
nand U8617 (N_8617,N_8488,N_8370);
nand U8618 (N_8618,N_8479,N_8395);
nand U8619 (N_8619,N_8269,N_8342);
or U8620 (N_8620,N_8329,N_8416);
nand U8621 (N_8621,N_8456,N_8470);
xor U8622 (N_8622,N_8283,N_8424);
and U8623 (N_8623,N_8307,N_8262);
or U8624 (N_8624,N_8264,N_8257);
and U8625 (N_8625,N_8479,N_8471);
nand U8626 (N_8626,N_8417,N_8488);
nor U8627 (N_8627,N_8324,N_8404);
or U8628 (N_8628,N_8275,N_8322);
xnor U8629 (N_8629,N_8266,N_8436);
and U8630 (N_8630,N_8355,N_8309);
and U8631 (N_8631,N_8432,N_8476);
or U8632 (N_8632,N_8465,N_8389);
or U8633 (N_8633,N_8447,N_8370);
nor U8634 (N_8634,N_8391,N_8467);
or U8635 (N_8635,N_8319,N_8461);
or U8636 (N_8636,N_8377,N_8251);
and U8637 (N_8637,N_8288,N_8469);
nor U8638 (N_8638,N_8477,N_8348);
xor U8639 (N_8639,N_8353,N_8428);
nand U8640 (N_8640,N_8291,N_8381);
nand U8641 (N_8641,N_8340,N_8254);
or U8642 (N_8642,N_8253,N_8410);
or U8643 (N_8643,N_8409,N_8472);
xor U8644 (N_8644,N_8253,N_8353);
xnor U8645 (N_8645,N_8265,N_8320);
nor U8646 (N_8646,N_8326,N_8315);
or U8647 (N_8647,N_8270,N_8395);
or U8648 (N_8648,N_8478,N_8332);
and U8649 (N_8649,N_8298,N_8282);
nor U8650 (N_8650,N_8386,N_8398);
nand U8651 (N_8651,N_8442,N_8352);
xnor U8652 (N_8652,N_8264,N_8319);
nand U8653 (N_8653,N_8381,N_8361);
nand U8654 (N_8654,N_8372,N_8483);
nor U8655 (N_8655,N_8339,N_8473);
or U8656 (N_8656,N_8424,N_8413);
xor U8657 (N_8657,N_8264,N_8289);
nand U8658 (N_8658,N_8285,N_8440);
xnor U8659 (N_8659,N_8287,N_8496);
nor U8660 (N_8660,N_8377,N_8373);
or U8661 (N_8661,N_8272,N_8351);
or U8662 (N_8662,N_8478,N_8343);
xnor U8663 (N_8663,N_8414,N_8443);
or U8664 (N_8664,N_8272,N_8298);
nand U8665 (N_8665,N_8317,N_8309);
nand U8666 (N_8666,N_8269,N_8370);
nand U8667 (N_8667,N_8352,N_8253);
nor U8668 (N_8668,N_8300,N_8308);
or U8669 (N_8669,N_8498,N_8276);
or U8670 (N_8670,N_8400,N_8381);
or U8671 (N_8671,N_8360,N_8410);
or U8672 (N_8672,N_8395,N_8365);
or U8673 (N_8673,N_8299,N_8444);
or U8674 (N_8674,N_8445,N_8495);
nor U8675 (N_8675,N_8285,N_8463);
xor U8676 (N_8676,N_8429,N_8278);
and U8677 (N_8677,N_8385,N_8424);
nor U8678 (N_8678,N_8327,N_8365);
xnor U8679 (N_8679,N_8431,N_8325);
xnor U8680 (N_8680,N_8285,N_8430);
or U8681 (N_8681,N_8370,N_8260);
xor U8682 (N_8682,N_8440,N_8272);
nand U8683 (N_8683,N_8472,N_8318);
and U8684 (N_8684,N_8330,N_8293);
xnor U8685 (N_8685,N_8326,N_8320);
and U8686 (N_8686,N_8465,N_8269);
nand U8687 (N_8687,N_8392,N_8458);
nor U8688 (N_8688,N_8411,N_8307);
or U8689 (N_8689,N_8495,N_8435);
or U8690 (N_8690,N_8288,N_8304);
nand U8691 (N_8691,N_8419,N_8493);
xnor U8692 (N_8692,N_8397,N_8354);
nor U8693 (N_8693,N_8314,N_8343);
nand U8694 (N_8694,N_8369,N_8452);
xor U8695 (N_8695,N_8271,N_8250);
xor U8696 (N_8696,N_8339,N_8382);
or U8697 (N_8697,N_8442,N_8274);
xnor U8698 (N_8698,N_8292,N_8276);
nand U8699 (N_8699,N_8430,N_8258);
or U8700 (N_8700,N_8287,N_8365);
nand U8701 (N_8701,N_8396,N_8447);
and U8702 (N_8702,N_8310,N_8320);
nand U8703 (N_8703,N_8444,N_8474);
nor U8704 (N_8704,N_8340,N_8463);
nor U8705 (N_8705,N_8321,N_8360);
or U8706 (N_8706,N_8291,N_8455);
and U8707 (N_8707,N_8407,N_8297);
xor U8708 (N_8708,N_8282,N_8400);
or U8709 (N_8709,N_8368,N_8413);
nor U8710 (N_8710,N_8468,N_8322);
xor U8711 (N_8711,N_8402,N_8449);
nand U8712 (N_8712,N_8446,N_8263);
xor U8713 (N_8713,N_8357,N_8487);
nor U8714 (N_8714,N_8344,N_8300);
or U8715 (N_8715,N_8404,N_8450);
nor U8716 (N_8716,N_8406,N_8472);
or U8717 (N_8717,N_8273,N_8285);
nor U8718 (N_8718,N_8449,N_8432);
nand U8719 (N_8719,N_8375,N_8332);
or U8720 (N_8720,N_8257,N_8478);
nor U8721 (N_8721,N_8325,N_8366);
or U8722 (N_8722,N_8357,N_8354);
nand U8723 (N_8723,N_8349,N_8292);
xnor U8724 (N_8724,N_8483,N_8303);
nand U8725 (N_8725,N_8310,N_8255);
or U8726 (N_8726,N_8367,N_8251);
nor U8727 (N_8727,N_8287,N_8430);
nor U8728 (N_8728,N_8430,N_8340);
nand U8729 (N_8729,N_8411,N_8409);
or U8730 (N_8730,N_8275,N_8395);
xor U8731 (N_8731,N_8253,N_8485);
xnor U8732 (N_8732,N_8490,N_8323);
xor U8733 (N_8733,N_8252,N_8484);
xor U8734 (N_8734,N_8306,N_8281);
or U8735 (N_8735,N_8347,N_8482);
xor U8736 (N_8736,N_8468,N_8489);
or U8737 (N_8737,N_8468,N_8482);
or U8738 (N_8738,N_8433,N_8293);
xnor U8739 (N_8739,N_8352,N_8381);
and U8740 (N_8740,N_8299,N_8309);
xor U8741 (N_8741,N_8419,N_8263);
or U8742 (N_8742,N_8320,N_8446);
and U8743 (N_8743,N_8493,N_8400);
nand U8744 (N_8744,N_8312,N_8374);
nand U8745 (N_8745,N_8334,N_8314);
and U8746 (N_8746,N_8261,N_8259);
nor U8747 (N_8747,N_8303,N_8306);
or U8748 (N_8748,N_8262,N_8297);
nand U8749 (N_8749,N_8348,N_8288);
nor U8750 (N_8750,N_8709,N_8612);
nor U8751 (N_8751,N_8615,N_8683);
and U8752 (N_8752,N_8671,N_8562);
and U8753 (N_8753,N_8554,N_8698);
xor U8754 (N_8754,N_8600,N_8670);
nand U8755 (N_8755,N_8694,N_8599);
xnor U8756 (N_8756,N_8542,N_8500);
nand U8757 (N_8757,N_8731,N_8602);
or U8758 (N_8758,N_8588,N_8524);
xnor U8759 (N_8759,N_8652,N_8641);
and U8760 (N_8760,N_8638,N_8665);
or U8761 (N_8761,N_8623,N_8664);
nand U8762 (N_8762,N_8642,N_8536);
xnor U8763 (N_8763,N_8589,N_8501);
and U8764 (N_8764,N_8593,N_8620);
nand U8765 (N_8765,N_8676,N_8630);
nor U8766 (N_8766,N_8617,N_8726);
nand U8767 (N_8767,N_8537,N_8702);
xor U8768 (N_8768,N_8513,N_8648);
and U8769 (N_8769,N_8685,N_8616);
and U8770 (N_8770,N_8658,N_8687);
nand U8771 (N_8771,N_8636,N_8545);
xor U8772 (N_8772,N_8637,N_8523);
nor U8773 (N_8773,N_8696,N_8667);
xnor U8774 (N_8774,N_8669,N_8580);
or U8775 (N_8775,N_8723,N_8565);
or U8776 (N_8776,N_8511,N_8604);
nand U8777 (N_8777,N_8730,N_8732);
or U8778 (N_8778,N_8508,N_8740);
nor U8779 (N_8779,N_8745,N_8681);
or U8780 (N_8780,N_8520,N_8531);
and U8781 (N_8781,N_8635,N_8724);
nor U8782 (N_8782,N_8729,N_8693);
and U8783 (N_8783,N_8690,N_8557);
nor U8784 (N_8784,N_8680,N_8514);
nand U8785 (N_8785,N_8643,N_8556);
nor U8786 (N_8786,N_8522,N_8597);
xnor U8787 (N_8787,N_8647,N_8639);
nand U8788 (N_8788,N_8708,N_8549);
nor U8789 (N_8789,N_8573,N_8572);
or U8790 (N_8790,N_8587,N_8558);
or U8791 (N_8791,N_8733,N_8738);
xnor U8792 (N_8792,N_8575,N_8744);
xnor U8793 (N_8793,N_8674,N_8555);
nor U8794 (N_8794,N_8656,N_8586);
nand U8795 (N_8795,N_8598,N_8735);
or U8796 (N_8796,N_8613,N_8528);
nand U8797 (N_8797,N_8530,N_8649);
nand U8798 (N_8798,N_8594,N_8629);
nor U8799 (N_8799,N_8546,N_8748);
nand U8800 (N_8800,N_8521,N_8715);
nor U8801 (N_8801,N_8653,N_8734);
and U8802 (N_8802,N_8574,N_8736);
and U8803 (N_8803,N_8577,N_8743);
xor U8804 (N_8804,N_8673,N_8532);
nor U8805 (N_8805,N_8699,N_8739);
xnor U8806 (N_8806,N_8644,N_8509);
and U8807 (N_8807,N_8526,N_8675);
or U8808 (N_8808,N_8553,N_8679);
xor U8809 (N_8809,N_8608,N_8607);
nor U8810 (N_8810,N_8678,N_8654);
and U8811 (N_8811,N_8728,N_8579);
xnor U8812 (N_8812,N_8633,N_8512);
or U8813 (N_8813,N_8660,N_8591);
or U8814 (N_8814,N_8716,N_8663);
xnor U8815 (N_8815,N_8567,N_8601);
or U8816 (N_8816,N_8668,N_8645);
nand U8817 (N_8817,N_8606,N_8625);
nand U8818 (N_8818,N_8640,N_8628);
or U8819 (N_8819,N_8703,N_8506);
xnor U8820 (N_8820,N_8560,N_8510);
and U8821 (N_8821,N_8650,N_8627);
or U8822 (N_8822,N_8634,N_8552);
or U8823 (N_8823,N_8610,N_8692);
nor U8824 (N_8824,N_8571,N_8614);
nand U8825 (N_8825,N_8596,N_8540);
nor U8826 (N_8826,N_8700,N_8551);
and U8827 (N_8827,N_8619,N_8541);
or U8828 (N_8828,N_8559,N_8659);
and U8829 (N_8829,N_8618,N_8725);
xor U8830 (N_8830,N_8503,N_8535);
or U8831 (N_8831,N_8543,N_8563);
and U8832 (N_8832,N_8622,N_8583);
and U8833 (N_8833,N_8561,N_8672);
nor U8834 (N_8834,N_8547,N_8718);
xor U8835 (N_8835,N_8646,N_8713);
or U8836 (N_8836,N_8626,N_8706);
nor U8837 (N_8837,N_8651,N_8719);
nor U8838 (N_8838,N_8504,N_8666);
nor U8839 (N_8839,N_8507,N_8689);
or U8840 (N_8840,N_8568,N_8662);
nor U8841 (N_8841,N_8576,N_8564);
xor U8842 (N_8842,N_8595,N_8632);
and U8843 (N_8843,N_8727,N_8722);
or U8844 (N_8844,N_8686,N_8533);
or U8845 (N_8845,N_8684,N_8519);
nor U8846 (N_8846,N_8717,N_8749);
xnor U8847 (N_8847,N_8720,N_8603);
nor U8848 (N_8848,N_8677,N_8621);
nor U8849 (N_8849,N_8582,N_8691);
xor U8850 (N_8850,N_8712,N_8548);
xor U8851 (N_8851,N_8534,N_8611);
xor U8852 (N_8852,N_8516,N_8711);
xor U8853 (N_8853,N_8544,N_8688);
xnor U8854 (N_8854,N_8529,N_8581);
and U8855 (N_8855,N_8742,N_8527);
nand U8856 (N_8856,N_8505,N_8585);
or U8857 (N_8857,N_8747,N_8661);
nor U8858 (N_8858,N_8655,N_8525);
and U8859 (N_8859,N_8746,N_8682);
nand U8860 (N_8860,N_8704,N_8705);
xnor U8861 (N_8861,N_8584,N_8569);
nand U8862 (N_8862,N_8609,N_8697);
or U8863 (N_8863,N_8737,N_8741);
xnor U8864 (N_8864,N_8515,N_8624);
nor U8865 (N_8865,N_8517,N_8570);
nor U8866 (N_8866,N_8714,N_8539);
xor U8867 (N_8867,N_8590,N_8721);
nand U8868 (N_8868,N_8538,N_8518);
xor U8869 (N_8869,N_8502,N_8657);
or U8870 (N_8870,N_8550,N_8707);
nor U8871 (N_8871,N_8605,N_8631);
xor U8872 (N_8872,N_8578,N_8592);
nor U8873 (N_8873,N_8695,N_8701);
and U8874 (N_8874,N_8710,N_8566);
nand U8875 (N_8875,N_8648,N_8714);
nor U8876 (N_8876,N_8565,N_8719);
and U8877 (N_8877,N_8519,N_8630);
nor U8878 (N_8878,N_8610,N_8512);
and U8879 (N_8879,N_8556,N_8658);
and U8880 (N_8880,N_8636,N_8538);
nand U8881 (N_8881,N_8583,N_8686);
nor U8882 (N_8882,N_8624,N_8648);
xnor U8883 (N_8883,N_8523,N_8718);
or U8884 (N_8884,N_8600,N_8678);
nor U8885 (N_8885,N_8720,N_8507);
and U8886 (N_8886,N_8571,N_8633);
nor U8887 (N_8887,N_8556,N_8624);
or U8888 (N_8888,N_8625,N_8543);
nor U8889 (N_8889,N_8608,N_8702);
or U8890 (N_8890,N_8720,N_8508);
nand U8891 (N_8891,N_8689,N_8661);
nor U8892 (N_8892,N_8711,N_8529);
and U8893 (N_8893,N_8638,N_8585);
and U8894 (N_8894,N_8696,N_8505);
or U8895 (N_8895,N_8602,N_8599);
nand U8896 (N_8896,N_8741,N_8691);
nand U8897 (N_8897,N_8632,N_8679);
nand U8898 (N_8898,N_8507,N_8719);
xor U8899 (N_8899,N_8694,N_8653);
nand U8900 (N_8900,N_8741,N_8552);
nand U8901 (N_8901,N_8525,N_8652);
or U8902 (N_8902,N_8727,N_8706);
and U8903 (N_8903,N_8545,N_8598);
nor U8904 (N_8904,N_8552,N_8565);
nor U8905 (N_8905,N_8565,N_8639);
xnor U8906 (N_8906,N_8591,N_8619);
nand U8907 (N_8907,N_8502,N_8709);
nor U8908 (N_8908,N_8505,N_8710);
nor U8909 (N_8909,N_8733,N_8708);
xor U8910 (N_8910,N_8670,N_8514);
nor U8911 (N_8911,N_8620,N_8707);
nand U8912 (N_8912,N_8743,N_8547);
and U8913 (N_8913,N_8519,N_8646);
or U8914 (N_8914,N_8630,N_8597);
or U8915 (N_8915,N_8508,N_8512);
nor U8916 (N_8916,N_8590,N_8503);
xnor U8917 (N_8917,N_8658,N_8549);
and U8918 (N_8918,N_8633,N_8668);
nand U8919 (N_8919,N_8717,N_8677);
and U8920 (N_8920,N_8654,N_8672);
xnor U8921 (N_8921,N_8674,N_8747);
nor U8922 (N_8922,N_8658,N_8713);
nor U8923 (N_8923,N_8554,N_8556);
or U8924 (N_8924,N_8520,N_8590);
or U8925 (N_8925,N_8713,N_8665);
and U8926 (N_8926,N_8539,N_8509);
nor U8927 (N_8927,N_8595,N_8612);
nand U8928 (N_8928,N_8588,N_8600);
xor U8929 (N_8929,N_8714,N_8640);
nor U8930 (N_8930,N_8589,N_8653);
nand U8931 (N_8931,N_8617,N_8561);
and U8932 (N_8932,N_8509,N_8650);
or U8933 (N_8933,N_8545,N_8588);
xnor U8934 (N_8934,N_8695,N_8565);
xor U8935 (N_8935,N_8714,N_8526);
and U8936 (N_8936,N_8596,N_8720);
or U8937 (N_8937,N_8737,N_8534);
or U8938 (N_8938,N_8565,N_8562);
xor U8939 (N_8939,N_8623,N_8713);
nor U8940 (N_8940,N_8688,N_8626);
and U8941 (N_8941,N_8659,N_8542);
nand U8942 (N_8942,N_8731,N_8570);
nor U8943 (N_8943,N_8556,N_8711);
and U8944 (N_8944,N_8639,N_8650);
nor U8945 (N_8945,N_8662,N_8599);
and U8946 (N_8946,N_8520,N_8702);
or U8947 (N_8947,N_8701,N_8673);
nor U8948 (N_8948,N_8681,N_8543);
xnor U8949 (N_8949,N_8541,N_8649);
nand U8950 (N_8950,N_8569,N_8587);
xor U8951 (N_8951,N_8696,N_8690);
xnor U8952 (N_8952,N_8559,N_8614);
or U8953 (N_8953,N_8733,N_8526);
or U8954 (N_8954,N_8714,N_8683);
nand U8955 (N_8955,N_8689,N_8730);
or U8956 (N_8956,N_8541,N_8728);
or U8957 (N_8957,N_8673,N_8629);
and U8958 (N_8958,N_8719,N_8686);
xor U8959 (N_8959,N_8522,N_8589);
nand U8960 (N_8960,N_8508,N_8743);
and U8961 (N_8961,N_8568,N_8542);
and U8962 (N_8962,N_8524,N_8593);
xnor U8963 (N_8963,N_8705,N_8708);
xor U8964 (N_8964,N_8738,N_8616);
xnor U8965 (N_8965,N_8710,N_8629);
and U8966 (N_8966,N_8663,N_8729);
xnor U8967 (N_8967,N_8543,N_8715);
nor U8968 (N_8968,N_8727,N_8607);
xor U8969 (N_8969,N_8565,N_8607);
nor U8970 (N_8970,N_8669,N_8582);
nand U8971 (N_8971,N_8558,N_8690);
or U8972 (N_8972,N_8671,N_8536);
and U8973 (N_8973,N_8634,N_8561);
or U8974 (N_8974,N_8563,N_8654);
and U8975 (N_8975,N_8707,N_8667);
or U8976 (N_8976,N_8638,N_8683);
and U8977 (N_8977,N_8562,N_8532);
and U8978 (N_8978,N_8573,N_8594);
xnor U8979 (N_8979,N_8511,N_8517);
xnor U8980 (N_8980,N_8645,N_8733);
nor U8981 (N_8981,N_8741,N_8528);
or U8982 (N_8982,N_8607,N_8705);
nor U8983 (N_8983,N_8727,N_8505);
or U8984 (N_8984,N_8737,N_8547);
nand U8985 (N_8985,N_8614,N_8629);
or U8986 (N_8986,N_8504,N_8558);
nand U8987 (N_8987,N_8680,N_8663);
and U8988 (N_8988,N_8539,N_8658);
or U8989 (N_8989,N_8547,N_8667);
xor U8990 (N_8990,N_8621,N_8596);
xor U8991 (N_8991,N_8696,N_8590);
xor U8992 (N_8992,N_8636,N_8577);
nor U8993 (N_8993,N_8597,N_8628);
xnor U8994 (N_8994,N_8615,N_8573);
or U8995 (N_8995,N_8546,N_8553);
and U8996 (N_8996,N_8749,N_8673);
or U8997 (N_8997,N_8739,N_8634);
nor U8998 (N_8998,N_8555,N_8597);
nand U8999 (N_8999,N_8721,N_8509);
nand U9000 (N_9000,N_8930,N_8926);
or U9001 (N_9001,N_8750,N_8777);
nand U9002 (N_9002,N_8943,N_8849);
and U9003 (N_9003,N_8969,N_8887);
nand U9004 (N_9004,N_8973,N_8897);
or U9005 (N_9005,N_8902,N_8863);
or U9006 (N_9006,N_8955,N_8964);
nand U9007 (N_9007,N_8835,N_8878);
xor U9008 (N_9008,N_8993,N_8776);
nand U9009 (N_9009,N_8894,N_8946);
nor U9010 (N_9010,N_8971,N_8982);
nor U9011 (N_9011,N_8758,N_8855);
xor U9012 (N_9012,N_8914,N_8960);
nand U9013 (N_9013,N_8788,N_8872);
and U9014 (N_9014,N_8841,N_8954);
xnor U9015 (N_9015,N_8842,N_8761);
nand U9016 (N_9016,N_8765,N_8986);
nand U9017 (N_9017,N_8988,N_8804);
and U9018 (N_9018,N_8965,N_8990);
nand U9019 (N_9019,N_8882,N_8942);
and U9020 (N_9020,N_8826,N_8778);
and U9021 (N_9021,N_8825,N_8931);
and U9022 (N_9022,N_8763,N_8848);
or U9023 (N_9023,N_8814,N_8807);
or U9024 (N_9024,N_8907,N_8769);
nor U9025 (N_9025,N_8781,N_8901);
or U9026 (N_9026,N_8991,N_8757);
nor U9027 (N_9027,N_8854,N_8805);
nor U9028 (N_9028,N_8967,N_8768);
xnor U9029 (N_9029,N_8868,N_8984);
nand U9030 (N_9030,N_8819,N_8839);
or U9031 (N_9031,N_8939,N_8808);
or U9032 (N_9032,N_8767,N_8795);
or U9033 (N_9033,N_8992,N_8922);
or U9034 (N_9034,N_8752,N_8802);
or U9035 (N_9035,N_8941,N_8916);
nand U9036 (N_9036,N_8970,N_8950);
nor U9037 (N_9037,N_8756,N_8856);
xor U9038 (N_9038,N_8785,N_8958);
and U9039 (N_9039,N_8952,N_8925);
or U9040 (N_9040,N_8775,N_8904);
or U9041 (N_9041,N_8770,N_8917);
nor U9042 (N_9042,N_8806,N_8811);
nor U9043 (N_9043,N_8797,N_8838);
nor U9044 (N_9044,N_8751,N_8869);
and U9045 (N_9045,N_8989,N_8885);
and U9046 (N_9046,N_8891,N_8800);
nand U9047 (N_9047,N_8913,N_8799);
or U9048 (N_9048,N_8923,N_8956);
nor U9049 (N_9049,N_8888,N_8821);
nor U9050 (N_9050,N_8772,N_8874);
nor U9051 (N_9051,N_8880,N_8790);
nand U9052 (N_9052,N_8918,N_8812);
nand U9053 (N_9053,N_8972,N_8915);
nand U9054 (N_9054,N_8783,N_8844);
or U9055 (N_9055,N_8822,N_8774);
nor U9056 (N_9056,N_8979,N_8793);
nand U9057 (N_9057,N_8817,N_8895);
or U9058 (N_9058,N_8762,N_8754);
or U9059 (N_9059,N_8779,N_8801);
nand U9060 (N_9060,N_8813,N_8846);
nor U9061 (N_9061,N_8999,N_8810);
xnor U9062 (N_9062,N_8995,N_8843);
nor U9063 (N_9063,N_8794,N_8796);
xnor U9064 (N_9064,N_8908,N_8924);
xnor U9065 (N_9065,N_8829,N_8851);
nand U9066 (N_9066,N_8753,N_8833);
nand U9067 (N_9067,N_8875,N_8938);
nor U9068 (N_9068,N_8823,N_8879);
or U9069 (N_9069,N_8935,N_8909);
or U9070 (N_9070,N_8962,N_8905);
and U9071 (N_9071,N_8830,N_8929);
and U9072 (N_9072,N_8867,N_8919);
and U9073 (N_9073,N_8974,N_8959);
or U9074 (N_9074,N_8877,N_8850);
xor U9075 (N_9075,N_8866,N_8957);
nor U9076 (N_9076,N_8994,N_8889);
and U9077 (N_9077,N_8865,N_8784);
nand U9078 (N_9078,N_8847,N_8996);
or U9079 (N_9079,N_8820,N_8983);
nand U9080 (N_9080,N_8827,N_8859);
nand U9081 (N_9081,N_8951,N_8818);
xor U9082 (N_9082,N_8831,N_8906);
and U9083 (N_9083,N_8928,N_8755);
xor U9084 (N_9084,N_8899,N_8787);
nor U9085 (N_9085,N_8764,N_8968);
and U9086 (N_9086,N_8857,N_8864);
nand U9087 (N_9087,N_8760,N_8873);
xnor U9088 (N_9088,N_8832,N_8886);
and U9089 (N_9089,N_8900,N_8860);
nor U9090 (N_9090,N_8798,N_8976);
xnor U9091 (N_9091,N_8948,N_8828);
nor U9092 (N_9092,N_8903,N_8816);
or U9093 (N_9093,N_8871,N_8949);
or U9094 (N_9094,N_8786,N_8858);
nor U9095 (N_9095,N_8981,N_8963);
nand U9096 (N_9096,N_8883,N_8920);
nor U9097 (N_9097,N_8782,N_8980);
nor U9098 (N_9098,N_8791,N_8853);
nand U9099 (N_9099,N_8884,N_8766);
xnor U9100 (N_9100,N_8947,N_8940);
or U9101 (N_9101,N_8932,N_8927);
nand U9102 (N_9102,N_8966,N_8896);
and U9103 (N_9103,N_8840,N_8862);
nand U9104 (N_9104,N_8945,N_8921);
or U9105 (N_9105,N_8834,N_8861);
xor U9106 (N_9106,N_8845,N_8944);
nor U9107 (N_9107,N_8997,N_8870);
or U9108 (N_9108,N_8898,N_8934);
xnor U9109 (N_9109,N_8910,N_8809);
or U9110 (N_9110,N_8893,N_8837);
nand U9111 (N_9111,N_8824,N_8937);
nand U9112 (N_9112,N_8876,N_8836);
or U9113 (N_9113,N_8977,N_8985);
or U9114 (N_9114,N_8890,N_8987);
or U9115 (N_9115,N_8998,N_8789);
and U9116 (N_9116,N_8852,N_8771);
nand U9117 (N_9117,N_8912,N_8933);
and U9118 (N_9118,N_8881,N_8936);
or U9119 (N_9119,N_8911,N_8975);
nand U9120 (N_9120,N_8803,N_8978);
and U9121 (N_9121,N_8953,N_8780);
or U9122 (N_9122,N_8773,N_8792);
xor U9123 (N_9123,N_8759,N_8892);
nor U9124 (N_9124,N_8961,N_8815);
nand U9125 (N_9125,N_8829,N_8926);
nor U9126 (N_9126,N_8947,N_8846);
nand U9127 (N_9127,N_8818,N_8851);
xor U9128 (N_9128,N_8898,N_8857);
nand U9129 (N_9129,N_8905,N_8840);
xor U9130 (N_9130,N_8815,N_8861);
xnor U9131 (N_9131,N_8963,N_8927);
nand U9132 (N_9132,N_8968,N_8794);
xnor U9133 (N_9133,N_8781,N_8758);
nor U9134 (N_9134,N_8785,N_8888);
nand U9135 (N_9135,N_8810,N_8831);
and U9136 (N_9136,N_8904,N_8982);
xor U9137 (N_9137,N_8893,N_8866);
or U9138 (N_9138,N_8813,N_8872);
nor U9139 (N_9139,N_8964,N_8992);
nand U9140 (N_9140,N_8863,N_8878);
or U9141 (N_9141,N_8976,N_8842);
nand U9142 (N_9142,N_8897,N_8833);
nand U9143 (N_9143,N_8846,N_8852);
or U9144 (N_9144,N_8766,N_8850);
xor U9145 (N_9145,N_8803,N_8991);
nor U9146 (N_9146,N_8767,N_8959);
or U9147 (N_9147,N_8864,N_8964);
and U9148 (N_9148,N_8849,N_8751);
and U9149 (N_9149,N_8902,N_8775);
or U9150 (N_9150,N_8877,N_8786);
or U9151 (N_9151,N_8808,N_8819);
nand U9152 (N_9152,N_8767,N_8766);
and U9153 (N_9153,N_8772,N_8935);
xor U9154 (N_9154,N_8875,N_8760);
xnor U9155 (N_9155,N_8780,N_8753);
nand U9156 (N_9156,N_8776,N_8822);
nand U9157 (N_9157,N_8831,N_8757);
or U9158 (N_9158,N_8900,N_8807);
nand U9159 (N_9159,N_8948,N_8856);
nand U9160 (N_9160,N_8879,N_8884);
and U9161 (N_9161,N_8786,N_8935);
nand U9162 (N_9162,N_8891,N_8921);
xor U9163 (N_9163,N_8892,N_8970);
and U9164 (N_9164,N_8925,N_8943);
nand U9165 (N_9165,N_8760,N_8850);
or U9166 (N_9166,N_8899,N_8879);
and U9167 (N_9167,N_8767,N_8802);
xor U9168 (N_9168,N_8810,N_8834);
or U9169 (N_9169,N_8841,N_8996);
nor U9170 (N_9170,N_8955,N_8913);
nor U9171 (N_9171,N_8941,N_8808);
xnor U9172 (N_9172,N_8847,N_8938);
or U9173 (N_9173,N_8929,N_8888);
and U9174 (N_9174,N_8864,N_8815);
nand U9175 (N_9175,N_8957,N_8770);
nand U9176 (N_9176,N_8811,N_8922);
xor U9177 (N_9177,N_8921,N_8885);
xor U9178 (N_9178,N_8813,N_8818);
or U9179 (N_9179,N_8922,N_8993);
or U9180 (N_9180,N_8955,N_8872);
nor U9181 (N_9181,N_8884,N_8750);
nor U9182 (N_9182,N_8843,N_8784);
xor U9183 (N_9183,N_8837,N_8801);
nand U9184 (N_9184,N_8792,N_8767);
or U9185 (N_9185,N_8851,N_8833);
and U9186 (N_9186,N_8939,N_8962);
xnor U9187 (N_9187,N_8818,N_8819);
nor U9188 (N_9188,N_8971,N_8939);
nor U9189 (N_9189,N_8797,N_8927);
and U9190 (N_9190,N_8864,N_8853);
nand U9191 (N_9191,N_8901,N_8974);
nor U9192 (N_9192,N_8965,N_8930);
nand U9193 (N_9193,N_8770,N_8796);
or U9194 (N_9194,N_8963,N_8766);
xnor U9195 (N_9195,N_8971,N_8870);
nand U9196 (N_9196,N_8876,N_8916);
and U9197 (N_9197,N_8906,N_8756);
xor U9198 (N_9198,N_8853,N_8996);
xnor U9199 (N_9199,N_8950,N_8797);
nor U9200 (N_9200,N_8903,N_8958);
nand U9201 (N_9201,N_8920,N_8809);
and U9202 (N_9202,N_8961,N_8757);
and U9203 (N_9203,N_8845,N_8884);
or U9204 (N_9204,N_8999,N_8808);
nor U9205 (N_9205,N_8805,N_8756);
nor U9206 (N_9206,N_8990,N_8906);
or U9207 (N_9207,N_8886,N_8995);
nand U9208 (N_9208,N_8755,N_8776);
xnor U9209 (N_9209,N_8798,N_8928);
or U9210 (N_9210,N_8991,N_8945);
xnor U9211 (N_9211,N_8937,N_8997);
or U9212 (N_9212,N_8978,N_8944);
xor U9213 (N_9213,N_8984,N_8845);
or U9214 (N_9214,N_8892,N_8962);
or U9215 (N_9215,N_8788,N_8889);
or U9216 (N_9216,N_8921,N_8983);
and U9217 (N_9217,N_8923,N_8855);
nand U9218 (N_9218,N_8908,N_8752);
and U9219 (N_9219,N_8863,N_8875);
xor U9220 (N_9220,N_8906,N_8752);
xnor U9221 (N_9221,N_8780,N_8826);
and U9222 (N_9222,N_8792,N_8764);
and U9223 (N_9223,N_8886,N_8981);
xnor U9224 (N_9224,N_8905,N_8765);
xnor U9225 (N_9225,N_8866,N_8916);
xnor U9226 (N_9226,N_8761,N_8874);
nor U9227 (N_9227,N_8797,N_8973);
or U9228 (N_9228,N_8992,N_8779);
nand U9229 (N_9229,N_8863,N_8793);
nand U9230 (N_9230,N_8870,N_8831);
or U9231 (N_9231,N_8767,N_8883);
nor U9232 (N_9232,N_8954,N_8915);
or U9233 (N_9233,N_8765,N_8938);
xnor U9234 (N_9234,N_8777,N_8901);
xor U9235 (N_9235,N_8822,N_8836);
xor U9236 (N_9236,N_8967,N_8830);
nor U9237 (N_9237,N_8801,N_8764);
nand U9238 (N_9238,N_8806,N_8857);
xor U9239 (N_9239,N_8765,N_8755);
or U9240 (N_9240,N_8773,N_8756);
or U9241 (N_9241,N_8790,N_8765);
xnor U9242 (N_9242,N_8804,N_8946);
nor U9243 (N_9243,N_8787,N_8867);
nor U9244 (N_9244,N_8762,N_8766);
and U9245 (N_9245,N_8860,N_8889);
xor U9246 (N_9246,N_8951,N_8907);
nor U9247 (N_9247,N_8760,N_8938);
and U9248 (N_9248,N_8814,N_8977);
xor U9249 (N_9249,N_8901,N_8869);
or U9250 (N_9250,N_9174,N_9157);
xor U9251 (N_9251,N_9228,N_9035);
xor U9252 (N_9252,N_9217,N_9224);
xnor U9253 (N_9253,N_9072,N_9191);
and U9254 (N_9254,N_9088,N_9207);
nor U9255 (N_9255,N_9069,N_9091);
xor U9256 (N_9256,N_9179,N_9019);
and U9257 (N_9257,N_9182,N_9189);
or U9258 (N_9258,N_9233,N_9194);
xor U9259 (N_9259,N_9083,N_9203);
nor U9260 (N_9260,N_9075,N_9043);
nor U9261 (N_9261,N_9108,N_9038);
nor U9262 (N_9262,N_9080,N_9167);
or U9263 (N_9263,N_9138,N_9246);
and U9264 (N_9264,N_9085,N_9014);
xnor U9265 (N_9265,N_9172,N_9020);
nor U9266 (N_9266,N_9219,N_9016);
or U9267 (N_9267,N_9052,N_9081);
xnor U9268 (N_9268,N_9047,N_9235);
nand U9269 (N_9269,N_9158,N_9036);
and U9270 (N_9270,N_9198,N_9055);
or U9271 (N_9271,N_9141,N_9037);
and U9272 (N_9272,N_9197,N_9031);
nor U9273 (N_9273,N_9238,N_9153);
xnor U9274 (N_9274,N_9135,N_9044);
or U9275 (N_9275,N_9146,N_9236);
xnor U9276 (N_9276,N_9165,N_9160);
or U9277 (N_9277,N_9053,N_9034);
nand U9278 (N_9278,N_9022,N_9032);
nand U9279 (N_9279,N_9005,N_9173);
xnor U9280 (N_9280,N_9000,N_9121);
or U9281 (N_9281,N_9216,N_9008);
nand U9282 (N_9282,N_9161,N_9186);
xor U9283 (N_9283,N_9087,N_9248);
or U9284 (N_9284,N_9015,N_9009);
nor U9285 (N_9285,N_9247,N_9188);
xnor U9286 (N_9286,N_9006,N_9245);
or U9287 (N_9287,N_9195,N_9115);
and U9288 (N_9288,N_9120,N_9028);
nand U9289 (N_9289,N_9192,N_9097);
or U9290 (N_9290,N_9017,N_9106);
nor U9291 (N_9291,N_9113,N_9090);
nor U9292 (N_9292,N_9159,N_9098);
nand U9293 (N_9293,N_9112,N_9012);
nand U9294 (N_9294,N_9078,N_9229);
nor U9295 (N_9295,N_9070,N_9241);
nand U9296 (N_9296,N_9211,N_9045);
nand U9297 (N_9297,N_9209,N_9025);
nor U9298 (N_9298,N_9249,N_9059);
and U9299 (N_9299,N_9007,N_9178);
xnor U9300 (N_9300,N_9024,N_9027);
nor U9301 (N_9301,N_9201,N_9134);
or U9302 (N_9302,N_9234,N_9122);
nor U9303 (N_9303,N_9086,N_9154);
nand U9304 (N_9304,N_9130,N_9230);
and U9305 (N_9305,N_9058,N_9004);
and U9306 (N_9306,N_9033,N_9125);
or U9307 (N_9307,N_9049,N_9118);
xor U9308 (N_9308,N_9223,N_9114);
or U9309 (N_9309,N_9119,N_9079);
or U9310 (N_9310,N_9185,N_9151);
and U9311 (N_9311,N_9076,N_9101);
and U9312 (N_9312,N_9023,N_9102);
xnor U9313 (N_9313,N_9239,N_9042);
and U9314 (N_9314,N_9140,N_9066);
nor U9315 (N_9315,N_9084,N_9218);
nand U9316 (N_9316,N_9123,N_9104);
xnor U9317 (N_9317,N_9061,N_9215);
nor U9318 (N_9318,N_9107,N_9171);
nor U9319 (N_9319,N_9155,N_9176);
and U9320 (N_9320,N_9202,N_9082);
nand U9321 (N_9321,N_9030,N_9149);
and U9322 (N_9322,N_9204,N_9210);
nor U9323 (N_9323,N_9213,N_9221);
or U9324 (N_9324,N_9063,N_9060);
nand U9325 (N_9325,N_9109,N_9093);
xnor U9326 (N_9326,N_9242,N_9150);
nand U9327 (N_9327,N_9029,N_9089);
nand U9328 (N_9328,N_9205,N_9222);
or U9329 (N_9329,N_9162,N_9099);
and U9330 (N_9330,N_9244,N_9183);
nand U9331 (N_9331,N_9056,N_9240);
nor U9332 (N_9332,N_9065,N_9147);
xnor U9333 (N_9333,N_9111,N_9184);
xor U9334 (N_9334,N_9095,N_9116);
nor U9335 (N_9335,N_9011,N_9040);
xor U9336 (N_9336,N_9021,N_9094);
nand U9337 (N_9337,N_9026,N_9139);
or U9338 (N_9338,N_9187,N_9190);
xnor U9339 (N_9339,N_9067,N_9226);
or U9340 (N_9340,N_9133,N_9092);
or U9341 (N_9341,N_9227,N_9010);
nor U9342 (N_9342,N_9193,N_9220);
nand U9343 (N_9343,N_9144,N_9152);
or U9344 (N_9344,N_9145,N_9050);
nor U9345 (N_9345,N_9142,N_9206);
or U9346 (N_9346,N_9175,N_9051);
nor U9347 (N_9347,N_9166,N_9117);
nand U9348 (N_9348,N_9127,N_9143);
nor U9349 (N_9349,N_9100,N_9199);
xor U9350 (N_9350,N_9105,N_9163);
and U9351 (N_9351,N_9137,N_9148);
nor U9352 (N_9352,N_9181,N_9126);
or U9353 (N_9353,N_9243,N_9013);
and U9354 (N_9354,N_9074,N_9168);
nor U9355 (N_9355,N_9073,N_9136);
or U9356 (N_9356,N_9156,N_9231);
nor U9357 (N_9357,N_9039,N_9212);
nor U9358 (N_9358,N_9048,N_9071);
nand U9359 (N_9359,N_9068,N_9164);
nor U9360 (N_9360,N_9103,N_9132);
or U9361 (N_9361,N_9170,N_9128);
nor U9362 (N_9362,N_9196,N_9131);
nand U9363 (N_9363,N_9180,N_9208);
or U9364 (N_9364,N_9110,N_9003);
and U9365 (N_9365,N_9057,N_9018);
or U9366 (N_9366,N_9001,N_9002);
and U9367 (N_9367,N_9124,N_9096);
nor U9368 (N_9368,N_9062,N_9054);
nand U9369 (N_9369,N_9237,N_9225);
or U9370 (N_9370,N_9129,N_9232);
nand U9371 (N_9371,N_9077,N_9064);
and U9372 (N_9372,N_9200,N_9177);
nand U9373 (N_9373,N_9214,N_9041);
nor U9374 (N_9374,N_9169,N_9046);
nor U9375 (N_9375,N_9068,N_9043);
nor U9376 (N_9376,N_9000,N_9031);
and U9377 (N_9377,N_9038,N_9033);
nor U9378 (N_9378,N_9124,N_9121);
nor U9379 (N_9379,N_9057,N_9166);
or U9380 (N_9380,N_9195,N_9055);
or U9381 (N_9381,N_9020,N_9106);
nand U9382 (N_9382,N_9081,N_9237);
nor U9383 (N_9383,N_9187,N_9058);
nor U9384 (N_9384,N_9233,N_9147);
or U9385 (N_9385,N_9048,N_9110);
nor U9386 (N_9386,N_9150,N_9081);
or U9387 (N_9387,N_9187,N_9159);
or U9388 (N_9388,N_9075,N_9169);
and U9389 (N_9389,N_9015,N_9213);
nor U9390 (N_9390,N_9242,N_9235);
nand U9391 (N_9391,N_9110,N_9072);
or U9392 (N_9392,N_9084,N_9188);
nand U9393 (N_9393,N_9023,N_9219);
or U9394 (N_9394,N_9236,N_9220);
nor U9395 (N_9395,N_9121,N_9022);
nor U9396 (N_9396,N_9086,N_9024);
and U9397 (N_9397,N_9101,N_9005);
or U9398 (N_9398,N_9213,N_9193);
or U9399 (N_9399,N_9051,N_9115);
xor U9400 (N_9400,N_9177,N_9166);
nand U9401 (N_9401,N_9093,N_9203);
xor U9402 (N_9402,N_9073,N_9122);
nand U9403 (N_9403,N_9063,N_9080);
or U9404 (N_9404,N_9225,N_9015);
nand U9405 (N_9405,N_9060,N_9218);
or U9406 (N_9406,N_9130,N_9194);
or U9407 (N_9407,N_9049,N_9225);
or U9408 (N_9408,N_9144,N_9233);
and U9409 (N_9409,N_9162,N_9234);
nand U9410 (N_9410,N_9138,N_9170);
nand U9411 (N_9411,N_9023,N_9029);
and U9412 (N_9412,N_9189,N_9055);
xor U9413 (N_9413,N_9155,N_9211);
xnor U9414 (N_9414,N_9049,N_9221);
nand U9415 (N_9415,N_9006,N_9126);
and U9416 (N_9416,N_9060,N_9224);
xor U9417 (N_9417,N_9179,N_9045);
nand U9418 (N_9418,N_9096,N_9095);
nor U9419 (N_9419,N_9223,N_9037);
nor U9420 (N_9420,N_9068,N_9087);
or U9421 (N_9421,N_9136,N_9113);
or U9422 (N_9422,N_9239,N_9084);
nand U9423 (N_9423,N_9175,N_9189);
and U9424 (N_9424,N_9148,N_9044);
nor U9425 (N_9425,N_9234,N_9064);
and U9426 (N_9426,N_9166,N_9157);
or U9427 (N_9427,N_9011,N_9172);
and U9428 (N_9428,N_9020,N_9080);
or U9429 (N_9429,N_9240,N_9204);
and U9430 (N_9430,N_9193,N_9020);
xor U9431 (N_9431,N_9103,N_9236);
nor U9432 (N_9432,N_9230,N_9041);
nor U9433 (N_9433,N_9131,N_9160);
and U9434 (N_9434,N_9085,N_9106);
or U9435 (N_9435,N_9015,N_9140);
and U9436 (N_9436,N_9112,N_9167);
or U9437 (N_9437,N_9106,N_9054);
or U9438 (N_9438,N_9138,N_9189);
nand U9439 (N_9439,N_9133,N_9216);
xnor U9440 (N_9440,N_9041,N_9004);
and U9441 (N_9441,N_9241,N_9194);
xor U9442 (N_9442,N_9111,N_9035);
or U9443 (N_9443,N_9050,N_9169);
and U9444 (N_9444,N_9072,N_9106);
and U9445 (N_9445,N_9006,N_9124);
xor U9446 (N_9446,N_9219,N_9220);
nand U9447 (N_9447,N_9192,N_9161);
and U9448 (N_9448,N_9202,N_9111);
nor U9449 (N_9449,N_9108,N_9225);
and U9450 (N_9450,N_9217,N_9116);
nand U9451 (N_9451,N_9082,N_9186);
xnor U9452 (N_9452,N_9234,N_9097);
nand U9453 (N_9453,N_9082,N_9172);
and U9454 (N_9454,N_9008,N_9075);
nor U9455 (N_9455,N_9199,N_9214);
xnor U9456 (N_9456,N_9049,N_9047);
and U9457 (N_9457,N_9194,N_9196);
nand U9458 (N_9458,N_9017,N_9232);
xnor U9459 (N_9459,N_9078,N_9005);
or U9460 (N_9460,N_9170,N_9132);
nor U9461 (N_9461,N_9044,N_9189);
nor U9462 (N_9462,N_9100,N_9122);
xnor U9463 (N_9463,N_9098,N_9237);
xor U9464 (N_9464,N_9090,N_9183);
or U9465 (N_9465,N_9032,N_9171);
nand U9466 (N_9466,N_9090,N_9043);
nor U9467 (N_9467,N_9237,N_9091);
nand U9468 (N_9468,N_9117,N_9223);
and U9469 (N_9469,N_9065,N_9088);
and U9470 (N_9470,N_9234,N_9130);
and U9471 (N_9471,N_9166,N_9054);
xnor U9472 (N_9472,N_9011,N_9042);
nor U9473 (N_9473,N_9179,N_9155);
nand U9474 (N_9474,N_9013,N_9233);
and U9475 (N_9475,N_9245,N_9097);
or U9476 (N_9476,N_9169,N_9170);
and U9477 (N_9477,N_9229,N_9242);
nand U9478 (N_9478,N_9037,N_9111);
nand U9479 (N_9479,N_9161,N_9053);
and U9480 (N_9480,N_9094,N_9231);
nor U9481 (N_9481,N_9019,N_9033);
xor U9482 (N_9482,N_9019,N_9185);
nand U9483 (N_9483,N_9007,N_9213);
and U9484 (N_9484,N_9247,N_9021);
xnor U9485 (N_9485,N_9214,N_9115);
or U9486 (N_9486,N_9101,N_9159);
nor U9487 (N_9487,N_9055,N_9178);
and U9488 (N_9488,N_9104,N_9226);
or U9489 (N_9489,N_9034,N_9128);
or U9490 (N_9490,N_9210,N_9125);
nand U9491 (N_9491,N_9103,N_9155);
or U9492 (N_9492,N_9096,N_9109);
nor U9493 (N_9493,N_9056,N_9101);
and U9494 (N_9494,N_9100,N_9242);
and U9495 (N_9495,N_9053,N_9043);
nor U9496 (N_9496,N_9242,N_9044);
xnor U9497 (N_9497,N_9171,N_9025);
or U9498 (N_9498,N_9229,N_9073);
xnor U9499 (N_9499,N_9169,N_9137);
nor U9500 (N_9500,N_9411,N_9437);
nand U9501 (N_9501,N_9396,N_9265);
and U9502 (N_9502,N_9412,N_9467);
nor U9503 (N_9503,N_9340,N_9284);
xnor U9504 (N_9504,N_9408,N_9471);
xnor U9505 (N_9505,N_9404,N_9489);
or U9506 (N_9506,N_9370,N_9261);
nand U9507 (N_9507,N_9497,N_9345);
xor U9508 (N_9508,N_9277,N_9323);
or U9509 (N_9509,N_9273,N_9400);
and U9510 (N_9510,N_9389,N_9348);
nand U9511 (N_9511,N_9254,N_9440);
or U9512 (N_9512,N_9468,N_9259);
nor U9513 (N_9513,N_9304,N_9379);
or U9514 (N_9514,N_9260,N_9496);
nor U9515 (N_9515,N_9485,N_9465);
nand U9516 (N_9516,N_9448,N_9495);
and U9517 (N_9517,N_9391,N_9354);
or U9518 (N_9518,N_9449,N_9480);
or U9519 (N_9519,N_9403,N_9319);
xnor U9520 (N_9520,N_9463,N_9452);
or U9521 (N_9521,N_9294,N_9472);
xor U9522 (N_9522,N_9331,N_9338);
xor U9523 (N_9523,N_9470,N_9446);
or U9524 (N_9524,N_9336,N_9368);
nor U9525 (N_9525,N_9315,N_9325);
and U9526 (N_9526,N_9482,N_9416);
xnor U9527 (N_9527,N_9267,N_9447);
nand U9528 (N_9528,N_9382,N_9387);
and U9529 (N_9529,N_9414,N_9381);
and U9530 (N_9530,N_9364,N_9429);
xnor U9531 (N_9531,N_9433,N_9327);
nor U9532 (N_9532,N_9291,N_9475);
and U9533 (N_9533,N_9314,N_9450);
nand U9534 (N_9534,N_9431,N_9349);
xnor U9535 (N_9535,N_9380,N_9445);
nor U9536 (N_9536,N_9322,N_9316);
and U9537 (N_9537,N_9324,N_9295);
and U9538 (N_9538,N_9286,N_9378);
nand U9539 (N_9539,N_9312,N_9410);
or U9540 (N_9540,N_9306,N_9406);
nor U9541 (N_9541,N_9462,N_9283);
and U9542 (N_9542,N_9432,N_9487);
and U9543 (N_9543,N_9441,N_9385);
or U9544 (N_9544,N_9330,N_9430);
nand U9545 (N_9545,N_9363,N_9255);
xnor U9546 (N_9546,N_9442,N_9320);
or U9547 (N_9547,N_9454,N_9332);
or U9548 (N_9548,N_9456,N_9317);
xnor U9549 (N_9549,N_9374,N_9444);
xor U9550 (N_9550,N_9402,N_9268);
nand U9551 (N_9551,N_9401,N_9460);
nand U9552 (N_9552,N_9303,N_9490);
xnor U9553 (N_9553,N_9399,N_9419);
and U9554 (N_9554,N_9455,N_9326);
nor U9555 (N_9555,N_9285,N_9308);
nor U9556 (N_9556,N_9427,N_9371);
or U9557 (N_9557,N_9494,N_9421);
nor U9558 (N_9558,N_9499,N_9328);
nand U9559 (N_9559,N_9409,N_9388);
nand U9560 (N_9560,N_9334,N_9453);
and U9561 (N_9561,N_9392,N_9293);
nand U9562 (N_9562,N_9300,N_9253);
nor U9563 (N_9563,N_9281,N_9266);
or U9564 (N_9564,N_9282,N_9358);
nor U9565 (N_9565,N_9257,N_9420);
and U9566 (N_9566,N_9461,N_9376);
and U9567 (N_9567,N_9263,N_9434);
nand U9568 (N_9568,N_9279,N_9262);
xnor U9569 (N_9569,N_9313,N_9436);
xnor U9570 (N_9570,N_9466,N_9426);
nand U9571 (N_9571,N_9302,N_9366);
nand U9572 (N_9572,N_9483,N_9318);
or U9573 (N_9573,N_9258,N_9439);
xnor U9574 (N_9574,N_9407,N_9476);
nor U9575 (N_9575,N_9251,N_9435);
and U9576 (N_9576,N_9355,N_9360);
nand U9577 (N_9577,N_9367,N_9464);
nor U9578 (N_9578,N_9390,N_9393);
and U9579 (N_9579,N_9275,N_9350);
or U9580 (N_9580,N_9491,N_9335);
xor U9581 (N_9581,N_9305,N_9369);
or U9582 (N_9582,N_9469,N_9484);
nand U9583 (N_9583,N_9428,N_9457);
nor U9584 (N_9584,N_9290,N_9337);
xnor U9585 (N_9585,N_9280,N_9347);
and U9586 (N_9586,N_9352,N_9375);
nor U9587 (N_9587,N_9359,N_9343);
or U9588 (N_9588,N_9289,N_9270);
or U9589 (N_9589,N_9271,N_9288);
or U9590 (N_9590,N_9373,N_9297);
or U9591 (N_9591,N_9477,N_9362);
or U9592 (N_9592,N_9310,N_9473);
nand U9593 (N_9593,N_9397,N_9311);
nor U9594 (N_9594,N_9346,N_9321);
or U9595 (N_9595,N_9492,N_9413);
nor U9596 (N_9596,N_9274,N_9478);
or U9597 (N_9597,N_9341,N_9398);
xor U9598 (N_9598,N_9386,N_9342);
xnor U9599 (N_9599,N_9339,N_9301);
nor U9600 (N_9600,N_9353,N_9451);
nand U9601 (N_9601,N_9383,N_9493);
or U9602 (N_9602,N_9299,N_9479);
or U9603 (N_9603,N_9309,N_9298);
nand U9604 (N_9604,N_9423,N_9372);
and U9605 (N_9605,N_9272,N_9264);
nor U9606 (N_9606,N_9438,N_9422);
nand U9607 (N_9607,N_9292,N_9252);
xnor U9608 (N_9608,N_9361,N_9256);
xnor U9609 (N_9609,N_9351,N_9329);
nor U9610 (N_9610,N_9356,N_9394);
nor U9611 (N_9611,N_9486,N_9417);
and U9612 (N_9612,N_9287,N_9384);
or U9613 (N_9613,N_9395,N_9269);
nor U9614 (N_9614,N_9296,N_9307);
xnor U9615 (N_9615,N_9415,N_9250);
xnor U9616 (N_9616,N_9425,N_9344);
nor U9617 (N_9617,N_9333,N_9377);
nor U9618 (N_9618,N_9357,N_9278);
nor U9619 (N_9619,N_9405,N_9443);
nand U9620 (N_9620,N_9418,N_9481);
xor U9621 (N_9621,N_9488,N_9458);
nand U9622 (N_9622,N_9498,N_9365);
nor U9623 (N_9623,N_9459,N_9424);
or U9624 (N_9624,N_9276,N_9474);
nor U9625 (N_9625,N_9452,N_9432);
and U9626 (N_9626,N_9258,N_9255);
and U9627 (N_9627,N_9371,N_9455);
or U9628 (N_9628,N_9416,N_9250);
nor U9629 (N_9629,N_9425,N_9392);
or U9630 (N_9630,N_9331,N_9339);
nor U9631 (N_9631,N_9396,N_9373);
nor U9632 (N_9632,N_9445,N_9319);
and U9633 (N_9633,N_9490,N_9344);
xnor U9634 (N_9634,N_9410,N_9278);
xor U9635 (N_9635,N_9444,N_9251);
and U9636 (N_9636,N_9250,N_9322);
nand U9637 (N_9637,N_9425,N_9428);
xnor U9638 (N_9638,N_9478,N_9467);
or U9639 (N_9639,N_9409,N_9436);
xnor U9640 (N_9640,N_9349,N_9328);
nor U9641 (N_9641,N_9416,N_9272);
or U9642 (N_9642,N_9390,N_9299);
and U9643 (N_9643,N_9313,N_9418);
xnor U9644 (N_9644,N_9252,N_9290);
and U9645 (N_9645,N_9286,N_9250);
or U9646 (N_9646,N_9457,N_9447);
nor U9647 (N_9647,N_9340,N_9303);
nor U9648 (N_9648,N_9370,N_9411);
nand U9649 (N_9649,N_9324,N_9338);
or U9650 (N_9650,N_9361,N_9309);
xor U9651 (N_9651,N_9295,N_9300);
and U9652 (N_9652,N_9298,N_9464);
nand U9653 (N_9653,N_9255,N_9372);
or U9654 (N_9654,N_9402,N_9406);
xor U9655 (N_9655,N_9313,N_9364);
xnor U9656 (N_9656,N_9321,N_9286);
xnor U9657 (N_9657,N_9325,N_9303);
nor U9658 (N_9658,N_9288,N_9289);
and U9659 (N_9659,N_9259,N_9363);
xnor U9660 (N_9660,N_9348,N_9346);
and U9661 (N_9661,N_9443,N_9415);
nor U9662 (N_9662,N_9327,N_9406);
and U9663 (N_9663,N_9331,N_9399);
or U9664 (N_9664,N_9281,N_9325);
nor U9665 (N_9665,N_9467,N_9491);
nand U9666 (N_9666,N_9268,N_9333);
xnor U9667 (N_9667,N_9490,N_9453);
xor U9668 (N_9668,N_9333,N_9387);
or U9669 (N_9669,N_9428,N_9365);
nand U9670 (N_9670,N_9478,N_9286);
nand U9671 (N_9671,N_9424,N_9289);
xor U9672 (N_9672,N_9416,N_9268);
and U9673 (N_9673,N_9468,N_9268);
or U9674 (N_9674,N_9405,N_9419);
xnor U9675 (N_9675,N_9460,N_9421);
or U9676 (N_9676,N_9361,N_9253);
or U9677 (N_9677,N_9468,N_9457);
and U9678 (N_9678,N_9448,N_9315);
nor U9679 (N_9679,N_9261,N_9293);
xnor U9680 (N_9680,N_9269,N_9250);
nor U9681 (N_9681,N_9303,N_9262);
or U9682 (N_9682,N_9434,N_9428);
nor U9683 (N_9683,N_9255,N_9348);
nor U9684 (N_9684,N_9329,N_9397);
or U9685 (N_9685,N_9349,N_9293);
xor U9686 (N_9686,N_9485,N_9337);
xnor U9687 (N_9687,N_9488,N_9418);
or U9688 (N_9688,N_9310,N_9439);
or U9689 (N_9689,N_9373,N_9345);
nand U9690 (N_9690,N_9387,N_9378);
and U9691 (N_9691,N_9449,N_9286);
nor U9692 (N_9692,N_9361,N_9294);
xnor U9693 (N_9693,N_9412,N_9354);
and U9694 (N_9694,N_9314,N_9466);
nor U9695 (N_9695,N_9446,N_9442);
nand U9696 (N_9696,N_9352,N_9412);
xor U9697 (N_9697,N_9471,N_9383);
and U9698 (N_9698,N_9323,N_9442);
and U9699 (N_9699,N_9416,N_9274);
and U9700 (N_9700,N_9334,N_9326);
nand U9701 (N_9701,N_9311,N_9262);
or U9702 (N_9702,N_9291,N_9396);
and U9703 (N_9703,N_9279,N_9422);
xor U9704 (N_9704,N_9311,N_9359);
or U9705 (N_9705,N_9375,N_9278);
and U9706 (N_9706,N_9347,N_9323);
and U9707 (N_9707,N_9419,N_9288);
nand U9708 (N_9708,N_9446,N_9347);
nand U9709 (N_9709,N_9264,N_9406);
xnor U9710 (N_9710,N_9347,N_9295);
and U9711 (N_9711,N_9459,N_9250);
xnor U9712 (N_9712,N_9272,N_9456);
or U9713 (N_9713,N_9368,N_9457);
nor U9714 (N_9714,N_9457,N_9291);
nor U9715 (N_9715,N_9338,N_9406);
or U9716 (N_9716,N_9294,N_9436);
or U9717 (N_9717,N_9251,N_9427);
nor U9718 (N_9718,N_9327,N_9330);
and U9719 (N_9719,N_9286,N_9465);
nand U9720 (N_9720,N_9446,N_9450);
xnor U9721 (N_9721,N_9420,N_9380);
and U9722 (N_9722,N_9429,N_9325);
nand U9723 (N_9723,N_9466,N_9276);
nand U9724 (N_9724,N_9354,N_9281);
or U9725 (N_9725,N_9273,N_9394);
nor U9726 (N_9726,N_9448,N_9464);
xor U9727 (N_9727,N_9321,N_9260);
or U9728 (N_9728,N_9418,N_9449);
nand U9729 (N_9729,N_9406,N_9308);
nor U9730 (N_9730,N_9254,N_9387);
or U9731 (N_9731,N_9287,N_9345);
or U9732 (N_9732,N_9396,N_9477);
nand U9733 (N_9733,N_9481,N_9270);
or U9734 (N_9734,N_9341,N_9254);
xnor U9735 (N_9735,N_9381,N_9371);
nand U9736 (N_9736,N_9407,N_9325);
or U9737 (N_9737,N_9285,N_9258);
or U9738 (N_9738,N_9346,N_9459);
or U9739 (N_9739,N_9480,N_9407);
xnor U9740 (N_9740,N_9335,N_9477);
and U9741 (N_9741,N_9349,N_9442);
and U9742 (N_9742,N_9279,N_9266);
or U9743 (N_9743,N_9283,N_9351);
xnor U9744 (N_9744,N_9385,N_9464);
xnor U9745 (N_9745,N_9494,N_9453);
and U9746 (N_9746,N_9277,N_9408);
and U9747 (N_9747,N_9479,N_9349);
xnor U9748 (N_9748,N_9316,N_9283);
nor U9749 (N_9749,N_9399,N_9267);
and U9750 (N_9750,N_9661,N_9510);
xor U9751 (N_9751,N_9603,N_9692);
or U9752 (N_9752,N_9589,N_9610);
and U9753 (N_9753,N_9573,N_9636);
and U9754 (N_9754,N_9513,N_9709);
and U9755 (N_9755,N_9731,N_9644);
nand U9756 (N_9756,N_9745,N_9529);
nand U9757 (N_9757,N_9722,N_9602);
xnor U9758 (N_9758,N_9665,N_9574);
nor U9759 (N_9759,N_9627,N_9534);
or U9760 (N_9760,N_9648,N_9605);
or U9761 (N_9761,N_9645,N_9555);
xnor U9762 (N_9762,N_9683,N_9614);
or U9763 (N_9763,N_9626,N_9580);
nand U9764 (N_9764,N_9712,N_9638);
or U9765 (N_9765,N_9635,N_9507);
and U9766 (N_9766,N_9640,N_9564);
or U9767 (N_9767,N_9651,N_9595);
and U9768 (N_9768,N_9549,N_9578);
nor U9769 (N_9769,N_9524,N_9613);
and U9770 (N_9770,N_9526,N_9681);
or U9771 (N_9771,N_9667,N_9705);
xnor U9772 (N_9772,N_9678,N_9568);
xor U9773 (N_9773,N_9515,N_9565);
or U9774 (N_9774,N_9743,N_9634);
nor U9775 (N_9775,N_9695,N_9521);
nand U9776 (N_9776,N_9547,N_9542);
or U9777 (N_9777,N_9706,N_9536);
or U9778 (N_9778,N_9622,N_9567);
and U9779 (N_9779,N_9700,N_9673);
nand U9780 (N_9780,N_9530,N_9562);
nor U9781 (N_9781,N_9749,N_9672);
xor U9782 (N_9782,N_9646,N_9724);
or U9783 (N_9783,N_9747,N_9693);
or U9784 (N_9784,N_9615,N_9734);
nor U9785 (N_9785,N_9611,N_9554);
nand U9786 (N_9786,N_9561,N_9556);
xnor U9787 (N_9787,N_9713,N_9512);
or U9788 (N_9788,N_9525,N_9608);
xnor U9789 (N_9789,N_9650,N_9502);
and U9790 (N_9790,N_9514,N_9500);
xnor U9791 (N_9791,N_9694,N_9623);
nand U9792 (N_9792,N_9716,N_9730);
nand U9793 (N_9793,N_9620,N_9548);
and U9794 (N_9794,N_9617,N_9559);
or U9795 (N_9795,N_9541,N_9563);
xnor U9796 (N_9796,N_9552,N_9641);
or U9797 (N_9797,N_9582,N_9566);
nand U9798 (N_9798,N_9600,N_9660);
or U9799 (N_9799,N_9629,N_9686);
or U9800 (N_9800,N_9719,N_9590);
or U9801 (N_9801,N_9643,N_9717);
nor U9802 (N_9802,N_9710,N_9720);
and U9803 (N_9803,N_9704,N_9726);
or U9804 (N_9804,N_9517,N_9744);
or U9805 (N_9805,N_9715,N_9735);
xor U9806 (N_9806,N_9732,N_9505);
and U9807 (N_9807,N_9729,N_9532);
nand U9808 (N_9808,N_9733,N_9511);
xor U9809 (N_9809,N_9684,N_9642);
xnor U9810 (N_9810,N_9699,N_9689);
xor U9811 (N_9811,N_9668,N_9691);
and U9812 (N_9812,N_9551,N_9696);
xor U9813 (N_9813,N_9663,N_9609);
or U9814 (N_9814,N_9658,N_9736);
and U9815 (N_9815,N_9633,N_9560);
or U9816 (N_9816,N_9543,N_9569);
xor U9817 (N_9817,N_9528,N_9599);
or U9818 (N_9818,N_9588,N_9682);
and U9819 (N_9819,N_9674,N_9708);
xor U9820 (N_9820,N_9737,N_9619);
nand U9821 (N_9821,N_9680,N_9702);
xor U9822 (N_9822,N_9523,N_9746);
xnor U9823 (N_9823,N_9698,N_9557);
nand U9824 (N_9824,N_9508,N_9740);
or U9825 (N_9825,N_9607,N_9649);
or U9826 (N_9826,N_9718,N_9533);
nor U9827 (N_9827,N_9657,N_9503);
and U9828 (N_9828,N_9637,N_9516);
and U9829 (N_9829,N_9625,N_9520);
and U9830 (N_9830,N_9669,N_9553);
nand U9831 (N_9831,N_9538,N_9519);
xnor U9832 (N_9832,N_9654,N_9630);
and U9833 (N_9833,N_9628,N_9666);
nand U9834 (N_9834,N_9537,N_9583);
nor U9835 (N_9835,N_9527,N_9585);
xor U9836 (N_9836,N_9575,N_9741);
or U9837 (N_9837,N_9687,N_9518);
nand U9838 (N_9838,N_9631,N_9738);
nand U9839 (N_9839,N_9586,N_9545);
nor U9840 (N_9840,N_9621,N_9723);
or U9841 (N_9841,N_9577,N_9664);
nand U9842 (N_9842,N_9604,N_9504);
xnor U9843 (N_9843,N_9587,N_9612);
nand U9844 (N_9844,N_9618,N_9688);
xnor U9845 (N_9845,N_9725,N_9670);
nor U9846 (N_9846,N_9632,N_9539);
nand U9847 (N_9847,N_9739,N_9748);
xor U9848 (N_9848,N_9727,N_9616);
and U9849 (N_9849,N_9703,N_9711);
xnor U9850 (N_9850,N_9597,N_9506);
nand U9851 (N_9851,N_9581,N_9676);
nand U9852 (N_9852,N_9659,N_9697);
xor U9853 (N_9853,N_9594,N_9606);
xor U9854 (N_9854,N_9593,N_9584);
or U9855 (N_9855,N_9596,N_9509);
xnor U9856 (N_9856,N_9653,N_9592);
nor U9857 (N_9857,N_9571,N_9531);
nand U9858 (N_9858,N_9685,N_9591);
or U9859 (N_9859,N_9647,N_9550);
nand U9860 (N_9860,N_9707,N_9624);
or U9861 (N_9861,N_9721,N_9576);
and U9862 (N_9862,N_9579,N_9714);
nor U9863 (N_9863,N_9546,N_9656);
and U9864 (N_9864,N_9675,N_9652);
xor U9865 (N_9865,N_9677,N_9535);
or U9866 (N_9866,N_9558,N_9570);
and U9867 (N_9867,N_9540,N_9662);
or U9868 (N_9868,N_9598,N_9728);
nor U9869 (N_9869,N_9639,N_9522);
or U9870 (N_9870,N_9671,N_9601);
xnor U9871 (N_9871,N_9572,N_9501);
xnor U9872 (N_9872,N_9742,N_9679);
nand U9873 (N_9873,N_9655,N_9544);
and U9874 (N_9874,N_9701,N_9690);
and U9875 (N_9875,N_9599,N_9633);
xor U9876 (N_9876,N_9683,N_9586);
and U9877 (N_9877,N_9642,N_9741);
nor U9878 (N_9878,N_9632,N_9595);
nand U9879 (N_9879,N_9626,N_9513);
nand U9880 (N_9880,N_9563,N_9579);
xor U9881 (N_9881,N_9578,N_9709);
nand U9882 (N_9882,N_9588,N_9721);
nand U9883 (N_9883,N_9563,N_9736);
nand U9884 (N_9884,N_9509,N_9517);
or U9885 (N_9885,N_9532,N_9535);
or U9886 (N_9886,N_9681,N_9517);
nand U9887 (N_9887,N_9561,N_9660);
nor U9888 (N_9888,N_9543,N_9661);
xor U9889 (N_9889,N_9631,N_9617);
or U9890 (N_9890,N_9652,N_9566);
nand U9891 (N_9891,N_9585,N_9565);
xnor U9892 (N_9892,N_9596,N_9588);
nor U9893 (N_9893,N_9518,N_9664);
or U9894 (N_9894,N_9695,N_9657);
nand U9895 (N_9895,N_9533,N_9579);
xnor U9896 (N_9896,N_9523,N_9678);
nor U9897 (N_9897,N_9708,N_9587);
nor U9898 (N_9898,N_9656,N_9737);
and U9899 (N_9899,N_9696,N_9704);
nand U9900 (N_9900,N_9664,N_9665);
nor U9901 (N_9901,N_9662,N_9730);
or U9902 (N_9902,N_9597,N_9567);
and U9903 (N_9903,N_9573,N_9555);
nor U9904 (N_9904,N_9735,N_9622);
nor U9905 (N_9905,N_9639,N_9682);
nor U9906 (N_9906,N_9717,N_9567);
or U9907 (N_9907,N_9501,N_9535);
nor U9908 (N_9908,N_9586,N_9543);
or U9909 (N_9909,N_9515,N_9669);
nor U9910 (N_9910,N_9631,N_9701);
and U9911 (N_9911,N_9725,N_9594);
xnor U9912 (N_9912,N_9666,N_9678);
nor U9913 (N_9913,N_9594,N_9645);
nand U9914 (N_9914,N_9674,N_9642);
and U9915 (N_9915,N_9714,N_9736);
xor U9916 (N_9916,N_9636,N_9560);
nand U9917 (N_9917,N_9564,N_9665);
nor U9918 (N_9918,N_9562,N_9678);
xor U9919 (N_9919,N_9622,N_9666);
nand U9920 (N_9920,N_9566,N_9689);
nor U9921 (N_9921,N_9538,N_9500);
and U9922 (N_9922,N_9594,N_9549);
xnor U9923 (N_9923,N_9718,N_9505);
xnor U9924 (N_9924,N_9721,N_9651);
and U9925 (N_9925,N_9582,N_9528);
nand U9926 (N_9926,N_9510,N_9721);
nand U9927 (N_9927,N_9604,N_9699);
and U9928 (N_9928,N_9570,N_9556);
and U9929 (N_9929,N_9611,N_9503);
nand U9930 (N_9930,N_9656,N_9512);
and U9931 (N_9931,N_9726,N_9574);
or U9932 (N_9932,N_9710,N_9717);
or U9933 (N_9933,N_9545,N_9521);
nand U9934 (N_9934,N_9659,N_9614);
nor U9935 (N_9935,N_9609,N_9541);
or U9936 (N_9936,N_9661,N_9716);
or U9937 (N_9937,N_9674,N_9558);
xnor U9938 (N_9938,N_9707,N_9666);
nand U9939 (N_9939,N_9523,N_9687);
and U9940 (N_9940,N_9688,N_9518);
and U9941 (N_9941,N_9590,N_9566);
or U9942 (N_9942,N_9701,N_9630);
xnor U9943 (N_9943,N_9505,N_9740);
nor U9944 (N_9944,N_9638,N_9627);
or U9945 (N_9945,N_9628,N_9680);
nor U9946 (N_9946,N_9541,N_9558);
nand U9947 (N_9947,N_9634,N_9654);
or U9948 (N_9948,N_9706,N_9649);
xnor U9949 (N_9949,N_9702,N_9632);
and U9950 (N_9950,N_9577,N_9586);
and U9951 (N_9951,N_9605,N_9589);
and U9952 (N_9952,N_9533,N_9527);
and U9953 (N_9953,N_9667,N_9556);
nand U9954 (N_9954,N_9662,N_9580);
nor U9955 (N_9955,N_9717,N_9503);
and U9956 (N_9956,N_9587,N_9549);
xnor U9957 (N_9957,N_9720,N_9701);
and U9958 (N_9958,N_9537,N_9584);
nand U9959 (N_9959,N_9582,N_9642);
nand U9960 (N_9960,N_9683,N_9682);
and U9961 (N_9961,N_9670,N_9507);
xnor U9962 (N_9962,N_9605,N_9521);
and U9963 (N_9963,N_9705,N_9561);
xnor U9964 (N_9964,N_9641,N_9635);
nor U9965 (N_9965,N_9583,N_9500);
and U9966 (N_9966,N_9609,N_9531);
nor U9967 (N_9967,N_9545,N_9569);
and U9968 (N_9968,N_9660,N_9505);
xor U9969 (N_9969,N_9550,N_9736);
and U9970 (N_9970,N_9700,N_9631);
nor U9971 (N_9971,N_9734,N_9689);
nor U9972 (N_9972,N_9561,N_9522);
nand U9973 (N_9973,N_9717,N_9714);
nor U9974 (N_9974,N_9565,N_9551);
xnor U9975 (N_9975,N_9651,N_9690);
and U9976 (N_9976,N_9509,N_9739);
xor U9977 (N_9977,N_9734,N_9610);
nand U9978 (N_9978,N_9502,N_9581);
xnor U9979 (N_9979,N_9676,N_9574);
nor U9980 (N_9980,N_9693,N_9572);
xnor U9981 (N_9981,N_9513,N_9569);
nor U9982 (N_9982,N_9581,N_9568);
xor U9983 (N_9983,N_9603,N_9601);
xor U9984 (N_9984,N_9522,N_9512);
nor U9985 (N_9985,N_9640,N_9514);
nor U9986 (N_9986,N_9572,N_9547);
and U9987 (N_9987,N_9710,N_9533);
xor U9988 (N_9988,N_9628,N_9511);
or U9989 (N_9989,N_9502,N_9512);
xnor U9990 (N_9990,N_9599,N_9611);
nand U9991 (N_9991,N_9714,N_9742);
and U9992 (N_9992,N_9574,N_9541);
nand U9993 (N_9993,N_9729,N_9539);
and U9994 (N_9994,N_9542,N_9524);
and U9995 (N_9995,N_9706,N_9596);
and U9996 (N_9996,N_9546,N_9682);
nand U9997 (N_9997,N_9532,N_9725);
xnor U9998 (N_9998,N_9623,N_9510);
and U9999 (N_9999,N_9634,N_9564);
nor U10000 (N_10000,N_9802,N_9798);
nor U10001 (N_10001,N_9990,N_9836);
and U10002 (N_10002,N_9769,N_9835);
or U10003 (N_10003,N_9796,N_9892);
xnor U10004 (N_10004,N_9811,N_9823);
and U10005 (N_10005,N_9900,N_9801);
nor U10006 (N_10006,N_9807,N_9943);
and U10007 (N_10007,N_9767,N_9956);
xnor U10008 (N_10008,N_9987,N_9934);
xor U10009 (N_10009,N_9809,N_9978);
nand U10010 (N_10010,N_9783,N_9780);
xnor U10011 (N_10011,N_9760,N_9996);
or U10012 (N_10012,N_9989,N_9949);
nand U10013 (N_10013,N_9937,N_9763);
or U10014 (N_10014,N_9813,N_9812);
xor U10015 (N_10015,N_9974,N_9895);
and U10016 (N_10016,N_9926,N_9848);
xnor U10017 (N_10017,N_9877,N_9961);
nand U10018 (N_10018,N_9818,N_9947);
or U10019 (N_10019,N_9750,N_9994);
nand U10020 (N_10020,N_9817,N_9893);
xnor U10021 (N_10021,N_9983,N_9858);
or U10022 (N_10022,N_9757,N_9821);
xor U10023 (N_10023,N_9843,N_9850);
nor U10024 (N_10024,N_9753,N_9846);
or U10025 (N_10025,N_9953,N_9918);
or U10026 (N_10026,N_9762,N_9912);
xor U10027 (N_10027,N_9905,N_9768);
or U10028 (N_10028,N_9864,N_9884);
and U10029 (N_10029,N_9880,N_9857);
or U10030 (N_10030,N_9970,N_9828);
nor U10031 (N_10031,N_9794,N_9787);
or U10032 (N_10032,N_9792,N_9882);
xnor U10033 (N_10033,N_9826,N_9932);
xnor U10034 (N_10034,N_9906,N_9904);
or U10035 (N_10035,N_9907,N_9940);
xnor U10036 (N_10036,N_9921,N_9842);
xor U10037 (N_10037,N_9825,N_9751);
and U10038 (N_10038,N_9863,N_9942);
xor U10039 (N_10039,N_9824,N_9764);
nor U10040 (N_10040,N_9831,N_9916);
nor U10041 (N_10041,N_9952,N_9804);
or U10042 (N_10042,N_9955,N_9833);
xor U10043 (N_10043,N_9992,N_9883);
and U10044 (N_10044,N_9861,N_9946);
nor U10045 (N_10045,N_9856,N_9908);
nor U10046 (N_10046,N_9982,N_9964);
nor U10047 (N_10047,N_9944,N_9951);
xor U10048 (N_10048,N_9776,N_9939);
or U10049 (N_10049,N_9841,N_9967);
and U10050 (N_10050,N_9997,N_9933);
or U10051 (N_10051,N_9795,N_9866);
nor U10052 (N_10052,N_9765,N_9847);
or U10053 (N_10053,N_9920,N_9781);
nor U10054 (N_10054,N_9868,N_9993);
or U10055 (N_10055,N_9957,N_9761);
or U10056 (N_10056,N_9985,N_9919);
or U10057 (N_10057,N_9991,N_9976);
or U10058 (N_10058,N_9815,N_9894);
or U10059 (N_10059,N_9984,N_9810);
nand U10060 (N_10060,N_9851,N_9928);
nor U10061 (N_10061,N_9754,N_9988);
xnor U10062 (N_10062,N_9786,N_9936);
nand U10063 (N_10063,N_9859,N_9797);
or U10064 (N_10064,N_9779,N_9845);
or U10065 (N_10065,N_9816,N_9938);
nand U10066 (N_10066,N_9924,N_9980);
xnor U10067 (N_10067,N_9909,N_9948);
or U10068 (N_10068,N_9929,N_9903);
or U10069 (N_10069,N_9844,N_9925);
nand U10070 (N_10070,N_9840,N_9962);
nor U10071 (N_10071,N_9910,N_9897);
nor U10072 (N_10072,N_9775,N_9838);
and U10073 (N_10073,N_9782,N_9899);
xor U10074 (N_10074,N_9777,N_9945);
xnor U10075 (N_10075,N_9881,N_9986);
nand U10076 (N_10076,N_9865,N_9879);
or U10077 (N_10077,N_9902,N_9885);
nand U10078 (N_10078,N_9771,N_9873);
xnor U10079 (N_10079,N_9791,N_9875);
nor U10080 (N_10080,N_9959,N_9898);
nor U10081 (N_10081,N_9788,N_9832);
nor U10082 (N_10082,N_9888,N_9837);
xor U10083 (N_10083,N_9886,N_9758);
xor U10084 (N_10084,N_9772,N_9871);
and U10085 (N_10085,N_9820,N_9773);
nor U10086 (N_10086,N_9774,N_9914);
and U10087 (N_10087,N_9806,N_9849);
nand U10088 (N_10088,N_9935,N_9852);
and U10089 (N_10089,N_9950,N_9822);
and U10090 (N_10090,N_9834,N_9805);
and U10091 (N_10091,N_9759,N_9887);
nor U10092 (N_10092,N_9869,N_9917);
nor U10093 (N_10093,N_9790,N_9930);
xor U10094 (N_10094,N_9941,N_9874);
nand U10095 (N_10095,N_9789,N_9855);
nor U10096 (N_10096,N_9870,N_9814);
and U10097 (N_10097,N_9799,N_9922);
or U10098 (N_10098,N_9829,N_9927);
or U10099 (N_10099,N_9878,N_9913);
nand U10100 (N_10100,N_9911,N_9965);
and U10101 (N_10101,N_9839,N_9931);
and U10102 (N_10102,N_9972,N_9891);
nor U10103 (N_10103,N_9819,N_9979);
xnor U10104 (N_10104,N_9901,N_9808);
nor U10105 (N_10105,N_9977,N_9889);
or U10106 (N_10106,N_9784,N_9973);
or U10107 (N_10107,N_9890,N_9860);
and U10108 (N_10108,N_9755,N_9766);
or U10109 (N_10109,N_9999,N_9923);
nor U10110 (N_10110,N_9872,N_9915);
nor U10111 (N_10111,N_9975,N_9756);
or U10112 (N_10112,N_9770,N_9778);
nor U10113 (N_10113,N_9862,N_9830);
or U10114 (N_10114,N_9785,N_9800);
xor U10115 (N_10115,N_9958,N_9803);
and U10116 (N_10116,N_9960,N_9968);
nor U10117 (N_10117,N_9966,N_9969);
nor U10118 (N_10118,N_9752,N_9854);
or U10119 (N_10119,N_9981,N_9998);
or U10120 (N_10120,N_9793,N_9954);
or U10121 (N_10121,N_9963,N_9876);
or U10122 (N_10122,N_9827,N_9867);
nand U10123 (N_10123,N_9853,N_9971);
and U10124 (N_10124,N_9896,N_9995);
nand U10125 (N_10125,N_9948,N_9817);
nor U10126 (N_10126,N_9888,N_9905);
xnor U10127 (N_10127,N_9915,N_9888);
xor U10128 (N_10128,N_9844,N_9792);
or U10129 (N_10129,N_9899,N_9818);
or U10130 (N_10130,N_9793,N_9900);
and U10131 (N_10131,N_9912,N_9863);
and U10132 (N_10132,N_9931,N_9791);
nand U10133 (N_10133,N_9990,N_9903);
xnor U10134 (N_10134,N_9789,N_9896);
and U10135 (N_10135,N_9837,N_9999);
nor U10136 (N_10136,N_9868,N_9829);
or U10137 (N_10137,N_9825,N_9859);
or U10138 (N_10138,N_9787,N_9858);
and U10139 (N_10139,N_9782,N_9948);
or U10140 (N_10140,N_9849,N_9768);
or U10141 (N_10141,N_9902,N_9789);
or U10142 (N_10142,N_9833,N_9900);
nor U10143 (N_10143,N_9824,N_9920);
and U10144 (N_10144,N_9869,N_9879);
and U10145 (N_10145,N_9991,N_9875);
or U10146 (N_10146,N_9877,N_9939);
nor U10147 (N_10147,N_9798,N_9978);
or U10148 (N_10148,N_9791,N_9804);
nand U10149 (N_10149,N_9851,N_9903);
and U10150 (N_10150,N_9828,N_9884);
or U10151 (N_10151,N_9812,N_9880);
nand U10152 (N_10152,N_9863,N_9828);
nand U10153 (N_10153,N_9796,N_9915);
and U10154 (N_10154,N_9873,N_9985);
and U10155 (N_10155,N_9987,N_9806);
nand U10156 (N_10156,N_9887,N_9861);
nor U10157 (N_10157,N_9885,N_9903);
and U10158 (N_10158,N_9908,N_9938);
and U10159 (N_10159,N_9939,N_9946);
or U10160 (N_10160,N_9976,N_9767);
nor U10161 (N_10161,N_9929,N_9770);
nor U10162 (N_10162,N_9803,N_9751);
xnor U10163 (N_10163,N_9817,N_9854);
or U10164 (N_10164,N_9790,N_9903);
nand U10165 (N_10165,N_9792,N_9996);
nor U10166 (N_10166,N_9914,N_9977);
nand U10167 (N_10167,N_9761,N_9902);
and U10168 (N_10168,N_9861,N_9874);
xnor U10169 (N_10169,N_9754,N_9935);
or U10170 (N_10170,N_9956,N_9959);
nor U10171 (N_10171,N_9848,N_9981);
and U10172 (N_10172,N_9848,N_9910);
xnor U10173 (N_10173,N_9979,N_9807);
nor U10174 (N_10174,N_9861,N_9849);
and U10175 (N_10175,N_9841,N_9793);
xnor U10176 (N_10176,N_9949,N_9942);
xor U10177 (N_10177,N_9880,N_9993);
or U10178 (N_10178,N_9989,N_9799);
nand U10179 (N_10179,N_9976,N_9898);
xor U10180 (N_10180,N_9976,N_9899);
and U10181 (N_10181,N_9944,N_9978);
or U10182 (N_10182,N_9852,N_9932);
and U10183 (N_10183,N_9807,N_9881);
xor U10184 (N_10184,N_9896,N_9767);
nor U10185 (N_10185,N_9898,N_9870);
nand U10186 (N_10186,N_9845,N_9921);
and U10187 (N_10187,N_9841,N_9968);
nand U10188 (N_10188,N_9924,N_9888);
nand U10189 (N_10189,N_9972,N_9813);
or U10190 (N_10190,N_9941,N_9948);
nor U10191 (N_10191,N_9900,N_9827);
nor U10192 (N_10192,N_9858,N_9829);
xor U10193 (N_10193,N_9828,N_9951);
xor U10194 (N_10194,N_9951,N_9878);
or U10195 (N_10195,N_9782,N_9976);
or U10196 (N_10196,N_9943,N_9776);
xnor U10197 (N_10197,N_9869,N_9788);
or U10198 (N_10198,N_9870,N_9979);
xor U10199 (N_10199,N_9824,N_9931);
nor U10200 (N_10200,N_9850,N_9753);
xor U10201 (N_10201,N_9982,N_9966);
nor U10202 (N_10202,N_9779,N_9936);
or U10203 (N_10203,N_9968,N_9785);
nor U10204 (N_10204,N_9789,N_9894);
xnor U10205 (N_10205,N_9822,N_9815);
xnor U10206 (N_10206,N_9978,N_9892);
xnor U10207 (N_10207,N_9805,N_9877);
xor U10208 (N_10208,N_9795,N_9801);
nor U10209 (N_10209,N_9831,N_9917);
nand U10210 (N_10210,N_9880,N_9909);
or U10211 (N_10211,N_9817,N_9907);
nor U10212 (N_10212,N_9985,N_9790);
xnor U10213 (N_10213,N_9796,N_9919);
xnor U10214 (N_10214,N_9908,N_9873);
and U10215 (N_10215,N_9879,N_9891);
nor U10216 (N_10216,N_9798,N_9944);
xor U10217 (N_10217,N_9910,N_9847);
nand U10218 (N_10218,N_9754,N_9887);
nand U10219 (N_10219,N_9815,N_9851);
and U10220 (N_10220,N_9945,N_9761);
or U10221 (N_10221,N_9816,N_9856);
nand U10222 (N_10222,N_9859,N_9974);
nand U10223 (N_10223,N_9859,N_9758);
xnor U10224 (N_10224,N_9908,N_9945);
or U10225 (N_10225,N_9882,N_9928);
nor U10226 (N_10226,N_9860,N_9933);
or U10227 (N_10227,N_9776,N_9875);
nand U10228 (N_10228,N_9783,N_9778);
nor U10229 (N_10229,N_9959,N_9764);
and U10230 (N_10230,N_9965,N_9798);
xnor U10231 (N_10231,N_9857,N_9850);
nand U10232 (N_10232,N_9815,N_9950);
xnor U10233 (N_10233,N_9782,N_9916);
xnor U10234 (N_10234,N_9857,N_9778);
or U10235 (N_10235,N_9850,N_9863);
or U10236 (N_10236,N_9997,N_9911);
nand U10237 (N_10237,N_9802,N_9870);
xor U10238 (N_10238,N_9937,N_9965);
xor U10239 (N_10239,N_9838,N_9944);
xor U10240 (N_10240,N_9761,N_9922);
nor U10241 (N_10241,N_9829,N_9844);
xnor U10242 (N_10242,N_9780,N_9901);
and U10243 (N_10243,N_9811,N_9830);
xor U10244 (N_10244,N_9875,N_9753);
nor U10245 (N_10245,N_9910,N_9974);
and U10246 (N_10246,N_9925,N_9752);
or U10247 (N_10247,N_9761,N_9884);
nor U10248 (N_10248,N_9753,N_9871);
or U10249 (N_10249,N_9995,N_9815);
xnor U10250 (N_10250,N_10079,N_10242);
or U10251 (N_10251,N_10012,N_10014);
xnor U10252 (N_10252,N_10180,N_10123);
and U10253 (N_10253,N_10068,N_10111);
and U10254 (N_10254,N_10228,N_10036);
and U10255 (N_10255,N_10131,N_10065);
and U10256 (N_10256,N_10201,N_10247);
xnor U10257 (N_10257,N_10216,N_10053);
nor U10258 (N_10258,N_10207,N_10233);
nor U10259 (N_10259,N_10006,N_10052);
and U10260 (N_10260,N_10025,N_10210);
xor U10261 (N_10261,N_10167,N_10114);
xnor U10262 (N_10262,N_10077,N_10175);
nor U10263 (N_10263,N_10090,N_10191);
nand U10264 (N_10264,N_10059,N_10085);
xor U10265 (N_10265,N_10100,N_10154);
or U10266 (N_10266,N_10092,N_10110);
or U10267 (N_10267,N_10027,N_10064);
nor U10268 (N_10268,N_10023,N_10058);
or U10269 (N_10269,N_10098,N_10245);
nor U10270 (N_10270,N_10187,N_10151);
nand U10271 (N_10271,N_10196,N_10209);
nor U10272 (N_10272,N_10190,N_10057);
nor U10273 (N_10273,N_10115,N_10109);
xor U10274 (N_10274,N_10135,N_10072);
nand U10275 (N_10275,N_10222,N_10044);
xnor U10276 (N_10276,N_10112,N_10067);
nand U10277 (N_10277,N_10129,N_10140);
xor U10278 (N_10278,N_10192,N_10125);
nand U10279 (N_10279,N_10198,N_10083);
or U10280 (N_10280,N_10087,N_10020);
or U10281 (N_10281,N_10062,N_10105);
xnor U10282 (N_10282,N_10226,N_10005);
and U10283 (N_10283,N_10047,N_10091);
and U10284 (N_10284,N_10214,N_10069);
nand U10285 (N_10285,N_10134,N_10162);
or U10286 (N_10286,N_10074,N_10035);
or U10287 (N_10287,N_10004,N_10204);
xor U10288 (N_10288,N_10136,N_10238);
or U10289 (N_10289,N_10021,N_10249);
or U10290 (N_10290,N_10063,N_10119);
xor U10291 (N_10291,N_10080,N_10248);
nand U10292 (N_10292,N_10128,N_10193);
or U10293 (N_10293,N_10246,N_10102);
and U10294 (N_10294,N_10212,N_10026);
nand U10295 (N_10295,N_10078,N_10173);
nor U10296 (N_10296,N_10039,N_10009);
nand U10297 (N_10297,N_10197,N_10073);
nor U10298 (N_10298,N_10213,N_10060);
xor U10299 (N_10299,N_10008,N_10095);
xor U10300 (N_10300,N_10041,N_10202);
xor U10301 (N_10301,N_10132,N_10164);
nand U10302 (N_10302,N_10042,N_10051);
and U10303 (N_10303,N_10241,N_10031);
or U10304 (N_10304,N_10148,N_10024);
xnor U10305 (N_10305,N_10094,N_10130);
nor U10306 (N_10306,N_10161,N_10169);
or U10307 (N_10307,N_10243,N_10182);
nand U10308 (N_10308,N_10231,N_10118);
nand U10309 (N_10309,N_10108,N_10200);
or U10310 (N_10310,N_10103,N_10055);
nand U10311 (N_10311,N_10218,N_10019);
or U10312 (N_10312,N_10106,N_10208);
nand U10313 (N_10313,N_10240,N_10040);
and U10314 (N_10314,N_10244,N_10217);
xnor U10315 (N_10315,N_10194,N_10230);
and U10316 (N_10316,N_10116,N_10152);
xor U10317 (N_10317,N_10237,N_10121);
nor U10318 (N_10318,N_10104,N_10015);
and U10319 (N_10319,N_10185,N_10029);
nand U10320 (N_10320,N_10211,N_10168);
nand U10321 (N_10321,N_10163,N_10143);
or U10322 (N_10322,N_10045,N_10120);
nand U10323 (N_10323,N_10165,N_10007);
and U10324 (N_10324,N_10166,N_10050);
nor U10325 (N_10325,N_10232,N_10221);
and U10326 (N_10326,N_10219,N_10127);
nand U10327 (N_10327,N_10113,N_10234);
and U10328 (N_10328,N_10195,N_10158);
nand U10329 (N_10329,N_10093,N_10013);
xor U10330 (N_10330,N_10066,N_10199);
xnor U10331 (N_10331,N_10002,N_10137);
or U10332 (N_10332,N_10084,N_10149);
nor U10333 (N_10333,N_10033,N_10082);
or U10334 (N_10334,N_10122,N_10049);
nor U10335 (N_10335,N_10043,N_10178);
or U10336 (N_10336,N_10205,N_10117);
or U10337 (N_10337,N_10146,N_10223);
or U10338 (N_10338,N_10086,N_10177);
or U10339 (N_10339,N_10088,N_10181);
nand U10340 (N_10340,N_10070,N_10139);
xnor U10341 (N_10341,N_10028,N_10096);
and U10342 (N_10342,N_10157,N_10133);
xor U10343 (N_10343,N_10153,N_10046);
nand U10344 (N_10344,N_10101,N_10016);
and U10345 (N_10345,N_10038,N_10075);
xor U10346 (N_10346,N_10147,N_10126);
nand U10347 (N_10347,N_10022,N_10107);
or U10348 (N_10348,N_10076,N_10215);
and U10349 (N_10349,N_10145,N_10037);
xor U10350 (N_10350,N_10048,N_10225);
nand U10351 (N_10351,N_10089,N_10001);
xnor U10352 (N_10352,N_10138,N_10189);
nand U10353 (N_10353,N_10097,N_10054);
and U10354 (N_10354,N_10056,N_10010);
xnor U10355 (N_10355,N_10170,N_10183);
and U10356 (N_10356,N_10011,N_10071);
and U10357 (N_10357,N_10171,N_10155);
or U10358 (N_10358,N_10099,N_10159);
or U10359 (N_10359,N_10186,N_10142);
and U10360 (N_10360,N_10176,N_10160);
nand U10361 (N_10361,N_10061,N_10124);
nor U10362 (N_10362,N_10206,N_10229);
nor U10363 (N_10363,N_10236,N_10184);
nor U10364 (N_10364,N_10220,N_10239);
xor U10365 (N_10365,N_10235,N_10179);
or U10366 (N_10366,N_10018,N_10003);
and U10367 (N_10367,N_10034,N_10156);
and U10368 (N_10368,N_10188,N_10081);
or U10369 (N_10369,N_10141,N_10144);
and U10370 (N_10370,N_10172,N_10032);
and U10371 (N_10371,N_10203,N_10174);
or U10372 (N_10372,N_10000,N_10224);
or U10373 (N_10373,N_10150,N_10017);
xnor U10374 (N_10374,N_10030,N_10227);
xor U10375 (N_10375,N_10017,N_10097);
nand U10376 (N_10376,N_10022,N_10244);
nor U10377 (N_10377,N_10156,N_10002);
nor U10378 (N_10378,N_10053,N_10131);
and U10379 (N_10379,N_10189,N_10067);
and U10380 (N_10380,N_10018,N_10093);
nor U10381 (N_10381,N_10185,N_10072);
nand U10382 (N_10382,N_10110,N_10125);
xnor U10383 (N_10383,N_10225,N_10203);
xor U10384 (N_10384,N_10077,N_10168);
or U10385 (N_10385,N_10079,N_10046);
nor U10386 (N_10386,N_10102,N_10192);
or U10387 (N_10387,N_10197,N_10043);
or U10388 (N_10388,N_10011,N_10066);
xor U10389 (N_10389,N_10182,N_10037);
and U10390 (N_10390,N_10009,N_10139);
nor U10391 (N_10391,N_10019,N_10029);
and U10392 (N_10392,N_10158,N_10156);
xor U10393 (N_10393,N_10125,N_10061);
or U10394 (N_10394,N_10148,N_10010);
nor U10395 (N_10395,N_10210,N_10013);
nand U10396 (N_10396,N_10101,N_10241);
and U10397 (N_10397,N_10212,N_10158);
nand U10398 (N_10398,N_10161,N_10043);
or U10399 (N_10399,N_10047,N_10168);
and U10400 (N_10400,N_10176,N_10011);
and U10401 (N_10401,N_10030,N_10212);
nor U10402 (N_10402,N_10036,N_10022);
or U10403 (N_10403,N_10030,N_10115);
nand U10404 (N_10404,N_10071,N_10172);
and U10405 (N_10405,N_10243,N_10153);
xnor U10406 (N_10406,N_10183,N_10202);
xor U10407 (N_10407,N_10244,N_10156);
nand U10408 (N_10408,N_10175,N_10152);
or U10409 (N_10409,N_10171,N_10085);
and U10410 (N_10410,N_10160,N_10039);
nand U10411 (N_10411,N_10050,N_10000);
or U10412 (N_10412,N_10161,N_10152);
nand U10413 (N_10413,N_10051,N_10249);
and U10414 (N_10414,N_10070,N_10039);
and U10415 (N_10415,N_10105,N_10066);
nand U10416 (N_10416,N_10181,N_10029);
and U10417 (N_10417,N_10236,N_10034);
and U10418 (N_10418,N_10213,N_10021);
xnor U10419 (N_10419,N_10118,N_10249);
xor U10420 (N_10420,N_10200,N_10062);
xor U10421 (N_10421,N_10046,N_10098);
xor U10422 (N_10422,N_10157,N_10033);
nor U10423 (N_10423,N_10141,N_10108);
nand U10424 (N_10424,N_10019,N_10092);
nand U10425 (N_10425,N_10009,N_10052);
and U10426 (N_10426,N_10210,N_10003);
or U10427 (N_10427,N_10040,N_10151);
nand U10428 (N_10428,N_10184,N_10182);
nor U10429 (N_10429,N_10134,N_10194);
and U10430 (N_10430,N_10111,N_10102);
xnor U10431 (N_10431,N_10009,N_10044);
and U10432 (N_10432,N_10062,N_10114);
or U10433 (N_10433,N_10152,N_10242);
nor U10434 (N_10434,N_10208,N_10243);
nand U10435 (N_10435,N_10151,N_10235);
or U10436 (N_10436,N_10020,N_10209);
nor U10437 (N_10437,N_10167,N_10056);
xnor U10438 (N_10438,N_10142,N_10028);
and U10439 (N_10439,N_10053,N_10069);
or U10440 (N_10440,N_10208,N_10056);
xnor U10441 (N_10441,N_10094,N_10100);
and U10442 (N_10442,N_10150,N_10144);
or U10443 (N_10443,N_10050,N_10178);
or U10444 (N_10444,N_10071,N_10004);
nand U10445 (N_10445,N_10057,N_10129);
nand U10446 (N_10446,N_10017,N_10039);
or U10447 (N_10447,N_10056,N_10247);
nor U10448 (N_10448,N_10093,N_10196);
or U10449 (N_10449,N_10014,N_10113);
or U10450 (N_10450,N_10133,N_10009);
nand U10451 (N_10451,N_10021,N_10167);
or U10452 (N_10452,N_10057,N_10189);
nor U10453 (N_10453,N_10030,N_10208);
and U10454 (N_10454,N_10030,N_10124);
or U10455 (N_10455,N_10079,N_10156);
or U10456 (N_10456,N_10047,N_10078);
nor U10457 (N_10457,N_10213,N_10249);
and U10458 (N_10458,N_10162,N_10131);
nor U10459 (N_10459,N_10082,N_10225);
nor U10460 (N_10460,N_10171,N_10166);
nand U10461 (N_10461,N_10031,N_10076);
or U10462 (N_10462,N_10222,N_10105);
nand U10463 (N_10463,N_10239,N_10194);
nand U10464 (N_10464,N_10119,N_10207);
nand U10465 (N_10465,N_10187,N_10132);
or U10466 (N_10466,N_10048,N_10078);
nand U10467 (N_10467,N_10032,N_10191);
or U10468 (N_10468,N_10191,N_10003);
nand U10469 (N_10469,N_10244,N_10106);
xnor U10470 (N_10470,N_10018,N_10168);
and U10471 (N_10471,N_10049,N_10223);
nand U10472 (N_10472,N_10045,N_10160);
and U10473 (N_10473,N_10049,N_10167);
and U10474 (N_10474,N_10155,N_10008);
nor U10475 (N_10475,N_10038,N_10057);
xnor U10476 (N_10476,N_10104,N_10077);
xor U10477 (N_10477,N_10086,N_10007);
or U10478 (N_10478,N_10210,N_10002);
nand U10479 (N_10479,N_10181,N_10122);
or U10480 (N_10480,N_10007,N_10063);
nor U10481 (N_10481,N_10241,N_10248);
xor U10482 (N_10482,N_10176,N_10109);
or U10483 (N_10483,N_10161,N_10091);
xor U10484 (N_10484,N_10156,N_10151);
nor U10485 (N_10485,N_10037,N_10088);
nor U10486 (N_10486,N_10118,N_10077);
nand U10487 (N_10487,N_10172,N_10192);
or U10488 (N_10488,N_10179,N_10162);
xor U10489 (N_10489,N_10023,N_10130);
xnor U10490 (N_10490,N_10039,N_10087);
and U10491 (N_10491,N_10092,N_10151);
or U10492 (N_10492,N_10018,N_10213);
or U10493 (N_10493,N_10091,N_10111);
nor U10494 (N_10494,N_10175,N_10133);
nor U10495 (N_10495,N_10238,N_10214);
nor U10496 (N_10496,N_10011,N_10226);
nor U10497 (N_10497,N_10191,N_10179);
xor U10498 (N_10498,N_10003,N_10041);
xor U10499 (N_10499,N_10138,N_10067);
nand U10500 (N_10500,N_10404,N_10316);
xor U10501 (N_10501,N_10420,N_10493);
or U10502 (N_10502,N_10481,N_10289);
or U10503 (N_10503,N_10498,N_10334);
or U10504 (N_10504,N_10441,N_10415);
nand U10505 (N_10505,N_10308,N_10407);
xnor U10506 (N_10506,N_10479,N_10497);
or U10507 (N_10507,N_10409,N_10421);
and U10508 (N_10508,N_10355,N_10259);
nor U10509 (N_10509,N_10450,N_10480);
or U10510 (N_10510,N_10358,N_10344);
nand U10511 (N_10511,N_10368,N_10466);
and U10512 (N_10512,N_10485,N_10430);
nor U10513 (N_10513,N_10406,N_10326);
nand U10514 (N_10514,N_10490,N_10268);
xnor U10515 (N_10515,N_10295,N_10284);
or U10516 (N_10516,N_10291,N_10294);
xnor U10517 (N_10517,N_10317,N_10455);
nand U10518 (N_10518,N_10427,N_10474);
or U10519 (N_10519,N_10258,N_10297);
and U10520 (N_10520,N_10448,N_10390);
or U10521 (N_10521,N_10413,N_10496);
nor U10522 (N_10522,N_10449,N_10387);
nand U10523 (N_10523,N_10462,N_10276);
and U10524 (N_10524,N_10264,N_10440);
xor U10525 (N_10525,N_10352,N_10431);
and U10526 (N_10526,N_10353,N_10408);
xor U10527 (N_10527,N_10381,N_10312);
nand U10528 (N_10528,N_10321,N_10262);
nor U10529 (N_10529,N_10320,N_10301);
nand U10530 (N_10530,N_10345,N_10444);
nor U10531 (N_10531,N_10454,N_10476);
nor U10532 (N_10532,N_10475,N_10460);
or U10533 (N_10533,N_10482,N_10278);
and U10534 (N_10534,N_10477,N_10438);
or U10535 (N_10535,N_10456,N_10329);
xnor U10536 (N_10536,N_10467,N_10332);
or U10537 (N_10537,N_10279,N_10377);
nor U10538 (N_10538,N_10275,N_10434);
or U10539 (N_10539,N_10311,N_10389);
nor U10540 (N_10540,N_10388,N_10324);
nor U10541 (N_10541,N_10269,N_10280);
nand U10542 (N_10542,N_10288,N_10260);
nand U10543 (N_10543,N_10299,N_10364);
or U10544 (N_10544,N_10298,N_10370);
or U10545 (N_10545,N_10419,N_10447);
and U10546 (N_10546,N_10402,N_10399);
or U10547 (N_10547,N_10470,N_10486);
nand U10548 (N_10548,N_10302,N_10433);
xor U10549 (N_10549,N_10263,N_10397);
xnor U10550 (N_10550,N_10256,N_10471);
nand U10551 (N_10551,N_10322,N_10310);
nand U10552 (N_10552,N_10250,N_10376);
or U10553 (N_10553,N_10484,N_10341);
and U10554 (N_10554,N_10338,N_10453);
xor U10555 (N_10555,N_10361,N_10369);
xor U10556 (N_10556,N_10380,N_10357);
nor U10557 (N_10557,N_10468,N_10267);
or U10558 (N_10558,N_10451,N_10461);
xnor U10559 (N_10559,N_10285,N_10305);
xor U10560 (N_10560,N_10383,N_10348);
nor U10561 (N_10561,N_10394,N_10346);
xnor U10562 (N_10562,N_10432,N_10281);
nor U10563 (N_10563,N_10417,N_10422);
nand U10564 (N_10564,N_10391,N_10253);
or U10565 (N_10565,N_10292,N_10273);
and U10566 (N_10566,N_10499,N_10405);
or U10567 (N_10567,N_10379,N_10435);
nor U10568 (N_10568,N_10403,N_10360);
xor U10569 (N_10569,N_10314,N_10365);
nor U10570 (N_10570,N_10489,N_10495);
nor U10571 (N_10571,N_10335,N_10429);
nor U10572 (N_10572,N_10296,N_10330);
or U10573 (N_10573,N_10488,N_10473);
nor U10574 (N_10574,N_10266,N_10392);
and U10575 (N_10575,N_10411,N_10319);
nand U10576 (N_10576,N_10272,N_10342);
or U10577 (N_10577,N_10463,N_10439);
nand U10578 (N_10578,N_10286,N_10437);
or U10579 (N_10579,N_10374,N_10293);
nor U10580 (N_10580,N_10382,N_10414);
or U10581 (N_10581,N_10478,N_10412);
nor U10582 (N_10582,N_10323,N_10339);
nor U10583 (N_10583,N_10359,N_10303);
or U10584 (N_10584,N_10337,N_10343);
nor U10585 (N_10585,N_10315,N_10452);
nand U10586 (N_10586,N_10347,N_10401);
xor U10587 (N_10587,N_10325,N_10363);
nor U10588 (N_10588,N_10261,N_10464);
or U10589 (N_10589,N_10410,N_10252);
nor U10590 (N_10590,N_10328,N_10265);
xnor U10591 (N_10591,N_10426,N_10457);
and U10592 (N_10592,N_10400,N_10386);
xnor U10593 (N_10593,N_10396,N_10251);
or U10594 (N_10594,N_10459,N_10270);
or U10595 (N_10595,N_10255,N_10443);
nor U10596 (N_10596,N_10425,N_10416);
nor U10597 (N_10597,N_10327,N_10366);
nor U10598 (N_10598,N_10436,N_10398);
nand U10599 (N_10599,N_10306,N_10340);
nand U10600 (N_10600,N_10304,N_10349);
and U10601 (N_10601,N_10336,N_10469);
nand U10602 (N_10602,N_10445,N_10290);
nand U10603 (N_10603,N_10307,N_10442);
nor U10604 (N_10604,N_10483,N_10492);
nor U10605 (N_10605,N_10384,N_10313);
nand U10606 (N_10606,N_10418,N_10283);
or U10607 (N_10607,N_10351,N_10282);
or U10608 (N_10608,N_10487,N_10472);
nand U10609 (N_10609,N_10424,N_10354);
nand U10610 (N_10610,N_10318,N_10423);
or U10611 (N_10611,N_10309,N_10257);
nor U10612 (N_10612,N_10375,N_10494);
nand U10613 (N_10613,N_10362,N_10395);
nand U10614 (N_10614,N_10277,N_10446);
nor U10615 (N_10615,N_10373,N_10385);
and U10616 (N_10616,N_10333,N_10350);
xnor U10617 (N_10617,N_10491,N_10274);
xnor U10618 (N_10618,N_10393,N_10465);
or U10619 (N_10619,N_10458,N_10287);
and U10620 (N_10620,N_10378,N_10271);
or U10621 (N_10621,N_10300,N_10254);
nand U10622 (N_10622,N_10331,N_10372);
nand U10623 (N_10623,N_10428,N_10371);
nor U10624 (N_10624,N_10356,N_10367);
or U10625 (N_10625,N_10319,N_10481);
xnor U10626 (N_10626,N_10380,N_10471);
or U10627 (N_10627,N_10498,N_10430);
or U10628 (N_10628,N_10462,N_10289);
nand U10629 (N_10629,N_10318,N_10424);
xor U10630 (N_10630,N_10431,N_10476);
xnor U10631 (N_10631,N_10348,N_10304);
or U10632 (N_10632,N_10465,N_10272);
and U10633 (N_10633,N_10486,N_10327);
and U10634 (N_10634,N_10341,N_10426);
xnor U10635 (N_10635,N_10340,N_10302);
nor U10636 (N_10636,N_10300,N_10477);
nand U10637 (N_10637,N_10352,N_10423);
or U10638 (N_10638,N_10324,N_10322);
nor U10639 (N_10639,N_10322,N_10314);
and U10640 (N_10640,N_10400,N_10445);
and U10641 (N_10641,N_10341,N_10336);
xnor U10642 (N_10642,N_10466,N_10250);
nor U10643 (N_10643,N_10339,N_10288);
or U10644 (N_10644,N_10279,N_10406);
or U10645 (N_10645,N_10316,N_10356);
nor U10646 (N_10646,N_10489,N_10474);
nor U10647 (N_10647,N_10317,N_10306);
or U10648 (N_10648,N_10282,N_10356);
xor U10649 (N_10649,N_10391,N_10272);
nand U10650 (N_10650,N_10371,N_10264);
and U10651 (N_10651,N_10306,N_10444);
xor U10652 (N_10652,N_10427,N_10399);
or U10653 (N_10653,N_10423,N_10366);
xor U10654 (N_10654,N_10485,N_10296);
xor U10655 (N_10655,N_10439,N_10312);
or U10656 (N_10656,N_10355,N_10439);
nor U10657 (N_10657,N_10422,N_10472);
and U10658 (N_10658,N_10283,N_10451);
and U10659 (N_10659,N_10387,N_10268);
xor U10660 (N_10660,N_10347,N_10409);
and U10661 (N_10661,N_10394,N_10365);
xor U10662 (N_10662,N_10352,N_10258);
xnor U10663 (N_10663,N_10432,N_10418);
and U10664 (N_10664,N_10337,N_10283);
or U10665 (N_10665,N_10405,N_10290);
or U10666 (N_10666,N_10472,N_10401);
nand U10667 (N_10667,N_10299,N_10413);
nand U10668 (N_10668,N_10484,N_10345);
and U10669 (N_10669,N_10345,N_10257);
nor U10670 (N_10670,N_10389,N_10484);
and U10671 (N_10671,N_10295,N_10376);
nor U10672 (N_10672,N_10428,N_10366);
nor U10673 (N_10673,N_10293,N_10393);
xor U10674 (N_10674,N_10421,N_10487);
xnor U10675 (N_10675,N_10407,N_10460);
nand U10676 (N_10676,N_10419,N_10411);
and U10677 (N_10677,N_10494,N_10262);
and U10678 (N_10678,N_10346,N_10462);
xor U10679 (N_10679,N_10492,N_10449);
and U10680 (N_10680,N_10282,N_10419);
nor U10681 (N_10681,N_10332,N_10305);
and U10682 (N_10682,N_10412,N_10317);
xnor U10683 (N_10683,N_10326,N_10418);
nor U10684 (N_10684,N_10499,N_10408);
or U10685 (N_10685,N_10285,N_10323);
nor U10686 (N_10686,N_10287,N_10422);
xor U10687 (N_10687,N_10315,N_10382);
xnor U10688 (N_10688,N_10294,N_10293);
xnor U10689 (N_10689,N_10400,N_10417);
xor U10690 (N_10690,N_10397,N_10420);
nand U10691 (N_10691,N_10271,N_10405);
nand U10692 (N_10692,N_10303,N_10299);
nand U10693 (N_10693,N_10369,N_10262);
xnor U10694 (N_10694,N_10312,N_10394);
nand U10695 (N_10695,N_10403,N_10269);
nor U10696 (N_10696,N_10380,N_10438);
and U10697 (N_10697,N_10390,N_10433);
or U10698 (N_10698,N_10319,N_10412);
nor U10699 (N_10699,N_10291,N_10428);
xnor U10700 (N_10700,N_10329,N_10489);
nand U10701 (N_10701,N_10251,N_10310);
or U10702 (N_10702,N_10428,N_10442);
nor U10703 (N_10703,N_10276,N_10355);
or U10704 (N_10704,N_10268,N_10266);
or U10705 (N_10705,N_10464,N_10357);
and U10706 (N_10706,N_10318,N_10374);
and U10707 (N_10707,N_10390,N_10254);
xnor U10708 (N_10708,N_10283,N_10358);
or U10709 (N_10709,N_10357,N_10388);
or U10710 (N_10710,N_10356,N_10457);
nor U10711 (N_10711,N_10272,N_10373);
nand U10712 (N_10712,N_10458,N_10439);
xor U10713 (N_10713,N_10435,N_10273);
xor U10714 (N_10714,N_10379,N_10276);
xnor U10715 (N_10715,N_10263,N_10353);
xor U10716 (N_10716,N_10304,N_10482);
nand U10717 (N_10717,N_10394,N_10470);
nor U10718 (N_10718,N_10324,N_10449);
nand U10719 (N_10719,N_10362,N_10403);
nor U10720 (N_10720,N_10279,N_10412);
xnor U10721 (N_10721,N_10485,N_10360);
xor U10722 (N_10722,N_10318,N_10473);
or U10723 (N_10723,N_10434,N_10488);
and U10724 (N_10724,N_10254,N_10417);
nand U10725 (N_10725,N_10291,N_10383);
and U10726 (N_10726,N_10414,N_10317);
xnor U10727 (N_10727,N_10377,N_10440);
xnor U10728 (N_10728,N_10420,N_10315);
or U10729 (N_10729,N_10408,N_10435);
nand U10730 (N_10730,N_10404,N_10481);
or U10731 (N_10731,N_10283,N_10263);
or U10732 (N_10732,N_10432,N_10324);
nand U10733 (N_10733,N_10468,N_10449);
nand U10734 (N_10734,N_10275,N_10450);
xnor U10735 (N_10735,N_10373,N_10285);
nor U10736 (N_10736,N_10491,N_10371);
or U10737 (N_10737,N_10418,N_10275);
nand U10738 (N_10738,N_10334,N_10399);
or U10739 (N_10739,N_10362,N_10457);
and U10740 (N_10740,N_10324,N_10313);
nand U10741 (N_10741,N_10280,N_10336);
nor U10742 (N_10742,N_10278,N_10399);
xor U10743 (N_10743,N_10465,N_10397);
xnor U10744 (N_10744,N_10369,N_10327);
nor U10745 (N_10745,N_10270,N_10482);
or U10746 (N_10746,N_10387,N_10482);
or U10747 (N_10747,N_10268,N_10409);
or U10748 (N_10748,N_10427,N_10482);
nand U10749 (N_10749,N_10358,N_10491);
nor U10750 (N_10750,N_10509,N_10654);
nand U10751 (N_10751,N_10727,N_10650);
xnor U10752 (N_10752,N_10596,N_10632);
and U10753 (N_10753,N_10630,N_10656);
nand U10754 (N_10754,N_10700,N_10637);
xor U10755 (N_10755,N_10663,N_10601);
nand U10756 (N_10756,N_10728,N_10722);
nor U10757 (N_10757,N_10502,N_10693);
nor U10758 (N_10758,N_10530,N_10683);
nand U10759 (N_10759,N_10746,N_10518);
and U10760 (N_10760,N_10730,N_10582);
and U10761 (N_10761,N_10735,N_10616);
or U10762 (N_10762,N_10617,N_10598);
xor U10763 (N_10763,N_10606,N_10723);
and U10764 (N_10764,N_10521,N_10576);
and U10765 (N_10765,N_10716,N_10622);
nor U10766 (N_10766,N_10652,N_10563);
nand U10767 (N_10767,N_10707,N_10545);
and U10768 (N_10768,N_10520,N_10741);
or U10769 (N_10769,N_10548,N_10615);
and U10770 (N_10770,N_10748,N_10558);
nor U10771 (N_10771,N_10564,N_10519);
xnor U10772 (N_10772,N_10666,N_10568);
and U10773 (N_10773,N_10706,N_10685);
nand U10774 (N_10774,N_10638,N_10523);
nor U10775 (N_10775,N_10710,N_10726);
xnor U10776 (N_10776,N_10613,N_10567);
nand U10777 (N_10777,N_10584,N_10665);
xor U10778 (N_10778,N_10745,N_10577);
and U10779 (N_10779,N_10697,N_10543);
nor U10780 (N_10780,N_10633,N_10549);
and U10781 (N_10781,N_10565,N_10566);
nor U10782 (N_10782,N_10588,N_10668);
nand U10783 (N_10783,N_10537,N_10614);
nand U10784 (N_10784,N_10525,N_10714);
and U10785 (N_10785,N_10609,N_10587);
or U10786 (N_10786,N_10699,N_10736);
xor U10787 (N_10787,N_10590,N_10725);
xnor U10788 (N_10788,N_10667,N_10634);
nor U10789 (N_10789,N_10661,N_10738);
nor U10790 (N_10790,N_10664,N_10692);
nand U10791 (N_10791,N_10660,N_10522);
xor U10792 (N_10792,N_10625,N_10684);
and U10793 (N_10793,N_10734,N_10635);
or U10794 (N_10794,N_10554,N_10593);
or U10795 (N_10795,N_10508,N_10511);
xnor U10796 (N_10796,N_10611,N_10573);
nand U10797 (N_10797,N_10680,N_10636);
and U10798 (N_10798,N_10688,N_10533);
or U10799 (N_10799,N_10704,N_10690);
and U10800 (N_10800,N_10505,N_10708);
and U10801 (N_10801,N_10687,N_10541);
nor U10802 (N_10802,N_10709,N_10589);
or U10803 (N_10803,N_10737,N_10662);
nor U10804 (N_10804,N_10671,N_10631);
or U10805 (N_10805,N_10569,N_10628);
nand U10806 (N_10806,N_10643,N_10619);
nand U10807 (N_10807,N_10642,N_10743);
nor U10808 (N_10808,N_10645,N_10550);
nor U10809 (N_10809,N_10552,N_10527);
or U10810 (N_10810,N_10681,N_10560);
and U10811 (N_10811,N_10653,N_10695);
xnor U10812 (N_10812,N_10592,N_10513);
nand U10813 (N_10813,N_10618,N_10682);
or U10814 (N_10814,N_10649,N_10532);
nand U10815 (N_10815,N_10524,N_10719);
nand U10816 (N_10816,N_10534,N_10640);
nor U10817 (N_10817,N_10526,N_10544);
nand U10818 (N_10818,N_10540,N_10585);
xnor U10819 (N_10819,N_10657,N_10651);
xor U10820 (N_10820,N_10574,N_10639);
nand U10821 (N_10821,N_10553,N_10712);
or U10822 (N_10822,N_10749,N_10506);
nor U10823 (N_10823,N_10655,N_10612);
nor U10824 (N_10824,N_10648,N_10731);
xnor U10825 (N_10825,N_10627,N_10696);
nand U10826 (N_10826,N_10647,N_10594);
nand U10827 (N_10827,N_10512,N_10705);
nand U10828 (N_10828,N_10501,N_10604);
xnor U10829 (N_10829,N_10718,N_10547);
nand U10830 (N_10830,N_10583,N_10691);
or U10831 (N_10831,N_10602,N_10717);
xnor U10832 (N_10832,N_10703,N_10620);
nand U10833 (N_10833,N_10535,N_10621);
or U10834 (N_10834,N_10644,N_10739);
or U10835 (N_10835,N_10675,N_10733);
or U10836 (N_10836,N_10581,N_10740);
xor U10837 (N_10837,N_10546,N_10686);
and U10838 (N_10838,N_10579,N_10729);
and U10839 (N_10839,N_10603,N_10698);
nand U10840 (N_10840,N_10669,N_10597);
xor U10841 (N_10841,N_10559,N_10595);
xor U10842 (N_10842,N_10561,N_10702);
or U10843 (N_10843,N_10721,N_10676);
nand U10844 (N_10844,N_10711,N_10673);
xor U10845 (N_10845,N_10591,N_10542);
or U10846 (N_10846,N_10578,N_10529);
or U10847 (N_10847,N_10551,N_10677);
or U10848 (N_10848,N_10580,N_10678);
nand U10849 (N_10849,N_10538,N_10646);
xor U10850 (N_10850,N_10624,N_10742);
xnor U10851 (N_10851,N_10605,N_10510);
nor U10852 (N_10852,N_10747,N_10629);
nand U10853 (N_10853,N_10623,N_10572);
xor U10854 (N_10854,N_10575,N_10528);
nor U10855 (N_10855,N_10536,N_10500);
or U10856 (N_10856,N_10608,N_10556);
and U10857 (N_10857,N_10570,N_10599);
nor U10858 (N_10858,N_10713,N_10600);
or U10859 (N_10859,N_10586,N_10715);
nand U10860 (N_10860,N_10503,N_10571);
and U10861 (N_10861,N_10607,N_10514);
nand U10862 (N_10862,N_10557,N_10517);
xnor U10863 (N_10863,N_10659,N_10679);
nand U10864 (N_10864,N_10626,N_10724);
and U10865 (N_10865,N_10610,N_10531);
and U10866 (N_10866,N_10689,N_10504);
nor U10867 (N_10867,N_10516,N_10539);
nand U10868 (N_10868,N_10515,N_10641);
or U10869 (N_10869,N_10507,N_10720);
xor U10870 (N_10870,N_10562,N_10732);
nor U10871 (N_10871,N_10701,N_10670);
or U10872 (N_10872,N_10744,N_10555);
nor U10873 (N_10873,N_10672,N_10694);
xnor U10874 (N_10874,N_10674,N_10658);
nor U10875 (N_10875,N_10595,N_10511);
nand U10876 (N_10876,N_10601,N_10619);
nor U10877 (N_10877,N_10624,N_10589);
nand U10878 (N_10878,N_10616,N_10632);
xnor U10879 (N_10879,N_10592,N_10736);
nor U10880 (N_10880,N_10632,N_10608);
nand U10881 (N_10881,N_10572,N_10621);
and U10882 (N_10882,N_10521,N_10656);
nor U10883 (N_10883,N_10546,N_10676);
or U10884 (N_10884,N_10611,N_10729);
xnor U10885 (N_10885,N_10559,N_10536);
xor U10886 (N_10886,N_10600,N_10632);
or U10887 (N_10887,N_10712,N_10648);
or U10888 (N_10888,N_10646,N_10711);
and U10889 (N_10889,N_10581,N_10530);
or U10890 (N_10890,N_10617,N_10694);
nor U10891 (N_10891,N_10575,N_10560);
nor U10892 (N_10892,N_10547,N_10721);
nor U10893 (N_10893,N_10537,N_10749);
xor U10894 (N_10894,N_10641,N_10526);
and U10895 (N_10895,N_10665,N_10541);
or U10896 (N_10896,N_10688,N_10623);
nor U10897 (N_10897,N_10533,N_10693);
nand U10898 (N_10898,N_10542,N_10681);
nand U10899 (N_10899,N_10641,N_10669);
nand U10900 (N_10900,N_10509,N_10740);
xnor U10901 (N_10901,N_10636,N_10664);
nor U10902 (N_10902,N_10728,N_10547);
nand U10903 (N_10903,N_10506,N_10643);
and U10904 (N_10904,N_10618,N_10538);
nand U10905 (N_10905,N_10521,N_10584);
or U10906 (N_10906,N_10516,N_10633);
or U10907 (N_10907,N_10582,N_10643);
nand U10908 (N_10908,N_10699,N_10747);
xor U10909 (N_10909,N_10717,N_10595);
or U10910 (N_10910,N_10656,N_10579);
xnor U10911 (N_10911,N_10667,N_10745);
nor U10912 (N_10912,N_10536,N_10667);
xnor U10913 (N_10913,N_10555,N_10718);
nand U10914 (N_10914,N_10619,N_10625);
or U10915 (N_10915,N_10661,N_10601);
nor U10916 (N_10916,N_10628,N_10523);
nand U10917 (N_10917,N_10712,N_10556);
nand U10918 (N_10918,N_10692,N_10549);
or U10919 (N_10919,N_10603,N_10655);
xor U10920 (N_10920,N_10601,N_10568);
xnor U10921 (N_10921,N_10614,N_10638);
or U10922 (N_10922,N_10558,N_10650);
xor U10923 (N_10923,N_10642,N_10547);
nand U10924 (N_10924,N_10505,N_10718);
or U10925 (N_10925,N_10529,N_10672);
nor U10926 (N_10926,N_10601,N_10611);
or U10927 (N_10927,N_10613,N_10591);
xnor U10928 (N_10928,N_10647,N_10563);
nor U10929 (N_10929,N_10535,N_10522);
and U10930 (N_10930,N_10608,N_10714);
or U10931 (N_10931,N_10702,N_10570);
or U10932 (N_10932,N_10507,N_10673);
or U10933 (N_10933,N_10739,N_10681);
nand U10934 (N_10934,N_10671,N_10519);
nor U10935 (N_10935,N_10565,N_10629);
nand U10936 (N_10936,N_10737,N_10576);
and U10937 (N_10937,N_10639,N_10626);
nand U10938 (N_10938,N_10550,N_10663);
xnor U10939 (N_10939,N_10599,N_10736);
nand U10940 (N_10940,N_10592,N_10704);
nand U10941 (N_10941,N_10544,N_10513);
and U10942 (N_10942,N_10566,N_10560);
or U10943 (N_10943,N_10511,N_10533);
nor U10944 (N_10944,N_10610,N_10517);
nand U10945 (N_10945,N_10565,N_10542);
nor U10946 (N_10946,N_10716,N_10709);
nand U10947 (N_10947,N_10636,N_10502);
nand U10948 (N_10948,N_10663,N_10688);
nand U10949 (N_10949,N_10709,N_10689);
xor U10950 (N_10950,N_10543,N_10500);
and U10951 (N_10951,N_10686,N_10671);
or U10952 (N_10952,N_10681,N_10647);
or U10953 (N_10953,N_10618,N_10600);
nor U10954 (N_10954,N_10506,N_10636);
and U10955 (N_10955,N_10714,N_10609);
xor U10956 (N_10956,N_10521,N_10581);
nor U10957 (N_10957,N_10736,N_10545);
or U10958 (N_10958,N_10585,N_10528);
xnor U10959 (N_10959,N_10638,N_10630);
and U10960 (N_10960,N_10725,N_10675);
and U10961 (N_10961,N_10746,N_10542);
nor U10962 (N_10962,N_10511,N_10550);
and U10963 (N_10963,N_10743,N_10676);
nor U10964 (N_10964,N_10543,N_10638);
nand U10965 (N_10965,N_10540,N_10688);
or U10966 (N_10966,N_10577,N_10547);
xnor U10967 (N_10967,N_10579,N_10738);
and U10968 (N_10968,N_10675,N_10615);
nand U10969 (N_10969,N_10534,N_10695);
nand U10970 (N_10970,N_10506,N_10726);
nand U10971 (N_10971,N_10602,N_10710);
or U10972 (N_10972,N_10520,N_10708);
and U10973 (N_10973,N_10505,N_10517);
nor U10974 (N_10974,N_10562,N_10622);
and U10975 (N_10975,N_10530,N_10569);
xnor U10976 (N_10976,N_10531,N_10592);
nand U10977 (N_10977,N_10541,N_10572);
and U10978 (N_10978,N_10729,N_10665);
or U10979 (N_10979,N_10599,N_10609);
and U10980 (N_10980,N_10686,N_10568);
and U10981 (N_10981,N_10549,N_10589);
or U10982 (N_10982,N_10700,N_10581);
xnor U10983 (N_10983,N_10719,N_10609);
xor U10984 (N_10984,N_10606,N_10704);
or U10985 (N_10985,N_10744,N_10515);
nor U10986 (N_10986,N_10525,N_10737);
xor U10987 (N_10987,N_10689,N_10565);
and U10988 (N_10988,N_10549,N_10675);
nand U10989 (N_10989,N_10508,N_10611);
and U10990 (N_10990,N_10615,N_10659);
and U10991 (N_10991,N_10611,N_10516);
or U10992 (N_10992,N_10678,N_10589);
nor U10993 (N_10993,N_10664,N_10639);
or U10994 (N_10994,N_10559,N_10720);
xor U10995 (N_10995,N_10514,N_10596);
nor U10996 (N_10996,N_10710,N_10723);
or U10997 (N_10997,N_10556,N_10668);
and U10998 (N_10998,N_10537,N_10534);
or U10999 (N_10999,N_10550,N_10680);
or U11000 (N_11000,N_10802,N_10780);
nand U11001 (N_11001,N_10821,N_10874);
nor U11002 (N_11002,N_10972,N_10947);
or U11003 (N_11003,N_10966,N_10978);
or U11004 (N_11004,N_10960,N_10888);
nor U11005 (N_11005,N_10954,N_10827);
nor U11006 (N_11006,N_10863,N_10779);
nor U11007 (N_11007,N_10769,N_10828);
or U11008 (N_11008,N_10886,N_10813);
nand U11009 (N_11009,N_10911,N_10762);
nor U11010 (N_11010,N_10822,N_10905);
and U11011 (N_11011,N_10868,N_10943);
nand U11012 (N_11012,N_10935,N_10789);
nand U11013 (N_11013,N_10936,N_10791);
xor U11014 (N_11014,N_10852,N_10873);
nand U11015 (N_11015,N_10851,N_10800);
and U11016 (N_11016,N_10837,N_10958);
or U11017 (N_11017,N_10765,N_10910);
xnor U11018 (N_11018,N_10806,N_10914);
or U11019 (N_11019,N_10767,N_10871);
nor U11020 (N_11020,N_10772,N_10781);
nor U11021 (N_11021,N_10901,N_10792);
nor U11022 (N_11022,N_10809,N_10866);
or U11023 (N_11023,N_10971,N_10816);
xnor U11024 (N_11024,N_10934,N_10766);
nor U11025 (N_11025,N_10782,N_10930);
xnor U11026 (N_11026,N_10788,N_10758);
or U11027 (N_11027,N_10970,N_10784);
and U11028 (N_11028,N_10992,N_10820);
nor U11029 (N_11029,N_10961,N_10949);
and U11030 (N_11030,N_10962,N_10754);
or U11031 (N_11031,N_10778,N_10948);
or U11032 (N_11032,N_10804,N_10940);
nand U11033 (N_11033,N_10869,N_10879);
xnor U11034 (N_11034,N_10959,N_10920);
nand U11035 (N_11035,N_10773,N_10944);
or U11036 (N_11036,N_10927,N_10897);
nor U11037 (N_11037,N_10808,N_10892);
or U11038 (N_11038,N_10835,N_10777);
nand U11039 (N_11039,N_10753,N_10755);
or U11040 (N_11040,N_10880,N_10933);
nor U11041 (N_11041,N_10896,N_10803);
xor U11042 (N_11042,N_10975,N_10845);
xor U11043 (N_11043,N_10951,N_10801);
and U11044 (N_11044,N_10928,N_10774);
and U11045 (N_11045,N_10977,N_10841);
nor U11046 (N_11046,N_10831,N_10840);
and U11047 (N_11047,N_10956,N_10775);
nor U11048 (N_11048,N_10955,N_10846);
xor U11049 (N_11049,N_10854,N_10924);
and U11050 (N_11050,N_10946,N_10857);
xor U11051 (N_11051,N_10937,N_10786);
xor U11052 (N_11052,N_10993,N_10756);
nand U11053 (N_11053,N_10922,N_10923);
nand U11054 (N_11054,N_10843,N_10858);
nand U11055 (N_11055,N_10900,N_10825);
nand U11056 (N_11056,N_10763,N_10995);
or U11057 (N_11057,N_10895,N_10760);
and U11058 (N_11058,N_10872,N_10881);
nor U11059 (N_11059,N_10997,N_10771);
nor U11060 (N_11060,N_10824,N_10941);
xnor U11061 (N_11061,N_10985,N_10893);
nor U11062 (N_11062,N_10898,N_10829);
and U11063 (N_11063,N_10987,N_10797);
nand U11064 (N_11064,N_10812,N_10850);
xnor U11065 (N_11065,N_10832,N_10902);
or U11066 (N_11066,N_10885,N_10776);
nor U11067 (N_11067,N_10899,N_10830);
nor U11068 (N_11068,N_10810,N_10826);
or U11069 (N_11069,N_10882,N_10976);
xnor U11070 (N_11070,N_10847,N_10844);
nand U11071 (N_11071,N_10834,N_10968);
nand U11072 (N_11072,N_10906,N_10998);
or U11073 (N_11073,N_10999,N_10926);
or U11074 (N_11074,N_10953,N_10918);
or U11075 (N_11075,N_10790,N_10921);
or U11076 (N_11076,N_10761,N_10931);
or U11077 (N_11077,N_10982,N_10836);
xor U11078 (N_11078,N_10752,N_10853);
or U11079 (N_11079,N_10981,N_10796);
nor U11080 (N_11080,N_10856,N_10963);
nand U11081 (N_11081,N_10991,N_10855);
xnor U11082 (N_11082,N_10979,N_10864);
or U11083 (N_11083,N_10793,N_10913);
and U11084 (N_11084,N_10823,N_10915);
or U11085 (N_11085,N_10795,N_10964);
nand U11086 (N_11086,N_10884,N_10785);
or U11087 (N_11087,N_10794,N_10870);
nand U11088 (N_11088,N_10818,N_10988);
nand U11089 (N_11089,N_10942,N_10890);
and U11090 (N_11090,N_10807,N_10996);
or U11091 (N_11091,N_10757,N_10908);
and U11092 (N_11092,N_10903,N_10783);
nor U11093 (N_11093,N_10887,N_10990);
nand U11094 (N_11094,N_10878,N_10967);
nor U11095 (N_11095,N_10939,N_10994);
and U11096 (N_11096,N_10877,N_10799);
nand U11097 (N_11097,N_10919,N_10815);
nand U11098 (N_11098,N_10833,N_10989);
nand U11099 (N_11099,N_10945,N_10787);
or U11100 (N_11100,N_10980,N_10865);
or U11101 (N_11101,N_10805,N_10969);
nand U11102 (N_11102,N_10965,N_10986);
xnor U11103 (N_11103,N_10875,N_10848);
nand U11104 (N_11104,N_10932,N_10952);
nand U11105 (N_11105,N_10889,N_10819);
nor U11106 (N_11106,N_10891,N_10811);
nor U11107 (N_11107,N_10912,N_10751);
and U11108 (N_11108,N_10859,N_10907);
nor U11109 (N_11109,N_10957,N_10984);
xnor U11110 (N_11110,N_10838,N_10814);
nor U11111 (N_11111,N_10867,N_10938);
and U11112 (N_11112,N_10917,N_10876);
nand U11113 (N_11113,N_10770,N_10916);
nand U11114 (N_11114,N_10839,N_10861);
nand U11115 (N_11115,N_10849,N_10983);
or U11116 (N_11116,N_10909,N_10842);
or U11117 (N_11117,N_10950,N_10860);
nor U11118 (N_11118,N_10929,N_10798);
nand U11119 (N_11119,N_10764,N_10904);
xnor U11120 (N_11120,N_10925,N_10768);
or U11121 (N_11121,N_10894,N_10817);
or U11122 (N_11122,N_10974,N_10883);
nor U11123 (N_11123,N_10759,N_10973);
and U11124 (N_11124,N_10862,N_10750);
nor U11125 (N_11125,N_10815,N_10877);
nand U11126 (N_11126,N_10870,N_10961);
and U11127 (N_11127,N_10937,N_10771);
xnor U11128 (N_11128,N_10954,N_10856);
nor U11129 (N_11129,N_10751,N_10872);
or U11130 (N_11130,N_10978,N_10800);
or U11131 (N_11131,N_10948,N_10974);
nor U11132 (N_11132,N_10897,N_10919);
xnor U11133 (N_11133,N_10973,N_10958);
and U11134 (N_11134,N_10807,N_10887);
nor U11135 (N_11135,N_10924,N_10977);
xor U11136 (N_11136,N_10914,N_10792);
or U11137 (N_11137,N_10816,N_10857);
and U11138 (N_11138,N_10970,N_10920);
nand U11139 (N_11139,N_10876,N_10856);
nand U11140 (N_11140,N_10861,N_10867);
and U11141 (N_11141,N_10952,N_10950);
and U11142 (N_11142,N_10865,N_10796);
nand U11143 (N_11143,N_10954,N_10821);
or U11144 (N_11144,N_10876,N_10830);
or U11145 (N_11145,N_10752,N_10779);
nand U11146 (N_11146,N_10902,N_10980);
nor U11147 (N_11147,N_10793,N_10880);
xor U11148 (N_11148,N_10768,N_10897);
or U11149 (N_11149,N_10787,N_10808);
nand U11150 (N_11150,N_10833,N_10755);
nor U11151 (N_11151,N_10817,N_10997);
xor U11152 (N_11152,N_10795,N_10846);
and U11153 (N_11153,N_10912,N_10879);
nand U11154 (N_11154,N_10925,N_10848);
nor U11155 (N_11155,N_10808,N_10952);
xor U11156 (N_11156,N_10830,N_10924);
nor U11157 (N_11157,N_10917,N_10891);
xor U11158 (N_11158,N_10893,N_10873);
xor U11159 (N_11159,N_10784,N_10873);
nor U11160 (N_11160,N_10837,N_10954);
and U11161 (N_11161,N_10867,N_10907);
xnor U11162 (N_11162,N_10865,N_10911);
or U11163 (N_11163,N_10907,N_10755);
and U11164 (N_11164,N_10815,N_10807);
xor U11165 (N_11165,N_10821,N_10834);
xnor U11166 (N_11166,N_10814,N_10953);
and U11167 (N_11167,N_10781,N_10998);
and U11168 (N_11168,N_10915,N_10862);
and U11169 (N_11169,N_10849,N_10937);
xnor U11170 (N_11170,N_10931,N_10804);
xnor U11171 (N_11171,N_10804,N_10951);
and U11172 (N_11172,N_10908,N_10864);
and U11173 (N_11173,N_10949,N_10810);
nand U11174 (N_11174,N_10837,N_10754);
nor U11175 (N_11175,N_10889,N_10981);
xor U11176 (N_11176,N_10797,N_10988);
or U11177 (N_11177,N_10777,N_10846);
xor U11178 (N_11178,N_10860,N_10772);
and U11179 (N_11179,N_10934,N_10977);
and U11180 (N_11180,N_10900,N_10997);
nand U11181 (N_11181,N_10934,N_10860);
or U11182 (N_11182,N_10882,N_10810);
and U11183 (N_11183,N_10899,N_10895);
or U11184 (N_11184,N_10899,N_10841);
nand U11185 (N_11185,N_10855,N_10950);
or U11186 (N_11186,N_10970,N_10971);
xor U11187 (N_11187,N_10819,N_10949);
xnor U11188 (N_11188,N_10980,N_10897);
or U11189 (N_11189,N_10930,N_10901);
and U11190 (N_11190,N_10843,N_10900);
xnor U11191 (N_11191,N_10833,N_10812);
or U11192 (N_11192,N_10851,N_10761);
nand U11193 (N_11193,N_10915,N_10852);
xor U11194 (N_11194,N_10866,N_10796);
nor U11195 (N_11195,N_10773,N_10931);
nand U11196 (N_11196,N_10825,N_10758);
nand U11197 (N_11197,N_10762,N_10934);
or U11198 (N_11198,N_10949,N_10875);
and U11199 (N_11199,N_10952,N_10978);
or U11200 (N_11200,N_10753,N_10935);
and U11201 (N_11201,N_10817,N_10991);
xnor U11202 (N_11202,N_10788,N_10838);
nor U11203 (N_11203,N_10787,N_10977);
nor U11204 (N_11204,N_10765,N_10943);
or U11205 (N_11205,N_10961,N_10832);
nor U11206 (N_11206,N_10878,N_10846);
nor U11207 (N_11207,N_10980,N_10890);
or U11208 (N_11208,N_10974,N_10922);
or U11209 (N_11209,N_10847,N_10854);
nor U11210 (N_11210,N_10891,N_10885);
nand U11211 (N_11211,N_10921,N_10819);
nand U11212 (N_11212,N_10790,N_10959);
nand U11213 (N_11213,N_10833,N_10841);
and U11214 (N_11214,N_10968,N_10765);
nor U11215 (N_11215,N_10806,N_10850);
and U11216 (N_11216,N_10852,N_10790);
or U11217 (N_11217,N_10959,N_10967);
nand U11218 (N_11218,N_10981,N_10759);
nand U11219 (N_11219,N_10856,N_10941);
and U11220 (N_11220,N_10874,N_10851);
and U11221 (N_11221,N_10896,N_10810);
nand U11222 (N_11222,N_10939,N_10803);
nand U11223 (N_11223,N_10796,N_10803);
or U11224 (N_11224,N_10934,N_10819);
nor U11225 (N_11225,N_10786,N_10842);
nand U11226 (N_11226,N_10889,N_10772);
or U11227 (N_11227,N_10943,N_10763);
nor U11228 (N_11228,N_10756,N_10936);
xor U11229 (N_11229,N_10954,N_10977);
nand U11230 (N_11230,N_10880,N_10847);
or U11231 (N_11231,N_10838,N_10810);
xor U11232 (N_11232,N_10861,N_10855);
nand U11233 (N_11233,N_10913,N_10962);
xnor U11234 (N_11234,N_10785,N_10858);
and U11235 (N_11235,N_10765,N_10868);
nor U11236 (N_11236,N_10782,N_10895);
nand U11237 (N_11237,N_10813,N_10903);
or U11238 (N_11238,N_10918,N_10903);
nor U11239 (N_11239,N_10882,N_10787);
xor U11240 (N_11240,N_10970,N_10867);
nor U11241 (N_11241,N_10767,N_10913);
nor U11242 (N_11242,N_10897,N_10888);
xnor U11243 (N_11243,N_10786,N_10851);
nor U11244 (N_11244,N_10828,N_10895);
nor U11245 (N_11245,N_10912,N_10904);
nor U11246 (N_11246,N_10804,N_10917);
nand U11247 (N_11247,N_10848,N_10919);
or U11248 (N_11248,N_10858,N_10996);
and U11249 (N_11249,N_10873,N_10992);
nor U11250 (N_11250,N_11123,N_11128);
xor U11251 (N_11251,N_11007,N_11178);
nor U11252 (N_11252,N_11088,N_11195);
or U11253 (N_11253,N_11192,N_11236);
and U11254 (N_11254,N_11229,N_11155);
or U11255 (N_11255,N_11005,N_11147);
nor U11256 (N_11256,N_11230,N_11019);
and U11257 (N_11257,N_11196,N_11182);
and U11258 (N_11258,N_11074,N_11045);
nand U11259 (N_11259,N_11145,N_11190);
or U11260 (N_11260,N_11063,N_11110);
xnor U11261 (N_11261,N_11030,N_11079);
nand U11262 (N_11262,N_11012,N_11173);
nand U11263 (N_11263,N_11223,N_11218);
and U11264 (N_11264,N_11133,N_11002);
xor U11265 (N_11265,N_11070,N_11058);
or U11266 (N_11266,N_11086,N_11177);
nand U11267 (N_11267,N_11038,N_11067);
nand U11268 (N_11268,N_11206,N_11244);
nand U11269 (N_11269,N_11227,N_11224);
nand U11270 (N_11270,N_11141,N_11150);
and U11271 (N_11271,N_11017,N_11109);
nand U11272 (N_11272,N_11202,N_11097);
nor U11273 (N_11273,N_11162,N_11077);
nand U11274 (N_11274,N_11127,N_11120);
nand U11275 (N_11275,N_11129,N_11132);
nor U11276 (N_11276,N_11217,N_11095);
nor U11277 (N_11277,N_11170,N_11199);
nor U11278 (N_11278,N_11146,N_11083);
or U11279 (N_11279,N_11187,N_11093);
and U11280 (N_11280,N_11204,N_11113);
xnor U11281 (N_11281,N_11158,N_11241);
nand U11282 (N_11282,N_11062,N_11025);
or U11283 (N_11283,N_11137,N_11075);
nor U11284 (N_11284,N_11211,N_11131);
or U11285 (N_11285,N_11050,N_11144);
nor U11286 (N_11286,N_11048,N_11176);
or U11287 (N_11287,N_11189,N_11152);
nor U11288 (N_11288,N_11232,N_11226);
and U11289 (N_11289,N_11210,N_11043);
nor U11290 (N_11290,N_11186,N_11164);
or U11291 (N_11291,N_11175,N_11034);
and U11292 (N_11292,N_11234,N_11157);
or U11293 (N_11293,N_11064,N_11087);
nor U11294 (N_11294,N_11181,N_11049);
nor U11295 (N_11295,N_11193,N_11011);
nand U11296 (N_11296,N_11082,N_11235);
nor U11297 (N_11297,N_11142,N_11015);
or U11298 (N_11298,N_11035,N_11054);
xnor U11299 (N_11299,N_11056,N_11108);
nor U11300 (N_11300,N_11243,N_11183);
xnor U11301 (N_11301,N_11040,N_11102);
nand U11302 (N_11302,N_11148,N_11208);
nor U11303 (N_11303,N_11174,N_11059);
nand U11304 (N_11304,N_11238,N_11167);
and U11305 (N_11305,N_11246,N_11140);
nor U11306 (N_11306,N_11160,N_11130);
or U11307 (N_11307,N_11159,N_11231);
nor U11308 (N_11308,N_11184,N_11008);
nor U11309 (N_11309,N_11249,N_11240);
xnor U11310 (N_11310,N_11004,N_11122);
and U11311 (N_11311,N_11239,N_11169);
or U11312 (N_11312,N_11091,N_11194);
nand U11313 (N_11313,N_11185,N_11242);
or U11314 (N_11314,N_11103,N_11151);
nand U11315 (N_11315,N_11046,N_11179);
nor U11316 (N_11316,N_11111,N_11221);
or U11317 (N_11317,N_11000,N_11018);
or U11318 (N_11318,N_11171,N_11166);
nor U11319 (N_11319,N_11135,N_11006);
and U11320 (N_11320,N_11247,N_11071);
nor U11321 (N_11321,N_11057,N_11220);
or U11322 (N_11322,N_11134,N_11037);
nand U11323 (N_11323,N_11115,N_11216);
xnor U11324 (N_11324,N_11219,N_11016);
and U11325 (N_11325,N_11112,N_11089);
nor U11326 (N_11326,N_11069,N_11020);
or U11327 (N_11327,N_11248,N_11154);
xnor U11328 (N_11328,N_11201,N_11022);
nand U11329 (N_11329,N_11098,N_11096);
nand U11330 (N_11330,N_11126,N_11139);
nand U11331 (N_11331,N_11027,N_11153);
xnor U11332 (N_11332,N_11014,N_11191);
nand U11333 (N_11333,N_11041,N_11081);
nand U11334 (N_11334,N_11055,N_11036);
and U11335 (N_11335,N_11117,N_11149);
and U11336 (N_11336,N_11010,N_11053);
xor U11337 (N_11337,N_11031,N_11104);
nand U11338 (N_11338,N_11094,N_11084);
xnor U11339 (N_11339,N_11068,N_11021);
nand U11340 (N_11340,N_11228,N_11033);
nand U11341 (N_11341,N_11119,N_11090);
nand U11342 (N_11342,N_11209,N_11163);
and U11343 (N_11343,N_11052,N_11051);
nor U11344 (N_11344,N_11107,N_11165);
nand U11345 (N_11345,N_11101,N_11197);
and U11346 (N_11346,N_11013,N_11207);
and U11347 (N_11347,N_11225,N_11237);
xor U11348 (N_11348,N_11042,N_11125);
nand U11349 (N_11349,N_11124,N_11214);
xnor U11350 (N_11350,N_11203,N_11001);
xnor U11351 (N_11351,N_11143,N_11072);
nor U11352 (N_11352,N_11205,N_11039);
nor U11353 (N_11353,N_11100,N_11136);
or U11354 (N_11354,N_11023,N_11121);
xnor U11355 (N_11355,N_11073,N_11114);
and U11356 (N_11356,N_11106,N_11061);
and U11357 (N_11357,N_11105,N_11212);
or U11358 (N_11358,N_11078,N_11080);
nand U11359 (N_11359,N_11116,N_11076);
nor U11360 (N_11360,N_11180,N_11060);
or U11361 (N_11361,N_11138,N_11198);
and U11362 (N_11362,N_11065,N_11029);
nor U11363 (N_11363,N_11222,N_11233);
nor U11364 (N_11364,N_11003,N_11009);
and U11365 (N_11365,N_11032,N_11085);
nor U11366 (N_11366,N_11024,N_11245);
nor U11367 (N_11367,N_11026,N_11188);
and U11368 (N_11368,N_11044,N_11118);
or U11369 (N_11369,N_11047,N_11213);
nor U11370 (N_11370,N_11172,N_11099);
nand U11371 (N_11371,N_11168,N_11066);
or U11372 (N_11372,N_11161,N_11028);
nor U11373 (N_11373,N_11215,N_11156);
and U11374 (N_11374,N_11092,N_11200);
and U11375 (N_11375,N_11079,N_11171);
and U11376 (N_11376,N_11087,N_11204);
nand U11377 (N_11377,N_11152,N_11195);
nand U11378 (N_11378,N_11197,N_11133);
and U11379 (N_11379,N_11123,N_11174);
or U11380 (N_11380,N_11015,N_11140);
xor U11381 (N_11381,N_11052,N_11188);
nor U11382 (N_11382,N_11164,N_11050);
nand U11383 (N_11383,N_11202,N_11078);
nor U11384 (N_11384,N_11003,N_11195);
nor U11385 (N_11385,N_11217,N_11228);
and U11386 (N_11386,N_11047,N_11187);
xnor U11387 (N_11387,N_11205,N_11019);
nand U11388 (N_11388,N_11015,N_11106);
or U11389 (N_11389,N_11187,N_11162);
xnor U11390 (N_11390,N_11191,N_11113);
and U11391 (N_11391,N_11036,N_11053);
xor U11392 (N_11392,N_11249,N_11188);
nand U11393 (N_11393,N_11223,N_11137);
nand U11394 (N_11394,N_11026,N_11033);
nor U11395 (N_11395,N_11137,N_11076);
xnor U11396 (N_11396,N_11218,N_11092);
nor U11397 (N_11397,N_11203,N_11110);
and U11398 (N_11398,N_11036,N_11245);
or U11399 (N_11399,N_11103,N_11100);
nand U11400 (N_11400,N_11191,N_11100);
nor U11401 (N_11401,N_11132,N_11081);
or U11402 (N_11402,N_11081,N_11236);
nor U11403 (N_11403,N_11105,N_11010);
or U11404 (N_11404,N_11112,N_11186);
nor U11405 (N_11405,N_11082,N_11091);
nor U11406 (N_11406,N_11099,N_11153);
and U11407 (N_11407,N_11248,N_11037);
or U11408 (N_11408,N_11141,N_11168);
or U11409 (N_11409,N_11164,N_11020);
nor U11410 (N_11410,N_11120,N_11001);
nand U11411 (N_11411,N_11118,N_11242);
xnor U11412 (N_11412,N_11134,N_11044);
nand U11413 (N_11413,N_11002,N_11009);
and U11414 (N_11414,N_11047,N_11128);
and U11415 (N_11415,N_11050,N_11001);
nor U11416 (N_11416,N_11197,N_11001);
and U11417 (N_11417,N_11027,N_11056);
nor U11418 (N_11418,N_11186,N_11064);
nor U11419 (N_11419,N_11049,N_11200);
and U11420 (N_11420,N_11233,N_11106);
xor U11421 (N_11421,N_11204,N_11061);
or U11422 (N_11422,N_11242,N_11132);
xnor U11423 (N_11423,N_11060,N_11227);
nand U11424 (N_11424,N_11131,N_11102);
nand U11425 (N_11425,N_11182,N_11192);
or U11426 (N_11426,N_11045,N_11128);
or U11427 (N_11427,N_11160,N_11210);
nand U11428 (N_11428,N_11175,N_11003);
or U11429 (N_11429,N_11164,N_11143);
nand U11430 (N_11430,N_11157,N_11097);
xnor U11431 (N_11431,N_11096,N_11057);
nor U11432 (N_11432,N_11142,N_11074);
xor U11433 (N_11433,N_11137,N_11143);
nor U11434 (N_11434,N_11207,N_11049);
xor U11435 (N_11435,N_11079,N_11159);
nor U11436 (N_11436,N_11111,N_11162);
xnor U11437 (N_11437,N_11017,N_11073);
xor U11438 (N_11438,N_11065,N_11212);
or U11439 (N_11439,N_11058,N_11135);
nor U11440 (N_11440,N_11201,N_11075);
nor U11441 (N_11441,N_11141,N_11147);
and U11442 (N_11442,N_11127,N_11166);
nor U11443 (N_11443,N_11089,N_11118);
or U11444 (N_11444,N_11086,N_11230);
nand U11445 (N_11445,N_11245,N_11029);
nor U11446 (N_11446,N_11019,N_11111);
or U11447 (N_11447,N_11067,N_11202);
nor U11448 (N_11448,N_11137,N_11035);
nand U11449 (N_11449,N_11025,N_11063);
nor U11450 (N_11450,N_11046,N_11239);
nand U11451 (N_11451,N_11212,N_11010);
or U11452 (N_11452,N_11168,N_11163);
and U11453 (N_11453,N_11214,N_11149);
nor U11454 (N_11454,N_11105,N_11214);
xnor U11455 (N_11455,N_11198,N_11175);
nor U11456 (N_11456,N_11171,N_11225);
nand U11457 (N_11457,N_11098,N_11012);
nand U11458 (N_11458,N_11190,N_11170);
or U11459 (N_11459,N_11116,N_11135);
nand U11460 (N_11460,N_11142,N_11249);
nand U11461 (N_11461,N_11047,N_11186);
xor U11462 (N_11462,N_11129,N_11028);
nor U11463 (N_11463,N_11004,N_11029);
and U11464 (N_11464,N_11106,N_11096);
nor U11465 (N_11465,N_11089,N_11035);
nand U11466 (N_11466,N_11214,N_11234);
and U11467 (N_11467,N_11115,N_11036);
xor U11468 (N_11468,N_11218,N_11147);
and U11469 (N_11469,N_11233,N_11213);
nor U11470 (N_11470,N_11242,N_11096);
nand U11471 (N_11471,N_11228,N_11141);
or U11472 (N_11472,N_11117,N_11053);
or U11473 (N_11473,N_11191,N_11125);
and U11474 (N_11474,N_11128,N_11114);
nand U11475 (N_11475,N_11176,N_11215);
nor U11476 (N_11476,N_11132,N_11075);
or U11477 (N_11477,N_11105,N_11136);
or U11478 (N_11478,N_11219,N_11028);
xor U11479 (N_11479,N_11012,N_11193);
and U11480 (N_11480,N_11105,N_11167);
nor U11481 (N_11481,N_11215,N_11031);
nor U11482 (N_11482,N_11201,N_11157);
nand U11483 (N_11483,N_11032,N_11036);
and U11484 (N_11484,N_11008,N_11038);
nor U11485 (N_11485,N_11111,N_11117);
xnor U11486 (N_11486,N_11114,N_11224);
and U11487 (N_11487,N_11205,N_11086);
nor U11488 (N_11488,N_11073,N_11129);
and U11489 (N_11489,N_11123,N_11001);
and U11490 (N_11490,N_11160,N_11010);
nand U11491 (N_11491,N_11181,N_11237);
or U11492 (N_11492,N_11022,N_11044);
and U11493 (N_11493,N_11204,N_11011);
nand U11494 (N_11494,N_11181,N_11092);
or U11495 (N_11495,N_11245,N_11015);
and U11496 (N_11496,N_11111,N_11043);
nor U11497 (N_11497,N_11201,N_11211);
or U11498 (N_11498,N_11063,N_11068);
and U11499 (N_11499,N_11187,N_11212);
nor U11500 (N_11500,N_11262,N_11303);
and U11501 (N_11501,N_11486,N_11452);
or U11502 (N_11502,N_11320,N_11355);
and U11503 (N_11503,N_11354,N_11348);
nand U11504 (N_11504,N_11461,N_11498);
xnor U11505 (N_11505,N_11270,N_11383);
or U11506 (N_11506,N_11328,N_11479);
and U11507 (N_11507,N_11390,N_11329);
and U11508 (N_11508,N_11279,N_11424);
or U11509 (N_11509,N_11269,N_11305);
or U11510 (N_11510,N_11284,N_11398);
or U11511 (N_11511,N_11497,N_11457);
xnor U11512 (N_11512,N_11492,N_11381);
nand U11513 (N_11513,N_11473,N_11391);
nor U11514 (N_11514,N_11370,N_11451);
nand U11515 (N_11515,N_11433,N_11425);
or U11516 (N_11516,N_11322,N_11491);
or U11517 (N_11517,N_11293,N_11323);
xnor U11518 (N_11518,N_11394,N_11475);
xor U11519 (N_11519,N_11325,N_11476);
nor U11520 (N_11520,N_11306,N_11442);
nand U11521 (N_11521,N_11407,N_11487);
nand U11522 (N_11522,N_11488,N_11459);
or U11523 (N_11523,N_11256,N_11401);
nor U11524 (N_11524,N_11389,N_11330);
nand U11525 (N_11525,N_11312,N_11367);
nand U11526 (N_11526,N_11444,N_11404);
nand U11527 (N_11527,N_11335,N_11484);
nand U11528 (N_11528,N_11410,N_11400);
or U11529 (N_11529,N_11275,N_11485);
and U11530 (N_11530,N_11298,N_11291);
and U11531 (N_11531,N_11469,N_11481);
nand U11532 (N_11532,N_11336,N_11307);
and U11533 (N_11533,N_11326,N_11324);
or U11534 (N_11534,N_11439,N_11477);
xor U11535 (N_11535,N_11464,N_11447);
or U11536 (N_11536,N_11285,N_11357);
nor U11537 (N_11537,N_11358,N_11294);
nor U11538 (N_11538,N_11387,N_11392);
nor U11539 (N_11539,N_11490,N_11427);
xnor U11540 (N_11540,N_11482,N_11434);
xor U11541 (N_11541,N_11277,N_11265);
nand U11542 (N_11542,N_11345,N_11251);
or U11543 (N_11543,N_11397,N_11319);
nand U11544 (N_11544,N_11493,N_11409);
nand U11545 (N_11545,N_11454,N_11455);
and U11546 (N_11546,N_11456,N_11463);
nand U11547 (N_11547,N_11352,N_11347);
nor U11548 (N_11548,N_11449,N_11349);
nand U11549 (N_11549,N_11386,N_11418);
xor U11550 (N_11550,N_11467,N_11302);
and U11551 (N_11551,N_11308,N_11403);
nand U11552 (N_11552,N_11384,N_11458);
nor U11553 (N_11553,N_11268,N_11462);
and U11554 (N_11554,N_11402,N_11317);
nand U11555 (N_11555,N_11376,N_11252);
or U11556 (N_11556,N_11271,N_11263);
xnor U11557 (N_11557,N_11421,N_11304);
nand U11558 (N_11558,N_11261,N_11250);
and U11559 (N_11559,N_11411,N_11416);
nand U11560 (N_11560,N_11315,N_11286);
nor U11561 (N_11561,N_11369,N_11292);
nor U11562 (N_11562,N_11441,N_11267);
or U11563 (N_11563,N_11489,N_11373);
or U11564 (N_11564,N_11408,N_11273);
or U11565 (N_11565,N_11353,N_11350);
and U11566 (N_11566,N_11254,N_11295);
and U11567 (N_11567,N_11422,N_11260);
nand U11568 (N_11568,N_11280,N_11287);
and U11569 (N_11569,N_11382,N_11346);
or U11570 (N_11570,N_11496,N_11474);
nand U11571 (N_11571,N_11314,N_11344);
nor U11572 (N_11572,N_11316,N_11470);
and U11573 (N_11573,N_11289,N_11440);
nor U11574 (N_11574,N_11297,N_11412);
nor U11575 (N_11575,N_11415,N_11313);
xnor U11576 (N_11576,N_11374,N_11378);
and U11577 (N_11577,N_11342,N_11300);
xnor U11578 (N_11578,N_11311,N_11272);
and U11579 (N_11579,N_11423,N_11333);
nor U11580 (N_11580,N_11443,N_11274);
or U11581 (N_11581,N_11290,N_11362);
and U11582 (N_11582,N_11395,N_11377);
xnor U11583 (N_11583,N_11379,N_11436);
and U11584 (N_11584,N_11478,N_11366);
xor U11585 (N_11585,N_11253,N_11426);
xor U11586 (N_11586,N_11375,N_11446);
or U11587 (N_11587,N_11468,N_11417);
and U11588 (N_11588,N_11371,N_11399);
nand U11589 (N_11589,N_11343,N_11396);
and U11590 (N_11590,N_11419,N_11296);
xnor U11591 (N_11591,N_11445,N_11321);
xor U11592 (N_11592,N_11420,N_11495);
xor U11593 (N_11593,N_11299,N_11356);
xor U11594 (N_11594,N_11431,N_11310);
nor U11595 (N_11595,N_11483,N_11453);
and U11596 (N_11596,N_11282,N_11258);
xnor U11597 (N_11597,N_11332,N_11337);
xnor U11598 (N_11598,N_11435,N_11361);
nand U11599 (N_11599,N_11288,N_11494);
nand U11600 (N_11600,N_11359,N_11405);
nor U11601 (N_11601,N_11406,N_11365);
nand U11602 (N_11602,N_11429,N_11301);
nor U11603 (N_11603,N_11460,N_11372);
nor U11604 (N_11604,N_11428,N_11480);
or U11605 (N_11605,N_11341,N_11380);
or U11606 (N_11606,N_11472,N_11388);
nor U11607 (N_11607,N_11257,N_11499);
nor U11608 (N_11608,N_11334,N_11264);
or U11609 (N_11609,N_11327,N_11255);
or U11610 (N_11610,N_11331,N_11385);
and U11611 (N_11611,N_11339,N_11368);
xor U11612 (N_11612,N_11259,N_11414);
xor U11613 (N_11613,N_11471,N_11413);
nand U11614 (N_11614,N_11450,N_11276);
and U11615 (N_11615,N_11364,N_11318);
xor U11616 (N_11616,N_11466,N_11393);
nor U11617 (N_11617,N_11360,N_11338);
or U11618 (N_11618,N_11438,N_11363);
nor U11619 (N_11619,N_11465,N_11266);
nand U11620 (N_11620,N_11432,N_11309);
or U11621 (N_11621,N_11278,N_11351);
and U11622 (N_11622,N_11437,N_11340);
or U11623 (N_11623,N_11430,N_11283);
xnor U11624 (N_11624,N_11281,N_11448);
nand U11625 (N_11625,N_11428,N_11468);
or U11626 (N_11626,N_11488,N_11338);
nand U11627 (N_11627,N_11327,N_11443);
xor U11628 (N_11628,N_11269,N_11471);
or U11629 (N_11629,N_11477,N_11355);
xor U11630 (N_11630,N_11371,N_11424);
xnor U11631 (N_11631,N_11307,N_11357);
xnor U11632 (N_11632,N_11256,N_11311);
nand U11633 (N_11633,N_11371,N_11365);
nor U11634 (N_11634,N_11440,N_11344);
or U11635 (N_11635,N_11404,N_11488);
and U11636 (N_11636,N_11456,N_11368);
nor U11637 (N_11637,N_11320,N_11493);
xnor U11638 (N_11638,N_11344,N_11373);
or U11639 (N_11639,N_11340,N_11480);
nand U11640 (N_11640,N_11499,N_11379);
or U11641 (N_11641,N_11464,N_11310);
nor U11642 (N_11642,N_11302,N_11367);
and U11643 (N_11643,N_11412,N_11430);
and U11644 (N_11644,N_11351,N_11419);
nand U11645 (N_11645,N_11360,N_11380);
xor U11646 (N_11646,N_11303,N_11304);
nand U11647 (N_11647,N_11407,N_11292);
nor U11648 (N_11648,N_11448,N_11430);
and U11649 (N_11649,N_11394,N_11441);
nand U11650 (N_11650,N_11251,N_11471);
nand U11651 (N_11651,N_11320,N_11465);
and U11652 (N_11652,N_11481,N_11364);
xnor U11653 (N_11653,N_11382,N_11316);
nand U11654 (N_11654,N_11334,N_11350);
nor U11655 (N_11655,N_11460,N_11451);
and U11656 (N_11656,N_11297,N_11302);
xor U11657 (N_11657,N_11459,N_11406);
nor U11658 (N_11658,N_11420,N_11440);
or U11659 (N_11659,N_11331,N_11462);
nor U11660 (N_11660,N_11462,N_11265);
and U11661 (N_11661,N_11284,N_11330);
and U11662 (N_11662,N_11350,N_11452);
nor U11663 (N_11663,N_11397,N_11269);
or U11664 (N_11664,N_11324,N_11464);
xor U11665 (N_11665,N_11270,N_11404);
or U11666 (N_11666,N_11263,N_11424);
and U11667 (N_11667,N_11264,N_11483);
or U11668 (N_11668,N_11308,N_11417);
xor U11669 (N_11669,N_11450,N_11269);
or U11670 (N_11670,N_11336,N_11480);
and U11671 (N_11671,N_11281,N_11428);
nor U11672 (N_11672,N_11453,N_11489);
nand U11673 (N_11673,N_11256,N_11384);
and U11674 (N_11674,N_11413,N_11317);
or U11675 (N_11675,N_11436,N_11329);
xor U11676 (N_11676,N_11312,N_11422);
xor U11677 (N_11677,N_11405,N_11479);
xor U11678 (N_11678,N_11283,N_11397);
xor U11679 (N_11679,N_11413,N_11440);
nand U11680 (N_11680,N_11390,N_11286);
and U11681 (N_11681,N_11271,N_11398);
or U11682 (N_11682,N_11296,N_11378);
nand U11683 (N_11683,N_11421,N_11389);
or U11684 (N_11684,N_11357,N_11454);
or U11685 (N_11685,N_11275,N_11482);
and U11686 (N_11686,N_11255,N_11448);
nor U11687 (N_11687,N_11298,N_11420);
or U11688 (N_11688,N_11286,N_11354);
xnor U11689 (N_11689,N_11274,N_11361);
or U11690 (N_11690,N_11477,N_11360);
nand U11691 (N_11691,N_11392,N_11277);
nor U11692 (N_11692,N_11366,N_11394);
and U11693 (N_11693,N_11361,N_11289);
xor U11694 (N_11694,N_11295,N_11458);
or U11695 (N_11695,N_11370,N_11313);
nand U11696 (N_11696,N_11283,N_11451);
or U11697 (N_11697,N_11295,N_11419);
nor U11698 (N_11698,N_11441,N_11397);
or U11699 (N_11699,N_11344,N_11383);
nand U11700 (N_11700,N_11280,N_11435);
nor U11701 (N_11701,N_11440,N_11360);
or U11702 (N_11702,N_11490,N_11280);
and U11703 (N_11703,N_11287,N_11345);
nand U11704 (N_11704,N_11476,N_11268);
nor U11705 (N_11705,N_11273,N_11370);
and U11706 (N_11706,N_11321,N_11344);
and U11707 (N_11707,N_11357,N_11334);
nand U11708 (N_11708,N_11419,N_11305);
nor U11709 (N_11709,N_11373,N_11368);
nor U11710 (N_11710,N_11291,N_11499);
or U11711 (N_11711,N_11314,N_11254);
or U11712 (N_11712,N_11472,N_11490);
and U11713 (N_11713,N_11301,N_11319);
nor U11714 (N_11714,N_11446,N_11382);
xor U11715 (N_11715,N_11304,N_11449);
nand U11716 (N_11716,N_11386,N_11341);
and U11717 (N_11717,N_11260,N_11391);
nor U11718 (N_11718,N_11407,N_11382);
xnor U11719 (N_11719,N_11258,N_11341);
or U11720 (N_11720,N_11364,N_11385);
nand U11721 (N_11721,N_11399,N_11279);
and U11722 (N_11722,N_11360,N_11482);
and U11723 (N_11723,N_11477,N_11491);
xnor U11724 (N_11724,N_11369,N_11481);
xor U11725 (N_11725,N_11261,N_11275);
nand U11726 (N_11726,N_11451,N_11479);
and U11727 (N_11727,N_11406,N_11367);
nor U11728 (N_11728,N_11477,N_11259);
nand U11729 (N_11729,N_11416,N_11450);
xnor U11730 (N_11730,N_11370,N_11436);
nor U11731 (N_11731,N_11405,N_11319);
nor U11732 (N_11732,N_11361,N_11275);
xor U11733 (N_11733,N_11276,N_11363);
nand U11734 (N_11734,N_11279,N_11446);
nand U11735 (N_11735,N_11352,N_11421);
and U11736 (N_11736,N_11372,N_11396);
xor U11737 (N_11737,N_11489,N_11487);
and U11738 (N_11738,N_11485,N_11262);
and U11739 (N_11739,N_11285,N_11493);
xor U11740 (N_11740,N_11320,N_11492);
or U11741 (N_11741,N_11477,N_11456);
or U11742 (N_11742,N_11357,N_11278);
xor U11743 (N_11743,N_11448,N_11307);
nor U11744 (N_11744,N_11263,N_11323);
and U11745 (N_11745,N_11287,N_11477);
nand U11746 (N_11746,N_11404,N_11449);
nor U11747 (N_11747,N_11445,N_11498);
xor U11748 (N_11748,N_11389,N_11351);
xor U11749 (N_11749,N_11279,N_11480);
nor U11750 (N_11750,N_11654,N_11600);
xnor U11751 (N_11751,N_11519,N_11527);
xnor U11752 (N_11752,N_11659,N_11642);
nand U11753 (N_11753,N_11554,N_11535);
nand U11754 (N_11754,N_11517,N_11672);
nand U11755 (N_11755,N_11606,N_11692);
nand U11756 (N_11756,N_11520,N_11604);
nor U11757 (N_11757,N_11631,N_11562);
nor U11758 (N_11758,N_11703,N_11731);
and U11759 (N_11759,N_11670,N_11643);
nand U11760 (N_11760,N_11619,N_11586);
and U11761 (N_11761,N_11663,N_11638);
nor U11762 (N_11762,N_11500,N_11669);
nand U11763 (N_11763,N_11577,N_11656);
and U11764 (N_11764,N_11684,N_11709);
xnor U11765 (N_11765,N_11641,N_11514);
nor U11766 (N_11766,N_11698,N_11734);
and U11767 (N_11767,N_11637,N_11532);
nor U11768 (N_11768,N_11602,N_11745);
nand U11769 (N_11769,N_11658,N_11726);
xor U11770 (N_11770,N_11609,N_11722);
nor U11771 (N_11771,N_11572,N_11627);
or U11772 (N_11772,N_11615,N_11617);
nand U11773 (N_11773,N_11714,N_11537);
and U11774 (N_11774,N_11727,N_11538);
and U11775 (N_11775,N_11723,N_11569);
or U11776 (N_11776,N_11743,N_11547);
or U11777 (N_11777,N_11650,N_11634);
nand U11778 (N_11778,N_11725,N_11705);
nor U11779 (N_11779,N_11584,N_11673);
nand U11780 (N_11780,N_11647,N_11581);
xor U11781 (N_11781,N_11608,N_11607);
or U11782 (N_11782,N_11729,N_11689);
nand U11783 (N_11783,N_11561,N_11591);
and U11784 (N_11784,N_11605,N_11702);
nor U11785 (N_11785,N_11624,N_11628);
and U11786 (N_11786,N_11644,N_11680);
or U11787 (N_11787,N_11597,N_11635);
nand U11788 (N_11788,N_11601,N_11622);
xor U11789 (N_11789,N_11664,N_11735);
xor U11790 (N_11790,N_11671,N_11616);
nor U11791 (N_11791,N_11748,N_11536);
nand U11792 (N_11792,N_11529,N_11696);
or U11793 (N_11793,N_11549,N_11582);
and U11794 (N_11794,N_11585,N_11590);
nand U11795 (N_11795,N_11704,N_11739);
nand U11796 (N_11796,N_11686,N_11575);
xor U11797 (N_11797,N_11630,N_11700);
and U11798 (N_11798,N_11510,N_11742);
or U11799 (N_11799,N_11556,N_11530);
nor U11800 (N_11800,N_11645,N_11687);
xor U11801 (N_11801,N_11675,N_11716);
xnor U11802 (N_11802,N_11545,N_11515);
xor U11803 (N_11803,N_11533,N_11712);
nand U11804 (N_11804,N_11603,N_11540);
nand U11805 (N_11805,N_11576,N_11657);
nand U11806 (N_11806,N_11667,N_11564);
nor U11807 (N_11807,N_11525,N_11541);
xnor U11808 (N_11808,N_11639,N_11553);
or U11809 (N_11809,N_11690,N_11694);
or U11810 (N_11810,N_11508,N_11701);
or U11811 (N_11811,N_11550,N_11587);
xnor U11812 (N_11812,N_11507,N_11640);
nand U11813 (N_11813,N_11524,N_11625);
and U11814 (N_11814,N_11632,N_11599);
or U11815 (N_11815,N_11559,N_11578);
nor U11816 (N_11816,N_11691,N_11614);
and U11817 (N_11817,N_11522,N_11646);
or U11818 (N_11818,N_11523,N_11555);
xnor U11819 (N_11819,N_11502,N_11678);
nor U11820 (N_11820,N_11588,N_11621);
nand U11821 (N_11821,N_11706,N_11679);
or U11822 (N_11822,N_11746,N_11717);
or U11823 (N_11823,N_11676,N_11503);
and U11824 (N_11824,N_11543,N_11668);
or U11825 (N_11825,N_11573,N_11688);
nand U11826 (N_11826,N_11720,N_11580);
xnor U11827 (N_11827,N_11548,N_11501);
xor U11828 (N_11828,N_11633,N_11516);
and U11829 (N_11829,N_11677,N_11736);
nor U11830 (N_11830,N_11740,N_11651);
or U11831 (N_11831,N_11560,N_11749);
and U11832 (N_11832,N_11737,N_11674);
nand U11833 (N_11833,N_11552,N_11693);
nor U11834 (N_11834,N_11539,N_11504);
nand U11835 (N_11835,N_11521,N_11526);
xor U11836 (N_11836,N_11741,N_11653);
nor U11837 (N_11837,N_11662,N_11595);
nor U11838 (N_11838,N_11563,N_11666);
xnor U11839 (N_11839,N_11593,N_11505);
xnor U11840 (N_11840,N_11509,N_11683);
and U11841 (N_11841,N_11682,N_11747);
nand U11842 (N_11842,N_11744,N_11506);
or U11843 (N_11843,N_11574,N_11660);
nor U11844 (N_11844,N_11629,N_11568);
and U11845 (N_11845,N_11710,N_11613);
nand U11846 (N_11846,N_11618,N_11707);
nor U11847 (N_11847,N_11649,N_11655);
nand U11848 (N_11848,N_11695,N_11699);
nand U11849 (N_11849,N_11626,N_11610);
nor U11850 (N_11850,N_11697,N_11732);
xor U11851 (N_11851,N_11512,N_11721);
and U11852 (N_11852,N_11531,N_11665);
nor U11853 (N_11853,N_11518,N_11708);
and U11854 (N_11854,N_11513,N_11579);
xnor U11855 (N_11855,N_11620,N_11636);
nor U11856 (N_11856,N_11596,N_11583);
nand U11857 (N_11857,N_11648,N_11719);
and U11858 (N_11858,N_11570,N_11589);
xnor U11859 (N_11859,N_11728,N_11681);
and U11860 (N_11860,N_11528,N_11718);
and U11861 (N_11861,N_11567,N_11652);
nor U11862 (N_11862,N_11598,N_11566);
and U11863 (N_11863,N_11557,N_11571);
nand U11864 (N_11864,N_11594,N_11713);
xnor U11865 (N_11865,N_11711,N_11730);
and U11866 (N_11866,N_11542,N_11733);
nand U11867 (N_11867,N_11661,N_11612);
or U11868 (N_11868,N_11544,N_11534);
or U11869 (N_11869,N_11558,N_11511);
xor U11870 (N_11870,N_11715,N_11685);
or U11871 (N_11871,N_11724,N_11565);
or U11872 (N_11872,N_11611,N_11592);
nor U11873 (N_11873,N_11551,N_11738);
xor U11874 (N_11874,N_11546,N_11623);
nand U11875 (N_11875,N_11638,N_11654);
nand U11876 (N_11876,N_11710,N_11639);
xnor U11877 (N_11877,N_11727,N_11503);
or U11878 (N_11878,N_11586,N_11578);
xnor U11879 (N_11879,N_11746,N_11580);
nor U11880 (N_11880,N_11573,N_11736);
or U11881 (N_11881,N_11700,N_11606);
or U11882 (N_11882,N_11691,N_11676);
and U11883 (N_11883,N_11675,N_11523);
xor U11884 (N_11884,N_11555,N_11731);
nor U11885 (N_11885,N_11537,N_11521);
nor U11886 (N_11886,N_11625,N_11617);
or U11887 (N_11887,N_11650,N_11637);
nand U11888 (N_11888,N_11579,N_11514);
nor U11889 (N_11889,N_11532,N_11501);
or U11890 (N_11890,N_11541,N_11699);
and U11891 (N_11891,N_11737,N_11527);
nor U11892 (N_11892,N_11607,N_11503);
or U11893 (N_11893,N_11523,N_11608);
or U11894 (N_11894,N_11554,N_11727);
xor U11895 (N_11895,N_11710,N_11620);
or U11896 (N_11896,N_11732,N_11736);
and U11897 (N_11897,N_11578,N_11661);
xnor U11898 (N_11898,N_11671,N_11639);
xor U11899 (N_11899,N_11528,N_11521);
or U11900 (N_11900,N_11512,N_11553);
and U11901 (N_11901,N_11512,N_11637);
nor U11902 (N_11902,N_11615,N_11725);
and U11903 (N_11903,N_11526,N_11685);
xnor U11904 (N_11904,N_11529,N_11747);
and U11905 (N_11905,N_11513,N_11556);
or U11906 (N_11906,N_11739,N_11673);
and U11907 (N_11907,N_11645,N_11569);
nor U11908 (N_11908,N_11645,N_11658);
or U11909 (N_11909,N_11571,N_11634);
or U11910 (N_11910,N_11504,N_11540);
nand U11911 (N_11911,N_11519,N_11742);
nand U11912 (N_11912,N_11737,N_11563);
and U11913 (N_11913,N_11683,N_11705);
or U11914 (N_11914,N_11534,N_11734);
or U11915 (N_11915,N_11593,N_11535);
xnor U11916 (N_11916,N_11609,N_11661);
nor U11917 (N_11917,N_11645,N_11643);
nor U11918 (N_11918,N_11603,N_11732);
or U11919 (N_11919,N_11719,N_11602);
nor U11920 (N_11920,N_11502,N_11605);
and U11921 (N_11921,N_11733,N_11684);
and U11922 (N_11922,N_11711,N_11691);
xnor U11923 (N_11923,N_11598,N_11679);
nand U11924 (N_11924,N_11625,N_11643);
nor U11925 (N_11925,N_11683,N_11531);
xnor U11926 (N_11926,N_11537,N_11652);
nor U11927 (N_11927,N_11734,N_11514);
nor U11928 (N_11928,N_11746,N_11660);
or U11929 (N_11929,N_11573,N_11567);
and U11930 (N_11930,N_11708,N_11687);
nand U11931 (N_11931,N_11720,N_11514);
or U11932 (N_11932,N_11505,N_11587);
and U11933 (N_11933,N_11546,N_11622);
or U11934 (N_11934,N_11693,N_11730);
xor U11935 (N_11935,N_11563,N_11551);
xnor U11936 (N_11936,N_11690,N_11725);
and U11937 (N_11937,N_11658,N_11516);
nor U11938 (N_11938,N_11675,N_11562);
nor U11939 (N_11939,N_11654,N_11575);
and U11940 (N_11940,N_11693,N_11635);
or U11941 (N_11941,N_11509,N_11608);
and U11942 (N_11942,N_11677,N_11649);
xnor U11943 (N_11943,N_11601,N_11602);
xor U11944 (N_11944,N_11702,N_11615);
nand U11945 (N_11945,N_11720,N_11567);
and U11946 (N_11946,N_11583,N_11566);
or U11947 (N_11947,N_11741,N_11712);
nand U11948 (N_11948,N_11534,N_11671);
xnor U11949 (N_11949,N_11501,N_11682);
nor U11950 (N_11950,N_11681,N_11541);
nand U11951 (N_11951,N_11603,N_11672);
and U11952 (N_11952,N_11745,N_11651);
and U11953 (N_11953,N_11729,N_11676);
nand U11954 (N_11954,N_11604,N_11515);
nor U11955 (N_11955,N_11540,N_11660);
nor U11956 (N_11956,N_11728,N_11657);
xor U11957 (N_11957,N_11568,N_11630);
xnor U11958 (N_11958,N_11557,N_11525);
nand U11959 (N_11959,N_11672,N_11697);
and U11960 (N_11960,N_11609,N_11713);
xor U11961 (N_11961,N_11685,N_11524);
nand U11962 (N_11962,N_11559,N_11730);
xor U11963 (N_11963,N_11571,N_11577);
nor U11964 (N_11964,N_11728,N_11742);
xor U11965 (N_11965,N_11628,N_11519);
nand U11966 (N_11966,N_11553,N_11570);
nand U11967 (N_11967,N_11540,N_11516);
xnor U11968 (N_11968,N_11736,N_11596);
nand U11969 (N_11969,N_11610,N_11736);
nand U11970 (N_11970,N_11578,N_11697);
and U11971 (N_11971,N_11610,N_11599);
xor U11972 (N_11972,N_11690,N_11630);
nor U11973 (N_11973,N_11724,N_11722);
nor U11974 (N_11974,N_11607,N_11631);
xnor U11975 (N_11975,N_11672,N_11636);
nor U11976 (N_11976,N_11615,N_11550);
xnor U11977 (N_11977,N_11716,N_11545);
xnor U11978 (N_11978,N_11653,N_11646);
xor U11979 (N_11979,N_11506,N_11504);
nor U11980 (N_11980,N_11680,N_11699);
xor U11981 (N_11981,N_11713,N_11532);
xnor U11982 (N_11982,N_11649,N_11513);
nand U11983 (N_11983,N_11540,N_11629);
and U11984 (N_11984,N_11736,N_11592);
or U11985 (N_11985,N_11649,N_11524);
xnor U11986 (N_11986,N_11716,N_11544);
and U11987 (N_11987,N_11536,N_11679);
nand U11988 (N_11988,N_11661,N_11510);
nor U11989 (N_11989,N_11658,N_11531);
nor U11990 (N_11990,N_11746,N_11620);
nor U11991 (N_11991,N_11700,N_11726);
xor U11992 (N_11992,N_11646,N_11591);
nor U11993 (N_11993,N_11531,N_11673);
nor U11994 (N_11994,N_11587,N_11723);
nor U11995 (N_11995,N_11638,N_11571);
nor U11996 (N_11996,N_11723,N_11676);
and U11997 (N_11997,N_11731,N_11572);
nand U11998 (N_11998,N_11588,N_11607);
xnor U11999 (N_11999,N_11573,N_11526);
or U12000 (N_12000,N_11903,N_11802);
nor U12001 (N_12001,N_11933,N_11870);
nand U12002 (N_12002,N_11765,N_11914);
nand U12003 (N_12003,N_11869,N_11992);
or U12004 (N_12004,N_11985,N_11763);
nand U12005 (N_12005,N_11976,N_11959);
xor U12006 (N_12006,N_11904,N_11817);
xnor U12007 (N_12007,N_11857,N_11779);
xnor U12008 (N_12008,N_11885,N_11814);
and U12009 (N_12009,N_11986,N_11878);
and U12010 (N_12010,N_11922,N_11831);
xnor U12011 (N_12011,N_11911,N_11773);
xnor U12012 (N_12012,N_11811,N_11859);
or U12013 (N_12013,N_11786,N_11908);
nand U12014 (N_12014,N_11792,N_11955);
nand U12015 (N_12015,N_11767,N_11788);
nand U12016 (N_12016,N_11810,N_11828);
xnor U12017 (N_12017,N_11842,N_11925);
or U12018 (N_12018,N_11907,N_11915);
or U12019 (N_12019,N_11896,N_11938);
and U12020 (N_12020,N_11989,N_11930);
or U12021 (N_12021,N_11919,N_11755);
nand U12022 (N_12022,N_11929,N_11939);
or U12023 (N_12023,N_11999,N_11797);
xnor U12024 (N_12024,N_11854,N_11968);
nand U12025 (N_12025,N_11761,N_11826);
xnor U12026 (N_12026,N_11863,N_11754);
and U12027 (N_12027,N_11762,N_11991);
and U12028 (N_12028,N_11946,N_11993);
or U12029 (N_12029,N_11935,N_11988);
and U12030 (N_12030,N_11884,N_11981);
xor U12031 (N_12031,N_11990,N_11972);
and U12032 (N_12032,N_11781,N_11830);
and U12033 (N_12033,N_11920,N_11950);
xnor U12034 (N_12034,N_11888,N_11756);
nand U12035 (N_12035,N_11759,N_11836);
nor U12036 (N_12036,N_11974,N_11867);
or U12037 (N_12037,N_11956,N_11924);
or U12038 (N_12038,N_11898,N_11926);
xor U12039 (N_12039,N_11790,N_11980);
nand U12040 (N_12040,N_11760,N_11832);
nor U12041 (N_12041,N_11835,N_11958);
nor U12042 (N_12042,N_11983,N_11900);
xnor U12043 (N_12043,N_11882,N_11808);
or U12044 (N_12044,N_11960,N_11780);
or U12045 (N_12045,N_11847,N_11949);
nand U12046 (N_12046,N_11962,N_11818);
nor U12047 (N_12047,N_11771,N_11772);
and U12048 (N_12048,N_11775,N_11758);
and U12049 (N_12049,N_11953,N_11864);
and U12050 (N_12050,N_11873,N_11901);
and U12051 (N_12051,N_11902,N_11899);
nor U12052 (N_12052,N_11931,N_11913);
nand U12053 (N_12053,N_11945,N_11894);
xor U12054 (N_12054,N_11851,N_11909);
nor U12055 (N_12055,N_11905,N_11838);
and U12056 (N_12056,N_11998,N_11752);
or U12057 (N_12057,N_11751,N_11969);
xnor U12058 (N_12058,N_11928,N_11805);
and U12059 (N_12059,N_11753,N_11979);
nand U12060 (N_12060,N_11778,N_11812);
xor U12061 (N_12061,N_11889,N_11875);
xnor U12062 (N_12062,N_11840,N_11943);
or U12063 (N_12063,N_11833,N_11871);
xnor U12064 (N_12064,N_11820,N_11809);
xnor U12065 (N_12065,N_11803,N_11819);
nand U12066 (N_12066,N_11793,N_11927);
nand U12067 (N_12067,N_11879,N_11963);
or U12068 (N_12068,N_11977,N_11954);
nor U12069 (N_12069,N_11937,N_11944);
and U12070 (N_12070,N_11881,N_11839);
or U12071 (N_12071,N_11934,N_11975);
nand U12072 (N_12072,N_11997,N_11941);
and U12073 (N_12073,N_11964,N_11917);
or U12074 (N_12074,N_11942,N_11855);
nand U12075 (N_12075,N_11893,N_11852);
or U12076 (N_12076,N_11895,N_11984);
nand U12077 (N_12077,N_11806,N_11799);
nor U12078 (N_12078,N_11957,N_11843);
and U12079 (N_12079,N_11789,N_11823);
nor U12080 (N_12080,N_11890,N_11872);
or U12081 (N_12081,N_11916,N_11766);
nor U12082 (N_12082,N_11800,N_11829);
nor U12083 (N_12083,N_11807,N_11825);
nor U12084 (N_12084,N_11866,N_11785);
and U12085 (N_12085,N_11824,N_11850);
xnor U12086 (N_12086,N_11845,N_11834);
or U12087 (N_12087,N_11844,N_11967);
nor U12088 (N_12088,N_11961,N_11876);
and U12089 (N_12089,N_11798,N_11995);
nor U12090 (N_12090,N_11978,N_11880);
and U12091 (N_12091,N_11770,N_11848);
xor U12092 (N_12092,N_11764,N_11952);
or U12093 (N_12093,N_11906,N_11791);
nand U12094 (N_12094,N_11783,N_11892);
or U12095 (N_12095,N_11891,N_11860);
xnor U12096 (N_12096,N_11973,N_11971);
xnor U12097 (N_12097,N_11856,N_11970);
nor U12098 (N_12098,N_11822,N_11868);
and U12099 (N_12099,N_11858,N_11951);
or U12100 (N_12100,N_11815,N_11768);
nor U12101 (N_12101,N_11936,N_11769);
nand U12102 (N_12102,N_11947,N_11923);
or U12103 (N_12103,N_11849,N_11966);
nand U12104 (N_12104,N_11784,N_11846);
nor U12105 (N_12105,N_11787,N_11965);
nand U12106 (N_12106,N_11782,N_11921);
nor U12107 (N_12107,N_11794,N_11897);
nand U12108 (N_12108,N_11795,N_11821);
or U12109 (N_12109,N_11887,N_11940);
xor U12110 (N_12110,N_11837,N_11996);
xnor U12111 (N_12111,N_11816,N_11948);
nor U12112 (N_12112,N_11874,N_11883);
and U12113 (N_12113,N_11912,N_11987);
nor U12114 (N_12114,N_11982,N_11877);
and U12115 (N_12115,N_11757,N_11865);
nor U12116 (N_12116,N_11910,N_11853);
nor U12117 (N_12117,N_11841,N_11750);
or U12118 (N_12118,N_11813,N_11777);
nor U12119 (N_12119,N_11776,N_11827);
and U12120 (N_12120,N_11932,N_11801);
nor U12121 (N_12121,N_11994,N_11774);
xor U12122 (N_12122,N_11804,N_11918);
xnor U12123 (N_12123,N_11886,N_11862);
and U12124 (N_12124,N_11861,N_11796);
nand U12125 (N_12125,N_11866,N_11857);
nor U12126 (N_12126,N_11795,N_11792);
nor U12127 (N_12127,N_11857,N_11862);
and U12128 (N_12128,N_11861,N_11858);
nand U12129 (N_12129,N_11766,N_11992);
xnor U12130 (N_12130,N_11840,N_11862);
and U12131 (N_12131,N_11849,N_11957);
nor U12132 (N_12132,N_11946,N_11917);
and U12133 (N_12133,N_11808,N_11999);
nand U12134 (N_12134,N_11802,N_11860);
or U12135 (N_12135,N_11902,N_11908);
or U12136 (N_12136,N_11750,N_11802);
and U12137 (N_12137,N_11879,N_11826);
and U12138 (N_12138,N_11771,N_11997);
and U12139 (N_12139,N_11864,N_11992);
xor U12140 (N_12140,N_11976,N_11871);
or U12141 (N_12141,N_11899,N_11924);
nor U12142 (N_12142,N_11805,N_11807);
or U12143 (N_12143,N_11815,N_11802);
and U12144 (N_12144,N_11879,N_11822);
nand U12145 (N_12145,N_11967,N_11821);
and U12146 (N_12146,N_11809,N_11834);
or U12147 (N_12147,N_11820,N_11976);
and U12148 (N_12148,N_11773,N_11792);
or U12149 (N_12149,N_11861,N_11896);
xnor U12150 (N_12150,N_11837,N_11867);
nand U12151 (N_12151,N_11804,N_11759);
nand U12152 (N_12152,N_11766,N_11871);
xnor U12153 (N_12153,N_11908,N_11825);
nor U12154 (N_12154,N_11884,N_11853);
nand U12155 (N_12155,N_11811,N_11803);
xnor U12156 (N_12156,N_11762,N_11959);
xor U12157 (N_12157,N_11769,N_11954);
nor U12158 (N_12158,N_11961,N_11754);
and U12159 (N_12159,N_11807,N_11904);
nor U12160 (N_12160,N_11860,N_11958);
nand U12161 (N_12161,N_11811,N_11923);
or U12162 (N_12162,N_11781,N_11755);
xnor U12163 (N_12163,N_11840,N_11884);
nand U12164 (N_12164,N_11791,N_11761);
nand U12165 (N_12165,N_11986,N_11937);
xnor U12166 (N_12166,N_11752,N_11931);
nor U12167 (N_12167,N_11858,N_11986);
and U12168 (N_12168,N_11804,N_11801);
and U12169 (N_12169,N_11840,N_11779);
xor U12170 (N_12170,N_11966,N_11881);
and U12171 (N_12171,N_11854,N_11921);
nand U12172 (N_12172,N_11766,N_11844);
nor U12173 (N_12173,N_11756,N_11895);
xnor U12174 (N_12174,N_11869,N_11865);
nor U12175 (N_12175,N_11789,N_11764);
nor U12176 (N_12176,N_11824,N_11810);
and U12177 (N_12177,N_11766,N_11791);
xnor U12178 (N_12178,N_11750,N_11851);
nand U12179 (N_12179,N_11892,N_11884);
xnor U12180 (N_12180,N_11913,N_11870);
xnor U12181 (N_12181,N_11883,N_11868);
nor U12182 (N_12182,N_11981,N_11823);
nor U12183 (N_12183,N_11780,N_11772);
nand U12184 (N_12184,N_11770,N_11881);
and U12185 (N_12185,N_11974,N_11901);
or U12186 (N_12186,N_11901,N_11894);
xnor U12187 (N_12187,N_11818,N_11812);
and U12188 (N_12188,N_11903,N_11896);
and U12189 (N_12189,N_11872,N_11888);
and U12190 (N_12190,N_11818,N_11947);
xor U12191 (N_12191,N_11994,N_11938);
nand U12192 (N_12192,N_11980,N_11957);
and U12193 (N_12193,N_11895,N_11976);
and U12194 (N_12194,N_11943,N_11831);
xnor U12195 (N_12195,N_11762,N_11909);
or U12196 (N_12196,N_11751,N_11974);
or U12197 (N_12197,N_11968,N_11984);
nor U12198 (N_12198,N_11971,N_11989);
nand U12199 (N_12199,N_11809,N_11893);
nor U12200 (N_12200,N_11839,N_11840);
xor U12201 (N_12201,N_11861,N_11907);
nand U12202 (N_12202,N_11878,N_11854);
xor U12203 (N_12203,N_11859,N_11974);
nor U12204 (N_12204,N_11909,N_11827);
or U12205 (N_12205,N_11755,N_11870);
nor U12206 (N_12206,N_11915,N_11991);
and U12207 (N_12207,N_11846,N_11847);
or U12208 (N_12208,N_11939,N_11759);
nand U12209 (N_12209,N_11793,N_11877);
nor U12210 (N_12210,N_11925,N_11796);
nor U12211 (N_12211,N_11828,N_11858);
nor U12212 (N_12212,N_11874,N_11759);
nand U12213 (N_12213,N_11786,N_11953);
xor U12214 (N_12214,N_11889,N_11812);
nor U12215 (N_12215,N_11921,N_11802);
or U12216 (N_12216,N_11905,N_11788);
nand U12217 (N_12217,N_11990,N_11979);
xnor U12218 (N_12218,N_11792,N_11863);
or U12219 (N_12219,N_11872,N_11944);
nor U12220 (N_12220,N_11991,N_11919);
nor U12221 (N_12221,N_11999,N_11887);
xnor U12222 (N_12222,N_11834,N_11920);
nor U12223 (N_12223,N_11972,N_11955);
xnor U12224 (N_12224,N_11933,N_11940);
nor U12225 (N_12225,N_11783,N_11961);
nand U12226 (N_12226,N_11973,N_11855);
and U12227 (N_12227,N_11915,N_11804);
xnor U12228 (N_12228,N_11770,N_11817);
and U12229 (N_12229,N_11980,N_11984);
nor U12230 (N_12230,N_11772,N_11882);
nor U12231 (N_12231,N_11769,N_11889);
xor U12232 (N_12232,N_11862,N_11971);
and U12233 (N_12233,N_11759,N_11959);
nor U12234 (N_12234,N_11825,N_11967);
or U12235 (N_12235,N_11976,N_11939);
xor U12236 (N_12236,N_11992,N_11782);
nand U12237 (N_12237,N_11777,N_11869);
xnor U12238 (N_12238,N_11912,N_11945);
and U12239 (N_12239,N_11782,N_11761);
xor U12240 (N_12240,N_11807,N_11846);
xnor U12241 (N_12241,N_11883,N_11788);
and U12242 (N_12242,N_11804,N_11975);
nor U12243 (N_12243,N_11874,N_11839);
or U12244 (N_12244,N_11962,N_11779);
or U12245 (N_12245,N_11929,N_11790);
nor U12246 (N_12246,N_11954,N_11839);
xor U12247 (N_12247,N_11965,N_11799);
and U12248 (N_12248,N_11983,N_11877);
or U12249 (N_12249,N_11777,N_11882);
nand U12250 (N_12250,N_12144,N_12199);
or U12251 (N_12251,N_12083,N_12043);
and U12252 (N_12252,N_12078,N_12006);
nor U12253 (N_12253,N_12185,N_12056);
or U12254 (N_12254,N_12242,N_12062);
nand U12255 (N_12255,N_12073,N_12207);
or U12256 (N_12256,N_12081,N_12036);
and U12257 (N_12257,N_12241,N_12070);
nor U12258 (N_12258,N_12243,N_12063);
nand U12259 (N_12259,N_12152,N_12061);
nand U12260 (N_12260,N_12065,N_12216);
nand U12261 (N_12261,N_12112,N_12196);
xor U12262 (N_12262,N_12190,N_12197);
nand U12263 (N_12263,N_12131,N_12172);
xnor U12264 (N_12264,N_12118,N_12060);
xnor U12265 (N_12265,N_12004,N_12101);
nor U12266 (N_12266,N_12040,N_12170);
and U12267 (N_12267,N_12123,N_12219);
and U12268 (N_12268,N_12029,N_12168);
nor U12269 (N_12269,N_12008,N_12195);
xnor U12270 (N_12270,N_12104,N_12249);
nor U12271 (N_12271,N_12149,N_12092);
and U12272 (N_12272,N_12102,N_12133);
nor U12273 (N_12273,N_12163,N_12090);
or U12274 (N_12274,N_12137,N_12127);
xor U12275 (N_12275,N_12237,N_12119);
or U12276 (N_12276,N_12224,N_12244);
or U12277 (N_12277,N_12132,N_12212);
nor U12278 (N_12278,N_12179,N_12178);
and U12279 (N_12279,N_12174,N_12231);
or U12280 (N_12280,N_12009,N_12186);
or U12281 (N_12281,N_12171,N_12027);
nand U12282 (N_12282,N_12156,N_12136);
nor U12283 (N_12283,N_12176,N_12183);
xnor U12284 (N_12284,N_12228,N_12113);
nor U12285 (N_12285,N_12147,N_12015);
nand U12286 (N_12286,N_12210,N_12184);
xnor U12287 (N_12287,N_12018,N_12201);
nor U12288 (N_12288,N_12191,N_12005);
nor U12289 (N_12289,N_12048,N_12225);
and U12290 (N_12290,N_12103,N_12020);
nor U12291 (N_12291,N_12054,N_12044);
xnor U12292 (N_12292,N_12223,N_12106);
and U12293 (N_12293,N_12097,N_12026);
xor U12294 (N_12294,N_12138,N_12204);
xor U12295 (N_12295,N_12135,N_12175);
xor U12296 (N_12296,N_12116,N_12202);
xor U12297 (N_12297,N_12145,N_12213);
nor U12298 (N_12298,N_12235,N_12206);
xnor U12299 (N_12299,N_12182,N_12037);
or U12300 (N_12300,N_12014,N_12052);
xnor U12301 (N_12301,N_12130,N_12248);
nor U12302 (N_12302,N_12039,N_12177);
and U12303 (N_12303,N_12033,N_12158);
or U12304 (N_12304,N_12028,N_12167);
xnor U12305 (N_12305,N_12042,N_12074);
xnor U12306 (N_12306,N_12245,N_12120);
nor U12307 (N_12307,N_12222,N_12205);
or U12308 (N_12308,N_12087,N_12181);
nor U12309 (N_12309,N_12068,N_12208);
nor U12310 (N_12310,N_12002,N_12093);
nand U12311 (N_12311,N_12066,N_12236);
xnor U12312 (N_12312,N_12079,N_12082);
xnor U12313 (N_12313,N_12143,N_12076);
xnor U12314 (N_12314,N_12173,N_12069);
or U12315 (N_12315,N_12151,N_12150);
or U12316 (N_12316,N_12154,N_12214);
xor U12317 (N_12317,N_12215,N_12155);
nand U12318 (N_12318,N_12098,N_12217);
and U12319 (N_12319,N_12211,N_12059);
or U12320 (N_12320,N_12064,N_12053);
xnor U12321 (N_12321,N_12021,N_12058);
xor U12322 (N_12322,N_12166,N_12165);
nand U12323 (N_12323,N_12114,N_12134);
or U12324 (N_12324,N_12125,N_12221);
nor U12325 (N_12325,N_12072,N_12232);
or U12326 (N_12326,N_12031,N_12148);
xor U12327 (N_12327,N_12162,N_12038);
or U12328 (N_12328,N_12218,N_12055);
xnor U12329 (N_12329,N_12105,N_12227);
nand U12330 (N_12330,N_12025,N_12067);
nand U12331 (N_12331,N_12047,N_12091);
and U12332 (N_12332,N_12088,N_12084);
nor U12333 (N_12333,N_12140,N_12046);
xnor U12334 (N_12334,N_12071,N_12095);
nand U12335 (N_12335,N_12146,N_12209);
nor U12336 (N_12336,N_12159,N_12203);
nor U12337 (N_12337,N_12180,N_12234);
nand U12338 (N_12338,N_12000,N_12080);
nand U12339 (N_12339,N_12240,N_12188);
or U12340 (N_12340,N_12094,N_12077);
nand U12341 (N_12341,N_12086,N_12246);
nand U12342 (N_12342,N_12239,N_12193);
xnor U12343 (N_12343,N_12139,N_12189);
xor U12344 (N_12344,N_12200,N_12051);
nand U12345 (N_12345,N_12194,N_12024);
and U12346 (N_12346,N_12108,N_12022);
nor U12347 (N_12347,N_12198,N_12247);
nor U12348 (N_12348,N_12041,N_12085);
or U12349 (N_12349,N_12057,N_12107);
nor U12350 (N_12350,N_12192,N_12007);
nand U12351 (N_12351,N_12141,N_12030);
and U12352 (N_12352,N_12220,N_12035);
nand U12353 (N_12353,N_12032,N_12003);
or U12354 (N_12354,N_12121,N_12126);
nor U12355 (N_12355,N_12226,N_12023);
and U12356 (N_12356,N_12160,N_12096);
nand U12357 (N_12357,N_12010,N_12034);
nand U12358 (N_12358,N_12045,N_12128);
nand U12359 (N_12359,N_12153,N_12016);
xnor U12360 (N_12360,N_12075,N_12129);
and U12361 (N_12361,N_12230,N_12161);
xnor U12362 (N_12362,N_12169,N_12111);
and U12363 (N_12363,N_12115,N_12017);
xnor U12364 (N_12364,N_12012,N_12001);
nor U12365 (N_12365,N_12124,N_12089);
nor U12366 (N_12366,N_12122,N_12050);
or U12367 (N_12367,N_12142,N_12187);
or U12368 (N_12368,N_12110,N_12164);
xnor U12369 (N_12369,N_12229,N_12109);
or U12370 (N_12370,N_12013,N_12100);
nand U12371 (N_12371,N_12049,N_12238);
or U12372 (N_12372,N_12099,N_12011);
xor U12373 (N_12373,N_12019,N_12157);
and U12374 (N_12374,N_12117,N_12233);
xor U12375 (N_12375,N_12135,N_12055);
xor U12376 (N_12376,N_12248,N_12193);
nand U12377 (N_12377,N_12042,N_12148);
and U12378 (N_12378,N_12123,N_12201);
and U12379 (N_12379,N_12204,N_12115);
nand U12380 (N_12380,N_12079,N_12211);
or U12381 (N_12381,N_12064,N_12219);
xor U12382 (N_12382,N_12210,N_12147);
or U12383 (N_12383,N_12115,N_12207);
and U12384 (N_12384,N_12081,N_12030);
and U12385 (N_12385,N_12224,N_12213);
nand U12386 (N_12386,N_12151,N_12231);
and U12387 (N_12387,N_12154,N_12069);
nor U12388 (N_12388,N_12227,N_12163);
or U12389 (N_12389,N_12039,N_12069);
nand U12390 (N_12390,N_12101,N_12105);
xor U12391 (N_12391,N_12083,N_12028);
xnor U12392 (N_12392,N_12185,N_12072);
nand U12393 (N_12393,N_12101,N_12050);
nand U12394 (N_12394,N_12203,N_12057);
or U12395 (N_12395,N_12056,N_12180);
nor U12396 (N_12396,N_12102,N_12032);
or U12397 (N_12397,N_12086,N_12093);
and U12398 (N_12398,N_12047,N_12079);
xor U12399 (N_12399,N_12088,N_12160);
and U12400 (N_12400,N_12205,N_12040);
nand U12401 (N_12401,N_12171,N_12073);
nor U12402 (N_12402,N_12172,N_12074);
nand U12403 (N_12403,N_12026,N_12178);
and U12404 (N_12404,N_12189,N_12157);
xor U12405 (N_12405,N_12019,N_12128);
xnor U12406 (N_12406,N_12076,N_12003);
and U12407 (N_12407,N_12087,N_12033);
xor U12408 (N_12408,N_12220,N_12090);
nor U12409 (N_12409,N_12126,N_12144);
and U12410 (N_12410,N_12065,N_12220);
nor U12411 (N_12411,N_12192,N_12178);
nor U12412 (N_12412,N_12001,N_12055);
nor U12413 (N_12413,N_12228,N_12028);
or U12414 (N_12414,N_12010,N_12081);
nand U12415 (N_12415,N_12011,N_12016);
or U12416 (N_12416,N_12125,N_12106);
or U12417 (N_12417,N_12074,N_12043);
or U12418 (N_12418,N_12248,N_12135);
or U12419 (N_12419,N_12230,N_12174);
nand U12420 (N_12420,N_12062,N_12146);
xnor U12421 (N_12421,N_12133,N_12210);
nor U12422 (N_12422,N_12071,N_12198);
or U12423 (N_12423,N_12174,N_12239);
or U12424 (N_12424,N_12174,N_12077);
and U12425 (N_12425,N_12047,N_12055);
nor U12426 (N_12426,N_12240,N_12185);
nor U12427 (N_12427,N_12204,N_12105);
or U12428 (N_12428,N_12133,N_12040);
nor U12429 (N_12429,N_12106,N_12029);
nand U12430 (N_12430,N_12240,N_12051);
or U12431 (N_12431,N_12194,N_12203);
or U12432 (N_12432,N_12139,N_12137);
nor U12433 (N_12433,N_12020,N_12136);
and U12434 (N_12434,N_12106,N_12151);
or U12435 (N_12435,N_12231,N_12137);
or U12436 (N_12436,N_12116,N_12204);
nor U12437 (N_12437,N_12114,N_12071);
nor U12438 (N_12438,N_12211,N_12109);
or U12439 (N_12439,N_12209,N_12192);
and U12440 (N_12440,N_12063,N_12020);
nor U12441 (N_12441,N_12064,N_12038);
nor U12442 (N_12442,N_12121,N_12027);
and U12443 (N_12443,N_12017,N_12026);
xor U12444 (N_12444,N_12017,N_12083);
or U12445 (N_12445,N_12235,N_12202);
xor U12446 (N_12446,N_12238,N_12110);
or U12447 (N_12447,N_12216,N_12096);
nand U12448 (N_12448,N_12003,N_12062);
nand U12449 (N_12449,N_12175,N_12088);
or U12450 (N_12450,N_12196,N_12129);
or U12451 (N_12451,N_12030,N_12108);
xor U12452 (N_12452,N_12249,N_12158);
or U12453 (N_12453,N_12150,N_12018);
or U12454 (N_12454,N_12206,N_12168);
nor U12455 (N_12455,N_12230,N_12222);
nor U12456 (N_12456,N_12227,N_12088);
xnor U12457 (N_12457,N_12113,N_12232);
or U12458 (N_12458,N_12061,N_12238);
or U12459 (N_12459,N_12065,N_12201);
or U12460 (N_12460,N_12099,N_12218);
xnor U12461 (N_12461,N_12147,N_12017);
or U12462 (N_12462,N_12070,N_12189);
nor U12463 (N_12463,N_12010,N_12204);
or U12464 (N_12464,N_12115,N_12143);
and U12465 (N_12465,N_12070,N_12201);
xnor U12466 (N_12466,N_12016,N_12041);
xnor U12467 (N_12467,N_12222,N_12135);
xnor U12468 (N_12468,N_12225,N_12183);
and U12469 (N_12469,N_12249,N_12191);
xor U12470 (N_12470,N_12117,N_12039);
and U12471 (N_12471,N_12143,N_12110);
nand U12472 (N_12472,N_12136,N_12043);
xnor U12473 (N_12473,N_12101,N_12031);
or U12474 (N_12474,N_12097,N_12155);
or U12475 (N_12475,N_12069,N_12156);
nor U12476 (N_12476,N_12172,N_12183);
xor U12477 (N_12477,N_12149,N_12115);
xor U12478 (N_12478,N_12106,N_12166);
and U12479 (N_12479,N_12186,N_12047);
nor U12480 (N_12480,N_12177,N_12214);
and U12481 (N_12481,N_12042,N_12044);
and U12482 (N_12482,N_12131,N_12047);
xor U12483 (N_12483,N_12107,N_12014);
nand U12484 (N_12484,N_12064,N_12067);
nor U12485 (N_12485,N_12162,N_12204);
and U12486 (N_12486,N_12004,N_12217);
nand U12487 (N_12487,N_12141,N_12074);
or U12488 (N_12488,N_12207,N_12116);
xor U12489 (N_12489,N_12249,N_12132);
or U12490 (N_12490,N_12212,N_12170);
and U12491 (N_12491,N_12100,N_12068);
nor U12492 (N_12492,N_12020,N_12092);
or U12493 (N_12493,N_12037,N_12066);
xnor U12494 (N_12494,N_12114,N_12075);
nor U12495 (N_12495,N_12003,N_12069);
or U12496 (N_12496,N_12119,N_12004);
or U12497 (N_12497,N_12070,N_12039);
nor U12498 (N_12498,N_12003,N_12104);
or U12499 (N_12499,N_12083,N_12217);
nor U12500 (N_12500,N_12485,N_12347);
nand U12501 (N_12501,N_12294,N_12325);
or U12502 (N_12502,N_12457,N_12356);
nand U12503 (N_12503,N_12254,N_12368);
nor U12504 (N_12504,N_12260,N_12316);
and U12505 (N_12505,N_12322,N_12461);
or U12506 (N_12506,N_12374,N_12293);
nand U12507 (N_12507,N_12475,N_12450);
and U12508 (N_12508,N_12443,N_12494);
nand U12509 (N_12509,N_12497,N_12357);
nand U12510 (N_12510,N_12439,N_12292);
or U12511 (N_12511,N_12253,N_12392);
or U12512 (N_12512,N_12272,N_12299);
xor U12513 (N_12513,N_12403,N_12287);
nand U12514 (N_12514,N_12496,N_12452);
nor U12515 (N_12515,N_12381,N_12456);
and U12516 (N_12516,N_12335,N_12300);
xor U12517 (N_12517,N_12416,N_12409);
and U12518 (N_12518,N_12426,N_12404);
nand U12519 (N_12519,N_12408,N_12464);
nor U12520 (N_12520,N_12290,N_12307);
nand U12521 (N_12521,N_12481,N_12402);
nand U12522 (N_12522,N_12378,N_12281);
nor U12523 (N_12523,N_12435,N_12448);
or U12524 (N_12524,N_12442,N_12274);
nand U12525 (N_12525,N_12284,N_12495);
xor U12526 (N_12526,N_12359,N_12326);
or U12527 (N_12527,N_12479,N_12454);
xor U12528 (N_12528,N_12405,N_12472);
xnor U12529 (N_12529,N_12476,N_12343);
xor U12530 (N_12530,N_12327,N_12372);
and U12531 (N_12531,N_12469,N_12484);
nor U12532 (N_12532,N_12367,N_12470);
xnor U12533 (N_12533,N_12342,N_12463);
xnor U12534 (N_12534,N_12283,N_12425);
or U12535 (N_12535,N_12353,N_12473);
xor U12536 (N_12536,N_12362,N_12411);
or U12537 (N_12537,N_12398,N_12433);
nand U12538 (N_12538,N_12382,N_12477);
xor U12539 (N_12539,N_12380,N_12258);
or U12540 (N_12540,N_12266,N_12467);
xor U12541 (N_12541,N_12318,N_12345);
nor U12542 (N_12542,N_12465,N_12384);
nand U12543 (N_12543,N_12311,N_12455);
nand U12544 (N_12544,N_12360,N_12346);
nand U12545 (N_12545,N_12371,N_12332);
nor U12546 (N_12546,N_12369,N_12262);
and U12547 (N_12547,N_12490,N_12419);
xor U12548 (N_12548,N_12298,N_12333);
or U12549 (N_12549,N_12491,N_12478);
nand U12550 (N_12550,N_12257,N_12423);
xnor U12551 (N_12551,N_12460,N_12498);
and U12552 (N_12552,N_12317,N_12387);
xor U12553 (N_12553,N_12377,N_12256);
xor U12554 (N_12554,N_12483,N_12330);
nor U12555 (N_12555,N_12441,N_12418);
or U12556 (N_12556,N_12389,N_12487);
and U12557 (N_12557,N_12399,N_12269);
or U12558 (N_12558,N_12458,N_12414);
nand U12559 (N_12559,N_12492,N_12273);
xnor U12560 (N_12560,N_12310,N_12429);
xnor U12561 (N_12561,N_12361,N_12267);
or U12562 (N_12562,N_12275,N_12352);
xnor U12563 (N_12563,N_12393,N_12390);
nor U12564 (N_12564,N_12324,N_12431);
nor U12565 (N_12565,N_12339,N_12412);
nor U12566 (N_12566,N_12340,N_12305);
or U12567 (N_12567,N_12451,N_12410);
or U12568 (N_12568,N_12270,N_12264);
nand U12569 (N_12569,N_12391,N_12313);
nand U12570 (N_12570,N_12420,N_12474);
nor U12571 (N_12571,N_12251,N_12302);
or U12572 (N_12572,N_12468,N_12295);
or U12573 (N_12573,N_12444,N_12323);
nor U12574 (N_12574,N_12303,N_12289);
nor U12575 (N_12575,N_12364,N_12499);
xnor U12576 (N_12576,N_12376,N_12471);
nand U12577 (N_12577,N_12480,N_12355);
xor U12578 (N_12578,N_12268,N_12301);
xnor U12579 (N_12579,N_12459,N_12482);
or U12580 (N_12580,N_12438,N_12337);
or U12581 (N_12581,N_12328,N_12341);
nand U12582 (N_12582,N_12415,N_12383);
and U12583 (N_12583,N_12351,N_12331);
nand U12584 (N_12584,N_12489,N_12432);
nand U12585 (N_12585,N_12312,N_12440);
nand U12586 (N_12586,N_12385,N_12250);
xor U12587 (N_12587,N_12279,N_12379);
or U12588 (N_12588,N_12285,N_12308);
nor U12589 (N_12589,N_12348,N_12291);
nand U12590 (N_12590,N_12363,N_12280);
xnor U12591 (N_12591,N_12286,N_12255);
or U12592 (N_12592,N_12338,N_12413);
or U12593 (N_12593,N_12265,N_12306);
xnor U12594 (N_12594,N_12263,N_12373);
or U12595 (N_12595,N_12394,N_12336);
or U12596 (N_12596,N_12406,N_12397);
xor U12597 (N_12597,N_12309,N_12296);
nand U12598 (N_12598,N_12344,N_12428);
nor U12599 (N_12599,N_12350,N_12401);
xor U12600 (N_12600,N_12261,N_12288);
nand U12601 (N_12601,N_12488,N_12314);
or U12602 (N_12602,N_12445,N_12320);
nor U12603 (N_12603,N_12329,N_12462);
and U12604 (N_12604,N_12304,N_12271);
nor U12605 (N_12605,N_12493,N_12421);
nand U12606 (N_12606,N_12395,N_12277);
or U12607 (N_12607,N_12297,N_12334);
nand U12608 (N_12608,N_12375,N_12386);
nor U12609 (N_12609,N_12422,N_12278);
nor U12610 (N_12610,N_12349,N_12437);
nand U12611 (N_12611,N_12424,N_12396);
or U12612 (N_12612,N_12407,N_12400);
and U12613 (N_12613,N_12427,N_12276);
nor U12614 (N_12614,N_12319,N_12430);
nand U12615 (N_12615,N_12366,N_12449);
xnor U12616 (N_12616,N_12282,N_12388);
or U12617 (N_12617,N_12436,N_12417);
and U12618 (N_12618,N_12486,N_12315);
xnor U12619 (N_12619,N_12453,N_12446);
and U12620 (N_12620,N_12447,N_12434);
or U12621 (N_12621,N_12358,N_12252);
nor U12622 (N_12622,N_12259,N_12466);
or U12623 (N_12623,N_12321,N_12365);
nand U12624 (N_12624,N_12354,N_12370);
or U12625 (N_12625,N_12309,N_12369);
nand U12626 (N_12626,N_12291,N_12459);
and U12627 (N_12627,N_12350,N_12412);
nor U12628 (N_12628,N_12329,N_12472);
or U12629 (N_12629,N_12321,N_12395);
nand U12630 (N_12630,N_12452,N_12337);
xor U12631 (N_12631,N_12435,N_12270);
nand U12632 (N_12632,N_12282,N_12324);
xnor U12633 (N_12633,N_12488,N_12273);
or U12634 (N_12634,N_12456,N_12399);
nand U12635 (N_12635,N_12378,N_12413);
nor U12636 (N_12636,N_12496,N_12360);
xor U12637 (N_12637,N_12415,N_12295);
nand U12638 (N_12638,N_12452,N_12424);
xnor U12639 (N_12639,N_12483,N_12474);
nor U12640 (N_12640,N_12259,N_12338);
xor U12641 (N_12641,N_12434,N_12264);
nand U12642 (N_12642,N_12482,N_12292);
nor U12643 (N_12643,N_12419,N_12401);
nand U12644 (N_12644,N_12424,N_12288);
and U12645 (N_12645,N_12344,N_12486);
or U12646 (N_12646,N_12402,N_12412);
xnor U12647 (N_12647,N_12448,N_12283);
nor U12648 (N_12648,N_12412,N_12471);
nand U12649 (N_12649,N_12343,N_12354);
nand U12650 (N_12650,N_12335,N_12400);
xnor U12651 (N_12651,N_12375,N_12329);
and U12652 (N_12652,N_12262,N_12440);
xnor U12653 (N_12653,N_12295,N_12256);
nor U12654 (N_12654,N_12487,N_12290);
xnor U12655 (N_12655,N_12290,N_12490);
or U12656 (N_12656,N_12486,N_12499);
nand U12657 (N_12657,N_12499,N_12283);
or U12658 (N_12658,N_12455,N_12481);
nor U12659 (N_12659,N_12449,N_12255);
nand U12660 (N_12660,N_12274,N_12435);
nor U12661 (N_12661,N_12265,N_12380);
and U12662 (N_12662,N_12293,N_12452);
nor U12663 (N_12663,N_12318,N_12499);
xor U12664 (N_12664,N_12289,N_12315);
nand U12665 (N_12665,N_12367,N_12307);
or U12666 (N_12666,N_12301,N_12443);
nand U12667 (N_12667,N_12472,N_12481);
xor U12668 (N_12668,N_12281,N_12252);
and U12669 (N_12669,N_12380,N_12436);
nand U12670 (N_12670,N_12486,N_12331);
nor U12671 (N_12671,N_12314,N_12354);
nand U12672 (N_12672,N_12464,N_12300);
or U12673 (N_12673,N_12408,N_12436);
nand U12674 (N_12674,N_12417,N_12492);
nand U12675 (N_12675,N_12457,N_12271);
and U12676 (N_12676,N_12256,N_12267);
nand U12677 (N_12677,N_12316,N_12293);
nand U12678 (N_12678,N_12365,N_12323);
or U12679 (N_12679,N_12374,N_12272);
and U12680 (N_12680,N_12350,N_12455);
nand U12681 (N_12681,N_12428,N_12254);
or U12682 (N_12682,N_12261,N_12495);
and U12683 (N_12683,N_12453,N_12341);
and U12684 (N_12684,N_12387,N_12459);
xnor U12685 (N_12685,N_12483,N_12314);
xor U12686 (N_12686,N_12358,N_12457);
and U12687 (N_12687,N_12385,N_12338);
or U12688 (N_12688,N_12454,N_12295);
and U12689 (N_12689,N_12310,N_12477);
xnor U12690 (N_12690,N_12328,N_12269);
nand U12691 (N_12691,N_12426,N_12387);
and U12692 (N_12692,N_12335,N_12325);
nand U12693 (N_12693,N_12475,N_12260);
or U12694 (N_12694,N_12262,N_12323);
nor U12695 (N_12695,N_12492,N_12482);
and U12696 (N_12696,N_12267,N_12366);
and U12697 (N_12697,N_12284,N_12375);
nor U12698 (N_12698,N_12322,N_12468);
nand U12699 (N_12699,N_12345,N_12266);
nor U12700 (N_12700,N_12375,N_12463);
nand U12701 (N_12701,N_12269,N_12414);
xor U12702 (N_12702,N_12281,N_12276);
nor U12703 (N_12703,N_12448,N_12418);
nor U12704 (N_12704,N_12433,N_12461);
xor U12705 (N_12705,N_12264,N_12421);
xnor U12706 (N_12706,N_12407,N_12298);
and U12707 (N_12707,N_12356,N_12349);
and U12708 (N_12708,N_12431,N_12348);
nand U12709 (N_12709,N_12387,N_12381);
or U12710 (N_12710,N_12444,N_12396);
xnor U12711 (N_12711,N_12340,N_12350);
xnor U12712 (N_12712,N_12343,N_12253);
and U12713 (N_12713,N_12272,N_12435);
and U12714 (N_12714,N_12281,N_12345);
xor U12715 (N_12715,N_12491,N_12353);
xnor U12716 (N_12716,N_12418,N_12273);
nor U12717 (N_12717,N_12352,N_12354);
or U12718 (N_12718,N_12408,N_12456);
and U12719 (N_12719,N_12284,N_12291);
nand U12720 (N_12720,N_12371,N_12382);
xor U12721 (N_12721,N_12495,N_12474);
xor U12722 (N_12722,N_12448,N_12356);
and U12723 (N_12723,N_12298,N_12465);
nand U12724 (N_12724,N_12498,N_12294);
nand U12725 (N_12725,N_12467,N_12251);
nor U12726 (N_12726,N_12360,N_12431);
or U12727 (N_12727,N_12383,N_12452);
or U12728 (N_12728,N_12424,N_12463);
xnor U12729 (N_12729,N_12490,N_12384);
xnor U12730 (N_12730,N_12439,N_12416);
and U12731 (N_12731,N_12334,N_12482);
nor U12732 (N_12732,N_12472,N_12324);
nor U12733 (N_12733,N_12341,N_12309);
or U12734 (N_12734,N_12450,N_12383);
xnor U12735 (N_12735,N_12473,N_12335);
nor U12736 (N_12736,N_12355,N_12350);
nor U12737 (N_12737,N_12314,N_12300);
or U12738 (N_12738,N_12333,N_12254);
or U12739 (N_12739,N_12298,N_12429);
or U12740 (N_12740,N_12425,N_12442);
nor U12741 (N_12741,N_12380,N_12454);
nand U12742 (N_12742,N_12274,N_12403);
xor U12743 (N_12743,N_12400,N_12369);
or U12744 (N_12744,N_12360,N_12418);
xor U12745 (N_12745,N_12432,N_12470);
xnor U12746 (N_12746,N_12389,N_12476);
or U12747 (N_12747,N_12436,N_12255);
xor U12748 (N_12748,N_12391,N_12261);
nor U12749 (N_12749,N_12336,N_12471);
xor U12750 (N_12750,N_12646,N_12695);
xor U12751 (N_12751,N_12725,N_12692);
nand U12752 (N_12752,N_12539,N_12582);
nor U12753 (N_12753,N_12713,N_12500);
and U12754 (N_12754,N_12737,N_12586);
nand U12755 (N_12755,N_12532,N_12517);
nand U12756 (N_12756,N_12739,N_12508);
or U12757 (N_12757,N_12664,N_12667);
or U12758 (N_12758,N_12526,N_12738);
nand U12759 (N_12759,N_12729,N_12572);
or U12760 (N_12760,N_12510,N_12600);
nor U12761 (N_12761,N_12696,N_12732);
and U12762 (N_12762,N_12556,N_12565);
nand U12763 (N_12763,N_12523,N_12703);
nand U12764 (N_12764,N_12649,N_12598);
xor U12765 (N_12765,N_12727,N_12548);
xnor U12766 (N_12766,N_12679,N_12672);
nor U12767 (N_12767,N_12528,N_12519);
nand U12768 (N_12768,N_12531,N_12615);
or U12769 (N_12769,N_12693,N_12647);
nor U12770 (N_12770,N_12574,N_12515);
nand U12771 (N_12771,N_12663,N_12557);
and U12772 (N_12772,N_12516,N_12666);
and U12773 (N_12773,N_12563,N_12654);
or U12774 (N_12774,N_12733,N_12699);
nor U12775 (N_12775,N_12509,N_12669);
and U12776 (N_12776,N_12685,N_12564);
nor U12777 (N_12777,N_12512,N_12620);
xor U12778 (N_12778,N_12655,N_12577);
and U12779 (N_12779,N_12579,N_12723);
xor U12780 (N_12780,N_12540,N_12559);
nand U12781 (N_12781,N_12661,N_12637);
nand U12782 (N_12782,N_12588,N_12589);
nor U12783 (N_12783,N_12636,N_12627);
nand U12784 (N_12784,N_12622,N_12629);
and U12785 (N_12785,N_12625,N_12507);
or U12786 (N_12786,N_12529,N_12658);
or U12787 (N_12787,N_12665,N_12599);
and U12788 (N_12788,N_12734,N_12578);
or U12789 (N_12789,N_12660,N_12639);
or U12790 (N_12790,N_12594,N_12644);
and U12791 (N_12791,N_12705,N_12743);
nor U12792 (N_12792,N_12561,N_12682);
nand U12793 (N_12793,N_12538,N_12670);
or U12794 (N_12794,N_12533,N_12706);
or U12795 (N_12795,N_12688,N_12656);
xnor U12796 (N_12796,N_12716,N_12592);
and U12797 (N_12797,N_12676,N_12648);
or U12798 (N_12798,N_12616,N_12736);
or U12799 (N_12799,N_12580,N_12546);
nor U12800 (N_12800,N_12535,N_12575);
nor U12801 (N_12801,N_12748,N_12645);
and U12802 (N_12802,N_12534,N_12542);
and U12803 (N_12803,N_12651,N_12614);
or U12804 (N_12804,N_12721,N_12747);
nor U12805 (N_12805,N_12518,N_12501);
xnor U12806 (N_12806,N_12724,N_12605);
nor U12807 (N_12807,N_12746,N_12536);
xnor U12808 (N_12808,N_12584,N_12573);
or U12809 (N_12809,N_12544,N_12643);
or U12810 (N_12810,N_12617,N_12623);
nor U12811 (N_12811,N_12697,N_12630);
or U12812 (N_12812,N_12590,N_12680);
nor U12813 (N_12813,N_12612,N_12511);
nor U12814 (N_12814,N_12571,N_12671);
nor U12815 (N_12815,N_12562,N_12631);
xor U12816 (N_12816,N_12681,N_12502);
and U12817 (N_12817,N_12566,N_12677);
and U12818 (N_12818,N_12601,N_12744);
and U12819 (N_12819,N_12603,N_12583);
nor U12820 (N_12820,N_12555,N_12674);
nand U12821 (N_12821,N_12728,N_12570);
nand U12822 (N_12822,N_12690,N_12653);
nand U12823 (N_12823,N_12715,N_12726);
and U12824 (N_12824,N_12722,N_12608);
nand U12825 (N_12825,N_12708,N_12530);
xor U12826 (N_12826,N_12642,N_12668);
or U12827 (N_12827,N_12541,N_12550);
and U12828 (N_12828,N_12635,N_12652);
xor U12829 (N_12829,N_12545,N_12606);
and U12830 (N_12830,N_12662,N_12711);
nor U12831 (N_12831,N_12731,N_12552);
nand U12832 (N_12832,N_12522,N_12569);
nand U12833 (N_12833,N_12621,N_12611);
nor U12834 (N_12834,N_12741,N_12596);
or U12835 (N_12835,N_12700,N_12687);
or U12836 (N_12836,N_12597,N_12673);
nor U12837 (N_12837,N_12650,N_12525);
or U12838 (N_12838,N_12585,N_12587);
xnor U12839 (N_12839,N_12506,N_12593);
and U12840 (N_12840,N_12628,N_12520);
nand U12841 (N_12841,N_12707,N_12657);
nand U12842 (N_12842,N_12524,N_12521);
nand U12843 (N_12843,N_12735,N_12568);
and U12844 (N_12844,N_12609,N_12730);
nand U12845 (N_12845,N_12691,N_12619);
nor U12846 (N_12846,N_12720,N_12717);
or U12847 (N_12847,N_12638,N_12659);
and U12848 (N_12848,N_12610,N_12675);
xnor U12849 (N_12849,N_12634,N_12745);
or U12850 (N_12850,N_12701,N_12613);
and U12851 (N_12851,N_12549,N_12547);
nor U12852 (N_12852,N_12505,N_12543);
or U12853 (N_12853,N_12640,N_12633);
or U12854 (N_12854,N_12553,N_12576);
and U12855 (N_12855,N_12602,N_12527);
xor U12856 (N_12856,N_12513,N_12537);
and U12857 (N_12857,N_12740,N_12714);
and U12858 (N_12858,N_12719,N_12624);
xnor U12859 (N_12859,N_12704,N_12581);
or U12860 (N_12860,N_12710,N_12712);
and U12861 (N_12861,N_12641,N_12504);
nor U12862 (N_12862,N_12604,N_12718);
or U12863 (N_12863,N_12686,N_12683);
and U12864 (N_12864,N_12684,N_12694);
xnor U12865 (N_12865,N_12591,N_12607);
xnor U12866 (N_12866,N_12560,N_12567);
nor U12867 (N_12867,N_12618,N_12702);
and U12868 (N_12868,N_12595,N_12742);
or U12869 (N_12869,N_12551,N_12554);
and U12870 (N_12870,N_12709,N_12689);
nand U12871 (N_12871,N_12514,N_12626);
and U12872 (N_12872,N_12558,N_12698);
nor U12873 (N_12873,N_12632,N_12503);
and U12874 (N_12874,N_12749,N_12678);
and U12875 (N_12875,N_12707,N_12719);
xor U12876 (N_12876,N_12570,N_12582);
xnor U12877 (N_12877,N_12600,N_12699);
xor U12878 (N_12878,N_12719,N_12593);
nand U12879 (N_12879,N_12721,N_12548);
nor U12880 (N_12880,N_12655,N_12611);
and U12881 (N_12881,N_12625,N_12636);
or U12882 (N_12882,N_12503,N_12561);
xor U12883 (N_12883,N_12596,N_12667);
xor U12884 (N_12884,N_12637,N_12683);
or U12885 (N_12885,N_12563,N_12736);
xnor U12886 (N_12886,N_12698,N_12652);
or U12887 (N_12887,N_12610,N_12615);
nor U12888 (N_12888,N_12630,N_12618);
nor U12889 (N_12889,N_12711,N_12642);
nand U12890 (N_12890,N_12660,N_12543);
nand U12891 (N_12891,N_12671,N_12639);
nand U12892 (N_12892,N_12611,N_12519);
and U12893 (N_12893,N_12745,N_12676);
nor U12894 (N_12894,N_12553,N_12653);
or U12895 (N_12895,N_12714,N_12518);
xor U12896 (N_12896,N_12712,N_12660);
or U12897 (N_12897,N_12660,N_12686);
nor U12898 (N_12898,N_12696,N_12537);
nand U12899 (N_12899,N_12671,N_12596);
nand U12900 (N_12900,N_12602,N_12729);
and U12901 (N_12901,N_12688,N_12706);
xor U12902 (N_12902,N_12561,N_12610);
nor U12903 (N_12903,N_12749,N_12565);
or U12904 (N_12904,N_12650,N_12603);
nor U12905 (N_12905,N_12683,N_12733);
nor U12906 (N_12906,N_12508,N_12705);
nor U12907 (N_12907,N_12687,N_12537);
nor U12908 (N_12908,N_12630,N_12706);
and U12909 (N_12909,N_12592,N_12586);
nand U12910 (N_12910,N_12568,N_12514);
and U12911 (N_12911,N_12652,N_12622);
xnor U12912 (N_12912,N_12625,N_12718);
or U12913 (N_12913,N_12610,N_12531);
or U12914 (N_12914,N_12565,N_12720);
and U12915 (N_12915,N_12557,N_12677);
or U12916 (N_12916,N_12562,N_12515);
xor U12917 (N_12917,N_12679,N_12576);
and U12918 (N_12918,N_12700,N_12552);
nand U12919 (N_12919,N_12656,N_12743);
or U12920 (N_12920,N_12567,N_12543);
and U12921 (N_12921,N_12593,N_12536);
xnor U12922 (N_12922,N_12522,N_12662);
nor U12923 (N_12923,N_12725,N_12635);
and U12924 (N_12924,N_12729,N_12591);
xnor U12925 (N_12925,N_12516,N_12726);
and U12926 (N_12926,N_12577,N_12706);
nand U12927 (N_12927,N_12652,N_12688);
xor U12928 (N_12928,N_12590,N_12629);
nand U12929 (N_12929,N_12703,N_12718);
or U12930 (N_12930,N_12648,N_12543);
nor U12931 (N_12931,N_12599,N_12641);
and U12932 (N_12932,N_12605,N_12727);
nand U12933 (N_12933,N_12535,N_12537);
xor U12934 (N_12934,N_12718,N_12700);
and U12935 (N_12935,N_12654,N_12675);
or U12936 (N_12936,N_12560,N_12530);
nand U12937 (N_12937,N_12522,N_12743);
and U12938 (N_12938,N_12713,N_12620);
nor U12939 (N_12939,N_12693,N_12646);
and U12940 (N_12940,N_12737,N_12552);
or U12941 (N_12941,N_12569,N_12731);
nor U12942 (N_12942,N_12627,N_12560);
and U12943 (N_12943,N_12648,N_12744);
and U12944 (N_12944,N_12632,N_12648);
nor U12945 (N_12945,N_12524,N_12564);
or U12946 (N_12946,N_12666,N_12544);
xor U12947 (N_12947,N_12677,N_12507);
nand U12948 (N_12948,N_12612,N_12608);
and U12949 (N_12949,N_12579,N_12617);
and U12950 (N_12950,N_12609,N_12532);
nor U12951 (N_12951,N_12687,N_12716);
nand U12952 (N_12952,N_12555,N_12596);
xor U12953 (N_12953,N_12611,N_12648);
nor U12954 (N_12954,N_12554,N_12530);
xnor U12955 (N_12955,N_12533,N_12610);
and U12956 (N_12956,N_12673,N_12659);
xnor U12957 (N_12957,N_12654,N_12591);
and U12958 (N_12958,N_12510,N_12649);
or U12959 (N_12959,N_12509,N_12567);
nand U12960 (N_12960,N_12519,N_12550);
and U12961 (N_12961,N_12681,N_12518);
and U12962 (N_12962,N_12607,N_12514);
nor U12963 (N_12963,N_12502,N_12537);
or U12964 (N_12964,N_12561,N_12725);
and U12965 (N_12965,N_12654,N_12719);
nand U12966 (N_12966,N_12723,N_12630);
nand U12967 (N_12967,N_12658,N_12587);
nand U12968 (N_12968,N_12638,N_12547);
or U12969 (N_12969,N_12603,N_12641);
xnor U12970 (N_12970,N_12689,N_12607);
xor U12971 (N_12971,N_12542,N_12577);
nor U12972 (N_12972,N_12592,N_12729);
nand U12973 (N_12973,N_12566,N_12644);
xnor U12974 (N_12974,N_12672,N_12713);
nor U12975 (N_12975,N_12555,N_12653);
nand U12976 (N_12976,N_12629,N_12696);
nand U12977 (N_12977,N_12677,N_12636);
xor U12978 (N_12978,N_12550,N_12561);
nand U12979 (N_12979,N_12563,N_12701);
nor U12980 (N_12980,N_12514,N_12523);
nand U12981 (N_12981,N_12661,N_12662);
or U12982 (N_12982,N_12716,N_12662);
or U12983 (N_12983,N_12638,N_12663);
nor U12984 (N_12984,N_12705,N_12600);
nor U12985 (N_12985,N_12618,N_12559);
nand U12986 (N_12986,N_12729,N_12536);
xor U12987 (N_12987,N_12505,N_12559);
xnor U12988 (N_12988,N_12711,N_12599);
nor U12989 (N_12989,N_12506,N_12646);
and U12990 (N_12990,N_12703,N_12506);
or U12991 (N_12991,N_12506,N_12664);
nand U12992 (N_12992,N_12533,N_12683);
nand U12993 (N_12993,N_12704,N_12558);
or U12994 (N_12994,N_12521,N_12522);
or U12995 (N_12995,N_12696,N_12548);
or U12996 (N_12996,N_12694,N_12660);
xnor U12997 (N_12997,N_12650,N_12550);
or U12998 (N_12998,N_12709,N_12679);
nor U12999 (N_12999,N_12547,N_12739);
nor U13000 (N_13000,N_12843,N_12755);
and U13001 (N_13001,N_12796,N_12926);
nand U13002 (N_13002,N_12813,N_12827);
and U13003 (N_13003,N_12972,N_12801);
xnor U13004 (N_13004,N_12964,N_12971);
xor U13005 (N_13005,N_12780,N_12908);
nand U13006 (N_13006,N_12802,N_12951);
and U13007 (N_13007,N_12935,N_12818);
xnor U13008 (N_13008,N_12900,N_12820);
xnor U13009 (N_13009,N_12917,N_12873);
and U13010 (N_13010,N_12853,N_12916);
nor U13011 (N_13011,N_12757,N_12817);
and U13012 (N_13012,N_12913,N_12952);
nor U13013 (N_13013,N_12875,N_12904);
xnor U13014 (N_13014,N_12840,N_12884);
nand U13015 (N_13015,N_12980,N_12828);
nand U13016 (N_13016,N_12824,N_12992);
nor U13017 (N_13017,N_12805,N_12859);
nor U13018 (N_13018,N_12923,N_12830);
and U13019 (N_13019,N_12890,N_12922);
nand U13020 (N_13020,N_12928,N_12791);
nor U13021 (N_13021,N_12868,N_12879);
and U13022 (N_13022,N_12927,N_12940);
nor U13023 (N_13023,N_12774,N_12835);
or U13024 (N_13024,N_12938,N_12787);
xor U13025 (N_13025,N_12858,N_12999);
nor U13026 (N_13026,N_12931,N_12763);
xor U13027 (N_13027,N_12845,N_12960);
nor U13028 (N_13028,N_12867,N_12915);
xor U13029 (N_13029,N_12956,N_12885);
and U13030 (N_13030,N_12783,N_12982);
or U13031 (N_13031,N_12771,N_12969);
xor U13032 (N_13032,N_12932,N_12930);
xor U13033 (N_13033,N_12959,N_12761);
or U13034 (N_13034,N_12785,N_12881);
xnor U13035 (N_13035,N_12987,N_12997);
and U13036 (N_13036,N_12961,N_12897);
nor U13037 (N_13037,N_12955,N_12841);
xnor U13038 (N_13038,N_12754,N_12814);
or U13039 (N_13039,N_12750,N_12979);
nand U13040 (N_13040,N_12810,N_12962);
nand U13041 (N_13041,N_12883,N_12918);
and U13042 (N_13042,N_12949,N_12842);
and U13043 (N_13043,N_12872,N_12983);
or U13044 (N_13044,N_12948,N_12989);
nand U13045 (N_13045,N_12766,N_12793);
xnor U13046 (N_13046,N_12756,N_12770);
or U13047 (N_13047,N_12933,N_12986);
nand U13048 (N_13048,N_12823,N_12870);
nor U13049 (N_13049,N_12907,N_12804);
and U13050 (N_13050,N_12894,N_12806);
and U13051 (N_13051,N_12994,N_12963);
xnor U13052 (N_13052,N_12899,N_12795);
and U13053 (N_13053,N_12786,N_12919);
and U13054 (N_13054,N_12906,N_12968);
and U13055 (N_13055,N_12778,N_12798);
nand U13056 (N_13056,N_12874,N_12880);
nor U13057 (N_13057,N_12887,N_12993);
xnor U13058 (N_13058,N_12811,N_12844);
or U13059 (N_13059,N_12941,N_12839);
xor U13060 (N_13060,N_12779,N_12910);
nor U13061 (N_13061,N_12767,N_12914);
or U13062 (N_13062,N_12772,N_12769);
xor U13063 (N_13063,N_12996,N_12800);
nand U13064 (N_13064,N_12816,N_12808);
nand U13065 (N_13065,N_12762,N_12945);
and U13066 (N_13066,N_12865,N_12891);
and U13067 (N_13067,N_12975,N_12847);
or U13068 (N_13068,N_12998,N_12825);
and U13069 (N_13069,N_12849,N_12947);
or U13070 (N_13070,N_12995,N_12833);
nor U13071 (N_13071,N_12812,N_12792);
nor U13072 (N_13072,N_12892,N_12958);
or U13073 (N_13073,N_12777,N_12773);
xor U13074 (N_13074,N_12768,N_12782);
nor U13075 (N_13075,N_12936,N_12861);
or U13076 (N_13076,N_12909,N_12781);
nor U13077 (N_13077,N_12759,N_12834);
nor U13078 (N_13078,N_12966,N_12753);
nand U13079 (N_13079,N_12974,N_12856);
nor U13080 (N_13080,N_12882,N_12784);
xor U13081 (N_13081,N_12752,N_12889);
or U13082 (N_13082,N_12967,N_12826);
xnor U13083 (N_13083,N_12819,N_12850);
nand U13084 (N_13084,N_12985,N_12758);
xor U13085 (N_13085,N_12976,N_12898);
or U13086 (N_13086,N_12803,N_12886);
xnor U13087 (N_13087,N_12977,N_12807);
or U13088 (N_13088,N_12829,N_12765);
xor U13089 (N_13089,N_12981,N_12838);
nor U13090 (N_13090,N_12855,N_12944);
xor U13091 (N_13091,N_12866,N_12821);
xnor U13092 (N_13092,N_12937,N_12954);
and U13093 (N_13093,N_12878,N_12776);
nand U13094 (N_13094,N_12905,N_12920);
xnor U13095 (N_13095,N_12871,N_12901);
nor U13096 (N_13096,N_12903,N_12965);
nor U13097 (N_13097,N_12921,N_12854);
and U13098 (N_13098,N_12895,N_12876);
or U13099 (N_13099,N_12822,N_12877);
xor U13100 (N_13100,N_12809,N_12863);
and U13101 (N_13101,N_12831,N_12832);
xnor U13102 (N_13102,N_12925,N_12851);
nand U13103 (N_13103,N_12988,N_12764);
or U13104 (N_13104,N_12862,N_12751);
xor U13105 (N_13105,N_12837,N_12973);
xor U13106 (N_13106,N_12939,N_12797);
and U13107 (N_13107,N_12911,N_12864);
nand U13108 (N_13108,N_12815,N_12946);
nor U13109 (N_13109,N_12943,N_12990);
nor U13110 (N_13110,N_12789,N_12775);
xnor U13111 (N_13111,N_12934,N_12857);
xnor U13112 (N_13112,N_12846,N_12978);
nand U13113 (N_13113,N_12893,N_12788);
or U13114 (N_13114,N_12950,N_12860);
and U13115 (N_13115,N_12984,N_12799);
and U13116 (N_13116,N_12836,N_12848);
or U13117 (N_13117,N_12991,N_12760);
and U13118 (N_13118,N_12852,N_12902);
xor U13119 (N_13119,N_12953,N_12912);
or U13120 (N_13120,N_12790,N_12970);
nor U13121 (N_13121,N_12888,N_12896);
nand U13122 (N_13122,N_12869,N_12929);
or U13123 (N_13123,N_12957,N_12942);
nand U13124 (N_13124,N_12924,N_12794);
xnor U13125 (N_13125,N_12802,N_12824);
nand U13126 (N_13126,N_12907,N_12979);
xor U13127 (N_13127,N_12850,N_12800);
xor U13128 (N_13128,N_12806,N_12762);
and U13129 (N_13129,N_12895,N_12943);
nor U13130 (N_13130,N_12832,N_12946);
nand U13131 (N_13131,N_12926,N_12801);
nand U13132 (N_13132,N_12996,N_12831);
nand U13133 (N_13133,N_12871,N_12783);
xor U13134 (N_13134,N_12893,N_12967);
nor U13135 (N_13135,N_12842,N_12773);
xor U13136 (N_13136,N_12911,N_12991);
or U13137 (N_13137,N_12903,N_12871);
nand U13138 (N_13138,N_12948,N_12886);
xnor U13139 (N_13139,N_12771,N_12765);
and U13140 (N_13140,N_12783,N_12958);
and U13141 (N_13141,N_12781,N_12970);
and U13142 (N_13142,N_12921,N_12881);
and U13143 (N_13143,N_12835,N_12949);
nand U13144 (N_13144,N_12900,N_12931);
and U13145 (N_13145,N_12919,N_12856);
and U13146 (N_13146,N_12814,N_12854);
or U13147 (N_13147,N_12835,N_12974);
nand U13148 (N_13148,N_12827,N_12836);
nand U13149 (N_13149,N_12792,N_12872);
nand U13150 (N_13150,N_12924,N_12958);
xnor U13151 (N_13151,N_12981,N_12811);
and U13152 (N_13152,N_12815,N_12795);
nor U13153 (N_13153,N_12893,N_12765);
and U13154 (N_13154,N_12835,N_12929);
nand U13155 (N_13155,N_12816,N_12894);
nor U13156 (N_13156,N_12901,N_12977);
or U13157 (N_13157,N_12888,N_12866);
and U13158 (N_13158,N_12843,N_12863);
or U13159 (N_13159,N_12793,N_12773);
or U13160 (N_13160,N_12857,N_12762);
nand U13161 (N_13161,N_12888,N_12750);
nand U13162 (N_13162,N_12758,N_12950);
xnor U13163 (N_13163,N_12852,N_12971);
nor U13164 (N_13164,N_12906,N_12845);
or U13165 (N_13165,N_12937,N_12853);
nor U13166 (N_13166,N_12964,N_12918);
nor U13167 (N_13167,N_12815,N_12842);
and U13168 (N_13168,N_12870,N_12814);
and U13169 (N_13169,N_12853,N_12874);
nor U13170 (N_13170,N_12864,N_12958);
and U13171 (N_13171,N_12785,N_12981);
nor U13172 (N_13172,N_12857,N_12873);
and U13173 (N_13173,N_12902,N_12884);
and U13174 (N_13174,N_12838,N_12753);
or U13175 (N_13175,N_12766,N_12803);
and U13176 (N_13176,N_12755,N_12948);
nor U13177 (N_13177,N_12772,N_12849);
or U13178 (N_13178,N_12775,N_12948);
nand U13179 (N_13179,N_12991,N_12947);
and U13180 (N_13180,N_12892,N_12874);
nand U13181 (N_13181,N_12820,N_12905);
nand U13182 (N_13182,N_12774,N_12977);
and U13183 (N_13183,N_12911,N_12886);
and U13184 (N_13184,N_12801,N_12776);
xor U13185 (N_13185,N_12875,N_12804);
nand U13186 (N_13186,N_12785,N_12851);
nand U13187 (N_13187,N_12809,N_12920);
and U13188 (N_13188,N_12780,N_12861);
and U13189 (N_13189,N_12775,N_12991);
xnor U13190 (N_13190,N_12818,N_12763);
xor U13191 (N_13191,N_12921,N_12898);
xnor U13192 (N_13192,N_12932,N_12755);
or U13193 (N_13193,N_12765,N_12960);
nand U13194 (N_13194,N_12988,N_12849);
xor U13195 (N_13195,N_12996,N_12763);
and U13196 (N_13196,N_12789,N_12810);
and U13197 (N_13197,N_12867,N_12871);
or U13198 (N_13198,N_12878,N_12830);
and U13199 (N_13199,N_12855,N_12985);
nand U13200 (N_13200,N_12936,N_12891);
nand U13201 (N_13201,N_12769,N_12950);
nor U13202 (N_13202,N_12855,N_12913);
and U13203 (N_13203,N_12878,N_12992);
nand U13204 (N_13204,N_12964,N_12767);
or U13205 (N_13205,N_12977,N_12809);
or U13206 (N_13206,N_12851,N_12982);
and U13207 (N_13207,N_12751,N_12915);
nand U13208 (N_13208,N_12863,N_12845);
and U13209 (N_13209,N_12860,N_12972);
or U13210 (N_13210,N_12879,N_12835);
and U13211 (N_13211,N_12785,N_12928);
nand U13212 (N_13212,N_12911,N_12814);
and U13213 (N_13213,N_12833,N_12952);
nand U13214 (N_13214,N_12796,N_12916);
xor U13215 (N_13215,N_12766,N_12781);
nand U13216 (N_13216,N_12857,N_12832);
nor U13217 (N_13217,N_12808,N_12938);
or U13218 (N_13218,N_12884,N_12893);
or U13219 (N_13219,N_12778,N_12937);
and U13220 (N_13220,N_12975,N_12958);
nand U13221 (N_13221,N_12913,N_12889);
nand U13222 (N_13222,N_12869,N_12984);
or U13223 (N_13223,N_12984,N_12861);
and U13224 (N_13224,N_12938,N_12962);
and U13225 (N_13225,N_12862,N_12857);
or U13226 (N_13226,N_12830,N_12823);
nor U13227 (N_13227,N_12860,N_12850);
and U13228 (N_13228,N_12924,N_12875);
nor U13229 (N_13229,N_12789,N_12865);
nand U13230 (N_13230,N_12926,N_12883);
and U13231 (N_13231,N_12780,N_12798);
nor U13232 (N_13232,N_12799,N_12888);
or U13233 (N_13233,N_12831,N_12972);
or U13234 (N_13234,N_12831,N_12788);
xnor U13235 (N_13235,N_12880,N_12862);
nor U13236 (N_13236,N_12855,N_12867);
xnor U13237 (N_13237,N_12916,N_12941);
or U13238 (N_13238,N_12811,N_12781);
and U13239 (N_13239,N_12952,N_12904);
or U13240 (N_13240,N_12869,N_12943);
xor U13241 (N_13241,N_12821,N_12842);
or U13242 (N_13242,N_12950,N_12929);
and U13243 (N_13243,N_12833,N_12906);
nor U13244 (N_13244,N_12802,N_12980);
nor U13245 (N_13245,N_12974,N_12826);
or U13246 (N_13246,N_12819,N_12763);
and U13247 (N_13247,N_12826,N_12991);
or U13248 (N_13248,N_12757,N_12892);
nand U13249 (N_13249,N_12826,N_12892);
nand U13250 (N_13250,N_13165,N_13053);
nor U13251 (N_13251,N_13003,N_13075);
or U13252 (N_13252,N_13193,N_13178);
nor U13253 (N_13253,N_13226,N_13006);
and U13254 (N_13254,N_13026,N_13141);
nand U13255 (N_13255,N_13198,N_13190);
and U13256 (N_13256,N_13179,N_13248);
nor U13257 (N_13257,N_13132,N_13123);
and U13258 (N_13258,N_13192,N_13052);
or U13259 (N_13259,N_13022,N_13169);
nand U13260 (N_13260,N_13019,N_13078);
or U13261 (N_13261,N_13045,N_13105);
xnor U13262 (N_13262,N_13089,N_13103);
xnor U13263 (N_13263,N_13016,N_13166);
xor U13264 (N_13264,N_13100,N_13073);
or U13265 (N_13265,N_13180,N_13076);
and U13266 (N_13266,N_13015,N_13200);
xor U13267 (N_13267,N_13236,N_13098);
xor U13268 (N_13268,N_13229,N_13051);
or U13269 (N_13269,N_13168,N_13138);
and U13270 (N_13270,N_13159,N_13188);
or U13271 (N_13271,N_13243,N_13149);
nor U13272 (N_13272,N_13207,N_13066);
nor U13273 (N_13273,N_13143,N_13010);
nand U13274 (N_13274,N_13222,N_13114);
and U13275 (N_13275,N_13044,N_13212);
nor U13276 (N_13276,N_13218,N_13032);
xor U13277 (N_13277,N_13187,N_13118);
and U13278 (N_13278,N_13213,N_13217);
xor U13279 (N_13279,N_13077,N_13033);
and U13280 (N_13280,N_13202,N_13230);
nand U13281 (N_13281,N_13063,N_13086);
nand U13282 (N_13282,N_13119,N_13020);
nand U13283 (N_13283,N_13094,N_13203);
and U13284 (N_13284,N_13129,N_13151);
nand U13285 (N_13285,N_13241,N_13096);
or U13286 (N_13286,N_13081,N_13012);
xnor U13287 (N_13287,N_13001,N_13112);
or U13288 (N_13288,N_13087,N_13232);
nand U13289 (N_13289,N_13150,N_13201);
and U13290 (N_13290,N_13237,N_13133);
nor U13291 (N_13291,N_13054,N_13014);
or U13292 (N_13292,N_13195,N_13072);
and U13293 (N_13293,N_13153,N_13034);
nand U13294 (N_13294,N_13035,N_13139);
and U13295 (N_13295,N_13070,N_13172);
and U13296 (N_13296,N_13167,N_13244);
xor U13297 (N_13297,N_13131,N_13067);
xnor U13298 (N_13298,N_13102,N_13116);
nor U13299 (N_13299,N_13093,N_13204);
xor U13300 (N_13300,N_13161,N_13110);
nand U13301 (N_13301,N_13227,N_13005);
nor U13302 (N_13302,N_13109,N_13068);
xor U13303 (N_13303,N_13041,N_13108);
and U13304 (N_13304,N_13199,N_13158);
or U13305 (N_13305,N_13145,N_13206);
xnor U13306 (N_13306,N_13043,N_13029);
or U13307 (N_13307,N_13017,N_13249);
and U13308 (N_13308,N_13160,N_13059);
nor U13309 (N_13309,N_13128,N_13058);
nor U13310 (N_13310,N_13027,N_13121);
nand U13311 (N_13311,N_13231,N_13113);
nor U13312 (N_13312,N_13175,N_13173);
nor U13313 (N_13313,N_13009,N_13126);
xnor U13314 (N_13314,N_13211,N_13214);
nor U13315 (N_13315,N_13221,N_13071);
nand U13316 (N_13316,N_13127,N_13185);
and U13317 (N_13317,N_13194,N_13013);
nor U13318 (N_13318,N_13197,N_13162);
nand U13319 (N_13319,N_13239,N_13007);
nand U13320 (N_13320,N_13177,N_13082);
nor U13321 (N_13321,N_13042,N_13025);
or U13322 (N_13322,N_13124,N_13137);
nor U13323 (N_13323,N_13216,N_13233);
and U13324 (N_13324,N_13083,N_13021);
xor U13325 (N_13325,N_13140,N_13235);
and U13326 (N_13326,N_13208,N_13156);
or U13327 (N_13327,N_13215,N_13092);
nand U13328 (N_13328,N_13000,N_13189);
nand U13329 (N_13329,N_13101,N_13060);
xor U13330 (N_13330,N_13247,N_13023);
nor U13331 (N_13331,N_13040,N_13048);
nor U13332 (N_13332,N_13182,N_13245);
or U13333 (N_13333,N_13024,N_13135);
and U13334 (N_13334,N_13240,N_13142);
xnor U13335 (N_13335,N_13164,N_13008);
nand U13336 (N_13336,N_13111,N_13031);
nand U13337 (N_13337,N_13157,N_13064);
and U13338 (N_13338,N_13223,N_13062);
nor U13339 (N_13339,N_13039,N_13147);
and U13340 (N_13340,N_13011,N_13125);
nor U13341 (N_13341,N_13099,N_13028);
or U13342 (N_13342,N_13057,N_13036);
and U13343 (N_13343,N_13224,N_13107);
xnor U13344 (N_13344,N_13065,N_13205);
xnor U13345 (N_13345,N_13242,N_13069);
nand U13346 (N_13346,N_13183,N_13037);
nand U13347 (N_13347,N_13080,N_13209);
xnor U13348 (N_13348,N_13134,N_13246);
xor U13349 (N_13349,N_13152,N_13046);
xnor U13350 (N_13350,N_13038,N_13163);
xnor U13351 (N_13351,N_13084,N_13154);
or U13352 (N_13352,N_13181,N_13155);
and U13353 (N_13353,N_13079,N_13117);
or U13354 (N_13354,N_13146,N_13136);
or U13355 (N_13355,N_13106,N_13238);
nand U13356 (N_13356,N_13091,N_13191);
and U13357 (N_13357,N_13088,N_13170);
xnor U13358 (N_13358,N_13002,N_13030);
or U13359 (N_13359,N_13115,N_13004);
nand U13360 (N_13360,N_13196,N_13050);
xor U13361 (N_13361,N_13104,N_13228);
nand U13362 (N_13362,N_13122,N_13210);
or U13363 (N_13363,N_13234,N_13061);
nor U13364 (N_13364,N_13018,N_13049);
or U13365 (N_13365,N_13220,N_13176);
or U13366 (N_13366,N_13120,N_13144);
and U13367 (N_13367,N_13055,N_13186);
or U13368 (N_13368,N_13171,N_13219);
nor U13369 (N_13369,N_13184,N_13074);
or U13370 (N_13370,N_13174,N_13097);
xnor U13371 (N_13371,N_13148,N_13130);
xor U13372 (N_13372,N_13085,N_13225);
and U13373 (N_13373,N_13056,N_13047);
nor U13374 (N_13374,N_13090,N_13095);
nor U13375 (N_13375,N_13035,N_13022);
and U13376 (N_13376,N_13226,N_13235);
xnor U13377 (N_13377,N_13113,N_13180);
nor U13378 (N_13378,N_13120,N_13031);
and U13379 (N_13379,N_13218,N_13190);
nor U13380 (N_13380,N_13029,N_13154);
or U13381 (N_13381,N_13118,N_13151);
nand U13382 (N_13382,N_13173,N_13249);
nor U13383 (N_13383,N_13137,N_13195);
nor U13384 (N_13384,N_13064,N_13076);
and U13385 (N_13385,N_13245,N_13154);
and U13386 (N_13386,N_13232,N_13092);
nor U13387 (N_13387,N_13168,N_13203);
and U13388 (N_13388,N_13113,N_13143);
or U13389 (N_13389,N_13084,N_13215);
or U13390 (N_13390,N_13222,N_13241);
or U13391 (N_13391,N_13134,N_13219);
or U13392 (N_13392,N_13041,N_13224);
nor U13393 (N_13393,N_13087,N_13136);
and U13394 (N_13394,N_13234,N_13191);
nor U13395 (N_13395,N_13147,N_13001);
xnor U13396 (N_13396,N_13112,N_13024);
nor U13397 (N_13397,N_13241,N_13167);
nor U13398 (N_13398,N_13008,N_13174);
or U13399 (N_13399,N_13101,N_13104);
and U13400 (N_13400,N_13127,N_13087);
or U13401 (N_13401,N_13116,N_13240);
xnor U13402 (N_13402,N_13100,N_13242);
nor U13403 (N_13403,N_13211,N_13174);
and U13404 (N_13404,N_13013,N_13079);
or U13405 (N_13405,N_13150,N_13066);
or U13406 (N_13406,N_13003,N_13157);
and U13407 (N_13407,N_13167,N_13140);
and U13408 (N_13408,N_13215,N_13118);
nand U13409 (N_13409,N_13201,N_13119);
xor U13410 (N_13410,N_13154,N_13050);
and U13411 (N_13411,N_13226,N_13120);
nand U13412 (N_13412,N_13123,N_13041);
nand U13413 (N_13413,N_13234,N_13146);
xnor U13414 (N_13414,N_13177,N_13065);
nand U13415 (N_13415,N_13024,N_13001);
nor U13416 (N_13416,N_13044,N_13071);
nor U13417 (N_13417,N_13193,N_13079);
or U13418 (N_13418,N_13105,N_13155);
nor U13419 (N_13419,N_13246,N_13003);
or U13420 (N_13420,N_13228,N_13025);
or U13421 (N_13421,N_13205,N_13237);
or U13422 (N_13422,N_13182,N_13176);
nor U13423 (N_13423,N_13109,N_13059);
or U13424 (N_13424,N_13206,N_13171);
nor U13425 (N_13425,N_13096,N_13081);
nor U13426 (N_13426,N_13135,N_13241);
or U13427 (N_13427,N_13007,N_13037);
and U13428 (N_13428,N_13018,N_13159);
xnor U13429 (N_13429,N_13181,N_13152);
or U13430 (N_13430,N_13072,N_13171);
and U13431 (N_13431,N_13121,N_13025);
nor U13432 (N_13432,N_13119,N_13228);
xnor U13433 (N_13433,N_13198,N_13195);
or U13434 (N_13434,N_13187,N_13084);
nor U13435 (N_13435,N_13179,N_13171);
or U13436 (N_13436,N_13208,N_13222);
nand U13437 (N_13437,N_13068,N_13029);
and U13438 (N_13438,N_13092,N_13076);
or U13439 (N_13439,N_13249,N_13186);
nand U13440 (N_13440,N_13092,N_13123);
xnor U13441 (N_13441,N_13099,N_13163);
xnor U13442 (N_13442,N_13080,N_13083);
nand U13443 (N_13443,N_13120,N_13211);
nor U13444 (N_13444,N_13092,N_13235);
and U13445 (N_13445,N_13094,N_13075);
and U13446 (N_13446,N_13249,N_13095);
nand U13447 (N_13447,N_13100,N_13231);
nor U13448 (N_13448,N_13122,N_13216);
xnor U13449 (N_13449,N_13115,N_13007);
or U13450 (N_13450,N_13136,N_13133);
or U13451 (N_13451,N_13190,N_13015);
xnor U13452 (N_13452,N_13106,N_13047);
nand U13453 (N_13453,N_13233,N_13065);
nor U13454 (N_13454,N_13021,N_13012);
xor U13455 (N_13455,N_13086,N_13100);
and U13456 (N_13456,N_13206,N_13107);
and U13457 (N_13457,N_13207,N_13007);
nand U13458 (N_13458,N_13031,N_13177);
xnor U13459 (N_13459,N_13206,N_13057);
nor U13460 (N_13460,N_13028,N_13088);
or U13461 (N_13461,N_13185,N_13239);
xor U13462 (N_13462,N_13098,N_13040);
or U13463 (N_13463,N_13172,N_13228);
or U13464 (N_13464,N_13120,N_13143);
or U13465 (N_13465,N_13156,N_13158);
and U13466 (N_13466,N_13013,N_13131);
or U13467 (N_13467,N_13062,N_13011);
nor U13468 (N_13468,N_13029,N_13102);
xor U13469 (N_13469,N_13240,N_13077);
xor U13470 (N_13470,N_13101,N_13241);
nor U13471 (N_13471,N_13210,N_13192);
nor U13472 (N_13472,N_13033,N_13199);
nor U13473 (N_13473,N_13216,N_13115);
and U13474 (N_13474,N_13135,N_13157);
nand U13475 (N_13475,N_13132,N_13138);
xor U13476 (N_13476,N_13194,N_13041);
or U13477 (N_13477,N_13003,N_13055);
xor U13478 (N_13478,N_13145,N_13242);
nor U13479 (N_13479,N_13218,N_13024);
or U13480 (N_13480,N_13045,N_13226);
nand U13481 (N_13481,N_13207,N_13155);
and U13482 (N_13482,N_13143,N_13240);
and U13483 (N_13483,N_13189,N_13151);
or U13484 (N_13484,N_13245,N_13093);
nand U13485 (N_13485,N_13238,N_13204);
or U13486 (N_13486,N_13245,N_13243);
nor U13487 (N_13487,N_13011,N_13024);
nor U13488 (N_13488,N_13205,N_13167);
and U13489 (N_13489,N_13151,N_13234);
nand U13490 (N_13490,N_13219,N_13211);
or U13491 (N_13491,N_13042,N_13064);
or U13492 (N_13492,N_13160,N_13216);
nand U13493 (N_13493,N_13120,N_13033);
and U13494 (N_13494,N_13247,N_13011);
or U13495 (N_13495,N_13187,N_13002);
or U13496 (N_13496,N_13235,N_13026);
xor U13497 (N_13497,N_13042,N_13109);
nor U13498 (N_13498,N_13179,N_13169);
xnor U13499 (N_13499,N_13181,N_13082);
nand U13500 (N_13500,N_13364,N_13325);
nand U13501 (N_13501,N_13370,N_13338);
xnor U13502 (N_13502,N_13323,N_13394);
and U13503 (N_13503,N_13253,N_13282);
nor U13504 (N_13504,N_13342,N_13330);
nand U13505 (N_13505,N_13475,N_13358);
nor U13506 (N_13506,N_13402,N_13303);
xor U13507 (N_13507,N_13256,N_13318);
xnor U13508 (N_13508,N_13322,N_13365);
nor U13509 (N_13509,N_13388,N_13363);
xnor U13510 (N_13510,N_13422,N_13468);
nand U13511 (N_13511,N_13435,N_13446);
or U13512 (N_13512,N_13272,N_13430);
and U13513 (N_13513,N_13448,N_13336);
nand U13514 (N_13514,N_13382,N_13254);
nand U13515 (N_13515,N_13319,N_13310);
nor U13516 (N_13516,N_13437,N_13315);
nand U13517 (N_13517,N_13465,N_13384);
nand U13518 (N_13518,N_13295,N_13376);
nand U13519 (N_13519,N_13387,N_13467);
nor U13520 (N_13520,N_13423,N_13334);
and U13521 (N_13521,N_13415,N_13458);
nand U13522 (N_13522,N_13417,N_13317);
and U13523 (N_13523,N_13309,N_13476);
nor U13524 (N_13524,N_13487,N_13378);
nor U13525 (N_13525,N_13414,N_13287);
xor U13526 (N_13526,N_13486,N_13490);
nor U13527 (N_13527,N_13445,N_13447);
xor U13528 (N_13528,N_13259,N_13499);
nor U13529 (N_13529,N_13485,N_13369);
nand U13530 (N_13530,N_13297,N_13452);
or U13531 (N_13531,N_13328,N_13283);
xnor U13532 (N_13532,N_13301,N_13280);
nand U13533 (N_13533,N_13398,N_13492);
nand U13534 (N_13534,N_13366,N_13434);
xnor U13535 (N_13535,N_13260,N_13279);
nor U13536 (N_13536,N_13483,N_13353);
and U13537 (N_13537,N_13333,N_13292);
and U13538 (N_13538,N_13294,N_13305);
and U13539 (N_13539,N_13379,N_13290);
or U13540 (N_13540,N_13455,N_13472);
or U13541 (N_13541,N_13413,N_13493);
or U13542 (N_13542,N_13262,N_13329);
nand U13543 (N_13543,N_13479,N_13419);
xor U13544 (N_13544,N_13488,N_13278);
or U13545 (N_13545,N_13444,N_13339);
or U13546 (N_13546,N_13420,N_13450);
and U13547 (N_13547,N_13474,N_13425);
nand U13548 (N_13548,N_13346,N_13307);
or U13549 (N_13549,N_13274,N_13473);
or U13550 (N_13550,N_13288,N_13306);
or U13551 (N_13551,N_13314,N_13457);
and U13552 (N_13552,N_13498,N_13456);
nand U13553 (N_13553,N_13408,N_13374);
or U13554 (N_13554,N_13371,N_13271);
and U13555 (N_13555,N_13392,N_13257);
and U13556 (N_13556,N_13421,N_13316);
xnor U13557 (N_13557,N_13349,N_13407);
and U13558 (N_13558,N_13470,N_13404);
and U13559 (N_13559,N_13442,N_13480);
xor U13560 (N_13560,N_13321,N_13469);
and U13561 (N_13561,N_13296,N_13424);
nor U13562 (N_13562,N_13443,N_13350);
nor U13563 (N_13563,N_13357,N_13405);
xnor U13564 (N_13564,N_13362,N_13428);
nand U13565 (N_13565,N_13471,N_13386);
nor U13566 (N_13566,N_13289,N_13418);
and U13567 (N_13567,N_13453,N_13494);
and U13568 (N_13568,N_13416,N_13396);
nor U13569 (N_13569,N_13304,N_13466);
xnor U13570 (N_13570,N_13460,N_13343);
and U13571 (N_13571,N_13258,N_13263);
nor U13572 (N_13572,N_13373,N_13478);
and U13573 (N_13573,N_13348,N_13462);
nor U13574 (N_13574,N_13385,N_13451);
nand U13575 (N_13575,N_13463,N_13332);
nand U13576 (N_13576,N_13293,N_13335);
nor U13577 (N_13577,N_13308,N_13433);
or U13578 (N_13578,N_13352,N_13496);
and U13579 (N_13579,N_13432,N_13380);
or U13580 (N_13580,N_13497,N_13341);
and U13581 (N_13581,N_13381,N_13266);
and U13582 (N_13582,N_13397,N_13372);
and U13583 (N_13583,N_13354,N_13410);
xor U13584 (N_13584,N_13454,N_13267);
and U13585 (N_13585,N_13277,N_13383);
xnor U13586 (N_13586,N_13252,N_13284);
and U13587 (N_13587,N_13409,N_13298);
nand U13588 (N_13588,N_13440,N_13337);
and U13589 (N_13589,N_13355,N_13389);
or U13590 (N_13590,N_13411,N_13312);
or U13591 (N_13591,N_13461,N_13464);
nor U13592 (N_13592,N_13438,N_13436);
nor U13593 (N_13593,N_13300,N_13406);
or U13594 (N_13594,N_13481,N_13359);
xor U13595 (N_13595,N_13484,N_13400);
and U13596 (N_13596,N_13285,N_13347);
nand U13597 (N_13597,N_13491,N_13340);
and U13598 (N_13598,N_13269,N_13495);
nor U13599 (N_13599,N_13412,N_13361);
nand U13600 (N_13600,N_13401,N_13331);
or U13601 (N_13601,N_13320,N_13395);
xor U13602 (N_13602,N_13275,N_13276);
xnor U13603 (N_13603,N_13391,N_13281);
or U13604 (N_13604,N_13393,N_13250);
and U13605 (N_13605,N_13449,N_13268);
and U13606 (N_13606,N_13356,N_13324);
nor U13607 (N_13607,N_13368,N_13313);
xnor U13608 (N_13608,N_13431,N_13477);
xor U13609 (N_13609,N_13426,N_13327);
and U13610 (N_13610,N_13264,N_13482);
nand U13611 (N_13611,N_13367,N_13286);
or U13612 (N_13612,N_13302,N_13360);
xnor U13613 (N_13613,N_13427,N_13390);
and U13614 (N_13614,N_13429,N_13344);
or U13615 (N_13615,N_13441,N_13261);
nand U13616 (N_13616,N_13377,N_13291);
and U13617 (N_13617,N_13299,N_13403);
or U13618 (N_13618,N_13345,N_13270);
or U13619 (N_13619,N_13489,N_13255);
xor U13620 (N_13620,N_13459,N_13399);
nand U13621 (N_13621,N_13375,N_13439);
or U13622 (N_13622,N_13265,N_13326);
and U13623 (N_13623,N_13273,N_13311);
nor U13624 (N_13624,N_13251,N_13351);
xnor U13625 (N_13625,N_13343,N_13361);
nand U13626 (N_13626,N_13490,N_13291);
or U13627 (N_13627,N_13328,N_13300);
or U13628 (N_13628,N_13301,N_13471);
xor U13629 (N_13629,N_13354,N_13355);
nor U13630 (N_13630,N_13303,N_13311);
or U13631 (N_13631,N_13488,N_13401);
or U13632 (N_13632,N_13272,N_13464);
nor U13633 (N_13633,N_13264,N_13485);
nand U13634 (N_13634,N_13321,N_13460);
nor U13635 (N_13635,N_13382,N_13401);
nand U13636 (N_13636,N_13497,N_13462);
xor U13637 (N_13637,N_13414,N_13459);
nand U13638 (N_13638,N_13421,N_13463);
or U13639 (N_13639,N_13267,N_13293);
nor U13640 (N_13640,N_13321,N_13433);
or U13641 (N_13641,N_13369,N_13291);
or U13642 (N_13642,N_13439,N_13277);
xnor U13643 (N_13643,N_13392,N_13357);
xnor U13644 (N_13644,N_13343,N_13253);
nor U13645 (N_13645,N_13286,N_13254);
nand U13646 (N_13646,N_13485,N_13275);
and U13647 (N_13647,N_13465,N_13309);
or U13648 (N_13648,N_13286,N_13289);
xnor U13649 (N_13649,N_13256,N_13388);
or U13650 (N_13650,N_13346,N_13279);
or U13651 (N_13651,N_13277,N_13491);
or U13652 (N_13652,N_13494,N_13287);
nand U13653 (N_13653,N_13313,N_13438);
xor U13654 (N_13654,N_13346,N_13316);
and U13655 (N_13655,N_13283,N_13325);
and U13656 (N_13656,N_13393,N_13380);
nand U13657 (N_13657,N_13313,N_13304);
nand U13658 (N_13658,N_13436,N_13402);
xor U13659 (N_13659,N_13461,N_13317);
and U13660 (N_13660,N_13414,N_13461);
or U13661 (N_13661,N_13401,N_13306);
xor U13662 (N_13662,N_13270,N_13306);
xnor U13663 (N_13663,N_13483,N_13300);
xor U13664 (N_13664,N_13416,N_13451);
nor U13665 (N_13665,N_13330,N_13451);
nand U13666 (N_13666,N_13494,N_13286);
and U13667 (N_13667,N_13263,N_13356);
and U13668 (N_13668,N_13378,N_13278);
and U13669 (N_13669,N_13418,N_13349);
and U13670 (N_13670,N_13472,N_13257);
nand U13671 (N_13671,N_13250,N_13495);
nor U13672 (N_13672,N_13296,N_13374);
xor U13673 (N_13673,N_13480,N_13401);
xor U13674 (N_13674,N_13424,N_13326);
and U13675 (N_13675,N_13344,N_13461);
xnor U13676 (N_13676,N_13427,N_13304);
or U13677 (N_13677,N_13491,N_13444);
nand U13678 (N_13678,N_13367,N_13467);
xor U13679 (N_13679,N_13345,N_13283);
and U13680 (N_13680,N_13410,N_13284);
or U13681 (N_13681,N_13367,N_13385);
xor U13682 (N_13682,N_13258,N_13393);
nand U13683 (N_13683,N_13495,N_13451);
and U13684 (N_13684,N_13356,N_13450);
nand U13685 (N_13685,N_13255,N_13331);
xnor U13686 (N_13686,N_13396,N_13402);
nor U13687 (N_13687,N_13450,N_13263);
and U13688 (N_13688,N_13435,N_13406);
or U13689 (N_13689,N_13492,N_13362);
xnor U13690 (N_13690,N_13263,N_13459);
xor U13691 (N_13691,N_13442,N_13264);
nor U13692 (N_13692,N_13254,N_13299);
and U13693 (N_13693,N_13310,N_13296);
nor U13694 (N_13694,N_13457,N_13268);
nand U13695 (N_13695,N_13455,N_13300);
nand U13696 (N_13696,N_13331,N_13300);
xor U13697 (N_13697,N_13455,N_13418);
or U13698 (N_13698,N_13297,N_13305);
nand U13699 (N_13699,N_13309,N_13342);
xnor U13700 (N_13700,N_13469,N_13250);
xnor U13701 (N_13701,N_13463,N_13425);
nand U13702 (N_13702,N_13394,N_13377);
and U13703 (N_13703,N_13313,N_13355);
and U13704 (N_13704,N_13493,N_13475);
and U13705 (N_13705,N_13368,N_13383);
nand U13706 (N_13706,N_13313,N_13424);
xor U13707 (N_13707,N_13403,N_13428);
nand U13708 (N_13708,N_13358,N_13324);
nand U13709 (N_13709,N_13478,N_13381);
nor U13710 (N_13710,N_13338,N_13484);
or U13711 (N_13711,N_13368,N_13467);
and U13712 (N_13712,N_13411,N_13405);
xnor U13713 (N_13713,N_13285,N_13461);
nor U13714 (N_13714,N_13424,N_13421);
xnor U13715 (N_13715,N_13283,N_13347);
nor U13716 (N_13716,N_13379,N_13445);
or U13717 (N_13717,N_13345,N_13442);
nand U13718 (N_13718,N_13296,N_13371);
and U13719 (N_13719,N_13466,N_13277);
nand U13720 (N_13720,N_13423,N_13403);
xnor U13721 (N_13721,N_13442,N_13343);
nor U13722 (N_13722,N_13459,N_13440);
nand U13723 (N_13723,N_13487,N_13405);
nor U13724 (N_13724,N_13429,N_13400);
xor U13725 (N_13725,N_13406,N_13262);
xnor U13726 (N_13726,N_13322,N_13264);
nor U13727 (N_13727,N_13259,N_13334);
and U13728 (N_13728,N_13456,N_13389);
nor U13729 (N_13729,N_13431,N_13306);
xnor U13730 (N_13730,N_13430,N_13313);
nand U13731 (N_13731,N_13390,N_13421);
nand U13732 (N_13732,N_13350,N_13363);
nor U13733 (N_13733,N_13283,N_13259);
xnor U13734 (N_13734,N_13260,N_13451);
and U13735 (N_13735,N_13256,N_13327);
xnor U13736 (N_13736,N_13422,N_13329);
or U13737 (N_13737,N_13299,N_13441);
nor U13738 (N_13738,N_13311,N_13414);
xnor U13739 (N_13739,N_13403,N_13449);
nor U13740 (N_13740,N_13493,N_13250);
and U13741 (N_13741,N_13324,N_13476);
nor U13742 (N_13742,N_13405,N_13371);
nand U13743 (N_13743,N_13322,N_13276);
xor U13744 (N_13744,N_13429,N_13468);
xor U13745 (N_13745,N_13374,N_13402);
nand U13746 (N_13746,N_13467,N_13414);
nand U13747 (N_13747,N_13250,N_13463);
or U13748 (N_13748,N_13489,N_13475);
and U13749 (N_13749,N_13356,N_13280);
xnor U13750 (N_13750,N_13681,N_13583);
nand U13751 (N_13751,N_13646,N_13525);
nor U13752 (N_13752,N_13708,N_13587);
or U13753 (N_13753,N_13581,N_13580);
and U13754 (N_13754,N_13604,N_13704);
nor U13755 (N_13755,N_13615,N_13546);
nor U13756 (N_13756,N_13743,N_13624);
nand U13757 (N_13757,N_13632,N_13638);
xnor U13758 (N_13758,N_13713,N_13671);
xor U13759 (N_13759,N_13666,N_13723);
xnor U13760 (N_13760,N_13711,N_13538);
or U13761 (N_13761,N_13608,N_13503);
nand U13762 (N_13762,N_13688,N_13532);
and U13763 (N_13763,N_13717,N_13504);
nand U13764 (N_13764,N_13636,N_13652);
and U13765 (N_13765,N_13617,N_13545);
and U13766 (N_13766,N_13619,N_13517);
nor U13767 (N_13767,N_13676,N_13630);
or U13768 (N_13768,N_13643,N_13515);
xnor U13769 (N_13769,N_13639,N_13668);
or U13770 (N_13770,N_13728,N_13659);
or U13771 (N_13771,N_13578,N_13635);
and U13772 (N_13772,N_13718,N_13523);
nand U13773 (N_13773,N_13586,N_13606);
and U13774 (N_13774,N_13582,N_13536);
nand U13775 (N_13775,N_13575,N_13698);
or U13776 (N_13776,N_13500,N_13597);
and U13777 (N_13777,N_13518,N_13591);
nand U13778 (N_13778,N_13506,N_13610);
or U13779 (N_13779,N_13732,N_13640);
nor U13780 (N_13780,N_13634,N_13522);
and U13781 (N_13781,N_13707,N_13651);
xnor U13782 (N_13782,N_13528,N_13574);
or U13783 (N_13783,N_13527,N_13649);
xor U13784 (N_13784,N_13677,N_13702);
and U13785 (N_13785,N_13692,N_13740);
nand U13786 (N_13786,N_13594,N_13524);
nor U13787 (N_13787,N_13621,N_13508);
nand U13788 (N_13788,N_13648,N_13622);
nor U13789 (N_13789,N_13730,N_13516);
nor U13790 (N_13790,N_13706,N_13641);
and U13791 (N_13791,N_13678,N_13629);
nor U13792 (N_13792,N_13540,N_13694);
xor U13793 (N_13793,N_13560,N_13710);
or U13794 (N_13794,N_13609,N_13746);
xnor U13795 (N_13795,N_13612,N_13563);
and U13796 (N_13796,N_13644,N_13513);
xor U13797 (N_13797,N_13512,N_13555);
nor U13798 (N_13798,N_13533,N_13502);
or U13799 (N_13799,N_13534,N_13670);
or U13800 (N_13800,N_13565,N_13703);
nand U13801 (N_13801,N_13655,N_13675);
nand U13802 (N_13802,N_13544,N_13589);
and U13803 (N_13803,N_13726,N_13637);
xnor U13804 (N_13804,N_13673,N_13566);
nor U13805 (N_13805,N_13745,N_13600);
or U13806 (N_13806,N_13735,N_13664);
nor U13807 (N_13807,N_13531,N_13562);
xnor U13808 (N_13808,N_13611,N_13737);
xor U13809 (N_13809,N_13665,N_13537);
or U13810 (N_13810,N_13656,N_13557);
or U13811 (N_13811,N_13584,N_13722);
xor U13812 (N_13812,N_13667,N_13747);
and U13813 (N_13813,N_13660,N_13716);
nor U13814 (N_13814,N_13691,N_13559);
xor U13815 (N_13815,N_13653,N_13719);
xor U13816 (N_13816,N_13645,N_13507);
or U13817 (N_13817,N_13585,N_13521);
or U13818 (N_13818,N_13509,N_13680);
nand U13819 (N_13819,N_13647,N_13614);
and U13820 (N_13820,N_13542,N_13590);
nand U13821 (N_13821,N_13564,N_13588);
and U13822 (N_13822,N_13547,N_13535);
nor U13823 (N_13823,N_13724,N_13572);
and U13824 (N_13824,N_13720,N_13685);
and U13825 (N_13825,N_13567,N_13623);
nor U13826 (N_13826,N_13598,N_13744);
nand U13827 (N_13827,N_13618,N_13697);
and U13828 (N_13828,N_13558,N_13616);
and U13829 (N_13829,N_13749,N_13510);
nand U13830 (N_13830,N_13715,N_13501);
or U13831 (N_13831,N_13712,N_13550);
xnor U13832 (N_13832,N_13738,N_13593);
and U13833 (N_13833,N_13709,N_13576);
or U13834 (N_13834,N_13548,N_13739);
nand U13835 (N_13835,N_13736,N_13520);
xor U13836 (N_13836,N_13631,N_13734);
and U13837 (N_13837,N_13721,N_13689);
xnor U13838 (N_13838,N_13539,N_13603);
nand U13839 (N_13839,N_13733,N_13573);
and U13840 (N_13840,N_13505,N_13633);
or U13841 (N_13841,N_13687,N_13627);
xor U13842 (N_13842,N_13686,N_13601);
xnor U13843 (N_13843,N_13568,N_13551);
nor U13844 (N_13844,N_13553,N_13561);
xor U13845 (N_13845,N_13571,N_13674);
or U13846 (N_13846,N_13662,N_13741);
or U13847 (N_13847,N_13620,N_13683);
or U13848 (N_13848,N_13569,N_13654);
and U13849 (N_13849,N_13657,N_13663);
xor U13850 (N_13850,N_13595,N_13599);
nand U13851 (N_13851,N_13714,N_13699);
and U13852 (N_13852,N_13700,N_13695);
and U13853 (N_13853,N_13530,N_13748);
nand U13854 (N_13854,N_13725,N_13592);
and U13855 (N_13855,N_13696,N_13549);
and U13856 (N_13856,N_13658,N_13672);
nor U13857 (N_13857,N_13669,N_13742);
nand U13858 (N_13858,N_13519,N_13727);
nand U13859 (N_13859,N_13705,N_13529);
nor U13860 (N_13860,N_13729,N_13554);
or U13861 (N_13861,N_13605,N_13693);
or U13862 (N_13862,N_13684,N_13570);
nor U13863 (N_13863,N_13625,N_13690);
or U13864 (N_13864,N_13661,N_13731);
nor U13865 (N_13865,N_13613,N_13577);
and U13866 (N_13866,N_13541,N_13526);
nor U13867 (N_13867,N_13511,N_13596);
and U13868 (N_13868,N_13682,N_13628);
or U13869 (N_13869,N_13626,N_13556);
and U13870 (N_13870,N_13701,N_13543);
and U13871 (N_13871,N_13552,N_13607);
and U13872 (N_13872,N_13514,N_13642);
and U13873 (N_13873,N_13602,N_13650);
xnor U13874 (N_13874,N_13679,N_13579);
nor U13875 (N_13875,N_13566,N_13618);
xor U13876 (N_13876,N_13701,N_13557);
nor U13877 (N_13877,N_13692,N_13733);
or U13878 (N_13878,N_13626,N_13661);
or U13879 (N_13879,N_13675,N_13561);
or U13880 (N_13880,N_13633,N_13638);
nor U13881 (N_13881,N_13658,N_13630);
nor U13882 (N_13882,N_13699,N_13648);
and U13883 (N_13883,N_13716,N_13691);
and U13884 (N_13884,N_13736,N_13557);
xor U13885 (N_13885,N_13747,N_13507);
and U13886 (N_13886,N_13568,N_13668);
or U13887 (N_13887,N_13566,N_13569);
and U13888 (N_13888,N_13682,N_13585);
nand U13889 (N_13889,N_13706,N_13581);
xnor U13890 (N_13890,N_13526,N_13679);
xor U13891 (N_13891,N_13575,N_13649);
nand U13892 (N_13892,N_13560,N_13739);
or U13893 (N_13893,N_13569,N_13642);
or U13894 (N_13894,N_13533,N_13532);
and U13895 (N_13895,N_13612,N_13701);
and U13896 (N_13896,N_13711,N_13615);
or U13897 (N_13897,N_13672,N_13544);
and U13898 (N_13898,N_13590,N_13529);
and U13899 (N_13899,N_13544,N_13636);
nand U13900 (N_13900,N_13628,N_13687);
and U13901 (N_13901,N_13642,N_13700);
nand U13902 (N_13902,N_13571,N_13726);
nand U13903 (N_13903,N_13610,N_13545);
and U13904 (N_13904,N_13721,N_13594);
and U13905 (N_13905,N_13730,N_13623);
nor U13906 (N_13906,N_13731,N_13617);
nor U13907 (N_13907,N_13522,N_13576);
or U13908 (N_13908,N_13715,N_13716);
nor U13909 (N_13909,N_13744,N_13740);
nand U13910 (N_13910,N_13643,N_13605);
nand U13911 (N_13911,N_13519,N_13673);
and U13912 (N_13912,N_13660,N_13556);
xor U13913 (N_13913,N_13655,N_13526);
nand U13914 (N_13914,N_13558,N_13706);
or U13915 (N_13915,N_13521,N_13692);
xor U13916 (N_13916,N_13736,N_13535);
nor U13917 (N_13917,N_13701,N_13629);
xnor U13918 (N_13918,N_13513,N_13503);
nand U13919 (N_13919,N_13613,N_13703);
nand U13920 (N_13920,N_13613,N_13561);
nand U13921 (N_13921,N_13686,N_13539);
or U13922 (N_13922,N_13646,N_13726);
xnor U13923 (N_13923,N_13650,N_13697);
or U13924 (N_13924,N_13627,N_13673);
nand U13925 (N_13925,N_13544,N_13548);
nand U13926 (N_13926,N_13588,N_13696);
and U13927 (N_13927,N_13519,N_13706);
or U13928 (N_13928,N_13650,N_13739);
and U13929 (N_13929,N_13738,N_13511);
and U13930 (N_13930,N_13658,N_13629);
nand U13931 (N_13931,N_13667,N_13679);
or U13932 (N_13932,N_13635,N_13515);
nor U13933 (N_13933,N_13695,N_13696);
nand U13934 (N_13934,N_13720,N_13658);
xnor U13935 (N_13935,N_13712,N_13710);
xor U13936 (N_13936,N_13630,N_13616);
and U13937 (N_13937,N_13506,N_13566);
xnor U13938 (N_13938,N_13562,N_13609);
xor U13939 (N_13939,N_13699,N_13539);
nand U13940 (N_13940,N_13611,N_13580);
or U13941 (N_13941,N_13719,N_13623);
nand U13942 (N_13942,N_13668,N_13501);
xnor U13943 (N_13943,N_13717,N_13613);
xor U13944 (N_13944,N_13547,N_13640);
nand U13945 (N_13945,N_13576,N_13703);
nand U13946 (N_13946,N_13741,N_13678);
nand U13947 (N_13947,N_13536,N_13580);
xor U13948 (N_13948,N_13676,N_13703);
or U13949 (N_13949,N_13682,N_13503);
xnor U13950 (N_13950,N_13708,N_13696);
xor U13951 (N_13951,N_13663,N_13523);
or U13952 (N_13952,N_13542,N_13581);
or U13953 (N_13953,N_13723,N_13592);
or U13954 (N_13954,N_13663,N_13679);
and U13955 (N_13955,N_13722,N_13681);
or U13956 (N_13956,N_13571,N_13692);
or U13957 (N_13957,N_13691,N_13625);
nand U13958 (N_13958,N_13725,N_13580);
and U13959 (N_13959,N_13742,N_13576);
nand U13960 (N_13960,N_13517,N_13568);
and U13961 (N_13961,N_13737,N_13572);
and U13962 (N_13962,N_13586,N_13696);
nand U13963 (N_13963,N_13662,N_13695);
nand U13964 (N_13964,N_13587,N_13596);
nand U13965 (N_13965,N_13707,N_13704);
and U13966 (N_13966,N_13543,N_13554);
xnor U13967 (N_13967,N_13659,N_13693);
nand U13968 (N_13968,N_13596,N_13684);
xnor U13969 (N_13969,N_13543,N_13574);
nand U13970 (N_13970,N_13529,N_13691);
or U13971 (N_13971,N_13573,N_13664);
and U13972 (N_13972,N_13674,N_13743);
nand U13973 (N_13973,N_13556,N_13649);
nand U13974 (N_13974,N_13743,N_13558);
or U13975 (N_13975,N_13625,N_13603);
and U13976 (N_13976,N_13661,N_13614);
or U13977 (N_13977,N_13688,N_13540);
nor U13978 (N_13978,N_13728,N_13671);
or U13979 (N_13979,N_13545,N_13719);
xor U13980 (N_13980,N_13526,N_13613);
nor U13981 (N_13981,N_13655,N_13640);
nor U13982 (N_13982,N_13637,N_13672);
or U13983 (N_13983,N_13524,N_13592);
nor U13984 (N_13984,N_13663,N_13629);
xor U13985 (N_13985,N_13605,N_13745);
and U13986 (N_13986,N_13619,N_13578);
nand U13987 (N_13987,N_13641,N_13749);
or U13988 (N_13988,N_13506,N_13501);
and U13989 (N_13989,N_13676,N_13585);
or U13990 (N_13990,N_13614,N_13672);
nand U13991 (N_13991,N_13611,N_13712);
xnor U13992 (N_13992,N_13696,N_13516);
xnor U13993 (N_13993,N_13654,N_13638);
nand U13994 (N_13994,N_13657,N_13578);
nand U13995 (N_13995,N_13670,N_13526);
and U13996 (N_13996,N_13578,N_13666);
nor U13997 (N_13997,N_13597,N_13575);
and U13998 (N_13998,N_13613,N_13744);
xnor U13999 (N_13999,N_13651,N_13613);
xor U14000 (N_14000,N_13762,N_13979);
and U14001 (N_14001,N_13750,N_13909);
and U14002 (N_14002,N_13873,N_13930);
xor U14003 (N_14003,N_13799,N_13779);
or U14004 (N_14004,N_13995,N_13915);
xnor U14005 (N_14005,N_13870,N_13954);
and U14006 (N_14006,N_13842,N_13807);
or U14007 (N_14007,N_13927,N_13957);
nand U14008 (N_14008,N_13893,N_13876);
or U14009 (N_14009,N_13879,N_13908);
nor U14010 (N_14010,N_13999,N_13896);
nand U14011 (N_14011,N_13880,N_13850);
nor U14012 (N_14012,N_13751,N_13910);
and U14013 (N_14013,N_13785,N_13943);
xnor U14014 (N_14014,N_13795,N_13867);
or U14015 (N_14015,N_13757,N_13839);
nand U14016 (N_14016,N_13851,N_13941);
xor U14017 (N_14017,N_13970,N_13761);
xnor U14018 (N_14018,N_13900,N_13776);
and U14019 (N_14019,N_13860,N_13773);
nand U14020 (N_14020,N_13960,N_13774);
xor U14021 (N_14021,N_13986,N_13819);
nand U14022 (N_14022,N_13874,N_13760);
nor U14023 (N_14023,N_13801,N_13853);
nor U14024 (N_14024,N_13814,N_13822);
and U14025 (N_14025,N_13857,N_13899);
nor U14026 (N_14026,N_13856,N_13935);
xor U14027 (N_14027,N_13996,N_13987);
or U14028 (N_14028,N_13976,N_13800);
nor U14029 (N_14029,N_13961,N_13753);
nand U14030 (N_14030,N_13913,N_13938);
xnor U14031 (N_14031,N_13926,N_13984);
nand U14032 (N_14032,N_13902,N_13813);
nand U14033 (N_14033,N_13828,N_13759);
or U14034 (N_14034,N_13988,N_13796);
and U14035 (N_14035,N_13791,N_13824);
nand U14036 (N_14036,N_13977,N_13848);
and U14037 (N_14037,N_13883,N_13797);
and U14038 (N_14038,N_13964,N_13858);
xor U14039 (N_14039,N_13990,N_13821);
xor U14040 (N_14040,N_13985,N_13997);
nor U14041 (N_14041,N_13998,N_13865);
or U14042 (N_14042,N_13780,N_13837);
nand U14043 (N_14043,N_13875,N_13942);
or U14044 (N_14044,N_13830,N_13871);
and U14045 (N_14045,N_13792,N_13968);
nor U14046 (N_14046,N_13869,N_13916);
nand U14047 (N_14047,N_13804,N_13825);
xor U14048 (N_14048,N_13812,N_13790);
nor U14049 (N_14049,N_13993,N_13891);
nand U14050 (N_14050,N_13950,N_13854);
nand U14051 (N_14051,N_13934,N_13794);
nor U14052 (N_14052,N_13881,N_13843);
nand U14053 (N_14053,N_13864,N_13810);
nand U14054 (N_14054,N_13921,N_13754);
nand U14055 (N_14055,N_13962,N_13931);
xor U14056 (N_14056,N_13763,N_13906);
nor U14057 (N_14057,N_13835,N_13928);
or U14058 (N_14058,N_13823,N_13920);
nor U14059 (N_14059,N_13786,N_13844);
or U14060 (N_14060,N_13862,N_13783);
and U14061 (N_14061,N_13980,N_13940);
or U14062 (N_14062,N_13758,N_13831);
nor U14063 (N_14063,N_13885,N_13772);
nand U14064 (N_14064,N_13919,N_13861);
or U14065 (N_14065,N_13882,N_13847);
or U14066 (N_14066,N_13923,N_13973);
nor U14067 (N_14067,N_13949,N_13784);
nor U14068 (N_14068,N_13904,N_13992);
or U14069 (N_14069,N_13782,N_13922);
or U14070 (N_14070,N_13884,N_13767);
and U14071 (N_14071,N_13789,N_13894);
or U14072 (N_14072,N_13946,N_13981);
or U14073 (N_14073,N_13781,N_13868);
nand U14074 (N_14074,N_13877,N_13951);
and U14075 (N_14075,N_13972,N_13755);
nand U14076 (N_14076,N_13820,N_13852);
xnor U14077 (N_14077,N_13945,N_13966);
nand U14078 (N_14078,N_13897,N_13971);
or U14079 (N_14079,N_13793,N_13826);
or U14080 (N_14080,N_13939,N_13777);
and U14081 (N_14081,N_13770,N_13937);
nor U14082 (N_14082,N_13863,N_13788);
or U14083 (N_14083,N_13752,N_13849);
xnor U14084 (N_14084,N_13907,N_13989);
or U14085 (N_14085,N_13798,N_13969);
nand U14086 (N_14086,N_13771,N_13959);
nor U14087 (N_14087,N_13994,N_13914);
nor U14088 (N_14088,N_13889,N_13769);
nor U14089 (N_14089,N_13803,N_13905);
or U14090 (N_14090,N_13855,N_13808);
nor U14091 (N_14091,N_13809,N_13833);
xnor U14092 (N_14092,N_13918,N_13829);
nor U14093 (N_14093,N_13963,N_13787);
nand U14094 (N_14094,N_13958,N_13802);
or U14095 (N_14095,N_13840,N_13911);
nor U14096 (N_14096,N_13948,N_13947);
nor U14097 (N_14097,N_13929,N_13924);
nand U14098 (N_14098,N_13982,N_13838);
nor U14099 (N_14099,N_13917,N_13890);
or U14100 (N_14100,N_13815,N_13983);
nand U14101 (N_14101,N_13903,N_13932);
or U14102 (N_14102,N_13841,N_13859);
nand U14103 (N_14103,N_13836,N_13978);
and U14104 (N_14104,N_13944,N_13912);
and U14105 (N_14105,N_13925,N_13965);
or U14106 (N_14106,N_13975,N_13974);
nand U14107 (N_14107,N_13895,N_13845);
nand U14108 (N_14108,N_13887,N_13878);
and U14109 (N_14109,N_13811,N_13953);
nand U14110 (N_14110,N_13886,N_13775);
xor U14111 (N_14111,N_13765,N_13768);
xor U14112 (N_14112,N_13888,N_13832);
or U14113 (N_14113,N_13756,N_13817);
and U14114 (N_14114,N_13952,N_13955);
nand U14115 (N_14115,N_13805,N_13834);
nand U14116 (N_14116,N_13778,N_13967);
nor U14117 (N_14117,N_13991,N_13764);
nor U14118 (N_14118,N_13933,N_13827);
or U14119 (N_14119,N_13956,N_13898);
nand U14120 (N_14120,N_13816,N_13766);
and U14121 (N_14121,N_13818,N_13806);
and U14122 (N_14122,N_13892,N_13866);
nor U14123 (N_14123,N_13872,N_13901);
or U14124 (N_14124,N_13846,N_13936);
nor U14125 (N_14125,N_13996,N_13809);
nand U14126 (N_14126,N_13947,N_13858);
and U14127 (N_14127,N_13952,N_13798);
or U14128 (N_14128,N_13771,N_13987);
or U14129 (N_14129,N_13910,N_13860);
nand U14130 (N_14130,N_13926,N_13998);
nor U14131 (N_14131,N_13921,N_13903);
nor U14132 (N_14132,N_13907,N_13797);
xor U14133 (N_14133,N_13820,N_13985);
nand U14134 (N_14134,N_13808,N_13879);
xnor U14135 (N_14135,N_13795,N_13980);
and U14136 (N_14136,N_13935,N_13823);
nor U14137 (N_14137,N_13794,N_13942);
and U14138 (N_14138,N_13847,N_13918);
xor U14139 (N_14139,N_13752,N_13806);
xnor U14140 (N_14140,N_13895,N_13966);
nand U14141 (N_14141,N_13989,N_13958);
xnor U14142 (N_14142,N_13799,N_13843);
nor U14143 (N_14143,N_13804,N_13940);
or U14144 (N_14144,N_13968,N_13858);
nand U14145 (N_14145,N_13977,N_13987);
nor U14146 (N_14146,N_13878,N_13870);
xnor U14147 (N_14147,N_13811,N_13835);
nand U14148 (N_14148,N_13875,N_13816);
or U14149 (N_14149,N_13942,N_13815);
xor U14150 (N_14150,N_13853,N_13816);
nand U14151 (N_14151,N_13888,N_13937);
xor U14152 (N_14152,N_13830,N_13821);
xor U14153 (N_14153,N_13787,N_13971);
xnor U14154 (N_14154,N_13906,N_13967);
nor U14155 (N_14155,N_13773,N_13913);
or U14156 (N_14156,N_13919,N_13822);
nor U14157 (N_14157,N_13924,N_13905);
xnor U14158 (N_14158,N_13956,N_13825);
nand U14159 (N_14159,N_13834,N_13882);
xor U14160 (N_14160,N_13927,N_13844);
nor U14161 (N_14161,N_13819,N_13800);
and U14162 (N_14162,N_13848,N_13800);
and U14163 (N_14163,N_13795,N_13876);
nand U14164 (N_14164,N_13891,N_13856);
nor U14165 (N_14165,N_13757,N_13907);
or U14166 (N_14166,N_13951,N_13937);
and U14167 (N_14167,N_13780,N_13890);
nand U14168 (N_14168,N_13795,N_13919);
xnor U14169 (N_14169,N_13785,N_13930);
and U14170 (N_14170,N_13798,N_13850);
or U14171 (N_14171,N_13798,N_13770);
and U14172 (N_14172,N_13849,N_13850);
and U14173 (N_14173,N_13978,N_13917);
xor U14174 (N_14174,N_13887,N_13795);
nand U14175 (N_14175,N_13997,N_13795);
nand U14176 (N_14176,N_13962,N_13943);
and U14177 (N_14177,N_13983,N_13833);
nand U14178 (N_14178,N_13752,N_13943);
nor U14179 (N_14179,N_13934,N_13755);
xnor U14180 (N_14180,N_13751,N_13786);
xnor U14181 (N_14181,N_13861,N_13793);
nand U14182 (N_14182,N_13922,N_13989);
and U14183 (N_14183,N_13886,N_13758);
nor U14184 (N_14184,N_13896,N_13810);
and U14185 (N_14185,N_13808,N_13775);
and U14186 (N_14186,N_13796,N_13888);
xnor U14187 (N_14187,N_13807,N_13759);
and U14188 (N_14188,N_13930,N_13755);
xor U14189 (N_14189,N_13976,N_13776);
xnor U14190 (N_14190,N_13832,N_13775);
xor U14191 (N_14191,N_13887,N_13836);
or U14192 (N_14192,N_13758,N_13759);
or U14193 (N_14193,N_13960,N_13898);
and U14194 (N_14194,N_13844,N_13876);
nor U14195 (N_14195,N_13860,N_13987);
and U14196 (N_14196,N_13898,N_13995);
and U14197 (N_14197,N_13872,N_13966);
or U14198 (N_14198,N_13788,N_13760);
and U14199 (N_14199,N_13997,N_13930);
nand U14200 (N_14200,N_13914,N_13999);
nand U14201 (N_14201,N_13777,N_13988);
and U14202 (N_14202,N_13809,N_13842);
and U14203 (N_14203,N_13810,N_13867);
and U14204 (N_14204,N_13861,N_13959);
xnor U14205 (N_14205,N_13838,N_13880);
and U14206 (N_14206,N_13831,N_13950);
and U14207 (N_14207,N_13893,N_13868);
xnor U14208 (N_14208,N_13958,N_13967);
and U14209 (N_14209,N_13882,N_13777);
xnor U14210 (N_14210,N_13780,N_13970);
or U14211 (N_14211,N_13892,N_13834);
or U14212 (N_14212,N_13800,N_13809);
or U14213 (N_14213,N_13950,N_13862);
and U14214 (N_14214,N_13832,N_13874);
xor U14215 (N_14215,N_13949,N_13851);
xor U14216 (N_14216,N_13798,N_13822);
and U14217 (N_14217,N_13925,N_13831);
nor U14218 (N_14218,N_13888,N_13755);
xor U14219 (N_14219,N_13996,N_13759);
and U14220 (N_14220,N_13864,N_13858);
nand U14221 (N_14221,N_13915,N_13835);
and U14222 (N_14222,N_13769,N_13942);
and U14223 (N_14223,N_13810,N_13955);
nor U14224 (N_14224,N_13842,N_13760);
nand U14225 (N_14225,N_13994,N_13924);
and U14226 (N_14226,N_13824,N_13987);
or U14227 (N_14227,N_13924,N_13920);
nor U14228 (N_14228,N_13827,N_13865);
nand U14229 (N_14229,N_13803,N_13965);
or U14230 (N_14230,N_13882,N_13898);
nor U14231 (N_14231,N_13867,N_13964);
nor U14232 (N_14232,N_13884,N_13855);
and U14233 (N_14233,N_13824,N_13887);
and U14234 (N_14234,N_13833,N_13905);
xnor U14235 (N_14235,N_13997,N_13855);
and U14236 (N_14236,N_13901,N_13782);
xor U14237 (N_14237,N_13873,N_13874);
or U14238 (N_14238,N_13964,N_13869);
nand U14239 (N_14239,N_13782,N_13882);
or U14240 (N_14240,N_13782,N_13987);
nor U14241 (N_14241,N_13977,N_13899);
xor U14242 (N_14242,N_13777,N_13975);
or U14243 (N_14243,N_13826,N_13798);
or U14244 (N_14244,N_13946,N_13834);
nand U14245 (N_14245,N_13769,N_13888);
xnor U14246 (N_14246,N_13776,N_13946);
nand U14247 (N_14247,N_13996,N_13917);
or U14248 (N_14248,N_13750,N_13914);
or U14249 (N_14249,N_13863,N_13923);
xor U14250 (N_14250,N_14013,N_14137);
or U14251 (N_14251,N_14048,N_14159);
nand U14252 (N_14252,N_14024,N_14235);
and U14253 (N_14253,N_14094,N_14089);
and U14254 (N_14254,N_14043,N_14128);
and U14255 (N_14255,N_14219,N_14054);
nor U14256 (N_14256,N_14151,N_14226);
nor U14257 (N_14257,N_14100,N_14126);
and U14258 (N_14258,N_14225,N_14115);
nor U14259 (N_14259,N_14059,N_14158);
nand U14260 (N_14260,N_14178,N_14180);
nor U14261 (N_14261,N_14026,N_14058);
and U14262 (N_14262,N_14139,N_14217);
or U14263 (N_14263,N_14032,N_14082);
nand U14264 (N_14264,N_14042,N_14134);
or U14265 (N_14265,N_14101,N_14138);
nand U14266 (N_14266,N_14243,N_14209);
nand U14267 (N_14267,N_14006,N_14199);
and U14268 (N_14268,N_14197,N_14182);
xor U14269 (N_14269,N_14087,N_14008);
and U14270 (N_14270,N_14183,N_14073);
nor U14271 (N_14271,N_14143,N_14040);
xor U14272 (N_14272,N_14107,N_14000);
nand U14273 (N_14273,N_14039,N_14105);
or U14274 (N_14274,N_14085,N_14062);
nand U14275 (N_14275,N_14057,N_14152);
nand U14276 (N_14276,N_14228,N_14181);
xnor U14277 (N_14277,N_14116,N_14187);
xor U14278 (N_14278,N_14127,N_14122);
and U14279 (N_14279,N_14200,N_14034);
and U14280 (N_14280,N_14002,N_14078);
or U14281 (N_14281,N_14051,N_14175);
nand U14282 (N_14282,N_14046,N_14163);
nor U14283 (N_14283,N_14037,N_14146);
nor U14284 (N_14284,N_14130,N_14076);
nor U14285 (N_14285,N_14123,N_14055);
xor U14286 (N_14286,N_14171,N_14003);
xor U14287 (N_14287,N_14067,N_14213);
nand U14288 (N_14288,N_14030,N_14153);
xor U14289 (N_14289,N_14022,N_14244);
or U14290 (N_14290,N_14246,N_14157);
xor U14291 (N_14291,N_14207,N_14021);
and U14292 (N_14292,N_14227,N_14242);
or U14293 (N_14293,N_14079,N_14038);
nor U14294 (N_14294,N_14001,N_14149);
nor U14295 (N_14295,N_14113,N_14096);
nand U14296 (N_14296,N_14190,N_14177);
nand U14297 (N_14297,N_14035,N_14241);
nand U14298 (N_14298,N_14156,N_14004);
nand U14299 (N_14299,N_14248,N_14208);
or U14300 (N_14300,N_14086,N_14015);
or U14301 (N_14301,N_14170,N_14184);
nand U14302 (N_14302,N_14202,N_14220);
and U14303 (N_14303,N_14192,N_14154);
and U14304 (N_14304,N_14012,N_14135);
nand U14305 (N_14305,N_14230,N_14216);
nor U14306 (N_14306,N_14141,N_14104);
nor U14307 (N_14307,N_14052,N_14028);
or U14308 (N_14308,N_14131,N_14237);
xnor U14309 (N_14309,N_14047,N_14169);
or U14310 (N_14310,N_14165,N_14041);
and U14311 (N_14311,N_14162,N_14231);
or U14312 (N_14312,N_14009,N_14196);
nand U14313 (N_14313,N_14064,N_14091);
nand U14314 (N_14314,N_14108,N_14161);
and U14315 (N_14315,N_14110,N_14103);
nand U14316 (N_14316,N_14083,N_14011);
xor U14317 (N_14317,N_14172,N_14117);
nor U14318 (N_14318,N_14176,N_14097);
and U14319 (N_14319,N_14164,N_14204);
and U14320 (N_14320,N_14186,N_14068);
or U14321 (N_14321,N_14224,N_14179);
nand U14322 (N_14322,N_14088,N_14027);
xor U14323 (N_14323,N_14155,N_14121);
nor U14324 (N_14324,N_14095,N_14045);
nand U14325 (N_14325,N_14142,N_14066);
nor U14326 (N_14326,N_14185,N_14140);
or U14327 (N_14327,N_14191,N_14081);
nor U14328 (N_14328,N_14124,N_14023);
or U14329 (N_14329,N_14007,N_14238);
nand U14330 (N_14330,N_14071,N_14069);
nand U14331 (N_14331,N_14020,N_14150);
xor U14332 (N_14332,N_14025,N_14070);
xor U14333 (N_14333,N_14029,N_14019);
xor U14334 (N_14334,N_14173,N_14240);
nor U14335 (N_14335,N_14111,N_14132);
xor U14336 (N_14336,N_14206,N_14188);
or U14337 (N_14337,N_14072,N_14063);
or U14338 (N_14338,N_14160,N_14245);
or U14339 (N_14339,N_14093,N_14198);
and U14340 (N_14340,N_14234,N_14056);
xnor U14341 (N_14341,N_14017,N_14201);
and U14342 (N_14342,N_14044,N_14074);
and U14343 (N_14343,N_14147,N_14120);
or U14344 (N_14344,N_14014,N_14174);
or U14345 (N_14345,N_14053,N_14144);
xor U14346 (N_14346,N_14148,N_14136);
xnor U14347 (N_14347,N_14080,N_14212);
nand U14348 (N_14348,N_14221,N_14211);
nand U14349 (N_14349,N_14218,N_14061);
or U14350 (N_14350,N_14214,N_14102);
nand U14351 (N_14351,N_14249,N_14106);
and U14352 (N_14352,N_14223,N_14075);
nand U14353 (N_14353,N_14077,N_14114);
and U14354 (N_14354,N_14125,N_14166);
nand U14355 (N_14355,N_14215,N_14205);
and U14356 (N_14356,N_14049,N_14084);
and U14357 (N_14357,N_14112,N_14232);
and U14358 (N_14358,N_14189,N_14118);
and U14359 (N_14359,N_14133,N_14129);
nand U14360 (N_14360,N_14098,N_14060);
and U14361 (N_14361,N_14233,N_14247);
nand U14362 (N_14362,N_14167,N_14168);
nor U14363 (N_14363,N_14195,N_14018);
nand U14364 (N_14364,N_14092,N_14010);
nor U14365 (N_14365,N_14031,N_14222);
nor U14366 (N_14366,N_14090,N_14193);
and U14367 (N_14367,N_14239,N_14210);
xor U14368 (N_14368,N_14005,N_14236);
nor U14369 (N_14369,N_14145,N_14229);
and U14370 (N_14370,N_14099,N_14119);
xnor U14371 (N_14371,N_14203,N_14036);
nor U14372 (N_14372,N_14109,N_14016);
and U14373 (N_14373,N_14065,N_14050);
nor U14374 (N_14374,N_14194,N_14033);
or U14375 (N_14375,N_14028,N_14212);
nand U14376 (N_14376,N_14029,N_14204);
nand U14377 (N_14377,N_14034,N_14019);
xor U14378 (N_14378,N_14151,N_14213);
nand U14379 (N_14379,N_14207,N_14141);
or U14380 (N_14380,N_14137,N_14135);
nor U14381 (N_14381,N_14239,N_14121);
nand U14382 (N_14382,N_14033,N_14148);
and U14383 (N_14383,N_14096,N_14115);
nor U14384 (N_14384,N_14175,N_14161);
nor U14385 (N_14385,N_14030,N_14063);
nor U14386 (N_14386,N_14004,N_14211);
xor U14387 (N_14387,N_14196,N_14118);
xnor U14388 (N_14388,N_14151,N_14205);
nor U14389 (N_14389,N_14223,N_14090);
nand U14390 (N_14390,N_14204,N_14044);
nand U14391 (N_14391,N_14249,N_14059);
nand U14392 (N_14392,N_14242,N_14070);
nand U14393 (N_14393,N_14069,N_14168);
xnor U14394 (N_14394,N_14157,N_14046);
or U14395 (N_14395,N_14046,N_14082);
nor U14396 (N_14396,N_14150,N_14138);
xor U14397 (N_14397,N_14244,N_14217);
and U14398 (N_14398,N_14112,N_14107);
nor U14399 (N_14399,N_14186,N_14154);
or U14400 (N_14400,N_14041,N_14040);
xnor U14401 (N_14401,N_14156,N_14015);
xnor U14402 (N_14402,N_14209,N_14027);
xnor U14403 (N_14403,N_14189,N_14143);
xnor U14404 (N_14404,N_14018,N_14097);
xnor U14405 (N_14405,N_14038,N_14159);
and U14406 (N_14406,N_14031,N_14160);
and U14407 (N_14407,N_14090,N_14008);
or U14408 (N_14408,N_14122,N_14220);
nor U14409 (N_14409,N_14003,N_14230);
and U14410 (N_14410,N_14238,N_14139);
and U14411 (N_14411,N_14051,N_14160);
xor U14412 (N_14412,N_14148,N_14124);
nand U14413 (N_14413,N_14190,N_14026);
nand U14414 (N_14414,N_14034,N_14004);
and U14415 (N_14415,N_14205,N_14048);
and U14416 (N_14416,N_14110,N_14125);
xor U14417 (N_14417,N_14200,N_14201);
or U14418 (N_14418,N_14032,N_14138);
and U14419 (N_14419,N_14209,N_14062);
xnor U14420 (N_14420,N_14082,N_14231);
xnor U14421 (N_14421,N_14116,N_14022);
and U14422 (N_14422,N_14249,N_14081);
nor U14423 (N_14423,N_14045,N_14177);
and U14424 (N_14424,N_14061,N_14119);
or U14425 (N_14425,N_14224,N_14154);
or U14426 (N_14426,N_14203,N_14148);
and U14427 (N_14427,N_14046,N_14077);
xnor U14428 (N_14428,N_14197,N_14232);
or U14429 (N_14429,N_14154,N_14094);
and U14430 (N_14430,N_14144,N_14048);
and U14431 (N_14431,N_14003,N_14145);
and U14432 (N_14432,N_14044,N_14139);
and U14433 (N_14433,N_14091,N_14150);
nand U14434 (N_14434,N_14087,N_14184);
xnor U14435 (N_14435,N_14059,N_14030);
nor U14436 (N_14436,N_14207,N_14070);
and U14437 (N_14437,N_14198,N_14011);
or U14438 (N_14438,N_14069,N_14246);
or U14439 (N_14439,N_14102,N_14049);
or U14440 (N_14440,N_14101,N_14133);
nand U14441 (N_14441,N_14244,N_14034);
xor U14442 (N_14442,N_14237,N_14113);
nand U14443 (N_14443,N_14125,N_14231);
xnor U14444 (N_14444,N_14071,N_14026);
nand U14445 (N_14445,N_14024,N_14109);
or U14446 (N_14446,N_14120,N_14135);
nor U14447 (N_14447,N_14132,N_14042);
and U14448 (N_14448,N_14155,N_14106);
or U14449 (N_14449,N_14016,N_14019);
nand U14450 (N_14450,N_14181,N_14185);
nor U14451 (N_14451,N_14005,N_14122);
and U14452 (N_14452,N_14225,N_14035);
nand U14453 (N_14453,N_14097,N_14245);
xor U14454 (N_14454,N_14132,N_14205);
or U14455 (N_14455,N_14099,N_14168);
nor U14456 (N_14456,N_14187,N_14242);
and U14457 (N_14457,N_14127,N_14090);
and U14458 (N_14458,N_14220,N_14245);
nor U14459 (N_14459,N_14233,N_14235);
nor U14460 (N_14460,N_14172,N_14071);
or U14461 (N_14461,N_14090,N_14097);
or U14462 (N_14462,N_14039,N_14133);
or U14463 (N_14463,N_14225,N_14024);
nor U14464 (N_14464,N_14059,N_14019);
nand U14465 (N_14465,N_14116,N_14189);
xor U14466 (N_14466,N_14098,N_14075);
xnor U14467 (N_14467,N_14221,N_14103);
or U14468 (N_14468,N_14237,N_14142);
nor U14469 (N_14469,N_14195,N_14104);
or U14470 (N_14470,N_14161,N_14097);
nor U14471 (N_14471,N_14107,N_14138);
nand U14472 (N_14472,N_14105,N_14144);
nand U14473 (N_14473,N_14211,N_14145);
nand U14474 (N_14474,N_14130,N_14098);
xor U14475 (N_14475,N_14035,N_14057);
or U14476 (N_14476,N_14041,N_14194);
and U14477 (N_14477,N_14170,N_14178);
xnor U14478 (N_14478,N_14041,N_14164);
xnor U14479 (N_14479,N_14220,N_14221);
nand U14480 (N_14480,N_14140,N_14205);
or U14481 (N_14481,N_14225,N_14047);
or U14482 (N_14482,N_14098,N_14031);
nor U14483 (N_14483,N_14249,N_14019);
or U14484 (N_14484,N_14049,N_14089);
xnor U14485 (N_14485,N_14240,N_14183);
nor U14486 (N_14486,N_14204,N_14056);
and U14487 (N_14487,N_14129,N_14094);
nand U14488 (N_14488,N_14238,N_14052);
or U14489 (N_14489,N_14147,N_14108);
xor U14490 (N_14490,N_14068,N_14078);
nor U14491 (N_14491,N_14214,N_14156);
or U14492 (N_14492,N_14012,N_14091);
or U14493 (N_14493,N_14208,N_14198);
nor U14494 (N_14494,N_14021,N_14099);
and U14495 (N_14495,N_14053,N_14217);
and U14496 (N_14496,N_14081,N_14045);
nand U14497 (N_14497,N_14131,N_14013);
and U14498 (N_14498,N_14154,N_14137);
and U14499 (N_14499,N_14177,N_14230);
nand U14500 (N_14500,N_14407,N_14485);
xor U14501 (N_14501,N_14412,N_14373);
xnor U14502 (N_14502,N_14411,N_14481);
or U14503 (N_14503,N_14325,N_14324);
and U14504 (N_14504,N_14387,N_14397);
nor U14505 (N_14505,N_14459,N_14454);
nand U14506 (N_14506,N_14429,N_14299);
nor U14507 (N_14507,N_14326,N_14408);
nor U14508 (N_14508,N_14361,N_14496);
or U14509 (N_14509,N_14266,N_14336);
xnor U14510 (N_14510,N_14443,N_14405);
xnor U14511 (N_14511,N_14448,N_14495);
xor U14512 (N_14512,N_14288,N_14271);
and U14513 (N_14513,N_14479,N_14269);
xnor U14514 (N_14514,N_14267,N_14254);
nand U14515 (N_14515,N_14497,N_14435);
nor U14516 (N_14516,N_14450,N_14270);
and U14517 (N_14517,N_14314,N_14418);
nand U14518 (N_14518,N_14434,N_14438);
xnor U14519 (N_14519,N_14331,N_14320);
nand U14520 (N_14520,N_14388,N_14430);
or U14521 (N_14521,N_14385,N_14253);
nand U14522 (N_14522,N_14306,N_14465);
and U14523 (N_14523,N_14251,N_14482);
or U14524 (N_14524,N_14364,N_14410);
nor U14525 (N_14525,N_14367,N_14303);
xnor U14526 (N_14526,N_14426,N_14280);
nand U14527 (N_14527,N_14451,N_14273);
nor U14528 (N_14528,N_14301,N_14396);
nand U14529 (N_14529,N_14480,N_14276);
nand U14530 (N_14530,N_14359,N_14258);
nand U14531 (N_14531,N_14492,N_14475);
nand U14532 (N_14532,N_14293,N_14460);
and U14533 (N_14533,N_14341,N_14441);
or U14534 (N_14534,N_14277,N_14366);
nand U14535 (N_14535,N_14349,N_14389);
and U14536 (N_14536,N_14468,N_14374);
or U14537 (N_14537,N_14309,N_14463);
xnor U14538 (N_14538,N_14308,N_14456);
xor U14539 (N_14539,N_14297,N_14256);
and U14540 (N_14540,N_14337,N_14488);
nor U14541 (N_14541,N_14310,N_14449);
xor U14542 (N_14542,N_14302,N_14398);
or U14543 (N_14543,N_14436,N_14285);
and U14544 (N_14544,N_14457,N_14313);
nand U14545 (N_14545,N_14427,N_14466);
nor U14546 (N_14546,N_14261,N_14327);
nor U14547 (N_14547,N_14440,N_14358);
and U14548 (N_14548,N_14334,N_14394);
and U14549 (N_14549,N_14379,N_14469);
nand U14550 (N_14550,N_14365,N_14363);
nand U14551 (N_14551,N_14347,N_14343);
and U14552 (N_14552,N_14339,N_14403);
nand U14553 (N_14553,N_14386,N_14432);
and U14554 (N_14554,N_14477,N_14292);
nand U14555 (N_14555,N_14345,N_14372);
xnor U14556 (N_14556,N_14452,N_14491);
and U14557 (N_14557,N_14294,N_14462);
xor U14558 (N_14558,N_14362,N_14317);
or U14559 (N_14559,N_14338,N_14458);
or U14560 (N_14560,N_14395,N_14272);
or U14561 (N_14561,N_14353,N_14470);
nor U14562 (N_14562,N_14255,N_14257);
or U14563 (N_14563,N_14259,N_14431);
xor U14564 (N_14564,N_14445,N_14400);
or U14565 (N_14565,N_14329,N_14490);
xnor U14566 (N_14566,N_14464,N_14473);
nand U14567 (N_14567,N_14305,N_14384);
and U14568 (N_14568,N_14422,N_14252);
nor U14569 (N_14569,N_14274,N_14498);
nand U14570 (N_14570,N_14378,N_14494);
or U14571 (N_14571,N_14442,N_14282);
and U14572 (N_14572,N_14278,N_14493);
and U14573 (N_14573,N_14298,N_14428);
xnor U14574 (N_14574,N_14368,N_14265);
xnor U14575 (N_14575,N_14419,N_14376);
or U14576 (N_14576,N_14381,N_14390);
or U14577 (N_14577,N_14439,N_14319);
or U14578 (N_14578,N_14402,N_14315);
and U14579 (N_14579,N_14332,N_14423);
and U14580 (N_14580,N_14321,N_14377);
nand U14581 (N_14581,N_14356,N_14291);
xnor U14582 (N_14582,N_14420,N_14289);
and U14583 (N_14583,N_14300,N_14401);
nand U14584 (N_14584,N_14416,N_14264);
nand U14585 (N_14585,N_14415,N_14421);
nor U14586 (N_14586,N_14263,N_14433);
and U14587 (N_14587,N_14287,N_14369);
nor U14588 (N_14588,N_14318,N_14323);
and U14589 (N_14589,N_14340,N_14478);
nand U14590 (N_14590,N_14330,N_14425);
and U14591 (N_14591,N_14467,N_14406);
nand U14592 (N_14592,N_14286,N_14455);
nor U14593 (N_14593,N_14447,N_14476);
nor U14594 (N_14594,N_14316,N_14371);
xnor U14595 (N_14595,N_14489,N_14380);
and U14596 (N_14596,N_14360,N_14304);
and U14597 (N_14597,N_14461,N_14486);
or U14598 (N_14598,N_14484,N_14472);
nand U14599 (N_14599,N_14296,N_14295);
and U14600 (N_14600,N_14382,N_14279);
and U14601 (N_14601,N_14348,N_14355);
nand U14602 (N_14602,N_14499,N_14413);
nor U14603 (N_14603,N_14283,N_14357);
xor U14604 (N_14604,N_14417,N_14311);
xor U14605 (N_14605,N_14312,N_14328);
nand U14606 (N_14606,N_14383,N_14453);
and U14607 (N_14607,N_14444,N_14414);
xnor U14608 (N_14608,N_14351,N_14409);
and U14609 (N_14609,N_14281,N_14370);
or U14610 (N_14610,N_14275,N_14268);
or U14611 (N_14611,N_14284,N_14354);
nand U14612 (N_14612,N_14424,N_14250);
xnor U14613 (N_14613,N_14290,N_14483);
and U14614 (N_14614,N_14307,N_14352);
nor U14615 (N_14615,N_14404,N_14392);
nor U14616 (N_14616,N_14399,N_14262);
nand U14617 (N_14617,N_14346,N_14487);
nor U14618 (N_14618,N_14260,N_14446);
and U14619 (N_14619,N_14335,N_14474);
xnor U14620 (N_14620,N_14471,N_14322);
xnor U14621 (N_14621,N_14350,N_14437);
or U14622 (N_14622,N_14391,N_14333);
nand U14623 (N_14623,N_14344,N_14342);
or U14624 (N_14624,N_14393,N_14375);
and U14625 (N_14625,N_14374,N_14345);
and U14626 (N_14626,N_14277,N_14396);
nor U14627 (N_14627,N_14429,N_14383);
and U14628 (N_14628,N_14483,N_14319);
or U14629 (N_14629,N_14313,N_14270);
nor U14630 (N_14630,N_14423,N_14266);
or U14631 (N_14631,N_14265,N_14454);
nand U14632 (N_14632,N_14320,N_14304);
or U14633 (N_14633,N_14318,N_14420);
nor U14634 (N_14634,N_14261,N_14482);
and U14635 (N_14635,N_14305,N_14353);
nand U14636 (N_14636,N_14327,N_14389);
nor U14637 (N_14637,N_14480,N_14375);
nor U14638 (N_14638,N_14377,N_14369);
or U14639 (N_14639,N_14407,N_14476);
nand U14640 (N_14640,N_14393,N_14398);
xor U14641 (N_14641,N_14417,N_14377);
nor U14642 (N_14642,N_14338,N_14362);
xnor U14643 (N_14643,N_14323,N_14328);
nor U14644 (N_14644,N_14478,N_14293);
nor U14645 (N_14645,N_14497,N_14404);
xnor U14646 (N_14646,N_14452,N_14332);
nand U14647 (N_14647,N_14495,N_14442);
and U14648 (N_14648,N_14346,N_14319);
xor U14649 (N_14649,N_14426,N_14369);
xor U14650 (N_14650,N_14280,N_14284);
nand U14651 (N_14651,N_14331,N_14338);
or U14652 (N_14652,N_14444,N_14486);
or U14653 (N_14653,N_14463,N_14283);
nand U14654 (N_14654,N_14437,N_14336);
and U14655 (N_14655,N_14417,N_14354);
xor U14656 (N_14656,N_14456,N_14284);
nor U14657 (N_14657,N_14443,N_14256);
or U14658 (N_14658,N_14327,N_14408);
and U14659 (N_14659,N_14438,N_14359);
nor U14660 (N_14660,N_14330,N_14395);
nor U14661 (N_14661,N_14253,N_14431);
nand U14662 (N_14662,N_14382,N_14266);
nor U14663 (N_14663,N_14344,N_14387);
xnor U14664 (N_14664,N_14470,N_14455);
nor U14665 (N_14665,N_14261,N_14274);
nor U14666 (N_14666,N_14332,N_14340);
nor U14667 (N_14667,N_14355,N_14451);
and U14668 (N_14668,N_14466,N_14269);
nor U14669 (N_14669,N_14298,N_14425);
xor U14670 (N_14670,N_14462,N_14279);
nor U14671 (N_14671,N_14496,N_14329);
or U14672 (N_14672,N_14266,N_14484);
nor U14673 (N_14673,N_14404,N_14363);
nor U14674 (N_14674,N_14385,N_14415);
and U14675 (N_14675,N_14268,N_14328);
or U14676 (N_14676,N_14474,N_14376);
nand U14677 (N_14677,N_14272,N_14475);
and U14678 (N_14678,N_14415,N_14443);
nor U14679 (N_14679,N_14341,N_14368);
nor U14680 (N_14680,N_14495,N_14474);
nor U14681 (N_14681,N_14288,N_14469);
nor U14682 (N_14682,N_14309,N_14420);
or U14683 (N_14683,N_14323,N_14280);
nor U14684 (N_14684,N_14371,N_14254);
xor U14685 (N_14685,N_14413,N_14489);
xnor U14686 (N_14686,N_14499,N_14349);
nor U14687 (N_14687,N_14268,N_14305);
nor U14688 (N_14688,N_14394,N_14438);
and U14689 (N_14689,N_14406,N_14271);
nor U14690 (N_14690,N_14490,N_14395);
xnor U14691 (N_14691,N_14355,N_14266);
nor U14692 (N_14692,N_14495,N_14281);
nand U14693 (N_14693,N_14476,N_14373);
nor U14694 (N_14694,N_14320,N_14462);
or U14695 (N_14695,N_14410,N_14368);
or U14696 (N_14696,N_14381,N_14481);
xnor U14697 (N_14697,N_14422,N_14298);
and U14698 (N_14698,N_14412,N_14392);
nor U14699 (N_14699,N_14323,N_14326);
xor U14700 (N_14700,N_14366,N_14252);
and U14701 (N_14701,N_14487,N_14459);
and U14702 (N_14702,N_14322,N_14372);
or U14703 (N_14703,N_14274,N_14437);
xor U14704 (N_14704,N_14314,N_14388);
nand U14705 (N_14705,N_14397,N_14276);
or U14706 (N_14706,N_14457,N_14279);
xnor U14707 (N_14707,N_14334,N_14298);
and U14708 (N_14708,N_14320,N_14258);
xnor U14709 (N_14709,N_14416,N_14417);
or U14710 (N_14710,N_14467,N_14310);
or U14711 (N_14711,N_14289,N_14305);
or U14712 (N_14712,N_14430,N_14351);
or U14713 (N_14713,N_14460,N_14396);
nor U14714 (N_14714,N_14409,N_14389);
or U14715 (N_14715,N_14327,N_14378);
nor U14716 (N_14716,N_14413,N_14424);
nor U14717 (N_14717,N_14316,N_14280);
nor U14718 (N_14718,N_14332,N_14375);
nor U14719 (N_14719,N_14414,N_14252);
nor U14720 (N_14720,N_14381,N_14449);
nor U14721 (N_14721,N_14367,N_14453);
and U14722 (N_14722,N_14308,N_14386);
or U14723 (N_14723,N_14297,N_14302);
nor U14724 (N_14724,N_14333,N_14470);
and U14725 (N_14725,N_14379,N_14428);
xor U14726 (N_14726,N_14335,N_14492);
or U14727 (N_14727,N_14297,N_14291);
nand U14728 (N_14728,N_14390,N_14334);
nor U14729 (N_14729,N_14320,N_14350);
xor U14730 (N_14730,N_14303,N_14321);
nor U14731 (N_14731,N_14363,N_14298);
or U14732 (N_14732,N_14454,N_14453);
xnor U14733 (N_14733,N_14476,N_14484);
nand U14734 (N_14734,N_14490,N_14493);
nor U14735 (N_14735,N_14294,N_14263);
and U14736 (N_14736,N_14489,N_14352);
and U14737 (N_14737,N_14328,N_14387);
and U14738 (N_14738,N_14288,N_14266);
nor U14739 (N_14739,N_14458,N_14277);
xor U14740 (N_14740,N_14263,N_14396);
nor U14741 (N_14741,N_14453,N_14403);
nor U14742 (N_14742,N_14420,N_14337);
nor U14743 (N_14743,N_14255,N_14352);
or U14744 (N_14744,N_14296,N_14471);
and U14745 (N_14745,N_14386,N_14381);
xnor U14746 (N_14746,N_14275,N_14301);
xnor U14747 (N_14747,N_14385,N_14254);
and U14748 (N_14748,N_14294,N_14451);
nand U14749 (N_14749,N_14395,N_14250);
and U14750 (N_14750,N_14669,N_14532);
and U14751 (N_14751,N_14585,N_14717);
nand U14752 (N_14752,N_14715,N_14681);
and U14753 (N_14753,N_14539,N_14619);
nand U14754 (N_14754,N_14725,N_14566);
nand U14755 (N_14755,N_14616,N_14579);
xnor U14756 (N_14756,N_14576,N_14559);
nand U14757 (N_14757,N_14500,N_14688);
and U14758 (N_14758,N_14660,N_14560);
or U14759 (N_14759,N_14695,N_14561);
xor U14760 (N_14760,N_14544,N_14718);
nand U14761 (N_14761,N_14605,N_14513);
nor U14762 (N_14762,N_14656,N_14700);
nor U14763 (N_14763,N_14506,N_14541);
or U14764 (N_14764,N_14524,N_14708);
nor U14765 (N_14765,N_14522,N_14680);
nor U14766 (N_14766,N_14535,N_14683);
nand U14767 (N_14767,N_14567,N_14523);
or U14768 (N_14768,N_14531,N_14729);
nand U14769 (N_14769,N_14594,N_14657);
or U14770 (N_14770,N_14623,N_14546);
nand U14771 (N_14771,N_14586,N_14595);
or U14772 (N_14772,N_14554,N_14597);
nand U14773 (N_14773,N_14732,N_14687);
nand U14774 (N_14774,N_14658,N_14525);
and U14775 (N_14775,N_14550,N_14599);
nand U14776 (N_14776,N_14507,N_14721);
xor U14777 (N_14777,N_14650,N_14592);
nand U14778 (N_14778,N_14588,N_14611);
nand U14779 (N_14779,N_14565,N_14583);
and U14780 (N_14780,N_14555,N_14728);
nor U14781 (N_14781,N_14644,N_14590);
nand U14782 (N_14782,N_14502,N_14711);
nor U14783 (N_14783,N_14724,N_14572);
nor U14784 (N_14784,N_14543,N_14664);
or U14785 (N_14785,N_14519,N_14662);
nand U14786 (N_14786,N_14659,N_14747);
and U14787 (N_14787,N_14686,N_14508);
nor U14788 (N_14788,N_14704,N_14614);
or U14789 (N_14789,N_14604,N_14581);
nand U14790 (N_14790,N_14549,N_14661);
and U14791 (N_14791,N_14719,N_14749);
nor U14792 (N_14792,N_14629,N_14625);
nor U14793 (N_14793,N_14564,N_14591);
and U14794 (N_14794,N_14568,N_14690);
and U14795 (N_14795,N_14505,N_14639);
or U14796 (N_14796,N_14510,N_14557);
nand U14797 (N_14797,N_14638,N_14726);
and U14798 (N_14798,N_14563,N_14624);
xor U14799 (N_14799,N_14735,N_14736);
and U14800 (N_14800,N_14710,N_14696);
nor U14801 (N_14801,N_14533,N_14636);
nand U14802 (N_14802,N_14530,N_14642);
nand U14803 (N_14803,N_14635,N_14528);
nor U14804 (N_14804,N_14622,N_14621);
nor U14805 (N_14805,N_14677,N_14734);
and U14806 (N_14806,N_14655,N_14534);
nor U14807 (N_14807,N_14640,N_14692);
and U14808 (N_14808,N_14698,N_14529);
nor U14809 (N_14809,N_14628,N_14504);
or U14810 (N_14810,N_14620,N_14731);
nor U14811 (N_14811,N_14733,N_14648);
and U14812 (N_14812,N_14521,N_14612);
nor U14813 (N_14813,N_14551,N_14679);
nand U14814 (N_14814,N_14697,N_14503);
or U14815 (N_14815,N_14702,N_14615);
or U14816 (N_14816,N_14509,N_14675);
xnor U14817 (N_14817,N_14699,N_14518);
xor U14818 (N_14818,N_14527,N_14577);
nand U14819 (N_14819,N_14632,N_14740);
xnor U14820 (N_14820,N_14608,N_14501);
and U14821 (N_14821,N_14556,N_14601);
or U14822 (N_14822,N_14512,N_14516);
nand U14823 (N_14823,N_14654,N_14693);
nand U14824 (N_14824,N_14553,N_14670);
and U14825 (N_14825,N_14709,N_14653);
nor U14826 (N_14826,N_14743,N_14575);
nor U14827 (N_14827,N_14671,N_14584);
or U14828 (N_14828,N_14649,N_14589);
nor U14829 (N_14829,N_14598,N_14515);
nand U14830 (N_14830,N_14637,N_14730);
nand U14831 (N_14831,N_14691,N_14547);
nand U14832 (N_14832,N_14600,N_14582);
nand U14833 (N_14833,N_14537,N_14744);
nor U14834 (N_14834,N_14526,N_14552);
xnor U14835 (N_14835,N_14727,N_14517);
nor U14836 (N_14836,N_14705,N_14722);
nor U14837 (N_14837,N_14651,N_14746);
xor U14838 (N_14838,N_14536,N_14573);
xor U14839 (N_14839,N_14706,N_14684);
nand U14840 (N_14840,N_14720,N_14627);
or U14841 (N_14841,N_14742,N_14748);
or U14842 (N_14842,N_14665,N_14646);
nor U14843 (N_14843,N_14542,N_14666);
xnor U14844 (N_14844,N_14689,N_14558);
nor U14845 (N_14845,N_14538,N_14682);
xor U14846 (N_14846,N_14574,N_14667);
xnor U14847 (N_14847,N_14737,N_14676);
xor U14848 (N_14848,N_14703,N_14712);
nor U14849 (N_14849,N_14641,N_14741);
xor U14850 (N_14850,N_14645,N_14607);
and U14851 (N_14851,N_14685,N_14602);
nor U14852 (N_14852,N_14603,N_14609);
nor U14853 (N_14853,N_14569,N_14618);
or U14854 (N_14854,N_14694,N_14606);
and U14855 (N_14855,N_14634,N_14745);
nor U14856 (N_14856,N_14714,N_14570);
xnor U14857 (N_14857,N_14562,N_14548);
xnor U14858 (N_14858,N_14578,N_14626);
xor U14859 (N_14859,N_14663,N_14596);
or U14860 (N_14860,N_14593,N_14514);
or U14861 (N_14861,N_14701,N_14571);
or U14862 (N_14862,N_14739,N_14668);
and U14863 (N_14863,N_14647,N_14673);
nand U14864 (N_14864,N_14545,N_14723);
xnor U14865 (N_14865,N_14738,N_14707);
xnor U14866 (N_14866,N_14520,N_14613);
xnor U14867 (N_14867,N_14674,N_14716);
nor U14868 (N_14868,N_14633,N_14540);
or U14869 (N_14869,N_14643,N_14672);
xor U14870 (N_14870,N_14713,N_14630);
xor U14871 (N_14871,N_14610,N_14587);
nand U14872 (N_14872,N_14617,N_14511);
nor U14873 (N_14873,N_14678,N_14580);
and U14874 (N_14874,N_14652,N_14631);
nand U14875 (N_14875,N_14525,N_14639);
nand U14876 (N_14876,N_14718,N_14553);
nand U14877 (N_14877,N_14666,N_14576);
and U14878 (N_14878,N_14702,N_14574);
xnor U14879 (N_14879,N_14712,N_14612);
nor U14880 (N_14880,N_14530,N_14567);
nand U14881 (N_14881,N_14561,N_14538);
nor U14882 (N_14882,N_14565,N_14719);
xnor U14883 (N_14883,N_14745,N_14522);
nand U14884 (N_14884,N_14527,N_14518);
nand U14885 (N_14885,N_14617,N_14672);
and U14886 (N_14886,N_14517,N_14648);
nor U14887 (N_14887,N_14609,N_14552);
or U14888 (N_14888,N_14597,N_14616);
or U14889 (N_14889,N_14521,N_14507);
xor U14890 (N_14890,N_14593,N_14688);
nand U14891 (N_14891,N_14588,N_14678);
or U14892 (N_14892,N_14628,N_14578);
xnor U14893 (N_14893,N_14649,N_14677);
xnor U14894 (N_14894,N_14637,N_14608);
nand U14895 (N_14895,N_14619,N_14738);
nand U14896 (N_14896,N_14734,N_14656);
xor U14897 (N_14897,N_14597,N_14601);
or U14898 (N_14898,N_14645,N_14552);
and U14899 (N_14899,N_14651,N_14654);
nand U14900 (N_14900,N_14646,N_14614);
nand U14901 (N_14901,N_14617,N_14581);
or U14902 (N_14902,N_14735,N_14667);
nor U14903 (N_14903,N_14594,N_14660);
and U14904 (N_14904,N_14727,N_14719);
or U14905 (N_14905,N_14691,N_14692);
and U14906 (N_14906,N_14535,N_14630);
and U14907 (N_14907,N_14706,N_14629);
xor U14908 (N_14908,N_14696,N_14624);
nor U14909 (N_14909,N_14733,N_14727);
nand U14910 (N_14910,N_14607,N_14732);
xor U14911 (N_14911,N_14740,N_14611);
or U14912 (N_14912,N_14741,N_14708);
and U14913 (N_14913,N_14704,N_14641);
nand U14914 (N_14914,N_14520,N_14596);
and U14915 (N_14915,N_14668,N_14505);
or U14916 (N_14916,N_14559,N_14741);
or U14917 (N_14917,N_14671,N_14610);
and U14918 (N_14918,N_14624,N_14627);
or U14919 (N_14919,N_14597,N_14602);
or U14920 (N_14920,N_14739,N_14721);
or U14921 (N_14921,N_14621,N_14581);
xor U14922 (N_14922,N_14665,N_14659);
or U14923 (N_14923,N_14541,N_14525);
xnor U14924 (N_14924,N_14551,N_14636);
xor U14925 (N_14925,N_14708,N_14609);
nor U14926 (N_14926,N_14554,N_14740);
xnor U14927 (N_14927,N_14517,N_14647);
nor U14928 (N_14928,N_14583,N_14701);
nand U14929 (N_14929,N_14581,N_14601);
nand U14930 (N_14930,N_14535,N_14666);
nand U14931 (N_14931,N_14511,N_14716);
nand U14932 (N_14932,N_14501,N_14538);
nand U14933 (N_14933,N_14508,N_14747);
or U14934 (N_14934,N_14674,N_14604);
or U14935 (N_14935,N_14547,N_14620);
nor U14936 (N_14936,N_14549,N_14603);
or U14937 (N_14937,N_14650,N_14529);
or U14938 (N_14938,N_14724,N_14733);
nor U14939 (N_14939,N_14542,N_14635);
and U14940 (N_14940,N_14724,N_14502);
xnor U14941 (N_14941,N_14598,N_14622);
or U14942 (N_14942,N_14575,N_14646);
or U14943 (N_14943,N_14736,N_14605);
nor U14944 (N_14944,N_14636,N_14676);
nand U14945 (N_14945,N_14748,N_14624);
xor U14946 (N_14946,N_14605,N_14611);
xnor U14947 (N_14947,N_14578,N_14534);
nor U14948 (N_14948,N_14572,N_14732);
or U14949 (N_14949,N_14523,N_14503);
xor U14950 (N_14950,N_14501,N_14601);
nor U14951 (N_14951,N_14730,N_14538);
or U14952 (N_14952,N_14503,N_14558);
or U14953 (N_14953,N_14729,N_14699);
nor U14954 (N_14954,N_14590,N_14591);
or U14955 (N_14955,N_14581,N_14623);
xor U14956 (N_14956,N_14637,N_14538);
or U14957 (N_14957,N_14747,N_14688);
nor U14958 (N_14958,N_14595,N_14539);
and U14959 (N_14959,N_14541,N_14707);
xor U14960 (N_14960,N_14608,N_14739);
xor U14961 (N_14961,N_14525,N_14501);
or U14962 (N_14962,N_14606,N_14648);
or U14963 (N_14963,N_14505,N_14636);
or U14964 (N_14964,N_14546,N_14648);
and U14965 (N_14965,N_14585,N_14693);
nand U14966 (N_14966,N_14669,N_14576);
and U14967 (N_14967,N_14675,N_14601);
and U14968 (N_14968,N_14734,N_14544);
or U14969 (N_14969,N_14605,N_14594);
xnor U14970 (N_14970,N_14696,N_14632);
and U14971 (N_14971,N_14728,N_14667);
nor U14972 (N_14972,N_14749,N_14506);
and U14973 (N_14973,N_14707,N_14521);
xor U14974 (N_14974,N_14544,N_14740);
xnor U14975 (N_14975,N_14508,N_14535);
xnor U14976 (N_14976,N_14744,N_14681);
xor U14977 (N_14977,N_14731,N_14722);
and U14978 (N_14978,N_14518,N_14717);
or U14979 (N_14979,N_14581,N_14661);
xor U14980 (N_14980,N_14664,N_14705);
and U14981 (N_14981,N_14693,N_14676);
xor U14982 (N_14982,N_14516,N_14704);
nor U14983 (N_14983,N_14569,N_14589);
and U14984 (N_14984,N_14609,N_14560);
xor U14985 (N_14985,N_14603,N_14682);
nor U14986 (N_14986,N_14636,N_14711);
and U14987 (N_14987,N_14547,N_14571);
nand U14988 (N_14988,N_14544,N_14551);
xor U14989 (N_14989,N_14558,N_14654);
nand U14990 (N_14990,N_14749,N_14670);
nand U14991 (N_14991,N_14639,N_14647);
nor U14992 (N_14992,N_14628,N_14743);
xor U14993 (N_14993,N_14597,N_14733);
nand U14994 (N_14994,N_14569,N_14723);
or U14995 (N_14995,N_14670,N_14738);
and U14996 (N_14996,N_14655,N_14577);
and U14997 (N_14997,N_14652,N_14541);
or U14998 (N_14998,N_14659,N_14657);
nand U14999 (N_14999,N_14632,N_14714);
nor UO_0 (O_0,N_14802,N_14791);
and UO_1 (O_1,N_14772,N_14845);
nand UO_2 (O_2,N_14858,N_14953);
nand UO_3 (O_3,N_14971,N_14911);
nor UO_4 (O_4,N_14918,N_14872);
and UO_5 (O_5,N_14927,N_14904);
nor UO_6 (O_6,N_14805,N_14917);
or UO_7 (O_7,N_14929,N_14877);
nand UO_8 (O_8,N_14771,N_14849);
or UO_9 (O_9,N_14826,N_14905);
and UO_10 (O_10,N_14921,N_14869);
xor UO_11 (O_11,N_14989,N_14922);
or UO_12 (O_12,N_14874,N_14897);
or UO_13 (O_13,N_14907,N_14956);
or UO_14 (O_14,N_14835,N_14761);
xnor UO_15 (O_15,N_14993,N_14962);
xnor UO_16 (O_16,N_14836,N_14892);
and UO_17 (O_17,N_14999,N_14964);
nor UO_18 (O_18,N_14759,N_14972);
and UO_19 (O_19,N_14886,N_14768);
nand UO_20 (O_20,N_14803,N_14983);
or UO_21 (O_21,N_14899,N_14843);
xor UO_22 (O_22,N_14920,N_14878);
or UO_23 (O_23,N_14873,N_14808);
nor UO_24 (O_24,N_14861,N_14955);
and UO_25 (O_25,N_14850,N_14949);
xnor UO_26 (O_26,N_14903,N_14751);
and UO_27 (O_27,N_14839,N_14821);
xnor UO_28 (O_28,N_14887,N_14965);
and UO_29 (O_29,N_14851,N_14984);
and UO_30 (O_30,N_14875,N_14994);
or UO_31 (O_31,N_14818,N_14941);
nand UO_32 (O_32,N_14856,N_14752);
nor UO_33 (O_33,N_14963,N_14770);
nor UO_34 (O_34,N_14909,N_14944);
or UO_35 (O_35,N_14975,N_14914);
nand UO_36 (O_36,N_14754,N_14978);
nand UO_37 (O_37,N_14789,N_14884);
xnor UO_38 (O_38,N_14915,N_14837);
xor UO_39 (O_39,N_14866,N_14782);
or UO_40 (O_40,N_14982,N_14912);
or UO_41 (O_41,N_14783,N_14823);
nand UO_42 (O_42,N_14868,N_14779);
and UO_43 (O_43,N_14812,N_14902);
nor UO_44 (O_44,N_14801,N_14906);
xnor UO_45 (O_45,N_14847,N_14937);
or UO_46 (O_46,N_14774,N_14908);
xnor UO_47 (O_47,N_14781,N_14763);
and UO_48 (O_48,N_14926,N_14940);
nor UO_49 (O_49,N_14936,N_14952);
nand UO_50 (O_50,N_14777,N_14829);
or UO_51 (O_51,N_14784,N_14811);
nor UO_52 (O_52,N_14852,N_14996);
or UO_53 (O_53,N_14894,N_14797);
and UO_54 (O_54,N_14998,N_14976);
nand UO_55 (O_55,N_14825,N_14961);
or UO_56 (O_56,N_14788,N_14833);
nand UO_57 (O_57,N_14824,N_14848);
and UO_58 (O_58,N_14819,N_14795);
xor UO_59 (O_59,N_14991,N_14986);
nor UO_60 (O_60,N_14932,N_14854);
or UO_61 (O_61,N_14910,N_14959);
nand UO_62 (O_62,N_14809,N_14780);
nor UO_63 (O_63,N_14753,N_14890);
nor UO_64 (O_64,N_14974,N_14860);
or UO_65 (O_65,N_14773,N_14947);
nor UO_66 (O_66,N_14924,N_14841);
xnor UO_67 (O_67,N_14977,N_14787);
or UO_68 (O_68,N_14804,N_14762);
nand UO_69 (O_69,N_14951,N_14756);
or UO_70 (O_70,N_14838,N_14997);
xnor UO_71 (O_71,N_14880,N_14816);
and UO_72 (O_72,N_14969,N_14806);
xor UO_73 (O_73,N_14867,N_14883);
or UO_74 (O_74,N_14948,N_14966);
nor UO_75 (O_75,N_14980,N_14815);
nand UO_76 (O_76,N_14817,N_14992);
nand UO_77 (O_77,N_14985,N_14798);
or UO_78 (O_78,N_14960,N_14946);
xnor UO_79 (O_79,N_14925,N_14785);
nand UO_80 (O_80,N_14935,N_14794);
xnor UO_81 (O_81,N_14765,N_14973);
xor UO_82 (O_82,N_14786,N_14990);
xnor UO_83 (O_83,N_14755,N_14876);
xnor UO_84 (O_84,N_14827,N_14981);
nor UO_85 (O_85,N_14931,N_14810);
and UO_86 (O_86,N_14919,N_14865);
xor UO_87 (O_87,N_14813,N_14913);
or UO_88 (O_88,N_14928,N_14750);
or UO_89 (O_89,N_14893,N_14954);
and UO_90 (O_90,N_14855,N_14830);
xnor UO_91 (O_91,N_14933,N_14834);
or UO_92 (O_92,N_14846,N_14842);
nand UO_93 (O_93,N_14840,N_14776);
nor UO_94 (O_94,N_14831,N_14853);
nand UO_95 (O_95,N_14968,N_14945);
and UO_96 (O_96,N_14881,N_14967);
and UO_97 (O_97,N_14970,N_14820);
nand UO_98 (O_98,N_14870,N_14882);
and UO_99 (O_99,N_14988,N_14895);
and UO_100 (O_100,N_14862,N_14942);
nor UO_101 (O_101,N_14930,N_14828);
and UO_102 (O_102,N_14943,N_14950);
nand UO_103 (O_103,N_14934,N_14995);
and UO_104 (O_104,N_14885,N_14857);
nor UO_105 (O_105,N_14822,N_14979);
xor UO_106 (O_106,N_14916,N_14958);
xor UO_107 (O_107,N_14799,N_14864);
xnor UO_108 (O_108,N_14987,N_14863);
nor UO_109 (O_109,N_14859,N_14767);
and UO_110 (O_110,N_14790,N_14923);
or UO_111 (O_111,N_14879,N_14792);
and UO_112 (O_112,N_14889,N_14775);
xnor UO_113 (O_113,N_14814,N_14957);
nor UO_114 (O_114,N_14796,N_14888);
xor UO_115 (O_115,N_14901,N_14891);
or UO_116 (O_116,N_14757,N_14800);
and UO_117 (O_117,N_14807,N_14900);
nor UO_118 (O_118,N_14758,N_14896);
or UO_119 (O_119,N_14769,N_14844);
or UO_120 (O_120,N_14939,N_14793);
or UO_121 (O_121,N_14898,N_14832);
or UO_122 (O_122,N_14871,N_14778);
nor UO_123 (O_123,N_14760,N_14766);
nand UO_124 (O_124,N_14938,N_14764);
nor UO_125 (O_125,N_14973,N_14805);
nand UO_126 (O_126,N_14866,N_14787);
nor UO_127 (O_127,N_14775,N_14956);
or UO_128 (O_128,N_14947,N_14989);
and UO_129 (O_129,N_14854,N_14832);
or UO_130 (O_130,N_14825,N_14979);
nand UO_131 (O_131,N_14794,N_14950);
nand UO_132 (O_132,N_14759,N_14800);
or UO_133 (O_133,N_14841,N_14901);
and UO_134 (O_134,N_14977,N_14968);
or UO_135 (O_135,N_14762,N_14982);
nor UO_136 (O_136,N_14913,N_14756);
and UO_137 (O_137,N_14885,N_14892);
and UO_138 (O_138,N_14759,N_14939);
nand UO_139 (O_139,N_14940,N_14797);
or UO_140 (O_140,N_14854,N_14947);
nand UO_141 (O_141,N_14855,N_14932);
xor UO_142 (O_142,N_14866,N_14948);
nor UO_143 (O_143,N_14807,N_14769);
or UO_144 (O_144,N_14989,N_14921);
nor UO_145 (O_145,N_14971,N_14976);
nand UO_146 (O_146,N_14779,N_14873);
and UO_147 (O_147,N_14982,N_14819);
nand UO_148 (O_148,N_14759,N_14956);
xnor UO_149 (O_149,N_14950,N_14946);
xnor UO_150 (O_150,N_14881,N_14842);
and UO_151 (O_151,N_14795,N_14757);
xnor UO_152 (O_152,N_14920,N_14947);
xnor UO_153 (O_153,N_14968,N_14881);
and UO_154 (O_154,N_14886,N_14943);
or UO_155 (O_155,N_14908,N_14970);
nand UO_156 (O_156,N_14970,N_14991);
xnor UO_157 (O_157,N_14753,N_14914);
and UO_158 (O_158,N_14750,N_14816);
nand UO_159 (O_159,N_14923,N_14803);
nand UO_160 (O_160,N_14822,N_14945);
or UO_161 (O_161,N_14781,N_14814);
nor UO_162 (O_162,N_14964,N_14785);
xnor UO_163 (O_163,N_14756,N_14774);
xnor UO_164 (O_164,N_14981,N_14814);
and UO_165 (O_165,N_14938,N_14769);
nand UO_166 (O_166,N_14851,N_14926);
nand UO_167 (O_167,N_14777,N_14763);
or UO_168 (O_168,N_14877,N_14782);
and UO_169 (O_169,N_14767,N_14932);
and UO_170 (O_170,N_14830,N_14876);
nand UO_171 (O_171,N_14791,N_14995);
and UO_172 (O_172,N_14862,N_14941);
xnor UO_173 (O_173,N_14764,N_14920);
or UO_174 (O_174,N_14755,N_14877);
and UO_175 (O_175,N_14810,N_14794);
xnor UO_176 (O_176,N_14758,N_14880);
nor UO_177 (O_177,N_14956,N_14833);
or UO_178 (O_178,N_14836,N_14819);
nand UO_179 (O_179,N_14983,N_14999);
or UO_180 (O_180,N_14879,N_14795);
nand UO_181 (O_181,N_14930,N_14904);
xnor UO_182 (O_182,N_14782,N_14869);
or UO_183 (O_183,N_14822,N_14954);
xnor UO_184 (O_184,N_14807,N_14798);
nand UO_185 (O_185,N_14865,N_14875);
or UO_186 (O_186,N_14750,N_14804);
xor UO_187 (O_187,N_14998,N_14963);
or UO_188 (O_188,N_14996,N_14955);
or UO_189 (O_189,N_14846,N_14784);
and UO_190 (O_190,N_14857,N_14767);
nor UO_191 (O_191,N_14793,N_14955);
and UO_192 (O_192,N_14993,N_14791);
nand UO_193 (O_193,N_14824,N_14856);
nor UO_194 (O_194,N_14767,N_14852);
xor UO_195 (O_195,N_14966,N_14871);
and UO_196 (O_196,N_14936,N_14946);
xnor UO_197 (O_197,N_14919,N_14774);
or UO_198 (O_198,N_14921,N_14844);
xnor UO_199 (O_199,N_14854,N_14815);
xnor UO_200 (O_200,N_14955,N_14981);
xor UO_201 (O_201,N_14820,N_14787);
xor UO_202 (O_202,N_14838,N_14930);
or UO_203 (O_203,N_14939,N_14976);
nor UO_204 (O_204,N_14772,N_14897);
nand UO_205 (O_205,N_14819,N_14897);
nor UO_206 (O_206,N_14805,N_14888);
or UO_207 (O_207,N_14980,N_14936);
xor UO_208 (O_208,N_14840,N_14918);
nor UO_209 (O_209,N_14910,N_14828);
xor UO_210 (O_210,N_14784,N_14853);
nor UO_211 (O_211,N_14854,N_14781);
xor UO_212 (O_212,N_14968,N_14771);
or UO_213 (O_213,N_14873,N_14957);
nand UO_214 (O_214,N_14819,N_14766);
xnor UO_215 (O_215,N_14817,N_14993);
nor UO_216 (O_216,N_14754,N_14949);
nor UO_217 (O_217,N_14958,N_14878);
nand UO_218 (O_218,N_14954,N_14982);
and UO_219 (O_219,N_14980,N_14963);
or UO_220 (O_220,N_14831,N_14842);
xnor UO_221 (O_221,N_14836,N_14769);
xor UO_222 (O_222,N_14764,N_14777);
nor UO_223 (O_223,N_14904,N_14771);
or UO_224 (O_224,N_14964,N_14893);
nand UO_225 (O_225,N_14847,N_14969);
and UO_226 (O_226,N_14807,N_14965);
nor UO_227 (O_227,N_14902,N_14952);
xor UO_228 (O_228,N_14934,N_14933);
or UO_229 (O_229,N_14891,N_14859);
and UO_230 (O_230,N_14946,N_14874);
nand UO_231 (O_231,N_14793,N_14964);
and UO_232 (O_232,N_14861,N_14918);
and UO_233 (O_233,N_14931,N_14973);
and UO_234 (O_234,N_14811,N_14849);
and UO_235 (O_235,N_14943,N_14896);
nor UO_236 (O_236,N_14956,N_14765);
and UO_237 (O_237,N_14799,N_14862);
and UO_238 (O_238,N_14755,N_14993);
and UO_239 (O_239,N_14946,N_14816);
nand UO_240 (O_240,N_14860,N_14925);
nor UO_241 (O_241,N_14874,N_14825);
xnor UO_242 (O_242,N_14915,N_14984);
nor UO_243 (O_243,N_14974,N_14980);
xor UO_244 (O_244,N_14782,N_14963);
nand UO_245 (O_245,N_14895,N_14757);
and UO_246 (O_246,N_14937,N_14928);
and UO_247 (O_247,N_14941,N_14853);
and UO_248 (O_248,N_14994,N_14830);
nand UO_249 (O_249,N_14824,N_14949);
and UO_250 (O_250,N_14776,N_14806);
or UO_251 (O_251,N_14890,N_14938);
nor UO_252 (O_252,N_14861,N_14804);
nand UO_253 (O_253,N_14814,N_14796);
nand UO_254 (O_254,N_14763,N_14857);
xor UO_255 (O_255,N_14985,N_14933);
nand UO_256 (O_256,N_14866,N_14915);
or UO_257 (O_257,N_14846,N_14920);
xnor UO_258 (O_258,N_14822,N_14809);
xnor UO_259 (O_259,N_14786,N_14971);
xnor UO_260 (O_260,N_14813,N_14824);
or UO_261 (O_261,N_14849,N_14920);
nand UO_262 (O_262,N_14849,N_14826);
and UO_263 (O_263,N_14792,N_14779);
nor UO_264 (O_264,N_14915,N_14855);
nand UO_265 (O_265,N_14908,N_14769);
and UO_266 (O_266,N_14802,N_14950);
or UO_267 (O_267,N_14838,N_14904);
xor UO_268 (O_268,N_14911,N_14772);
nand UO_269 (O_269,N_14793,N_14959);
nand UO_270 (O_270,N_14896,N_14989);
nand UO_271 (O_271,N_14872,N_14987);
and UO_272 (O_272,N_14933,N_14770);
and UO_273 (O_273,N_14896,N_14860);
xnor UO_274 (O_274,N_14979,N_14955);
nor UO_275 (O_275,N_14968,N_14925);
nor UO_276 (O_276,N_14916,N_14921);
nand UO_277 (O_277,N_14956,N_14810);
or UO_278 (O_278,N_14930,N_14850);
or UO_279 (O_279,N_14944,N_14940);
and UO_280 (O_280,N_14984,N_14875);
or UO_281 (O_281,N_14923,N_14849);
nand UO_282 (O_282,N_14963,N_14854);
nand UO_283 (O_283,N_14934,N_14932);
nand UO_284 (O_284,N_14897,N_14891);
nor UO_285 (O_285,N_14892,N_14775);
xor UO_286 (O_286,N_14963,N_14929);
nand UO_287 (O_287,N_14825,N_14921);
xor UO_288 (O_288,N_14904,N_14877);
nand UO_289 (O_289,N_14998,N_14899);
nand UO_290 (O_290,N_14826,N_14881);
nor UO_291 (O_291,N_14929,N_14807);
nor UO_292 (O_292,N_14801,N_14841);
nand UO_293 (O_293,N_14807,N_14804);
nor UO_294 (O_294,N_14782,N_14803);
nor UO_295 (O_295,N_14804,N_14806);
nand UO_296 (O_296,N_14818,N_14957);
and UO_297 (O_297,N_14924,N_14809);
xor UO_298 (O_298,N_14898,N_14765);
and UO_299 (O_299,N_14829,N_14854);
and UO_300 (O_300,N_14882,N_14789);
nand UO_301 (O_301,N_14766,N_14991);
or UO_302 (O_302,N_14936,N_14758);
nor UO_303 (O_303,N_14848,N_14877);
or UO_304 (O_304,N_14980,N_14837);
nand UO_305 (O_305,N_14980,N_14916);
and UO_306 (O_306,N_14815,N_14895);
nor UO_307 (O_307,N_14906,N_14819);
nor UO_308 (O_308,N_14825,N_14938);
and UO_309 (O_309,N_14918,N_14979);
or UO_310 (O_310,N_14943,N_14766);
and UO_311 (O_311,N_14767,N_14765);
nand UO_312 (O_312,N_14831,N_14820);
and UO_313 (O_313,N_14960,N_14978);
xor UO_314 (O_314,N_14843,N_14904);
or UO_315 (O_315,N_14838,N_14914);
xor UO_316 (O_316,N_14970,N_14837);
and UO_317 (O_317,N_14908,N_14953);
and UO_318 (O_318,N_14969,N_14866);
xnor UO_319 (O_319,N_14939,N_14753);
and UO_320 (O_320,N_14889,N_14994);
and UO_321 (O_321,N_14898,N_14814);
nand UO_322 (O_322,N_14869,N_14879);
and UO_323 (O_323,N_14901,N_14982);
and UO_324 (O_324,N_14799,N_14895);
xor UO_325 (O_325,N_14918,N_14926);
nor UO_326 (O_326,N_14775,N_14824);
or UO_327 (O_327,N_14813,N_14874);
xnor UO_328 (O_328,N_14975,N_14843);
or UO_329 (O_329,N_14877,N_14867);
and UO_330 (O_330,N_14899,N_14858);
xor UO_331 (O_331,N_14895,N_14857);
nor UO_332 (O_332,N_14838,N_14830);
and UO_333 (O_333,N_14889,N_14837);
xnor UO_334 (O_334,N_14781,N_14949);
nor UO_335 (O_335,N_14824,N_14860);
and UO_336 (O_336,N_14849,N_14837);
nor UO_337 (O_337,N_14966,N_14785);
and UO_338 (O_338,N_14788,N_14767);
nor UO_339 (O_339,N_14887,N_14924);
nand UO_340 (O_340,N_14967,N_14948);
xnor UO_341 (O_341,N_14889,N_14840);
and UO_342 (O_342,N_14831,N_14756);
nand UO_343 (O_343,N_14814,N_14926);
nand UO_344 (O_344,N_14837,N_14956);
nor UO_345 (O_345,N_14831,N_14778);
or UO_346 (O_346,N_14968,N_14756);
and UO_347 (O_347,N_14847,N_14839);
nor UO_348 (O_348,N_14765,N_14842);
and UO_349 (O_349,N_14911,N_14983);
nor UO_350 (O_350,N_14862,N_14972);
nor UO_351 (O_351,N_14878,N_14969);
nor UO_352 (O_352,N_14808,N_14862);
xor UO_353 (O_353,N_14793,N_14991);
and UO_354 (O_354,N_14829,N_14996);
xnor UO_355 (O_355,N_14907,N_14883);
nand UO_356 (O_356,N_14822,N_14902);
nand UO_357 (O_357,N_14853,N_14817);
and UO_358 (O_358,N_14809,N_14975);
or UO_359 (O_359,N_14774,N_14836);
nor UO_360 (O_360,N_14877,N_14756);
nor UO_361 (O_361,N_14790,N_14972);
and UO_362 (O_362,N_14870,N_14768);
and UO_363 (O_363,N_14776,N_14824);
xnor UO_364 (O_364,N_14759,N_14945);
and UO_365 (O_365,N_14969,N_14889);
nor UO_366 (O_366,N_14865,N_14768);
nand UO_367 (O_367,N_14997,N_14946);
xor UO_368 (O_368,N_14983,N_14777);
nand UO_369 (O_369,N_14799,N_14917);
nand UO_370 (O_370,N_14758,N_14785);
xor UO_371 (O_371,N_14805,N_14991);
and UO_372 (O_372,N_14809,N_14999);
or UO_373 (O_373,N_14998,N_14964);
and UO_374 (O_374,N_14966,N_14877);
or UO_375 (O_375,N_14942,N_14859);
and UO_376 (O_376,N_14906,N_14956);
and UO_377 (O_377,N_14891,N_14967);
and UO_378 (O_378,N_14939,N_14970);
nor UO_379 (O_379,N_14825,N_14884);
nor UO_380 (O_380,N_14836,N_14945);
nor UO_381 (O_381,N_14996,N_14907);
and UO_382 (O_382,N_14855,N_14839);
nand UO_383 (O_383,N_14771,N_14764);
nand UO_384 (O_384,N_14929,N_14927);
nor UO_385 (O_385,N_14846,N_14831);
and UO_386 (O_386,N_14863,N_14877);
nor UO_387 (O_387,N_14785,N_14794);
nand UO_388 (O_388,N_14793,N_14835);
nand UO_389 (O_389,N_14936,N_14969);
and UO_390 (O_390,N_14753,N_14936);
or UO_391 (O_391,N_14853,N_14844);
nand UO_392 (O_392,N_14797,N_14772);
nand UO_393 (O_393,N_14881,N_14890);
nor UO_394 (O_394,N_14915,N_14938);
or UO_395 (O_395,N_14792,N_14990);
and UO_396 (O_396,N_14756,N_14994);
nand UO_397 (O_397,N_14921,N_14881);
nor UO_398 (O_398,N_14864,N_14961);
nor UO_399 (O_399,N_14886,N_14770);
or UO_400 (O_400,N_14817,N_14908);
and UO_401 (O_401,N_14753,N_14845);
xnor UO_402 (O_402,N_14856,N_14786);
nand UO_403 (O_403,N_14934,N_14825);
nand UO_404 (O_404,N_14925,N_14984);
and UO_405 (O_405,N_14983,N_14870);
nor UO_406 (O_406,N_14997,N_14973);
nand UO_407 (O_407,N_14972,N_14800);
nor UO_408 (O_408,N_14884,N_14770);
xnor UO_409 (O_409,N_14972,N_14812);
and UO_410 (O_410,N_14843,N_14915);
and UO_411 (O_411,N_14960,N_14871);
or UO_412 (O_412,N_14955,N_14993);
and UO_413 (O_413,N_14838,N_14898);
xor UO_414 (O_414,N_14750,N_14832);
xnor UO_415 (O_415,N_14806,N_14837);
nor UO_416 (O_416,N_14958,N_14793);
or UO_417 (O_417,N_14896,N_14799);
nand UO_418 (O_418,N_14815,N_14940);
or UO_419 (O_419,N_14890,N_14768);
nor UO_420 (O_420,N_14799,N_14885);
and UO_421 (O_421,N_14763,N_14846);
and UO_422 (O_422,N_14834,N_14993);
xor UO_423 (O_423,N_14785,N_14814);
xor UO_424 (O_424,N_14867,N_14825);
xor UO_425 (O_425,N_14891,N_14836);
or UO_426 (O_426,N_14969,N_14989);
xnor UO_427 (O_427,N_14778,N_14789);
xor UO_428 (O_428,N_14908,N_14823);
xnor UO_429 (O_429,N_14798,N_14989);
nand UO_430 (O_430,N_14785,N_14957);
and UO_431 (O_431,N_14779,N_14818);
and UO_432 (O_432,N_14963,N_14939);
nor UO_433 (O_433,N_14779,N_14884);
nand UO_434 (O_434,N_14892,N_14895);
nor UO_435 (O_435,N_14936,N_14778);
and UO_436 (O_436,N_14939,N_14765);
or UO_437 (O_437,N_14935,N_14787);
xor UO_438 (O_438,N_14979,N_14862);
xor UO_439 (O_439,N_14886,N_14942);
nor UO_440 (O_440,N_14817,N_14935);
or UO_441 (O_441,N_14992,N_14814);
or UO_442 (O_442,N_14993,N_14932);
nand UO_443 (O_443,N_14774,N_14867);
nor UO_444 (O_444,N_14964,N_14877);
xnor UO_445 (O_445,N_14783,N_14809);
nor UO_446 (O_446,N_14764,N_14776);
or UO_447 (O_447,N_14769,N_14781);
or UO_448 (O_448,N_14778,N_14811);
nor UO_449 (O_449,N_14825,N_14873);
nor UO_450 (O_450,N_14823,N_14856);
nand UO_451 (O_451,N_14842,N_14979);
nor UO_452 (O_452,N_14987,N_14865);
and UO_453 (O_453,N_14970,N_14921);
nor UO_454 (O_454,N_14981,N_14896);
and UO_455 (O_455,N_14765,N_14945);
nand UO_456 (O_456,N_14924,N_14921);
xor UO_457 (O_457,N_14981,N_14889);
or UO_458 (O_458,N_14904,N_14880);
or UO_459 (O_459,N_14906,N_14835);
nor UO_460 (O_460,N_14841,N_14796);
or UO_461 (O_461,N_14977,N_14828);
xor UO_462 (O_462,N_14845,N_14872);
or UO_463 (O_463,N_14807,N_14812);
nand UO_464 (O_464,N_14835,N_14975);
and UO_465 (O_465,N_14794,N_14819);
nor UO_466 (O_466,N_14956,N_14904);
or UO_467 (O_467,N_14851,N_14799);
nor UO_468 (O_468,N_14876,N_14892);
nand UO_469 (O_469,N_14980,N_14817);
nor UO_470 (O_470,N_14827,N_14944);
or UO_471 (O_471,N_14837,N_14841);
and UO_472 (O_472,N_14934,N_14782);
nor UO_473 (O_473,N_14981,N_14859);
or UO_474 (O_474,N_14992,N_14819);
or UO_475 (O_475,N_14858,N_14836);
and UO_476 (O_476,N_14964,N_14768);
nand UO_477 (O_477,N_14816,N_14949);
and UO_478 (O_478,N_14796,N_14811);
nor UO_479 (O_479,N_14994,N_14896);
and UO_480 (O_480,N_14949,N_14882);
xnor UO_481 (O_481,N_14928,N_14760);
xnor UO_482 (O_482,N_14892,N_14787);
xor UO_483 (O_483,N_14994,N_14921);
nor UO_484 (O_484,N_14929,N_14804);
and UO_485 (O_485,N_14920,N_14803);
and UO_486 (O_486,N_14985,N_14982);
nor UO_487 (O_487,N_14978,N_14768);
and UO_488 (O_488,N_14983,N_14856);
nand UO_489 (O_489,N_14898,N_14833);
and UO_490 (O_490,N_14863,N_14946);
nor UO_491 (O_491,N_14966,N_14993);
nand UO_492 (O_492,N_14858,N_14796);
nor UO_493 (O_493,N_14811,N_14819);
nand UO_494 (O_494,N_14988,N_14951);
xnor UO_495 (O_495,N_14843,N_14838);
nor UO_496 (O_496,N_14839,N_14931);
nor UO_497 (O_497,N_14909,N_14829);
nand UO_498 (O_498,N_14910,N_14990);
nand UO_499 (O_499,N_14928,N_14934);
or UO_500 (O_500,N_14754,N_14959);
and UO_501 (O_501,N_14840,N_14781);
nand UO_502 (O_502,N_14973,N_14874);
nor UO_503 (O_503,N_14822,N_14812);
xor UO_504 (O_504,N_14861,N_14750);
nor UO_505 (O_505,N_14902,N_14784);
or UO_506 (O_506,N_14965,N_14939);
nand UO_507 (O_507,N_14873,N_14956);
nor UO_508 (O_508,N_14936,N_14904);
nor UO_509 (O_509,N_14879,N_14878);
or UO_510 (O_510,N_14810,N_14874);
nor UO_511 (O_511,N_14938,N_14869);
or UO_512 (O_512,N_14878,N_14828);
xor UO_513 (O_513,N_14977,N_14799);
xnor UO_514 (O_514,N_14793,N_14894);
and UO_515 (O_515,N_14999,N_14778);
nand UO_516 (O_516,N_14977,N_14815);
xnor UO_517 (O_517,N_14892,N_14987);
and UO_518 (O_518,N_14922,N_14897);
xor UO_519 (O_519,N_14926,N_14750);
and UO_520 (O_520,N_14924,N_14799);
or UO_521 (O_521,N_14985,N_14986);
or UO_522 (O_522,N_14964,N_14755);
nand UO_523 (O_523,N_14847,N_14976);
xnor UO_524 (O_524,N_14758,N_14938);
nor UO_525 (O_525,N_14888,N_14862);
or UO_526 (O_526,N_14842,N_14770);
and UO_527 (O_527,N_14869,N_14935);
nor UO_528 (O_528,N_14806,N_14977);
and UO_529 (O_529,N_14962,N_14976);
xor UO_530 (O_530,N_14996,N_14983);
nor UO_531 (O_531,N_14857,N_14992);
and UO_532 (O_532,N_14960,N_14807);
nor UO_533 (O_533,N_14908,N_14888);
nand UO_534 (O_534,N_14953,N_14907);
or UO_535 (O_535,N_14756,N_14815);
nand UO_536 (O_536,N_14882,N_14775);
nor UO_537 (O_537,N_14790,N_14945);
xor UO_538 (O_538,N_14883,N_14858);
nor UO_539 (O_539,N_14865,N_14798);
nand UO_540 (O_540,N_14893,N_14832);
nand UO_541 (O_541,N_14965,N_14968);
and UO_542 (O_542,N_14942,N_14866);
and UO_543 (O_543,N_14891,N_14846);
nor UO_544 (O_544,N_14966,N_14905);
and UO_545 (O_545,N_14972,N_14947);
and UO_546 (O_546,N_14832,N_14927);
nor UO_547 (O_547,N_14865,N_14756);
nor UO_548 (O_548,N_14874,N_14849);
or UO_549 (O_549,N_14875,N_14964);
nor UO_550 (O_550,N_14777,N_14966);
nor UO_551 (O_551,N_14819,N_14775);
or UO_552 (O_552,N_14916,N_14842);
xor UO_553 (O_553,N_14768,N_14855);
and UO_554 (O_554,N_14979,N_14872);
nand UO_555 (O_555,N_14868,N_14842);
nor UO_556 (O_556,N_14798,N_14918);
xnor UO_557 (O_557,N_14906,N_14927);
nor UO_558 (O_558,N_14868,N_14946);
nor UO_559 (O_559,N_14806,N_14909);
nor UO_560 (O_560,N_14884,N_14860);
xnor UO_561 (O_561,N_14986,N_14989);
nor UO_562 (O_562,N_14888,N_14768);
nor UO_563 (O_563,N_14951,N_14919);
nand UO_564 (O_564,N_14800,N_14790);
nor UO_565 (O_565,N_14900,N_14878);
nor UO_566 (O_566,N_14808,N_14936);
nor UO_567 (O_567,N_14751,N_14958);
or UO_568 (O_568,N_14823,N_14889);
nand UO_569 (O_569,N_14870,N_14941);
nor UO_570 (O_570,N_14818,N_14915);
or UO_571 (O_571,N_14856,N_14886);
and UO_572 (O_572,N_14864,N_14995);
nor UO_573 (O_573,N_14952,N_14844);
or UO_574 (O_574,N_14878,N_14853);
nand UO_575 (O_575,N_14826,N_14909);
xnor UO_576 (O_576,N_14902,N_14819);
nand UO_577 (O_577,N_14993,N_14777);
and UO_578 (O_578,N_14756,N_14889);
and UO_579 (O_579,N_14822,N_14986);
nor UO_580 (O_580,N_14929,N_14940);
xor UO_581 (O_581,N_14963,N_14806);
nor UO_582 (O_582,N_14895,N_14869);
xor UO_583 (O_583,N_14934,N_14819);
xor UO_584 (O_584,N_14961,N_14831);
xnor UO_585 (O_585,N_14780,N_14818);
nor UO_586 (O_586,N_14922,N_14800);
xor UO_587 (O_587,N_14855,N_14832);
or UO_588 (O_588,N_14786,N_14894);
xor UO_589 (O_589,N_14904,N_14984);
or UO_590 (O_590,N_14956,N_14883);
and UO_591 (O_591,N_14889,N_14839);
or UO_592 (O_592,N_14794,N_14944);
nor UO_593 (O_593,N_14770,N_14882);
and UO_594 (O_594,N_14800,N_14765);
or UO_595 (O_595,N_14858,N_14805);
or UO_596 (O_596,N_14967,N_14827);
xor UO_597 (O_597,N_14959,N_14886);
nand UO_598 (O_598,N_14789,N_14787);
xnor UO_599 (O_599,N_14864,N_14815);
or UO_600 (O_600,N_14822,N_14774);
or UO_601 (O_601,N_14824,N_14980);
and UO_602 (O_602,N_14805,N_14861);
nor UO_603 (O_603,N_14995,N_14917);
and UO_604 (O_604,N_14884,N_14976);
xnor UO_605 (O_605,N_14845,N_14951);
and UO_606 (O_606,N_14792,N_14817);
and UO_607 (O_607,N_14923,N_14871);
nand UO_608 (O_608,N_14783,N_14794);
nand UO_609 (O_609,N_14951,N_14820);
nand UO_610 (O_610,N_14827,N_14801);
xor UO_611 (O_611,N_14966,N_14892);
or UO_612 (O_612,N_14790,N_14839);
or UO_613 (O_613,N_14922,N_14756);
or UO_614 (O_614,N_14881,N_14767);
nand UO_615 (O_615,N_14942,N_14933);
nor UO_616 (O_616,N_14864,N_14940);
nand UO_617 (O_617,N_14898,N_14906);
nand UO_618 (O_618,N_14799,N_14770);
and UO_619 (O_619,N_14837,N_14800);
xor UO_620 (O_620,N_14989,N_14790);
and UO_621 (O_621,N_14985,N_14796);
nor UO_622 (O_622,N_14965,N_14916);
and UO_623 (O_623,N_14838,N_14986);
nand UO_624 (O_624,N_14944,N_14933);
nand UO_625 (O_625,N_14957,N_14938);
xnor UO_626 (O_626,N_14855,N_14871);
nor UO_627 (O_627,N_14984,N_14989);
and UO_628 (O_628,N_14889,N_14898);
or UO_629 (O_629,N_14932,N_14848);
or UO_630 (O_630,N_14953,N_14888);
and UO_631 (O_631,N_14996,N_14859);
or UO_632 (O_632,N_14872,N_14900);
nand UO_633 (O_633,N_14904,N_14965);
nor UO_634 (O_634,N_14954,N_14754);
or UO_635 (O_635,N_14975,N_14955);
and UO_636 (O_636,N_14885,N_14793);
nand UO_637 (O_637,N_14971,N_14761);
and UO_638 (O_638,N_14821,N_14972);
nor UO_639 (O_639,N_14751,N_14839);
nor UO_640 (O_640,N_14846,N_14786);
xnor UO_641 (O_641,N_14892,N_14763);
xor UO_642 (O_642,N_14907,N_14817);
nand UO_643 (O_643,N_14787,N_14811);
nand UO_644 (O_644,N_14889,N_14916);
nor UO_645 (O_645,N_14895,N_14751);
xnor UO_646 (O_646,N_14827,N_14922);
or UO_647 (O_647,N_14963,N_14919);
nor UO_648 (O_648,N_14785,N_14946);
or UO_649 (O_649,N_14780,N_14829);
xnor UO_650 (O_650,N_14878,N_14989);
or UO_651 (O_651,N_14927,N_14858);
or UO_652 (O_652,N_14760,N_14839);
or UO_653 (O_653,N_14851,N_14853);
or UO_654 (O_654,N_14944,N_14879);
nor UO_655 (O_655,N_14918,N_14848);
nor UO_656 (O_656,N_14957,N_14757);
nand UO_657 (O_657,N_14812,N_14866);
nor UO_658 (O_658,N_14813,N_14827);
nand UO_659 (O_659,N_14874,N_14902);
xor UO_660 (O_660,N_14932,N_14944);
or UO_661 (O_661,N_14936,N_14819);
nand UO_662 (O_662,N_14946,N_14757);
nor UO_663 (O_663,N_14800,N_14901);
nand UO_664 (O_664,N_14856,N_14845);
nand UO_665 (O_665,N_14947,N_14988);
nor UO_666 (O_666,N_14764,N_14950);
nor UO_667 (O_667,N_14933,N_14880);
nor UO_668 (O_668,N_14903,N_14992);
xor UO_669 (O_669,N_14815,N_14948);
and UO_670 (O_670,N_14972,N_14908);
nor UO_671 (O_671,N_14873,N_14756);
and UO_672 (O_672,N_14875,N_14787);
nor UO_673 (O_673,N_14806,N_14759);
nand UO_674 (O_674,N_14782,N_14816);
and UO_675 (O_675,N_14880,N_14907);
or UO_676 (O_676,N_14877,N_14835);
nand UO_677 (O_677,N_14807,N_14990);
and UO_678 (O_678,N_14811,N_14950);
nor UO_679 (O_679,N_14874,N_14943);
or UO_680 (O_680,N_14852,N_14887);
and UO_681 (O_681,N_14884,N_14807);
nor UO_682 (O_682,N_14850,N_14755);
xor UO_683 (O_683,N_14857,N_14949);
nand UO_684 (O_684,N_14942,N_14764);
xnor UO_685 (O_685,N_14960,N_14795);
xnor UO_686 (O_686,N_14921,N_14993);
nand UO_687 (O_687,N_14891,N_14874);
nor UO_688 (O_688,N_14780,N_14860);
xnor UO_689 (O_689,N_14770,N_14889);
and UO_690 (O_690,N_14907,N_14831);
nand UO_691 (O_691,N_14811,N_14973);
and UO_692 (O_692,N_14956,N_14914);
and UO_693 (O_693,N_14750,N_14847);
xnor UO_694 (O_694,N_14835,N_14988);
or UO_695 (O_695,N_14917,N_14897);
nor UO_696 (O_696,N_14857,N_14872);
and UO_697 (O_697,N_14925,N_14981);
nand UO_698 (O_698,N_14821,N_14989);
and UO_699 (O_699,N_14930,N_14818);
nand UO_700 (O_700,N_14967,N_14884);
or UO_701 (O_701,N_14823,N_14937);
xnor UO_702 (O_702,N_14766,N_14809);
xor UO_703 (O_703,N_14754,N_14921);
nand UO_704 (O_704,N_14975,N_14984);
nor UO_705 (O_705,N_14880,N_14949);
and UO_706 (O_706,N_14902,N_14780);
xor UO_707 (O_707,N_14819,N_14980);
or UO_708 (O_708,N_14873,N_14882);
and UO_709 (O_709,N_14802,N_14819);
nor UO_710 (O_710,N_14774,N_14899);
nor UO_711 (O_711,N_14955,N_14791);
nand UO_712 (O_712,N_14895,N_14856);
xnor UO_713 (O_713,N_14932,N_14873);
and UO_714 (O_714,N_14880,N_14813);
nand UO_715 (O_715,N_14839,N_14930);
and UO_716 (O_716,N_14785,N_14927);
nand UO_717 (O_717,N_14769,N_14832);
or UO_718 (O_718,N_14950,N_14871);
xnor UO_719 (O_719,N_14855,N_14803);
or UO_720 (O_720,N_14908,N_14800);
and UO_721 (O_721,N_14865,N_14780);
xnor UO_722 (O_722,N_14977,N_14775);
xnor UO_723 (O_723,N_14876,N_14832);
nand UO_724 (O_724,N_14811,N_14866);
nand UO_725 (O_725,N_14786,N_14836);
nor UO_726 (O_726,N_14801,N_14971);
nor UO_727 (O_727,N_14865,N_14851);
or UO_728 (O_728,N_14835,N_14812);
or UO_729 (O_729,N_14895,N_14959);
or UO_730 (O_730,N_14951,N_14993);
nor UO_731 (O_731,N_14919,N_14931);
xnor UO_732 (O_732,N_14921,N_14981);
nand UO_733 (O_733,N_14871,N_14828);
nand UO_734 (O_734,N_14753,N_14924);
and UO_735 (O_735,N_14973,N_14847);
nor UO_736 (O_736,N_14862,N_14828);
and UO_737 (O_737,N_14766,N_14931);
nand UO_738 (O_738,N_14891,N_14860);
and UO_739 (O_739,N_14859,N_14781);
and UO_740 (O_740,N_14847,N_14972);
xor UO_741 (O_741,N_14751,N_14880);
or UO_742 (O_742,N_14985,N_14983);
or UO_743 (O_743,N_14802,N_14977);
nor UO_744 (O_744,N_14822,N_14891);
nor UO_745 (O_745,N_14885,N_14775);
and UO_746 (O_746,N_14864,N_14886);
nand UO_747 (O_747,N_14978,N_14924);
and UO_748 (O_748,N_14835,N_14780);
and UO_749 (O_749,N_14903,N_14896);
nor UO_750 (O_750,N_14869,N_14962);
nor UO_751 (O_751,N_14884,N_14861);
nor UO_752 (O_752,N_14999,N_14969);
or UO_753 (O_753,N_14852,N_14783);
nor UO_754 (O_754,N_14944,N_14857);
xor UO_755 (O_755,N_14937,N_14871);
nand UO_756 (O_756,N_14885,N_14845);
or UO_757 (O_757,N_14880,N_14775);
and UO_758 (O_758,N_14953,N_14940);
or UO_759 (O_759,N_14886,N_14931);
nor UO_760 (O_760,N_14782,N_14971);
xor UO_761 (O_761,N_14994,N_14969);
nand UO_762 (O_762,N_14913,N_14918);
nor UO_763 (O_763,N_14987,N_14763);
xor UO_764 (O_764,N_14816,N_14906);
nand UO_765 (O_765,N_14786,N_14779);
xor UO_766 (O_766,N_14835,N_14936);
nand UO_767 (O_767,N_14808,N_14773);
nor UO_768 (O_768,N_14949,N_14761);
xor UO_769 (O_769,N_14779,N_14810);
and UO_770 (O_770,N_14914,N_14833);
xor UO_771 (O_771,N_14805,N_14996);
nor UO_772 (O_772,N_14969,N_14885);
nand UO_773 (O_773,N_14937,N_14851);
nor UO_774 (O_774,N_14885,N_14777);
or UO_775 (O_775,N_14847,N_14808);
and UO_776 (O_776,N_14936,N_14972);
xor UO_777 (O_777,N_14967,N_14918);
nor UO_778 (O_778,N_14884,N_14907);
and UO_779 (O_779,N_14929,N_14881);
xor UO_780 (O_780,N_14774,N_14906);
and UO_781 (O_781,N_14933,N_14909);
nand UO_782 (O_782,N_14860,N_14871);
xor UO_783 (O_783,N_14931,N_14963);
nand UO_784 (O_784,N_14765,N_14970);
xor UO_785 (O_785,N_14898,N_14792);
nand UO_786 (O_786,N_14832,N_14794);
nand UO_787 (O_787,N_14843,N_14969);
nand UO_788 (O_788,N_14881,N_14859);
and UO_789 (O_789,N_14850,N_14753);
nand UO_790 (O_790,N_14854,N_14814);
or UO_791 (O_791,N_14964,N_14753);
or UO_792 (O_792,N_14845,N_14882);
nor UO_793 (O_793,N_14894,N_14926);
and UO_794 (O_794,N_14999,N_14897);
xnor UO_795 (O_795,N_14879,N_14987);
or UO_796 (O_796,N_14846,N_14946);
or UO_797 (O_797,N_14882,N_14961);
nor UO_798 (O_798,N_14800,N_14884);
and UO_799 (O_799,N_14857,N_14836);
nor UO_800 (O_800,N_14855,N_14861);
or UO_801 (O_801,N_14790,N_14943);
and UO_802 (O_802,N_14868,N_14752);
nand UO_803 (O_803,N_14882,N_14934);
xor UO_804 (O_804,N_14931,N_14945);
or UO_805 (O_805,N_14957,N_14934);
xnor UO_806 (O_806,N_14947,N_14838);
nor UO_807 (O_807,N_14939,N_14803);
or UO_808 (O_808,N_14991,N_14962);
nor UO_809 (O_809,N_14789,N_14945);
nor UO_810 (O_810,N_14854,N_14971);
and UO_811 (O_811,N_14810,N_14924);
xnor UO_812 (O_812,N_14851,N_14785);
xnor UO_813 (O_813,N_14935,N_14919);
or UO_814 (O_814,N_14991,N_14781);
nor UO_815 (O_815,N_14877,N_14947);
xnor UO_816 (O_816,N_14951,N_14973);
and UO_817 (O_817,N_14901,N_14844);
nor UO_818 (O_818,N_14894,N_14899);
nor UO_819 (O_819,N_14829,N_14804);
nand UO_820 (O_820,N_14817,N_14978);
or UO_821 (O_821,N_14937,N_14950);
xor UO_822 (O_822,N_14909,N_14926);
nor UO_823 (O_823,N_14877,N_14775);
and UO_824 (O_824,N_14773,N_14918);
nand UO_825 (O_825,N_14930,N_14830);
nand UO_826 (O_826,N_14831,N_14947);
and UO_827 (O_827,N_14941,N_14803);
nor UO_828 (O_828,N_14835,N_14880);
and UO_829 (O_829,N_14954,N_14988);
nand UO_830 (O_830,N_14919,N_14835);
xor UO_831 (O_831,N_14891,N_14910);
nor UO_832 (O_832,N_14808,N_14887);
nand UO_833 (O_833,N_14790,N_14872);
nand UO_834 (O_834,N_14755,N_14863);
and UO_835 (O_835,N_14795,N_14983);
and UO_836 (O_836,N_14810,N_14994);
and UO_837 (O_837,N_14899,N_14912);
or UO_838 (O_838,N_14781,N_14829);
nor UO_839 (O_839,N_14828,N_14980);
and UO_840 (O_840,N_14923,N_14792);
xnor UO_841 (O_841,N_14928,N_14861);
nand UO_842 (O_842,N_14849,N_14932);
or UO_843 (O_843,N_14912,N_14789);
and UO_844 (O_844,N_14839,N_14954);
xor UO_845 (O_845,N_14810,N_14881);
and UO_846 (O_846,N_14881,N_14992);
xnor UO_847 (O_847,N_14975,N_14970);
xor UO_848 (O_848,N_14980,N_14790);
nor UO_849 (O_849,N_14956,N_14931);
or UO_850 (O_850,N_14853,N_14956);
xnor UO_851 (O_851,N_14883,N_14978);
nor UO_852 (O_852,N_14830,N_14785);
xnor UO_853 (O_853,N_14937,N_14817);
and UO_854 (O_854,N_14804,N_14884);
xor UO_855 (O_855,N_14948,N_14807);
nor UO_856 (O_856,N_14939,N_14990);
or UO_857 (O_857,N_14882,N_14941);
nor UO_858 (O_858,N_14785,N_14995);
nand UO_859 (O_859,N_14934,N_14994);
xor UO_860 (O_860,N_14837,N_14908);
nor UO_861 (O_861,N_14896,N_14846);
xnor UO_862 (O_862,N_14933,N_14966);
nand UO_863 (O_863,N_14897,N_14787);
nor UO_864 (O_864,N_14824,N_14829);
or UO_865 (O_865,N_14900,N_14753);
or UO_866 (O_866,N_14874,N_14809);
nand UO_867 (O_867,N_14981,N_14952);
nand UO_868 (O_868,N_14861,N_14797);
nor UO_869 (O_869,N_14794,N_14958);
nor UO_870 (O_870,N_14881,N_14937);
or UO_871 (O_871,N_14930,N_14807);
nor UO_872 (O_872,N_14810,N_14802);
or UO_873 (O_873,N_14828,N_14861);
nor UO_874 (O_874,N_14786,N_14998);
nand UO_875 (O_875,N_14914,N_14883);
xor UO_876 (O_876,N_14762,N_14923);
and UO_877 (O_877,N_14820,N_14934);
nand UO_878 (O_878,N_14814,N_14869);
or UO_879 (O_879,N_14991,N_14770);
nand UO_880 (O_880,N_14783,N_14814);
and UO_881 (O_881,N_14857,N_14986);
xor UO_882 (O_882,N_14945,N_14893);
and UO_883 (O_883,N_14862,N_14951);
or UO_884 (O_884,N_14938,N_14962);
nor UO_885 (O_885,N_14770,N_14914);
nand UO_886 (O_886,N_14946,N_14963);
xor UO_887 (O_887,N_14835,N_14788);
nor UO_888 (O_888,N_14825,N_14975);
xnor UO_889 (O_889,N_14930,N_14986);
or UO_890 (O_890,N_14820,N_14780);
xnor UO_891 (O_891,N_14966,N_14873);
nand UO_892 (O_892,N_14839,N_14834);
nand UO_893 (O_893,N_14971,N_14883);
or UO_894 (O_894,N_14985,N_14807);
xor UO_895 (O_895,N_14756,N_14982);
and UO_896 (O_896,N_14823,N_14791);
and UO_897 (O_897,N_14832,N_14755);
nor UO_898 (O_898,N_14783,N_14856);
nor UO_899 (O_899,N_14822,N_14791);
nand UO_900 (O_900,N_14887,N_14835);
or UO_901 (O_901,N_14792,N_14861);
or UO_902 (O_902,N_14933,N_14953);
and UO_903 (O_903,N_14976,N_14890);
or UO_904 (O_904,N_14977,N_14952);
and UO_905 (O_905,N_14913,N_14908);
or UO_906 (O_906,N_14760,N_14903);
nor UO_907 (O_907,N_14789,N_14785);
nor UO_908 (O_908,N_14950,N_14834);
nand UO_909 (O_909,N_14987,N_14935);
xnor UO_910 (O_910,N_14776,N_14898);
and UO_911 (O_911,N_14782,N_14967);
nor UO_912 (O_912,N_14902,N_14760);
nand UO_913 (O_913,N_14921,N_14855);
nor UO_914 (O_914,N_14883,N_14895);
xnor UO_915 (O_915,N_14844,N_14905);
or UO_916 (O_916,N_14765,N_14892);
xnor UO_917 (O_917,N_14815,N_14797);
nand UO_918 (O_918,N_14989,N_14967);
nand UO_919 (O_919,N_14954,N_14807);
or UO_920 (O_920,N_14997,N_14860);
and UO_921 (O_921,N_14878,N_14970);
nand UO_922 (O_922,N_14851,N_14931);
and UO_923 (O_923,N_14857,N_14883);
xor UO_924 (O_924,N_14957,N_14951);
nor UO_925 (O_925,N_14926,N_14933);
nor UO_926 (O_926,N_14832,N_14941);
or UO_927 (O_927,N_14753,N_14790);
and UO_928 (O_928,N_14772,N_14990);
and UO_929 (O_929,N_14941,N_14754);
xnor UO_930 (O_930,N_14882,N_14809);
nand UO_931 (O_931,N_14833,N_14928);
and UO_932 (O_932,N_14813,N_14820);
nor UO_933 (O_933,N_14986,N_14886);
nand UO_934 (O_934,N_14839,N_14849);
and UO_935 (O_935,N_14823,N_14923);
xor UO_936 (O_936,N_14980,N_14954);
xor UO_937 (O_937,N_14800,N_14941);
nand UO_938 (O_938,N_14821,N_14880);
nor UO_939 (O_939,N_14919,N_14930);
and UO_940 (O_940,N_14991,N_14819);
or UO_941 (O_941,N_14759,N_14928);
xnor UO_942 (O_942,N_14829,N_14766);
nand UO_943 (O_943,N_14824,N_14875);
and UO_944 (O_944,N_14863,N_14934);
xor UO_945 (O_945,N_14916,N_14878);
or UO_946 (O_946,N_14951,N_14882);
xor UO_947 (O_947,N_14907,N_14833);
nor UO_948 (O_948,N_14941,N_14962);
and UO_949 (O_949,N_14787,N_14895);
and UO_950 (O_950,N_14849,N_14903);
nand UO_951 (O_951,N_14787,N_14795);
xnor UO_952 (O_952,N_14904,N_14890);
and UO_953 (O_953,N_14983,N_14973);
nor UO_954 (O_954,N_14976,N_14887);
nand UO_955 (O_955,N_14824,N_14797);
and UO_956 (O_956,N_14888,N_14864);
nor UO_957 (O_957,N_14946,N_14750);
nor UO_958 (O_958,N_14834,N_14824);
or UO_959 (O_959,N_14851,N_14786);
and UO_960 (O_960,N_14921,N_14810);
and UO_961 (O_961,N_14982,N_14993);
nor UO_962 (O_962,N_14770,N_14901);
xnor UO_963 (O_963,N_14940,N_14997);
or UO_964 (O_964,N_14893,N_14751);
xnor UO_965 (O_965,N_14793,N_14822);
and UO_966 (O_966,N_14841,N_14939);
nand UO_967 (O_967,N_14998,N_14956);
or UO_968 (O_968,N_14750,N_14978);
xnor UO_969 (O_969,N_14931,N_14903);
xor UO_970 (O_970,N_14864,N_14980);
and UO_971 (O_971,N_14942,N_14788);
and UO_972 (O_972,N_14933,N_14868);
nand UO_973 (O_973,N_14861,N_14871);
and UO_974 (O_974,N_14776,N_14854);
xnor UO_975 (O_975,N_14771,N_14911);
nand UO_976 (O_976,N_14916,N_14751);
and UO_977 (O_977,N_14918,N_14782);
nor UO_978 (O_978,N_14986,N_14995);
nand UO_979 (O_979,N_14931,N_14838);
nand UO_980 (O_980,N_14856,N_14997);
nand UO_981 (O_981,N_14789,N_14795);
nor UO_982 (O_982,N_14954,N_14905);
nor UO_983 (O_983,N_14890,N_14932);
and UO_984 (O_984,N_14849,N_14885);
nor UO_985 (O_985,N_14777,N_14894);
or UO_986 (O_986,N_14795,N_14852);
xnor UO_987 (O_987,N_14826,N_14935);
nor UO_988 (O_988,N_14826,N_14971);
or UO_989 (O_989,N_14894,N_14971);
nand UO_990 (O_990,N_14824,N_14756);
nand UO_991 (O_991,N_14940,N_14791);
xor UO_992 (O_992,N_14838,N_14789);
or UO_993 (O_993,N_14992,N_14998);
and UO_994 (O_994,N_14975,N_14774);
xnor UO_995 (O_995,N_14952,N_14992);
and UO_996 (O_996,N_14864,N_14756);
xnor UO_997 (O_997,N_14932,N_14912);
nor UO_998 (O_998,N_14786,N_14755);
nand UO_999 (O_999,N_14959,N_14786);
nor UO_1000 (O_1000,N_14786,N_14833);
nor UO_1001 (O_1001,N_14800,N_14761);
nand UO_1002 (O_1002,N_14956,N_14850);
or UO_1003 (O_1003,N_14888,N_14887);
or UO_1004 (O_1004,N_14755,N_14911);
nand UO_1005 (O_1005,N_14837,N_14987);
or UO_1006 (O_1006,N_14788,N_14817);
xor UO_1007 (O_1007,N_14801,N_14985);
and UO_1008 (O_1008,N_14953,N_14823);
and UO_1009 (O_1009,N_14840,N_14880);
nand UO_1010 (O_1010,N_14769,N_14918);
nand UO_1011 (O_1011,N_14994,N_14751);
nor UO_1012 (O_1012,N_14980,N_14992);
nand UO_1013 (O_1013,N_14766,N_14913);
nand UO_1014 (O_1014,N_14925,N_14886);
or UO_1015 (O_1015,N_14757,N_14840);
or UO_1016 (O_1016,N_14799,N_14980);
nor UO_1017 (O_1017,N_14771,N_14973);
or UO_1018 (O_1018,N_14935,N_14762);
nor UO_1019 (O_1019,N_14791,N_14967);
nor UO_1020 (O_1020,N_14798,N_14991);
or UO_1021 (O_1021,N_14793,N_14862);
or UO_1022 (O_1022,N_14917,N_14915);
nor UO_1023 (O_1023,N_14810,N_14847);
and UO_1024 (O_1024,N_14775,N_14805);
or UO_1025 (O_1025,N_14840,N_14876);
and UO_1026 (O_1026,N_14863,N_14916);
xnor UO_1027 (O_1027,N_14920,N_14923);
xnor UO_1028 (O_1028,N_14874,N_14999);
xnor UO_1029 (O_1029,N_14793,N_14839);
or UO_1030 (O_1030,N_14858,N_14956);
nor UO_1031 (O_1031,N_14862,N_14931);
nand UO_1032 (O_1032,N_14948,N_14883);
nand UO_1033 (O_1033,N_14763,N_14947);
xnor UO_1034 (O_1034,N_14886,N_14944);
or UO_1035 (O_1035,N_14822,N_14927);
nor UO_1036 (O_1036,N_14948,N_14933);
nand UO_1037 (O_1037,N_14844,N_14807);
or UO_1038 (O_1038,N_14785,N_14836);
or UO_1039 (O_1039,N_14944,N_14905);
or UO_1040 (O_1040,N_14923,N_14891);
or UO_1041 (O_1041,N_14865,N_14844);
nand UO_1042 (O_1042,N_14876,N_14897);
or UO_1043 (O_1043,N_14829,N_14966);
and UO_1044 (O_1044,N_14934,N_14805);
nor UO_1045 (O_1045,N_14762,N_14782);
and UO_1046 (O_1046,N_14940,N_14930);
nand UO_1047 (O_1047,N_14759,N_14760);
nand UO_1048 (O_1048,N_14775,N_14933);
nor UO_1049 (O_1049,N_14970,N_14760);
nand UO_1050 (O_1050,N_14832,N_14809);
and UO_1051 (O_1051,N_14946,N_14826);
nand UO_1052 (O_1052,N_14871,N_14924);
nand UO_1053 (O_1053,N_14788,N_14787);
xor UO_1054 (O_1054,N_14905,N_14906);
nand UO_1055 (O_1055,N_14968,N_14810);
nand UO_1056 (O_1056,N_14943,N_14911);
xor UO_1057 (O_1057,N_14774,N_14754);
xor UO_1058 (O_1058,N_14985,N_14925);
nor UO_1059 (O_1059,N_14952,N_14895);
xnor UO_1060 (O_1060,N_14752,N_14876);
nor UO_1061 (O_1061,N_14775,N_14905);
nand UO_1062 (O_1062,N_14777,N_14797);
and UO_1063 (O_1063,N_14849,N_14864);
and UO_1064 (O_1064,N_14884,N_14985);
nand UO_1065 (O_1065,N_14951,N_14877);
xnor UO_1066 (O_1066,N_14788,N_14852);
nand UO_1067 (O_1067,N_14864,N_14833);
nor UO_1068 (O_1068,N_14828,N_14750);
nor UO_1069 (O_1069,N_14796,N_14924);
nand UO_1070 (O_1070,N_14855,N_14751);
and UO_1071 (O_1071,N_14859,N_14928);
nand UO_1072 (O_1072,N_14883,N_14796);
nor UO_1073 (O_1073,N_14893,N_14823);
nor UO_1074 (O_1074,N_14836,N_14751);
or UO_1075 (O_1075,N_14752,N_14916);
nand UO_1076 (O_1076,N_14828,N_14809);
nor UO_1077 (O_1077,N_14976,N_14985);
nand UO_1078 (O_1078,N_14962,N_14997);
nor UO_1079 (O_1079,N_14783,N_14907);
xnor UO_1080 (O_1080,N_14846,N_14961);
nor UO_1081 (O_1081,N_14874,N_14867);
and UO_1082 (O_1082,N_14795,N_14881);
or UO_1083 (O_1083,N_14816,N_14790);
or UO_1084 (O_1084,N_14868,N_14879);
xor UO_1085 (O_1085,N_14889,N_14936);
and UO_1086 (O_1086,N_14937,N_14828);
xnor UO_1087 (O_1087,N_14872,N_14884);
xor UO_1088 (O_1088,N_14928,N_14812);
nand UO_1089 (O_1089,N_14856,N_14870);
or UO_1090 (O_1090,N_14871,N_14887);
nor UO_1091 (O_1091,N_14800,N_14781);
nand UO_1092 (O_1092,N_14974,N_14864);
and UO_1093 (O_1093,N_14781,N_14951);
nor UO_1094 (O_1094,N_14778,N_14922);
nor UO_1095 (O_1095,N_14773,N_14926);
nor UO_1096 (O_1096,N_14958,N_14970);
and UO_1097 (O_1097,N_14757,N_14802);
nand UO_1098 (O_1098,N_14949,N_14856);
nand UO_1099 (O_1099,N_14874,N_14783);
or UO_1100 (O_1100,N_14813,N_14878);
xnor UO_1101 (O_1101,N_14969,N_14852);
or UO_1102 (O_1102,N_14900,N_14854);
and UO_1103 (O_1103,N_14857,N_14899);
nor UO_1104 (O_1104,N_14841,N_14826);
and UO_1105 (O_1105,N_14944,N_14989);
or UO_1106 (O_1106,N_14935,N_14962);
or UO_1107 (O_1107,N_14890,N_14992);
and UO_1108 (O_1108,N_14894,N_14875);
or UO_1109 (O_1109,N_14823,N_14772);
nor UO_1110 (O_1110,N_14859,N_14802);
or UO_1111 (O_1111,N_14841,N_14914);
and UO_1112 (O_1112,N_14882,N_14807);
xor UO_1113 (O_1113,N_14978,N_14887);
and UO_1114 (O_1114,N_14955,N_14765);
nor UO_1115 (O_1115,N_14831,N_14813);
xor UO_1116 (O_1116,N_14822,N_14919);
or UO_1117 (O_1117,N_14893,N_14918);
nor UO_1118 (O_1118,N_14998,N_14984);
and UO_1119 (O_1119,N_14918,N_14771);
or UO_1120 (O_1120,N_14769,N_14952);
nand UO_1121 (O_1121,N_14923,N_14892);
nor UO_1122 (O_1122,N_14893,N_14852);
or UO_1123 (O_1123,N_14795,N_14826);
nor UO_1124 (O_1124,N_14807,N_14906);
xnor UO_1125 (O_1125,N_14796,N_14988);
nand UO_1126 (O_1126,N_14873,N_14992);
xnor UO_1127 (O_1127,N_14770,N_14812);
xnor UO_1128 (O_1128,N_14773,N_14893);
xor UO_1129 (O_1129,N_14774,N_14934);
or UO_1130 (O_1130,N_14903,N_14864);
nand UO_1131 (O_1131,N_14755,N_14802);
nand UO_1132 (O_1132,N_14859,N_14861);
and UO_1133 (O_1133,N_14909,N_14827);
nor UO_1134 (O_1134,N_14890,N_14993);
and UO_1135 (O_1135,N_14939,N_14846);
and UO_1136 (O_1136,N_14935,N_14910);
nor UO_1137 (O_1137,N_14985,N_14759);
or UO_1138 (O_1138,N_14839,N_14791);
nor UO_1139 (O_1139,N_14776,N_14766);
or UO_1140 (O_1140,N_14979,N_14905);
or UO_1141 (O_1141,N_14810,N_14824);
nand UO_1142 (O_1142,N_14789,N_14814);
nor UO_1143 (O_1143,N_14999,N_14879);
and UO_1144 (O_1144,N_14791,N_14818);
or UO_1145 (O_1145,N_14910,N_14866);
or UO_1146 (O_1146,N_14867,N_14912);
xnor UO_1147 (O_1147,N_14955,N_14974);
nor UO_1148 (O_1148,N_14972,N_14823);
nand UO_1149 (O_1149,N_14960,N_14954);
xnor UO_1150 (O_1150,N_14778,N_14891);
nor UO_1151 (O_1151,N_14993,N_14770);
nand UO_1152 (O_1152,N_14974,N_14887);
or UO_1153 (O_1153,N_14855,N_14976);
nand UO_1154 (O_1154,N_14792,N_14912);
nand UO_1155 (O_1155,N_14829,N_14778);
or UO_1156 (O_1156,N_14891,N_14849);
nor UO_1157 (O_1157,N_14976,N_14864);
xor UO_1158 (O_1158,N_14796,N_14917);
nand UO_1159 (O_1159,N_14988,N_14880);
and UO_1160 (O_1160,N_14969,N_14793);
xnor UO_1161 (O_1161,N_14991,N_14964);
and UO_1162 (O_1162,N_14832,N_14784);
or UO_1163 (O_1163,N_14948,N_14984);
nor UO_1164 (O_1164,N_14886,N_14843);
and UO_1165 (O_1165,N_14798,N_14821);
and UO_1166 (O_1166,N_14798,N_14886);
nand UO_1167 (O_1167,N_14781,N_14773);
nor UO_1168 (O_1168,N_14794,N_14968);
or UO_1169 (O_1169,N_14791,N_14992);
xor UO_1170 (O_1170,N_14776,N_14791);
xor UO_1171 (O_1171,N_14988,N_14834);
and UO_1172 (O_1172,N_14992,N_14939);
nor UO_1173 (O_1173,N_14801,N_14766);
or UO_1174 (O_1174,N_14828,N_14791);
xor UO_1175 (O_1175,N_14974,N_14966);
nor UO_1176 (O_1176,N_14893,N_14924);
or UO_1177 (O_1177,N_14932,N_14986);
nor UO_1178 (O_1178,N_14932,N_14978);
nor UO_1179 (O_1179,N_14986,N_14900);
nand UO_1180 (O_1180,N_14981,N_14976);
and UO_1181 (O_1181,N_14844,N_14964);
xnor UO_1182 (O_1182,N_14822,N_14847);
nand UO_1183 (O_1183,N_14791,N_14912);
and UO_1184 (O_1184,N_14766,N_14920);
and UO_1185 (O_1185,N_14805,N_14932);
and UO_1186 (O_1186,N_14898,N_14829);
nand UO_1187 (O_1187,N_14803,N_14751);
nor UO_1188 (O_1188,N_14786,N_14787);
xnor UO_1189 (O_1189,N_14873,N_14958);
and UO_1190 (O_1190,N_14966,N_14899);
nand UO_1191 (O_1191,N_14804,N_14775);
and UO_1192 (O_1192,N_14845,N_14750);
xnor UO_1193 (O_1193,N_14928,N_14992);
and UO_1194 (O_1194,N_14856,N_14872);
and UO_1195 (O_1195,N_14900,N_14750);
nor UO_1196 (O_1196,N_14952,N_14896);
and UO_1197 (O_1197,N_14842,N_14804);
nor UO_1198 (O_1198,N_14913,N_14888);
or UO_1199 (O_1199,N_14944,N_14843);
and UO_1200 (O_1200,N_14813,N_14947);
nand UO_1201 (O_1201,N_14994,N_14900);
or UO_1202 (O_1202,N_14989,N_14927);
xnor UO_1203 (O_1203,N_14955,N_14851);
xnor UO_1204 (O_1204,N_14877,N_14994);
nand UO_1205 (O_1205,N_14777,N_14888);
nor UO_1206 (O_1206,N_14795,N_14966);
nor UO_1207 (O_1207,N_14998,N_14808);
nand UO_1208 (O_1208,N_14979,N_14771);
xor UO_1209 (O_1209,N_14822,N_14757);
nor UO_1210 (O_1210,N_14781,N_14978);
or UO_1211 (O_1211,N_14913,N_14912);
or UO_1212 (O_1212,N_14911,N_14867);
and UO_1213 (O_1213,N_14949,N_14971);
and UO_1214 (O_1214,N_14897,N_14985);
and UO_1215 (O_1215,N_14929,N_14973);
nor UO_1216 (O_1216,N_14876,N_14917);
nor UO_1217 (O_1217,N_14977,N_14791);
or UO_1218 (O_1218,N_14988,N_14992);
nand UO_1219 (O_1219,N_14996,N_14958);
xor UO_1220 (O_1220,N_14784,N_14891);
nand UO_1221 (O_1221,N_14753,N_14843);
and UO_1222 (O_1222,N_14803,N_14847);
or UO_1223 (O_1223,N_14763,N_14751);
or UO_1224 (O_1224,N_14890,N_14834);
nand UO_1225 (O_1225,N_14768,N_14894);
xnor UO_1226 (O_1226,N_14865,N_14980);
or UO_1227 (O_1227,N_14809,N_14969);
nand UO_1228 (O_1228,N_14809,N_14994);
xnor UO_1229 (O_1229,N_14895,N_14973);
nor UO_1230 (O_1230,N_14873,N_14807);
xnor UO_1231 (O_1231,N_14898,N_14885);
nor UO_1232 (O_1232,N_14839,N_14858);
and UO_1233 (O_1233,N_14831,N_14994);
nand UO_1234 (O_1234,N_14832,N_14948);
or UO_1235 (O_1235,N_14867,N_14792);
xnor UO_1236 (O_1236,N_14971,N_14948);
nor UO_1237 (O_1237,N_14784,N_14796);
and UO_1238 (O_1238,N_14910,N_14776);
nand UO_1239 (O_1239,N_14897,N_14829);
nand UO_1240 (O_1240,N_14795,N_14953);
and UO_1241 (O_1241,N_14957,N_14983);
nand UO_1242 (O_1242,N_14821,N_14771);
or UO_1243 (O_1243,N_14807,N_14829);
or UO_1244 (O_1244,N_14875,N_14838);
or UO_1245 (O_1245,N_14879,N_14765);
nand UO_1246 (O_1246,N_14799,N_14899);
xnor UO_1247 (O_1247,N_14951,N_14937);
nand UO_1248 (O_1248,N_14960,N_14760);
xnor UO_1249 (O_1249,N_14872,N_14930);
xnor UO_1250 (O_1250,N_14810,N_14755);
xor UO_1251 (O_1251,N_14894,N_14885);
nand UO_1252 (O_1252,N_14826,N_14965);
xnor UO_1253 (O_1253,N_14819,N_14907);
xor UO_1254 (O_1254,N_14844,N_14925);
and UO_1255 (O_1255,N_14772,N_14767);
or UO_1256 (O_1256,N_14760,N_14804);
xor UO_1257 (O_1257,N_14830,N_14845);
or UO_1258 (O_1258,N_14923,N_14921);
xor UO_1259 (O_1259,N_14998,N_14851);
nand UO_1260 (O_1260,N_14927,N_14996);
and UO_1261 (O_1261,N_14983,N_14830);
or UO_1262 (O_1262,N_14824,N_14750);
nor UO_1263 (O_1263,N_14836,N_14956);
xnor UO_1264 (O_1264,N_14765,N_14911);
nor UO_1265 (O_1265,N_14791,N_14870);
xnor UO_1266 (O_1266,N_14953,N_14980);
xnor UO_1267 (O_1267,N_14822,N_14871);
xor UO_1268 (O_1268,N_14752,N_14962);
nor UO_1269 (O_1269,N_14924,N_14797);
or UO_1270 (O_1270,N_14876,N_14894);
nand UO_1271 (O_1271,N_14880,N_14817);
nor UO_1272 (O_1272,N_14756,N_14809);
xnor UO_1273 (O_1273,N_14812,N_14955);
nor UO_1274 (O_1274,N_14963,N_14800);
or UO_1275 (O_1275,N_14876,N_14990);
and UO_1276 (O_1276,N_14773,N_14819);
nand UO_1277 (O_1277,N_14813,N_14990);
nor UO_1278 (O_1278,N_14972,N_14915);
and UO_1279 (O_1279,N_14793,N_14947);
xor UO_1280 (O_1280,N_14881,N_14759);
and UO_1281 (O_1281,N_14974,N_14936);
and UO_1282 (O_1282,N_14926,N_14911);
nor UO_1283 (O_1283,N_14993,N_14808);
or UO_1284 (O_1284,N_14976,N_14964);
or UO_1285 (O_1285,N_14996,N_14865);
nor UO_1286 (O_1286,N_14903,N_14790);
or UO_1287 (O_1287,N_14967,N_14850);
xnor UO_1288 (O_1288,N_14939,N_14884);
and UO_1289 (O_1289,N_14999,N_14842);
nor UO_1290 (O_1290,N_14770,N_14776);
and UO_1291 (O_1291,N_14885,N_14862);
nor UO_1292 (O_1292,N_14785,N_14987);
nor UO_1293 (O_1293,N_14913,N_14952);
or UO_1294 (O_1294,N_14806,N_14912);
xor UO_1295 (O_1295,N_14775,N_14951);
nand UO_1296 (O_1296,N_14788,N_14855);
and UO_1297 (O_1297,N_14947,N_14824);
xor UO_1298 (O_1298,N_14930,N_14766);
and UO_1299 (O_1299,N_14957,N_14914);
nand UO_1300 (O_1300,N_14901,N_14872);
or UO_1301 (O_1301,N_14929,N_14987);
and UO_1302 (O_1302,N_14861,N_14802);
xor UO_1303 (O_1303,N_14978,N_14943);
xnor UO_1304 (O_1304,N_14845,N_14909);
or UO_1305 (O_1305,N_14760,N_14823);
xor UO_1306 (O_1306,N_14760,N_14772);
nand UO_1307 (O_1307,N_14876,N_14916);
nand UO_1308 (O_1308,N_14941,N_14938);
xor UO_1309 (O_1309,N_14876,N_14925);
nor UO_1310 (O_1310,N_14983,N_14917);
and UO_1311 (O_1311,N_14766,N_14782);
nor UO_1312 (O_1312,N_14781,N_14780);
and UO_1313 (O_1313,N_14803,N_14943);
or UO_1314 (O_1314,N_14918,N_14948);
xor UO_1315 (O_1315,N_14920,N_14882);
xnor UO_1316 (O_1316,N_14930,N_14756);
nand UO_1317 (O_1317,N_14818,N_14953);
nor UO_1318 (O_1318,N_14960,N_14852);
or UO_1319 (O_1319,N_14782,N_14911);
or UO_1320 (O_1320,N_14907,N_14986);
nand UO_1321 (O_1321,N_14791,N_14866);
nor UO_1322 (O_1322,N_14758,N_14841);
nor UO_1323 (O_1323,N_14986,N_14788);
nand UO_1324 (O_1324,N_14767,N_14843);
and UO_1325 (O_1325,N_14773,N_14821);
nor UO_1326 (O_1326,N_14961,N_14821);
nor UO_1327 (O_1327,N_14758,N_14750);
xnor UO_1328 (O_1328,N_14990,N_14967);
nand UO_1329 (O_1329,N_14992,N_14895);
and UO_1330 (O_1330,N_14913,N_14914);
nand UO_1331 (O_1331,N_14991,N_14940);
xor UO_1332 (O_1332,N_14834,N_14924);
nor UO_1333 (O_1333,N_14996,N_14810);
and UO_1334 (O_1334,N_14818,N_14966);
nor UO_1335 (O_1335,N_14863,N_14801);
nand UO_1336 (O_1336,N_14878,N_14945);
xor UO_1337 (O_1337,N_14909,N_14783);
or UO_1338 (O_1338,N_14769,N_14763);
and UO_1339 (O_1339,N_14883,N_14806);
and UO_1340 (O_1340,N_14797,N_14931);
xnor UO_1341 (O_1341,N_14810,N_14859);
nor UO_1342 (O_1342,N_14820,N_14981);
xnor UO_1343 (O_1343,N_14814,N_14881);
nor UO_1344 (O_1344,N_14885,N_14829);
and UO_1345 (O_1345,N_14955,N_14959);
xor UO_1346 (O_1346,N_14907,N_14850);
or UO_1347 (O_1347,N_14920,N_14981);
nand UO_1348 (O_1348,N_14777,N_14947);
nand UO_1349 (O_1349,N_14779,N_14932);
and UO_1350 (O_1350,N_14994,N_14785);
nand UO_1351 (O_1351,N_14774,N_14802);
or UO_1352 (O_1352,N_14832,N_14760);
nor UO_1353 (O_1353,N_14885,N_14903);
nand UO_1354 (O_1354,N_14797,N_14963);
nor UO_1355 (O_1355,N_14846,N_14864);
nand UO_1356 (O_1356,N_14773,N_14770);
or UO_1357 (O_1357,N_14831,N_14967);
xnor UO_1358 (O_1358,N_14915,N_14997);
nor UO_1359 (O_1359,N_14760,N_14835);
or UO_1360 (O_1360,N_14756,N_14918);
and UO_1361 (O_1361,N_14850,N_14781);
nand UO_1362 (O_1362,N_14894,N_14783);
nand UO_1363 (O_1363,N_14964,N_14860);
nand UO_1364 (O_1364,N_14838,N_14810);
nor UO_1365 (O_1365,N_14986,N_14993);
nand UO_1366 (O_1366,N_14866,N_14802);
xor UO_1367 (O_1367,N_14891,N_14941);
nor UO_1368 (O_1368,N_14998,N_14795);
nor UO_1369 (O_1369,N_14810,N_14914);
xnor UO_1370 (O_1370,N_14840,N_14787);
and UO_1371 (O_1371,N_14921,N_14840);
and UO_1372 (O_1372,N_14914,N_14876);
or UO_1373 (O_1373,N_14918,N_14991);
nand UO_1374 (O_1374,N_14815,N_14991);
nor UO_1375 (O_1375,N_14840,N_14805);
or UO_1376 (O_1376,N_14852,N_14940);
or UO_1377 (O_1377,N_14789,N_14856);
xor UO_1378 (O_1378,N_14912,N_14931);
xnor UO_1379 (O_1379,N_14845,N_14775);
and UO_1380 (O_1380,N_14906,N_14912);
nor UO_1381 (O_1381,N_14922,N_14832);
and UO_1382 (O_1382,N_14916,N_14755);
nor UO_1383 (O_1383,N_14866,N_14902);
or UO_1384 (O_1384,N_14889,N_14824);
and UO_1385 (O_1385,N_14993,N_14917);
or UO_1386 (O_1386,N_14778,N_14955);
and UO_1387 (O_1387,N_14977,N_14753);
and UO_1388 (O_1388,N_14895,N_14754);
nand UO_1389 (O_1389,N_14763,N_14924);
or UO_1390 (O_1390,N_14782,N_14790);
nor UO_1391 (O_1391,N_14847,N_14768);
nand UO_1392 (O_1392,N_14874,N_14831);
or UO_1393 (O_1393,N_14846,N_14875);
or UO_1394 (O_1394,N_14966,N_14797);
xor UO_1395 (O_1395,N_14940,N_14835);
nand UO_1396 (O_1396,N_14932,N_14806);
and UO_1397 (O_1397,N_14955,N_14753);
and UO_1398 (O_1398,N_14923,N_14784);
xor UO_1399 (O_1399,N_14873,N_14883);
xor UO_1400 (O_1400,N_14929,N_14813);
or UO_1401 (O_1401,N_14836,N_14822);
or UO_1402 (O_1402,N_14754,N_14909);
and UO_1403 (O_1403,N_14927,N_14994);
and UO_1404 (O_1404,N_14814,N_14793);
nand UO_1405 (O_1405,N_14761,N_14750);
nor UO_1406 (O_1406,N_14899,N_14765);
nand UO_1407 (O_1407,N_14910,N_14849);
nand UO_1408 (O_1408,N_14955,N_14956);
nand UO_1409 (O_1409,N_14752,N_14898);
and UO_1410 (O_1410,N_14905,N_14878);
xor UO_1411 (O_1411,N_14811,N_14840);
nand UO_1412 (O_1412,N_14929,N_14821);
or UO_1413 (O_1413,N_14795,N_14964);
xor UO_1414 (O_1414,N_14971,N_14780);
nor UO_1415 (O_1415,N_14828,N_14844);
and UO_1416 (O_1416,N_14973,N_14855);
and UO_1417 (O_1417,N_14752,N_14991);
nand UO_1418 (O_1418,N_14907,N_14911);
xnor UO_1419 (O_1419,N_14784,N_14771);
or UO_1420 (O_1420,N_14834,N_14910);
nand UO_1421 (O_1421,N_14904,N_14900);
or UO_1422 (O_1422,N_14757,N_14903);
nor UO_1423 (O_1423,N_14934,N_14797);
xnor UO_1424 (O_1424,N_14962,N_14841);
or UO_1425 (O_1425,N_14957,N_14835);
and UO_1426 (O_1426,N_14768,N_14995);
or UO_1427 (O_1427,N_14976,N_14853);
or UO_1428 (O_1428,N_14855,N_14818);
xor UO_1429 (O_1429,N_14934,N_14793);
and UO_1430 (O_1430,N_14971,N_14897);
nand UO_1431 (O_1431,N_14857,N_14828);
nand UO_1432 (O_1432,N_14939,N_14917);
nor UO_1433 (O_1433,N_14931,N_14927);
xnor UO_1434 (O_1434,N_14776,N_14998);
xnor UO_1435 (O_1435,N_14921,N_14783);
nand UO_1436 (O_1436,N_14796,N_14751);
nand UO_1437 (O_1437,N_14963,N_14995);
xnor UO_1438 (O_1438,N_14814,N_14886);
xor UO_1439 (O_1439,N_14879,N_14906);
and UO_1440 (O_1440,N_14976,N_14817);
or UO_1441 (O_1441,N_14879,N_14880);
or UO_1442 (O_1442,N_14867,N_14891);
and UO_1443 (O_1443,N_14898,N_14969);
and UO_1444 (O_1444,N_14807,N_14945);
or UO_1445 (O_1445,N_14817,N_14975);
nand UO_1446 (O_1446,N_14759,N_14790);
nand UO_1447 (O_1447,N_14927,N_14778);
nand UO_1448 (O_1448,N_14751,N_14960);
nor UO_1449 (O_1449,N_14924,N_14849);
xor UO_1450 (O_1450,N_14941,N_14920);
and UO_1451 (O_1451,N_14986,N_14814);
or UO_1452 (O_1452,N_14838,N_14894);
nor UO_1453 (O_1453,N_14854,N_14907);
xor UO_1454 (O_1454,N_14762,N_14942);
and UO_1455 (O_1455,N_14816,N_14807);
nand UO_1456 (O_1456,N_14831,N_14807);
nor UO_1457 (O_1457,N_14942,N_14984);
nor UO_1458 (O_1458,N_14859,N_14758);
xnor UO_1459 (O_1459,N_14932,N_14808);
and UO_1460 (O_1460,N_14784,N_14982);
nand UO_1461 (O_1461,N_14898,N_14986);
nor UO_1462 (O_1462,N_14821,N_14994);
and UO_1463 (O_1463,N_14819,N_14975);
xor UO_1464 (O_1464,N_14847,N_14917);
or UO_1465 (O_1465,N_14869,N_14820);
xor UO_1466 (O_1466,N_14853,N_14839);
or UO_1467 (O_1467,N_14982,N_14997);
nand UO_1468 (O_1468,N_14899,N_14980);
nor UO_1469 (O_1469,N_14992,N_14937);
xor UO_1470 (O_1470,N_14779,N_14894);
nand UO_1471 (O_1471,N_14978,N_14939);
or UO_1472 (O_1472,N_14972,N_14921);
or UO_1473 (O_1473,N_14966,N_14970);
xor UO_1474 (O_1474,N_14828,N_14829);
xor UO_1475 (O_1475,N_14991,N_14808);
nand UO_1476 (O_1476,N_14908,N_14993);
nand UO_1477 (O_1477,N_14966,N_14976);
nand UO_1478 (O_1478,N_14880,N_14906);
xnor UO_1479 (O_1479,N_14784,N_14858);
xor UO_1480 (O_1480,N_14866,N_14879);
nand UO_1481 (O_1481,N_14820,N_14936);
or UO_1482 (O_1482,N_14833,N_14794);
or UO_1483 (O_1483,N_14963,N_14829);
xor UO_1484 (O_1484,N_14873,N_14877);
xor UO_1485 (O_1485,N_14909,N_14907);
nand UO_1486 (O_1486,N_14816,N_14979);
or UO_1487 (O_1487,N_14884,N_14778);
xor UO_1488 (O_1488,N_14812,N_14827);
xor UO_1489 (O_1489,N_14975,N_14971);
nand UO_1490 (O_1490,N_14845,N_14802);
nor UO_1491 (O_1491,N_14964,N_14775);
nand UO_1492 (O_1492,N_14954,N_14913);
xor UO_1493 (O_1493,N_14824,N_14893);
nand UO_1494 (O_1494,N_14903,N_14816);
nor UO_1495 (O_1495,N_14752,N_14953);
nand UO_1496 (O_1496,N_14819,N_14900);
or UO_1497 (O_1497,N_14824,N_14765);
or UO_1498 (O_1498,N_14924,N_14992);
xor UO_1499 (O_1499,N_14905,N_14824);
and UO_1500 (O_1500,N_14969,N_14872);
nor UO_1501 (O_1501,N_14775,N_14795);
nor UO_1502 (O_1502,N_14942,N_14982);
xnor UO_1503 (O_1503,N_14975,N_14761);
nand UO_1504 (O_1504,N_14836,N_14798);
or UO_1505 (O_1505,N_14822,N_14885);
or UO_1506 (O_1506,N_14998,N_14962);
nand UO_1507 (O_1507,N_14885,N_14986);
xnor UO_1508 (O_1508,N_14786,N_14865);
or UO_1509 (O_1509,N_14959,N_14965);
nor UO_1510 (O_1510,N_14785,N_14884);
and UO_1511 (O_1511,N_14905,N_14768);
or UO_1512 (O_1512,N_14967,N_14996);
and UO_1513 (O_1513,N_14787,N_14923);
xor UO_1514 (O_1514,N_14984,N_14852);
and UO_1515 (O_1515,N_14842,N_14824);
nor UO_1516 (O_1516,N_14843,N_14771);
and UO_1517 (O_1517,N_14902,N_14813);
or UO_1518 (O_1518,N_14854,N_14984);
nor UO_1519 (O_1519,N_14950,N_14851);
xnor UO_1520 (O_1520,N_14820,N_14975);
nor UO_1521 (O_1521,N_14842,N_14950);
or UO_1522 (O_1522,N_14765,N_14851);
xnor UO_1523 (O_1523,N_14994,N_14990);
nor UO_1524 (O_1524,N_14805,N_14981);
or UO_1525 (O_1525,N_14806,N_14773);
xnor UO_1526 (O_1526,N_14958,N_14945);
or UO_1527 (O_1527,N_14768,N_14860);
and UO_1528 (O_1528,N_14807,N_14865);
nor UO_1529 (O_1529,N_14850,N_14768);
xnor UO_1530 (O_1530,N_14846,N_14869);
and UO_1531 (O_1531,N_14817,N_14953);
and UO_1532 (O_1532,N_14870,N_14915);
or UO_1533 (O_1533,N_14975,N_14757);
nor UO_1534 (O_1534,N_14966,N_14798);
or UO_1535 (O_1535,N_14754,N_14975);
nand UO_1536 (O_1536,N_14815,N_14952);
nand UO_1537 (O_1537,N_14823,N_14845);
nand UO_1538 (O_1538,N_14953,N_14994);
or UO_1539 (O_1539,N_14864,N_14856);
or UO_1540 (O_1540,N_14777,N_14802);
or UO_1541 (O_1541,N_14979,N_14780);
xnor UO_1542 (O_1542,N_14784,N_14871);
xor UO_1543 (O_1543,N_14762,N_14924);
and UO_1544 (O_1544,N_14884,N_14994);
or UO_1545 (O_1545,N_14751,N_14878);
nor UO_1546 (O_1546,N_14850,N_14759);
xnor UO_1547 (O_1547,N_14777,N_14840);
xor UO_1548 (O_1548,N_14806,N_14814);
nand UO_1549 (O_1549,N_14756,N_14929);
and UO_1550 (O_1550,N_14963,N_14818);
nand UO_1551 (O_1551,N_14905,N_14919);
nor UO_1552 (O_1552,N_14934,N_14806);
and UO_1553 (O_1553,N_14778,N_14967);
nand UO_1554 (O_1554,N_14918,N_14951);
nand UO_1555 (O_1555,N_14825,N_14791);
nor UO_1556 (O_1556,N_14912,N_14954);
or UO_1557 (O_1557,N_14821,N_14910);
and UO_1558 (O_1558,N_14811,N_14777);
nor UO_1559 (O_1559,N_14764,N_14894);
or UO_1560 (O_1560,N_14934,N_14847);
xor UO_1561 (O_1561,N_14890,N_14805);
and UO_1562 (O_1562,N_14796,N_14792);
and UO_1563 (O_1563,N_14931,N_14827);
and UO_1564 (O_1564,N_14821,N_14794);
and UO_1565 (O_1565,N_14799,N_14812);
nand UO_1566 (O_1566,N_14907,N_14897);
nor UO_1567 (O_1567,N_14966,N_14917);
or UO_1568 (O_1568,N_14902,N_14824);
nand UO_1569 (O_1569,N_14755,N_14995);
nand UO_1570 (O_1570,N_14794,N_14776);
nand UO_1571 (O_1571,N_14801,N_14950);
and UO_1572 (O_1572,N_14884,N_14969);
or UO_1573 (O_1573,N_14781,N_14801);
xor UO_1574 (O_1574,N_14953,N_14996);
xor UO_1575 (O_1575,N_14994,N_14802);
and UO_1576 (O_1576,N_14913,N_14814);
nor UO_1577 (O_1577,N_14997,N_14771);
nor UO_1578 (O_1578,N_14962,N_14840);
or UO_1579 (O_1579,N_14925,N_14969);
nor UO_1580 (O_1580,N_14999,N_14823);
or UO_1581 (O_1581,N_14757,N_14796);
xnor UO_1582 (O_1582,N_14922,N_14817);
xor UO_1583 (O_1583,N_14995,N_14760);
or UO_1584 (O_1584,N_14758,N_14952);
nand UO_1585 (O_1585,N_14965,N_14761);
nand UO_1586 (O_1586,N_14997,N_14755);
nor UO_1587 (O_1587,N_14983,N_14845);
nand UO_1588 (O_1588,N_14932,N_14905);
nand UO_1589 (O_1589,N_14920,N_14916);
nand UO_1590 (O_1590,N_14978,N_14794);
xor UO_1591 (O_1591,N_14899,N_14761);
nand UO_1592 (O_1592,N_14820,N_14913);
nand UO_1593 (O_1593,N_14801,N_14887);
xor UO_1594 (O_1594,N_14800,N_14924);
nor UO_1595 (O_1595,N_14754,N_14938);
nor UO_1596 (O_1596,N_14929,N_14783);
xor UO_1597 (O_1597,N_14914,N_14818);
xor UO_1598 (O_1598,N_14836,N_14875);
and UO_1599 (O_1599,N_14808,N_14787);
or UO_1600 (O_1600,N_14824,N_14781);
and UO_1601 (O_1601,N_14973,N_14750);
nand UO_1602 (O_1602,N_14922,N_14813);
and UO_1603 (O_1603,N_14972,N_14973);
and UO_1604 (O_1604,N_14913,N_14815);
and UO_1605 (O_1605,N_14794,N_14982);
or UO_1606 (O_1606,N_14778,N_14873);
or UO_1607 (O_1607,N_14855,N_14859);
nand UO_1608 (O_1608,N_14953,N_14928);
or UO_1609 (O_1609,N_14891,N_14791);
and UO_1610 (O_1610,N_14992,N_14811);
xnor UO_1611 (O_1611,N_14836,N_14841);
and UO_1612 (O_1612,N_14937,N_14987);
xnor UO_1613 (O_1613,N_14941,N_14831);
nor UO_1614 (O_1614,N_14844,N_14800);
xnor UO_1615 (O_1615,N_14782,N_14888);
nor UO_1616 (O_1616,N_14769,N_14896);
nor UO_1617 (O_1617,N_14798,N_14806);
and UO_1618 (O_1618,N_14878,N_14933);
and UO_1619 (O_1619,N_14878,N_14975);
and UO_1620 (O_1620,N_14992,N_14763);
xor UO_1621 (O_1621,N_14988,N_14767);
and UO_1622 (O_1622,N_14827,N_14961);
and UO_1623 (O_1623,N_14860,N_14986);
and UO_1624 (O_1624,N_14817,N_14775);
nand UO_1625 (O_1625,N_14842,N_14921);
nor UO_1626 (O_1626,N_14874,N_14953);
nor UO_1627 (O_1627,N_14794,N_14915);
xnor UO_1628 (O_1628,N_14926,N_14808);
and UO_1629 (O_1629,N_14862,N_14787);
xnor UO_1630 (O_1630,N_14991,N_14807);
xnor UO_1631 (O_1631,N_14999,N_14945);
or UO_1632 (O_1632,N_14897,N_14865);
nand UO_1633 (O_1633,N_14808,N_14753);
or UO_1634 (O_1634,N_14905,N_14920);
nor UO_1635 (O_1635,N_14856,N_14994);
nor UO_1636 (O_1636,N_14955,N_14776);
nor UO_1637 (O_1637,N_14763,N_14784);
or UO_1638 (O_1638,N_14797,N_14935);
nor UO_1639 (O_1639,N_14796,N_14840);
nand UO_1640 (O_1640,N_14795,N_14804);
nor UO_1641 (O_1641,N_14885,N_14753);
nor UO_1642 (O_1642,N_14981,N_14855);
xnor UO_1643 (O_1643,N_14768,N_14957);
and UO_1644 (O_1644,N_14922,N_14750);
nor UO_1645 (O_1645,N_14942,N_14974);
and UO_1646 (O_1646,N_14831,N_14808);
nand UO_1647 (O_1647,N_14980,N_14881);
or UO_1648 (O_1648,N_14836,N_14903);
nor UO_1649 (O_1649,N_14799,N_14866);
or UO_1650 (O_1650,N_14866,N_14987);
nor UO_1651 (O_1651,N_14825,N_14933);
nand UO_1652 (O_1652,N_14857,N_14878);
or UO_1653 (O_1653,N_14950,N_14817);
nand UO_1654 (O_1654,N_14921,N_14879);
and UO_1655 (O_1655,N_14755,N_14846);
nand UO_1656 (O_1656,N_14993,N_14751);
nand UO_1657 (O_1657,N_14906,N_14991);
nand UO_1658 (O_1658,N_14816,N_14920);
nand UO_1659 (O_1659,N_14878,N_14821);
nor UO_1660 (O_1660,N_14926,N_14943);
xnor UO_1661 (O_1661,N_14937,N_14774);
nand UO_1662 (O_1662,N_14783,N_14889);
xor UO_1663 (O_1663,N_14873,N_14988);
or UO_1664 (O_1664,N_14862,N_14956);
nor UO_1665 (O_1665,N_14848,N_14829);
nand UO_1666 (O_1666,N_14820,N_14795);
xor UO_1667 (O_1667,N_14952,N_14798);
nand UO_1668 (O_1668,N_14932,N_14774);
and UO_1669 (O_1669,N_14841,N_14996);
or UO_1670 (O_1670,N_14984,N_14945);
nand UO_1671 (O_1671,N_14996,N_14895);
nor UO_1672 (O_1672,N_14902,N_14863);
and UO_1673 (O_1673,N_14942,N_14928);
and UO_1674 (O_1674,N_14768,N_14759);
nor UO_1675 (O_1675,N_14981,N_14877);
xor UO_1676 (O_1676,N_14957,N_14798);
nand UO_1677 (O_1677,N_14836,N_14986);
and UO_1678 (O_1678,N_14945,N_14788);
or UO_1679 (O_1679,N_14988,N_14966);
xnor UO_1680 (O_1680,N_14874,N_14834);
and UO_1681 (O_1681,N_14982,N_14796);
and UO_1682 (O_1682,N_14978,N_14860);
or UO_1683 (O_1683,N_14806,N_14922);
nor UO_1684 (O_1684,N_14820,N_14963);
nand UO_1685 (O_1685,N_14874,N_14824);
xor UO_1686 (O_1686,N_14764,N_14769);
nand UO_1687 (O_1687,N_14860,N_14807);
or UO_1688 (O_1688,N_14962,N_14802);
xor UO_1689 (O_1689,N_14920,N_14815);
xor UO_1690 (O_1690,N_14973,N_14799);
nand UO_1691 (O_1691,N_14797,N_14859);
xor UO_1692 (O_1692,N_14991,N_14839);
nor UO_1693 (O_1693,N_14928,N_14819);
nor UO_1694 (O_1694,N_14796,N_14825);
or UO_1695 (O_1695,N_14922,N_14921);
nand UO_1696 (O_1696,N_14983,N_14936);
or UO_1697 (O_1697,N_14970,N_14851);
or UO_1698 (O_1698,N_14992,N_14953);
or UO_1699 (O_1699,N_14845,N_14780);
or UO_1700 (O_1700,N_14862,N_14850);
nor UO_1701 (O_1701,N_14952,N_14894);
or UO_1702 (O_1702,N_14926,N_14854);
nor UO_1703 (O_1703,N_14780,N_14842);
nor UO_1704 (O_1704,N_14877,N_14776);
or UO_1705 (O_1705,N_14840,N_14964);
xnor UO_1706 (O_1706,N_14792,N_14986);
nor UO_1707 (O_1707,N_14758,N_14753);
nand UO_1708 (O_1708,N_14977,N_14766);
nor UO_1709 (O_1709,N_14961,N_14970);
or UO_1710 (O_1710,N_14936,N_14831);
or UO_1711 (O_1711,N_14796,N_14990);
and UO_1712 (O_1712,N_14883,N_14972);
nand UO_1713 (O_1713,N_14974,N_14960);
and UO_1714 (O_1714,N_14764,N_14851);
nand UO_1715 (O_1715,N_14934,N_14821);
and UO_1716 (O_1716,N_14996,N_14979);
and UO_1717 (O_1717,N_14889,N_14753);
nor UO_1718 (O_1718,N_14807,N_14758);
nand UO_1719 (O_1719,N_14840,N_14847);
and UO_1720 (O_1720,N_14762,N_14884);
nor UO_1721 (O_1721,N_14834,N_14774);
xor UO_1722 (O_1722,N_14859,N_14813);
or UO_1723 (O_1723,N_14922,N_14772);
nor UO_1724 (O_1724,N_14889,N_14772);
xnor UO_1725 (O_1725,N_14774,N_14997);
and UO_1726 (O_1726,N_14846,N_14780);
and UO_1727 (O_1727,N_14926,N_14925);
nand UO_1728 (O_1728,N_14839,N_14877);
and UO_1729 (O_1729,N_14900,N_14847);
xnor UO_1730 (O_1730,N_14895,N_14968);
nor UO_1731 (O_1731,N_14865,N_14979);
xnor UO_1732 (O_1732,N_14976,N_14984);
nor UO_1733 (O_1733,N_14953,N_14865);
or UO_1734 (O_1734,N_14980,N_14927);
nand UO_1735 (O_1735,N_14974,N_14846);
and UO_1736 (O_1736,N_14953,N_14913);
xnor UO_1737 (O_1737,N_14939,N_14967);
nor UO_1738 (O_1738,N_14906,N_14769);
nor UO_1739 (O_1739,N_14795,N_14821);
nand UO_1740 (O_1740,N_14806,N_14829);
or UO_1741 (O_1741,N_14805,N_14954);
or UO_1742 (O_1742,N_14972,N_14967);
nand UO_1743 (O_1743,N_14932,N_14820);
or UO_1744 (O_1744,N_14888,N_14857);
and UO_1745 (O_1745,N_14963,N_14874);
nor UO_1746 (O_1746,N_14799,N_14909);
xor UO_1747 (O_1747,N_14969,N_14942);
or UO_1748 (O_1748,N_14887,N_14786);
nor UO_1749 (O_1749,N_14800,N_14826);
nand UO_1750 (O_1750,N_14964,N_14959);
nand UO_1751 (O_1751,N_14941,N_14959);
and UO_1752 (O_1752,N_14775,N_14844);
or UO_1753 (O_1753,N_14760,N_14866);
xnor UO_1754 (O_1754,N_14786,N_14785);
or UO_1755 (O_1755,N_14967,N_14830);
nand UO_1756 (O_1756,N_14900,N_14873);
nor UO_1757 (O_1757,N_14918,N_14959);
and UO_1758 (O_1758,N_14786,N_14909);
or UO_1759 (O_1759,N_14858,N_14789);
nor UO_1760 (O_1760,N_14794,N_14948);
or UO_1761 (O_1761,N_14904,N_14909);
nand UO_1762 (O_1762,N_14918,N_14896);
xnor UO_1763 (O_1763,N_14776,N_14882);
nand UO_1764 (O_1764,N_14874,N_14986);
xnor UO_1765 (O_1765,N_14892,N_14814);
or UO_1766 (O_1766,N_14862,N_14939);
nor UO_1767 (O_1767,N_14776,N_14771);
xor UO_1768 (O_1768,N_14886,N_14871);
nor UO_1769 (O_1769,N_14753,N_14784);
and UO_1770 (O_1770,N_14941,N_14926);
nor UO_1771 (O_1771,N_14885,N_14918);
nand UO_1772 (O_1772,N_14777,N_14821);
nand UO_1773 (O_1773,N_14849,N_14999);
or UO_1774 (O_1774,N_14921,N_14778);
xor UO_1775 (O_1775,N_14903,N_14858);
nand UO_1776 (O_1776,N_14818,N_14971);
nor UO_1777 (O_1777,N_14798,N_14900);
nor UO_1778 (O_1778,N_14750,N_14794);
nor UO_1779 (O_1779,N_14842,N_14920);
nand UO_1780 (O_1780,N_14796,N_14865);
or UO_1781 (O_1781,N_14941,N_14797);
nor UO_1782 (O_1782,N_14892,N_14898);
nand UO_1783 (O_1783,N_14795,N_14765);
or UO_1784 (O_1784,N_14865,N_14955);
and UO_1785 (O_1785,N_14819,N_14941);
or UO_1786 (O_1786,N_14950,N_14786);
nand UO_1787 (O_1787,N_14979,N_14958);
or UO_1788 (O_1788,N_14758,N_14886);
nor UO_1789 (O_1789,N_14872,N_14773);
nor UO_1790 (O_1790,N_14999,N_14831);
nor UO_1791 (O_1791,N_14958,N_14884);
nand UO_1792 (O_1792,N_14992,N_14999);
nor UO_1793 (O_1793,N_14908,N_14797);
or UO_1794 (O_1794,N_14902,N_14959);
nand UO_1795 (O_1795,N_14993,N_14894);
nor UO_1796 (O_1796,N_14829,N_14962);
nor UO_1797 (O_1797,N_14821,N_14833);
or UO_1798 (O_1798,N_14848,N_14784);
nor UO_1799 (O_1799,N_14809,N_14785);
and UO_1800 (O_1800,N_14860,N_14790);
nand UO_1801 (O_1801,N_14867,N_14929);
xnor UO_1802 (O_1802,N_14916,N_14869);
and UO_1803 (O_1803,N_14969,N_14941);
nand UO_1804 (O_1804,N_14804,N_14964);
or UO_1805 (O_1805,N_14868,N_14839);
nor UO_1806 (O_1806,N_14753,N_14923);
xnor UO_1807 (O_1807,N_14952,N_14874);
xor UO_1808 (O_1808,N_14839,N_14777);
and UO_1809 (O_1809,N_14775,N_14797);
xnor UO_1810 (O_1810,N_14862,N_14820);
nand UO_1811 (O_1811,N_14983,N_14840);
or UO_1812 (O_1812,N_14975,N_14959);
xor UO_1813 (O_1813,N_14968,N_14856);
or UO_1814 (O_1814,N_14845,N_14814);
or UO_1815 (O_1815,N_14936,N_14801);
xnor UO_1816 (O_1816,N_14973,N_14964);
xor UO_1817 (O_1817,N_14771,N_14788);
or UO_1818 (O_1818,N_14975,N_14879);
nand UO_1819 (O_1819,N_14929,N_14925);
or UO_1820 (O_1820,N_14875,N_14804);
nor UO_1821 (O_1821,N_14967,N_14814);
nor UO_1822 (O_1822,N_14772,N_14777);
nand UO_1823 (O_1823,N_14955,N_14805);
nor UO_1824 (O_1824,N_14951,N_14831);
xor UO_1825 (O_1825,N_14970,N_14752);
nor UO_1826 (O_1826,N_14927,N_14967);
nand UO_1827 (O_1827,N_14750,N_14792);
xor UO_1828 (O_1828,N_14753,N_14765);
nand UO_1829 (O_1829,N_14835,N_14928);
and UO_1830 (O_1830,N_14973,N_14905);
nand UO_1831 (O_1831,N_14795,N_14908);
or UO_1832 (O_1832,N_14821,N_14960);
xnor UO_1833 (O_1833,N_14912,N_14869);
xor UO_1834 (O_1834,N_14970,N_14755);
nand UO_1835 (O_1835,N_14877,N_14783);
nor UO_1836 (O_1836,N_14945,N_14957);
nand UO_1837 (O_1837,N_14900,N_14870);
nor UO_1838 (O_1838,N_14829,N_14799);
or UO_1839 (O_1839,N_14977,N_14975);
nor UO_1840 (O_1840,N_14804,N_14848);
xor UO_1841 (O_1841,N_14784,N_14915);
xor UO_1842 (O_1842,N_14980,N_14957);
nor UO_1843 (O_1843,N_14899,N_14803);
nor UO_1844 (O_1844,N_14926,N_14838);
nand UO_1845 (O_1845,N_14840,N_14828);
nand UO_1846 (O_1846,N_14901,N_14991);
and UO_1847 (O_1847,N_14959,N_14946);
xor UO_1848 (O_1848,N_14844,N_14891);
or UO_1849 (O_1849,N_14849,N_14777);
nand UO_1850 (O_1850,N_14877,N_14809);
or UO_1851 (O_1851,N_14808,N_14838);
xnor UO_1852 (O_1852,N_14923,N_14938);
nand UO_1853 (O_1853,N_14759,N_14952);
and UO_1854 (O_1854,N_14801,N_14753);
and UO_1855 (O_1855,N_14914,N_14948);
and UO_1856 (O_1856,N_14802,N_14970);
xnor UO_1857 (O_1857,N_14974,N_14838);
and UO_1858 (O_1858,N_14828,N_14774);
nand UO_1859 (O_1859,N_14788,N_14827);
and UO_1860 (O_1860,N_14962,N_14773);
and UO_1861 (O_1861,N_14957,N_14827);
nor UO_1862 (O_1862,N_14790,N_14844);
nor UO_1863 (O_1863,N_14761,N_14879);
or UO_1864 (O_1864,N_14767,N_14750);
xor UO_1865 (O_1865,N_14828,N_14779);
nor UO_1866 (O_1866,N_14878,N_14799);
nand UO_1867 (O_1867,N_14827,N_14839);
or UO_1868 (O_1868,N_14954,N_14925);
and UO_1869 (O_1869,N_14865,N_14916);
xor UO_1870 (O_1870,N_14904,N_14902);
xor UO_1871 (O_1871,N_14878,N_14843);
nand UO_1872 (O_1872,N_14868,N_14875);
and UO_1873 (O_1873,N_14886,N_14775);
xnor UO_1874 (O_1874,N_14860,N_14802);
or UO_1875 (O_1875,N_14869,N_14891);
nand UO_1876 (O_1876,N_14909,N_14755);
xor UO_1877 (O_1877,N_14865,N_14794);
nor UO_1878 (O_1878,N_14942,N_14832);
and UO_1879 (O_1879,N_14800,N_14977);
and UO_1880 (O_1880,N_14902,N_14798);
or UO_1881 (O_1881,N_14905,N_14871);
nand UO_1882 (O_1882,N_14876,N_14808);
nor UO_1883 (O_1883,N_14778,N_14802);
nand UO_1884 (O_1884,N_14900,N_14876);
and UO_1885 (O_1885,N_14955,N_14941);
nand UO_1886 (O_1886,N_14831,N_14908);
nand UO_1887 (O_1887,N_14769,N_14867);
or UO_1888 (O_1888,N_14785,N_14850);
and UO_1889 (O_1889,N_14956,N_14897);
nor UO_1890 (O_1890,N_14866,N_14992);
nor UO_1891 (O_1891,N_14896,N_14797);
and UO_1892 (O_1892,N_14885,N_14995);
or UO_1893 (O_1893,N_14874,N_14910);
or UO_1894 (O_1894,N_14892,N_14778);
nor UO_1895 (O_1895,N_14895,N_14989);
nor UO_1896 (O_1896,N_14888,N_14940);
nor UO_1897 (O_1897,N_14986,N_14765);
xnor UO_1898 (O_1898,N_14965,N_14828);
or UO_1899 (O_1899,N_14752,N_14835);
or UO_1900 (O_1900,N_14946,N_14773);
or UO_1901 (O_1901,N_14841,N_14858);
or UO_1902 (O_1902,N_14919,N_14925);
or UO_1903 (O_1903,N_14997,N_14758);
nand UO_1904 (O_1904,N_14867,N_14889);
and UO_1905 (O_1905,N_14771,N_14988);
xnor UO_1906 (O_1906,N_14842,N_14872);
xor UO_1907 (O_1907,N_14848,N_14816);
and UO_1908 (O_1908,N_14984,N_14829);
nand UO_1909 (O_1909,N_14996,N_14999);
xor UO_1910 (O_1910,N_14769,N_14860);
nand UO_1911 (O_1911,N_14796,N_14970);
and UO_1912 (O_1912,N_14904,N_14794);
nand UO_1913 (O_1913,N_14771,N_14840);
or UO_1914 (O_1914,N_14889,N_14754);
xor UO_1915 (O_1915,N_14864,N_14852);
or UO_1916 (O_1916,N_14928,N_14809);
and UO_1917 (O_1917,N_14938,N_14796);
nor UO_1918 (O_1918,N_14792,N_14869);
nand UO_1919 (O_1919,N_14875,N_14879);
nand UO_1920 (O_1920,N_14996,N_14812);
nand UO_1921 (O_1921,N_14936,N_14854);
or UO_1922 (O_1922,N_14786,N_14895);
or UO_1923 (O_1923,N_14932,N_14948);
nand UO_1924 (O_1924,N_14880,N_14800);
xnor UO_1925 (O_1925,N_14909,N_14914);
xnor UO_1926 (O_1926,N_14849,N_14835);
or UO_1927 (O_1927,N_14963,N_14987);
nand UO_1928 (O_1928,N_14856,N_14800);
xor UO_1929 (O_1929,N_14776,N_14850);
nand UO_1930 (O_1930,N_14841,N_14943);
nor UO_1931 (O_1931,N_14797,N_14960);
and UO_1932 (O_1932,N_14825,N_14987);
nand UO_1933 (O_1933,N_14940,N_14822);
nand UO_1934 (O_1934,N_14767,N_14944);
or UO_1935 (O_1935,N_14882,N_14988);
xnor UO_1936 (O_1936,N_14785,N_14861);
nor UO_1937 (O_1937,N_14806,N_14769);
xor UO_1938 (O_1938,N_14915,N_14833);
or UO_1939 (O_1939,N_14963,N_14906);
or UO_1940 (O_1940,N_14888,N_14809);
nand UO_1941 (O_1941,N_14911,N_14938);
and UO_1942 (O_1942,N_14839,N_14969);
nand UO_1943 (O_1943,N_14968,N_14914);
nor UO_1944 (O_1944,N_14922,N_14781);
xnor UO_1945 (O_1945,N_14979,N_14880);
or UO_1946 (O_1946,N_14805,N_14896);
and UO_1947 (O_1947,N_14956,N_14821);
nand UO_1948 (O_1948,N_14810,N_14905);
or UO_1949 (O_1949,N_14752,N_14952);
nor UO_1950 (O_1950,N_14959,N_14967);
xnor UO_1951 (O_1951,N_14907,N_14859);
nor UO_1952 (O_1952,N_14936,N_14869);
and UO_1953 (O_1953,N_14924,N_14995);
nand UO_1954 (O_1954,N_14851,N_14814);
xnor UO_1955 (O_1955,N_14834,N_14926);
xnor UO_1956 (O_1956,N_14882,N_14886);
or UO_1957 (O_1957,N_14790,N_14788);
xnor UO_1958 (O_1958,N_14894,N_14818);
nand UO_1959 (O_1959,N_14842,N_14849);
xnor UO_1960 (O_1960,N_14950,N_14865);
or UO_1961 (O_1961,N_14942,N_14812);
nand UO_1962 (O_1962,N_14766,N_14891);
and UO_1963 (O_1963,N_14981,N_14969);
nor UO_1964 (O_1964,N_14915,N_14885);
nand UO_1965 (O_1965,N_14908,N_14987);
or UO_1966 (O_1966,N_14850,N_14889);
nand UO_1967 (O_1967,N_14752,N_14768);
nand UO_1968 (O_1968,N_14920,N_14808);
nor UO_1969 (O_1969,N_14985,N_14895);
xor UO_1970 (O_1970,N_14966,N_14983);
nor UO_1971 (O_1971,N_14899,N_14909);
or UO_1972 (O_1972,N_14987,N_14862);
and UO_1973 (O_1973,N_14832,N_14823);
nand UO_1974 (O_1974,N_14897,N_14845);
and UO_1975 (O_1975,N_14873,N_14941);
xnor UO_1976 (O_1976,N_14985,N_14908);
xnor UO_1977 (O_1977,N_14989,N_14900);
or UO_1978 (O_1978,N_14932,N_14812);
nor UO_1979 (O_1979,N_14854,N_14959);
nor UO_1980 (O_1980,N_14757,N_14773);
nand UO_1981 (O_1981,N_14912,N_14988);
xor UO_1982 (O_1982,N_14844,N_14785);
or UO_1983 (O_1983,N_14956,N_14967);
nand UO_1984 (O_1984,N_14958,N_14759);
and UO_1985 (O_1985,N_14863,N_14791);
or UO_1986 (O_1986,N_14975,N_14874);
or UO_1987 (O_1987,N_14869,N_14823);
xor UO_1988 (O_1988,N_14931,N_14898);
or UO_1989 (O_1989,N_14785,N_14813);
nand UO_1990 (O_1990,N_14924,N_14751);
nand UO_1991 (O_1991,N_14914,N_14777);
and UO_1992 (O_1992,N_14942,N_14805);
or UO_1993 (O_1993,N_14798,N_14787);
nor UO_1994 (O_1994,N_14803,N_14940);
xor UO_1995 (O_1995,N_14925,N_14910);
and UO_1996 (O_1996,N_14808,N_14834);
and UO_1997 (O_1997,N_14883,N_14921);
xor UO_1998 (O_1998,N_14751,N_14882);
xor UO_1999 (O_1999,N_14960,N_14825);
endmodule