module basic_1000_10000_1500_5_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_429,In_684);
nand U1 (N_1,In_352,In_765);
or U2 (N_2,In_496,In_308);
xor U3 (N_3,In_115,In_87);
and U4 (N_4,In_390,In_17);
nor U5 (N_5,In_416,In_111);
and U6 (N_6,In_642,In_340);
and U7 (N_7,In_224,In_967);
or U8 (N_8,In_217,In_623);
or U9 (N_9,In_43,In_332);
nand U10 (N_10,In_13,In_246);
and U11 (N_11,In_710,In_715);
nand U12 (N_12,In_92,In_854);
and U13 (N_13,In_508,In_221);
and U14 (N_14,In_786,In_940);
and U15 (N_15,In_24,In_640);
nand U16 (N_16,In_159,In_910);
or U17 (N_17,In_191,In_842);
or U18 (N_18,In_874,In_401);
or U19 (N_19,In_970,In_793);
nor U20 (N_20,In_904,In_353);
or U21 (N_21,In_120,In_804);
nand U22 (N_22,In_718,In_732);
nand U23 (N_23,In_659,In_47);
or U24 (N_24,In_431,In_286);
and U25 (N_25,In_238,In_346);
or U26 (N_26,In_862,In_649);
or U27 (N_27,In_222,In_38);
or U28 (N_28,In_951,In_744);
and U29 (N_29,In_397,In_543);
nor U30 (N_30,In_262,In_564);
nor U31 (N_31,In_116,In_957);
nor U32 (N_32,In_986,In_303);
and U33 (N_33,In_822,In_214);
and U34 (N_34,In_810,In_199);
and U35 (N_35,In_954,In_667);
and U36 (N_36,In_441,In_1);
or U37 (N_37,In_448,In_607);
and U38 (N_38,In_805,In_472);
and U39 (N_39,In_408,In_840);
nor U40 (N_40,In_628,In_81);
xnor U41 (N_41,In_655,In_535);
nor U42 (N_42,In_178,In_557);
nand U43 (N_43,In_894,In_702);
nor U44 (N_44,In_155,In_174);
nand U45 (N_45,In_194,In_838);
nand U46 (N_46,In_296,In_121);
nor U47 (N_47,In_622,In_530);
or U48 (N_48,In_414,In_922);
and U49 (N_49,In_196,In_741);
or U50 (N_50,In_562,In_551);
and U51 (N_51,In_432,In_438);
or U52 (N_52,In_109,In_25);
and U53 (N_53,In_11,In_489);
nor U54 (N_54,In_887,In_897);
nand U55 (N_55,In_687,In_434);
and U56 (N_56,In_698,In_189);
nor U57 (N_57,In_639,In_405);
and U58 (N_58,In_375,In_934);
and U59 (N_59,In_924,In_572);
nor U60 (N_60,In_658,In_594);
or U61 (N_61,In_892,In_516);
and U62 (N_62,In_169,In_506);
nand U63 (N_63,In_23,In_634);
nand U64 (N_64,In_880,In_373);
or U65 (N_65,In_371,In_125);
nor U66 (N_66,In_550,In_998);
and U67 (N_67,In_705,In_925);
nor U68 (N_68,In_5,In_674);
nor U69 (N_69,In_792,In_439);
nand U70 (N_70,In_150,In_226);
nand U71 (N_71,In_604,In_457);
and U72 (N_72,In_392,In_421);
nor U73 (N_73,In_680,In_19);
xnor U74 (N_74,In_118,In_500);
or U75 (N_75,In_866,In_966);
or U76 (N_76,In_367,In_102);
nand U77 (N_77,In_832,In_336);
or U78 (N_78,In_219,In_532);
or U79 (N_79,In_22,In_955);
nor U80 (N_80,In_76,In_475);
and U81 (N_81,In_959,In_830);
or U82 (N_82,In_858,In_253);
nor U83 (N_83,In_578,In_278);
nor U84 (N_84,In_657,In_859);
or U85 (N_85,In_341,In_536);
or U86 (N_86,In_9,In_153);
and U87 (N_87,In_776,In_268);
or U88 (N_88,In_446,In_818);
nor U89 (N_89,In_15,In_724);
or U90 (N_90,In_101,In_701);
and U91 (N_91,In_476,In_135);
and U92 (N_92,In_146,In_759);
nand U93 (N_93,In_54,In_933);
or U94 (N_94,In_415,In_798);
and U95 (N_95,In_568,In_394);
and U96 (N_96,In_179,In_398);
and U97 (N_97,In_388,In_351);
and U98 (N_98,In_84,In_495);
nand U99 (N_99,In_236,In_983);
or U100 (N_100,In_85,In_378);
and U101 (N_101,In_198,In_615);
nor U102 (N_102,In_225,In_624);
and U103 (N_103,In_257,In_952);
nand U104 (N_104,In_345,In_730);
and U105 (N_105,In_216,In_212);
or U106 (N_106,In_743,In_613);
nand U107 (N_107,In_771,In_826);
and U108 (N_108,In_309,In_368);
and U109 (N_109,In_449,In_784);
nor U110 (N_110,In_91,In_295);
nand U111 (N_111,In_200,In_526);
or U112 (N_112,In_164,In_294);
nand U113 (N_113,In_946,In_455);
or U114 (N_114,In_413,In_546);
nor U115 (N_115,In_736,In_689);
or U116 (N_116,In_911,In_89);
and U117 (N_117,In_334,In_105);
nor U118 (N_118,In_94,In_239);
nor U119 (N_119,In_329,In_721);
or U120 (N_120,In_139,In_355);
nand U121 (N_121,In_941,In_699);
and U122 (N_122,In_708,In_704);
or U123 (N_123,In_44,In_507);
nand U124 (N_124,In_188,In_377);
nand U125 (N_125,In_809,In_787);
or U126 (N_126,In_611,In_206);
nor U127 (N_127,In_50,In_240);
nand U128 (N_128,In_918,In_923);
nand U129 (N_129,In_6,In_494);
or U130 (N_130,In_513,In_981);
nand U131 (N_131,In_32,In_993);
nor U132 (N_132,In_962,In_618);
and U133 (N_133,In_877,In_462);
nor U134 (N_134,In_453,In_220);
or U135 (N_135,In_151,In_133);
and U136 (N_136,In_127,In_168);
or U137 (N_137,In_289,In_785);
or U138 (N_138,In_267,In_907);
nand U139 (N_139,In_936,In_208);
or U140 (N_140,In_540,In_354);
nand U141 (N_141,In_204,In_347);
nor U142 (N_142,In_906,In_523);
and U143 (N_143,In_511,In_487);
nand U144 (N_144,In_28,In_987);
and U145 (N_145,In_359,In_534);
nor U146 (N_146,In_531,In_777);
nand U147 (N_147,In_181,In_423);
nand U148 (N_148,In_361,In_323);
and U149 (N_149,In_600,In_590);
nand U150 (N_150,In_638,In_313);
nand U151 (N_151,In_833,In_707);
nor U152 (N_152,In_606,In_447);
and U153 (N_153,In_547,In_984);
and U154 (N_154,In_114,In_130);
or U155 (N_155,In_661,In_849);
and U156 (N_156,In_678,In_813);
and U157 (N_157,In_422,In_893);
or U158 (N_158,In_860,In_348);
nand U159 (N_159,In_648,In_841);
or U160 (N_160,In_265,In_808);
nor U161 (N_161,In_861,In_524);
or U162 (N_162,In_790,In_128);
and U163 (N_163,In_688,In_463);
nor U164 (N_164,In_890,In_258);
or U165 (N_165,In_737,In_83);
and U166 (N_166,In_542,In_509);
nor U167 (N_167,In_310,In_856);
and U168 (N_168,In_305,In_868);
or U169 (N_169,In_14,In_938);
or U170 (N_170,In_95,In_297);
or U171 (N_171,In_502,In_773);
nand U172 (N_172,In_396,In_33);
and U173 (N_173,In_287,In_888);
nor U174 (N_174,In_298,In_58);
or U175 (N_175,In_620,In_454);
nor U176 (N_176,In_331,In_68);
nor U177 (N_177,In_37,In_276);
nor U178 (N_178,In_205,In_691);
and U179 (N_179,In_451,In_758);
or U180 (N_180,In_791,In_949);
or U181 (N_181,In_160,In_66);
and U182 (N_182,In_364,In_619);
nor U183 (N_183,In_393,In_775);
and U184 (N_184,In_385,In_270);
nor U185 (N_185,In_503,In_283);
and U186 (N_186,In_458,In_67);
nor U187 (N_187,In_968,In_749);
and U188 (N_188,In_709,In_126);
nor U189 (N_189,In_321,In_990);
nor U190 (N_190,In_681,In_977);
nand U191 (N_191,In_141,In_827);
nor U192 (N_192,In_132,In_450);
nand U193 (N_193,In_110,In_851);
nand U194 (N_194,In_703,In_609);
nand U195 (N_195,In_197,In_444);
nand U196 (N_196,In_603,In_601);
nand U197 (N_197,In_343,In_113);
or U198 (N_198,In_260,In_72);
and U199 (N_199,In_467,In_3);
and U200 (N_200,In_520,In_559);
nor U201 (N_201,In_663,In_73);
nor U202 (N_202,In_403,In_104);
nand U203 (N_203,In_525,In_549);
or U204 (N_204,In_35,In_100);
or U205 (N_205,In_145,In_815);
nor U206 (N_206,In_241,In_468);
nor U207 (N_207,In_51,In_825);
and U208 (N_208,In_484,In_190);
nand U209 (N_209,In_249,In_60);
nor U210 (N_210,In_210,In_685);
nor U211 (N_211,In_519,In_598);
nand U212 (N_212,In_745,In_356);
or U213 (N_213,In_576,In_716);
nor U214 (N_214,In_529,In_614);
nand U215 (N_215,In_602,In_218);
and U216 (N_216,In_522,In_53);
and U217 (N_217,In_693,In_544);
or U218 (N_218,In_728,In_428);
nor U219 (N_219,In_548,In_912);
nor U220 (N_220,In_586,In_560);
and U221 (N_221,In_686,In_0);
and U222 (N_222,In_376,In_909);
or U223 (N_223,In_848,In_124);
nor U224 (N_224,In_409,In_875);
and U225 (N_225,In_333,In_882);
nand U226 (N_226,In_473,In_610);
and U227 (N_227,In_751,In_989);
nand U228 (N_228,In_596,In_588);
or U229 (N_229,In_232,In_436);
and U230 (N_230,In_725,In_235);
nor U231 (N_231,In_485,In_641);
nor U232 (N_232,In_886,In_872);
and U233 (N_233,In_692,In_668);
and U234 (N_234,In_669,In_733);
or U235 (N_235,In_706,In_322);
nor U236 (N_236,In_574,In_209);
nand U237 (N_237,In_311,In_411);
nor U238 (N_238,In_39,In_795);
and U239 (N_239,In_261,In_779);
or U240 (N_240,In_646,In_746);
or U241 (N_241,In_651,In_896);
xor U242 (N_242,In_148,In_913);
and U243 (N_243,In_811,In_407);
nor U244 (N_244,In_597,In_683);
xnor U245 (N_245,In_871,In_553);
nor U246 (N_246,In_55,In_505);
or U247 (N_247,In_635,In_788);
nor U248 (N_248,In_521,In_342);
nor U249 (N_249,In_142,In_820);
nand U250 (N_250,In_850,In_433);
and U251 (N_251,In_819,In_335);
or U252 (N_252,In_935,In_99);
nand U253 (N_253,In_554,In_138);
nor U254 (N_254,In_427,In_93);
nand U255 (N_255,In_486,In_677);
nand U256 (N_256,In_713,In_481);
nand U257 (N_257,In_493,In_279);
nor U258 (N_258,In_477,In_783);
or U259 (N_259,In_982,In_916);
and U260 (N_260,In_325,In_381);
and U261 (N_261,In_592,In_799);
nand U262 (N_262,In_837,In_917);
xor U263 (N_263,In_327,In_581);
nor U264 (N_264,In_171,In_137);
or U265 (N_265,In_571,In_630);
nand U266 (N_266,In_660,In_836);
and U267 (N_267,In_230,In_821);
nand U268 (N_268,In_664,In_424);
nor U269 (N_269,In_344,In_972);
and U270 (N_270,In_565,In_229);
nor U271 (N_271,In_61,In_470);
and U272 (N_272,In_170,In_695);
nor U273 (N_273,In_65,In_299);
nand U274 (N_274,In_443,In_490);
nand U275 (N_275,In_869,In_491);
nand U276 (N_276,In_326,In_929);
nor U277 (N_277,In_264,In_243);
or U278 (N_278,In_625,In_202);
nand U279 (N_279,In_895,In_337);
nor U280 (N_280,In_173,In_994);
nand U281 (N_281,In_976,In_274);
nand U282 (N_282,In_781,In_752);
or U283 (N_283,In_57,In_379);
and U284 (N_284,In_437,In_307);
nor U285 (N_285,In_979,In_845);
nor U286 (N_286,In_175,In_48);
nand U287 (N_287,In_154,In_460);
xnor U288 (N_288,In_931,In_847);
and U289 (N_289,In_247,In_63);
and U290 (N_290,In_653,In_662);
or U291 (N_291,In_514,In_165);
nor U292 (N_292,In_528,In_269);
nand U293 (N_293,In_816,In_193);
nand U294 (N_294,In_480,In_814);
and U295 (N_295,In_723,In_797);
or U296 (N_296,In_45,In_829);
and U297 (N_297,In_304,In_20);
nand U298 (N_298,In_865,In_10);
nor U299 (N_299,In_971,In_762);
nor U300 (N_300,In_694,In_645);
nor U301 (N_301,In_584,In_177);
or U302 (N_302,In_90,In_315);
and U303 (N_303,In_273,In_533);
or U304 (N_304,In_629,In_734);
or U305 (N_305,In_144,In_839);
or U306 (N_306,In_82,In_380);
or U307 (N_307,In_26,In_612);
and U308 (N_308,In_88,In_419);
nand U309 (N_309,In_608,In_942);
or U310 (N_310,In_266,In_566);
nand U311 (N_311,In_201,In_969);
nand U312 (N_312,In_927,In_497);
nand U313 (N_313,In_747,In_162);
nor U314 (N_314,In_459,In_478);
and U315 (N_315,In_537,In_147);
and U316 (N_316,In_250,In_69);
nand U317 (N_317,In_761,In_158);
nand U318 (N_318,In_255,In_654);
and U319 (N_319,In_233,In_275);
nand U320 (N_320,In_31,In_471);
nor U321 (N_321,In_711,In_482);
nand U322 (N_322,In_103,In_7);
or U323 (N_323,In_328,In_558);
nand U324 (N_324,In_958,In_2);
and U325 (N_325,In_182,In_445);
nor U326 (N_326,In_318,In_418);
nor U327 (N_327,In_567,In_726);
nor U328 (N_328,In_186,In_400);
nor U329 (N_329,In_231,In_140);
or U330 (N_330,In_357,In_627);
or U331 (N_331,In_254,In_636);
or U332 (N_332,In_316,In_504);
nor U333 (N_333,In_290,In_756);
or U334 (N_334,In_853,In_782);
or U335 (N_335,In_425,In_831);
or U336 (N_336,In_474,In_245);
and U337 (N_337,In_374,In_555);
or U338 (N_338,In_948,In_314);
and U339 (N_339,In_926,In_985);
and U340 (N_340,In_330,In_79);
nand U341 (N_341,In_965,In_774);
nand U342 (N_342,In_452,In_722);
or U343 (N_343,In_339,In_843);
or U344 (N_344,In_49,In_945);
nor U345 (N_345,In_96,In_617);
and U346 (N_346,In_857,In_300);
and U347 (N_347,In_263,In_288);
or U348 (N_348,In_123,In_873);
and U349 (N_349,In_369,In_56);
nand U350 (N_350,In_442,In_690);
or U351 (N_351,In_891,In_997);
or U352 (N_352,In_563,In_98);
nand U353 (N_353,In_36,In_280);
and U354 (N_354,In_71,In_855);
or U355 (N_355,In_338,In_914);
nand U356 (N_356,In_763,In_697);
nor U357 (N_357,In_995,In_134);
or U358 (N_358,In_616,In_956);
or U359 (N_359,In_675,In_350);
or U360 (N_360,In_589,In_973);
nand U361 (N_361,In_767,In_676);
nor U362 (N_362,In_870,In_696);
nor U363 (N_363,In_915,In_881);
nand U364 (N_364,In_930,In_921);
or U365 (N_365,In_682,In_256);
nor U366 (N_366,In_964,In_920);
and U367 (N_367,In_883,In_932);
nor U368 (N_368,In_714,In_391);
and U369 (N_369,In_992,In_386);
and U370 (N_370,In_515,In_172);
or U371 (N_371,In_570,In_817);
and U372 (N_372,In_320,In_950);
or U373 (N_373,In_975,In_62);
nor U374 (N_374,In_632,In_492);
or U375 (N_375,In_770,In_406);
or U376 (N_376,In_980,In_947);
nor U377 (N_377,In_876,In_129);
nand U378 (N_378,In_720,In_878);
nand U379 (N_379,In_780,In_595);
or U380 (N_380,In_108,In_835);
nand U381 (N_381,In_652,In_277);
nor U382 (N_382,In_889,In_937);
xnor U383 (N_383,In_78,In_928);
nor U384 (N_384,In_244,In_301);
nor U385 (N_385,In_372,In_74);
nor U386 (N_386,In_12,In_27);
nor U387 (N_387,In_647,In_410);
and U388 (N_388,In_16,In_131);
nand U389 (N_389,In_852,In_748);
or U390 (N_390,In_621,In_203);
nor U391 (N_391,In_884,In_580);
and U392 (N_392,In_802,In_349);
nand U393 (N_393,In_953,In_898);
nand U394 (N_394,In_456,In_901);
or U395 (N_395,In_86,In_97);
or U396 (N_396,In_626,In_52);
or U397 (N_397,In_382,In_302);
nand U398 (N_398,In_885,In_324);
nor U399 (N_399,In_974,In_903);
nand U400 (N_400,In_631,In_806);
nor U401 (N_401,In_633,In_430);
nand U402 (N_402,In_479,In_389);
and U403 (N_403,In_117,In_605);
nand U404 (N_404,In_729,In_41);
or U405 (N_405,In_807,In_213);
or U406 (N_406,In_383,In_545);
nor U407 (N_407,In_944,In_465);
or U408 (N_408,In_469,In_823);
nor U409 (N_409,In_293,In_402);
and U410 (N_410,In_237,In_319);
or U411 (N_411,In_228,In_180);
or U412 (N_412,In_517,In_281);
and U413 (N_413,In_306,In_242);
nor U414 (N_414,In_824,In_387);
nor U415 (N_415,In_999,In_136);
nor U416 (N_416,In_195,In_988);
nand U417 (N_417,In_666,In_665);
nor U418 (N_418,In_252,In_963);
nand U419 (N_419,In_864,In_719);
and U420 (N_420,In_899,In_8);
or U421 (N_421,In_905,In_643);
nor U422 (N_422,In_156,In_152);
nor U423 (N_423,In_766,In_234);
nor U424 (N_424,In_753,In_754);
nand U425 (N_425,In_556,In_742);
or U426 (N_426,In_583,In_561);
nand U427 (N_427,In_259,In_656);
and U428 (N_428,In_64,In_960);
or U429 (N_429,In_670,In_757);
nor U430 (N_430,In_769,In_360);
nor U431 (N_431,In_582,In_184);
nand U432 (N_432,In_363,In_75);
or U433 (N_433,In_122,In_637);
nor U434 (N_434,In_908,In_575);
or U435 (N_435,In_18,In_498);
nand U436 (N_436,In_284,In_362);
and U437 (N_437,In_834,In_466);
and U438 (N_438,In_538,In_501);
nor U439 (N_439,In_4,In_731);
and U440 (N_440,In_579,In_107);
nand U441 (N_441,In_464,In_755);
nor U442 (N_442,In_772,In_317);
or U443 (N_443,In_527,In_846);
and U444 (N_444,In_166,In_573);
or U445 (N_445,In_712,In_30);
or U446 (N_446,In_143,In_800);
nor U447 (N_447,In_900,In_46);
or U448 (N_448,In_163,In_569);
or U449 (N_449,In_176,In_812);
nand U450 (N_450,In_483,In_420);
and U451 (N_451,In_215,In_370);
nand U452 (N_452,In_59,In_417);
and U453 (N_453,In_768,In_863);
or U454 (N_454,In_978,In_943);
or U455 (N_455,In_844,In_440);
or U456 (N_456,In_735,In_587);
nand U457 (N_457,In_285,In_211);
or U458 (N_458,In_801,In_778);
nor U459 (N_459,In_727,In_77);
nand U460 (N_460,In_591,In_599);
nor U461 (N_461,In_902,In_700);
nor U462 (N_462,In_112,In_384);
nand U463 (N_463,In_512,In_585);
and U464 (N_464,In_412,In_404);
nand U465 (N_465,In_996,In_291);
or U466 (N_466,In_518,In_679);
or U467 (N_467,In_740,In_185);
nor U468 (N_468,In_939,In_499);
nand U469 (N_469,In_879,In_510);
or U470 (N_470,In_764,In_577);
nand U471 (N_471,In_717,In_867);
nor U472 (N_472,In_803,In_42);
or U473 (N_473,In_282,In_919);
and U474 (N_474,In_358,In_435);
and U475 (N_475,In_593,In_365);
and U476 (N_476,In_760,In_40);
or U477 (N_477,In_991,In_426);
nand U478 (N_478,In_119,In_738);
nor U479 (N_479,In_541,In_366);
nor U480 (N_480,In_828,In_673);
or U481 (N_481,In_248,In_292);
or U482 (N_482,In_70,In_106);
nor U483 (N_483,In_223,In_34);
nor U484 (N_484,In_157,In_312);
or U485 (N_485,In_488,In_750);
or U486 (N_486,In_739,In_395);
xor U487 (N_487,In_21,In_789);
or U488 (N_488,In_796,In_29);
xnor U489 (N_489,In_399,In_461);
nand U490 (N_490,In_80,In_671);
xor U491 (N_491,In_227,In_272);
and U492 (N_492,In_161,In_650);
and U493 (N_493,In_251,In_207);
nor U494 (N_494,In_187,In_183);
nor U495 (N_495,In_794,In_539);
nand U496 (N_496,In_644,In_167);
or U497 (N_497,In_672,In_271);
and U498 (N_498,In_961,In_149);
nor U499 (N_499,In_192,In_552);
and U500 (N_500,In_121,In_172);
nand U501 (N_501,In_391,In_294);
nand U502 (N_502,In_154,In_820);
or U503 (N_503,In_241,In_32);
nor U504 (N_504,In_81,In_522);
nor U505 (N_505,In_925,In_840);
nor U506 (N_506,In_472,In_336);
nand U507 (N_507,In_909,In_523);
nand U508 (N_508,In_696,In_835);
and U509 (N_509,In_270,In_818);
nor U510 (N_510,In_540,In_895);
nor U511 (N_511,In_923,In_82);
or U512 (N_512,In_157,In_862);
nor U513 (N_513,In_873,In_900);
nand U514 (N_514,In_319,In_243);
nand U515 (N_515,In_408,In_634);
nor U516 (N_516,In_161,In_132);
nand U517 (N_517,In_986,In_242);
or U518 (N_518,In_629,In_740);
and U519 (N_519,In_774,In_148);
nand U520 (N_520,In_920,In_547);
nor U521 (N_521,In_560,In_14);
or U522 (N_522,In_360,In_721);
xor U523 (N_523,In_386,In_788);
nand U524 (N_524,In_271,In_650);
and U525 (N_525,In_803,In_682);
and U526 (N_526,In_612,In_61);
nor U527 (N_527,In_910,In_884);
nor U528 (N_528,In_6,In_527);
nand U529 (N_529,In_727,In_889);
nor U530 (N_530,In_909,In_354);
and U531 (N_531,In_183,In_381);
and U532 (N_532,In_452,In_497);
nor U533 (N_533,In_342,In_720);
nor U534 (N_534,In_297,In_955);
and U535 (N_535,In_3,In_226);
and U536 (N_536,In_932,In_509);
nand U537 (N_537,In_194,In_769);
nand U538 (N_538,In_932,In_284);
and U539 (N_539,In_453,In_674);
nor U540 (N_540,In_47,In_472);
nor U541 (N_541,In_380,In_303);
nor U542 (N_542,In_17,In_897);
or U543 (N_543,In_81,In_835);
nand U544 (N_544,In_406,In_393);
nand U545 (N_545,In_649,In_322);
nand U546 (N_546,In_842,In_245);
or U547 (N_547,In_706,In_417);
or U548 (N_548,In_373,In_533);
and U549 (N_549,In_94,In_431);
nand U550 (N_550,In_915,In_600);
nor U551 (N_551,In_728,In_344);
or U552 (N_552,In_952,In_286);
nor U553 (N_553,In_796,In_193);
nor U554 (N_554,In_129,In_372);
nor U555 (N_555,In_480,In_740);
or U556 (N_556,In_918,In_674);
nor U557 (N_557,In_149,In_705);
or U558 (N_558,In_158,In_5);
and U559 (N_559,In_497,In_391);
nor U560 (N_560,In_785,In_57);
nand U561 (N_561,In_232,In_384);
nor U562 (N_562,In_710,In_337);
nand U563 (N_563,In_968,In_581);
or U564 (N_564,In_971,In_842);
and U565 (N_565,In_157,In_7);
nor U566 (N_566,In_821,In_85);
or U567 (N_567,In_351,In_547);
nand U568 (N_568,In_717,In_358);
or U569 (N_569,In_727,In_778);
nand U570 (N_570,In_267,In_414);
nand U571 (N_571,In_31,In_221);
or U572 (N_572,In_504,In_17);
nor U573 (N_573,In_958,In_400);
and U574 (N_574,In_575,In_253);
or U575 (N_575,In_906,In_319);
nor U576 (N_576,In_877,In_833);
and U577 (N_577,In_26,In_714);
nor U578 (N_578,In_76,In_322);
nand U579 (N_579,In_509,In_303);
or U580 (N_580,In_270,In_566);
or U581 (N_581,In_318,In_193);
or U582 (N_582,In_878,In_583);
or U583 (N_583,In_564,In_376);
nor U584 (N_584,In_508,In_490);
nand U585 (N_585,In_410,In_845);
nor U586 (N_586,In_425,In_68);
and U587 (N_587,In_985,In_290);
or U588 (N_588,In_978,In_380);
nand U589 (N_589,In_89,In_646);
nor U590 (N_590,In_13,In_935);
nand U591 (N_591,In_276,In_238);
and U592 (N_592,In_64,In_472);
or U593 (N_593,In_239,In_803);
nor U594 (N_594,In_299,In_49);
nand U595 (N_595,In_656,In_702);
or U596 (N_596,In_170,In_405);
nand U597 (N_597,In_223,In_338);
nor U598 (N_598,In_738,In_331);
and U599 (N_599,In_487,In_235);
nand U600 (N_600,In_371,In_728);
nand U601 (N_601,In_359,In_196);
and U602 (N_602,In_812,In_893);
nor U603 (N_603,In_488,In_838);
nor U604 (N_604,In_871,In_472);
nand U605 (N_605,In_447,In_106);
and U606 (N_606,In_927,In_290);
nor U607 (N_607,In_302,In_56);
or U608 (N_608,In_831,In_462);
nor U609 (N_609,In_275,In_801);
nor U610 (N_610,In_487,In_34);
nand U611 (N_611,In_69,In_500);
nor U612 (N_612,In_489,In_982);
and U613 (N_613,In_622,In_201);
and U614 (N_614,In_923,In_372);
or U615 (N_615,In_492,In_994);
and U616 (N_616,In_818,In_328);
nand U617 (N_617,In_872,In_640);
nor U618 (N_618,In_165,In_0);
and U619 (N_619,In_254,In_56);
nand U620 (N_620,In_551,In_632);
nor U621 (N_621,In_974,In_228);
nand U622 (N_622,In_80,In_729);
or U623 (N_623,In_464,In_289);
nor U624 (N_624,In_260,In_676);
nand U625 (N_625,In_952,In_940);
nor U626 (N_626,In_903,In_298);
nand U627 (N_627,In_861,In_709);
nand U628 (N_628,In_265,In_394);
or U629 (N_629,In_195,In_303);
or U630 (N_630,In_558,In_204);
or U631 (N_631,In_929,In_64);
nand U632 (N_632,In_970,In_550);
or U633 (N_633,In_867,In_142);
and U634 (N_634,In_88,In_371);
nor U635 (N_635,In_178,In_985);
nand U636 (N_636,In_960,In_771);
and U637 (N_637,In_303,In_382);
nand U638 (N_638,In_677,In_575);
nand U639 (N_639,In_470,In_504);
nand U640 (N_640,In_958,In_893);
nand U641 (N_641,In_544,In_871);
nor U642 (N_642,In_111,In_813);
nand U643 (N_643,In_630,In_207);
or U644 (N_644,In_706,In_795);
xnor U645 (N_645,In_597,In_674);
and U646 (N_646,In_292,In_631);
nor U647 (N_647,In_672,In_671);
nor U648 (N_648,In_912,In_990);
and U649 (N_649,In_710,In_116);
nor U650 (N_650,In_493,In_291);
and U651 (N_651,In_734,In_793);
and U652 (N_652,In_414,In_73);
or U653 (N_653,In_66,In_525);
nor U654 (N_654,In_454,In_408);
and U655 (N_655,In_455,In_317);
or U656 (N_656,In_973,In_23);
nor U657 (N_657,In_187,In_127);
or U658 (N_658,In_875,In_801);
and U659 (N_659,In_35,In_753);
nor U660 (N_660,In_725,In_216);
or U661 (N_661,In_256,In_659);
or U662 (N_662,In_282,In_681);
nand U663 (N_663,In_848,In_602);
nor U664 (N_664,In_408,In_206);
nand U665 (N_665,In_780,In_897);
or U666 (N_666,In_614,In_469);
or U667 (N_667,In_690,In_909);
nand U668 (N_668,In_303,In_60);
or U669 (N_669,In_211,In_280);
nand U670 (N_670,In_174,In_823);
and U671 (N_671,In_948,In_377);
and U672 (N_672,In_798,In_981);
nor U673 (N_673,In_160,In_790);
nand U674 (N_674,In_784,In_465);
nor U675 (N_675,In_556,In_261);
nand U676 (N_676,In_457,In_869);
nand U677 (N_677,In_408,In_611);
nand U678 (N_678,In_698,In_726);
nor U679 (N_679,In_508,In_132);
and U680 (N_680,In_735,In_691);
and U681 (N_681,In_925,In_756);
nand U682 (N_682,In_319,In_192);
or U683 (N_683,In_607,In_430);
or U684 (N_684,In_905,In_667);
nand U685 (N_685,In_836,In_969);
nand U686 (N_686,In_372,In_156);
nor U687 (N_687,In_982,In_308);
or U688 (N_688,In_410,In_305);
and U689 (N_689,In_416,In_785);
and U690 (N_690,In_512,In_810);
nor U691 (N_691,In_654,In_843);
or U692 (N_692,In_668,In_172);
and U693 (N_693,In_409,In_91);
nand U694 (N_694,In_628,In_60);
or U695 (N_695,In_991,In_968);
nand U696 (N_696,In_910,In_767);
and U697 (N_697,In_120,In_521);
or U698 (N_698,In_2,In_915);
or U699 (N_699,In_266,In_716);
nor U700 (N_700,In_487,In_266);
or U701 (N_701,In_588,In_676);
nor U702 (N_702,In_692,In_656);
and U703 (N_703,In_435,In_513);
and U704 (N_704,In_997,In_588);
and U705 (N_705,In_343,In_388);
nor U706 (N_706,In_683,In_495);
and U707 (N_707,In_628,In_88);
nor U708 (N_708,In_517,In_186);
and U709 (N_709,In_579,In_827);
xor U710 (N_710,In_230,In_37);
nor U711 (N_711,In_716,In_83);
nand U712 (N_712,In_151,In_432);
and U713 (N_713,In_408,In_225);
nor U714 (N_714,In_241,In_17);
nand U715 (N_715,In_180,In_101);
nor U716 (N_716,In_314,In_853);
nand U717 (N_717,In_509,In_879);
nand U718 (N_718,In_294,In_990);
nand U719 (N_719,In_434,In_521);
and U720 (N_720,In_657,In_654);
and U721 (N_721,In_848,In_611);
xor U722 (N_722,In_533,In_672);
nand U723 (N_723,In_132,In_832);
and U724 (N_724,In_982,In_408);
or U725 (N_725,In_638,In_347);
and U726 (N_726,In_214,In_450);
nor U727 (N_727,In_120,In_278);
nor U728 (N_728,In_271,In_234);
or U729 (N_729,In_38,In_880);
nor U730 (N_730,In_661,In_663);
nand U731 (N_731,In_916,In_225);
and U732 (N_732,In_965,In_9);
nand U733 (N_733,In_799,In_166);
nor U734 (N_734,In_969,In_672);
xnor U735 (N_735,In_112,In_544);
and U736 (N_736,In_451,In_508);
or U737 (N_737,In_490,In_828);
nor U738 (N_738,In_769,In_524);
nand U739 (N_739,In_892,In_537);
or U740 (N_740,In_245,In_91);
nor U741 (N_741,In_82,In_349);
nand U742 (N_742,In_321,In_269);
and U743 (N_743,In_957,In_698);
nand U744 (N_744,In_592,In_441);
nor U745 (N_745,In_623,In_669);
nand U746 (N_746,In_617,In_730);
nand U747 (N_747,In_294,In_62);
nand U748 (N_748,In_87,In_35);
nor U749 (N_749,In_834,In_990);
and U750 (N_750,In_704,In_89);
and U751 (N_751,In_120,In_151);
or U752 (N_752,In_751,In_475);
and U753 (N_753,In_175,In_158);
nand U754 (N_754,In_2,In_900);
and U755 (N_755,In_711,In_349);
or U756 (N_756,In_973,In_9);
or U757 (N_757,In_383,In_346);
or U758 (N_758,In_395,In_657);
nor U759 (N_759,In_339,In_615);
nor U760 (N_760,In_947,In_608);
and U761 (N_761,In_192,In_84);
nor U762 (N_762,In_234,In_197);
nand U763 (N_763,In_559,In_622);
nand U764 (N_764,In_570,In_552);
nor U765 (N_765,In_311,In_801);
or U766 (N_766,In_922,In_295);
and U767 (N_767,In_70,In_934);
nand U768 (N_768,In_444,In_678);
and U769 (N_769,In_794,In_368);
or U770 (N_770,In_393,In_433);
and U771 (N_771,In_917,In_765);
and U772 (N_772,In_682,In_894);
or U773 (N_773,In_530,In_359);
or U774 (N_774,In_658,In_313);
nand U775 (N_775,In_380,In_775);
and U776 (N_776,In_246,In_708);
nand U777 (N_777,In_251,In_726);
and U778 (N_778,In_930,In_979);
or U779 (N_779,In_617,In_359);
nand U780 (N_780,In_702,In_263);
and U781 (N_781,In_502,In_313);
nand U782 (N_782,In_970,In_474);
and U783 (N_783,In_395,In_614);
and U784 (N_784,In_297,In_567);
or U785 (N_785,In_291,In_203);
nor U786 (N_786,In_868,In_613);
nand U787 (N_787,In_702,In_491);
nor U788 (N_788,In_430,In_768);
or U789 (N_789,In_906,In_970);
or U790 (N_790,In_354,In_223);
or U791 (N_791,In_612,In_187);
nand U792 (N_792,In_842,In_209);
nor U793 (N_793,In_842,In_617);
and U794 (N_794,In_304,In_971);
nand U795 (N_795,In_224,In_999);
nor U796 (N_796,In_93,In_831);
nor U797 (N_797,In_441,In_571);
nand U798 (N_798,In_932,In_243);
and U799 (N_799,In_248,In_74);
or U800 (N_800,In_619,In_730);
or U801 (N_801,In_877,In_75);
nor U802 (N_802,In_816,In_655);
and U803 (N_803,In_179,In_209);
nor U804 (N_804,In_385,In_630);
and U805 (N_805,In_93,In_497);
nand U806 (N_806,In_731,In_406);
nand U807 (N_807,In_659,In_714);
and U808 (N_808,In_953,In_357);
nand U809 (N_809,In_250,In_185);
and U810 (N_810,In_57,In_123);
nor U811 (N_811,In_160,In_71);
nand U812 (N_812,In_761,In_560);
nand U813 (N_813,In_338,In_778);
nor U814 (N_814,In_430,In_321);
nor U815 (N_815,In_660,In_150);
or U816 (N_816,In_811,In_537);
nor U817 (N_817,In_517,In_519);
nor U818 (N_818,In_550,In_431);
nand U819 (N_819,In_638,In_654);
and U820 (N_820,In_893,In_855);
xor U821 (N_821,In_611,In_734);
or U822 (N_822,In_641,In_116);
nor U823 (N_823,In_265,In_989);
or U824 (N_824,In_238,In_818);
or U825 (N_825,In_658,In_113);
nor U826 (N_826,In_922,In_143);
or U827 (N_827,In_658,In_836);
xnor U828 (N_828,In_813,In_300);
or U829 (N_829,In_50,In_729);
nand U830 (N_830,In_715,In_701);
nor U831 (N_831,In_231,In_755);
nor U832 (N_832,In_882,In_231);
nor U833 (N_833,In_231,In_724);
nor U834 (N_834,In_545,In_107);
nor U835 (N_835,In_538,In_252);
and U836 (N_836,In_246,In_624);
and U837 (N_837,In_279,In_836);
nor U838 (N_838,In_265,In_618);
and U839 (N_839,In_672,In_196);
nand U840 (N_840,In_608,In_365);
or U841 (N_841,In_39,In_553);
and U842 (N_842,In_793,In_764);
nor U843 (N_843,In_440,In_284);
nor U844 (N_844,In_743,In_337);
and U845 (N_845,In_240,In_51);
or U846 (N_846,In_214,In_371);
and U847 (N_847,In_151,In_380);
or U848 (N_848,In_946,In_641);
or U849 (N_849,In_969,In_223);
nand U850 (N_850,In_234,In_942);
nand U851 (N_851,In_694,In_611);
nor U852 (N_852,In_376,In_828);
nor U853 (N_853,In_425,In_1);
nand U854 (N_854,In_659,In_900);
nor U855 (N_855,In_229,In_920);
and U856 (N_856,In_860,In_620);
and U857 (N_857,In_66,In_767);
nand U858 (N_858,In_661,In_62);
xor U859 (N_859,In_408,In_278);
and U860 (N_860,In_159,In_76);
nor U861 (N_861,In_581,In_990);
and U862 (N_862,In_287,In_111);
nor U863 (N_863,In_187,In_834);
nand U864 (N_864,In_331,In_141);
or U865 (N_865,In_989,In_115);
or U866 (N_866,In_101,In_95);
and U867 (N_867,In_943,In_78);
nor U868 (N_868,In_504,In_140);
nand U869 (N_869,In_705,In_200);
nor U870 (N_870,In_122,In_776);
and U871 (N_871,In_776,In_907);
nor U872 (N_872,In_780,In_183);
and U873 (N_873,In_953,In_991);
nor U874 (N_874,In_378,In_842);
or U875 (N_875,In_477,In_737);
and U876 (N_876,In_412,In_597);
or U877 (N_877,In_842,In_683);
or U878 (N_878,In_725,In_350);
nor U879 (N_879,In_601,In_978);
and U880 (N_880,In_344,In_918);
nand U881 (N_881,In_651,In_827);
nand U882 (N_882,In_747,In_837);
and U883 (N_883,In_356,In_584);
nand U884 (N_884,In_331,In_634);
and U885 (N_885,In_810,In_389);
nor U886 (N_886,In_521,In_495);
and U887 (N_887,In_390,In_370);
and U888 (N_888,In_355,In_952);
nor U889 (N_889,In_241,In_751);
nand U890 (N_890,In_530,In_627);
and U891 (N_891,In_461,In_44);
nor U892 (N_892,In_891,In_711);
or U893 (N_893,In_416,In_442);
nand U894 (N_894,In_753,In_947);
xor U895 (N_895,In_80,In_219);
nor U896 (N_896,In_357,In_685);
nor U897 (N_897,In_641,In_152);
nor U898 (N_898,In_265,In_518);
and U899 (N_899,In_451,In_417);
nor U900 (N_900,In_241,In_73);
nor U901 (N_901,In_352,In_331);
nand U902 (N_902,In_476,In_138);
and U903 (N_903,In_740,In_583);
or U904 (N_904,In_881,In_206);
nor U905 (N_905,In_389,In_117);
and U906 (N_906,In_886,In_404);
and U907 (N_907,In_138,In_664);
nor U908 (N_908,In_709,In_763);
or U909 (N_909,In_715,In_924);
nor U910 (N_910,In_780,In_725);
nor U911 (N_911,In_581,In_679);
or U912 (N_912,In_64,In_510);
nand U913 (N_913,In_114,In_265);
and U914 (N_914,In_647,In_882);
and U915 (N_915,In_615,In_599);
or U916 (N_916,In_346,In_263);
nand U917 (N_917,In_3,In_496);
nand U918 (N_918,In_263,In_612);
and U919 (N_919,In_436,In_495);
and U920 (N_920,In_739,In_536);
nor U921 (N_921,In_717,In_108);
xor U922 (N_922,In_695,In_373);
or U923 (N_923,In_127,In_927);
and U924 (N_924,In_61,In_901);
or U925 (N_925,In_675,In_353);
or U926 (N_926,In_102,In_38);
nand U927 (N_927,In_103,In_833);
and U928 (N_928,In_241,In_368);
nor U929 (N_929,In_90,In_489);
nand U930 (N_930,In_677,In_438);
or U931 (N_931,In_885,In_236);
or U932 (N_932,In_921,In_192);
nand U933 (N_933,In_213,In_533);
nand U934 (N_934,In_256,In_184);
nor U935 (N_935,In_392,In_785);
nand U936 (N_936,In_161,In_882);
and U937 (N_937,In_702,In_546);
and U938 (N_938,In_906,In_228);
nand U939 (N_939,In_518,In_595);
nand U940 (N_940,In_649,In_532);
xor U941 (N_941,In_225,In_58);
or U942 (N_942,In_778,In_879);
nand U943 (N_943,In_209,In_840);
nand U944 (N_944,In_563,In_606);
nand U945 (N_945,In_100,In_587);
and U946 (N_946,In_124,In_855);
and U947 (N_947,In_687,In_173);
or U948 (N_948,In_725,In_487);
or U949 (N_949,In_372,In_833);
nor U950 (N_950,In_293,In_460);
nand U951 (N_951,In_891,In_389);
and U952 (N_952,In_192,In_545);
or U953 (N_953,In_428,In_344);
and U954 (N_954,In_44,In_638);
nand U955 (N_955,In_551,In_170);
or U956 (N_956,In_513,In_389);
or U957 (N_957,In_581,In_29);
nand U958 (N_958,In_163,In_290);
nand U959 (N_959,In_653,In_87);
or U960 (N_960,In_968,In_828);
and U961 (N_961,In_939,In_980);
or U962 (N_962,In_768,In_985);
and U963 (N_963,In_582,In_11);
and U964 (N_964,In_428,In_305);
or U965 (N_965,In_440,In_32);
nand U966 (N_966,In_658,In_852);
and U967 (N_967,In_290,In_161);
and U968 (N_968,In_127,In_938);
nand U969 (N_969,In_238,In_438);
and U970 (N_970,In_2,In_101);
nand U971 (N_971,In_955,In_708);
and U972 (N_972,In_185,In_317);
nand U973 (N_973,In_303,In_942);
or U974 (N_974,In_839,In_1);
and U975 (N_975,In_450,In_575);
nor U976 (N_976,In_813,In_804);
nor U977 (N_977,In_528,In_202);
and U978 (N_978,In_169,In_733);
or U979 (N_979,In_737,In_690);
nand U980 (N_980,In_290,In_976);
nor U981 (N_981,In_884,In_231);
nand U982 (N_982,In_378,In_564);
or U983 (N_983,In_411,In_968);
nand U984 (N_984,In_157,In_364);
nor U985 (N_985,In_442,In_63);
and U986 (N_986,In_50,In_183);
nor U987 (N_987,In_460,In_869);
or U988 (N_988,In_438,In_422);
nor U989 (N_989,In_40,In_685);
or U990 (N_990,In_829,In_895);
nand U991 (N_991,In_267,In_100);
or U992 (N_992,In_940,In_274);
or U993 (N_993,In_934,In_2);
or U994 (N_994,In_787,In_86);
and U995 (N_995,In_423,In_723);
nor U996 (N_996,In_406,In_475);
or U997 (N_997,In_367,In_734);
nor U998 (N_998,In_7,In_581);
nor U999 (N_999,In_616,In_300);
nand U1000 (N_1000,In_224,In_775);
or U1001 (N_1001,In_934,In_380);
and U1002 (N_1002,In_634,In_259);
and U1003 (N_1003,In_659,In_979);
and U1004 (N_1004,In_45,In_329);
nand U1005 (N_1005,In_907,In_890);
and U1006 (N_1006,In_575,In_497);
nand U1007 (N_1007,In_230,In_700);
and U1008 (N_1008,In_93,In_345);
or U1009 (N_1009,In_521,In_298);
or U1010 (N_1010,In_793,In_244);
and U1011 (N_1011,In_617,In_500);
nand U1012 (N_1012,In_186,In_507);
nor U1013 (N_1013,In_99,In_8);
nand U1014 (N_1014,In_665,In_515);
nand U1015 (N_1015,In_185,In_197);
and U1016 (N_1016,In_228,In_201);
and U1017 (N_1017,In_727,In_990);
nand U1018 (N_1018,In_529,In_890);
nor U1019 (N_1019,In_195,In_21);
and U1020 (N_1020,In_35,In_846);
nand U1021 (N_1021,In_150,In_179);
or U1022 (N_1022,In_240,In_528);
nor U1023 (N_1023,In_174,In_446);
and U1024 (N_1024,In_887,In_588);
and U1025 (N_1025,In_77,In_890);
or U1026 (N_1026,In_360,In_444);
nor U1027 (N_1027,In_501,In_700);
nand U1028 (N_1028,In_873,In_381);
nor U1029 (N_1029,In_559,In_890);
nand U1030 (N_1030,In_958,In_546);
nand U1031 (N_1031,In_999,In_635);
and U1032 (N_1032,In_193,In_157);
or U1033 (N_1033,In_47,In_49);
nor U1034 (N_1034,In_847,In_790);
or U1035 (N_1035,In_16,In_191);
nor U1036 (N_1036,In_664,In_193);
or U1037 (N_1037,In_18,In_401);
nand U1038 (N_1038,In_193,In_894);
and U1039 (N_1039,In_539,In_86);
nor U1040 (N_1040,In_248,In_97);
and U1041 (N_1041,In_43,In_866);
or U1042 (N_1042,In_95,In_377);
or U1043 (N_1043,In_605,In_544);
nor U1044 (N_1044,In_680,In_663);
or U1045 (N_1045,In_627,In_904);
and U1046 (N_1046,In_233,In_151);
nor U1047 (N_1047,In_11,In_534);
or U1048 (N_1048,In_723,In_909);
or U1049 (N_1049,In_583,In_424);
and U1050 (N_1050,In_129,In_323);
nor U1051 (N_1051,In_126,In_544);
nor U1052 (N_1052,In_642,In_671);
or U1053 (N_1053,In_676,In_284);
nand U1054 (N_1054,In_959,In_594);
nand U1055 (N_1055,In_750,In_159);
or U1056 (N_1056,In_504,In_847);
and U1057 (N_1057,In_798,In_618);
or U1058 (N_1058,In_679,In_520);
nand U1059 (N_1059,In_873,In_679);
and U1060 (N_1060,In_114,In_483);
and U1061 (N_1061,In_268,In_232);
or U1062 (N_1062,In_629,In_492);
or U1063 (N_1063,In_468,In_232);
nor U1064 (N_1064,In_248,In_58);
nor U1065 (N_1065,In_999,In_673);
nor U1066 (N_1066,In_519,In_514);
and U1067 (N_1067,In_384,In_535);
nand U1068 (N_1068,In_442,In_338);
or U1069 (N_1069,In_136,In_914);
and U1070 (N_1070,In_111,In_432);
nand U1071 (N_1071,In_331,In_915);
nor U1072 (N_1072,In_133,In_625);
and U1073 (N_1073,In_57,In_241);
and U1074 (N_1074,In_956,In_506);
nand U1075 (N_1075,In_776,In_151);
nand U1076 (N_1076,In_997,In_375);
or U1077 (N_1077,In_887,In_907);
and U1078 (N_1078,In_411,In_820);
and U1079 (N_1079,In_88,In_132);
and U1080 (N_1080,In_565,In_548);
nor U1081 (N_1081,In_593,In_325);
and U1082 (N_1082,In_479,In_349);
or U1083 (N_1083,In_241,In_985);
and U1084 (N_1084,In_455,In_125);
nor U1085 (N_1085,In_936,In_673);
or U1086 (N_1086,In_976,In_172);
and U1087 (N_1087,In_710,In_654);
or U1088 (N_1088,In_5,In_305);
or U1089 (N_1089,In_957,In_219);
or U1090 (N_1090,In_116,In_183);
nor U1091 (N_1091,In_310,In_950);
xor U1092 (N_1092,In_172,In_70);
nor U1093 (N_1093,In_501,In_656);
or U1094 (N_1094,In_786,In_393);
nand U1095 (N_1095,In_210,In_375);
or U1096 (N_1096,In_375,In_719);
nor U1097 (N_1097,In_853,In_921);
or U1098 (N_1098,In_499,In_103);
nand U1099 (N_1099,In_205,In_709);
nor U1100 (N_1100,In_897,In_950);
and U1101 (N_1101,In_83,In_731);
nor U1102 (N_1102,In_945,In_407);
and U1103 (N_1103,In_22,In_726);
nor U1104 (N_1104,In_97,In_565);
nand U1105 (N_1105,In_351,In_454);
and U1106 (N_1106,In_627,In_548);
nand U1107 (N_1107,In_992,In_677);
nor U1108 (N_1108,In_77,In_320);
and U1109 (N_1109,In_17,In_905);
nor U1110 (N_1110,In_987,In_301);
and U1111 (N_1111,In_343,In_157);
nor U1112 (N_1112,In_895,In_162);
nor U1113 (N_1113,In_663,In_326);
nor U1114 (N_1114,In_510,In_321);
nor U1115 (N_1115,In_965,In_184);
and U1116 (N_1116,In_663,In_90);
nand U1117 (N_1117,In_793,In_673);
xnor U1118 (N_1118,In_214,In_440);
nor U1119 (N_1119,In_907,In_505);
or U1120 (N_1120,In_548,In_996);
and U1121 (N_1121,In_615,In_522);
nand U1122 (N_1122,In_919,In_44);
nor U1123 (N_1123,In_677,In_331);
and U1124 (N_1124,In_651,In_233);
nand U1125 (N_1125,In_676,In_894);
and U1126 (N_1126,In_286,In_756);
or U1127 (N_1127,In_215,In_727);
and U1128 (N_1128,In_27,In_168);
or U1129 (N_1129,In_317,In_141);
and U1130 (N_1130,In_579,In_559);
nand U1131 (N_1131,In_509,In_275);
nor U1132 (N_1132,In_885,In_637);
nor U1133 (N_1133,In_867,In_482);
and U1134 (N_1134,In_110,In_519);
nor U1135 (N_1135,In_945,In_96);
nor U1136 (N_1136,In_113,In_879);
nand U1137 (N_1137,In_390,In_547);
nand U1138 (N_1138,In_581,In_702);
nor U1139 (N_1139,In_818,In_136);
or U1140 (N_1140,In_779,In_293);
and U1141 (N_1141,In_729,In_51);
or U1142 (N_1142,In_800,In_917);
or U1143 (N_1143,In_531,In_589);
nand U1144 (N_1144,In_209,In_555);
nand U1145 (N_1145,In_883,In_198);
nand U1146 (N_1146,In_304,In_881);
or U1147 (N_1147,In_64,In_269);
or U1148 (N_1148,In_755,In_792);
or U1149 (N_1149,In_555,In_807);
and U1150 (N_1150,In_864,In_985);
nand U1151 (N_1151,In_329,In_863);
and U1152 (N_1152,In_863,In_346);
or U1153 (N_1153,In_431,In_607);
nand U1154 (N_1154,In_227,In_275);
nand U1155 (N_1155,In_988,In_898);
nor U1156 (N_1156,In_86,In_403);
nand U1157 (N_1157,In_955,In_164);
or U1158 (N_1158,In_443,In_623);
nor U1159 (N_1159,In_918,In_212);
and U1160 (N_1160,In_60,In_694);
nor U1161 (N_1161,In_325,In_542);
nand U1162 (N_1162,In_193,In_401);
nand U1163 (N_1163,In_98,In_328);
nor U1164 (N_1164,In_566,In_419);
nand U1165 (N_1165,In_832,In_937);
nor U1166 (N_1166,In_670,In_549);
nand U1167 (N_1167,In_768,In_536);
or U1168 (N_1168,In_335,In_899);
and U1169 (N_1169,In_998,In_969);
nand U1170 (N_1170,In_56,In_273);
or U1171 (N_1171,In_646,In_893);
or U1172 (N_1172,In_599,In_788);
nand U1173 (N_1173,In_163,In_284);
and U1174 (N_1174,In_92,In_15);
or U1175 (N_1175,In_657,In_170);
and U1176 (N_1176,In_440,In_992);
or U1177 (N_1177,In_413,In_237);
nor U1178 (N_1178,In_740,In_112);
nand U1179 (N_1179,In_759,In_426);
or U1180 (N_1180,In_735,In_680);
or U1181 (N_1181,In_70,In_698);
nand U1182 (N_1182,In_249,In_478);
and U1183 (N_1183,In_705,In_278);
and U1184 (N_1184,In_476,In_816);
nand U1185 (N_1185,In_394,In_94);
nand U1186 (N_1186,In_633,In_402);
and U1187 (N_1187,In_110,In_120);
or U1188 (N_1188,In_523,In_573);
nand U1189 (N_1189,In_812,In_638);
nand U1190 (N_1190,In_595,In_465);
or U1191 (N_1191,In_673,In_729);
nor U1192 (N_1192,In_649,In_158);
and U1193 (N_1193,In_181,In_784);
and U1194 (N_1194,In_456,In_72);
and U1195 (N_1195,In_243,In_157);
and U1196 (N_1196,In_634,In_76);
and U1197 (N_1197,In_58,In_454);
or U1198 (N_1198,In_898,In_571);
or U1199 (N_1199,In_795,In_130);
nor U1200 (N_1200,In_187,In_352);
nand U1201 (N_1201,In_990,In_993);
and U1202 (N_1202,In_137,In_479);
nor U1203 (N_1203,In_765,In_256);
or U1204 (N_1204,In_818,In_156);
and U1205 (N_1205,In_182,In_649);
or U1206 (N_1206,In_948,In_356);
or U1207 (N_1207,In_429,In_798);
or U1208 (N_1208,In_132,In_169);
nor U1209 (N_1209,In_744,In_539);
or U1210 (N_1210,In_296,In_954);
or U1211 (N_1211,In_167,In_570);
nor U1212 (N_1212,In_790,In_551);
and U1213 (N_1213,In_109,In_331);
and U1214 (N_1214,In_896,In_933);
and U1215 (N_1215,In_714,In_965);
nand U1216 (N_1216,In_301,In_440);
nor U1217 (N_1217,In_235,In_421);
and U1218 (N_1218,In_156,In_557);
nand U1219 (N_1219,In_626,In_105);
and U1220 (N_1220,In_188,In_609);
and U1221 (N_1221,In_446,In_462);
nor U1222 (N_1222,In_118,In_233);
nor U1223 (N_1223,In_392,In_23);
and U1224 (N_1224,In_136,In_438);
nor U1225 (N_1225,In_782,In_592);
and U1226 (N_1226,In_443,In_267);
and U1227 (N_1227,In_246,In_7);
or U1228 (N_1228,In_60,In_167);
or U1229 (N_1229,In_161,In_766);
nand U1230 (N_1230,In_68,In_243);
nand U1231 (N_1231,In_53,In_542);
or U1232 (N_1232,In_36,In_393);
and U1233 (N_1233,In_638,In_623);
nand U1234 (N_1234,In_923,In_228);
nor U1235 (N_1235,In_47,In_712);
nor U1236 (N_1236,In_443,In_561);
nor U1237 (N_1237,In_81,In_418);
nor U1238 (N_1238,In_231,In_493);
and U1239 (N_1239,In_655,In_603);
nand U1240 (N_1240,In_3,In_907);
or U1241 (N_1241,In_305,In_126);
and U1242 (N_1242,In_630,In_619);
nor U1243 (N_1243,In_488,In_694);
or U1244 (N_1244,In_452,In_824);
nor U1245 (N_1245,In_469,In_0);
nor U1246 (N_1246,In_408,In_651);
nor U1247 (N_1247,In_502,In_154);
and U1248 (N_1248,In_205,In_166);
nor U1249 (N_1249,In_70,In_731);
nand U1250 (N_1250,In_428,In_250);
nor U1251 (N_1251,In_986,In_947);
nand U1252 (N_1252,In_357,In_242);
nor U1253 (N_1253,In_899,In_322);
and U1254 (N_1254,In_307,In_915);
and U1255 (N_1255,In_324,In_284);
nand U1256 (N_1256,In_297,In_798);
and U1257 (N_1257,In_589,In_77);
nor U1258 (N_1258,In_701,In_305);
and U1259 (N_1259,In_256,In_118);
nor U1260 (N_1260,In_31,In_304);
and U1261 (N_1261,In_633,In_659);
nand U1262 (N_1262,In_664,In_273);
nand U1263 (N_1263,In_425,In_86);
and U1264 (N_1264,In_840,In_520);
and U1265 (N_1265,In_109,In_853);
nand U1266 (N_1266,In_944,In_756);
nor U1267 (N_1267,In_829,In_565);
or U1268 (N_1268,In_187,In_820);
nor U1269 (N_1269,In_600,In_400);
nor U1270 (N_1270,In_219,In_840);
and U1271 (N_1271,In_754,In_670);
nand U1272 (N_1272,In_428,In_953);
and U1273 (N_1273,In_295,In_691);
nand U1274 (N_1274,In_567,In_553);
nand U1275 (N_1275,In_567,In_593);
nor U1276 (N_1276,In_978,In_377);
and U1277 (N_1277,In_235,In_602);
nand U1278 (N_1278,In_770,In_196);
or U1279 (N_1279,In_765,In_930);
nand U1280 (N_1280,In_344,In_352);
and U1281 (N_1281,In_983,In_714);
or U1282 (N_1282,In_867,In_714);
or U1283 (N_1283,In_459,In_351);
nand U1284 (N_1284,In_78,In_643);
nor U1285 (N_1285,In_675,In_365);
nand U1286 (N_1286,In_233,In_177);
nand U1287 (N_1287,In_389,In_486);
nor U1288 (N_1288,In_379,In_633);
nor U1289 (N_1289,In_238,In_290);
nor U1290 (N_1290,In_476,In_432);
nor U1291 (N_1291,In_715,In_778);
or U1292 (N_1292,In_111,In_970);
or U1293 (N_1293,In_564,In_795);
nand U1294 (N_1294,In_163,In_240);
or U1295 (N_1295,In_132,In_51);
or U1296 (N_1296,In_690,In_285);
nand U1297 (N_1297,In_666,In_80);
and U1298 (N_1298,In_138,In_256);
nand U1299 (N_1299,In_459,In_762);
and U1300 (N_1300,In_728,In_370);
nand U1301 (N_1301,In_630,In_711);
or U1302 (N_1302,In_573,In_608);
nor U1303 (N_1303,In_17,In_41);
nor U1304 (N_1304,In_934,In_489);
nand U1305 (N_1305,In_906,In_807);
or U1306 (N_1306,In_332,In_472);
or U1307 (N_1307,In_38,In_350);
or U1308 (N_1308,In_5,In_693);
nand U1309 (N_1309,In_471,In_51);
or U1310 (N_1310,In_411,In_401);
nor U1311 (N_1311,In_973,In_434);
and U1312 (N_1312,In_237,In_341);
nand U1313 (N_1313,In_839,In_404);
or U1314 (N_1314,In_374,In_55);
and U1315 (N_1315,In_475,In_498);
nor U1316 (N_1316,In_927,In_64);
nor U1317 (N_1317,In_894,In_699);
and U1318 (N_1318,In_252,In_449);
nor U1319 (N_1319,In_737,In_801);
nand U1320 (N_1320,In_172,In_438);
and U1321 (N_1321,In_624,In_254);
nand U1322 (N_1322,In_448,In_472);
or U1323 (N_1323,In_168,In_714);
or U1324 (N_1324,In_100,In_796);
nand U1325 (N_1325,In_341,In_71);
or U1326 (N_1326,In_672,In_18);
or U1327 (N_1327,In_342,In_760);
nand U1328 (N_1328,In_377,In_813);
nand U1329 (N_1329,In_685,In_413);
and U1330 (N_1330,In_32,In_420);
nand U1331 (N_1331,In_513,In_824);
or U1332 (N_1332,In_397,In_778);
or U1333 (N_1333,In_937,In_380);
nand U1334 (N_1334,In_857,In_85);
or U1335 (N_1335,In_785,In_431);
nor U1336 (N_1336,In_989,In_42);
nand U1337 (N_1337,In_657,In_289);
nor U1338 (N_1338,In_7,In_400);
nand U1339 (N_1339,In_636,In_946);
or U1340 (N_1340,In_420,In_549);
or U1341 (N_1341,In_729,In_771);
or U1342 (N_1342,In_48,In_100);
and U1343 (N_1343,In_748,In_144);
and U1344 (N_1344,In_83,In_290);
and U1345 (N_1345,In_670,In_583);
nand U1346 (N_1346,In_915,In_594);
and U1347 (N_1347,In_205,In_295);
nor U1348 (N_1348,In_532,In_31);
or U1349 (N_1349,In_286,In_773);
or U1350 (N_1350,In_520,In_17);
and U1351 (N_1351,In_316,In_432);
nor U1352 (N_1352,In_585,In_601);
and U1353 (N_1353,In_406,In_270);
nor U1354 (N_1354,In_897,In_74);
or U1355 (N_1355,In_118,In_14);
nand U1356 (N_1356,In_203,In_211);
nor U1357 (N_1357,In_754,In_354);
nand U1358 (N_1358,In_528,In_180);
nor U1359 (N_1359,In_497,In_191);
nand U1360 (N_1360,In_916,In_120);
nand U1361 (N_1361,In_468,In_163);
or U1362 (N_1362,In_634,In_779);
nand U1363 (N_1363,In_679,In_197);
nor U1364 (N_1364,In_386,In_131);
nor U1365 (N_1365,In_48,In_198);
nor U1366 (N_1366,In_384,In_164);
nor U1367 (N_1367,In_961,In_514);
nand U1368 (N_1368,In_681,In_958);
and U1369 (N_1369,In_483,In_552);
nand U1370 (N_1370,In_514,In_114);
xnor U1371 (N_1371,In_176,In_819);
nor U1372 (N_1372,In_993,In_992);
nor U1373 (N_1373,In_317,In_681);
nand U1374 (N_1374,In_605,In_962);
and U1375 (N_1375,In_756,In_848);
and U1376 (N_1376,In_772,In_325);
or U1377 (N_1377,In_198,In_395);
nand U1378 (N_1378,In_857,In_610);
nand U1379 (N_1379,In_385,In_94);
and U1380 (N_1380,In_513,In_48);
and U1381 (N_1381,In_281,In_913);
and U1382 (N_1382,In_301,In_49);
nand U1383 (N_1383,In_912,In_541);
nor U1384 (N_1384,In_928,In_597);
and U1385 (N_1385,In_810,In_184);
nand U1386 (N_1386,In_20,In_118);
nand U1387 (N_1387,In_107,In_731);
nand U1388 (N_1388,In_888,In_264);
or U1389 (N_1389,In_688,In_100);
and U1390 (N_1390,In_328,In_11);
nor U1391 (N_1391,In_189,In_844);
nand U1392 (N_1392,In_330,In_26);
nor U1393 (N_1393,In_494,In_178);
and U1394 (N_1394,In_872,In_14);
and U1395 (N_1395,In_664,In_741);
nand U1396 (N_1396,In_18,In_267);
and U1397 (N_1397,In_612,In_970);
nand U1398 (N_1398,In_960,In_74);
nand U1399 (N_1399,In_296,In_795);
or U1400 (N_1400,In_658,In_688);
or U1401 (N_1401,In_297,In_561);
nor U1402 (N_1402,In_374,In_698);
nand U1403 (N_1403,In_509,In_568);
and U1404 (N_1404,In_206,In_113);
or U1405 (N_1405,In_735,In_330);
nand U1406 (N_1406,In_112,In_887);
or U1407 (N_1407,In_41,In_93);
or U1408 (N_1408,In_757,In_72);
nor U1409 (N_1409,In_765,In_225);
or U1410 (N_1410,In_982,In_831);
nor U1411 (N_1411,In_464,In_893);
or U1412 (N_1412,In_725,In_2);
and U1413 (N_1413,In_829,In_474);
nor U1414 (N_1414,In_797,In_128);
nand U1415 (N_1415,In_744,In_805);
nor U1416 (N_1416,In_708,In_980);
nor U1417 (N_1417,In_908,In_4);
nor U1418 (N_1418,In_249,In_511);
and U1419 (N_1419,In_438,In_867);
nor U1420 (N_1420,In_153,In_231);
or U1421 (N_1421,In_792,In_183);
nor U1422 (N_1422,In_591,In_269);
xor U1423 (N_1423,In_750,In_151);
nand U1424 (N_1424,In_378,In_393);
and U1425 (N_1425,In_520,In_83);
xor U1426 (N_1426,In_986,In_24);
nand U1427 (N_1427,In_304,In_75);
nand U1428 (N_1428,In_184,In_592);
or U1429 (N_1429,In_300,In_740);
or U1430 (N_1430,In_152,In_945);
nand U1431 (N_1431,In_458,In_353);
and U1432 (N_1432,In_307,In_709);
or U1433 (N_1433,In_176,In_144);
nand U1434 (N_1434,In_445,In_916);
or U1435 (N_1435,In_388,In_559);
or U1436 (N_1436,In_5,In_394);
nand U1437 (N_1437,In_317,In_764);
nor U1438 (N_1438,In_329,In_827);
nand U1439 (N_1439,In_819,In_316);
and U1440 (N_1440,In_997,In_7);
or U1441 (N_1441,In_722,In_803);
or U1442 (N_1442,In_945,In_944);
nor U1443 (N_1443,In_238,In_414);
nand U1444 (N_1444,In_663,In_565);
and U1445 (N_1445,In_8,In_4);
or U1446 (N_1446,In_118,In_357);
nand U1447 (N_1447,In_323,In_446);
nand U1448 (N_1448,In_341,In_475);
or U1449 (N_1449,In_426,In_768);
and U1450 (N_1450,In_609,In_262);
nor U1451 (N_1451,In_748,In_947);
or U1452 (N_1452,In_644,In_970);
and U1453 (N_1453,In_922,In_409);
nor U1454 (N_1454,In_477,In_245);
and U1455 (N_1455,In_183,In_576);
or U1456 (N_1456,In_671,In_954);
and U1457 (N_1457,In_955,In_805);
or U1458 (N_1458,In_640,In_40);
nand U1459 (N_1459,In_618,In_272);
nand U1460 (N_1460,In_314,In_266);
and U1461 (N_1461,In_889,In_124);
nor U1462 (N_1462,In_568,In_850);
nand U1463 (N_1463,In_561,In_955);
or U1464 (N_1464,In_147,In_593);
nand U1465 (N_1465,In_456,In_880);
nand U1466 (N_1466,In_160,In_909);
nand U1467 (N_1467,In_654,In_11);
nand U1468 (N_1468,In_464,In_50);
nand U1469 (N_1469,In_248,In_37);
nand U1470 (N_1470,In_174,In_812);
nor U1471 (N_1471,In_885,In_926);
nor U1472 (N_1472,In_709,In_670);
nor U1473 (N_1473,In_126,In_289);
nand U1474 (N_1474,In_584,In_994);
nand U1475 (N_1475,In_507,In_122);
and U1476 (N_1476,In_35,In_969);
nand U1477 (N_1477,In_306,In_805);
or U1478 (N_1478,In_858,In_814);
or U1479 (N_1479,In_994,In_969);
nor U1480 (N_1480,In_900,In_555);
or U1481 (N_1481,In_656,In_53);
or U1482 (N_1482,In_752,In_622);
nor U1483 (N_1483,In_837,In_277);
nor U1484 (N_1484,In_357,In_311);
and U1485 (N_1485,In_741,In_577);
nand U1486 (N_1486,In_993,In_380);
nand U1487 (N_1487,In_416,In_687);
nand U1488 (N_1488,In_529,In_713);
and U1489 (N_1489,In_153,In_766);
nor U1490 (N_1490,In_605,In_115);
nor U1491 (N_1491,In_342,In_873);
nand U1492 (N_1492,In_151,In_530);
or U1493 (N_1493,In_855,In_413);
and U1494 (N_1494,In_360,In_282);
nor U1495 (N_1495,In_447,In_291);
nor U1496 (N_1496,In_42,In_221);
nor U1497 (N_1497,In_397,In_480);
or U1498 (N_1498,In_859,In_850);
nor U1499 (N_1499,In_81,In_344);
nor U1500 (N_1500,In_59,In_432);
or U1501 (N_1501,In_674,In_333);
or U1502 (N_1502,In_117,In_866);
nor U1503 (N_1503,In_291,In_211);
or U1504 (N_1504,In_751,In_499);
nor U1505 (N_1505,In_653,In_94);
or U1506 (N_1506,In_624,In_424);
nand U1507 (N_1507,In_46,In_451);
or U1508 (N_1508,In_247,In_996);
nor U1509 (N_1509,In_492,In_992);
nand U1510 (N_1510,In_394,In_150);
or U1511 (N_1511,In_236,In_422);
nand U1512 (N_1512,In_261,In_451);
nand U1513 (N_1513,In_700,In_885);
nand U1514 (N_1514,In_412,In_403);
or U1515 (N_1515,In_725,In_267);
or U1516 (N_1516,In_392,In_153);
or U1517 (N_1517,In_520,In_541);
or U1518 (N_1518,In_242,In_150);
nor U1519 (N_1519,In_868,In_860);
and U1520 (N_1520,In_369,In_917);
and U1521 (N_1521,In_210,In_664);
or U1522 (N_1522,In_419,In_826);
or U1523 (N_1523,In_263,In_531);
and U1524 (N_1524,In_947,In_843);
or U1525 (N_1525,In_947,In_501);
nand U1526 (N_1526,In_845,In_475);
nand U1527 (N_1527,In_119,In_837);
and U1528 (N_1528,In_304,In_219);
and U1529 (N_1529,In_346,In_867);
and U1530 (N_1530,In_940,In_180);
and U1531 (N_1531,In_788,In_664);
nand U1532 (N_1532,In_304,In_587);
nand U1533 (N_1533,In_596,In_530);
and U1534 (N_1534,In_729,In_388);
nand U1535 (N_1535,In_496,In_762);
nand U1536 (N_1536,In_434,In_965);
and U1537 (N_1537,In_908,In_432);
nor U1538 (N_1538,In_764,In_449);
and U1539 (N_1539,In_620,In_769);
nand U1540 (N_1540,In_263,In_96);
and U1541 (N_1541,In_946,In_338);
and U1542 (N_1542,In_881,In_508);
nand U1543 (N_1543,In_701,In_65);
and U1544 (N_1544,In_253,In_568);
nor U1545 (N_1545,In_775,In_315);
or U1546 (N_1546,In_247,In_470);
nor U1547 (N_1547,In_916,In_44);
and U1548 (N_1548,In_249,In_304);
and U1549 (N_1549,In_715,In_785);
nand U1550 (N_1550,In_322,In_29);
and U1551 (N_1551,In_242,In_806);
nor U1552 (N_1552,In_687,In_412);
nor U1553 (N_1553,In_476,In_963);
nand U1554 (N_1554,In_613,In_550);
xnor U1555 (N_1555,In_19,In_64);
xnor U1556 (N_1556,In_163,In_278);
nor U1557 (N_1557,In_94,In_293);
nand U1558 (N_1558,In_198,In_706);
or U1559 (N_1559,In_553,In_573);
and U1560 (N_1560,In_535,In_162);
nand U1561 (N_1561,In_976,In_293);
nand U1562 (N_1562,In_77,In_20);
or U1563 (N_1563,In_593,In_572);
and U1564 (N_1564,In_984,In_787);
and U1565 (N_1565,In_593,In_470);
nand U1566 (N_1566,In_952,In_723);
nor U1567 (N_1567,In_558,In_785);
or U1568 (N_1568,In_741,In_206);
nor U1569 (N_1569,In_567,In_202);
nor U1570 (N_1570,In_221,In_478);
nand U1571 (N_1571,In_618,In_287);
nor U1572 (N_1572,In_487,In_660);
nor U1573 (N_1573,In_749,In_691);
or U1574 (N_1574,In_699,In_194);
and U1575 (N_1575,In_849,In_747);
and U1576 (N_1576,In_979,In_804);
and U1577 (N_1577,In_999,In_518);
xor U1578 (N_1578,In_5,In_908);
or U1579 (N_1579,In_352,In_676);
nor U1580 (N_1580,In_327,In_670);
nand U1581 (N_1581,In_549,In_318);
or U1582 (N_1582,In_495,In_324);
and U1583 (N_1583,In_277,In_458);
nor U1584 (N_1584,In_988,In_754);
nand U1585 (N_1585,In_998,In_847);
nand U1586 (N_1586,In_292,In_548);
nand U1587 (N_1587,In_368,In_322);
nor U1588 (N_1588,In_159,In_838);
and U1589 (N_1589,In_759,In_897);
or U1590 (N_1590,In_270,In_551);
and U1591 (N_1591,In_30,In_246);
nand U1592 (N_1592,In_338,In_387);
and U1593 (N_1593,In_409,In_233);
or U1594 (N_1594,In_126,In_476);
and U1595 (N_1595,In_401,In_30);
nor U1596 (N_1596,In_174,In_889);
nand U1597 (N_1597,In_490,In_168);
nand U1598 (N_1598,In_457,In_838);
and U1599 (N_1599,In_242,In_268);
nor U1600 (N_1600,In_711,In_861);
or U1601 (N_1601,In_366,In_688);
nor U1602 (N_1602,In_681,In_59);
and U1603 (N_1603,In_614,In_79);
nor U1604 (N_1604,In_688,In_936);
or U1605 (N_1605,In_161,In_992);
nor U1606 (N_1606,In_896,In_821);
nand U1607 (N_1607,In_674,In_788);
xor U1608 (N_1608,In_976,In_876);
or U1609 (N_1609,In_291,In_927);
nand U1610 (N_1610,In_559,In_576);
and U1611 (N_1611,In_798,In_102);
and U1612 (N_1612,In_504,In_169);
and U1613 (N_1613,In_624,In_301);
nand U1614 (N_1614,In_345,In_681);
nor U1615 (N_1615,In_72,In_668);
nor U1616 (N_1616,In_203,In_908);
or U1617 (N_1617,In_445,In_433);
nor U1618 (N_1618,In_777,In_163);
nand U1619 (N_1619,In_376,In_677);
nand U1620 (N_1620,In_612,In_867);
nor U1621 (N_1621,In_345,In_44);
nor U1622 (N_1622,In_738,In_563);
or U1623 (N_1623,In_421,In_957);
or U1624 (N_1624,In_174,In_881);
and U1625 (N_1625,In_698,In_289);
and U1626 (N_1626,In_670,In_95);
nor U1627 (N_1627,In_645,In_27);
and U1628 (N_1628,In_530,In_438);
or U1629 (N_1629,In_154,In_970);
nand U1630 (N_1630,In_598,In_468);
nand U1631 (N_1631,In_189,In_107);
nor U1632 (N_1632,In_217,In_856);
or U1633 (N_1633,In_809,In_359);
nand U1634 (N_1634,In_875,In_679);
nor U1635 (N_1635,In_347,In_904);
or U1636 (N_1636,In_321,In_600);
and U1637 (N_1637,In_280,In_951);
nor U1638 (N_1638,In_326,In_192);
and U1639 (N_1639,In_680,In_548);
and U1640 (N_1640,In_296,In_489);
and U1641 (N_1641,In_590,In_266);
or U1642 (N_1642,In_686,In_657);
or U1643 (N_1643,In_213,In_595);
nand U1644 (N_1644,In_571,In_601);
nor U1645 (N_1645,In_646,In_666);
and U1646 (N_1646,In_808,In_520);
nand U1647 (N_1647,In_359,In_177);
and U1648 (N_1648,In_207,In_740);
and U1649 (N_1649,In_396,In_831);
nor U1650 (N_1650,In_247,In_707);
and U1651 (N_1651,In_164,In_281);
and U1652 (N_1652,In_105,In_145);
nor U1653 (N_1653,In_114,In_570);
and U1654 (N_1654,In_768,In_450);
nand U1655 (N_1655,In_47,In_426);
nor U1656 (N_1656,In_276,In_877);
and U1657 (N_1657,In_574,In_792);
nand U1658 (N_1658,In_836,In_752);
and U1659 (N_1659,In_889,In_740);
nor U1660 (N_1660,In_946,In_473);
xnor U1661 (N_1661,In_383,In_939);
and U1662 (N_1662,In_42,In_420);
or U1663 (N_1663,In_631,In_235);
and U1664 (N_1664,In_455,In_468);
nand U1665 (N_1665,In_92,In_9);
nand U1666 (N_1666,In_350,In_131);
nand U1667 (N_1667,In_726,In_45);
nand U1668 (N_1668,In_13,In_91);
and U1669 (N_1669,In_368,In_192);
or U1670 (N_1670,In_518,In_320);
and U1671 (N_1671,In_984,In_159);
or U1672 (N_1672,In_903,In_607);
nand U1673 (N_1673,In_957,In_19);
and U1674 (N_1674,In_287,In_135);
nor U1675 (N_1675,In_684,In_77);
nand U1676 (N_1676,In_709,In_226);
nand U1677 (N_1677,In_704,In_155);
and U1678 (N_1678,In_257,In_772);
nand U1679 (N_1679,In_947,In_862);
and U1680 (N_1680,In_990,In_205);
nor U1681 (N_1681,In_153,In_570);
or U1682 (N_1682,In_552,In_952);
nor U1683 (N_1683,In_843,In_667);
or U1684 (N_1684,In_72,In_632);
and U1685 (N_1685,In_360,In_318);
nand U1686 (N_1686,In_467,In_971);
or U1687 (N_1687,In_601,In_215);
or U1688 (N_1688,In_779,In_438);
nor U1689 (N_1689,In_82,In_2);
and U1690 (N_1690,In_832,In_956);
or U1691 (N_1691,In_508,In_303);
or U1692 (N_1692,In_300,In_341);
nor U1693 (N_1693,In_822,In_35);
nor U1694 (N_1694,In_266,In_505);
or U1695 (N_1695,In_98,In_873);
nand U1696 (N_1696,In_897,In_349);
and U1697 (N_1697,In_35,In_166);
and U1698 (N_1698,In_875,In_262);
or U1699 (N_1699,In_513,In_9);
and U1700 (N_1700,In_761,In_189);
and U1701 (N_1701,In_531,In_706);
nand U1702 (N_1702,In_56,In_597);
nor U1703 (N_1703,In_776,In_933);
nor U1704 (N_1704,In_24,In_762);
and U1705 (N_1705,In_682,In_340);
or U1706 (N_1706,In_776,In_838);
and U1707 (N_1707,In_215,In_389);
nand U1708 (N_1708,In_228,In_17);
and U1709 (N_1709,In_903,In_598);
or U1710 (N_1710,In_699,In_145);
nor U1711 (N_1711,In_949,In_777);
or U1712 (N_1712,In_718,In_918);
xnor U1713 (N_1713,In_118,In_698);
and U1714 (N_1714,In_716,In_319);
nor U1715 (N_1715,In_181,In_24);
and U1716 (N_1716,In_243,In_972);
or U1717 (N_1717,In_415,In_946);
nand U1718 (N_1718,In_664,In_721);
and U1719 (N_1719,In_889,In_239);
nand U1720 (N_1720,In_438,In_978);
and U1721 (N_1721,In_118,In_242);
nand U1722 (N_1722,In_550,In_661);
nand U1723 (N_1723,In_136,In_817);
and U1724 (N_1724,In_285,In_71);
and U1725 (N_1725,In_452,In_82);
nor U1726 (N_1726,In_444,In_802);
nand U1727 (N_1727,In_978,In_965);
nor U1728 (N_1728,In_49,In_851);
or U1729 (N_1729,In_553,In_521);
and U1730 (N_1730,In_151,In_572);
nor U1731 (N_1731,In_401,In_555);
and U1732 (N_1732,In_779,In_877);
or U1733 (N_1733,In_895,In_231);
or U1734 (N_1734,In_103,In_861);
and U1735 (N_1735,In_298,In_809);
nor U1736 (N_1736,In_24,In_61);
nor U1737 (N_1737,In_557,In_562);
or U1738 (N_1738,In_643,In_181);
nor U1739 (N_1739,In_921,In_195);
and U1740 (N_1740,In_784,In_518);
nor U1741 (N_1741,In_681,In_428);
nand U1742 (N_1742,In_226,In_428);
or U1743 (N_1743,In_48,In_362);
and U1744 (N_1744,In_815,In_945);
or U1745 (N_1745,In_411,In_979);
nand U1746 (N_1746,In_194,In_743);
or U1747 (N_1747,In_41,In_109);
or U1748 (N_1748,In_594,In_152);
nand U1749 (N_1749,In_600,In_44);
or U1750 (N_1750,In_179,In_666);
nand U1751 (N_1751,In_164,In_212);
or U1752 (N_1752,In_382,In_45);
and U1753 (N_1753,In_36,In_577);
nand U1754 (N_1754,In_695,In_654);
and U1755 (N_1755,In_863,In_609);
nand U1756 (N_1756,In_423,In_201);
and U1757 (N_1757,In_215,In_67);
nor U1758 (N_1758,In_26,In_496);
nor U1759 (N_1759,In_647,In_746);
nand U1760 (N_1760,In_232,In_547);
and U1761 (N_1761,In_737,In_241);
or U1762 (N_1762,In_782,In_147);
nand U1763 (N_1763,In_162,In_595);
or U1764 (N_1764,In_349,In_113);
or U1765 (N_1765,In_478,In_448);
or U1766 (N_1766,In_875,In_850);
nand U1767 (N_1767,In_720,In_66);
and U1768 (N_1768,In_195,In_517);
nand U1769 (N_1769,In_251,In_312);
and U1770 (N_1770,In_26,In_514);
nand U1771 (N_1771,In_443,In_125);
nand U1772 (N_1772,In_447,In_744);
or U1773 (N_1773,In_901,In_622);
and U1774 (N_1774,In_803,In_691);
nand U1775 (N_1775,In_221,In_356);
xnor U1776 (N_1776,In_817,In_381);
or U1777 (N_1777,In_750,In_876);
nand U1778 (N_1778,In_499,In_106);
or U1779 (N_1779,In_511,In_497);
and U1780 (N_1780,In_980,In_555);
or U1781 (N_1781,In_699,In_950);
nand U1782 (N_1782,In_15,In_180);
nor U1783 (N_1783,In_721,In_681);
or U1784 (N_1784,In_947,In_59);
or U1785 (N_1785,In_918,In_268);
and U1786 (N_1786,In_836,In_404);
and U1787 (N_1787,In_839,In_293);
nand U1788 (N_1788,In_558,In_84);
nand U1789 (N_1789,In_912,In_358);
and U1790 (N_1790,In_477,In_531);
nor U1791 (N_1791,In_384,In_174);
or U1792 (N_1792,In_680,In_376);
or U1793 (N_1793,In_309,In_816);
nor U1794 (N_1794,In_917,In_125);
or U1795 (N_1795,In_440,In_86);
and U1796 (N_1796,In_54,In_865);
nand U1797 (N_1797,In_660,In_563);
or U1798 (N_1798,In_952,In_451);
and U1799 (N_1799,In_803,In_797);
or U1800 (N_1800,In_955,In_521);
nand U1801 (N_1801,In_490,In_384);
or U1802 (N_1802,In_34,In_949);
nand U1803 (N_1803,In_337,In_902);
nand U1804 (N_1804,In_463,In_672);
nand U1805 (N_1805,In_176,In_592);
or U1806 (N_1806,In_947,In_216);
and U1807 (N_1807,In_449,In_94);
nor U1808 (N_1808,In_888,In_148);
nand U1809 (N_1809,In_209,In_866);
nor U1810 (N_1810,In_367,In_547);
nand U1811 (N_1811,In_784,In_644);
nand U1812 (N_1812,In_883,In_359);
nand U1813 (N_1813,In_218,In_723);
or U1814 (N_1814,In_83,In_817);
nand U1815 (N_1815,In_331,In_904);
and U1816 (N_1816,In_825,In_732);
nand U1817 (N_1817,In_878,In_567);
and U1818 (N_1818,In_828,In_935);
nor U1819 (N_1819,In_877,In_217);
nor U1820 (N_1820,In_656,In_545);
and U1821 (N_1821,In_576,In_895);
nor U1822 (N_1822,In_578,In_819);
and U1823 (N_1823,In_684,In_716);
and U1824 (N_1824,In_327,In_20);
nand U1825 (N_1825,In_28,In_650);
or U1826 (N_1826,In_690,In_513);
and U1827 (N_1827,In_486,In_96);
or U1828 (N_1828,In_89,In_843);
or U1829 (N_1829,In_123,In_919);
nand U1830 (N_1830,In_726,In_670);
nand U1831 (N_1831,In_967,In_725);
or U1832 (N_1832,In_741,In_932);
or U1833 (N_1833,In_38,In_779);
nor U1834 (N_1834,In_335,In_864);
and U1835 (N_1835,In_876,In_789);
nand U1836 (N_1836,In_89,In_95);
or U1837 (N_1837,In_33,In_246);
or U1838 (N_1838,In_965,In_545);
or U1839 (N_1839,In_419,In_418);
and U1840 (N_1840,In_592,In_11);
nor U1841 (N_1841,In_386,In_98);
or U1842 (N_1842,In_172,In_247);
or U1843 (N_1843,In_106,In_966);
and U1844 (N_1844,In_41,In_836);
or U1845 (N_1845,In_320,In_704);
and U1846 (N_1846,In_703,In_237);
nand U1847 (N_1847,In_764,In_944);
nor U1848 (N_1848,In_356,In_608);
nand U1849 (N_1849,In_905,In_211);
nand U1850 (N_1850,In_760,In_902);
nor U1851 (N_1851,In_535,In_757);
or U1852 (N_1852,In_852,In_933);
and U1853 (N_1853,In_369,In_604);
nor U1854 (N_1854,In_206,In_360);
nor U1855 (N_1855,In_174,In_90);
nor U1856 (N_1856,In_117,In_500);
nand U1857 (N_1857,In_443,In_118);
nor U1858 (N_1858,In_195,In_44);
nor U1859 (N_1859,In_539,In_2);
and U1860 (N_1860,In_439,In_796);
nand U1861 (N_1861,In_473,In_482);
nand U1862 (N_1862,In_511,In_795);
and U1863 (N_1863,In_184,In_201);
nand U1864 (N_1864,In_336,In_627);
or U1865 (N_1865,In_418,In_916);
or U1866 (N_1866,In_880,In_944);
nor U1867 (N_1867,In_876,In_338);
or U1868 (N_1868,In_310,In_495);
and U1869 (N_1869,In_585,In_92);
and U1870 (N_1870,In_366,In_577);
nand U1871 (N_1871,In_357,In_542);
nor U1872 (N_1872,In_149,In_523);
or U1873 (N_1873,In_793,In_608);
and U1874 (N_1874,In_484,In_738);
or U1875 (N_1875,In_465,In_167);
and U1876 (N_1876,In_133,In_263);
nand U1877 (N_1877,In_379,In_897);
and U1878 (N_1878,In_504,In_261);
nand U1879 (N_1879,In_191,In_96);
nand U1880 (N_1880,In_717,In_893);
nand U1881 (N_1881,In_963,In_586);
nor U1882 (N_1882,In_113,In_60);
and U1883 (N_1883,In_959,In_947);
nand U1884 (N_1884,In_767,In_20);
and U1885 (N_1885,In_925,In_807);
xnor U1886 (N_1886,In_686,In_531);
or U1887 (N_1887,In_830,In_51);
nor U1888 (N_1888,In_402,In_170);
and U1889 (N_1889,In_391,In_846);
nand U1890 (N_1890,In_272,In_228);
and U1891 (N_1891,In_152,In_682);
nor U1892 (N_1892,In_145,In_649);
and U1893 (N_1893,In_837,In_322);
nor U1894 (N_1894,In_293,In_982);
and U1895 (N_1895,In_674,In_215);
nor U1896 (N_1896,In_21,In_589);
nand U1897 (N_1897,In_705,In_518);
nor U1898 (N_1898,In_638,In_505);
nor U1899 (N_1899,In_350,In_474);
and U1900 (N_1900,In_535,In_97);
nor U1901 (N_1901,In_83,In_927);
or U1902 (N_1902,In_241,In_252);
nor U1903 (N_1903,In_452,In_385);
or U1904 (N_1904,In_682,In_178);
nand U1905 (N_1905,In_926,In_805);
and U1906 (N_1906,In_616,In_996);
and U1907 (N_1907,In_679,In_174);
xor U1908 (N_1908,In_485,In_698);
nand U1909 (N_1909,In_539,In_114);
and U1910 (N_1910,In_714,In_35);
or U1911 (N_1911,In_851,In_354);
nor U1912 (N_1912,In_863,In_245);
and U1913 (N_1913,In_316,In_607);
nand U1914 (N_1914,In_775,In_694);
nor U1915 (N_1915,In_142,In_310);
and U1916 (N_1916,In_507,In_812);
and U1917 (N_1917,In_453,In_51);
nor U1918 (N_1918,In_833,In_316);
nand U1919 (N_1919,In_695,In_218);
nand U1920 (N_1920,In_36,In_728);
nand U1921 (N_1921,In_363,In_498);
nor U1922 (N_1922,In_243,In_955);
nor U1923 (N_1923,In_374,In_701);
or U1924 (N_1924,In_986,In_30);
and U1925 (N_1925,In_550,In_315);
or U1926 (N_1926,In_223,In_452);
and U1927 (N_1927,In_273,In_829);
and U1928 (N_1928,In_310,In_425);
nand U1929 (N_1929,In_99,In_286);
or U1930 (N_1930,In_540,In_204);
or U1931 (N_1931,In_47,In_35);
and U1932 (N_1932,In_703,In_722);
or U1933 (N_1933,In_430,In_325);
nor U1934 (N_1934,In_127,In_970);
and U1935 (N_1935,In_500,In_96);
and U1936 (N_1936,In_781,In_289);
nor U1937 (N_1937,In_898,In_101);
nor U1938 (N_1938,In_932,In_36);
and U1939 (N_1939,In_11,In_773);
nand U1940 (N_1940,In_832,In_866);
nor U1941 (N_1941,In_648,In_268);
nor U1942 (N_1942,In_241,In_128);
nor U1943 (N_1943,In_822,In_369);
and U1944 (N_1944,In_761,In_33);
and U1945 (N_1945,In_572,In_731);
nand U1946 (N_1946,In_878,In_91);
nand U1947 (N_1947,In_552,In_919);
and U1948 (N_1948,In_43,In_757);
nand U1949 (N_1949,In_947,In_880);
and U1950 (N_1950,In_188,In_7);
or U1951 (N_1951,In_662,In_588);
and U1952 (N_1952,In_486,In_317);
nand U1953 (N_1953,In_307,In_202);
nor U1954 (N_1954,In_943,In_384);
and U1955 (N_1955,In_690,In_784);
and U1956 (N_1956,In_172,In_257);
nor U1957 (N_1957,In_877,In_848);
or U1958 (N_1958,In_246,In_234);
nor U1959 (N_1959,In_769,In_438);
or U1960 (N_1960,In_70,In_877);
and U1961 (N_1961,In_505,In_595);
and U1962 (N_1962,In_714,In_66);
or U1963 (N_1963,In_991,In_60);
xor U1964 (N_1964,In_149,In_353);
nor U1965 (N_1965,In_583,In_923);
and U1966 (N_1966,In_992,In_514);
and U1967 (N_1967,In_670,In_308);
nand U1968 (N_1968,In_359,In_903);
nand U1969 (N_1969,In_364,In_3);
or U1970 (N_1970,In_639,In_285);
or U1971 (N_1971,In_4,In_392);
nand U1972 (N_1972,In_35,In_809);
nand U1973 (N_1973,In_439,In_710);
and U1974 (N_1974,In_937,In_961);
or U1975 (N_1975,In_654,In_291);
or U1976 (N_1976,In_584,In_241);
or U1977 (N_1977,In_413,In_719);
and U1978 (N_1978,In_34,In_514);
and U1979 (N_1979,In_785,In_471);
and U1980 (N_1980,In_101,In_716);
nor U1981 (N_1981,In_924,In_325);
nand U1982 (N_1982,In_248,In_491);
nand U1983 (N_1983,In_567,In_746);
and U1984 (N_1984,In_197,In_861);
nand U1985 (N_1985,In_985,In_342);
nor U1986 (N_1986,In_178,In_19);
nor U1987 (N_1987,In_71,In_188);
nor U1988 (N_1988,In_12,In_709);
or U1989 (N_1989,In_454,In_121);
or U1990 (N_1990,In_831,In_742);
nand U1991 (N_1991,In_870,In_774);
or U1992 (N_1992,In_902,In_882);
nor U1993 (N_1993,In_377,In_523);
or U1994 (N_1994,In_918,In_876);
or U1995 (N_1995,In_259,In_499);
and U1996 (N_1996,In_598,In_416);
and U1997 (N_1997,In_141,In_903);
or U1998 (N_1998,In_458,In_688);
nor U1999 (N_1999,In_99,In_643);
and U2000 (N_2000,N_1339,N_345);
and U2001 (N_2001,N_1312,N_1909);
nand U2002 (N_2002,N_1875,N_1021);
and U2003 (N_2003,N_54,N_1180);
nand U2004 (N_2004,N_1902,N_1888);
and U2005 (N_2005,N_656,N_1401);
nor U2006 (N_2006,N_1452,N_752);
or U2007 (N_2007,N_1911,N_1137);
or U2008 (N_2008,N_1956,N_1067);
or U2009 (N_2009,N_1567,N_1157);
nor U2010 (N_2010,N_1172,N_1214);
or U2011 (N_2011,N_1359,N_171);
nand U2012 (N_2012,N_1018,N_1672);
nor U2013 (N_2013,N_1476,N_1616);
nand U2014 (N_2014,N_1127,N_1299);
nand U2015 (N_2015,N_1224,N_1729);
nor U2016 (N_2016,N_1637,N_238);
and U2017 (N_2017,N_747,N_914);
nor U2018 (N_2018,N_1140,N_204);
nor U2019 (N_2019,N_966,N_1763);
or U2020 (N_2020,N_1201,N_1785);
and U2021 (N_2021,N_550,N_323);
and U2022 (N_2022,N_1838,N_277);
and U2023 (N_2023,N_210,N_577);
nor U2024 (N_2024,N_1411,N_1091);
nor U2025 (N_2025,N_181,N_406);
and U2026 (N_2026,N_307,N_1030);
or U2027 (N_2027,N_1707,N_1602);
nor U2028 (N_2028,N_1044,N_1383);
or U2029 (N_2029,N_160,N_1207);
and U2030 (N_2030,N_251,N_197);
nand U2031 (N_2031,N_214,N_1151);
nand U2032 (N_2032,N_1378,N_498);
and U2033 (N_2033,N_33,N_514);
nor U2034 (N_2034,N_292,N_1527);
nor U2035 (N_2035,N_22,N_756);
nand U2036 (N_2036,N_749,N_949);
or U2037 (N_2037,N_567,N_103);
or U2038 (N_2038,N_132,N_542);
nor U2039 (N_2039,N_173,N_396);
and U2040 (N_2040,N_1495,N_1356);
and U2041 (N_2041,N_738,N_1494);
nand U2042 (N_2042,N_1417,N_1566);
xor U2043 (N_2043,N_1898,N_740);
nor U2044 (N_2044,N_1100,N_1295);
and U2045 (N_2045,N_1065,N_19);
nor U2046 (N_2046,N_748,N_604);
and U2047 (N_2047,N_872,N_658);
and U2048 (N_2048,N_458,N_881);
nand U2049 (N_2049,N_285,N_1914);
and U2050 (N_2050,N_1355,N_31);
nor U2051 (N_2051,N_1661,N_1505);
or U2052 (N_2052,N_534,N_140);
and U2053 (N_2053,N_1499,N_408);
nor U2054 (N_2054,N_1473,N_954);
nor U2055 (N_2055,N_1697,N_660);
or U2056 (N_2056,N_1215,N_1235);
or U2057 (N_2057,N_1249,N_967);
nor U2058 (N_2058,N_957,N_502);
and U2059 (N_2059,N_1415,N_681);
nor U2060 (N_2060,N_1904,N_597);
nand U2061 (N_2061,N_179,N_1714);
nand U2062 (N_2062,N_1639,N_308);
nor U2063 (N_2063,N_1492,N_1809);
and U2064 (N_2064,N_1574,N_212);
nor U2065 (N_2065,N_875,N_1803);
nor U2066 (N_2066,N_229,N_1485);
or U2067 (N_2067,N_236,N_1075);
and U2068 (N_2068,N_325,N_1549);
nor U2069 (N_2069,N_1974,N_1354);
and U2070 (N_2070,N_221,N_338);
nand U2071 (N_2071,N_1597,N_719);
and U2072 (N_2072,N_1063,N_378);
nor U2073 (N_2073,N_669,N_1525);
nand U2074 (N_2074,N_1621,N_402);
or U2075 (N_2075,N_692,N_1744);
nand U2076 (N_2076,N_168,N_578);
nand U2077 (N_2077,N_1122,N_541);
nand U2078 (N_2078,N_1040,N_1456);
and U2079 (N_2079,N_1852,N_1942);
or U2080 (N_2080,N_1572,N_813);
nor U2081 (N_2081,N_1885,N_241);
nand U2082 (N_2082,N_1160,N_815);
and U2083 (N_2083,N_932,N_1404);
nor U2084 (N_2084,N_1928,N_1291);
or U2085 (N_2085,N_1773,N_150);
or U2086 (N_2086,N_265,N_650);
nor U2087 (N_2087,N_1442,N_1728);
nand U2088 (N_2088,N_226,N_1691);
nand U2089 (N_2089,N_1614,N_979);
nand U2090 (N_2090,N_1571,N_1144);
or U2091 (N_2091,N_939,N_1937);
or U2092 (N_2092,N_1818,N_1892);
and U2093 (N_2093,N_1568,N_1821);
or U2094 (N_2094,N_1406,N_341);
nor U2095 (N_2095,N_699,N_610);
nor U2096 (N_2096,N_721,N_97);
and U2097 (N_2097,N_1430,N_614);
nand U2098 (N_2098,N_1438,N_143);
or U2099 (N_2099,N_486,N_905);
or U2100 (N_2100,N_1164,N_958);
nor U2101 (N_2101,N_1074,N_574);
or U2102 (N_2102,N_470,N_503);
nand U2103 (N_2103,N_987,N_829);
nor U2104 (N_2104,N_400,N_394);
nor U2105 (N_2105,N_1273,N_1258);
nor U2106 (N_2106,N_924,N_1623);
nand U2107 (N_2107,N_1519,N_1675);
nor U2108 (N_2108,N_1446,N_1987);
or U2109 (N_2109,N_781,N_484);
and U2110 (N_2110,N_831,N_1545);
nand U2111 (N_2111,N_1622,N_778);
nand U2112 (N_2112,N_224,N_1244);
and U2113 (N_2113,N_446,N_342);
nor U2114 (N_2114,N_675,N_488);
and U2115 (N_2115,N_951,N_1783);
and U2116 (N_2116,N_475,N_1382);
and U2117 (N_2117,N_148,N_1003);
nor U2118 (N_2118,N_439,N_499);
or U2119 (N_2119,N_1116,N_18);
nor U2120 (N_2120,N_569,N_363);
nor U2121 (N_2121,N_1613,N_459);
nor U2122 (N_2122,N_1373,N_870);
and U2123 (N_2123,N_690,N_844);
nor U2124 (N_2124,N_476,N_1789);
nor U2125 (N_2125,N_588,N_672);
nor U2126 (N_2126,N_931,N_727);
nand U2127 (N_2127,N_1179,N_3);
nand U2128 (N_2128,N_14,N_773);
nor U2129 (N_2129,N_595,N_843);
nor U2130 (N_2130,N_964,N_633);
and U2131 (N_2131,N_665,N_388);
or U2132 (N_2132,N_465,N_1477);
xnor U2133 (N_2133,N_1688,N_1192);
nor U2134 (N_2134,N_1762,N_217);
nor U2135 (N_2135,N_48,N_1706);
nor U2136 (N_2136,N_134,N_1015);
and U2137 (N_2137,N_1115,N_1200);
nor U2138 (N_2138,N_1606,N_1757);
or U2139 (N_2139,N_131,N_1325);
and U2140 (N_2140,N_348,N_852);
and U2141 (N_2141,N_69,N_1197);
and U2142 (N_2142,N_1285,N_1288);
and U2143 (N_2143,N_575,N_1223);
nand U2144 (N_2144,N_1548,N_1882);
or U2145 (N_2145,N_70,N_1472);
or U2146 (N_2146,N_27,N_1580);
or U2147 (N_2147,N_860,N_1528);
nand U2148 (N_2148,N_1129,N_1610);
xnor U2149 (N_2149,N_1588,N_823);
nand U2150 (N_2150,N_1377,N_1700);
and U2151 (N_2151,N_728,N_935);
or U2152 (N_2152,N_274,N_203);
or U2153 (N_2153,N_1752,N_1256);
and U2154 (N_2154,N_929,N_840);
and U2155 (N_2155,N_587,N_771);
nor U2156 (N_2156,N_1195,N_188);
nand U2157 (N_2157,N_1212,N_869);
and U2158 (N_2158,N_1118,N_413);
or U2159 (N_2159,N_118,N_871);
and U2160 (N_2160,N_1049,N_1768);
or U2161 (N_2161,N_834,N_1252);
and U2162 (N_2162,N_456,N_846);
nand U2163 (N_2163,N_627,N_215);
or U2164 (N_2164,N_1275,N_15);
nor U2165 (N_2165,N_0,N_1418);
or U2166 (N_2166,N_1884,N_1802);
nand U2167 (N_2167,N_921,N_1635);
nor U2168 (N_2168,N_910,N_237);
nand U2169 (N_2169,N_1664,N_260);
nor U2170 (N_2170,N_1967,N_735);
nor U2171 (N_2171,N_1736,N_1400);
nand U2172 (N_2172,N_85,N_1931);
and U2173 (N_2173,N_189,N_1371);
nand U2174 (N_2174,N_89,N_809);
nand U2175 (N_2175,N_438,N_1008);
and U2176 (N_2176,N_1703,N_376);
or U2177 (N_2177,N_1958,N_725);
nor U2178 (N_2178,N_377,N_75);
nor U2179 (N_2179,N_20,N_1631);
nor U2180 (N_2180,N_828,N_379);
or U2181 (N_2181,N_1844,N_1829);
or U2182 (N_2182,N_1169,N_1426);
nor U2183 (N_2183,N_99,N_947);
and U2184 (N_2184,N_700,N_1464);
and U2185 (N_2185,N_1301,N_13);
nor U2186 (N_2186,N_718,N_362);
or U2187 (N_2187,N_422,N_1257);
or U2188 (N_2188,N_1489,N_1715);
or U2189 (N_2189,N_741,N_1072);
nor U2190 (N_2190,N_1685,N_246);
nor U2191 (N_2191,N_712,N_290);
or U2192 (N_2192,N_873,N_1658);
nand U2193 (N_2193,N_1579,N_688);
or U2194 (N_2194,N_248,N_1670);
nand U2195 (N_2195,N_57,N_1858);
nand U2196 (N_2196,N_982,N_205);
and U2197 (N_2197,N_454,N_1813);
nand U2198 (N_2198,N_1088,N_1936);
and U2199 (N_2199,N_1727,N_1893);
or U2200 (N_2200,N_415,N_1319);
and U2201 (N_2201,N_1510,N_1165);
nor U2202 (N_2202,N_1791,N_1334);
or U2203 (N_2203,N_1268,N_758);
nand U2204 (N_2204,N_30,N_591);
and U2205 (N_2205,N_287,N_51);
or U2206 (N_2206,N_509,N_293);
or U2207 (N_2207,N_783,N_1598);
and U2208 (N_2208,N_360,N_1361);
nand U2209 (N_2209,N_1923,N_862);
nor U2210 (N_2210,N_1384,N_350);
or U2211 (N_2211,N_737,N_62);
and U2212 (N_2212,N_1994,N_745);
nand U2213 (N_2213,N_1500,N_1905);
and U2214 (N_2214,N_676,N_332);
nand U2215 (N_2215,N_156,N_880);
nor U2216 (N_2216,N_1376,N_11);
nand U2217 (N_2217,N_616,N_144);
and U2218 (N_2218,N_1191,N_1663);
xor U2219 (N_2219,N_866,N_1344);
or U2220 (N_2220,N_1808,N_938);
and U2221 (N_2221,N_1081,N_762);
and U2222 (N_2222,N_418,N_1463);
and U2223 (N_2223,N_649,N_1996);
nor U2224 (N_2224,N_785,N_1038);
nand U2225 (N_2225,N_984,N_1094);
nor U2226 (N_2226,N_992,N_1540);
and U2227 (N_2227,N_1053,N_1759);
nand U2228 (N_2228,N_301,N_108);
nand U2229 (N_2229,N_281,N_1963);
nor U2230 (N_2230,N_708,N_1997);
nor U2231 (N_2231,N_733,N_1513);
or U2232 (N_2232,N_1812,N_1991);
or U2233 (N_2233,N_1145,N_874);
nor U2234 (N_2234,N_55,N_1704);
nand U2235 (N_2235,N_784,N_1462);
or U2236 (N_2236,N_1424,N_768);
and U2237 (N_2237,N_1303,N_1222);
and U2238 (N_2238,N_1925,N_1047);
and U2239 (N_2239,N_1381,N_1872);
or U2240 (N_2240,N_1913,N_253);
nor U2241 (N_2241,N_1238,N_1391);
or U2242 (N_2242,N_1086,N_1010);
or U2243 (N_2243,N_1447,N_1427);
nand U2244 (N_2244,N_539,N_538);
nand U2245 (N_2245,N_732,N_995);
or U2246 (N_2246,N_172,N_1874);
nand U2247 (N_2247,N_1321,N_651);
nand U2248 (N_2248,N_1612,N_1867);
or U2249 (N_2249,N_84,N_1877);
nor U2250 (N_2250,N_601,N_1971);
nor U2251 (N_2251,N_1428,N_1363);
or U2252 (N_2252,N_1595,N_1042);
or U2253 (N_2253,N_190,N_280);
nor U2254 (N_2254,N_1113,N_29);
or U2255 (N_2255,N_410,N_1521);
and U2256 (N_2256,N_522,N_1205);
nor U2257 (N_2257,N_117,N_303);
xor U2258 (N_2258,N_384,N_368);
or U2259 (N_2259,N_1724,N_295);
or U2260 (N_2260,N_1246,N_437);
nand U2261 (N_2261,N_1405,N_311);
nand U2262 (N_2262,N_107,N_1501);
and U2263 (N_2263,N_1362,N_1920);
or U2264 (N_2264,N_1776,N_1403);
or U2265 (N_2265,N_1058,N_417);
or U2266 (N_2266,N_657,N_937);
and U2267 (N_2267,N_716,N_1856);
nand U2268 (N_2268,N_1467,N_1175);
and U2269 (N_2269,N_1883,N_1340);
nand U2270 (N_2270,N_157,N_792);
or U2271 (N_2271,N_1850,N_276);
nor U2272 (N_2272,N_1769,N_485);
and U2273 (N_2273,N_1313,N_623);
and U2274 (N_2274,N_339,N_6);
nand U2275 (N_2275,N_349,N_1608);
nor U2276 (N_2276,N_463,N_477);
and U2277 (N_2277,N_1307,N_492);
nor U2278 (N_2278,N_1147,N_1270);
and U2279 (N_2279,N_1202,N_1276);
and U2280 (N_2280,N_506,N_808);
or U2281 (N_2281,N_892,N_606);
or U2282 (N_2282,N_666,N_533);
or U2283 (N_2283,N_1385,N_1799);
and U2284 (N_2284,N_1332,N_590);
nor U2285 (N_2285,N_1203,N_1233);
and U2286 (N_2286,N_1474,N_472);
nand U2287 (N_2287,N_1109,N_557);
nor U2288 (N_2288,N_1734,N_1629);
nor U2289 (N_2289,N_664,N_739);
and U2290 (N_2290,N_1643,N_1782);
or U2291 (N_2291,N_867,N_1692);
or U2292 (N_2292,N_1228,N_309);
nand U2293 (N_2293,N_894,N_1972);
and U2294 (N_2294,N_1742,N_136);
nand U2295 (N_2295,N_802,N_983);
and U2296 (N_2296,N_646,N_1369);
nor U2297 (N_2297,N_1399,N_1988);
and U2298 (N_2298,N_1265,N_1620);
or U2299 (N_2299,N_1226,N_826);
and U2300 (N_2300,N_1482,N_1443);
and U2301 (N_2301,N_162,N_491);
nand U2302 (N_2302,N_1287,N_970);
nor U2303 (N_2303,N_1817,N_1037);
nand U2304 (N_2304,N_701,N_1266);
or U2305 (N_2305,N_803,N_1459);
or U2306 (N_2306,N_640,N_192);
or U2307 (N_2307,N_562,N_1824);
or U2308 (N_2308,N_1669,N_1576);
and U2309 (N_2309,N_155,N_639);
and U2310 (N_2310,N_1792,N_464);
or U2311 (N_2311,N_674,N_1043);
and U2312 (N_2312,N_1078,N_959);
nand U2313 (N_2313,N_754,N_796);
and U2314 (N_2314,N_1444,N_93);
nor U2315 (N_2315,N_1645,N_72);
and U2316 (N_2316,N_1950,N_523);
and U2317 (N_2317,N_1733,N_202);
nand U2318 (N_2318,N_1564,N_1740);
nand U2319 (N_2319,N_1448,N_1896);
nor U2320 (N_2320,N_1601,N_1712);
nor U2321 (N_2321,N_1333,N_1341);
nand U2322 (N_2322,N_351,N_952);
or U2323 (N_2323,N_806,N_908);
nand U2324 (N_2324,N_724,N_429);
or U2325 (N_2325,N_495,N_1007);
nor U2326 (N_2326,N_507,N_1819);
nor U2327 (N_2327,N_256,N_988);
or U2328 (N_2328,N_1360,N_1751);
nor U2329 (N_2329,N_1502,N_1563);
and U2330 (N_2330,N_367,N_1136);
and U2331 (N_2331,N_252,N_884);
or U2332 (N_2332,N_49,N_483);
nand U2333 (N_2333,N_1310,N_960);
nand U2334 (N_2334,N_1880,N_1586);
or U2335 (N_2335,N_1055,N_1627);
nand U2336 (N_2336,N_4,N_1085);
and U2337 (N_2337,N_1358,N_381);
nand U2338 (N_2338,N_1283,N_366);
nor U2339 (N_2339,N_1573,N_1717);
nand U2340 (N_2340,N_1076,N_1922);
or U2341 (N_2341,N_294,N_705);
nand U2342 (N_2342,N_299,N_1000);
nor U2343 (N_2343,N_310,N_573);
nor U2344 (N_2344,N_397,N_1365);
nor U2345 (N_2345,N_1408,N_556);
nand U2346 (N_2346,N_426,N_865);
nand U2347 (N_2347,N_146,N_184);
nand U2348 (N_2348,N_279,N_167);
and U2349 (N_2349,N_1992,N_347);
and U2350 (N_2350,N_1646,N_1322);
or U2351 (N_2351,N_609,N_1798);
nor U2352 (N_2352,N_930,N_153);
or U2353 (N_2353,N_23,N_1132);
nor U2354 (N_2354,N_1368,N_1357);
and U2355 (N_2355,N_767,N_1772);
or U2356 (N_2356,N_1335,N_1183);
and U2357 (N_2357,N_673,N_878);
and U2358 (N_2358,N_450,N_133);
nor U2359 (N_2359,N_1533,N_1243);
nand U2360 (N_2360,N_1536,N_1407);
xor U2361 (N_2361,N_312,N_239);
and U2362 (N_2362,N_1957,N_558);
nand U2363 (N_2363,N_824,N_331);
nor U2364 (N_2364,N_469,N_876);
nor U2365 (N_2365,N_1578,N_1711);
or U2366 (N_2366,N_1916,N_26);
and U2367 (N_2367,N_457,N_1594);
and U2368 (N_2368,N_602,N_1626);
and U2369 (N_2369,N_693,N_838);
or U2370 (N_2370,N_644,N_326);
and U2371 (N_2371,N_489,N_985);
nand U2372 (N_2372,N_1073,N_71);
nor U2373 (N_2373,N_1114,N_289);
and U2374 (N_2374,N_1120,N_928);
and U2375 (N_2375,N_755,N_857);
nand U2376 (N_2376,N_302,N_135);
nor U2377 (N_2377,N_1035,N_405);
and U2378 (N_2378,N_36,N_1979);
or U2379 (N_2379,N_104,N_1119);
nor U2380 (N_2380,N_1271,N_592);
nand U2381 (N_2381,N_443,N_1414);
or U2382 (N_2382,N_1927,N_1966);
and U2383 (N_2383,N_87,N_206);
and U2384 (N_2384,N_1932,N_743);
and U2385 (N_2385,N_127,N_1306);
nand U2386 (N_2386,N_1587,N_720);
or U2387 (N_2387,N_670,N_1952);
nand U2388 (N_2388,N_1498,N_77);
and U2389 (N_2389,N_1810,N_1032);
or U2390 (N_2390,N_1014,N_327);
nand U2391 (N_2391,N_335,N_56);
and U2392 (N_2392,N_998,N_1353);
or U2393 (N_2393,N_624,N_1557);
or U2394 (N_2394,N_353,N_1603);
xnor U2395 (N_2395,N_125,N_915);
nor U2396 (N_2396,N_511,N_393);
or U2397 (N_2397,N_37,N_41);
nor U2398 (N_2398,N_1242,N_1861);
xor U2399 (N_2399,N_820,N_1240);
and U2400 (N_2400,N_449,N_1515);
or U2401 (N_2401,N_1849,N_1552);
or U2402 (N_2402,N_515,N_1251);
nor U2403 (N_2403,N_1778,N_631);
nand U2404 (N_2404,N_106,N_355);
nand U2405 (N_2405,N_1221,N_365);
and U2406 (N_2406,N_272,N_543);
or U2407 (N_2407,N_1668,N_1981);
or U2408 (N_2408,N_687,N_683);
and U2409 (N_2409,N_975,N_770);
nor U2410 (N_2410,N_1698,N_1260);
or U2411 (N_2411,N_1189,N_52);
nand U2412 (N_2412,N_1723,N_1701);
and U2413 (N_2413,N_1190,N_283);
or U2414 (N_2414,N_635,N_686);
nand U2415 (N_2415,N_731,N_1025);
or U2416 (N_2416,N_1644,N_321);
nand U2417 (N_2417,N_659,N_1143);
and U2418 (N_2418,N_909,N_1300);
or U2419 (N_2419,N_637,N_536);
nand U2420 (N_2420,N_176,N_744);
and U2421 (N_2421,N_1217,N_1518);
nor U2422 (N_2422,N_1943,N_1968);
or U2423 (N_2423,N_1951,N_1478);
and U2424 (N_2424,N_10,N_1863);
nand U2425 (N_2425,N_128,N_1379);
and U2426 (N_2426,N_1774,N_1370);
and U2427 (N_2427,N_1346,N_1767);
nand U2428 (N_2428,N_1350,N_1537);
or U2429 (N_2429,N_284,N_521);
and U2430 (N_2430,N_661,N_1835);
nor U2431 (N_2431,N_1546,N_1864);
nor U2432 (N_2432,N_612,N_158);
nor U2433 (N_2433,N_750,N_1338);
or U2434 (N_2434,N_1879,N_1080);
nor U2435 (N_2435,N_401,N_1033);
nand U2436 (N_2436,N_1386,N_1771);
nand U2437 (N_2437,N_1915,N_518);
nand U2438 (N_2438,N_1176,N_371);
and U2439 (N_2439,N_599,N_1794);
and U2440 (N_2440,N_940,N_1907);
nand U2441 (N_2441,N_1367,N_1681);
nand U2442 (N_2442,N_1503,N_546);
nand U2443 (N_2443,N_1390,N_1102);
or U2444 (N_2444,N_490,N_566);
nor U2445 (N_2445,N_1811,N_517);
and U2446 (N_2446,N_399,N_473);
and U2447 (N_2447,N_789,N_1781);
nor U2448 (N_2448,N_1009,N_1577);
and U2449 (N_2449,N_1901,N_1899);
or U2450 (N_2450,N_298,N_262);
nor U2451 (N_2451,N_1199,N_17);
or U2452 (N_2452,N_1402,N_1099);
xnor U2453 (N_2453,N_1820,N_1001);
or U2454 (N_2454,N_1617,N_1570);
nand U2455 (N_2455,N_906,N_370);
nor U2456 (N_2456,N_39,N_1416);
nand U2457 (N_2457,N_430,N_1830);
and U2458 (N_2458,N_504,N_1775);
and U2459 (N_2459,N_1947,N_1345);
or U2460 (N_2460,N_668,N_943);
nor U2461 (N_2461,N_313,N_1648);
and U2462 (N_2462,N_1064,N_111);
nor U2463 (N_2463,N_80,N_1554);
nor U2464 (N_2464,N_200,N_1990);
or U2465 (N_2465,N_1130,N_549);
nor U2466 (N_2466,N_1933,N_1910);
nand U2467 (N_2467,N_545,N_497);
or U2468 (N_2468,N_764,N_1722);
nand U2469 (N_2469,N_1929,N_554);
nand U2470 (N_2470,N_16,N_782);
nand U2471 (N_2471,N_730,N_95);
nor U2472 (N_2472,N_1890,N_726);
nand U2473 (N_2473,N_1410,N_1112);
and U2474 (N_2474,N_583,N_1998);
or U2475 (N_2475,N_1453,N_548);
or U2476 (N_2476,N_191,N_1174);
nor U2477 (N_2477,N_316,N_1654);
nor U2478 (N_2478,N_1329,N_629);
or U2479 (N_2479,N_1435,N_934);
and U2480 (N_2480,N_814,N_715);
nor U2481 (N_2481,N_859,N_1077);
and U2482 (N_2482,N_500,N_942);
nand U2483 (N_2483,N_594,N_1618);
and U2484 (N_2484,N_1708,N_1156);
nor U2485 (N_2485,N_968,N_1054);
and U2486 (N_2486,N_1297,N_263);
nand U2487 (N_2487,N_1068,N_965);
and U2488 (N_2488,N_1280,N_1969);
and U2489 (N_2489,N_1764,N_530);
nor U2490 (N_2490,N_547,N_220);
nand U2491 (N_2491,N_47,N_479);
and U2492 (N_2492,N_174,N_1153);
and U2493 (N_2493,N_1924,N_1107);
and U2494 (N_2494,N_621,N_1134);
or U2495 (N_2495,N_1676,N_1539);
and U2496 (N_2496,N_839,N_207);
nor U2497 (N_2497,N_1342,N_21);
or U2498 (N_2498,N_1739,N_305);
nand U2499 (N_2499,N_462,N_1272);
nand U2500 (N_2500,N_787,N_9);
or U2501 (N_2501,N_1218,N_833);
nand U2502 (N_2502,N_291,N_1241);
nor U2503 (N_2503,N_1866,N_1475);
or U2504 (N_2504,N_1150,N_387);
and U2505 (N_2505,N_1823,N_710);
or U2506 (N_2506,N_1504,N_1625);
or U2507 (N_2507,N_790,N_442);
and U2508 (N_2508,N_455,N_1826);
and U2509 (N_2509,N_90,N_424);
or U2510 (N_2510,N_671,N_185);
nor U2511 (N_2511,N_297,N_1793);
nor U2512 (N_2512,N_734,N_1050);
and U2513 (N_2513,N_1556,N_1483);
nand U2514 (N_2514,N_794,N_1709);
and U2515 (N_2515,N_1683,N_195);
or U2516 (N_2516,N_1634,N_386);
and U2517 (N_2517,N_182,N_343);
nor U2518 (N_2518,N_1187,N_1286);
or U2519 (N_2519,N_266,N_516);
nand U2520 (N_2520,N_222,N_568);
and U2521 (N_2521,N_78,N_1309);
nor U2522 (N_2522,N_1016,N_193);
nor U2523 (N_2523,N_1196,N_837);
nor U2524 (N_2524,N_1749,N_1831);
nand U2525 (N_2525,N_1281,N_482);
nor U2526 (N_2526,N_1229,N_1431);
xnor U2527 (N_2527,N_432,N_433);
nand U2528 (N_2528,N_227,N_1039);
nand U2529 (N_2529,N_452,N_1308);
nand U2530 (N_2530,N_1182,N_801);
and U2531 (N_2531,N_1656,N_1982);
or U2532 (N_2532,N_1264,N_969);
nor U2533 (N_2533,N_1524,N_1959);
or U2534 (N_2534,N_1761,N_1397);
or U2535 (N_2535,N_769,N_798);
and U2536 (N_2536,N_65,N_795);
nand U2537 (N_2537,N_416,N_382);
nor U2538 (N_2538,N_1946,N_1805);
nor U2539 (N_2539,N_1349,N_1457);
nand U2540 (N_2540,N_563,N_520);
nand U2541 (N_2541,N_895,N_1029);
nor U2542 (N_2542,N_1135,N_717);
or U2543 (N_2543,N_1930,N_1886);
nor U2544 (N_2544,N_1420,N_1259);
or U2545 (N_2545,N_1352,N_1652);
xor U2546 (N_2546,N_1364,N_1581);
and U2547 (N_2547,N_1986,N_1034);
and U2548 (N_2548,N_585,N_1184);
and U2549 (N_2549,N_1938,N_800);
or U2550 (N_2550,N_444,N_43);
or U2551 (N_2551,N_352,N_1327);
nand U2552 (N_2552,N_1833,N_936);
and U2553 (N_2553,N_1750,N_825);
nor U2554 (N_2554,N_913,N_1095);
or U2555 (N_2555,N_535,N_1891);
nor U2556 (N_2556,N_625,N_555);
or U2557 (N_2557,N_944,N_1393);
nor U2558 (N_2558,N_34,N_1547);
and U2559 (N_2559,N_1248,N_1939);
nand U2560 (N_2560,N_1028,N_441);
and U2561 (N_2561,N_336,N_907);
nand U2562 (N_2562,N_1111,N_1619);
nand U2563 (N_2563,N_1278,N_863);
nor U2564 (N_2564,N_1225,N_120);
and U2565 (N_2565,N_494,N_922);
or U2566 (N_2566,N_244,N_1731);
and U2567 (N_2567,N_999,N_380);
or U2568 (N_2568,N_1284,N_1465);
nand U2569 (N_2569,N_234,N_630);
and U2570 (N_2570,N_505,N_1961);
and U2571 (N_2571,N_561,N_1006);
nor U2572 (N_2572,N_753,N_1841);
nor U2573 (N_2573,N_404,N_1522);
or U2574 (N_2574,N_1784,N_42);
and U2575 (N_2575,N_689,N_990);
xor U2576 (N_2576,N_1279,N_1906);
or U2577 (N_2577,N_1213,N_851);
and U2578 (N_2578,N_1869,N_912);
nor U2579 (N_2579,N_1900,N_729);
or U2580 (N_2580,N_791,N_1396);
nor U2581 (N_2581,N_704,N_46);
and U2582 (N_2582,N_1128,N_412);
nand U2583 (N_2583,N_154,N_1870);
or U2584 (N_2584,N_961,N_1056);
and U2585 (N_2585,N_1640,N_1089);
nand U2586 (N_2586,N_1314,N_208);
nand U2587 (N_2587,N_1070,N_364);
and U2588 (N_2588,N_245,N_1674);
or U2589 (N_2589,N_580,N_551);
nand U2590 (N_2590,N_58,N_528);
and U2591 (N_2591,N_819,N_1741);
or U2592 (N_2592,N_1735,N_50);
or U2593 (N_2593,N_579,N_861);
or U2594 (N_2594,N_1738,N_1315);
nor U2595 (N_2595,N_344,N_53);
nor U2596 (N_2596,N_956,N_1516);
or U2597 (N_2597,N_1903,N_1526);
nor U2598 (N_2598,N_925,N_175);
nor U2599 (N_2599,N_340,N_1490);
and U2600 (N_2600,N_1868,N_166);
nand U2601 (N_2601,N_1152,N_1779);
and U2602 (N_2602,N_804,N_946);
and U2603 (N_2603,N_902,N_403);
and U2604 (N_2604,N_974,N_864);
and U2605 (N_2605,N_1743,N_685);
xor U2606 (N_2606,N_565,N_1746);
and U2607 (N_2607,N_526,N_199);
nor U2608 (N_2608,N_1269,N_149);
or U2609 (N_2609,N_1919,N_447);
and U2610 (N_2610,N_38,N_64);
or U2611 (N_2611,N_1261,N_1484);
nor U2612 (N_2612,N_1263,N_1211);
or U2613 (N_2613,N_1985,N_1206);
and U2614 (N_2614,N_1993,N_1935);
or U2615 (N_2615,N_1983,N_35);
nand U2616 (N_2616,N_453,N_1324);
or U2617 (N_2617,N_774,N_1517);
nor U2618 (N_2618,N_638,N_994);
and U2619 (N_2619,N_916,N_165);
or U2620 (N_2620,N_1026,N_847);
nor U2621 (N_2621,N_529,N_122);
and U2622 (N_2622,N_392,N_1673);
nor U2623 (N_2623,N_1277,N_1012);
nor U2624 (N_2624,N_1666,N_357);
nand U2625 (N_2625,N_811,N_508);
and U2626 (N_2626,N_196,N_642);
or U2627 (N_2627,N_1842,N_346);
and U2628 (N_2628,N_268,N_841);
xor U2629 (N_2629,N_445,N_1973);
nor U2630 (N_2630,N_1511,N_1162);
and U2631 (N_2631,N_560,N_559);
nor U2632 (N_2632,N_850,N_1599);
nor U2633 (N_2633,N_1455,N_1471);
and U2634 (N_2634,N_1048,N_853);
nand U2635 (N_2635,N_589,N_61);
nand U2636 (N_2636,N_436,N_848);
and U2637 (N_2637,N_1745,N_1984);
nor U2638 (N_2638,N_1454,N_1975);
nor U2639 (N_2639,N_391,N_1780);
nand U2640 (N_2640,N_897,N_159);
nand U2641 (N_2641,N_763,N_955);
nor U2642 (N_2642,N_243,N_92);
or U2643 (N_2643,N_1592,N_330);
nor U2644 (N_2644,N_1469,N_1194);
and U2645 (N_2645,N_678,N_948);
and U2646 (N_2646,N_977,N_608);
and U2647 (N_2647,N_766,N_232);
or U2648 (N_2648,N_1719,N_296);
or U2649 (N_2649,N_1694,N_655);
nor U2650 (N_2650,N_1655,N_1154);
or U2651 (N_2651,N_468,N_1139);
nand U2652 (N_2652,N_1705,N_114);
and U2653 (N_2653,N_911,N_1142);
nand U2654 (N_2654,N_194,N_901);
nand U2655 (N_2655,N_2,N_372);
nand U2656 (N_2656,N_1721,N_259);
nor U2657 (N_2657,N_1660,N_231);
nand U2658 (N_2658,N_1834,N_44);
xor U2659 (N_2659,N_1098,N_270);
or U2660 (N_2660,N_600,N_779);
nor U2661 (N_2661,N_1977,N_395);
and U2662 (N_2662,N_1908,N_1395);
nand U2663 (N_2663,N_318,N_971);
nand U2664 (N_2664,N_66,N_1330);
and U2665 (N_2665,N_257,N_1210);
nand U2666 (N_2666,N_267,N_1433);
or U2667 (N_2667,N_677,N_1331);
and U2668 (N_2668,N_1641,N_540);
nand U2669 (N_2669,N_1845,N_88);
nor U2670 (N_2670,N_1837,N_1045);
xnor U2671 (N_2671,N_835,N_324);
nor U2672 (N_2672,N_478,N_73);
and U2673 (N_2673,N_1801,N_1921);
nand U2674 (N_2674,N_596,N_1185);
or U2675 (N_2675,N_1814,N_564);
and U2676 (N_2676,N_885,N_581);
and U2677 (N_2677,N_1732,N_1693);
and U2678 (N_2678,N_1188,N_1274);
nor U2679 (N_2679,N_1380,N_628);
nor U2680 (N_2680,N_1155,N_1535);
and U2681 (N_2681,N_1158,N_1677);
nor U2682 (N_2682,N_714,N_1827);
nand U2683 (N_2683,N_1103,N_696);
nand U2684 (N_2684,N_1057,N_1389);
or U2685 (N_2685,N_1101,N_1531);
nor U2686 (N_2686,N_1421,N_1236);
and U2687 (N_2687,N_1550,N_703);
and U2688 (N_2688,N_337,N_45);
nor U2689 (N_2689,N_1591,N_883);
nor U2690 (N_2690,N_1177,N_79);
and U2691 (N_2691,N_904,N_121);
or U2692 (N_2692,N_1293,N_1855);
and U2693 (N_2693,N_1881,N_1138);
nand U2694 (N_2694,N_315,N_354);
nor U2695 (N_2695,N_1730,N_105);
nor U2696 (N_2696,N_1096,N_933);
or U2697 (N_2697,N_8,N_138);
and U2698 (N_2698,N_1198,N_1710);
and U2699 (N_2699,N_201,N_1159);
and U2700 (N_2700,N_626,N_1149);
nand U2701 (N_2701,N_1419,N_319);
and U2702 (N_2702,N_369,N_1822);
nor U2703 (N_2703,N_1294,N_1398);
nand U2704 (N_2704,N_481,N_1851);
and U2705 (N_2705,N_611,N_1328);
nor U2706 (N_2706,N_1004,N_1748);
nand U2707 (N_2707,N_411,N_918);
and U2708 (N_2708,N_512,N_1450);
or U2709 (N_2709,N_1161,N_1104);
or U2710 (N_2710,N_1121,N_1239);
nand U2711 (N_2711,N_1832,N_141);
and U2712 (N_2712,N_67,N_1529);
and U2713 (N_2713,N_1859,N_209);
nand U2714 (N_2714,N_652,N_1036);
nor U2715 (N_2715,N_211,N_1804);
or U2716 (N_2716,N_607,N_5);
and U2717 (N_2717,N_1041,N_691);
or U2718 (N_2718,N_1876,N_1227);
or U2719 (N_2719,N_1131,N_1167);
nor U2720 (N_2720,N_1871,N_1093);
nor U2721 (N_2721,N_1878,N_358);
nand U2722 (N_2722,N_684,N_314);
and U2723 (N_2723,N_219,N_1336);
or U2724 (N_2724,N_634,N_553);
or U2725 (N_2725,N_868,N_1846);
and U2726 (N_2726,N_261,N_586);
nor U2727 (N_2727,N_329,N_1964);
nand U2728 (N_2728,N_1737,N_765);
nand U2729 (N_2729,N_1166,N_1839);
nor U2730 (N_2730,N_328,N_582);
and U2731 (N_2731,N_1434,N_788);
nand U2732 (N_2732,N_1788,N_1388);
or U2733 (N_2733,N_1609,N_1105);
or U2734 (N_2734,N_1059,N_617);
or U2735 (N_2735,N_1375,N_694);
or U2736 (N_2736,N_1087,N_1432);
nor U2737 (N_2737,N_82,N_1289);
nand U2738 (N_2738,N_761,N_1512);
and U2739 (N_2739,N_927,N_230);
nor U2740 (N_2740,N_827,N_1253);
nor U2741 (N_2741,N_124,N_695);
nand U2742 (N_2742,N_1497,N_1052);
or U2743 (N_2743,N_1978,N_1051);
nand U2744 (N_2744,N_273,N_919);
nor U2745 (N_2745,N_183,N_1024);
nand U2746 (N_2746,N_1659,N_1005);
nor U2747 (N_2747,N_213,N_780);
or U2748 (N_2748,N_1326,N_759);
nand U2749 (N_2749,N_1060,N_1254);
or U2750 (N_2750,N_1019,N_613);
nand U2751 (N_2751,N_1520,N_474);
and U2752 (N_2752,N_1912,N_1695);
or U2753 (N_2753,N_1604,N_991);
nor U2754 (N_2754,N_1953,N_1084);
nand U2755 (N_2755,N_451,N_435);
and U2756 (N_2756,N_7,N_1671);
and U2757 (N_2757,N_1665,N_757);
and U2758 (N_2758,N_1231,N_414);
nor U2759 (N_2759,N_1593,N_83);
xnor U2760 (N_2760,N_1797,N_1662);
or U2761 (N_2761,N_178,N_1204);
and U2762 (N_2762,N_1351,N_1023);
or U2763 (N_2763,N_1815,N_1061);
nand U2764 (N_2764,N_1219,N_1374);
nor U2765 (N_2765,N_1995,N_1647);
nand U2766 (N_2766,N_247,N_1917);
nand U2767 (N_2767,N_1479,N_1079);
or U2768 (N_2768,N_641,N_1926);
nor U2769 (N_2769,N_632,N_1106);
nor U2770 (N_2770,N_1423,N_1680);
or U2771 (N_2771,N_425,N_1562);
nor U2772 (N_2772,N_1394,N_1110);
nor U2773 (N_2773,N_1970,N_249);
nand U2774 (N_2774,N_1125,N_186);
nor U2775 (N_2775,N_1317,N_793);
nand U2776 (N_2776,N_320,N_1148);
or U2777 (N_2777,N_855,N_501);
and U2778 (N_2778,N_496,N_645);
and U2779 (N_2779,N_306,N_471);
or U2780 (N_2780,N_98,N_648);
nor U2781 (N_2781,N_1292,N_407);
nand U2782 (N_2782,N_899,N_1699);
nand U2783 (N_2783,N_170,N_810);
nor U2784 (N_2784,N_1777,N_879);
nor U2785 (N_2785,N_304,N_112);
nand U2786 (N_2786,N_282,N_799);
nor U2787 (N_2787,N_603,N_996);
nand U2788 (N_2788,N_679,N_1316);
or U2789 (N_2789,N_1895,N_920);
nand U2790 (N_2790,N_1027,N_1532);
and U2791 (N_2791,N_1097,N_1765);
and U2792 (N_2792,N_1569,N_830);
or U2793 (N_2793,N_1667,N_373);
nand U2794 (N_2794,N_419,N_643);
and U2795 (N_2795,N_663,N_1304);
nand U2796 (N_2796,N_434,N_1760);
and U2797 (N_2797,N_102,N_1770);
and U2798 (N_2798,N_593,N_1684);
or U2799 (N_2799,N_1262,N_145);
and U2800 (N_2800,N_1558,N_1559);
nor U2801 (N_2801,N_886,N_775);
nand U2802 (N_2802,N_1848,N_1696);
or U2803 (N_2803,N_1590,N_1487);
nand U2804 (N_2804,N_889,N_619);
or U2805 (N_2805,N_1062,N_552);
nand U2806 (N_2806,N_1560,N_1146);
or U2807 (N_2807,N_926,N_1302);
and U2808 (N_2808,N_1071,N_1245);
and U2809 (N_2809,N_1689,N_989);
xor U2810 (N_2810,N_1208,N_1486);
and U2811 (N_2811,N_524,N_1541);
or U2812 (N_2812,N_1954,N_1237);
nor U2813 (N_2813,N_877,N_1551);
nor U2814 (N_2814,N_271,N_1323);
nand U2815 (N_2815,N_240,N_1305);
or U2816 (N_2816,N_123,N_269);
nor U2817 (N_2817,N_1941,N_1282);
nor U2818 (N_2818,N_1543,N_254);
or U2819 (N_2819,N_383,N_1766);
nand U2820 (N_2820,N_1488,N_1451);
nand U2821 (N_2821,N_1650,N_807);
or U2822 (N_2822,N_776,N_1439);
or U2823 (N_2823,N_572,N_1754);
nor U2824 (N_2824,N_1865,N_1318);
and U2825 (N_2825,N_1755,N_1565);
and U2826 (N_2826,N_1247,N_334);
nor U2827 (N_2827,N_1702,N_1460);
and U2828 (N_2828,N_1847,N_1853);
nand U2829 (N_2829,N_1948,N_101);
nor U2830 (N_2830,N_152,N_385);
nor U2831 (N_2831,N_1686,N_1347);
nor U2832 (N_2832,N_1679,N_1806);
nor U2833 (N_2833,N_713,N_1756);
nand U2834 (N_2834,N_1636,N_923);
and U2835 (N_2835,N_615,N_1753);
nand U2836 (N_2836,N_1255,N_945);
and U2837 (N_2837,N_86,N_711);
or U2838 (N_2838,N_570,N_59);
or U2839 (N_2839,N_962,N_682);
and U2840 (N_2840,N_161,N_941);
and U2841 (N_2841,N_1082,N_1046);
and U2842 (N_2842,N_976,N_576);
or U2843 (N_2843,N_680,N_1690);
or U2844 (N_2844,N_1461,N_896);
nor U2845 (N_2845,N_1862,N_390);
nand U2846 (N_2846,N_250,N_1795);
nand U2847 (N_2847,N_63,N_760);
or U2848 (N_2848,N_917,N_1949);
nand U2849 (N_2849,N_647,N_742);
and U2850 (N_2850,N_264,N_1069);
and U2851 (N_2851,N_1372,N_440);
or U2852 (N_2852,N_431,N_1320);
nand U2853 (N_2853,N_1002,N_317);
nand U2854 (N_2854,N_1828,N_527);
and U2855 (N_2855,N_1296,N_832);
and U2856 (N_2856,N_1337,N_1630);
nor U2857 (N_2857,N_1090,N_1141);
or U2858 (N_2858,N_1530,N_1836);
nor U2859 (N_2859,N_1366,N_32);
nand U2860 (N_2860,N_448,N_772);
nor U2861 (N_2861,N_1960,N_427);
and U2862 (N_2862,N_110,N_537);
and U2863 (N_2863,N_1962,N_1944);
nor U2864 (N_2864,N_1493,N_654);
nand U2865 (N_2865,N_544,N_1600);
or U2866 (N_2866,N_1607,N_1682);
nor U2867 (N_2867,N_163,N_953);
and U2868 (N_2868,N_1514,N_1429);
or U2869 (N_2869,N_1653,N_1409);
or U2870 (N_2870,N_845,N_973);
nand U2871 (N_2871,N_139,N_1615);
nor U2872 (N_2872,N_216,N_618);
and U2873 (N_2873,N_1181,N_1209);
and U2874 (N_2874,N_1718,N_898);
and U2875 (N_2875,N_950,N_1918);
nand U2876 (N_2876,N_374,N_461);
nor U2877 (N_2877,N_1017,N_1584);
or U2878 (N_2878,N_225,N_1887);
nand U2879 (N_2879,N_1687,N_849);
or U2880 (N_2880,N_258,N_1999);
nand U2881 (N_2881,N_519,N_398);
and U2882 (N_2882,N_147,N_1011);
nand U2883 (N_2883,N_115,N_1873);
or U2884 (N_2884,N_94,N_1436);
nand U2885 (N_2885,N_1575,N_1343);
nor U2886 (N_2886,N_1544,N_1720);
nand U2887 (N_2887,N_698,N_242);
or U2888 (N_2888,N_1642,N_223);
nand U2889 (N_2889,N_1980,N_1534);
nor U2890 (N_2890,N_900,N_662);
and U2891 (N_2891,N_1583,N_1117);
nand U2892 (N_2892,N_1031,N_1230);
or U2893 (N_2893,N_1840,N_60);
xnor U2894 (N_2894,N_129,N_421);
and U2895 (N_2895,N_821,N_180);
or U2896 (N_2896,N_736,N_1624);
or U2897 (N_2897,N_466,N_389);
and U2898 (N_2898,N_1989,N_1807);
nand U2899 (N_2899,N_723,N_1538);
nor U2900 (N_2900,N_1,N_584);
nor U2901 (N_2901,N_1216,N_1445);
nand U2902 (N_2902,N_1250,N_130);
or U2903 (N_2903,N_888,N_1509);
nand U2904 (N_2904,N_198,N_531);
or U2905 (N_2905,N_1657,N_636);
or U2906 (N_2906,N_980,N_777);
nand U2907 (N_2907,N_1561,N_164);
and U2908 (N_2908,N_817,N_1611);
nand U2909 (N_2909,N_1596,N_126);
nand U2910 (N_2910,N_1458,N_1854);
nand U2911 (N_2911,N_812,N_1726);
nand U2912 (N_2912,N_1441,N_113);
nor U2913 (N_2913,N_1725,N_1413);
and U2914 (N_2914,N_1894,N_1633);
nand U2915 (N_2915,N_109,N_1437);
nand U2916 (N_2916,N_1392,N_854);
nand U2917 (N_2917,N_805,N_235);
and U2918 (N_2918,N_1816,N_423);
or U2919 (N_2919,N_667,N_1468);
nand U2920 (N_2920,N_1298,N_893);
nor U2921 (N_2921,N_1582,N_233);
and U2922 (N_2922,N_903,N_997);
or U2923 (N_2923,N_882,N_1412);
or U2924 (N_2924,N_1651,N_1083);
and U2925 (N_2925,N_858,N_322);
nor U2926 (N_2926,N_978,N_460);
and U2927 (N_2927,N_1267,N_375);
xor U2928 (N_2928,N_1171,N_1632);
or U2929 (N_2929,N_1387,N_1232);
nand U2930 (N_2930,N_1170,N_1787);
and U2931 (N_2931,N_91,N_1168);
nor U2932 (N_2932,N_169,N_1678);
nor U2933 (N_2933,N_487,N_1825);
nand U2934 (N_2934,N_119,N_1133);
nand U2935 (N_2935,N_598,N_1124);
or U2936 (N_2936,N_255,N_722);
nand U2937 (N_2937,N_1425,N_1178);
xor U2938 (N_2938,N_25,N_1508);
nand U2939 (N_2939,N_1123,N_1523);
nor U2940 (N_2940,N_228,N_1857);
or U2941 (N_2941,N_1440,N_12);
and U2942 (N_2942,N_1786,N_100);
nand U2943 (N_2943,N_1506,N_751);
nor U2944 (N_2944,N_963,N_1496);
nand U2945 (N_2945,N_890,N_116);
or U2946 (N_2946,N_1585,N_409);
or U2947 (N_2947,N_986,N_76);
and U2948 (N_2948,N_1193,N_653);
or U2949 (N_2949,N_1976,N_1940);
or U2950 (N_2950,N_1945,N_278);
and U2951 (N_2951,N_1234,N_1092);
nand U2952 (N_2952,N_359,N_288);
nand U2953 (N_2953,N_1605,N_1796);
nor U2954 (N_2954,N_1507,N_300);
and U2955 (N_2955,N_1860,N_74);
and U2956 (N_2956,N_68,N_1955);
nand U2957 (N_2957,N_137,N_707);
and U2958 (N_2958,N_1889,N_275);
xor U2959 (N_2959,N_177,N_1553);
and U2960 (N_2960,N_818,N_1422);
or U2961 (N_2961,N_1220,N_1491);
and U2962 (N_2962,N_493,N_1173);
nor U2963 (N_2963,N_816,N_1108);
and U2964 (N_2964,N_1163,N_842);
nand U2965 (N_2965,N_605,N_622);
or U2966 (N_2966,N_1747,N_1022);
nand U2967 (N_2967,N_467,N_218);
xor U2968 (N_2968,N_420,N_356);
nand U2969 (N_2969,N_620,N_1311);
or U2970 (N_2970,N_96,N_142);
or U2971 (N_2971,N_706,N_1800);
nand U2972 (N_2972,N_981,N_510);
and U2973 (N_2973,N_1713,N_993);
or U2974 (N_2974,N_709,N_1843);
or U2975 (N_2975,N_1790,N_856);
nand U2976 (N_2976,N_1628,N_187);
nand U2977 (N_2977,N_1638,N_480);
or U2978 (N_2978,N_24,N_822);
and U2979 (N_2979,N_1965,N_1186);
nand U2980 (N_2980,N_1934,N_1758);
or U2981 (N_2981,N_1649,N_1589);
and U2982 (N_2982,N_797,N_513);
nand U2983 (N_2983,N_702,N_1066);
or U2984 (N_2984,N_697,N_1449);
and U2985 (N_2985,N_891,N_1020);
nand U2986 (N_2986,N_1542,N_1480);
nor U2987 (N_2987,N_786,N_571);
nor U2988 (N_2988,N_1897,N_333);
or U2989 (N_2989,N_1481,N_1348);
and U2990 (N_2990,N_1126,N_40);
or U2991 (N_2991,N_836,N_1470);
nor U2992 (N_2992,N_361,N_1555);
and U2993 (N_2993,N_1013,N_532);
nor U2994 (N_2994,N_972,N_746);
and U2995 (N_2995,N_1290,N_286);
or U2996 (N_2996,N_28,N_887);
or U2997 (N_2997,N_1466,N_81);
nand U2998 (N_2998,N_1716,N_428);
nor U2999 (N_2999,N_151,N_525);
nor U3000 (N_3000,N_659,N_1458);
nand U3001 (N_3001,N_1136,N_1041);
nand U3002 (N_3002,N_1129,N_390);
nor U3003 (N_3003,N_164,N_934);
and U3004 (N_3004,N_1185,N_1023);
nand U3005 (N_3005,N_1247,N_1090);
or U3006 (N_3006,N_845,N_1578);
nor U3007 (N_3007,N_1693,N_1796);
nand U3008 (N_3008,N_1008,N_1649);
and U3009 (N_3009,N_713,N_199);
nor U3010 (N_3010,N_1037,N_1611);
nor U3011 (N_3011,N_1594,N_1667);
or U3012 (N_3012,N_1183,N_1832);
nor U3013 (N_3013,N_580,N_83);
and U3014 (N_3014,N_65,N_1372);
or U3015 (N_3015,N_1603,N_795);
and U3016 (N_3016,N_1760,N_1580);
or U3017 (N_3017,N_1848,N_1633);
or U3018 (N_3018,N_197,N_1305);
nand U3019 (N_3019,N_1173,N_1273);
or U3020 (N_3020,N_1902,N_1733);
nand U3021 (N_3021,N_585,N_1119);
nand U3022 (N_3022,N_346,N_4);
or U3023 (N_3023,N_1725,N_1442);
nor U3024 (N_3024,N_542,N_1802);
or U3025 (N_3025,N_658,N_747);
nand U3026 (N_3026,N_886,N_1580);
nand U3027 (N_3027,N_1370,N_1445);
nand U3028 (N_3028,N_1725,N_1550);
nor U3029 (N_3029,N_1086,N_1414);
or U3030 (N_3030,N_1412,N_1619);
nand U3031 (N_3031,N_847,N_780);
nor U3032 (N_3032,N_931,N_1217);
nor U3033 (N_3033,N_155,N_104);
xor U3034 (N_3034,N_1343,N_1814);
nand U3035 (N_3035,N_1410,N_229);
or U3036 (N_3036,N_1919,N_1600);
or U3037 (N_3037,N_1657,N_89);
nand U3038 (N_3038,N_1684,N_220);
nand U3039 (N_3039,N_903,N_192);
nor U3040 (N_3040,N_1959,N_868);
nand U3041 (N_3041,N_1702,N_869);
nand U3042 (N_3042,N_832,N_862);
and U3043 (N_3043,N_126,N_1823);
xor U3044 (N_3044,N_1125,N_1827);
or U3045 (N_3045,N_947,N_148);
or U3046 (N_3046,N_1003,N_1834);
nor U3047 (N_3047,N_841,N_1775);
and U3048 (N_3048,N_837,N_1581);
nand U3049 (N_3049,N_1600,N_436);
nor U3050 (N_3050,N_417,N_1840);
and U3051 (N_3051,N_422,N_943);
or U3052 (N_3052,N_1370,N_556);
and U3053 (N_3053,N_1156,N_1434);
and U3054 (N_3054,N_162,N_73);
and U3055 (N_3055,N_1288,N_841);
and U3056 (N_3056,N_1859,N_918);
and U3057 (N_3057,N_1040,N_1104);
nor U3058 (N_3058,N_1519,N_497);
nand U3059 (N_3059,N_1957,N_1000);
nand U3060 (N_3060,N_1679,N_308);
and U3061 (N_3061,N_630,N_685);
or U3062 (N_3062,N_533,N_1998);
or U3063 (N_3063,N_554,N_578);
nor U3064 (N_3064,N_1984,N_581);
or U3065 (N_3065,N_252,N_352);
nand U3066 (N_3066,N_1213,N_51);
nand U3067 (N_3067,N_1973,N_1243);
or U3068 (N_3068,N_1558,N_291);
nand U3069 (N_3069,N_56,N_315);
or U3070 (N_3070,N_1106,N_921);
or U3071 (N_3071,N_16,N_370);
or U3072 (N_3072,N_132,N_833);
nand U3073 (N_3073,N_1584,N_662);
nor U3074 (N_3074,N_457,N_926);
and U3075 (N_3075,N_1840,N_1039);
nor U3076 (N_3076,N_1417,N_1649);
nand U3077 (N_3077,N_1903,N_1813);
nand U3078 (N_3078,N_866,N_1356);
and U3079 (N_3079,N_1758,N_1157);
and U3080 (N_3080,N_1250,N_1118);
nor U3081 (N_3081,N_81,N_1086);
or U3082 (N_3082,N_132,N_972);
nor U3083 (N_3083,N_1981,N_1951);
nand U3084 (N_3084,N_415,N_883);
nand U3085 (N_3085,N_474,N_81);
nor U3086 (N_3086,N_695,N_982);
or U3087 (N_3087,N_1126,N_936);
or U3088 (N_3088,N_1689,N_1082);
or U3089 (N_3089,N_489,N_31);
nand U3090 (N_3090,N_286,N_1768);
and U3091 (N_3091,N_844,N_1603);
nand U3092 (N_3092,N_992,N_416);
or U3093 (N_3093,N_457,N_1770);
and U3094 (N_3094,N_1881,N_646);
nor U3095 (N_3095,N_1170,N_234);
or U3096 (N_3096,N_1603,N_650);
and U3097 (N_3097,N_1299,N_1486);
or U3098 (N_3098,N_1411,N_1945);
nand U3099 (N_3099,N_677,N_569);
or U3100 (N_3100,N_162,N_1485);
or U3101 (N_3101,N_1466,N_1735);
and U3102 (N_3102,N_928,N_211);
nor U3103 (N_3103,N_1961,N_460);
and U3104 (N_3104,N_1127,N_1220);
or U3105 (N_3105,N_1009,N_1088);
or U3106 (N_3106,N_984,N_1400);
or U3107 (N_3107,N_512,N_1751);
nor U3108 (N_3108,N_1374,N_1117);
xnor U3109 (N_3109,N_3,N_609);
or U3110 (N_3110,N_1534,N_1835);
or U3111 (N_3111,N_1813,N_1707);
nor U3112 (N_3112,N_1194,N_1363);
nand U3113 (N_3113,N_692,N_1047);
and U3114 (N_3114,N_255,N_244);
xor U3115 (N_3115,N_321,N_974);
and U3116 (N_3116,N_453,N_871);
nor U3117 (N_3117,N_1726,N_1380);
xnor U3118 (N_3118,N_1942,N_1756);
nand U3119 (N_3119,N_1666,N_816);
nor U3120 (N_3120,N_497,N_314);
nor U3121 (N_3121,N_1555,N_1218);
and U3122 (N_3122,N_1496,N_1830);
and U3123 (N_3123,N_232,N_257);
and U3124 (N_3124,N_1545,N_112);
or U3125 (N_3125,N_1442,N_592);
or U3126 (N_3126,N_124,N_410);
and U3127 (N_3127,N_1117,N_550);
xnor U3128 (N_3128,N_1217,N_1702);
nor U3129 (N_3129,N_169,N_1679);
nand U3130 (N_3130,N_1034,N_365);
and U3131 (N_3131,N_1248,N_667);
nand U3132 (N_3132,N_148,N_174);
and U3133 (N_3133,N_1714,N_1528);
and U3134 (N_3134,N_1116,N_1415);
or U3135 (N_3135,N_1816,N_708);
nand U3136 (N_3136,N_1118,N_1626);
nor U3137 (N_3137,N_1243,N_1847);
nor U3138 (N_3138,N_940,N_1418);
nand U3139 (N_3139,N_1242,N_1604);
nor U3140 (N_3140,N_526,N_252);
nor U3141 (N_3141,N_1714,N_1156);
nor U3142 (N_3142,N_1112,N_1927);
nor U3143 (N_3143,N_577,N_110);
nor U3144 (N_3144,N_1052,N_1007);
nand U3145 (N_3145,N_669,N_429);
nor U3146 (N_3146,N_1584,N_269);
and U3147 (N_3147,N_1274,N_1307);
or U3148 (N_3148,N_1094,N_1412);
and U3149 (N_3149,N_1411,N_833);
nor U3150 (N_3150,N_52,N_601);
and U3151 (N_3151,N_1876,N_1547);
nor U3152 (N_3152,N_27,N_296);
nor U3153 (N_3153,N_1568,N_841);
nor U3154 (N_3154,N_994,N_967);
or U3155 (N_3155,N_1868,N_222);
nor U3156 (N_3156,N_287,N_1164);
nor U3157 (N_3157,N_283,N_324);
or U3158 (N_3158,N_1556,N_849);
or U3159 (N_3159,N_1481,N_942);
or U3160 (N_3160,N_1913,N_428);
nand U3161 (N_3161,N_1124,N_1731);
nor U3162 (N_3162,N_236,N_1408);
or U3163 (N_3163,N_825,N_49);
or U3164 (N_3164,N_281,N_406);
and U3165 (N_3165,N_832,N_1881);
nand U3166 (N_3166,N_1390,N_453);
and U3167 (N_3167,N_898,N_1472);
nand U3168 (N_3168,N_831,N_1291);
or U3169 (N_3169,N_1155,N_1708);
nor U3170 (N_3170,N_444,N_1692);
or U3171 (N_3171,N_1395,N_1415);
or U3172 (N_3172,N_1833,N_1976);
or U3173 (N_3173,N_1900,N_813);
and U3174 (N_3174,N_1480,N_1617);
nand U3175 (N_3175,N_887,N_105);
or U3176 (N_3176,N_1687,N_1906);
nand U3177 (N_3177,N_1518,N_516);
or U3178 (N_3178,N_1780,N_781);
or U3179 (N_3179,N_1091,N_324);
nor U3180 (N_3180,N_1668,N_1963);
and U3181 (N_3181,N_1641,N_1893);
or U3182 (N_3182,N_573,N_618);
and U3183 (N_3183,N_777,N_1908);
xnor U3184 (N_3184,N_138,N_1284);
nor U3185 (N_3185,N_909,N_1191);
nand U3186 (N_3186,N_556,N_655);
nand U3187 (N_3187,N_883,N_41);
and U3188 (N_3188,N_846,N_451);
nor U3189 (N_3189,N_1777,N_909);
or U3190 (N_3190,N_1656,N_1891);
nor U3191 (N_3191,N_92,N_1626);
nand U3192 (N_3192,N_1019,N_411);
nor U3193 (N_3193,N_1063,N_47);
and U3194 (N_3194,N_1202,N_344);
or U3195 (N_3195,N_485,N_1631);
or U3196 (N_3196,N_191,N_1464);
and U3197 (N_3197,N_243,N_1551);
nor U3198 (N_3198,N_1192,N_318);
nand U3199 (N_3199,N_839,N_519);
nand U3200 (N_3200,N_854,N_819);
nor U3201 (N_3201,N_83,N_424);
and U3202 (N_3202,N_1575,N_1573);
nor U3203 (N_3203,N_740,N_282);
nor U3204 (N_3204,N_509,N_1190);
and U3205 (N_3205,N_711,N_324);
or U3206 (N_3206,N_1526,N_252);
nor U3207 (N_3207,N_1150,N_208);
nor U3208 (N_3208,N_1883,N_1043);
and U3209 (N_3209,N_553,N_1725);
nor U3210 (N_3210,N_989,N_1336);
or U3211 (N_3211,N_1847,N_618);
nand U3212 (N_3212,N_492,N_1231);
nor U3213 (N_3213,N_559,N_840);
and U3214 (N_3214,N_1792,N_1576);
nor U3215 (N_3215,N_931,N_1911);
nor U3216 (N_3216,N_420,N_1766);
nand U3217 (N_3217,N_1042,N_961);
and U3218 (N_3218,N_602,N_103);
nand U3219 (N_3219,N_1242,N_1330);
nand U3220 (N_3220,N_824,N_1);
and U3221 (N_3221,N_1315,N_681);
or U3222 (N_3222,N_1691,N_1926);
or U3223 (N_3223,N_258,N_269);
nor U3224 (N_3224,N_348,N_613);
and U3225 (N_3225,N_442,N_729);
and U3226 (N_3226,N_1195,N_974);
and U3227 (N_3227,N_1263,N_1200);
nor U3228 (N_3228,N_1597,N_198);
nor U3229 (N_3229,N_973,N_79);
or U3230 (N_3230,N_1254,N_1265);
nor U3231 (N_3231,N_886,N_1230);
or U3232 (N_3232,N_1693,N_1125);
nand U3233 (N_3233,N_18,N_1901);
or U3234 (N_3234,N_1418,N_272);
nor U3235 (N_3235,N_1147,N_664);
and U3236 (N_3236,N_672,N_1539);
and U3237 (N_3237,N_213,N_787);
or U3238 (N_3238,N_1231,N_1323);
or U3239 (N_3239,N_791,N_728);
nor U3240 (N_3240,N_10,N_296);
nor U3241 (N_3241,N_1088,N_378);
and U3242 (N_3242,N_709,N_654);
or U3243 (N_3243,N_1758,N_260);
or U3244 (N_3244,N_1457,N_433);
nand U3245 (N_3245,N_113,N_432);
or U3246 (N_3246,N_492,N_17);
nor U3247 (N_3247,N_1926,N_476);
and U3248 (N_3248,N_686,N_312);
nor U3249 (N_3249,N_857,N_1177);
xor U3250 (N_3250,N_1053,N_1148);
nand U3251 (N_3251,N_472,N_928);
or U3252 (N_3252,N_355,N_689);
and U3253 (N_3253,N_264,N_1445);
nor U3254 (N_3254,N_1795,N_981);
nor U3255 (N_3255,N_831,N_1890);
and U3256 (N_3256,N_1532,N_1654);
nor U3257 (N_3257,N_1902,N_745);
and U3258 (N_3258,N_333,N_1397);
or U3259 (N_3259,N_1738,N_1727);
nor U3260 (N_3260,N_184,N_1777);
nand U3261 (N_3261,N_1089,N_679);
nand U3262 (N_3262,N_1458,N_852);
nand U3263 (N_3263,N_1612,N_131);
or U3264 (N_3264,N_1100,N_816);
nor U3265 (N_3265,N_182,N_1488);
nand U3266 (N_3266,N_1899,N_952);
and U3267 (N_3267,N_1250,N_562);
xor U3268 (N_3268,N_311,N_794);
nand U3269 (N_3269,N_1368,N_1431);
or U3270 (N_3270,N_214,N_286);
and U3271 (N_3271,N_1669,N_1191);
nor U3272 (N_3272,N_849,N_1369);
xor U3273 (N_3273,N_998,N_1292);
nor U3274 (N_3274,N_894,N_1326);
and U3275 (N_3275,N_770,N_1104);
or U3276 (N_3276,N_1405,N_1779);
nor U3277 (N_3277,N_1837,N_164);
and U3278 (N_3278,N_1330,N_598);
nor U3279 (N_3279,N_282,N_21);
or U3280 (N_3280,N_210,N_1570);
nand U3281 (N_3281,N_868,N_554);
nor U3282 (N_3282,N_868,N_1951);
and U3283 (N_3283,N_1788,N_277);
nand U3284 (N_3284,N_976,N_1494);
and U3285 (N_3285,N_564,N_1960);
and U3286 (N_3286,N_1743,N_1534);
and U3287 (N_3287,N_1245,N_1869);
or U3288 (N_3288,N_217,N_1168);
nor U3289 (N_3289,N_1758,N_1057);
nand U3290 (N_3290,N_1632,N_668);
nor U3291 (N_3291,N_865,N_1384);
nor U3292 (N_3292,N_1074,N_1618);
and U3293 (N_3293,N_1701,N_1911);
nor U3294 (N_3294,N_1909,N_323);
and U3295 (N_3295,N_678,N_1115);
and U3296 (N_3296,N_35,N_817);
and U3297 (N_3297,N_100,N_516);
or U3298 (N_3298,N_662,N_672);
and U3299 (N_3299,N_1830,N_665);
and U3300 (N_3300,N_191,N_1361);
nor U3301 (N_3301,N_1291,N_641);
nand U3302 (N_3302,N_194,N_652);
or U3303 (N_3303,N_229,N_1157);
nand U3304 (N_3304,N_191,N_1843);
and U3305 (N_3305,N_551,N_1298);
nor U3306 (N_3306,N_1730,N_491);
and U3307 (N_3307,N_474,N_1992);
nor U3308 (N_3308,N_1274,N_1116);
or U3309 (N_3309,N_1645,N_1040);
nor U3310 (N_3310,N_1248,N_767);
xor U3311 (N_3311,N_1805,N_571);
and U3312 (N_3312,N_231,N_1328);
or U3313 (N_3313,N_1355,N_1532);
or U3314 (N_3314,N_64,N_884);
nor U3315 (N_3315,N_45,N_466);
and U3316 (N_3316,N_1134,N_1072);
nor U3317 (N_3317,N_194,N_909);
nand U3318 (N_3318,N_1523,N_1561);
and U3319 (N_3319,N_1969,N_697);
or U3320 (N_3320,N_770,N_133);
or U3321 (N_3321,N_624,N_1971);
nor U3322 (N_3322,N_148,N_995);
and U3323 (N_3323,N_1373,N_105);
and U3324 (N_3324,N_1013,N_1872);
and U3325 (N_3325,N_1539,N_954);
nand U3326 (N_3326,N_465,N_196);
or U3327 (N_3327,N_1069,N_1801);
nand U3328 (N_3328,N_1614,N_1946);
or U3329 (N_3329,N_1370,N_1195);
nand U3330 (N_3330,N_456,N_712);
and U3331 (N_3331,N_976,N_59);
or U3332 (N_3332,N_1760,N_1567);
or U3333 (N_3333,N_235,N_303);
and U3334 (N_3334,N_383,N_1321);
and U3335 (N_3335,N_668,N_72);
nor U3336 (N_3336,N_1691,N_678);
and U3337 (N_3337,N_293,N_1106);
nor U3338 (N_3338,N_850,N_1863);
and U3339 (N_3339,N_1542,N_608);
nor U3340 (N_3340,N_971,N_897);
or U3341 (N_3341,N_920,N_1330);
nand U3342 (N_3342,N_1620,N_1304);
nor U3343 (N_3343,N_1084,N_396);
or U3344 (N_3344,N_29,N_632);
or U3345 (N_3345,N_1075,N_479);
and U3346 (N_3346,N_1647,N_990);
nand U3347 (N_3347,N_1815,N_454);
nand U3348 (N_3348,N_778,N_644);
nand U3349 (N_3349,N_863,N_1794);
or U3350 (N_3350,N_1633,N_1829);
or U3351 (N_3351,N_503,N_335);
nand U3352 (N_3352,N_984,N_92);
or U3353 (N_3353,N_360,N_1721);
nand U3354 (N_3354,N_767,N_505);
and U3355 (N_3355,N_1875,N_1592);
nand U3356 (N_3356,N_648,N_565);
nor U3357 (N_3357,N_1443,N_824);
nand U3358 (N_3358,N_871,N_1456);
and U3359 (N_3359,N_1082,N_1485);
or U3360 (N_3360,N_1147,N_1482);
nor U3361 (N_3361,N_859,N_1532);
and U3362 (N_3362,N_952,N_723);
xor U3363 (N_3363,N_1611,N_1153);
or U3364 (N_3364,N_425,N_1068);
and U3365 (N_3365,N_130,N_1725);
nand U3366 (N_3366,N_1220,N_1551);
and U3367 (N_3367,N_1668,N_1126);
and U3368 (N_3368,N_1408,N_357);
nand U3369 (N_3369,N_306,N_1968);
and U3370 (N_3370,N_251,N_211);
nor U3371 (N_3371,N_1640,N_295);
or U3372 (N_3372,N_1665,N_1933);
or U3373 (N_3373,N_662,N_1333);
and U3374 (N_3374,N_1606,N_652);
or U3375 (N_3375,N_1802,N_444);
and U3376 (N_3376,N_1735,N_668);
or U3377 (N_3377,N_175,N_1900);
nand U3378 (N_3378,N_1501,N_1600);
nor U3379 (N_3379,N_1132,N_842);
or U3380 (N_3380,N_1954,N_837);
and U3381 (N_3381,N_1359,N_613);
and U3382 (N_3382,N_14,N_806);
and U3383 (N_3383,N_1200,N_894);
and U3384 (N_3384,N_1274,N_1785);
or U3385 (N_3385,N_511,N_688);
or U3386 (N_3386,N_986,N_788);
nand U3387 (N_3387,N_280,N_1345);
nand U3388 (N_3388,N_153,N_247);
nor U3389 (N_3389,N_1548,N_1024);
nand U3390 (N_3390,N_1808,N_1652);
nand U3391 (N_3391,N_1537,N_835);
nor U3392 (N_3392,N_542,N_1597);
nor U3393 (N_3393,N_0,N_889);
or U3394 (N_3394,N_1133,N_1593);
or U3395 (N_3395,N_75,N_957);
and U3396 (N_3396,N_549,N_642);
nor U3397 (N_3397,N_608,N_1253);
or U3398 (N_3398,N_889,N_1743);
nand U3399 (N_3399,N_968,N_1999);
or U3400 (N_3400,N_309,N_1319);
nand U3401 (N_3401,N_60,N_718);
or U3402 (N_3402,N_1976,N_1037);
nand U3403 (N_3403,N_1053,N_942);
or U3404 (N_3404,N_1366,N_963);
and U3405 (N_3405,N_1613,N_419);
nand U3406 (N_3406,N_768,N_1566);
or U3407 (N_3407,N_1588,N_561);
or U3408 (N_3408,N_1736,N_723);
and U3409 (N_3409,N_1837,N_1739);
and U3410 (N_3410,N_1437,N_1136);
nand U3411 (N_3411,N_1046,N_1608);
nand U3412 (N_3412,N_499,N_1364);
nor U3413 (N_3413,N_1446,N_1030);
nand U3414 (N_3414,N_1951,N_570);
or U3415 (N_3415,N_117,N_85);
and U3416 (N_3416,N_744,N_148);
or U3417 (N_3417,N_1342,N_1495);
and U3418 (N_3418,N_1065,N_1508);
nand U3419 (N_3419,N_328,N_245);
nand U3420 (N_3420,N_1902,N_1401);
nor U3421 (N_3421,N_66,N_559);
nor U3422 (N_3422,N_1785,N_219);
or U3423 (N_3423,N_1695,N_1566);
or U3424 (N_3424,N_1327,N_344);
and U3425 (N_3425,N_464,N_1708);
or U3426 (N_3426,N_1211,N_1984);
or U3427 (N_3427,N_853,N_445);
nand U3428 (N_3428,N_1777,N_563);
nor U3429 (N_3429,N_396,N_471);
nor U3430 (N_3430,N_84,N_1794);
and U3431 (N_3431,N_427,N_1529);
nor U3432 (N_3432,N_1339,N_1252);
nand U3433 (N_3433,N_376,N_512);
nor U3434 (N_3434,N_1,N_860);
nor U3435 (N_3435,N_1924,N_527);
nand U3436 (N_3436,N_1139,N_94);
nand U3437 (N_3437,N_111,N_747);
nand U3438 (N_3438,N_301,N_1837);
and U3439 (N_3439,N_1934,N_1795);
or U3440 (N_3440,N_950,N_18);
or U3441 (N_3441,N_113,N_576);
and U3442 (N_3442,N_883,N_1575);
and U3443 (N_3443,N_70,N_1746);
nand U3444 (N_3444,N_614,N_1241);
or U3445 (N_3445,N_1326,N_1395);
and U3446 (N_3446,N_431,N_1186);
nand U3447 (N_3447,N_825,N_635);
nand U3448 (N_3448,N_1362,N_635);
nand U3449 (N_3449,N_210,N_397);
or U3450 (N_3450,N_1034,N_122);
or U3451 (N_3451,N_654,N_1541);
and U3452 (N_3452,N_1414,N_1743);
nand U3453 (N_3453,N_441,N_1050);
and U3454 (N_3454,N_1704,N_1376);
and U3455 (N_3455,N_1408,N_721);
nor U3456 (N_3456,N_1040,N_824);
nor U3457 (N_3457,N_29,N_1435);
or U3458 (N_3458,N_1631,N_1847);
and U3459 (N_3459,N_966,N_173);
or U3460 (N_3460,N_1114,N_260);
nand U3461 (N_3461,N_1783,N_92);
or U3462 (N_3462,N_752,N_528);
nand U3463 (N_3463,N_1208,N_1405);
and U3464 (N_3464,N_1147,N_431);
nor U3465 (N_3465,N_625,N_764);
nor U3466 (N_3466,N_77,N_16);
nor U3467 (N_3467,N_1653,N_1793);
xnor U3468 (N_3468,N_107,N_596);
or U3469 (N_3469,N_854,N_136);
nor U3470 (N_3470,N_518,N_1482);
nor U3471 (N_3471,N_388,N_1003);
nor U3472 (N_3472,N_715,N_1986);
nand U3473 (N_3473,N_728,N_1735);
nand U3474 (N_3474,N_1189,N_822);
and U3475 (N_3475,N_517,N_1591);
and U3476 (N_3476,N_584,N_1646);
or U3477 (N_3477,N_978,N_454);
or U3478 (N_3478,N_610,N_1710);
nand U3479 (N_3479,N_181,N_775);
nor U3480 (N_3480,N_1738,N_404);
or U3481 (N_3481,N_442,N_316);
and U3482 (N_3482,N_1967,N_710);
nor U3483 (N_3483,N_1301,N_1549);
nand U3484 (N_3484,N_907,N_1757);
and U3485 (N_3485,N_1043,N_1657);
and U3486 (N_3486,N_82,N_357);
and U3487 (N_3487,N_78,N_1767);
nand U3488 (N_3488,N_815,N_1869);
nand U3489 (N_3489,N_251,N_873);
nor U3490 (N_3490,N_1981,N_1761);
or U3491 (N_3491,N_1183,N_799);
or U3492 (N_3492,N_1863,N_344);
or U3493 (N_3493,N_261,N_1676);
nand U3494 (N_3494,N_681,N_419);
nand U3495 (N_3495,N_481,N_391);
or U3496 (N_3496,N_1954,N_1770);
or U3497 (N_3497,N_1073,N_1172);
nor U3498 (N_3498,N_1174,N_531);
nand U3499 (N_3499,N_800,N_550);
nor U3500 (N_3500,N_1641,N_1652);
or U3501 (N_3501,N_1692,N_1681);
nor U3502 (N_3502,N_1265,N_32);
xnor U3503 (N_3503,N_920,N_628);
nand U3504 (N_3504,N_533,N_1605);
and U3505 (N_3505,N_1463,N_42);
nand U3506 (N_3506,N_941,N_1448);
or U3507 (N_3507,N_986,N_844);
and U3508 (N_3508,N_1367,N_743);
nor U3509 (N_3509,N_33,N_928);
nor U3510 (N_3510,N_11,N_1750);
nand U3511 (N_3511,N_1948,N_1245);
and U3512 (N_3512,N_1698,N_1996);
nor U3513 (N_3513,N_354,N_1868);
nor U3514 (N_3514,N_207,N_782);
and U3515 (N_3515,N_805,N_581);
or U3516 (N_3516,N_1035,N_1499);
and U3517 (N_3517,N_974,N_1177);
nor U3518 (N_3518,N_1561,N_1291);
nor U3519 (N_3519,N_405,N_1406);
nor U3520 (N_3520,N_1469,N_1948);
nand U3521 (N_3521,N_1919,N_1868);
and U3522 (N_3522,N_1690,N_375);
or U3523 (N_3523,N_976,N_1043);
or U3524 (N_3524,N_1072,N_56);
nor U3525 (N_3525,N_642,N_1058);
and U3526 (N_3526,N_1810,N_1317);
nor U3527 (N_3527,N_1843,N_1403);
and U3528 (N_3528,N_1206,N_1267);
and U3529 (N_3529,N_744,N_160);
or U3530 (N_3530,N_870,N_676);
nor U3531 (N_3531,N_1886,N_1240);
or U3532 (N_3532,N_1501,N_907);
or U3533 (N_3533,N_1143,N_1181);
nand U3534 (N_3534,N_863,N_1121);
and U3535 (N_3535,N_563,N_910);
nor U3536 (N_3536,N_361,N_1064);
xor U3537 (N_3537,N_481,N_345);
or U3538 (N_3538,N_250,N_1164);
nor U3539 (N_3539,N_180,N_51);
or U3540 (N_3540,N_933,N_1005);
nor U3541 (N_3541,N_1103,N_70);
or U3542 (N_3542,N_1388,N_542);
nand U3543 (N_3543,N_1862,N_59);
nor U3544 (N_3544,N_708,N_44);
nor U3545 (N_3545,N_1091,N_541);
and U3546 (N_3546,N_1807,N_1693);
and U3547 (N_3547,N_1302,N_1947);
nor U3548 (N_3548,N_1594,N_175);
nor U3549 (N_3549,N_80,N_1704);
nand U3550 (N_3550,N_1713,N_1599);
nor U3551 (N_3551,N_134,N_867);
or U3552 (N_3552,N_871,N_352);
and U3553 (N_3553,N_1818,N_1114);
nand U3554 (N_3554,N_416,N_476);
nor U3555 (N_3555,N_39,N_554);
or U3556 (N_3556,N_1666,N_488);
nor U3557 (N_3557,N_1702,N_597);
or U3558 (N_3558,N_1060,N_1917);
or U3559 (N_3559,N_573,N_839);
nor U3560 (N_3560,N_1530,N_77);
nor U3561 (N_3561,N_1811,N_195);
xnor U3562 (N_3562,N_1689,N_811);
nand U3563 (N_3563,N_1939,N_1491);
or U3564 (N_3564,N_1187,N_416);
or U3565 (N_3565,N_365,N_539);
nor U3566 (N_3566,N_1265,N_543);
and U3567 (N_3567,N_1983,N_1805);
and U3568 (N_3568,N_1098,N_1569);
nand U3569 (N_3569,N_1875,N_1724);
nand U3570 (N_3570,N_1147,N_413);
nand U3571 (N_3571,N_1127,N_1528);
nor U3572 (N_3572,N_887,N_223);
nand U3573 (N_3573,N_250,N_0);
nand U3574 (N_3574,N_1887,N_1858);
nand U3575 (N_3575,N_1486,N_786);
nand U3576 (N_3576,N_1806,N_112);
nand U3577 (N_3577,N_164,N_1107);
nor U3578 (N_3578,N_1680,N_1951);
nand U3579 (N_3579,N_420,N_215);
and U3580 (N_3580,N_931,N_985);
nand U3581 (N_3581,N_1316,N_1250);
or U3582 (N_3582,N_420,N_893);
nor U3583 (N_3583,N_1154,N_1141);
and U3584 (N_3584,N_197,N_1163);
or U3585 (N_3585,N_1999,N_1233);
nor U3586 (N_3586,N_1524,N_1213);
or U3587 (N_3587,N_573,N_449);
nand U3588 (N_3588,N_1668,N_1860);
nand U3589 (N_3589,N_1299,N_1722);
nor U3590 (N_3590,N_1854,N_1335);
and U3591 (N_3591,N_579,N_1958);
and U3592 (N_3592,N_1004,N_156);
and U3593 (N_3593,N_492,N_1852);
nor U3594 (N_3594,N_543,N_1088);
nor U3595 (N_3595,N_1035,N_536);
or U3596 (N_3596,N_411,N_1937);
or U3597 (N_3597,N_643,N_429);
and U3598 (N_3598,N_1927,N_974);
nand U3599 (N_3599,N_1292,N_1423);
nor U3600 (N_3600,N_597,N_1577);
nor U3601 (N_3601,N_371,N_1947);
and U3602 (N_3602,N_1696,N_1098);
and U3603 (N_3603,N_170,N_1192);
nor U3604 (N_3604,N_964,N_1058);
or U3605 (N_3605,N_458,N_1451);
or U3606 (N_3606,N_1524,N_1640);
and U3607 (N_3607,N_1302,N_1566);
nor U3608 (N_3608,N_983,N_1002);
or U3609 (N_3609,N_1263,N_1287);
nor U3610 (N_3610,N_1986,N_1838);
nand U3611 (N_3611,N_592,N_396);
or U3612 (N_3612,N_1471,N_537);
nand U3613 (N_3613,N_1240,N_1106);
nand U3614 (N_3614,N_1784,N_809);
nor U3615 (N_3615,N_978,N_1647);
or U3616 (N_3616,N_1935,N_874);
nor U3617 (N_3617,N_1362,N_1520);
and U3618 (N_3618,N_134,N_948);
or U3619 (N_3619,N_426,N_1903);
and U3620 (N_3620,N_436,N_454);
or U3621 (N_3621,N_806,N_1665);
xnor U3622 (N_3622,N_832,N_256);
and U3623 (N_3623,N_1468,N_29);
nor U3624 (N_3624,N_1299,N_1900);
and U3625 (N_3625,N_103,N_1135);
nand U3626 (N_3626,N_1304,N_1948);
nand U3627 (N_3627,N_1215,N_1923);
and U3628 (N_3628,N_1720,N_264);
or U3629 (N_3629,N_1546,N_1186);
or U3630 (N_3630,N_1801,N_1874);
nor U3631 (N_3631,N_597,N_1589);
nand U3632 (N_3632,N_1049,N_1305);
nor U3633 (N_3633,N_616,N_1068);
and U3634 (N_3634,N_1582,N_472);
nand U3635 (N_3635,N_356,N_1314);
nor U3636 (N_3636,N_223,N_843);
or U3637 (N_3637,N_274,N_1706);
and U3638 (N_3638,N_1343,N_1788);
nand U3639 (N_3639,N_1859,N_814);
and U3640 (N_3640,N_932,N_1672);
or U3641 (N_3641,N_1157,N_718);
nand U3642 (N_3642,N_727,N_459);
and U3643 (N_3643,N_1449,N_532);
and U3644 (N_3644,N_1282,N_752);
or U3645 (N_3645,N_194,N_5);
nand U3646 (N_3646,N_575,N_268);
nand U3647 (N_3647,N_92,N_1388);
nand U3648 (N_3648,N_1315,N_194);
or U3649 (N_3649,N_24,N_1385);
nand U3650 (N_3650,N_1944,N_853);
or U3651 (N_3651,N_1812,N_1437);
or U3652 (N_3652,N_1548,N_1663);
nor U3653 (N_3653,N_5,N_704);
or U3654 (N_3654,N_1044,N_625);
and U3655 (N_3655,N_1836,N_773);
nand U3656 (N_3656,N_1947,N_1229);
nand U3657 (N_3657,N_1751,N_1584);
nor U3658 (N_3658,N_484,N_1511);
and U3659 (N_3659,N_1476,N_1232);
and U3660 (N_3660,N_1608,N_355);
or U3661 (N_3661,N_740,N_482);
and U3662 (N_3662,N_435,N_1733);
nand U3663 (N_3663,N_944,N_1580);
or U3664 (N_3664,N_224,N_1615);
and U3665 (N_3665,N_725,N_502);
and U3666 (N_3666,N_520,N_1457);
and U3667 (N_3667,N_1985,N_1600);
or U3668 (N_3668,N_1755,N_1037);
nand U3669 (N_3669,N_1791,N_1757);
nand U3670 (N_3670,N_69,N_391);
or U3671 (N_3671,N_1623,N_57);
and U3672 (N_3672,N_386,N_1043);
nand U3673 (N_3673,N_719,N_1013);
or U3674 (N_3674,N_1709,N_1661);
nor U3675 (N_3675,N_1099,N_1925);
or U3676 (N_3676,N_618,N_466);
nor U3677 (N_3677,N_1765,N_924);
nor U3678 (N_3678,N_48,N_6);
and U3679 (N_3679,N_136,N_423);
nand U3680 (N_3680,N_1851,N_292);
or U3681 (N_3681,N_1003,N_1641);
and U3682 (N_3682,N_995,N_1770);
and U3683 (N_3683,N_42,N_1190);
nand U3684 (N_3684,N_1992,N_221);
or U3685 (N_3685,N_1578,N_213);
or U3686 (N_3686,N_408,N_1625);
or U3687 (N_3687,N_500,N_142);
and U3688 (N_3688,N_1850,N_1794);
nand U3689 (N_3689,N_562,N_1093);
nor U3690 (N_3690,N_930,N_1231);
nand U3691 (N_3691,N_1147,N_428);
nor U3692 (N_3692,N_569,N_1723);
nor U3693 (N_3693,N_308,N_1829);
nor U3694 (N_3694,N_1886,N_631);
and U3695 (N_3695,N_1368,N_270);
nor U3696 (N_3696,N_503,N_1546);
nand U3697 (N_3697,N_1618,N_1723);
or U3698 (N_3698,N_524,N_397);
and U3699 (N_3699,N_165,N_1845);
nor U3700 (N_3700,N_961,N_1398);
nor U3701 (N_3701,N_845,N_960);
nand U3702 (N_3702,N_194,N_13);
or U3703 (N_3703,N_134,N_549);
nand U3704 (N_3704,N_450,N_45);
or U3705 (N_3705,N_1906,N_999);
and U3706 (N_3706,N_593,N_952);
nand U3707 (N_3707,N_513,N_1876);
or U3708 (N_3708,N_721,N_981);
xor U3709 (N_3709,N_1658,N_727);
nand U3710 (N_3710,N_215,N_1490);
nand U3711 (N_3711,N_1527,N_561);
nor U3712 (N_3712,N_1643,N_883);
or U3713 (N_3713,N_1568,N_1723);
nand U3714 (N_3714,N_1217,N_1792);
nor U3715 (N_3715,N_1260,N_325);
nand U3716 (N_3716,N_1610,N_1971);
and U3717 (N_3717,N_444,N_1844);
nor U3718 (N_3718,N_306,N_1335);
or U3719 (N_3719,N_237,N_425);
and U3720 (N_3720,N_901,N_1725);
nand U3721 (N_3721,N_1141,N_1819);
or U3722 (N_3722,N_219,N_998);
nand U3723 (N_3723,N_582,N_600);
or U3724 (N_3724,N_1240,N_1762);
or U3725 (N_3725,N_894,N_256);
or U3726 (N_3726,N_931,N_1979);
and U3727 (N_3727,N_813,N_680);
xnor U3728 (N_3728,N_943,N_36);
xnor U3729 (N_3729,N_1980,N_1877);
and U3730 (N_3730,N_475,N_1356);
and U3731 (N_3731,N_98,N_1594);
and U3732 (N_3732,N_270,N_35);
and U3733 (N_3733,N_1746,N_400);
and U3734 (N_3734,N_1770,N_1044);
nand U3735 (N_3735,N_1657,N_1262);
or U3736 (N_3736,N_207,N_362);
nand U3737 (N_3737,N_619,N_1521);
and U3738 (N_3738,N_176,N_31);
nand U3739 (N_3739,N_1908,N_1450);
nand U3740 (N_3740,N_669,N_632);
and U3741 (N_3741,N_884,N_239);
nand U3742 (N_3742,N_898,N_695);
nor U3743 (N_3743,N_1479,N_1434);
or U3744 (N_3744,N_608,N_378);
and U3745 (N_3745,N_786,N_564);
nand U3746 (N_3746,N_393,N_1653);
nand U3747 (N_3747,N_338,N_823);
nor U3748 (N_3748,N_1126,N_1085);
and U3749 (N_3749,N_263,N_1482);
and U3750 (N_3750,N_509,N_1717);
nand U3751 (N_3751,N_1806,N_591);
or U3752 (N_3752,N_922,N_1562);
or U3753 (N_3753,N_111,N_1874);
nor U3754 (N_3754,N_400,N_1169);
and U3755 (N_3755,N_1889,N_1886);
and U3756 (N_3756,N_291,N_1327);
or U3757 (N_3757,N_103,N_614);
nor U3758 (N_3758,N_1974,N_1884);
nor U3759 (N_3759,N_624,N_623);
and U3760 (N_3760,N_1740,N_1073);
nor U3761 (N_3761,N_1394,N_13);
nand U3762 (N_3762,N_660,N_708);
and U3763 (N_3763,N_1207,N_745);
nand U3764 (N_3764,N_1436,N_87);
or U3765 (N_3765,N_894,N_1113);
or U3766 (N_3766,N_556,N_1737);
nand U3767 (N_3767,N_602,N_1152);
and U3768 (N_3768,N_303,N_1387);
and U3769 (N_3769,N_342,N_321);
nor U3770 (N_3770,N_660,N_524);
and U3771 (N_3771,N_454,N_274);
nand U3772 (N_3772,N_600,N_1123);
nor U3773 (N_3773,N_744,N_162);
nor U3774 (N_3774,N_381,N_5);
nand U3775 (N_3775,N_1118,N_209);
and U3776 (N_3776,N_1107,N_88);
nand U3777 (N_3777,N_804,N_113);
xnor U3778 (N_3778,N_1558,N_216);
nand U3779 (N_3779,N_1051,N_1347);
nor U3780 (N_3780,N_1049,N_1187);
and U3781 (N_3781,N_1265,N_706);
or U3782 (N_3782,N_613,N_1092);
or U3783 (N_3783,N_38,N_253);
xnor U3784 (N_3784,N_1797,N_1166);
and U3785 (N_3785,N_1030,N_1613);
or U3786 (N_3786,N_1039,N_1131);
nand U3787 (N_3787,N_605,N_1052);
or U3788 (N_3788,N_4,N_444);
or U3789 (N_3789,N_74,N_77);
nand U3790 (N_3790,N_651,N_1311);
nand U3791 (N_3791,N_394,N_1897);
nand U3792 (N_3792,N_1604,N_1442);
nand U3793 (N_3793,N_562,N_1412);
nand U3794 (N_3794,N_1348,N_139);
nor U3795 (N_3795,N_1985,N_1994);
or U3796 (N_3796,N_349,N_893);
nor U3797 (N_3797,N_698,N_1090);
nor U3798 (N_3798,N_1170,N_1219);
and U3799 (N_3799,N_218,N_624);
nor U3800 (N_3800,N_901,N_1216);
nor U3801 (N_3801,N_1512,N_1223);
or U3802 (N_3802,N_649,N_200);
nor U3803 (N_3803,N_159,N_984);
and U3804 (N_3804,N_1559,N_619);
or U3805 (N_3805,N_244,N_1566);
nor U3806 (N_3806,N_1344,N_1843);
or U3807 (N_3807,N_418,N_432);
nand U3808 (N_3808,N_473,N_520);
or U3809 (N_3809,N_897,N_219);
and U3810 (N_3810,N_1089,N_397);
nor U3811 (N_3811,N_709,N_1525);
or U3812 (N_3812,N_1853,N_4);
nand U3813 (N_3813,N_1053,N_1351);
or U3814 (N_3814,N_1093,N_427);
nand U3815 (N_3815,N_1985,N_159);
nor U3816 (N_3816,N_1725,N_763);
or U3817 (N_3817,N_389,N_970);
nand U3818 (N_3818,N_1551,N_701);
or U3819 (N_3819,N_1394,N_1350);
and U3820 (N_3820,N_767,N_1294);
and U3821 (N_3821,N_93,N_905);
nand U3822 (N_3822,N_1162,N_554);
nand U3823 (N_3823,N_853,N_1010);
nand U3824 (N_3824,N_1744,N_591);
nor U3825 (N_3825,N_1548,N_1600);
nor U3826 (N_3826,N_1845,N_1208);
or U3827 (N_3827,N_1449,N_1458);
or U3828 (N_3828,N_198,N_1947);
nand U3829 (N_3829,N_673,N_337);
or U3830 (N_3830,N_187,N_1667);
or U3831 (N_3831,N_1682,N_47);
nor U3832 (N_3832,N_42,N_1908);
nor U3833 (N_3833,N_88,N_1374);
nand U3834 (N_3834,N_692,N_1546);
and U3835 (N_3835,N_923,N_555);
nor U3836 (N_3836,N_259,N_1095);
or U3837 (N_3837,N_800,N_614);
nand U3838 (N_3838,N_20,N_1595);
and U3839 (N_3839,N_1091,N_14);
xnor U3840 (N_3840,N_694,N_1151);
nor U3841 (N_3841,N_700,N_223);
and U3842 (N_3842,N_931,N_1136);
nor U3843 (N_3843,N_1748,N_387);
nor U3844 (N_3844,N_1429,N_815);
nor U3845 (N_3845,N_1066,N_1613);
nor U3846 (N_3846,N_1985,N_224);
nor U3847 (N_3847,N_287,N_1271);
or U3848 (N_3848,N_1874,N_840);
nand U3849 (N_3849,N_625,N_743);
or U3850 (N_3850,N_316,N_1807);
and U3851 (N_3851,N_631,N_1609);
nand U3852 (N_3852,N_1885,N_650);
and U3853 (N_3853,N_347,N_1027);
and U3854 (N_3854,N_1830,N_1187);
and U3855 (N_3855,N_1347,N_1110);
nand U3856 (N_3856,N_48,N_969);
nor U3857 (N_3857,N_818,N_1139);
nand U3858 (N_3858,N_1578,N_1166);
or U3859 (N_3859,N_108,N_1081);
nor U3860 (N_3860,N_1457,N_562);
or U3861 (N_3861,N_1823,N_150);
and U3862 (N_3862,N_424,N_653);
nor U3863 (N_3863,N_1617,N_761);
nor U3864 (N_3864,N_1991,N_1088);
and U3865 (N_3865,N_826,N_1261);
and U3866 (N_3866,N_811,N_16);
nand U3867 (N_3867,N_576,N_199);
or U3868 (N_3868,N_1258,N_1500);
nor U3869 (N_3869,N_1059,N_175);
and U3870 (N_3870,N_1036,N_68);
or U3871 (N_3871,N_485,N_1012);
xor U3872 (N_3872,N_1473,N_1521);
and U3873 (N_3873,N_1503,N_348);
or U3874 (N_3874,N_1140,N_424);
nor U3875 (N_3875,N_20,N_790);
nand U3876 (N_3876,N_1209,N_799);
or U3877 (N_3877,N_45,N_729);
or U3878 (N_3878,N_1570,N_676);
or U3879 (N_3879,N_1249,N_782);
or U3880 (N_3880,N_1006,N_1469);
nand U3881 (N_3881,N_1563,N_813);
and U3882 (N_3882,N_707,N_291);
nand U3883 (N_3883,N_171,N_124);
and U3884 (N_3884,N_1122,N_1002);
or U3885 (N_3885,N_236,N_1455);
nor U3886 (N_3886,N_1761,N_1993);
or U3887 (N_3887,N_986,N_1754);
nand U3888 (N_3888,N_1127,N_779);
nor U3889 (N_3889,N_793,N_1644);
and U3890 (N_3890,N_1639,N_309);
nand U3891 (N_3891,N_352,N_916);
and U3892 (N_3892,N_1138,N_1227);
or U3893 (N_3893,N_1140,N_769);
and U3894 (N_3894,N_1732,N_1788);
and U3895 (N_3895,N_866,N_1559);
and U3896 (N_3896,N_933,N_1672);
xor U3897 (N_3897,N_1775,N_1415);
and U3898 (N_3898,N_377,N_8);
nand U3899 (N_3899,N_899,N_974);
and U3900 (N_3900,N_1112,N_406);
nor U3901 (N_3901,N_1567,N_1057);
nor U3902 (N_3902,N_1227,N_1063);
or U3903 (N_3903,N_175,N_502);
or U3904 (N_3904,N_1088,N_807);
and U3905 (N_3905,N_1943,N_1390);
nand U3906 (N_3906,N_1161,N_1677);
nand U3907 (N_3907,N_81,N_1135);
nand U3908 (N_3908,N_1140,N_1195);
and U3909 (N_3909,N_1148,N_1903);
nand U3910 (N_3910,N_1058,N_1245);
or U3911 (N_3911,N_1022,N_583);
nand U3912 (N_3912,N_1777,N_1206);
nand U3913 (N_3913,N_317,N_776);
and U3914 (N_3914,N_1442,N_21);
nand U3915 (N_3915,N_1657,N_1498);
and U3916 (N_3916,N_1529,N_171);
or U3917 (N_3917,N_415,N_1528);
or U3918 (N_3918,N_1369,N_335);
and U3919 (N_3919,N_1225,N_515);
or U3920 (N_3920,N_1394,N_1814);
and U3921 (N_3921,N_1903,N_304);
or U3922 (N_3922,N_312,N_28);
nor U3923 (N_3923,N_1070,N_203);
and U3924 (N_3924,N_114,N_468);
or U3925 (N_3925,N_491,N_1715);
and U3926 (N_3926,N_647,N_1792);
nand U3927 (N_3927,N_976,N_1039);
and U3928 (N_3928,N_874,N_1442);
nand U3929 (N_3929,N_1655,N_1119);
nand U3930 (N_3930,N_1948,N_626);
or U3931 (N_3931,N_1369,N_46);
nor U3932 (N_3932,N_580,N_350);
and U3933 (N_3933,N_1474,N_266);
or U3934 (N_3934,N_568,N_1143);
nand U3935 (N_3935,N_1425,N_1971);
nand U3936 (N_3936,N_492,N_1362);
nand U3937 (N_3937,N_728,N_432);
or U3938 (N_3938,N_1791,N_1269);
nand U3939 (N_3939,N_1003,N_38);
nand U3940 (N_3940,N_974,N_505);
nand U3941 (N_3941,N_831,N_1082);
and U3942 (N_3942,N_387,N_230);
or U3943 (N_3943,N_934,N_99);
nor U3944 (N_3944,N_1133,N_65);
nor U3945 (N_3945,N_664,N_69);
nand U3946 (N_3946,N_154,N_1945);
nor U3947 (N_3947,N_1462,N_893);
or U3948 (N_3948,N_674,N_722);
nor U3949 (N_3949,N_1722,N_1126);
and U3950 (N_3950,N_549,N_1458);
nor U3951 (N_3951,N_212,N_1206);
nand U3952 (N_3952,N_468,N_830);
nand U3953 (N_3953,N_989,N_1269);
and U3954 (N_3954,N_877,N_478);
nor U3955 (N_3955,N_141,N_1554);
and U3956 (N_3956,N_1257,N_1194);
nand U3957 (N_3957,N_1676,N_347);
or U3958 (N_3958,N_1026,N_1520);
nand U3959 (N_3959,N_287,N_577);
nor U3960 (N_3960,N_563,N_515);
nand U3961 (N_3961,N_1236,N_1565);
nor U3962 (N_3962,N_158,N_1521);
nor U3963 (N_3963,N_1833,N_1864);
nor U3964 (N_3964,N_1783,N_1725);
nand U3965 (N_3965,N_1553,N_94);
nand U3966 (N_3966,N_499,N_114);
or U3967 (N_3967,N_40,N_1203);
and U3968 (N_3968,N_608,N_321);
nand U3969 (N_3969,N_4,N_838);
and U3970 (N_3970,N_1097,N_1450);
or U3971 (N_3971,N_823,N_1300);
nor U3972 (N_3972,N_1928,N_748);
nor U3973 (N_3973,N_1940,N_793);
or U3974 (N_3974,N_818,N_205);
nand U3975 (N_3975,N_1789,N_1043);
nor U3976 (N_3976,N_513,N_207);
and U3977 (N_3977,N_1123,N_250);
nand U3978 (N_3978,N_1700,N_1078);
nand U3979 (N_3979,N_175,N_1481);
nor U3980 (N_3980,N_1583,N_619);
or U3981 (N_3981,N_403,N_1113);
nor U3982 (N_3982,N_1329,N_826);
nor U3983 (N_3983,N_75,N_1746);
or U3984 (N_3984,N_1129,N_1458);
nor U3985 (N_3985,N_30,N_40);
nor U3986 (N_3986,N_34,N_915);
nor U3987 (N_3987,N_704,N_624);
or U3988 (N_3988,N_1883,N_224);
and U3989 (N_3989,N_1158,N_1295);
or U3990 (N_3990,N_1124,N_1452);
and U3991 (N_3991,N_1225,N_1356);
or U3992 (N_3992,N_180,N_1743);
or U3993 (N_3993,N_250,N_193);
nor U3994 (N_3994,N_495,N_1737);
and U3995 (N_3995,N_1873,N_578);
and U3996 (N_3996,N_460,N_1404);
nor U3997 (N_3997,N_425,N_388);
or U3998 (N_3998,N_1121,N_880);
nor U3999 (N_3999,N_814,N_1965);
or U4000 (N_4000,N_3108,N_2819);
nand U4001 (N_4001,N_2483,N_3262);
nor U4002 (N_4002,N_3364,N_3204);
nand U4003 (N_4003,N_2833,N_3597);
or U4004 (N_4004,N_3988,N_2508);
nand U4005 (N_4005,N_2109,N_2762);
nand U4006 (N_4006,N_3451,N_3498);
nand U4007 (N_4007,N_2395,N_3112);
or U4008 (N_4008,N_3740,N_3678);
nand U4009 (N_4009,N_2836,N_2667);
and U4010 (N_4010,N_2357,N_2979);
or U4011 (N_4011,N_3341,N_3157);
nor U4012 (N_4012,N_3716,N_2329);
and U4013 (N_4013,N_2846,N_3943);
nand U4014 (N_4014,N_2513,N_2177);
nand U4015 (N_4015,N_2607,N_3055);
nand U4016 (N_4016,N_2563,N_2690);
and U4017 (N_4017,N_3193,N_3124);
nor U4018 (N_4018,N_3966,N_3032);
or U4019 (N_4019,N_3294,N_3166);
and U4020 (N_4020,N_3984,N_2258);
and U4021 (N_4021,N_2014,N_3615);
nor U4022 (N_4022,N_3800,N_2188);
nor U4023 (N_4023,N_2999,N_2000);
or U4024 (N_4024,N_3210,N_2479);
nand U4025 (N_4025,N_2981,N_3351);
and U4026 (N_4026,N_3776,N_2326);
nor U4027 (N_4027,N_2117,N_2151);
nand U4028 (N_4028,N_2487,N_3626);
nor U4029 (N_4029,N_3468,N_3192);
or U4030 (N_4030,N_3565,N_2063);
nand U4031 (N_4031,N_3066,N_2373);
nand U4032 (N_4032,N_3080,N_3391);
and U4033 (N_4033,N_3825,N_2535);
nand U4034 (N_4034,N_2438,N_3777);
nand U4035 (N_4035,N_3896,N_3334);
and U4036 (N_4036,N_2350,N_2295);
nand U4037 (N_4037,N_2983,N_2824);
or U4038 (N_4038,N_2577,N_3070);
nand U4039 (N_4039,N_3168,N_2921);
nand U4040 (N_4040,N_3995,N_2728);
nand U4041 (N_4041,N_2221,N_2495);
and U4042 (N_4042,N_2382,N_2428);
or U4043 (N_4043,N_3295,N_2924);
nor U4044 (N_4044,N_2472,N_3891);
nand U4045 (N_4045,N_3692,N_2333);
and U4046 (N_4046,N_2925,N_3301);
or U4047 (N_4047,N_2374,N_2920);
nand U4048 (N_4048,N_2414,N_2340);
xnor U4049 (N_4049,N_3296,N_2678);
nor U4050 (N_4050,N_3371,N_2792);
and U4051 (N_4051,N_2183,N_2356);
and U4052 (N_4052,N_2649,N_3337);
nor U4053 (N_4053,N_3932,N_3178);
or U4054 (N_4054,N_3452,N_3450);
or U4055 (N_4055,N_2615,N_3456);
or U4056 (N_4056,N_3017,N_2206);
and U4057 (N_4057,N_3233,N_2281);
nand U4058 (N_4058,N_3858,N_3768);
or U4059 (N_4059,N_2166,N_3964);
nor U4060 (N_4060,N_3038,N_2353);
and U4061 (N_4061,N_3815,N_3308);
and U4062 (N_4062,N_3485,N_2372);
nor U4063 (N_4063,N_2279,N_3472);
or U4064 (N_4064,N_3093,N_2631);
and U4065 (N_4065,N_2634,N_3167);
or U4066 (N_4066,N_2768,N_3189);
xor U4067 (N_4067,N_2599,N_3852);
xnor U4068 (N_4068,N_3562,N_2540);
and U4069 (N_4069,N_2155,N_2504);
or U4070 (N_4070,N_3689,N_2711);
or U4071 (N_4071,N_3957,N_2590);
and U4072 (N_4072,N_2572,N_2855);
nand U4073 (N_4073,N_2229,N_3673);
and U4074 (N_4074,N_3828,N_2400);
and U4075 (N_4075,N_2717,N_3770);
nand U4076 (N_4076,N_3547,N_2880);
and U4077 (N_4077,N_3090,N_2881);
or U4078 (N_4078,N_3203,N_2022);
nand U4079 (N_4079,N_3211,N_3475);
nor U4080 (N_4080,N_2888,N_3739);
or U4081 (N_4081,N_3526,N_3752);
xor U4082 (N_4082,N_2074,N_2804);
or U4083 (N_4083,N_2490,N_3188);
nand U4084 (N_4084,N_3937,N_3798);
nand U4085 (N_4085,N_2791,N_3874);
or U4086 (N_4086,N_3647,N_3466);
nand U4087 (N_4087,N_2664,N_2480);
or U4088 (N_4088,N_2906,N_3100);
nor U4089 (N_4089,N_2874,N_3171);
or U4090 (N_4090,N_3343,N_3328);
or U4091 (N_4091,N_2270,N_3924);
nand U4092 (N_4092,N_3951,N_3007);
or U4093 (N_4093,N_2110,N_3478);
nor U4094 (N_4094,N_3427,N_3159);
nand U4095 (N_4095,N_2628,N_2884);
nand U4096 (N_4096,N_3175,N_3011);
and U4097 (N_4097,N_3455,N_3771);
and U4098 (N_4098,N_3836,N_3015);
nand U4099 (N_4099,N_3434,N_3042);
or U4100 (N_4100,N_3715,N_2985);
and U4101 (N_4101,N_3627,N_3195);
and U4102 (N_4102,N_3417,N_3479);
nor U4103 (N_4103,N_3026,N_3483);
or U4104 (N_4104,N_2050,N_3454);
nand U4105 (N_4105,N_3558,N_3757);
or U4106 (N_4106,N_3528,N_2026);
nand U4107 (N_4107,N_3268,N_3551);
nand U4108 (N_4108,N_2271,N_2586);
and U4109 (N_4109,N_3614,N_3938);
or U4110 (N_4110,N_2324,N_2514);
nor U4111 (N_4111,N_3674,N_2658);
and U4112 (N_4112,N_2908,N_2524);
nand U4113 (N_4113,N_3082,N_2662);
and U4114 (N_4114,N_3552,N_3734);
and U4115 (N_4115,N_2486,N_2064);
nor U4116 (N_4116,N_3877,N_3516);
nand U4117 (N_4117,N_3145,N_3069);
and U4118 (N_4118,N_3254,N_2632);
nand U4119 (N_4119,N_3135,N_3470);
nand U4120 (N_4120,N_3506,N_3062);
and U4121 (N_4121,N_3230,N_3520);
and U4122 (N_4122,N_3256,N_2697);
and U4123 (N_4123,N_3396,N_3016);
and U4124 (N_4124,N_3875,N_3902);
or U4125 (N_4125,N_3708,N_3862);
nand U4126 (N_4126,N_2457,N_2995);
nand U4127 (N_4127,N_2986,N_3854);
and U4128 (N_4128,N_2292,N_3245);
or U4129 (N_4129,N_3095,N_3677);
and U4130 (N_4130,N_3824,N_2439);
and U4131 (N_4131,N_2788,N_3711);
nor U4132 (N_4132,N_2341,N_2700);
nand U4133 (N_4133,N_3817,N_3865);
and U4134 (N_4134,N_2045,N_2316);
nor U4135 (N_4135,N_2331,N_2927);
and U4136 (N_4136,N_2500,N_3765);
nand U4137 (N_4137,N_2515,N_2956);
nand U4138 (N_4138,N_2950,N_2467);
and U4139 (N_4139,N_2043,N_2748);
and U4140 (N_4140,N_3623,N_2501);
nor U4141 (N_4141,N_2407,N_2334);
nor U4142 (N_4142,N_3033,N_2683);
nand U4143 (N_4143,N_3098,N_2716);
and U4144 (N_4144,N_2012,N_2492);
or U4145 (N_4145,N_2548,N_2893);
nand U4146 (N_4146,N_2078,N_2592);
nand U4147 (N_4147,N_2912,N_3282);
nand U4148 (N_4148,N_3944,N_3651);
nor U4149 (N_4149,N_2798,N_2023);
nor U4150 (N_4150,N_2820,N_3056);
xnor U4151 (N_4151,N_2345,N_2759);
nor U4152 (N_4152,N_2097,N_3618);
nor U4153 (N_4153,N_2058,N_2431);
and U4154 (N_4154,N_3025,N_3164);
nor U4155 (N_4155,N_3586,N_3619);
nor U4156 (N_4156,N_3002,N_2093);
nand U4157 (N_4157,N_3888,N_3217);
and U4158 (N_4158,N_3109,N_2077);
or U4159 (N_4159,N_3652,N_3119);
nor U4160 (N_4160,N_3999,N_2130);
and U4161 (N_4161,N_2967,N_3650);
nor U4162 (N_4162,N_3832,N_2168);
and U4163 (N_4163,N_3685,N_2688);
and U4164 (N_4164,N_2449,N_2231);
and U4165 (N_4165,N_3027,N_2755);
and U4166 (N_4166,N_3049,N_3773);
nor U4167 (N_4167,N_3335,N_3247);
nand U4168 (N_4168,N_2567,N_2651);
nor U4169 (N_4169,N_2485,N_3496);
and U4170 (N_4170,N_3279,N_2913);
and U4171 (N_4171,N_2140,N_3052);
or U4172 (N_4172,N_3545,N_2558);
and U4173 (N_4173,N_3379,N_3887);
and U4174 (N_4174,N_2435,N_3732);
nand U4175 (N_4175,N_3550,N_3792);
nand U4176 (N_4176,N_3931,N_2866);
nand U4177 (N_4177,N_2537,N_3050);
nand U4178 (N_4178,N_3909,N_3664);
nand U4179 (N_4179,N_3244,N_3419);
nor U4180 (N_4180,N_3345,N_2723);
nand U4181 (N_4181,N_3841,N_2876);
nor U4182 (N_4182,N_3121,N_3681);
or U4183 (N_4183,N_2699,N_3487);
and U4184 (N_4184,N_2047,N_3515);
nand U4185 (N_4185,N_2510,N_3416);
nand U4186 (N_4186,N_2554,N_2703);
nand U4187 (N_4187,N_3907,N_2303);
nand U4188 (N_4188,N_3051,N_3220);
xnor U4189 (N_4189,N_2006,N_3393);
and U4190 (N_4190,N_3111,N_2989);
and U4191 (N_4191,N_3280,N_3004);
or U4192 (N_4192,N_2718,N_2656);
and U4193 (N_4193,N_2565,N_2245);
and U4194 (N_4194,N_2830,N_2247);
or U4195 (N_4195,N_2623,N_2060);
or U4196 (N_4196,N_3845,N_3805);
nor U4197 (N_4197,N_3727,N_3612);
or U4198 (N_4198,N_2860,N_3595);
or U4199 (N_4199,N_2436,N_3730);
and U4200 (N_4200,N_2570,N_2227);
or U4201 (N_4201,N_3949,N_3641);
nor U4202 (N_4202,N_3269,N_3956);
or U4203 (N_4203,N_3846,N_3926);
or U4204 (N_4204,N_3068,N_3563);
or U4205 (N_4205,N_2828,N_2765);
nand U4206 (N_4206,N_3772,N_2808);
and U4207 (N_4207,N_3258,N_2386);
and U4208 (N_4208,N_2477,N_3539);
and U4209 (N_4209,N_3952,N_2013);
nor U4210 (N_4210,N_3310,N_2637);
nand U4211 (N_4211,N_3617,N_3355);
xnor U4212 (N_4212,N_3074,N_2252);
or U4213 (N_4213,N_2276,N_2142);
nor U4214 (N_4214,N_3543,N_2630);
nor U4215 (N_4215,N_2195,N_2827);
nor U4216 (N_4216,N_3428,N_3813);
nand U4217 (N_4217,N_3215,N_3009);
nor U4218 (N_4218,N_2761,N_2729);
nor U4219 (N_4219,N_2257,N_3645);
and U4220 (N_4220,N_2266,N_2089);
nor U4221 (N_4221,N_2559,N_2458);
nand U4222 (N_4222,N_2564,N_2444);
nor U4223 (N_4223,N_3126,N_2926);
nand U4224 (N_4224,N_3546,N_3635);
nor U4225 (N_4225,N_3710,N_2922);
and U4226 (N_4226,N_3208,N_3243);
nand U4227 (N_4227,N_3231,N_2408);
nand U4228 (N_4228,N_3467,N_2299);
nand U4229 (N_4229,N_3138,N_3120);
or U4230 (N_4230,N_3514,N_2165);
or U4231 (N_4231,N_3239,N_3696);
and U4232 (N_4232,N_2298,N_3459);
or U4233 (N_4233,N_3075,N_3866);
nand U4234 (N_4234,N_3735,N_2560);
nand U4235 (N_4235,N_2362,N_2680);
and U4236 (N_4236,N_2143,N_2197);
or U4237 (N_4237,N_3209,N_2364);
xor U4238 (N_4238,N_2453,N_2790);
nand U4239 (N_4239,N_2405,N_3968);
and U4240 (N_4240,N_2498,N_3170);
nand U4241 (N_4241,N_3046,N_3591);
or U4242 (N_4242,N_2965,N_2192);
and U4243 (N_4243,N_2978,N_3580);
or U4244 (N_4244,N_3084,N_2346);
and U4245 (N_4245,N_3150,N_3018);
nand U4246 (N_4246,N_3658,N_3024);
or U4247 (N_4247,N_3912,N_2764);
and U4248 (N_4248,N_3198,N_2147);
and U4249 (N_4249,N_3453,N_3305);
and U4250 (N_4250,N_2531,N_2429);
or U4251 (N_4251,N_3923,N_2726);
or U4252 (N_4252,N_2332,N_3144);
nor U4253 (N_4253,N_3742,N_2953);
nand U4254 (N_4254,N_2131,N_3219);
nand U4255 (N_4255,N_2970,N_2267);
nor U4256 (N_4256,N_2389,N_2360);
or U4257 (N_4257,N_2361,N_3216);
nand U4258 (N_4258,N_3141,N_2621);
nor U4259 (N_4259,N_3870,N_2911);
or U4260 (N_4260,N_3373,N_2124);
and U4261 (N_4261,N_3290,N_3382);
or U4262 (N_4262,N_2571,N_3398);
and U4263 (N_4263,N_2280,N_3557);
nand U4264 (N_4264,N_2417,N_3094);
or U4265 (N_4265,N_3083,N_3319);
or U4266 (N_4266,N_2205,N_2239);
or U4267 (N_4267,N_2943,N_3747);
nor U4268 (N_4268,N_2425,N_3590);
nand U4269 (N_4269,N_3348,N_2907);
nand U4270 (N_4270,N_3861,N_3047);
nand U4271 (N_4271,N_3272,N_3504);
or U4272 (N_4272,N_2672,N_2122);
or U4273 (N_4273,N_2609,N_3534);
nor U4274 (N_4274,N_2568,N_2832);
and U4275 (N_4275,N_3281,N_2743);
nand U4276 (N_4276,N_3346,N_3723);
nand U4277 (N_4277,N_3575,N_3997);
nand U4278 (N_4278,N_2481,N_3941);
or U4279 (N_4279,N_3699,N_3174);
nand U4280 (N_4280,N_3899,N_2910);
or U4281 (N_4281,N_2075,N_2810);
or U4282 (N_4282,N_2541,N_2371);
or U4283 (N_4283,N_3202,N_3820);
nor U4284 (N_4284,N_3162,N_3911);
and U4285 (N_4285,N_3818,N_3021);
nand U4286 (N_4286,N_3679,N_2156);
nor U4287 (N_4287,N_3400,N_3477);
nor U4288 (N_4288,N_2975,N_3315);
or U4289 (N_4289,N_2167,N_2573);
or U4290 (N_4290,N_3199,N_2948);
or U4291 (N_4291,N_2737,N_3934);
and U4292 (N_4292,N_3140,N_3733);
and U4293 (N_4293,N_3835,N_2099);
nor U4294 (N_4294,N_2125,N_2521);
or U4295 (N_4295,N_2674,N_2980);
nand U4296 (N_4296,N_3424,N_3327);
nand U4297 (N_4297,N_3572,N_3163);
nand U4298 (N_4298,N_2469,N_2376);
nand U4299 (N_4299,N_2010,N_3057);
or U4300 (N_4300,N_2070,N_2136);
nor U4301 (N_4301,N_2735,N_3317);
or U4302 (N_4302,N_3333,N_3630);
nand U4303 (N_4303,N_2940,N_3632);
or U4304 (N_4304,N_2668,N_3972);
nor U4305 (N_4305,N_3123,N_3332);
or U4306 (N_4306,N_2952,N_3078);
nand U4307 (N_4307,N_3631,N_3063);
or U4308 (N_4308,N_3061,N_2308);
or U4309 (N_4309,N_2309,N_2344);
nor U4310 (N_4310,N_3712,N_2584);
nand U4311 (N_4311,N_3264,N_2964);
nor U4312 (N_4312,N_3497,N_2625);
nand U4313 (N_4313,N_3155,N_2133);
or U4314 (N_4314,N_3844,N_3936);
nand U4315 (N_4315,N_2135,N_3374);
and U4316 (N_4316,N_2960,N_2736);
nand U4317 (N_4317,N_2654,N_2640);
nand U4318 (N_4318,N_3358,N_3176);
nor U4319 (N_4319,N_2459,N_2098);
nor U4320 (N_4320,N_3851,N_2152);
or U4321 (N_4321,N_2217,N_2958);
nand U4322 (N_4322,N_3149,N_3392);
or U4323 (N_4323,N_3859,N_2604);
or U4324 (N_4324,N_2845,N_3616);
or U4325 (N_4325,N_2685,N_2352);
nand U4326 (N_4326,N_2311,N_2779);
nor U4327 (N_4327,N_3810,N_2244);
nor U4328 (N_4328,N_2007,N_3903);
nand U4329 (N_4329,N_2693,N_2201);
nor U4330 (N_4330,N_3698,N_2113);
nor U4331 (N_4331,N_2998,N_3435);
or U4332 (N_4332,N_3878,N_3147);
or U4333 (N_4333,N_3129,N_3043);
and U4334 (N_4334,N_2100,N_2932);
xnor U4335 (N_4335,N_2619,N_2992);
or U4336 (N_4336,N_3469,N_2610);
or U4337 (N_4337,N_3431,N_2566);
and U4338 (N_4338,N_3278,N_3422);
or U4339 (N_4339,N_2870,N_3745);
and U4340 (N_4340,N_2419,N_2862);
nor U4341 (N_4341,N_3649,N_2294);
nor U4342 (N_4342,N_3476,N_3753);
and U4343 (N_4343,N_2232,N_3790);
and U4344 (N_4344,N_3639,N_3177);
or U4345 (N_4345,N_3250,N_3389);
nand U4346 (N_4346,N_2593,N_2463);
or U4347 (N_4347,N_3114,N_2233);
nand U4348 (N_4348,N_3444,N_3235);
nand U4349 (N_4349,N_2079,N_3414);
nor U4350 (N_4350,N_2666,N_2781);
and U4351 (N_4351,N_2497,N_2416);
nor U4352 (N_4352,N_3816,N_2170);
nor U4353 (N_4353,N_3786,N_3657);
and U4354 (N_4354,N_2523,N_3751);
and U4355 (N_4355,N_2336,N_2796);
nand U4356 (N_4356,N_3253,N_3561);
and U4357 (N_4357,N_2543,N_3814);
nand U4358 (N_4358,N_2406,N_2744);
and U4359 (N_4359,N_2991,N_2440);
nand U4360 (N_4360,N_2795,N_2713);
and U4361 (N_4361,N_2088,N_3819);
nand U4362 (N_4362,N_3118,N_3829);
nand U4363 (N_4363,N_2923,N_2354);
nand U4364 (N_4364,N_3989,N_2659);
xor U4365 (N_4365,N_2062,N_2003);
nand U4366 (N_4366,N_3499,N_3541);
nor U4367 (N_4367,N_3830,N_2750);
or U4368 (N_4368,N_2044,N_2635);
or U4369 (N_4369,N_3969,N_2682);
or U4370 (N_4370,N_2782,N_2679);
or U4371 (N_4371,N_3206,N_2008);
nand U4372 (N_4372,N_2212,N_2724);
nand U4373 (N_4373,N_3843,N_3388);
and U4374 (N_4374,N_2885,N_2225);
nand U4375 (N_4375,N_2196,N_3736);
and U4376 (N_4376,N_2230,N_3640);
or U4377 (N_4377,N_3303,N_2802);
nand U4378 (N_4378,N_3743,N_3680);
nor U4379 (N_4379,N_3576,N_3697);
and U4380 (N_4380,N_2409,N_3058);
nor U4381 (N_4381,N_2054,N_2536);
nand U4382 (N_4382,N_3092,N_2947);
or U4383 (N_4383,N_3115,N_3318);
and U4384 (N_4384,N_3241,N_2652);
nor U4385 (N_4385,N_2256,N_2511);
xor U4386 (N_4386,N_2160,N_3205);
or U4387 (N_4387,N_2016,N_2085);
nor U4388 (N_4388,N_2650,N_3659);
xor U4389 (N_4389,N_2517,N_3655);
and U4390 (N_4390,N_2259,N_2770);
or U4391 (N_4391,N_3300,N_2096);
or U4392 (N_4392,N_2594,N_3913);
or U4393 (N_4393,N_2246,N_3802);
or U4394 (N_4394,N_2253,N_2460);
nor U4395 (N_4395,N_2909,N_3172);
and U4396 (N_4396,N_2576,N_2898);
and U4397 (N_4397,N_3023,N_2051);
nor U4398 (N_4398,N_2774,N_3967);
or U4399 (N_4399,N_3554,N_2194);
nor U4400 (N_4400,N_3789,N_3919);
and U4401 (N_4401,N_3156,N_2848);
and U4402 (N_4402,N_2042,N_2264);
and U4403 (N_4403,N_3411,N_2734);
and U4404 (N_4404,N_3935,N_3105);
nand U4405 (N_4405,N_2038,N_2398);
nor U4406 (N_4406,N_2284,N_2814);
and U4407 (N_4407,N_3432,N_3885);
and U4408 (N_4408,N_2754,N_3644);
nor U4409 (N_4409,N_2144,N_2185);
nor U4410 (N_4410,N_3755,N_3321);
and U4411 (N_4411,N_2187,N_2423);
nand U4412 (N_4412,N_3872,N_3306);
nor U4413 (N_4413,N_3323,N_3532);
or U4414 (N_4414,N_2214,N_3847);
and U4415 (N_4415,N_2516,N_2213);
or U4416 (N_4416,N_3508,N_3180);
or U4417 (N_4417,N_3660,N_2198);
xnor U4418 (N_4418,N_3707,N_2758);
and U4419 (N_4419,N_2901,N_2930);
nand U4420 (N_4420,N_3240,N_2265);
nor U4421 (N_4421,N_3408,N_2068);
and U4422 (N_4422,N_3249,N_2306);
nand U4423 (N_4423,N_3384,N_3667);
nand U4424 (N_4424,N_2268,N_2394);
or U4425 (N_4425,N_2203,N_3443);
nor U4426 (N_4426,N_3347,N_3194);
and U4427 (N_4427,N_2464,N_3460);
and U4428 (N_4428,N_2622,N_3717);
nor U4429 (N_4429,N_3151,N_3803);
nand U4430 (N_4430,N_3289,N_3420);
and U4431 (N_4431,N_3041,N_3251);
nand U4432 (N_4432,N_3158,N_2101);
and U4433 (N_4433,N_3555,N_2660);
nor U4434 (N_4434,N_2494,N_2073);
nand U4435 (N_4435,N_3304,N_3490);
or U4436 (N_4436,N_2966,N_3439);
nor U4437 (N_4437,N_3257,N_2455);
nand U4438 (N_4438,N_2208,N_3925);
nand U4439 (N_4439,N_3603,N_2972);
or U4440 (N_4440,N_2335,N_3676);
nand U4441 (N_4441,N_2020,N_3970);
nand U4442 (N_4442,N_2646,N_2243);
and U4443 (N_4443,N_2698,N_2274);
nand U4444 (N_4444,N_2793,N_2526);
or U4445 (N_4445,N_3850,N_3085);
or U4446 (N_4446,N_3383,N_2675);
nand U4447 (N_4447,N_2383,N_2301);
and U4448 (N_4448,N_2437,N_2653);
and U4449 (N_4449,N_2815,N_3928);
or U4450 (N_4450,N_2533,N_3737);
or U4451 (N_4451,N_2450,N_2493);
nor U4452 (N_4452,N_2411,N_2747);
and U4453 (N_4453,N_3585,N_2742);
nand U4454 (N_4454,N_3142,N_3746);
or U4455 (N_4455,N_3725,N_2310);
or U4456 (N_4456,N_3769,N_3381);
nand U4457 (N_4457,N_3482,N_3701);
nor U4458 (N_4458,N_3731,N_3399);
nand U4459 (N_4459,N_3402,N_2226);
and U4460 (N_4460,N_3329,N_3921);
and U4461 (N_4461,N_3812,N_3307);
nand U4462 (N_4462,N_2946,N_3895);
or U4463 (N_4463,N_3578,N_3495);
or U4464 (N_4464,N_2182,N_3625);
and U4465 (N_4465,N_2300,N_2083);
and U4466 (N_4466,N_2738,N_2442);
or U4467 (N_4467,N_3276,N_3376);
nor U4468 (N_4468,N_2773,N_3471);
or U4469 (N_4469,N_3946,N_2763);
nor U4470 (N_4470,N_3213,N_2067);
nor U4471 (N_4471,N_3407,N_2714);
or U4472 (N_4472,N_2696,N_3463);
and U4473 (N_4473,N_2994,N_2145);
nand U4474 (N_4474,N_3184,N_3505);
nor U4475 (N_4475,N_3285,N_3613);
nand U4476 (N_4476,N_2942,N_2199);
nand U4477 (N_4477,N_3705,N_3297);
nor U4478 (N_4478,N_3782,N_3133);
and U4479 (N_4479,N_3001,N_2399);
or U4480 (N_4480,N_3088,N_3336);
and U4481 (N_4481,N_3540,N_3491);
nand U4482 (N_4482,N_3446,N_3030);
and U4483 (N_4483,N_2263,N_2809);
nand U4484 (N_4484,N_3863,N_2677);
and U4485 (N_4485,N_2937,N_3275);
nor U4486 (N_4486,N_2587,N_3102);
and U4487 (N_4487,N_2171,N_2039);
or U4488 (N_4488,N_3394,N_3441);
and U4489 (N_4489,N_3299,N_2837);
and U4490 (N_4490,N_2138,N_2803);
or U4491 (N_4491,N_3236,N_3985);
and U4492 (N_4492,N_2001,N_3367);
or U4493 (N_4493,N_3353,N_3464);
and U4494 (N_4494,N_3287,N_2669);
nor U4495 (N_4495,N_2178,N_2278);
or U4496 (N_4496,N_2119,N_2894);
or U4497 (N_4497,N_2603,N_2250);
nor U4498 (N_4498,N_2890,N_3898);
nand U4499 (N_4499,N_3917,N_2385);
and U4500 (N_4500,N_3437,N_3654);
nand U4501 (N_4501,N_3606,N_3127);
and U4502 (N_4502,N_3182,N_2897);
and U4503 (N_4503,N_3976,N_2328);
nand U4504 (N_4504,N_2287,N_3530);
nor U4505 (N_4505,N_3900,N_3750);
nor U4506 (N_4506,N_3447,N_3788);
nor U4507 (N_4507,N_2816,N_3890);
nand U4508 (N_4508,N_2118,N_2286);
or U4509 (N_4509,N_2189,N_3638);
nand U4510 (N_4510,N_2752,N_2639);
and U4511 (N_4511,N_2325,N_2030);
nor U4512 (N_4512,N_2616,N_3791);
nand U4513 (N_4513,N_2347,N_2505);
nand U4514 (N_4514,N_3529,N_2596);
or U4515 (N_4515,N_3196,N_3502);
nor U4516 (N_4516,N_3190,N_3764);
or U4517 (N_4517,N_2432,N_3762);
xnor U4518 (N_4518,N_3867,N_2448);
and U4519 (N_4519,N_2892,N_3097);
or U4520 (N_4520,N_2825,N_3633);
and U4521 (N_4521,N_2291,N_3915);
and U4522 (N_4522,N_3811,N_2760);
nor U4523 (N_4523,N_2720,N_3774);
or U4524 (N_4524,N_3775,N_2011);
and U4525 (N_4525,N_3186,N_3533);
nand U4526 (N_4526,N_2692,N_2351);
nand U4527 (N_4527,N_3134,N_3034);
or U4528 (N_4528,N_3525,N_2869);
or U4529 (N_4529,N_3113,N_3978);
and U4530 (N_4530,N_2858,N_2172);
and U4531 (N_4531,N_3808,N_2905);
and U4532 (N_4532,N_3889,N_3688);
nor U4533 (N_4533,N_3728,N_3461);
and U4534 (N_4534,N_2663,N_2181);
nor U4535 (N_4535,N_2812,N_2919);
nor U4536 (N_4536,N_2381,N_2207);
and U4537 (N_4537,N_3356,N_2530);
nor U4538 (N_4538,N_2153,N_2465);
nor U4539 (N_4539,N_2041,N_2767);
and U4540 (N_4540,N_3512,N_2034);
nor U4541 (N_4541,N_2065,N_3212);
and U4542 (N_4542,N_3965,N_3265);
nor U4543 (N_4543,N_3395,N_3570);
nand U4544 (N_4544,N_3494,N_2162);
nor U4545 (N_4545,N_3973,N_3187);
nand U4546 (N_4546,N_3436,N_2273);
and U4547 (N_4547,N_3661,N_3766);
nor U4548 (N_4548,N_3795,N_3448);
nand U4549 (N_4549,N_3901,N_3884);
nor U4550 (N_4550,N_3440,N_2297);
nor U4551 (N_4551,N_2982,N_3523);
or U4552 (N_4552,N_3799,N_2209);
nor U4553 (N_4553,N_3741,N_2518);
nor U4554 (N_4554,N_3596,N_3325);
nor U4555 (N_4555,N_2161,N_2987);
and U4556 (N_4556,N_3489,N_3908);
nor U4557 (N_4557,N_2550,N_3320);
or U4558 (N_4558,N_3998,N_2169);
nand U4559 (N_4559,N_3064,N_3493);
nor U4560 (N_4560,N_2818,N_3784);
nand U4561 (N_4561,N_3474,N_3588);
nor U4562 (N_4562,N_2320,N_2072);
nand U4563 (N_4563,N_2864,N_2024);
nand U4564 (N_4564,N_2087,N_3706);
nor U4565 (N_4565,N_3686,N_2613);
nor U4566 (N_4566,N_2865,N_2661);
nor U4567 (N_4567,N_3390,N_3503);
nand U4568 (N_4568,N_3807,N_3488);
nor U4569 (N_4569,N_3822,N_3744);
nor U4570 (N_4570,N_2561,N_2402);
nor U4571 (N_4571,N_3759,N_2591);
or U4572 (N_4572,N_2102,N_2601);
nor U4573 (N_4573,N_2219,N_3675);
or U4574 (N_4574,N_3871,N_3605);
or U4575 (N_4575,N_3480,N_2037);
nand U4576 (N_4576,N_2141,N_3362);
or U4577 (N_4577,N_2052,N_3486);
nand U4578 (N_4578,N_2955,N_2049);
nand U4579 (N_4579,N_3286,N_3637);
or U4580 (N_4580,N_3473,N_3971);
and U4581 (N_4581,N_3309,N_3423);
and U4582 (N_4582,N_3324,N_2915);
and U4583 (N_4583,N_3081,N_2954);
nor U4584 (N_4584,N_2021,N_2705);
and U4585 (N_4585,N_3067,N_2150);
nor U4586 (N_4586,N_3892,N_2384);
and U4587 (N_4587,N_3783,N_2838);
and U4588 (N_4588,N_3629,N_2944);
or U4589 (N_4589,N_2648,N_2850);
or U4590 (N_4590,N_2789,N_2534);
nand U4591 (N_4591,N_3963,N_3013);
nor U4592 (N_4592,N_2694,N_2849);
and U4593 (N_4593,N_2959,N_3283);
or U4594 (N_4594,N_2002,N_2784);
nand U4595 (N_4595,N_3990,N_3173);
nand U4596 (N_4596,N_3339,N_3054);
and U4597 (N_4597,N_3255,N_2971);
or U4598 (N_4598,N_2397,N_3342);
nor U4599 (N_4599,N_2123,N_2896);
and U4600 (N_4600,N_2708,N_2421);
or U4601 (N_4601,N_3361,N_3940);
nor U4602 (N_4602,N_3039,N_3375);
or U4603 (N_4603,N_3700,N_3542);
xor U4604 (N_4604,N_3442,N_2193);
nor U4605 (N_4605,N_3794,N_3636);
or U4606 (N_4606,N_2426,N_2753);
nand U4607 (N_4607,N_2095,N_2200);
and U4608 (N_4608,N_2725,N_2806);
nor U4609 (N_4609,N_2641,N_2191);
or U4610 (N_4610,N_3797,N_2321);
or U4611 (N_4611,N_2180,N_3366);
and U4612 (N_4612,N_3292,N_3600);
or U4613 (N_4613,N_2470,N_3237);
or U4614 (N_4614,N_2681,N_3560);
and U4615 (N_4615,N_3036,N_3028);
and U4616 (N_4616,N_2476,N_2404);
or U4617 (N_4617,N_2028,N_3720);
or U4618 (N_4618,N_3221,N_3311);
nor U4619 (N_4619,N_2777,N_3179);
nand U4620 (N_4620,N_2433,N_2877);
nand U4621 (N_4621,N_2055,N_3756);
nor U4622 (N_4622,N_2914,N_3767);
or U4623 (N_4623,N_2380,N_2215);
nand U4624 (N_4624,N_2671,N_3122);
nor U4625 (N_4625,N_2305,N_2184);
nor U4626 (N_4626,N_3370,N_2019);
xnor U4627 (N_4627,N_2401,N_2275);
nand U4628 (N_4628,N_2468,N_3839);
and U4629 (N_4629,N_2454,N_3405);
or U4630 (N_4630,N_3548,N_2204);
nor U4631 (N_4631,N_3449,N_3224);
or U4632 (N_4632,N_2839,N_2488);
nor U4633 (N_4633,N_3838,N_3458);
nor U4634 (N_4634,N_2260,N_2471);
nor U4635 (N_4635,N_3232,N_2337);
and U4636 (N_4636,N_2313,N_2702);
nor U4637 (N_4637,N_2176,N_3996);
nor U4638 (N_4638,N_3277,N_3856);
or U4639 (N_4639,N_2424,N_3568);
xnor U4640 (N_4640,N_2626,N_3804);
nor U4641 (N_4641,N_3724,N_2120);
or U4642 (N_4642,N_2137,N_2314);
nand U4643 (N_4643,N_2612,N_2478);
nor U4644 (N_4644,N_3582,N_2581);
nand U4645 (N_4645,N_2392,N_2104);
nor U4646 (N_4646,N_3864,N_2422);
nor U4647 (N_4647,N_3012,N_2840);
nor U4648 (N_4648,N_2835,N_3942);
or U4649 (N_4649,N_2853,N_2918);
nor U4650 (N_4650,N_2164,N_3465);
and U4651 (N_4651,N_2282,N_3410);
nor U4652 (N_4652,N_2174,N_2315);
or U4653 (N_4653,N_2388,N_3922);
or U4654 (N_4654,N_3780,N_2069);
nor U4655 (N_4655,N_2883,N_2569);
nor U4656 (N_4656,N_3670,N_2740);
nor U4657 (N_4657,N_2778,N_3252);
or U4658 (N_4658,N_2032,N_2749);
and U4659 (N_4659,N_2733,N_3316);
nand U4660 (N_4660,N_2452,N_2624);
and U4661 (N_4661,N_2636,N_2643);
and U4662 (N_4662,N_2248,N_2031);
or U4663 (N_4663,N_2574,N_3648);
or U4664 (N_4664,N_2304,N_3601);
nand U4665 (N_4665,N_2216,N_3787);
and U4666 (N_4666,N_2249,N_2811);
and U4667 (N_4667,N_3669,N_3567);
and U4668 (N_4668,N_2928,N_3006);
or U4669 (N_4669,N_3368,N_2844);
nand U4670 (N_4670,N_2710,N_3161);
nor U4671 (N_4671,N_3894,N_2236);
nor U4672 (N_4672,N_3599,N_3293);
and U4673 (N_4673,N_3656,N_2086);
nand U4674 (N_4674,N_2701,N_3430);
nor U4675 (N_4675,N_3330,N_3418);
nand U4676 (N_4676,N_2413,N_3425);
and U4677 (N_4677,N_3008,N_3796);
and U4678 (N_4678,N_2415,N_2769);
nand U4679 (N_4679,N_2241,N_3693);
and U4680 (N_4680,N_3982,N_2941);
nor U4681 (N_4681,N_2756,N_3059);
nor U4682 (N_4682,N_3020,N_2629);
nand U4683 (N_4683,N_2555,N_2081);
xor U4684 (N_4684,N_2283,N_2842);
or U4685 (N_4685,N_2091,N_3298);
nor U4686 (N_4686,N_2132,N_3823);
and U4687 (N_4687,N_2801,N_3779);
and U4688 (N_4688,N_2358,N_2084);
nand U4689 (N_4689,N_3522,N_2546);
or U4690 (N_4690,N_3214,N_3905);
nor U4691 (N_4691,N_2369,N_2092);
or U4692 (N_4692,N_2445,N_2879);
nor U4693 (N_4693,N_2990,N_3881);
nand U4694 (N_4694,N_3228,N_3106);
nor U4695 (N_4695,N_2642,N_2595);
nand U4696 (N_4696,N_2721,N_3302);
nor U4697 (N_4697,N_3577,N_3748);
nand U4698 (N_4698,N_3608,N_2080);
and U4699 (N_4699,N_2993,N_2552);
or U4700 (N_4700,N_2403,N_2730);
nand U4701 (N_4701,N_2775,N_2611);
nand U4702 (N_4702,N_2647,N_2847);
nand U4703 (N_4703,N_3072,N_2891);
or U4704 (N_4704,N_3404,N_2645);
nor U4705 (N_4705,N_3259,N_2797);
xnor U4706 (N_4706,N_2542,N_3197);
and U4707 (N_4707,N_2843,N_2969);
nand U4708 (N_4708,N_2547,N_2348);
or U4709 (N_4709,N_3385,N_3139);
nand U4710 (N_4710,N_3222,N_2644);
and U4711 (N_4711,N_3359,N_2539);
and U4712 (N_4712,N_2945,N_3682);
nand U4713 (N_4713,N_3513,N_3729);
nor U4714 (N_4714,N_3604,N_3401);
nor U4715 (N_4715,N_2794,N_2105);
and U4716 (N_4716,N_3344,N_3263);
or U4717 (N_4717,N_2951,N_2528);
and U4718 (N_4718,N_2799,N_3939);
nand U4719 (N_4719,N_2420,N_3718);
nand U4720 (N_4720,N_3260,N_2108);
and U4721 (N_4721,N_3509,N_2822);
and U4722 (N_4722,N_3037,N_3010);
nand U4723 (N_4723,N_3987,N_2127);
and U4724 (N_4724,N_3853,N_2307);
nand U4725 (N_4725,N_3620,N_2589);
or U4726 (N_4726,N_2234,N_3672);
or U4727 (N_4727,N_2343,N_2556);
or U4728 (N_4728,N_3031,N_3386);
and U4729 (N_4729,N_2520,N_3426);
nor U4730 (N_4730,N_3950,N_3246);
nand U4731 (N_4731,N_3234,N_2115);
or U4732 (N_4732,N_3778,N_2159);
nand U4733 (N_4733,N_3372,N_3352);
and U4734 (N_4734,N_3200,N_3904);
nand U4735 (N_4735,N_3994,N_2627);
nor U4736 (N_4736,N_3261,N_2887);
nor U4737 (N_4737,N_2934,N_3849);
and U4738 (N_4738,N_2027,N_2338);
nand U4739 (N_4739,N_3869,N_3288);
nor U4740 (N_4740,N_2551,N_2503);
and U4741 (N_4741,N_2746,N_3136);
or U4742 (N_4742,N_2046,N_3242);
and U4743 (N_4743,N_3053,N_3048);
nor U4744 (N_4744,N_2443,N_3684);
nand U4745 (N_4745,N_3840,N_2963);
nand U4746 (N_4746,N_3897,N_2868);
and U4747 (N_4747,N_2418,N_2441);
and U4748 (N_4748,N_2997,N_3709);
nand U4749 (N_4749,N_2235,N_2807);
and U4750 (N_4750,N_2863,N_2238);
nand U4751 (N_4751,N_2618,N_3500);
and U4752 (N_4752,N_2066,N_3809);
or U4753 (N_4753,N_2851,N_2228);
or U4754 (N_4754,N_3722,N_3827);
and U4755 (N_4755,N_2029,N_3831);
nand U4756 (N_4756,N_3313,N_3338);
nand U4757 (N_4757,N_2218,N_3573);
nand U4758 (N_4758,N_2785,N_2496);
or U4759 (N_4759,N_2902,N_3274);
or U4760 (N_4760,N_3191,N_2579);
nor U4761 (N_4761,N_3983,N_3642);
and U4762 (N_4762,N_2549,N_3501);
nor U4763 (N_4763,N_2608,N_3227);
nor U4764 (N_4764,N_2507,N_3125);
or U4765 (N_4765,N_2583,N_3785);
nand U4766 (N_4766,N_3826,N_2323);
and U4767 (N_4767,N_3223,N_2522);
or U4768 (N_4768,N_2370,N_2786);
or U4769 (N_4769,N_2525,N_3610);
nor U4770 (N_4770,N_2377,N_2935);
nor U4771 (N_4771,N_2655,N_2766);
and U4772 (N_4772,N_3663,N_3116);
nand U4773 (N_4773,N_3598,N_3929);
and U4774 (N_4774,N_2968,N_2707);
and U4775 (N_4775,N_2757,N_3569);
nand U4776 (N_4776,N_2355,N_3079);
and U4777 (N_4777,N_3979,N_3665);
nand U4778 (N_4778,N_2290,N_3566);
nor U4779 (N_4779,N_3406,N_2834);
and U4780 (N_4780,N_2154,N_3185);
nand U4781 (N_4781,N_2871,N_2817);
nand U4782 (N_4782,N_3584,N_3713);
and U4783 (N_4783,N_2727,N_3687);
nor U4784 (N_4784,N_3876,N_2004);
or U4785 (N_4785,N_3266,N_3920);
nand U4786 (N_4786,N_3349,N_2285);
nand U4787 (N_4787,N_3099,N_2732);
and U4788 (N_4788,N_2988,N_3714);
and U4789 (N_4789,N_2359,N_2900);
nand U4790 (N_4790,N_2949,N_3535);
nand U4791 (N_4791,N_3517,N_3587);
nor U4792 (N_4792,N_3948,N_2367);
and U4793 (N_4793,N_3363,N_2499);
nand U4794 (N_4794,N_3806,N_3621);
and U4795 (N_4795,N_2873,N_3153);
nand U4796 (N_4796,N_3793,N_2875);
nor U4797 (N_4797,N_2854,N_3238);
or U4798 (N_4798,N_2339,N_3821);
or U4799 (N_4799,N_2741,N_3666);
nand U4800 (N_4800,N_2296,N_2220);
nand U4801 (N_4801,N_3690,N_2317);
and U4802 (N_4802,N_2829,N_2107);
and U4803 (N_4803,N_2129,N_3131);
nor U4804 (N_4804,N_3091,N_2739);
or U4805 (N_4805,N_2057,N_3914);
or U4806 (N_4806,N_2018,N_3104);
and U4807 (N_4807,N_2506,N_3354);
nor U4808 (N_4808,N_2434,N_3960);
nor U4809 (N_4809,N_2363,N_3089);
or U4810 (N_4810,N_3977,N_2904);
and U4811 (N_4811,N_2379,N_3549);
nor U4812 (N_4812,N_3527,N_3071);
and U4813 (N_4813,N_3609,N_3357);
nand U4814 (N_4814,N_3022,N_2823);
or U4815 (N_4815,N_2617,N_3607);
nand U4816 (N_4816,N_3622,N_2251);
nor U4817 (N_4817,N_2709,N_2390);
nor U4818 (N_4818,N_3218,N_2657);
and U4819 (N_4819,N_3040,N_2938);
nor U4820 (N_4820,N_3553,N_2605);
nor U4821 (N_4821,N_3992,N_3248);
nor U4822 (N_4822,N_3226,N_3524);
nand U4823 (N_4823,N_3882,N_3683);
or U4824 (N_4824,N_3945,N_2614);
and U4825 (N_4825,N_2712,N_3801);
and U4826 (N_4826,N_3270,N_2009);
nor U4827 (N_4827,N_2146,N_2210);
nand U4828 (N_4828,N_2015,N_2059);
and U4829 (N_4829,N_3594,N_3291);
nand U4830 (N_4830,N_3537,N_2179);
nand U4831 (N_4831,N_2186,N_3518);
and U4832 (N_4832,N_3646,N_3045);
nand U4833 (N_4833,N_3322,N_2446);
and U4834 (N_4834,N_2242,N_2704);
nor U4835 (N_4835,N_2475,N_2519);
or U4836 (N_4836,N_3077,N_2447);
or U4837 (N_4837,N_2886,N_2288);
nand U4838 (N_4838,N_2112,N_2852);
and U4839 (N_4839,N_2620,N_2538);
or U4840 (N_4840,N_3927,N_3860);
or U4841 (N_4841,N_2148,N_3029);
nand U4842 (N_4842,N_3035,N_3229);
nor U4843 (N_4843,N_3589,N_3910);
nand U4844 (N_4844,N_3146,N_3536);
nor U4845 (N_4845,N_3583,N_3409);
and U4846 (N_4846,N_3893,N_2262);
and U4847 (N_4847,N_2861,N_3117);
and U4848 (N_4848,N_2588,N_2116);
nor U4849 (N_4849,N_3702,N_2931);
nor U4850 (N_4850,N_3930,N_3438);
nor U4851 (N_4851,N_2783,N_2474);
and U4852 (N_4852,N_2509,N_3415);
and U4853 (N_4853,N_2254,N_2040);
or U4854 (N_4854,N_3719,N_2638);
and U4855 (N_4855,N_2240,N_2163);
and U4856 (N_4856,N_2996,N_2512);
nor U4857 (N_4857,N_2025,N_3169);
and U4858 (N_4858,N_3060,N_3873);
nor U4859 (N_4859,N_3857,N_2211);
and U4860 (N_4860,N_2557,N_2772);
or U4861 (N_4861,N_3868,N_3340);
or U4862 (N_4862,N_3592,N_3662);
or U4863 (N_4863,N_3763,N_2805);
or U4864 (N_4864,N_2410,N_3975);
and U4865 (N_4865,N_2106,N_3556);
nor U4866 (N_4866,N_3165,N_2826);
nand U4867 (N_4867,N_3916,N_2787);
and U4868 (N_4868,N_2771,N_2033);
or U4869 (N_4869,N_3445,N_2005);
nand U4870 (N_4870,N_3065,N_3634);
and U4871 (N_4871,N_2048,N_2327);
or U4872 (N_4872,N_3883,N_2456);
or U4873 (N_4873,N_3225,N_3691);
nor U4874 (N_4874,N_3993,N_3749);
or U4875 (N_4875,N_2917,N_2017);
nor U4876 (N_4876,N_2330,N_3761);
and U4877 (N_4877,N_3284,N_2831);
or U4878 (N_4878,N_3538,N_3152);
nor U4879 (N_4879,N_3326,N_2856);
or U4880 (N_4880,N_3201,N_2061);
and U4881 (N_4881,N_2859,N_2544);
nor U4882 (N_4882,N_2731,N_2158);
nor U4883 (N_4883,N_3267,N_3962);
or U4884 (N_4884,N_2553,N_3207);
or U4885 (N_4885,N_3544,N_2691);
xor U4886 (N_4886,N_3906,N_2289);
and U4887 (N_4887,N_3721,N_2056);
nand U4888 (N_4888,N_3760,N_2430);
and U4889 (N_4889,N_2597,N_2462);
nor U4890 (N_4890,N_2780,N_2393);
and U4891 (N_4891,N_3519,N_2821);
or U4892 (N_4892,N_2387,N_3624);
nand U4893 (N_4893,N_3073,N_3103);
nor U4894 (N_4894,N_2134,N_2878);
nor U4895 (N_4895,N_3365,N_3507);
nor U4896 (N_4896,N_3653,N_2482);
nor U4897 (N_4897,N_3433,N_3781);
and U4898 (N_4898,N_2562,N_3003);
nand U4899 (N_4899,N_2427,N_3754);
and U4900 (N_4900,N_3160,N_2578);
or U4901 (N_4901,N_2857,N_2223);
nand U4902 (N_4902,N_3981,N_2319);
or U4903 (N_4903,N_2378,N_3593);
and U4904 (N_4904,N_3511,N_3132);
nand U4905 (N_4905,N_3986,N_3369);
and U4906 (N_4906,N_3833,N_2368);
nand U4907 (N_4907,N_3564,N_3834);
nand U4908 (N_4908,N_3738,N_2800);
and U4909 (N_4909,N_2114,N_2580);
nand U4910 (N_4910,N_3574,N_3695);
nor U4911 (N_4911,N_3350,N_2157);
nand U4912 (N_4912,N_2776,N_3377);
nor U4913 (N_4913,N_3087,N_3848);
nor U4914 (N_4914,N_2277,N_2684);
or U4915 (N_4915,N_2293,N_3387);
nor U4916 (N_4916,N_2139,N_3137);
and U4917 (N_4917,N_3412,N_3271);
nor U4918 (N_4918,N_3331,N_3955);
or U4919 (N_4919,N_2224,N_3886);
or U4920 (N_4920,N_2575,N_3959);
nand U4921 (N_4921,N_3947,N_2933);
nor U4922 (N_4922,N_2585,N_3571);
nand U4923 (N_4923,N_2961,N_3101);
nand U4924 (N_4924,N_2375,N_2237);
nand U4925 (N_4925,N_2532,N_2071);
or U4926 (N_4926,N_3397,N_2175);
or U4927 (N_4927,N_2867,N_3668);
nand U4928 (N_4928,N_2676,N_2190);
nor U4929 (N_4929,N_2689,N_3880);
nand U4930 (N_4930,N_2895,N_3183);
nor U4931 (N_4931,N_2962,N_2939);
nand U4932 (N_4932,N_2529,N_2527);
and U4933 (N_4933,N_3953,N_2035);
nor U4934 (N_4934,N_2491,N_2366);
nand U4935 (N_4935,N_2665,N_2451);
nand U4936 (N_4936,N_2149,N_3378);
or U4937 (N_4937,N_3421,N_2222);
or U4938 (N_4938,N_2889,N_3429);
nor U4939 (N_4939,N_2396,N_2128);
and U4940 (N_4940,N_3628,N_3918);
nand U4941 (N_4941,N_2882,N_3510);
or U4942 (N_4942,N_2916,N_2670);
nand U4943 (N_4943,N_2673,N_3143);
nor U4944 (N_4944,N_2484,N_2813);
nor U4945 (N_4945,N_2412,N_3128);
and U4946 (N_4946,N_2318,N_3462);
nand U4947 (N_4947,N_2841,N_2686);
nor U4948 (N_4948,N_2103,N_2173);
nand U4949 (N_4949,N_3758,N_3991);
nand U4950 (N_4950,N_3019,N_3086);
nand U4951 (N_4951,N_2545,N_2082);
or U4952 (N_4952,N_3314,N_3602);
and U4953 (N_4953,N_3531,N_3837);
or U4954 (N_4954,N_2473,N_2633);
or U4955 (N_4955,N_2751,N_3694);
or U4956 (N_4956,N_3611,N_2461);
or U4957 (N_4957,N_2365,N_2202);
and U4958 (N_4958,N_3879,N_3076);
or U4959 (N_4959,N_2272,N_2090);
nand U4960 (N_4960,N_2977,N_2606);
or U4961 (N_4961,N_2342,N_2719);
or U4962 (N_4962,N_3110,N_3413);
nand U4963 (N_4963,N_3559,N_2929);
nor U4964 (N_4964,N_2598,N_3148);
or U4965 (N_4965,N_2899,N_2687);
and U4966 (N_4966,N_2582,N_2957);
nand U4967 (N_4967,N_2715,N_3273);
nor U4968 (N_4968,N_3726,N_3961);
and U4969 (N_4969,N_3181,N_3403);
nand U4970 (N_4970,N_3980,N_3154);
or U4971 (N_4971,N_3974,N_3581);
or U4972 (N_4972,N_3643,N_2121);
nand U4973 (N_4973,N_2976,N_3954);
nor U4974 (N_4974,N_3521,N_3704);
nor U4975 (N_4975,N_2973,N_3842);
and U4976 (N_4976,N_2094,N_2349);
nand U4977 (N_4977,N_3130,N_3096);
nor U4978 (N_4978,N_2745,N_3579);
nor U4979 (N_4979,N_2053,N_3703);
nand U4980 (N_4980,N_2722,N_3671);
nand U4981 (N_4981,N_2600,N_2322);
and U4982 (N_4982,N_3044,N_2312);
nor U4983 (N_4983,N_2974,N_3107);
nor U4984 (N_4984,N_3360,N_3958);
nand U4985 (N_4985,N_2076,N_2269);
nand U4986 (N_4986,N_3484,N_2126);
nor U4987 (N_4987,N_2872,N_3014);
nand U4988 (N_4988,N_2602,N_3312);
nand U4989 (N_4989,N_2261,N_2936);
and U4990 (N_4990,N_2489,N_3933);
nand U4991 (N_4991,N_2706,N_2502);
nand U4992 (N_4992,N_3457,N_3492);
nand U4993 (N_4993,N_2466,N_2111);
nor U4994 (N_4994,N_3005,N_2391);
nor U4995 (N_4995,N_3000,N_3855);
and U4996 (N_4996,N_3380,N_2903);
and U4997 (N_4997,N_2302,N_2036);
nor U4998 (N_4998,N_2255,N_2695);
nor U4999 (N_4999,N_2984,N_3481);
nor U5000 (N_5000,N_3438,N_2310);
nand U5001 (N_5001,N_3794,N_2667);
or U5002 (N_5002,N_3286,N_3925);
nor U5003 (N_5003,N_3730,N_2695);
nor U5004 (N_5004,N_2354,N_3675);
nand U5005 (N_5005,N_3663,N_3192);
xnor U5006 (N_5006,N_2804,N_2922);
and U5007 (N_5007,N_2527,N_3014);
or U5008 (N_5008,N_2028,N_2501);
or U5009 (N_5009,N_2012,N_2998);
xnor U5010 (N_5010,N_3041,N_2515);
or U5011 (N_5011,N_3348,N_3914);
nand U5012 (N_5012,N_2652,N_2347);
or U5013 (N_5013,N_2926,N_2514);
or U5014 (N_5014,N_2576,N_2770);
nand U5015 (N_5015,N_2107,N_3027);
and U5016 (N_5016,N_3536,N_3280);
or U5017 (N_5017,N_3750,N_2523);
or U5018 (N_5018,N_3148,N_2768);
nand U5019 (N_5019,N_3612,N_2545);
and U5020 (N_5020,N_3722,N_2418);
or U5021 (N_5021,N_3139,N_2638);
or U5022 (N_5022,N_3297,N_3929);
or U5023 (N_5023,N_2489,N_2110);
or U5024 (N_5024,N_3793,N_3004);
nor U5025 (N_5025,N_3046,N_3984);
nand U5026 (N_5026,N_3492,N_2139);
nand U5027 (N_5027,N_2696,N_3622);
or U5028 (N_5028,N_2381,N_2213);
nand U5029 (N_5029,N_2749,N_3182);
and U5030 (N_5030,N_2219,N_3592);
nor U5031 (N_5031,N_2112,N_2219);
xor U5032 (N_5032,N_2764,N_3465);
nand U5033 (N_5033,N_3935,N_3896);
and U5034 (N_5034,N_3748,N_2662);
nor U5035 (N_5035,N_3868,N_2676);
nor U5036 (N_5036,N_2778,N_2295);
or U5037 (N_5037,N_3737,N_3245);
and U5038 (N_5038,N_3166,N_3672);
nor U5039 (N_5039,N_2848,N_3117);
or U5040 (N_5040,N_3536,N_3764);
xor U5041 (N_5041,N_3703,N_3259);
nor U5042 (N_5042,N_2030,N_2804);
nand U5043 (N_5043,N_3330,N_3374);
nor U5044 (N_5044,N_3665,N_3637);
and U5045 (N_5045,N_2185,N_2155);
nor U5046 (N_5046,N_2709,N_3327);
nor U5047 (N_5047,N_2030,N_2781);
or U5048 (N_5048,N_2758,N_2566);
nor U5049 (N_5049,N_2147,N_2258);
or U5050 (N_5050,N_3566,N_2085);
nor U5051 (N_5051,N_3880,N_3624);
and U5052 (N_5052,N_3416,N_2171);
and U5053 (N_5053,N_3141,N_2962);
nor U5054 (N_5054,N_3259,N_2231);
and U5055 (N_5055,N_2977,N_2171);
or U5056 (N_5056,N_2652,N_2255);
nand U5057 (N_5057,N_3405,N_3421);
and U5058 (N_5058,N_2667,N_2751);
or U5059 (N_5059,N_3781,N_2893);
and U5060 (N_5060,N_2964,N_3763);
nor U5061 (N_5061,N_3915,N_2985);
or U5062 (N_5062,N_2506,N_3872);
nor U5063 (N_5063,N_2668,N_2091);
and U5064 (N_5064,N_2715,N_2632);
and U5065 (N_5065,N_3710,N_3178);
nor U5066 (N_5066,N_2240,N_3628);
or U5067 (N_5067,N_3661,N_2647);
nand U5068 (N_5068,N_3163,N_2268);
nor U5069 (N_5069,N_2552,N_2335);
nor U5070 (N_5070,N_3261,N_2291);
or U5071 (N_5071,N_2522,N_2644);
nand U5072 (N_5072,N_2664,N_2507);
nand U5073 (N_5073,N_3140,N_3208);
or U5074 (N_5074,N_3030,N_3279);
nand U5075 (N_5075,N_3682,N_2930);
nor U5076 (N_5076,N_3888,N_3087);
and U5077 (N_5077,N_2987,N_2966);
nand U5078 (N_5078,N_2219,N_2637);
or U5079 (N_5079,N_2596,N_2885);
and U5080 (N_5080,N_2269,N_2339);
or U5081 (N_5081,N_2795,N_2408);
and U5082 (N_5082,N_3593,N_2117);
and U5083 (N_5083,N_3725,N_2470);
and U5084 (N_5084,N_2283,N_2163);
nand U5085 (N_5085,N_3931,N_3249);
or U5086 (N_5086,N_2686,N_2570);
nor U5087 (N_5087,N_3227,N_2983);
or U5088 (N_5088,N_2189,N_2980);
nand U5089 (N_5089,N_2526,N_2091);
or U5090 (N_5090,N_2966,N_2997);
or U5091 (N_5091,N_2499,N_2950);
nand U5092 (N_5092,N_2521,N_3629);
and U5093 (N_5093,N_3292,N_2693);
nor U5094 (N_5094,N_3136,N_2391);
and U5095 (N_5095,N_3935,N_2791);
and U5096 (N_5096,N_3809,N_3424);
nand U5097 (N_5097,N_2788,N_2409);
nor U5098 (N_5098,N_3658,N_3196);
nor U5099 (N_5099,N_2450,N_2644);
nor U5100 (N_5100,N_2153,N_3517);
and U5101 (N_5101,N_2405,N_3045);
and U5102 (N_5102,N_2293,N_2239);
nor U5103 (N_5103,N_3955,N_3686);
and U5104 (N_5104,N_2572,N_2819);
and U5105 (N_5105,N_3712,N_2950);
nand U5106 (N_5106,N_3271,N_3518);
or U5107 (N_5107,N_2065,N_3382);
nor U5108 (N_5108,N_2298,N_3901);
nor U5109 (N_5109,N_3349,N_3637);
nor U5110 (N_5110,N_3596,N_2471);
nand U5111 (N_5111,N_3492,N_3831);
or U5112 (N_5112,N_2520,N_3941);
or U5113 (N_5113,N_3567,N_3007);
nand U5114 (N_5114,N_3394,N_3885);
nand U5115 (N_5115,N_2510,N_2868);
nor U5116 (N_5116,N_3972,N_2053);
nor U5117 (N_5117,N_3773,N_2928);
nand U5118 (N_5118,N_2579,N_3133);
nand U5119 (N_5119,N_2488,N_2576);
or U5120 (N_5120,N_2197,N_3526);
nor U5121 (N_5121,N_2418,N_2711);
nand U5122 (N_5122,N_3044,N_3917);
nor U5123 (N_5123,N_3329,N_2588);
and U5124 (N_5124,N_3267,N_2408);
nor U5125 (N_5125,N_2845,N_3690);
nand U5126 (N_5126,N_3657,N_3648);
nand U5127 (N_5127,N_3576,N_3711);
nor U5128 (N_5128,N_3725,N_3767);
nor U5129 (N_5129,N_3514,N_3973);
or U5130 (N_5130,N_3810,N_3560);
and U5131 (N_5131,N_2283,N_2307);
or U5132 (N_5132,N_3529,N_2769);
nand U5133 (N_5133,N_3981,N_2591);
or U5134 (N_5134,N_3556,N_3951);
nand U5135 (N_5135,N_3772,N_2390);
and U5136 (N_5136,N_3004,N_3199);
nor U5137 (N_5137,N_3348,N_3189);
or U5138 (N_5138,N_3293,N_3534);
and U5139 (N_5139,N_2461,N_2000);
and U5140 (N_5140,N_2672,N_2226);
nand U5141 (N_5141,N_3749,N_3223);
nand U5142 (N_5142,N_3033,N_3163);
and U5143 (N_5143,N_2607,N_2165);
nor U5144 (N_5144,N_2365,N_3334);
and U5145 (N_5145,N_2073,N_2732);
or U5146 (N_5146,N_2166,N_2110);
or U5147 (N_5147,N_2848,N_2949);
nor U5148 (N_5148,N_3368,N_3998);
nand U5149 (N_5149,N_2444,N_3190);
and U5150 (N_5150,N_2902,N_3303);
or U5151 (N_5151,N_2636,N_3087);
nand U5152 (N_5152,N_2397,N_3409);
nand U5153 (N_5153,N_2553,N_2297);
and U5154 (N_5154,N_3836,N_3662);
nand U5155 (N_5155,N_2722,N_2409);
xnor U5156 (N_5156,N_2373,N_3135);
and U5157 (N_5157,N_3307,N_2326);
nand U5158 (N_5158,N_3527,N_3895);
and U5159 (N_5159,N_3603,N_2864);
nand U5160 (N_5160,N_3787,N_2602);
nor U5161 (N_5161,N_3427,N_2718);
nor U5162 (N_5162,N_3226,N_2152);
or U5163 (N_5163,N_3693,N_2819);
or U5164 (N_5164,N_3346,N_2811);
nand U5165 (N_5165,N_2778,N_3489);
nor U5166 (N_5166,N_3775,N_2821);
or U5167 (N_5167,N_2349,N_3682);
nand U5168 (N_5168,N_3537,N_3105);
nand U5169 (N_5169,N_2387,N_2766);
nand U5170 (N_5170,N_2308,N_3510);
nand U5171 (N_5171,N_2195,N_3616);
nand U5172 (N_5172,N_2738,N_2765);
and U5173 (N_5173,N_2010,N_3854);
or U5174 (N_5174,N_2459,N_3429);
nand U5175 (N_5175,N_2129,N_2111);
nand U5176 (N_5176,N_2723,N_3358);
nor U5177 (N_5177,N_2384,N_3214);
and U5178 (N_5178,N_3115,N_2312);
and U5179 (N_5179,N_2497,N_2590);
or U5180 (N_5180,N_3593,N_2978);
or U5181 (N_5181,N_3637,N_2125);
nand U5182 (N_5182,N_2992,N_3513);
nor U5183 (N_5183,N_2709,N_2359);
nor U5184 (N_5184,N_2549,N_2507);
nor U5185 (N_5185,N_2154,N_3133);
and U5186 (N_5186,N_2320,N_3617);
or U5187 (N_5187,N_2802,N_2421);
or U5188 (N_5188,N_2545,N_2255);
and U5189 (N_5189,N_3424,N_2552);
nor U5190 (N_5190,N_2037,N_2080);
nand U5191 (N_5191,N_3424,N_3014);
nand U5192 (N_5192,N_3863,N_3073);
nor U5193 (N_5193,N_2609,N_3686);
nand U5194 (N_5194,N_2459,N_3257);
and U5195 (N_5195,N_3913,N_2744);
nor U5196 (N_5196,N_3888,N_2547);
or U5197 (N_5197,N_2062,N_2385);
nand U5198 (N_5198,N_3475,N_2095);
or U5199 (N_5199,N_2723,N_2160);
nand U5200 (N_5200,N_3998,N_3324);
and U5201 (N_5201,N_2108,N_3321);
or U5202 (N_5202,N_3387,N_3384);
and U5203 (N_5203,N_2047,N_2585);
nand U5204 (N_5204,N_3271,N_3801);
and U5205 (N_5205,N_3156,N_2556);
and U5206 (N_5206,N_3311,N_2703);
or U5207 (N_5207,N_3130,N_3170);
nand U5208 (N_5208,N_3470,N_3315);
nor U5209 (N_5209,N_2543,N_3516);
nor U5210 (N_5210,N_2948,N_2095);
or U5211 (N_5211,N_3875,N_2983);
nand U5212 (N_5212,N_2627,N_2436);
and U5213 (N_5213,N_2214,N_2564);
nor U5214 (N_5214,N_3076,N_2769);
xor U5215 (N_5215,N_2587,N_3678);
nor U5216 (N_5216,N_2135,N_3042);
nor U5217 (N_5217,N_3157,N_3948);
and U5218 (N_5218,N_3461,N_3294);
nor U5219 (N_5219,N_2492,N_2191);
nor U5220 (N_5220,N_3497,N_2671);
or U5221 (N_5221,N_3531,N_2577);
or U5222 (N_5222,N_2235,N_2262);
or U5223 (N_5223,N_2577,N_2913);
nor U5224 (N_5224,N_2380,N_2349);
and U5225 (N_5225,N_2958,N_2396);
or U5226 (N_5226,N_3960,N_2186);
or U5227 (N_5227,N_3928,N_2758);
or U5228 (N_5228,N_3556,N_3670);
or U5229 (N_5229,N_3196,N_3781);
nand U5230 (N_5230,N_2230,N_3353);
or U5231 (N_5231,N_3420,N_2613);
nor U5232 (N_5232,N_3441,N_2744);
or U5233 (N_5233,N_3522,N_2926);
nor U5234 (N_5234,N_2187,N_2058);
nand U5235 (N_5235,N_2749,N_3662);
nand U5236 (N_5236,N_3658,N_3434);
nand U5237 (N_5237,N_2615,N_2832);
nand U5238 (N_5238,N_2460,N_2812);
nand U5239 (N_5239,N_2884,N_3735);
or U5240 (N_5240,N_3388,N_3302);
or U5241 (N_5241,N_2686,N_2429);
nor U5242 (N_5242,N_2874,N_3427);
and U5243 (N_5243,N_3276,N_3565);
and U5244 (N_5244,N_3973,N_2655);
nand U5245 (N_5245,N_3138,N_2609);
or U5246 (N_5246,N_2083,N_2332);
xor U5247 (N_5247,N_2816,N_2264);
or U5248 (N_5248,N_2451,N_2575);
or U5249 (N_5249,N_2733,N_3294);
nand U5250 (N_5250,N_2333,N_2113);
nand U5251 (N_5251,N_2551,N_3938);
or U5252 (N_5252,N_2526,N_2461);
and U5253 (N_5253,N_3724,N_2565);
or U5254 (N_5254,N_3145,N_3504);
or U5255 (N_5255,N_2469,N_2488);
or U5256 (N_5256,N_3775,N_2383);
or U5257 (N_5257,N_3073,N_2729);
or U5258 (N_5258,N_2109,N_2209);
nor U5259 (N_5259,N_3990,N_2498);
nand U5260 (N_5260,N_3341,N_2578);
nand U5261 (N_5261,N_3186,N_3647);
nand U5262 (N_5262,N_2671,N_2222);
nand U5263 (N_5263,N_3840,N_3429);
or U5264 (N_5264,N_2878,N_2062);
or U5265 (N_5265,N_3885,N_2091);
or U5266 (N_5266,N_3281,N_3055);
nor U5267 (N_5267,N_2502,N_3657);
nand U5268 (N_5268,N_2700,N_3537);
nand U5269 (N_5269,N_3493,N_2858);
and U5270 (N_5270,N_3098,N_3910);
nor U5271 (N_5271,N_2527,N_3768);
nand U5272 (N_5272,N_2218,N_2869);
nor U5273 (N_5273,N_2190,N_3402);
or U5274 (N_5274,N_3360,N_3497);
and U5275 (N_5275,N_3814,N_2035);
and U5276 (N_5276,N_3019,N_3906);
and U5277 (N_5277,N_2179,N_2615);
nand U5278 (N_5278,N_2019,N_2982);
nand U5279 (N_5279,N_2301,N_3957);
nor U5280 (N_5280,N_3745,N_2460);
nor U5281 (N_5281,N_3809,N_3869);
nand U5282 (N_5282,N_3248,N_2241);
nor U5283 (N_5283,N_2817,N_3776);
nor U5284 (N_5284,N_3101,N_2093);
or U5285 (N_5285,N_2123,N_3146);
and U5286 (N_5286,N_2970,N_3851);
nand U5287 (N_5287,N_3511,N_2593);
and U5288 (N_5288,N_3929,N_3856);
or U5289 (N_5289,N_2420,N_2485);
and U5290 (N_5290,N_2724,N_2862);
nand U5291 (N_5291,N_2753,N_2947);
nor U5292 (N_5292,N_2544,N_2777);
nand U5293 (N_5293,N_2784,N_3629);
or U5294 (N_5294,N_2883,N_2423);
or U5295 (N_5295,N_2916,N_2421);
nand U5296 (N_5296,N_2769,N_2887);
nand U5297 (N_5297,N_3114,N_2172);
nor U5298 (N_5298,N_3066,N_2556);
nand U5299 (N_5299,N_2738,N_3269);
and U5300 (N_5300,N_2259,N_3378);
nor U5301 (N_5301,N_2410,N_2037);
or U5302 (N_5302,N_3545,N_3555);
and U5303 (N_5303,N_2543,N_2768);
nand U5304 (N_5304,N_3535,N_2242);
and U5305 (N_5305,N_3696,N_2959);
nor U5306 (N_5306,N_3119,N_3724);
or U5307 (N_5307,N_3064,N_3310);
and U5308 (N_5308,N_2959,N_2830);
nand U5309 (N_5309,N_2103,N_2016);
nor U5310 (N_5310,N_2495,N_2171);
or U5311 (N_5311,N_2096,N_3569);
nor U5312 (N_5312,N_2455,N_3018);
nand U5313 (N_5313,N_2270,N_2331);
or U5314 (N_5314,N_3606,N_3450);
nand U5315 (N_5315,N_2796,N_3971);
or U5316 (N_5316,N_3369,N_2594);
and U5317 (N_5317,N_2737,N_3787);
and U5318 (N_5318,N_2722,N_3796);
nor U5319 (N_5319,N_2636,N_3796);
nor U5320 (N_5320,N_3816,N_2330);
nor U5321 (N_5321,N_3158,N_3695);
or U5322 (N_5322,N_2318,N_2279);
and U5323 (N_5323,N_3180,N_2798);
or U5324 (N_5324,N_3866,N_2732);
or U5325 (N_5325,N_3257,N_2491);
nor U5326 (N_5326,N_3071,N_3112);
and U5327 (N_5327,N_3979,N_3169);
or U5328 (N_5328,N_3802,N_2635);
nor U5329 (N_5329,N_2210,N_3936);
nor U5330 (N_5330,N_3309,N_2510);
and U5331 (N_5331,N_3011,N_3430);
nor U5332 (N_5332,N_3653,N_3201);
and U5333 (N_5333,N_3512,N_3373);
or U5334 (N_5334,N_2611,N_2767);
or U5335 (N_5335,N_3050,N_3052);
or U5336 (N_5336,N_3689,N_2631);
or U5337 (N_5337,N_2371,N_2652);
and U5338 (N_5338,N_3339,N_3415);
nand U5339 (N_5339,N_2564,N_2814);
nand U5340 (N_5340,N_2955,N_3496);
nor U5341 (N_5341,N_3261,N_2374);
nand U5342 (N_5342,N_3045,N_2376);
and U5343 (N_5343,N_2018,N_2403);
nand U5344 (N_5344,N_3001,N_2536);
or U5345 (N_5345,N_2175,N_3665);
or U5346 (N_5346,N_3606,N_3458);
nor U5347 (N_5347,N_3145,N_3199);
or U5348 (N_5348,N_2445,N_3479);
nand U5349 (N_5349,N_3093,N_3799);
and U5350 (N_5350,N_2544,N_3456);
nand U5351 (N_5351,N_2855,N_3298);
nand U5352 (N_5352,N_3375,N_2460);
or U5353 (N_5353,N_2865,N_3290);
nor U5354 (N_5354,N_2531,N_2064);
and U5355 (N_5355,N_2495,N_3229);
nor U5356 (N_5356,N_2911,N_3973);
nand U5357 (N_5357,N_3978,N_3199);
or U5358 (N_5358,N_3372,N_3602);
nand U5359 (N_5359,N_3104,N_3247);
nand U5360 (N_5360,N_2309,N_2661);
nand U5361 (N_5361,N_3493,N_3697);
or U5362 (N_5362,N_3874,N_3718);
or U5363 (N_5363,N_2363,N_2321);
and U5364 (N_5364,N_2149,N_2443);
nor U5365 (N_5365,N_3991,N_3288);
nand U5366 (N_5366,N_2387,N_3492);
nor U5367 (N_5367,N_3766,N_3443);
and U5368 (N_5368,N_2659,N_3199);
nand U5369 (N_5369,N_2892,N_2814);
nor U5370 (N_5370,N_3141,N_2353);
or U5371 (N_5371,N_3694,N_2193);
or U5372 (N_5372,N_2446,N_2131);
or U5373 (N_5373,N_2698,N_2627);
and U5374 (N_5374,N_2468,N_3449);
or U5375 (N_5375,N_3554,N_3800);
nor U5376 (N_5376,N_3344,N_3495);
nand U5377 (N_5377,N_2620,N_3192);
nor U5378 (N_5378,N_3327,N_2079);
nand U5379 (N_5379,N_3062,N_3405);
or U5380 (N_5380,N_2714,N_2775);
nand U5381 (N_5381,N_3964,N_3501);
nand U5382 (N_5382,N_2013,N_2512);
and U5383 (N_5383,N_2018,N_3263);
or U5384 (N_5384,N_2076,N_2854);
and U5385 (N_5385,N_3176,N_3765);
nand U5386 (N_5386,N_2468,N_2503);
and U5387 (N_5387,N_2768,N_2807);
nor U5388 (N_5388,N_3412,N_3641);
nor U5389 (N_5389,N_3218,N_2388);
and U5390 (N_5390,N_3375,N_3555);
nand U5391 (N_5391,N_2234,N_3304);
nand U5392 (N_5392,N_2059,N_3409);
nand U5393 (N_5393,N_3463,N_2415);
nand U5394 (N_5394,N_2042,N_3465);
nor U5395 (N_5395,N_3379,N_2327);
nand U5396 (N_5396,N_3488,N_3363);
or U5397 (N_5397,N_3431,N_3485);
nor U5398 (N_5398,N_3607,N_2177);
and U5399 (N_5399,N_3551,N_3242);
nor U5400 (N_5400,N_2276,N_3432);
nand U5401 (N_5401,N_2105,N_3392);
nor U5402 (N_5402,N_3947,N_2652);
nand U5403 (N_5403,N_2689,N_3290);
nor U5404 (N_5404,N_3718,N_3254);
and U5405 (N_5405,N_3685,N_2012);
and U5406 (N_5406,N_2050,N_3095);
nor U5407 (N_5407,N_3577,N_2793);
and U5408 (N_5408,N_2792,N_2874);
and U5409 (N_5409,N_2689,N_2235);
or U5410 (N_5410,N_3984,N_3879);
and U5411 (N_5411,N_2259,N_3565);
and U5412 (N_5412,N_2512,N_2257);
xor U5413 (N_5413,N_3109,N_3060);
nor U5414 (N_5414,N_3314,N_3117);
or U5415 (N_5415,N_3342,N_3891);
nand U5416 (N_5416,N_3218,N_2325);
nand U5417 (N_5417,N_3408,N_3061);
nor U5418 (N_5418,N_3672,N_2519);
nor U5419 (N_5419,N_3107,N_3974);
nor U5420 (N_5420,N_2821,N_2224);
or U5421 (N_5421,N_2860,N_3940);
nand U5422 (N_5422,N_2366,N_3547);
nor U5423 (N_5423,N_2842,N_2440);
and U5424 (N_5424,N_3510,N_3691);
nor U5425 (N_5425,N_3067,N_2634);
nor U5426 (N_5426,N_3889,N_3761);
nand U5427 (N_5427,N_3615,N_2588);
nor U5428 (N_5428,N_3033,N_2194);
nand U5429 (N_5429,N_2087,N_3387);
nor U5430 (N_5430,N_2743,N_3522);
nand U5431 (N_5431,N_2687,N_3895);
and U5432 (N_5432,N_3442,N_2511);
nor U5433 (N_5433,N_3475,N_2055);
nor U5434 (N_5434,N_3552,N_2771);
and U5435 (N_5435,N_3126,N_3278);
nor U5436 (N_5436,N_3958,N_2516);
nand U5437 (N_5437,N_2990,N_2041);
nor U5438 (N_5438,N_3241,N_2825);
nor U5439 (N_5439,N_3790,N_3341);
nand U5440 (N_5440,N_3222,N_2478);
or U5441 (N_5441,N_2148,N_3051);
nor U5442 (N_5442,N_2819,N_2194);
or U5443 (N_5443,N_2286,N_3103);
nor U5444 (N_5444,N_2565,N_2033);
nand U5445 (N_5445,N_3076,N_3162);
nand U5446 (N_5446,N_2566,N_3929);
or U5447 (N_5447,N_2778,N_3600);
nand U5448 (N_5448,N_3365,N_2024);
and U5449 (N_5449,N_3942,N_2486);
and U5450 (N_5450,N_3346,N_3992);
or U5451 (N_5451,N_2243,N_2257);
nor U5452 (N_5452,N_2268,N_3692);
and U5453 (N_5453,N_3412,N_3182);
nor U5454 (N_5454,N_3182,N_3856);
or U5455 (N_5455,N_2323,N_3472);
and U5456 (N_5456,N_3510,N_3284);
or U5457 (N_5457,N_2139,N_2513);
nand U5458 (N_5458,N_2397,N_3631);
nand U5459 (N_5459,N_3297,N_3143);
nor U5460 (N_5460,N_3291,N_2525);
nand U5461 (N_5461,N_2629,N_3751);
or U5462 (N_5462,N_2708,N_2704);
and U5463 (N_5463,N_3475,N_3868);
nand U5464 (N_5464,N_3912,N_2371);
and U5465 (N_5465,N_3291,N_3303);
and U5466 (N_5466,N_2065,N_2119);
nor U5467 (N_5467,N_3506,N_3269);
nor U5468 (N_5468,N_2661,N_2481);
and U5469 (N_5469,N_3083,N_2379);
nand U5470 (N_5470,N_2012,N_3256);
nor U5471 (N_5471,N_3387,N_2568);
nor U5472 (N_5472,N_2363,N_2072);
nor U5473 (N_5473,N_3820,N_2208);
and U5474 (N_5474,N_2092,N_3174);
nand U5475 (N_5475,N_3831,N_2450);
or U5476 (N_5476,N_2477,N_2671);
and U5477 (N_5477,N_2480,N_2008);
nor U5478 (N_5478,N_2530,N_3012);
or U5479 (N_5479,N_2932,N_2025);
nor U5480 (N_5480,N_3086,N_2787);
nand U5481 (N_5481,N_2929,N_2299);
nand U5482 (N_5482,N_3396,N_2564);
nor U5483 (N_5483,N_3957,N_2117);
or U5484 (N_5484,N_2792,N_2766);
or U5485 (N_5485,N_2746,N_3389);
or U5486 (N_5486,N_3808,N_3185);
nand U5487 (N_5487,N_2295,N_2820);
or U5488 (N_5488,N_2993,N_3986);
or U5489 (N_5489,N_3539,N_3898);
or U5490 (N_5490,N_2130,N_2045);
and U5491 (N_5491,N_2633,N_2498);
nand U5492 (N_5492,N_2632,N_2488);
nor U5493 (N_5493,N_2680,N_3940);
or U5494 (N_5494,N_2694,N_3255);
and U5495 (N_5495,N_3345,N_2383);
and U5496 (N_5496,N_3122,N_3700);
and U5497 (N_5497,N_3957,N_3958);
nand U5498 (N_5498,N_2538,N_3589);
nand U5499 (N_5499,N_2299,N_3996);
or U5500 (N_5500,N_3176,N_3226);
or U5501 (N_5501,N_2170,N_2981);
nand U5502 (N_5502,N_2437,N_2040);
or U5503 (N_5503,N_3180,N_2672);
or U5504 (N_5504,N_2318,N_2010);
or U5505 (N_5505,N_2871,N_3035);
nand U5506 (N_5506,N_2989,N_3085);
nand U5507 (N_5507,N_3205,N_2727);
or U5508 (N_5508,N_3372,N_2178);
or U5509 (N_5509,N_3480,N_3787);
and U5510 (N_5510,N_3864,N_2750);
and U5511 (N_5511,N_3661,N_3206);
or U5512 (N_5512,N_3904,N_3085);
and U5513 (N_5513,N_2011,N_3211);
nor U5514 (N_5514,N_2448,N_2922);
and U5515 (N_5515,N_3656,N_2805);
nor U5516 (N_5516,N_2270,N_3042);
nand U5517 (N_5517,N_2425,N_3972);
nor U5518 (N_5518,N_3069,N_2154);
and U5519 (N_5519,N_3262,N_2901);
and U5520 (N_5520,N_2969,N_2296);
and U5521 (N_5521,N_3706,N_2527);
nor U5522 (N_5522,N_3617,N_2110);
nor U5523 (N_5523,N_3897,N_2278);
nand U5524 (N_5524,N_2719,N_2509);
nor U5525 (N_5525,N_3048,N_3964);
or U5526 (N_5526,N_2537,N_3454);
nand U5527 (N_5527,N_3734,N_3709);
and U5528 (N_5528,N_3901,N_2704);
and U5529 (N_5529,N_2943,N_3122);
or U5530 (N_5530,N_2134,N_3864);
or U5531 (N_5531,N_2976,N_2995);
nand U5532 (N_5532,N_2021,N_2786);
or U5533 (N_5533,N_3497,N_3252);
and U5534 (N_5534,N_2016,N_3634);
or U5535 (N_5535,N_3301,N_2710);
or U5536 (N_5536,N_2314,N_2100);
nor U5537 (N_5537,N_2274,N_2029);
nand U5538 (N_5538,N_3237,N_3200);
and U5539 (N_5539,N_3889,N_3510);
or U5540 (N_5540,N_2989,N_2759);
nand U5541 (N_5541,N_2084,N_2648);
or U5542 (N_5542,N_2534,N_3391);
nand U5543 (N_5543,N_3783,N_3523);
nor U5544 (N_5544,N_2081,N_2895);
and U5545 (N_5545,N_3699,N_2663);
nor U5546 (N_5546,N_2613,N_3462);
or U5547 (N_5547,N_3599,N_2574);
and U5548 (N_5548,N_3367,N_2299);
or U5549 (N_5549,N_2429,N_3521);
nor U5550 (N_5550,N_2710,N_3179);
nand U5551 (N_5551,N_2687,N_2385);
or U5552 (N_5552,N_2078,N_3540);
nor U5553 (N_5553,N_2037,N_2244);
nor U5554 (N_5554,N_3551,N_2761);
nor U5555 (N_5555,N_2607,N_2997);
nand U5556 (N_5556,N_2612,N_3763);
or U5557 (N_5557,N_3496,N_3998);
or U5558 (N_5558,N_3590,N_3941);
or U5559 (N_5559,N_2516,N_3800);
nor U5560 (N_5560,N_2186,N_3837);
nor U5561 (N_5561,N_2603,N_2321);
and U5562 (N_5562,N_3999,N_3121);
or U5563 (N_5563,N_2261,N_3940);
or U5564 (N_5564,N_2219,N_2681);
nand U5565 (N_5565,N_3395,N_2861);
nand U5566 (N_5566,N_2223,N_3599);
nand U5567 (N_5567,N_3237,N_3267);
nor U5568 (N_5568,N_3880,N_3008);
or U5569 (N_5569,N_3298,N_2505);
xnor U5570 (N_5570,N_3817,N_2091);
and U5571 (N_5571,N_3459,N_2015);
nor U5572 (N_5572,N_2272,N_2396);
nand U5573 (N_5573,N_2715,N_2786);
or U5574 (N_5574,N_3113,N_2476);
and U5575 (N_5575,N_2481,N_3394);
or U5576 (N_5576,N_3891,N_3652);
and U5577 (N_5577,N_2907,N_2753);
and U5578 (N_5578,N_3662,N_3301);
nor U5579 (N_5579,N_2000,N_3797);
and U5580 (N_5580,N_3289,N_2595);
and U5581 (N_5581,N_3921,N_2360);
or U5582 (N_5582,N_2205,N_3521);
nor U5583 (N_5583,N_2635,N_2806);
and U5584 (N_5584,N_2473,N_3307);
and U5585 (N_5585,N_3673,N_3523);
nor U5586 (N_5586,N_3472,N_2810);
or U5587 (N_5587,N_2656,N_3978);
and U5588 (N_5588,N_3178,N_3510);
nor U5589 (N_5589,N_3877,N_3053);
nand U5590 (N_5590,N_3308,N_2605);
and U5591 (N_5591,N_2203,N_3692);
nand U5592 (N_5592,N_2671,N_2145);
and U5593 (N_5593,N_2108,N_3109);
or U5594 (N_5594,N_3306,N_3173);
nand U5595 (N_5595,N_3459,N_2879);
or U5596 (N_5596,N_2257,N_3600);
or U5597 (N_5597,N_2592,N_3932);
and U5598 (N_5598,N_3673,N_3531);
nor U5599 (N_5599,N_2536,N_2738);
or U5600 (N_5600,N_3750,N_2983);
or U5601 (N_5601,N_2682,N_3755);
or U5602 (N_5602,N_3820,N_2296);
nor U5603 (N_5603,N_2941,N_3015);
nand U5604 (N_5604,N_3869,N_2066);
nor U5605 (N_5605,N_3902,N_2275);
or U5606 (N_5606,N_2274,N_3110);
nor U5607 (N_5607,N_2397,N_2575);
nand U5608 (N_5608,N_3506,N_3397);
nand U5609 (N_5609,N_3286,N_3593);
nand U5610 (N_5610,N_3650,N_2310);
nand U5611 (N_5611,N_3076,N_2315);
nand U5612 (N_5612,N_2519,N_2916);
nor U5613 (N_5613,N_2199,N_3136);
and U5614 (N_5614,N_2944,N_2506);
or U5615 (N_5615,N_2565,N_2025);
nor U5616 (N_5616,N_3081,N_3902);
and U5617 (N_5617,N_2074,N_3093);
or U5618 (N_5618,N_3350,N_2430);
and U5619 (N_5619,N_2081,N_3662);
nor U5620 (N_5620,N_2598,N_3862);
nor U5621 (N_5621,N_2844,N_2795);
nand U5622 (N_5622,N_3441,N_3396);
and U5623 (N_5623,N_2629,N_2412);
or U5624 (N_5624,N_2790,N_2759);
and U5625 (N_5625,N_3332,N_2504);
nor U5626 (N_5626,N_3831,N_2214);
or U5627 (N_5627,N_2723,N_2821);
or U5628 (N_5628,N_3500,N_3551);
nor U5629 (N_5629,N_3280,N_2965);
nand U5630 (N_5630,N_2642,N_2804);
nand U5631 (N_5631,N_3845,N_3932);
and U5632 (N_5632,N_3636,N_3901);
nor U5633 (N_5633,N_3919,N_3438);
nor U5634 (N_5634,N_3959,N_3696);
or U5635 (N_5635,N_3341,N_2341);
and U5636 (N_5636,N_3414,N_3999);
and U5637 (N_5637,N_3504,N_3149);
nor U5638 (N_5638,N_3870,N_3547);
or U5639 (N_5639,N_2991,N_2571);
nand U5640 (N_5640,N_3603,N_3642);
and U5641 (N_5641,N_2618,N_3676);
nand U5642 (N_5642,N_2840,N_2896);
nor U5643 (N_5643,N_3919,N_3181);
nor U5644 (N_5644,N_3729,N_3306);
and U5645 (N_5645,N_3091,N_3761);
nand U5646 (N_5646,N_2580,N_3164);
xor U5647 (N_5647,N_2161,N_3697);
nor U5648 (N_5648,N_3574,N_3793);
nand U5649 (N_5649,N_2489,N_3338);
nand U5650 (N_5650,N_2438,N_2235);
and U5651 (N_5651,N_3776,N_3539);
nor U5652 (N_5652,N_2469,N_2219);
and U5653 (N_5653,N_3257,N_3744);
nand U5654 (N_5654,N_3453,N_3937);
and U5655 (N_5655,N_2576,N_3900);
nand U5656 (N_5656,N_2705,N_3445);
nor U5657 (N_5657,N_2500,N_2466);
or U5658 (N_5658,N_3879,N_3972);
nor U5659 (N_5659,N_2257,N_2283);
and U5660 (N_5660,N_2755,N_3941);
nand U5661 (N_5661,N_3458,N_2489);
nand U5662 (N_5662,N_2089,N_2733);
nand U5663 (N_5663,N_3147,N_3210);
or U5664 (N_5664,N_2454,N_3168);
and U5665 (N_5665,N_3121,N_3146);
nor U5666 (N_5666,N_2950,N_3239);
nor U5667 (N_5667,N_2714,N_3206);
or U5668 (N_5668,N_3954,N_3545);
nand U5669 (N_5669,N_3477,N_3260);
nor U5670 (N_5670,N_3237,N_2179);
and U5671 (N_5671,N_3727,N_2954);
or U5672 (N_5672,N_3862,N_2283);
nand U5673 (N_5673,N_3176,N_2069);
nor U5674 (N_5674,N_2643,N_3920);
nor U5675 (N_5675,N_3366,N_2619);
and U5676 (N_5676,N_3662,N_3526);
and U5677 (N_5677,N_3658,N_2169);
or U5678 (N_5678,N_2566,N_3784);
xnor U5679 (N_5679,N_3802,N_2957);
or U5680 (N_5680,N_2315,N_3619);
nor U5681 (N_5681,N_3022,N_3825);
or U5682 (N_5682,N_2158,N_2457);
or U5683 (N_5683,N_2630,N_3417);
and U5684 (N_5684,N_2112,N_3194);
nand U5685 (N_5685,N_3947,N_2041);
and U5686 (N_5686,N_2626,N_3085);
or U5687 (N_5687,N_2587,N_3345);
nand U5688 (N_5688,N_3692,N_3752);
nor U5689 (N_5689,N_3392,N_2639);
nand U5690 (N_5690,N_3303,N_3422);
nor U5691 (N_5691,N_2900,N_2446);
or U5692 (N_5692,N_2209,N_2558);
or U5693 (N_5693,N_3234,N_2941);
nand U5694 (N_5694,N_2015,N_3048);
nand U5695 (N_5695,N_3760,N_3793);
nand U5696 (N_5696,N_3017,N_3537);
or U5697 (N_5697,N_2063,N_2527);
nor U5698 (N_5698,N_3051,N_3111);
and U5699 (N_5699,N_3307,N_2681);
nor U5700 (N_5700,N_3741,N_3242);
or U5701 (N_5701,N_3800,N_3597);
xor U5702 (N_5702,N_3374,N_3243);
nor U5703 (N_5703,N_3451,N_3031);
nor U5704 (N_5704,N_3093,N_3960);
nand U5705 (N_5705,N_3746,N_2957);
nor U5706 (N_5706,N_3505,N_2553);
nand U5707 (N_5707,N_3856,N_3428);
or U5708 (N_5708,N_2476,N_2385);
or U5709 (N_5709,N_3529,N_2813);
nor U5710 (N_5710,N_3451,N_3454);
nand U5711 (N_5711,N_3133,N_3916);
and U5712 (N_5712,N_2548,N_3588);
nand U5713 (N_5713,N_2385,N_3853);
or U5714 (N_5714,N_3118,N_3570);
and U5715 (N_5715,N_3394,N_2720);
and U5716 (N_5716,N_2543,N_2185);
nor U5717 (N_5717,N_2802,N_3179);
and U5718 (N_5718,N_2856,N_3249);
nor U5719 (N_5719,N_2542,N_2973);
nor U5720 (N_5720,N_3578,N_2643);
nor U5721 (N_5721,N_2789,N_3612);
nor U5722 (N_5722,N_2790,N_2738);
nor U5723 (N_5723,N_3536,N_2419);
or U5724 (N_5724,N_2245,N_2722);
nand U5725 (N_5725,N_2527,N_3952);
nand U5726 (N_5726,N_2856,N_3567);
and U5727 (N_5727,N_2170,N_3727);
and U5728 (N_5728,N_3429,N_2113);
and U5729 (N_5729,N_2339,N_2160);
or U5730 (N_5730,N_2844,N_3832);
nand U5731 (N_5731,N_3243,N_3267);
nand U5732 (N_5732,N_2893,N_2748);
nor U5733 (N_5733,N_3913,N_3184);
nor U5734 (N_5734,N_2096,N_2663);
or U5735 (N_5735,N_3196,N_3987);
or U5736 (N_5736,N_2238,N_3424);
and U5737 (N_5737,N_3406,N_3213);
nand U5738 (N_5738,N_3903,N_3105);
nor U5739 (N_5739,N_3402,N_3376);
nor U5740 (N_5740,N_2179,N_3596);
and U5741 (N_5741,N_2672,N_3702);
nand U5742 (N_5742,N_3863,N_3572);
nor U5743 (N_5743,N_3887,N_2208);
nand U5744 (N_5744,N_3391,N_2319);
and U5745 (N_5745,N_2917,N_3486);
nand U5746 (N_5746,N_3246,N_2100);
nand U5747 (N_5747,N_3544,N_2771);
and U5748 (N_5748,N_2811,N_3658);
or U5749 (N_5749,N_3947,N_3528);
nand U5750 (N_5750,N_2155,N_2790);
or U5751 (N_5751,N_3548,N_3373);
and U5752 (N_5752,N_3763,N_3357);
nand U5753 (N_5753,N_3037,N_2965);
nor U5754 (N_5754,N_3788,N_2394);
nor U5755 (N_5755,N_2562,N_3644);
nand U5756 (N_5756,N_3407,N_2847);
or U5757 (N_5757,N_3096,N_3017);
and U5758 (N_5758,N_2129,N_3189);
or U5759 (N_5759,N_3853,N_2406);
nor U5760 (N_5760,N_3619,N_2958);
or U5761 (N_5761,N_2064,N_3019);
nor U5762 (N_5762,N_2112,N_3770);
and U5763 (N_5763,N_2336,N_2516);
nor U5764 (N_5764,N_2891,N_2595);
nor U5765 (N_5765,N_2317,N_3597);
nand U5766 (N_5766,N_3264,N_3942);
nand U5767 (N_5767,N_2716,N_3899);
nand U5768 (N_5768,N_2399,N_3695);
nand U5769 (N_5769,N_3871,N_3951);
or U5770 (N_5770,N_2056,N_2278);
nor U5771 (N_5771,N_2189,N_2553);
nor U5772 (N_5772,N_2003,N_2161);
nor U5773 (N_5773,N_3882,N_3810);
nor U5774 (N_5774,N_2415,N_3815);
nor U5775 (N_5775,N_2160,N_3100);
nand U5776 (N_5776,N_2130,N_2627);
and U5777 (N_5777,N_2672,N_3044);
and U5778 (N_5778,N_2391,N_3201);
nand U5779 (N_5779,N_2954,N_2035);
and U5780 (N_5780,N_2883,N_3877);
nand U5781 (N_5781,N_3272,N_2549);
and U5782 (N_5782,N_2636,N_3470);
and U5783 (N_5783,N_2330,N_3539);
nor U5784 (N_5784,N_2222,N_3099);
nor U5785 (N_5785,N_3805,N_3190);
and U5786 (N_5786,N_2983,N_2975);
nand U5787 (N_5787,N_3980,N_2833);
or U5788 (N_5788,N_3663,N_2872);
and U5789 (N_5789,N_3749,N_3574);
or U5790 (N_5790,N_3720,N_3967);
nor U5791 (N_5791,N_2474,N_2273);
nor U5792 (N_5792,N_2995,N_3686);
nor U5793 (N_5793,N_3085,N_3416);
nand U5794 (N_5794,N_3857,N_3444);
nor U5795 (N_5795,N_2999,N_2417);
nand U5796 (N_5796,N_2361,N_3867);
or U5797 (N_5797,N_2873,N_3163);
or U5798 (N_5798,N_3440,N_3015);
nand U5799 (N_5799,N_3442,N_2904);
nor U5800 (N_5800,N_3634,N_2039);
nor U5801 (N_5801,N_2628,N_2330);
nor U5802 (N_5802,N_2972,N_3534);
or U5803 (N_5803,N_3955,N_2755);
nand U5804 (N_5804,N_2890,N_3748);
nor U5805 (N_5805,N_3622,N_2070);
and U5806 (N_5806,N_3904,N_3106);
nand U5807 (N_5807,N_2726,N_2731);
and U5808 (N_5808,N_3594,N_3778);
and U5809 (N_5809,N_3674,N_2981);
or U5810 (N_5810,N_2577,N_3447);
or U5811 (N_5811,N_3769,N_3807);
nand U5812 (N_5812,N_3838,N_2305);
and U5813 (N_5813,N_3802,N_3940);
and U5814 (N_5814,N_2221,N_2832);
nor U5815 (N_5815,N_3488,N_2252);
nand U5816 (N_5816,N_3346,N_3258);
nor U5817 (N_5817,N_2003,N_3473);
nand U5818 (N_5818,N_2009,N_2045);
xor U5819 (N_5819,N_2760,N_2477);
nor U5820 (N_5820,N_2780,N_2313);
or U5821 (N_5821,N_2881,N_2646);
nor U5822 (N_5822,N_2051,N_3254);
and U5823 (N_5823,N_2475,N_3359);
nand U5824 (N_5824,N_2784,N_3848);
and U5825 (N_5825,N_3178,N_2776);
or U5826 (N_5826,N_3813,N_3382);
and U5827 (N_5827,N_3849,N_2886);
or U5828 (N_5828,N_3525,N_2430);
nor U5829 (N_5829,N_3270,N_2688);
nand U5830 (N_5830,N_2563,N_2712);
and U5831 (N_5831,N_2756,N_2767);
nor U5832 (N_5832,N_3302,N_2436);
or U5833 (N_5833,N_3629,N_2483);
or U5834 (N_5834,N_2793,N_3769);
and U5835 (N_5835,N_2998,N_3469);
nor U5836 (N_5836,N_3463,N_3066);
nor U5837 (N_5837,N_3465,N_3405);
nand U5838 (N_5838,N_3075,N_3825);
or U5839 (N_5839,N_3864,N_3033);
and U5840 (N_5840,N_3378,N_2713);
nand U5841 (N_5841,N_3322,N_2056);
and U5842 (N_5842,N_3680,N_3022);
nor U5843 (N_5843,N_2203,N_3074);
or U5844 (N_5844,N_2077,N_2337);
nor U5845 (N_5845,N_3000,N_3704);
or U5846 (N_5846,N_2233,N_3704);
and U5847 (N_5847,N_2686,N_2281);
nand U5848 (N_5848,N_3245,N_2558);
nor U5849 (N_5849,N_3749,N_3522);
and U5850 (N_5850,N_2619,N_3248);
or U5851 (N_5851,N_2492,N_2399);
or U5852 (N_5852,N_2636,N_2572);
nor U5853 (N_5853,N_3872,N_3606);
or U5854 (N_5854,N_3417,N_2548);
nand U5855 (N_5855,N_2428,N_2929);
nand U5856 (N_5856,N_3423,N_2372);
nand U5857 (N_5857,N_3906,N_2137);
nand U5858 (N_5858,N_3978,N_2061);
nor U5859 (N_5859,N_3861,N_3092);
and U5860 (N_5860,N_3921,N_2015);
and U5861 (N_5861,N_3041,N_3912);
and U5862 (N_5862,N_2787,N_3990);
nand U5863 (N_5863,N_2707,N_3768);
nand U5864 (N_5864,N_3258,N_3962);
or U5865 (N_5865,N_3060,N_2448);
or U5866 (N_5866,N_3100,N_2910);
and U5867 (N_5867,N_3591,N_3844);
nand U5868 (N_5868,N_2662,N_2881);
or U5869 (N_5869,N_3168,N_3833);
and U5870 (N_5870,N_2238,N_2191);
or U5871 (N_5871,N_3133,N_3469);
and U5872 (N_5872,N_3054,N_3920);
and U5873 (N_5873,N_2134,N_2043);
and U5874 (N_5874,N_2103,N_3948);
nor U5875 (N_5875,N_3936,N_3135);
nor U5876 (N_5876,N_2336,N_3763);
nor U5877 (N_5877,N_3916,N_2294);
nor U5878 (N_5878,N_3362,N_2177);
nand U5879 (N_5879,N_2420,N_2750);
and U5880 (N_5880,N_3819,N_3064);
nor U5881 (N_5881,N_2801,N_2179);
or U5882 (N_5882,N_2645,N_3604);
nor U5883 (N_5883,N_2389,N_2272);
nor U5884 (N_5884,N_2397,N_3014);
nor U5885 (N_5885,N_2739,N_2161);
and U5886 (N_5886,N_2987,N_2550);
and U5887 (N_5887,N_3598,N_2447);
or U5888 (N_5888,N_2062,N_3940);
nand U5889 (N_5889,N_3364,N_3269);
or U5890 (N_5890,N_3567,N_2035);
and U5891 (N_5891,N_2384,N_2873);
and U5892 (N_5892,N_2763,N_3090);
and U5893 (N_5893,N_3962,N_3357);
or U5894 (N_5894,N_3891,N_2192);
or U5895 (N_5895,N_3675,N_2782);
nor U5896 (N_5896,N_3978,N_2002);
or U5897 (N_5897,N_3035,N_2035);
and U5898 (N_5898,N_2554,N_2798);
nor U5899 (N_5899,N_2499,N_3904);
nor U5900 (N_5900,N_3907,N_2500);
and U5901 (N_5901,N_3744,N_3729);
and U5902 (N_5902,N_2340,N_2793);
nand U5903 (N_5903,N_2219,N_2969);
nand U5904 (N_5904,N_2502,N_3299);
or U5905 (N_5905,N_2142,N_3654);
or U5906 (N_5906,N_3653,N_2449);
nor U5907 (N_5907,N_3866,N_2120);
nor U5908 (N_5908,N_3584,N_3972);
and U5909 (N_5909,N_3235,N_2222);
or U5910 (N_5910,N_3246,N_2288);
or U5911 (N_5911,N_2284,N_3164);
nand U5912 (N_5912,N_2097,N_3750);
or U5913 (N_5913,N_3606,N_3221);
or U5914 (N_5914,N_2627,N_2725);
nand U5915 (N_5915,N_2353,N_3244);
nor U5916 (N_5916,N_3392,N_3405);
and U5917 (N_5917,N_3420,N_2183);
and U5918 (N_5918,N_2994,N_2016);
and U5919 (N_5919,N_2143,N_3517);
nor U5920 (N_5920,N_3373,N_2211);
nand U5921 (N_5921,N_3306,N_3238);
and U5922 (N_5922,N_2567,N_3620);
nor U5923 (N_5923,N_2258,N_2075);
and U5924 (N_5924,N_2272,N_3042);
or U5925 (N_5925,N_2625,N_3167);
nor U5926 (N_5926,N_2950,N_2541);
nor U5927 (N_5927,N_2214,N_3502);
nor U5928 (N_5928,N_2962,N_3798);
and U5929 (N_5929,N_2243,N_2732);
and U5930 (N_5930,N_2717,N_2047);
or U5931 (N_5931,N_2421,N_2720);
and U5932 (N_5932,N_3581,N_2385);
nand U5933 (N_5933,N_3966,N_2005);
and U5934 (N_5934,N_2161,N_3912);
xnor U5935 (N_5935,N_3437,N_3304);
or U5936 (N_5936,N_3527,N_2244);
nor U5937 (N_5937,N_3280,N_2422);
and U5938 (N_5938,N_3713,N_3034);
or U5939 (N_5939,N_3231,N_3266);
or U5940 (N_5940,N_3639,N_3763);
and U5941 (N_5941,N_2417,N_2566);
and U5942 (N_5942,N_3836,N_3333);
nor U5943 (N_5943,N_3808,N_3756);
nor U5944 (N_5944,N_3658,N_2221);
nand U5945 (N_5945,N_3119,N_3107);
nand U5946 (N_5946,N_2815,N_3499);
nand U5947 (N_5947,N_3245,N_2154);
and U5948 (N_5948,N_2514,N_2269);
and U5949 (N_5949,N_3772,N_2458);
nor U5950 (N_5950,N_3035,N_3620);
and U5951 (N_5951,N_2329,N_2601);
nand U5952 (N_5952,N_2580,N_3508);
nand U5953 (N_5953,N_2092,N_3602);
nor U5954 (N_5954,N_2320,N_2723);
nor U5955 (N_5955,N_3647,N_2559);
or U5956 (N_5956,N_3737,N_3927);
nor U5957 (N_5957,N_2190,N_2059);
nand U5958 (N_5958,N_2426,N_3140);
nor U5959 (N_5959,N_3708,N_2032);
nor U5960 (N_5960,N_3165,N_2464);
nor U5961 (N_5961,N_3007,N_2867);
nand U5962 (N_5962,N_2904,N_3873);
and U5963 (N_5963,N_2645,N_2447);
or U5964 (N_5964,N_3730,N_2721);
or U5965 (N_5965,N_2455,N_3301);
nor U5966 (N_5966,N_3043,N_3161);
or U5967 (N_5967,N_2620,N_2185);
nor U5968 (N_5968,N_3232,N_3399);
and U5969 (N_5969,N_3331,N_2794);
and U5970 (N_5970,N_2520,N_3326);
and U5971 (N_5971,N_2419,N_2599);
nand U5972 (N_5972,N_2723,N_2013);
nand U5973 (N_5973,N_2830,N_3102);
and U5974 (N_5974,N_2445,N_3965);
or U5975 (N_5975,N_2347,N_2905);
nand U5976 (N_5976,N_2416,N_3809);
nor U5977 (N_5977,N_3785,N_2075);
nand U5978 (N_5978,N_3513,N_3090);
and U5979 (N_5979,N_2414,N_2308);
nor U5980 (N_5980,N_3772,N_2913);
and U5981 (N_5981,N_2673,N_3115);
and U5982 (N_5982,N_2230,N_2918);
and U5983 (N_5983,N_2302,N_2762);
or U5984 (N_5984,N_2638,N_3499);
and U5985 (N_5985,N_2670,N_2070);
nand U5986 (N_5986,N_2905,N_2423);
nor U5987 (N_5987,N_2148,N_2105);
or U5988 (N_5988,N_2386,N_2380);
or U5989 (N_5989,N_3823,N_3351);
and U5990 (N_5990,N_2223,N_2375);
nor U5991 (N_5991,N_2111,N_3948);
nor U5992 (N_5992,N_3577,N_2601);
xnor U5993 (N_5993,N_2522,N_3633);
and U5994 (N_5994,N_2829,N_2058);
and U5995 (N_5995,N_2953,N_2484);
or U5996 (N_5996,N_2506,N_2482);
and U5997 (N_5997,N_2631,N_2802);
and U5998 (N_5998,N_3895,N_3049);
nand U5999 (N_5999,N_2109,N_2727);
nand U6000 (N_6000,N_5719,N_4853);
nor U6001 (N_6001,N_5419,N_5332);
nor U6002 (N_6002,N_5802,N_4918);
nand U6003 (N_6003,N_5508,N_4609);
nor U6004 (N_6004,N_4723,N_4139);
nor U6005 (N_6005,N_5650,N_5918);
nor U6006 (N_6006,N_4223,N_4649);
nand U6007 (N_6007,N_4610,N_5180);
or U6008 (N_6008,N_5268,N_4745);
nor U6009 (N_6009,N_4237,N_4180);
or U6010 (N_6010,N_5424,N_4002);
or U6011 (N_6011,N_5727,N_5235);
nand U6012 (N_6012,N_5111,N_4955);
or U6013 (N_6013,N_5984,N_5136);
nor U6014 (N_6014,N_5524,N_4282);
xnor U6015 (N_6015,N_4784,N_5598);
and U6016 (N_6016,N_5916,N_4840);
nor U6017 (N_6017,N_4488,N_4615);
nor U6018 (N_6018,N_5676,N_5870);
and U6019 (N_6019,N_5474,N_4622);
nor U6020 (N_6020,N_5611,N_4938);
nor U6021 (N_6021,N_5317,N_5912);
and U6022 (N_6022,N_5612,N_5570);
nand U6023 (N_6023,N_5402,N_5485);
or U6024 (N_6024,N_4041,N_5737);
nor U6025 (N_6025,N_5473,N_4716);
or U6026 (N_6026,N_4545,N_4017);
or U6027 (N_6027,N_4508,N_5834);
nor U6028 (N_6028,N_5023,N_4846);
and U6029 (N_6029,N_5278,N_5955);
or U6030 (N_6030,N_4075,N_5569);
or U6031 (N_6031,N_5441,N_4318);
or U6032 (N_6032,N_5795,N_4176);
nor U6033 (N_6033,N_5519,N_5693);
or U6034 (N_6034,N_5456,N_4015);
or U6035 (N_6035,N_5208,N_4514);
or U6036 (N_6036,N_4877,N_5203);
nor U6037 (N_6037,N_5454,N_5100);
nand U6038 (N_6038,N_5705,N_4817);
nand U6039 (N_6039,N_4192,N_5828);
or U6040 (N_6040,N_4149,N_5274);
or U6041 (N_6041,N_5428,N_5156);
and U6042 (N_6042,N_5254,N_5489);
nor U6043 (N_6043,N_5507,N_4516);
nand U6044 (N_6044,N_5286,N_5889);
or U6045 (N_6045,N_5165,N_4263);
or U6046 (N_6046,N_4295,N_4327);
nor U6047 (N_6047,N_5991,N_5938);
nor U6048 (N_6048,N_5315,N_5123);
or U6049 (N_6049,N_5252,N_5401);
or U6050 (N_6050,N_4195,N_5781);
nor U6051 (N_6051,N_4573,N_5357);
nor U6052 (N_6052,N_5121,N_5723);
nor U6053 (N_6053,N_5396,N_5506);
nor U6054 (N_6054,N_4645,N_4110);
and U6055 (N_6055,N_5706,N_5417);
and U6056 (N_6056,N_5182,N_4504);
nand U6057 (N_6057,N_4602,N_5904);
or U6058 (N_6058,N_4688,N_5854);
nor U6059 (N_6059,N_4733,N_4048);
or U6060 (N_6060,N_5794,N_4813);
nor U6061 (N_6061,N_5391,N_5599);
and U6062 (N_6062,N_5627,N_4071);
and U6063 (N_6063,N_4505,N_4147);
or U6064 (N_6064,N_4683,N_5347);
or U6065 (N_6065,N_5899,N_4381);
nand U6066 (N_6066,N_5162,N_5699);
nand U6067 (N_6067,N_4168,N_4495);
or U6068 (N_6068,N_4666,N_4397);
nand U6069 (N_6069,N_5536,N_4083);
nor U6070 (N_6070,N_4445,N_4750);
nor U6071 (N_6071,N_5643,N_4399);
nand U6072 (N_6072,N_4629,N_5608);
nand U6073 (N_6073,N_4836,N_5697);
nor U6074 (N_6074,N_4668,N_5394);
nor U6075 (N_6075,N_5616,N_4103);
and U6076 (N_6076,N_5792,N_5059);
nor U6077 (N_6077,N_5537,N_4624);
or U6078 (N_6078,N_5558,N_4739);
or U6079 (N_6079,N_5092,N_4931);
or U6080 (N_6080,N_5110,N_5079);
nand U6081 (N_6081,N_4059,N_4014);
nor U6082 (N_6082,N_4358,N_5363);
or U6083 (N_6083,N_4751,N_4013);
and U6084 (N_6084,N_4845,N_4884);
nor U6085 (N_6085,N_5176,N_5886);
nor U6086 (N_6086,N_4788,N_4703);
nor U6087 (N_6087,N_5097,N_4022);
and U6088 (N_6088,N_5806,N_4670);
or U6089 (N_6089,N_5996,N_5484);
or U6090 (N_6090,N_5109,N_4419);
or U6091 (N_6091,N_5352,N_4903);
nor U6092 (N_6092,N_4216,N_5851);
and U6093 (N_6093,N_4033,N_5872);
and U6094 (N_6094,N_4979,N_5408);
nor U6095 (N_6095,N_5492,N_4264);
or U6096 (N_6096,N_4215,N_4581);
and U6097 (N_6097,N_4262,N_5166);
nand U6098 (N_6098,N_5201,N_5345);
and U6099 (N_6099,N_4672,N_5116);
nor U6100 (N_6100,N_5085,N_4679);
nand U6101 (N_6101,N_4606,N_5714);
nand U6102 (N_6102,N_4142,N_5452);
and U6103 (N_6103,N_4964,N_4309);
and U6104 (N_6104,N_5571,N_4208);
nand U6105 (N_6105,N_5768,N_4698);
and U6106 (N_6106,N_4321,N_4638);
and U6107 (N_6107,N_4541,N_5358);
and U6108 (N_6108,N_5024,N_4685);
or U6109 (N_6109,N_5873,N_4773);
xor U6110 (N_6110,N_5207,N_4589);
nor U6111 (N_6111,N_4842,N_4532);
or U6112 (N_6112,N_4651,N_5636);
and U6113 (N_6113,N_4108,N_5018);
nand U6114 (N_6114,N_5647,N_4693);
nor U6115 (N_6115,N_4772,N_4025);
nand U6116 (N_6116,N_4648,N_5135);
nand U6117 (N_6117,N_4521,N_5130);
and U6118 (N_6118,N_4061,N_5983);
and U6119 (N_6119,N_5917,N_5459);
or U6120 (N_6120,N_4667,N_4101);
and U6121 (N_6121,N_5529,N_5051);
and U6122 (N_6122,N_4409,N_4157);
and U6123 (N_6123,N_5739,N_5076);
nand U6124 (N_6124,N_4339,N_5838);
and U6125 (N_6125,N_5450,N_5583);
nor U6126 (N_6126,N_5189,N_4424);
and U6127 (N_6127,N_4114,N_5971);
nor U6128 (N_6128,N_4257,N_4565);
and U6129 (N_6129,N_4731,N_4276);
and U6130 (N_6130,N_4883,N_4961);
or U6131 (N_6131,N_4882,N_5762);
nor U6132 (N_6132,N_4383,N_5004);
or U6133 (N_6133,N_4815,N_5505);
and U6134 (N_6134,N_5497,N_4028);
nand U6135 (N_6135,N_4517,N_5354);
nor U6136 (N_6136,N_4193,N_5383);
and U6137 (N_6137,N_4133,N_5236);
nand U6138 (N_6138,N_5349,N_4362);
and U6139 (N_6139,N_4879,N_4953);
and U6140 (N_6140,N_5898,N_4039);
or U6141 (N_6141,N_5887,N_5979);
and U6142 (N_6142,N_4984,N_4600);
nand U6143 (N_6143,N_4839,N_5893);
nor U6144 (N_6144,N_4513,N_5368);
or U6145 (N_6145,N_5279,N_5057);
nor U6146 (N_6146,N_5206,N_4469);
nand U6147 (N_6147,N_4486,N_5879);
nand U6148 (N_6148,N_4368,N_4538);
or U6149 (N_6149,N_4084,N_4531);
nor U6150 (N_6150,N_5934,N_4416);
and U6151 (N_6151,N_4432,N_4669);
and U6152 (N_6152,N_5707,N_4554);
nand U6153 (N_6153,N_4909,N_4336);
nand U6154 (N_6154,N_4152,N_5037);
and U6155 (N_6155,N_5775,N_5796);
or U6156 (N_6156,N_4497,N_4639);
and U6157 (N_6157,N_4987,N_4222);
and U6158 (N_6158,N_5399,N_4914);
or U6159 (N_6159,N_4975,N_5052);
nand U6160 (N_6160,N_5393,N_5379);
or U6161 (N_6161,N_4427,N_5677);
or U6162 (N_6162,N_4352,N_4696);
or U6163 (N_6163,N_5602,N_5905);
and U6164 (N_6164,N_4981,N_4323);
or U6165 (N_6165,N_4047,N_5326);
nor U6166 (N_6166,N_4369,N_5062);
and U6167 (N_6167,N_4632,N_5324);
and U6168 (N_6168,N_5318,N_4546);
nand U6169 (N_6169,N_5193,N_4311);
nand U6170 (N_6170,N_5241,N_4198);
and U6171 (N_6171,N_5266,N_4908);
and U6172 (N_6172,N_5554,N_5303);
nand U6173 (N_6173,N_5360,N_4288);
nand U6174 (N_6174,N_4260,N_4475);
nor U6175 (N_6175,N_4125,N_5649);
nor U6176 (N_6176,N_4407,N_4332);
or U6177 (N_6177,N_4313,N_5029);
or U6178 (N_6178,N_5939,N_5852);
and U6179 (N_6179,N_4625,N_5095);
and U6180 (N_6180,N_5866,N_5048);
nand U6181 (N_6181,N_4951,N_5621);
nor U6182 (N_6182,N_4759,N_4359);
and U6183 (N_6183,N_5963,N_5703);
and U6184 (N_6184,N_4661,N_5653);
or U6185 (N_6185,N_4464,N_4361);
or U6186 (N_6186,N_4122,N_5986);
nor U6187 (N_6187,N_4206,N_4038);
and U6188 (N_6188,N_5339,N_4044);
and U6189 (N_6189,N_5483,N_4566);
nand U6190 (N_6190,N_5249,N_4138);
and U6191 (N_6191,N_4175,N_5531);
or U6192 (N_6192,N_4709,N_5751);
and U6193 (N_6193,N_5493,N_5977);
nor U6194 (N_6194,N_4869,N_4553);
or U6195 (N_6195,N_5875,N_4246);
nor U6196 (N_6196,N_5844,N_4753);
nand U6197 (N_6197,N_4034,N_5748);
or U6198 (N_6198,N_4927,N_4165);
or U6199 (N_6199,N_4824,N_5269);
nand U6200 (N_6200,N_4786,N_5259);
or U6201 (N_6201,N_5356,N_5125);
and U6202 (N_6202,N_5750,N_5058);
nand U6203 (N_6203,N_5388,N_5761);
and U6204 (N_6204,N_4895,N_5334);
nor U6205 (N_6205,N_5543,N_4776);
and U6206 (N_6206,N_4241,N_5535);
nand U6207 (N_6207,N_4894,N_5311);
or U6208 (N_6208,N_5847,N_4898);
nor U6209 (N_6209,N_4120,N_5798);
or U6210 (N_6210,N_5901,N_4076);
nor U6211 (N_6211,N_4476,N_5805);
or U6212 (N_6212,N_5897,N_5126);
nand U6213 (N_6213,N_4136,N_5829);
nor U6214 (N_6214,N_4522,N_4585);
and U6215 (N_6215,N_4983,N_5572);
nand U6216 (N_6216,N_4986,N_4460);
nand U6217 (N_6217,N_5435,N_5281);
or U6218 (N_6218,N_5831,N_5040);
or U6219 (N_6219,N_5623,N_5128);
nor U6220 (N_6220,N_5929,N_4158);
or U6221 (N_6221,N_4978,N_5528);
nor U6222 (N_6222,N_5378,N_5271);
or U6223 (N_6223,N_5858,N_4253);
nor U6224 (N_6224,N_4601,N_4082);
and U6225 (N_6225,N_5168,N_5691);
nand U6226 (N_6226,N_5782,N_5733);
or U6227 (N_6227,N_5876,N_4935);
or U6228 (N_6228,N_5370,N_4652);
nand U6229 (N_6229,N_4389,N_5477);
and U6230 (N_6230,N_5814,N_5453);
and U6231 (N_6231,N_5147,N_4112);
or U6232 (N_6232,N_5509,N_5908);
nand U6233 (N_6233,N_4375,N_5285);
or U6234 (N_6234,N_5812,N_5053);
and U6235 (N_6235,N_5803,N_5864);
nand U6236 (N_6236,N_4473,N_4963);
nor U6237 (N_6237,N_4635,N_5824);
or U6238 (N_6238,N_5752,N_5478);
nand U6239 (N_6239,N_4329,N_5362);
or U6240 (N_6240,N_4694,N_5142);
nor U6241 (N_6241,N_5465,N_4163);
nor U6242 (N_6242,N_4436,N_5436);
nor U6243 (N_6243,N_5118,N_5837);
nand U6244 (N_6244,N_4798,N_5581);
nor U6245 (N_6245,N_5250,N_5856);
or U6246 (N_6246,N_5578,N_5398);
nand U6247 (N_6247,N_5511,N_5213);
nand U6248 (N_6248,N_5019,N_5670);
or U6249 (N_6249,N_5124,N_5630);
and U6250 (N_6250,N_5496,N_5001);
and U6251 (N_6251,N_4428,N_4873);
nand U6252 (N_6252,N_4036,N_4132);
nand U6253 (N_6253,N_4921,N_4027);
or U6254 (N_6254,N_5395,N_5006);
and U6255 (N_6255,N_4293,N_5325);
nor U6256 (N_6256,N_5726,N_5439);
nand U6257 (N_6257,N_4370,N_5003);
nand U6258 (N_6258,N_5813,N_5800);
nand U6259 (N_6259,N_5718,N_5197);
and U6260 (N_6260,N_4185,N_4579);
and U6261 (N_6261,N_4200,N_4159);
nand U6262 (N_6262,N_4151,N_5686);
nand U6263 (N_6263,N_5954,N_5444);
nor U6264 (N_6264,N_4593,N_4535);
nand U6265 (N_6265,N_4063,N_4787);
and U6266 (N_6266,N_5545,N_4760);
nand U6267 (N_6267,N_4782,N_5300);
or U6268 (N_6268,N_5577,N_4220);
nand U6269 (N_6269,N_5961,N_5769);
nand U6270 (N_6270,N_5140,N_5822);
and U6271 (N_6271,N_5219,N_4333);
nand U6272 (N_6272,N_5045,N_5550);
nand U6273 (N_6273,N_5853,N_4548);
nand U6274 (N_6274,N_4173,N_4519);
nor U6275 (N_6275,N_5049,N_4586);
or U6276 (N_6276,N_4093,N_4924);
and U6277 (N_6277,N_5442,N_4385);
or U6278 (N_6278,N_4524,N_5731);
or U6279 (N_6279,N_5372,N_4660);
and U6280 (N_6280,N_5967,N_5797);
and U6281 (N_6281,N_5696,N_5468);
or U6282 (N_6282,N_5808,N_4144);
and U6283 (N_6283,N_4684,N_5947);
and U6284 (N_6284,N_5759,N_5475);
nor U6285 (N_6285,N_5171,N_4637);
or U6286 (N_6286,N_4490,N_5490);
and U6287 (N_6287,N_5425,N_4506);
nand U6288 (N_6288,N_4790,N_4785);
nand U6289 (N_6289,N_5287,N_5260);
xnor U6290 (N_6290,N_4796,N_5178);
nand U6291 (N_6291,N_5307,N_5482);
nand U6292 (N_6292,N_5629,N_5722);
xnor U6293 (N_6293,N_4450,N_5985);
xnor U6294 (N_6294,N_4008,N_4856);
and U6295 (N_6295,N_5626,N_4483);
and U6296 (N_6296,N_4492,N_4422);
nor U6297 (N_6297,N_4852,N_5212);
or U6298 (N_6298,N_4550,N_5498);
nor U6299 (N_6299,N_5253,N_5687);
and U6300 (N_6300,N_5839,N_4614);
and U6301 (N_6301,N_4973,N_5234);
nor U6302 (N_6302,N_5948,N_4991);
nand U6303 (N_6303,N_5031,N_5830);
nor U6304 (N_6304,N_5639,N_5720);
nor U6305 (N_6305,N_4674,N_5669);
nor U6306 (N_6306,N_4126,N_4265);
nor U6307 (N_6307,N_5292,N_5232);
nand U6308 (N_6308,N_5237,N_4677);
nor U6309 (N_6309,N_5290,N_4205);
nand U6310 (N_6310,N_5557,N_4518);
nand U6311 (N_6311,N_4993,N_5129);
or U6312 (N_6312,N_4347,N_5843);
nor U6313 (N_6313,N_5734,N_5749);
and U6314 (N_6314,N_4561,N_5277);
or U6315 (N_6315,N_5127,N_5426);
or U6316 (N_6316,N_4307,N_5502);
nand U6317 (N_6317,N_4653,N_5713);
or U6318 (N_6318,N_5868,N_4135);
and U6319 (N_6319,N_5273,N_4491);
nand U6320 (N_6320,N_4453,N_4418);
nand U6321 (N_6321,N_4062,N_5863);
and U6322 (N_6322,N_5527,N_4328);
nor U6323 (N_6323,N_4689,N_4079);
nor U6324 (N_6324,N_5933,N_4576);
nor U6325 (N_6325,N_4090,N_4820);
nand U6326 (N_6326,N_4229,N_4226);
nor U6327 (N_6327,N_4179,N_4727);
nand U6328 (N_6328,N_5950,N_4704);
or U6329 (N_6329,N_4421,N_5012);
nand U6330 (N_6330,N_5825,N_4687);
xnor U6331 (N_6331,N_4325,N_4899);
nand U6332 (N_6332,N_4354,N_5177);
or U6333 (N_6333,N_5291,N_4081);
nor U6334 (N_6334,N_4105,N_4254);
nor U6335 (N_6335,N_5648,N_5952);
and U6336 (N_6336,N_5298,N_5657);
or U6337 (N_6337,N_5584,N_4213);
nor U6338 (N_6338,N_4489,N_4943);
nor U6339 (N_6339,N_5910,N_4045);
nor U6340 (N_6340,N_5685,N_4634);
and U6341 (N_6341,N_5264,N_5978);
nor U6342 (N_6342,N_5728,N_5440);
nand U6343 (N_6343,N_4583,N_4074);
nor U6344 (N_6344,N_4512,N_4465);
nand U6345 (N_6345,N_5148,N_5161);
and U6346 (N_6346,N_5913,N_5862);
nor U6347 (N_6347,N_4713,N_5013);
or U6348 (N_6348,N_5596,N_4239);
and U6349 (N_6349,N_4697,N_5937);
nand U6350 (N_6350,N_5282,N_5522);
and U6351 (N_6351,N_4744,N_5245);
and U6352 (N_6352,N_4280,N_5674);
and U6353 (N_6353,N_4578,N_4503);
nand U6354 (N_6354,N_4340,N_4156);
nand U6355 (N_6355,N_5411,N_4757);
nand U6356 (N_6356,N_5087,N_4072);
and U6357 (N_6357,N_4060,N_5771);
or U6358 (N_6358,N_5267,N_5944);
and U6359 (N_6359,N_4259,N_5860);
and U6360 (N_6360,N_5380,N_4641);
or U6361 (N_6361,N_4306,N_4087);
or U6362 (N_6362,N_5054,N_5560);
and U6363 (N_6363,N_5702,N_5044);
nand U6364 (N_6364,N_4663,N_5431);
nand U6365 (N_6365,N_5688,N_4190);
or U6366 (N_6366,N_5359,N_5199);
and U6367 (N_6367,N_4722,N_5679);
or U6368 (N_6368,N_5840,N_4374);
nor U6369 (N_6369,N_5160,N_4337);
nand U6370 (N_6370,N_4429,N_5747);
nand U6371 (N_6371,N_5068,N_5516);
or U6372 (N_6372,N_5365,N_5382);
nor U6373 (N_6373,N_5772,N_4890);
and U6374 (N_6374,N_4218,N_5131);
nand U6375 (N_6375,N_5007,N_4099);
or U6376 (N_6376,N_5026,N_4848);
and U6377 (N_6377,N_4570,N_4888);
or U6378 (N_6378,N_5141,N_5500);
and U6379 (N_6379,N_5082,N_4952);
or U6380 (N_6380,N_5753,N_4113);
or U6381 (N_6381,N_4708,N_4148);
and U6382 (N_6382,N_5549,N_4803);
or U6383 (N_6383,N_4801,N_4119);
nand U6384 (N_6384,N_5151,N_5030);
and U6385 (N_6385,N_5144,N_5288);
nor U6386 (N_6386,N_5150,N_4243);
or U6387 (N_6387,N_4201,N_4838);
nor U6388 (N_6388,N_4043,N_5836);
nor U6389 (N_6389,N_5566,N_4247);
or U6390 (N_6390,N_5641,N_4974);
nand U6391 (N_6391,N_5107,N_5050);
nand U6392 (N_6392,N_5907,N_5099);
nor U6393 (N_6393,N_4720,N_5405);
nand U6394 (N_6394,N_5518,N_4092);
xnor U6395 (N_6395,N_5355,N_4472);
nand U6396 (N_6396,N_5538,N_5164);
or U6397 (N_6397,N_4699,N_4940);
nand U6398 (N_6398,N_5416,N_5962);
nand U6399 (N_6399,N_4391,N_4412);
and U6400 (N_6400,N_4402,N_4302);
or U6401 (N_6401,N_4233,N_5457);
nand U6402 (N_6402,N_5225,N_4665);
nor U6403 (N_6403,N_4050,N_5036);
or U6404 (N_6404,N_4829,N_4314);
nand U6405 (N_6405,N_5773,N_4764);
and U6406 (N_6406,N_4631,N_4242);
or U6407 (N_6407,N_4203,N_5039);
nor U6408 (N_6408,N_5544,N_5633);
nand U6409 (N_6409,N_4767,N_4559);
nor U6410 (N_6410,N_5385,N_4889);
nor U6411 (N_6411,N_5115,N_4843);
nand U6412 (N_6412,N_4988,N_4404);
and U6413 (N_6413,N_5548,N_4484);
nand U6414 (N_6414,N_4584,N_4948);
nand U6415 (N_6415,N_5846,N_5169);
nor U6416 (N_6416,N_4976,N_5038);
nand U6417 (N_6417,N_4673,N_5430);
and U6418 (N_6418,N_4171,N_5240);
nand U6419 (N_6419,N_5617,N_5390);
or U6420 (N_6420,N_4997,N_4187);
and U6421 (N_6421,N_5999,N_4249);
nor U6422 (N_6422,N_5790,N_4515);
nand U6423 (N_6423,N_4941,N_4875);
nor U6424 (N_6424,N_4662,N_5032);
nor U6425 (N_6425,N_5607,N_4982);
or U6426 (N_6426,N_5066,N_5681);
or U6427 (N_6427,N_5305,N_5888);
or U6428 (N_6428,N_4186,N_5936);
and U6429 (N_6429,N_4686,N_4556);
or U6430 (N_6430,N_5112,N_4998);
or U6431 (N_6431,N_5793,N_4807);
nor U6432 (N_6432,N_5754,N_5941);
nand U6433 (N_6433,N_5154,N_4181);
nor U6434 (N_6434,N_4442,N_5367);
and U6435 (N_6435,N_5083,N_4054);
nand U6436 (N_6436,N_4406,N_4344);
nand U6437 (N_6437,N_4134,N_5446);
or U6438 (N_6438,N_4240,N_5660);
nand U6439 (N_6439,N_4835,N_5982);
or U6440 (N_6440,N_5313,N_5559);
or U6441 (N_6441,N_4317,N_4870);
nor U6442 (N_6442,N_4740,N_4085);
and U6443 (N_6443,N_4202,N_5662);
nor U6444 (N_6444,N_5369,N_4496);
or U6445 (N_6445,N_4401,N_5479);
nor U6446 (N_6446,N_5423,N_5145);
nand U6447 (N_6447,N_5601,N_4454);
nand U6448 (N_6448,N_4819,N_5301);
and U6449 (N_6449,N_5070,N_4730);
or U6450 (N_6450,N_5224,N_5993);
nand U6451 (N_6451,N_4866,N_5086);
or U6452 (N_6452,N_5600,N_5959);
nor U6453 (N_6453,N_4452,N_4178);
nor U6454 (N_6454,N_4128,N_5920);
or U6455 (N_6455,N_5343,N_4335);
xor U6456 (N_6456,N_4066,N_5561);
or U6457 (N_6457,N_4056,N_5956);
and U6458 (N_6458,N_4070,N_4658);
and U6459 (N_6459,N_4117,N_5717);
nor U6460 (N_6460,N_5766,N_4956);
or U6461 (N_6461,N_5328,N_4906);
and U6462 (N_6462,N_5258,N_4826);
and U6463 (N_6463,N_4946,N_5221);
nor U6464 (N_6464,N_4474,N_4405);
or U6465 (N_6465,N_4905,N_4086);
and U6466 (N_6466,N_5471,N_5157);
and U6467 (N_6467,N_4960,N_5384);
nor U6468 (N_6468,N_4558,N_4771);
and U6469 (N_6469,N_5021,N_5895);
and U6470 (N_6470,N_5486,N_5783);
or U6471 (N_6471,N_4244,N_4547);
or U6472 (N_6472,N_5513,N_5780);
or U6473 (N_6473,N_5333,N_5585);
or U6474 (N_6474,N_4121,N_4737);
nand U6475 (N_6475,N_5758,N_4721);
nand U6476 (N_6476,N_5510,N_5063);
and U6477 (N_6477,N_5712,N_4590);
or U6478 (N_6478,N_5575,N_5742);
or U6479 (N_6479,N_4000,N_5521);
nand U6480 (N_6480,N_5077,N_5592);
and U6481 (N_6481,N_5034,N_4706);
or U6482 (N_6482,N_4777,N_4539);
nor U6483 (N_6483,N_5091,N_4357);
or U6484 (N_6484,N_4277,N_5882);
or U6485 (N_6485,N_5774,N_5460);
and U6486 (N_6486,N_5743,N_5849);
and U6487 (N_6487,N_4141,N_4816);
nand U6488 (N_6488,N_5715,N_5046);
or U6489 (N_6489,N_5244,N_4057);
and U6490 (N_6490,N_4734,N_4743);
nor U6491 (N_6491,N_5327,N_5418);
and U6492 (N_6492,N_5447,N_4832);
nor U6493 (N_6493,N_5943,N_4741);
nand U6494 (N_6494,N_5331,N_5562);
or U6495 (N_6495,N_5338,N_5185);
or U6496 (N_6496,N_5190,N_4732);
or U6497 (N_6497,N_4928,N_5081);
or U6498 (N_6498,N_4010,N_5906);
nand U6499 (N_6499,N_5407,N_4435);
or U6500 (N_6500,N_4718,N_5919);
xnor U6501 (N_6501,N_4269,N_4088);
nand U6502 (N_6502,N_5994,N_4860);
or U6503 (N_6503,N_5209,N_5655);
and U6504 (N_6504,N_5155,N_4289);
nor U6505 (N_6505,N_4793,N_5272);
nand U6506 (N_6506,N_5532,N_5815);
and U6507 (N_6507,N_4695,N_4236);
or U6508 (N_6508,N_4118,N_5953);
or U6509 (N_6509,N_4279,N_5845);
and U6510 (N_6510,N_5243,N_4507);
or U6511 (N_6511,N_5684,N_4562);
nor U6512 (N_6512,N_4482,N_5525);
or U6513 (N_6513,N_4457,N_5826);
and U6514 (N_6514,N_5586,N_4040);
nand U6515 (N_6515,N_4380,N_5312);
nand U6516 (N_6516,N_4885,N_4290);
or U6517 (N_6517,N_5179,N_5429);
or U6518 (N_6518,N_5414,N_4217);
and U6519 (N_6519,N_4612,N_4587);
xor U6520 (N_6520,N_4305,N_5659);
nand U6521 (N_6521,N_5512,N_4864);
or U6522 (N_6522,N_4922,N_4471);
nor U6523 (N_6523,N_4766,N_4598);
and U6524 (N_6524,N_5553,N_4011);
nand U6525 (N_6525,N_4752,N_5069);
nand U6526 (N_6526,N_4534,N_5694);
nand U6527 (N_6527,N_5476,N_4627);
or U6528 (N_6528,N_4725,N_5448);
nor U6529 (N_6529,N_5590,N_4341);
nor U6530 (N_6530,N_4502,N_5078);
xor U6531 (N_6531,N_4789,N_5187);
nand U6532 (N_6532,N_4447,N_5381);
nand U6533 (N_6533,N_4455,N_4959);
or U6534 (N_6534,N_5198,N_4904);
and U6535 (N_6535,N_4705,N_4129);
or U6536 (N_6536,N_5223,N_5567);
nor U6537 (N_6537,N_5646,N_4746);
and U6538 (N_6538,N_5074,N_5494);
nor U6539 (N_6539,N_5613,N_4274);
nor U6540 (N_6540,N_4901,N_4537);
nor U6541 (N_6541,N_4913,N_4387);
or U6542 (N_6542,N_5113,N_5818);
nand U6543 (N_6543,N_5481,N_4735);
and U6544 (N_6544,N_4494,N_5551);
and U6545 (N_6545,N_5064,N_4738);
nand U6546 (N_6546,N_5997,N_5745);
nand U6547 (N_6547,N_4330,N_5923);
and U6548 (N_6548,N_5700,N_5033);
nor U6549 (N_6549,N_4026,N_5819);
nand U6550 (N_6550,N_4462,N_4911);
or U6551 (N_6551,N_4150,N_5787);
and U6552 (N_6552,N_5624,N_4643);
xor U6553 (N_6553,N_4392,N_4939);
nand U6554 (N_6554,N_4499,N_5309);
nand U6555 (N_6555,N_4018,N_4795);
nor U6556 (N_6556,N_5547,N_4154);
nand U6557 (N_6557,N_5472,N_5132);
nor U6558 (N_6558,N_4792,N_5415);
nor U6559 (N_6559,N_5297,N_5785);
nor U6560 (N_6560,N_4287,N_5009);
nand U6561 (N_6561,N_4865,N_4234);
and U6562 (N_6562,N_4255,N_4153);
nand U6563 (N_6563,N_5823,N_4871);
nor U6564 (N_6564,N_4366,N_5911);
nand U6565 (N_6565,N_4726,N_4468);
or U6566 (N_6566,N_5642,N_5654);
nor U6567 (N_6567,N_4378,N_4571);
nand U6568 (N_6568,N_4710,N_5330);
nor U6569 (N_6569,N_4999,N_5088);
nor U6570 (N_6570,N_4207,N_5098);
and U6571 (N_6571,N_5564,N_5930);
nand U6572 (N_6572,N_5990,N_4613);
nand U6573 (N_6573,N_5361,N_4529);
nor U6574 (N_6574,N_4834,N_5143);
nor U6575 (N_6575,N_5663,N_5973);
nor U6576 (N_6576,N_4137,N_4647);
nand U6577 (N_6577,N_4676,N_4568);
nand U6578 (N_6578,N_5816,N_5914);
nor U6579 (N_6579,N_4467,N_5134);
or U6580 (N_6580,N_5503,N_4212);
nor U6581 (N_6581,N_4046,N_4299);
nor U6582 (N_6582,N_4408,N_4292);
nand U6583 (N_6583,N_5348,N_5931);
or U6584 (N_6584,N_5744,N_5975);
and U6585 (N_6585,N_4778,N_5094);
and U6586 (N_6586,N_4620,N_4949);
nor U6587 (N_6587,N_4009,N_4007);
nand U6588 (N_6588,N_5364,N_4273);
nor U6589 (N_6589,N_5885,N_5877);
or U6590 (N_6590,N_5117,N_4379);
or U6591 (N_6591,N_4214,N_5579);
nand U6592 (N_6592,N_4858,N_5022);
nor U6593 (N_6593,N_4481,N_5202);
nand U6594 (N_6594,N_4107,N_5989);
or U6595 (N_6595,N_5108,N_5196);
or U6596 (N_6596,N_4990,N_4925);
nor U6597 (N_6597,N_4278,N_5072);
or U6598 (N_6598,N_5765,N_4227);
nor U6599 (N_6599,N_4692,N_5344);
xor U6600 (N_6600,N_5283,N_4671);
or U6601 (N_6601,N_4847,N_4448);
nand U6602 (N_6602,N_5192,N_5632);
nand U6603 (N_6603,N_4967,N_4320);
or U6604 (N_6604,N_5329,N_5133);
and U6605 (N_6605,N_5615,N_4881);
or U6606 (N_6606,N_4441,N_5410);
or U6607 (N_6607,N_5645,N_5932);
nor U6608 (N_6608,N_5928,N_4920);
nor U6609 (N_6609,N_5488,N_4487);
nand U6610 (N_6610,N_5060,N_4294);
nor U6611 (N_6611,N_5409,N_4131);
nor U6612 (N_6612,N_5119,N_4825);
or U6613 (N_6613,N_4837,N_4526);
and U6614 (N_6614,N_4285,N_5041);
or U6615 (N_6615,N_4035,N_5306);
nand U6616 (N_6616,N_4823,N_4929);
or U6617 (N_6617,N_4224,N_4855);
nor U6618 (N_6618,N_5695,N_4607);
and U6619 (N_6619,N_4304,N_4162);
and U6620 (N_6620,N_4619,N_4880);
or U6621 (N_6621,N_4444,N_5071);
and U6622 (N_6622,N_4891,N_4711);
and U6623 (N_6623,N_5261,N_5859);
or U6624 (N_6624,N_4989,N_4794);
and U6625 (N_6625,N_5981,N_4560);
or U6626 (N_6626,N_4310,N_4995);
and U6627 (N_6627,N_5170,N_4985);
nand U6628 (N_6628,N_4768,N_5433);
and U6629 (N_6629,N_4962,N_5296);
nand U6630 (N_6630,N_4478,N_4650);
and U6631 (N_6631,N_4319,N_5588);
nor U6632 (N_6632,N_5976,N_4065);
nand U6633 (N_6633,N_4251,N_4360);
and U6634 (N_6634,N_4400,N_5316);
or U6635 (N_6635,N_4248,N_4595);
nor U6636 (N_6636,N_5682,N_4331);
nand U6637 (N_6637,N_4828,N_5709);
and U6638 (N_6638,N_4701,N_5779);
and U6639 (N_6639,N_5970,N_5740);
nand U6640 (N_6640,N_5958,N_5096);
and U6641 (N_6641,N_4833,N_5622);
nor U6642 (N_6642,N_5184,N_5738);
nor U6643 (N_6643,N_4230,N_4211);
and U6644 (N_6644,N_4197,N_5807);
nand U6645 (N_6645,N_4349,N_4396);
or U6646 (N_6646,N_4225,N_5960);
and U6647 (N_6647,N_4994,N_5397);
or U6648 (N_6648,N_4765,N_4183);
and U6649 (N_6649,N_5319,N_5992);
and U6650 (N_6650,N_5445,N_5055);
or U6651 (N_6651,N_5820,N_4433);
and U6652 (N_6652,N_5421,N_4199);
and U6653 (N_6653,N_4382,N_4417);
nand U6654 (N_6654,N_4267,N_4012);
nand U6655 (N_6655,N_4996,N_4947);
or U6656 (N_6656,N_4365,N_5861);
nor U6657 (N_6657,N_5891,N_5809);
nand U6658 (N_6658,N_5248,N_4896);
and U6659 (N_6659,N_4461,N_5591);
and U6660 (N_6660,N_4783,N_4897);
nor U6661 (N_6661,N_4501,N_5195);
and U6662 (N_6662,N_4682,N_4851);
or U6663 (N_6663,N_4567,N_4930);
and U6664 (N_6664,N_4655,N_4659);
or U6665 (N_6665,N_4563,N_5665);
and U6666 (N_6666,N_4749,N_5275);
and U6667 (N_6667,N_4523,N_5346);
nor U6668 (N_6668,N_5620,N_5320);
and U6669 (N_6669,N_4715,N_4572);
nand U6670 (N_6670,N_4603,N_5434);
nand U6671 (N_6671,N_5651,N_4334);
nand U6672 (N_6672,N_5881,N_5946);
and U6673 (N_6673,N_4169,N_5799);
nor U6674 (N_6674,N_4042,N_5289);
nor U6675 (N_6675,N_5741,N_5231);
or U6676 (N_6676,N_4530,N_4091);
nor U6677 (N_6677,N_5464,N_5942);
nor U6678 (N_6678,N_5949,N_5350);
and U6679 (N_6679,N_5940,N_4542);
or U6680 (N_6680,N_4067,N_5342);
and U6681 (N_6681,N_4123,N_5084);
nand U6682 (N_6682,N_4324,N_4937);
and U6683 (N_6683,N_4912,N_5015);
nand U6684 (N_6684,N_5101,N_5555);
nand U6685 (N_6685,N_4810,N_5903);
and U6686 (N_6686,N_4477,N_5167);
nor U6687 (N_6687,N_5210,N_5593);
nor U6688 (N_6688,N_4006,N_5480);
and U6689 (N_6689,N_4775,N_4616);
nand U6690 (N_6690,N_5972,N_4170);
nand U6691 (N_6691,N_4440,N_5680);
nor U6692 (N_6692,N_4954,N_4143);
nand U6693 (N_6693,N_4238,N_5466);
and U6694 (N_6694,N_4591,N_5073);
and U6695 (N_6695,N_5336,N_5438);
nand U6696 (N_6696,N_5106,N_5067);
nand U6697 (N_6697,N_5610,N_5957);
and U6698 (N_6698,N_5220,N_5314);
and U6699 (N_6699,N_4892,N_5103);
nor U6700 (N_6700,N_5546,N_4608);
or U6701 (N_6701,N_5413,N_4934);
nand U6702 (N_6702,N_5776,N_5238);
and U6703 (N_6703,N_5294,N_5595);
nor U6704 (N_6704,N_5463,N_5188);
xnor U6705 (N_6705,N_4761,N_5915);
nor U6706 (N_6706,N_4210,N_5308);
nand U6707 (N_6707,N_5848,N_5909);
nand U6708 (N_6708,N_5389,N_4822);
or U6709 (N_6709,N_4664,N_5756);
nor U6710 (N_6710,N_5159,N_4104);
or U6711 (N_6711,N_5878,N_5582);
or U6712 (N_6712,N_5689,N_4970);
nand U6713 (N_6713,N_5400,N_5386);
or U6714 (N_6714,N_4511,N_5678);
and U6715 (N_6715,N_5922,N_4256);
or U6716 (N_6716,N_4830,N_5215);
nand U6717 (N_6717,N_4130,N_4814);
and U6718 (N_6718,N_5974,N_4806);
nand U6719 (N_6719,N_4301,N_4353);
and U6720 (N_6720,N_4411,N_4748);
and U6721 (N_6721,N_4781,N_4714);
nor U6722 (N_6722,N_5900,N_5896);
nand U6723 (N_6723,N_4916,N_4016);
or U6724 (N_6724,N_4377,N_4969);
and U6725 (N_6725,N_4346,N_5995);
and U6726 (N_6726,N_5576,N_4958);
nor U6727 (N_6727,N_4763,N_5247);
or U6728 (N_6728,N_5568,N_4194);
or U6729 (N_6729,N_4430,N_5093);
nor U6730 (N_6730,N_4219,N_5138);
or U6731 (N_6731,N_4439,N_4657);
nor U6732 (N_6732,N_4862,N_4271);
nand U6733 (N_6733,N_4933,N_4425);
or U6734 (N_6734,N_4644,N_5299);
or U6735 (N_6735,N_5951,N_4742);
nor U6736 (N_6736,N_5832,N_4802);
and U6737 (N_6737,N_4235,N_4849);
or U6738 (N_6738,N_4116,N_5517);
nor U6739 (N_6739,N_5027,N_4250);
nand U6740 (N_6740,N_5387,N_4758);
nand U6741 (N_6741,N_5158,N_4326);
or U6742 (N_6742,N_4345,N_5675);
nor U6743 (N_6743,N_5227,N_4551);
nor U6744 (N_6744,N_5228,N_4388);
nand U6745 (N_6745,N_5884,N_5005);
nand U6746 (N_6746,N_4791,N_4755);
or U6747 (N_6747,N_4536,N_5841);
nand U6748 (N_6748,N_5392,N_5573);
nor U6749 (N_6749,N_4398,N_4373);
nand U6750 (N_6750,N_5353,N_4533);
nand U6751 (N_6751,N_4831,N_4636);
and U6752 (N_6752,N_5302,N_5628);
or U6753 (N_6753,N_4115,N_4068);
nor U6754 (N_6754,N_5181,N_5340);
nand U6755 (N_6755,N_5810,N_5683);
nand U6756 (N_6756,N_4423,N_4372);
nor U6757 (N_6757,N_4188,N_5789);
nor U6758 (N_6758,N_4527,N_4261);
nand U6759 (N_6759,N_5462,N_5609);
nor U6760 (N_6760,N_5175,N_5667);
and U6761 (N_6761,N_4191,N_5850);
nor U6762 (N_6762,N_4196,N_4167);
and U6763 (N_6763,N_5295,N_4599);
nor U6764 (N_6764,N_4756,N_5217);
or U6765 (N_6765,N_4109,N_5230);
or U6766 (N_6766,N_4160,N_5580);
nand U6767 (N_6767,N_5173,N_4681);
nor U6768 (N_6768,N_4004,N_5725);
nor U6769 (N_6769,N_4804,N_5233);
nand U6770 (N_6770,N_4395,N_5406);
or U6771 (N_6771,N_4555,N_5412);
and U6772 (N_6772,N_4640,N_5791);
or U6773 (N_6773,N_5603,N_5542);
nor U6774 (N_6774,N_5539,N_4204);
or U6775 (N_6775,N_4621,N_4003);
or U6776 (N_6776,N_5000,N_5604);
nor U6777 (N_6777,N_5341,N_4797);
nor U6778 (N_6778,N_5322,N_5708);
and U6779 (N_6779,N_5969,N_4977);
and U6780 (N_6780,N_5764,N_4617);
and U6781 (N_6781,N_4675,N_4808);
and U6782 (N_6782,N_5376,N_5216);
and U6783 (N_6783,N_4557,N_4945);
nor U6784 (N_6784,N_4342,N_4019);
nor U6785 (N_6785,N_5114,N_4438);
nor U6786 (N_6786,N_4915,N_4298);
and U6787 (N_6787,N_4272,N_4992);
or U6788 (N_6788,N_4097,N_4031);
and U6789 (N_6789,N_4437,N_5105);
and U6790 (N_6790,N_4367,N_5661);
nand U6791 (N_6791,N_5139,N_5945);
or U6792 (N_6792,N_4498,N_4355);
and U6793 (N_6793,N_5619,N_4702);
and U6794 (N_6794,N_5257,N_4569);
or U6795 (N_6795,N_5263,N_4393);
or U6796 (N_6796,N_5280,N_4592);
and U6797 (N_6797,N_5926,N_4077);
and U6798 (N_6798,N_4480,N_4932);
nand U6799 (N_6799,N_5625,N_5964);
or U6800 (N_6800,N_4451,N_4252);
nor U6801 (N_6801,N_5757,N_4887);
nor U6802 (N_6802,N_4161,N_4769);
nand U6803 (N_6803,N_5061,N_5469);
nand U6804 (N_6804,N_4874,N_5746);
nor U6805 (N_6805,N_4024,N_5634);
or U6806 (N_6806,N_5638,N_4500);
or U6807 (N_6807,N_4386,N_4762);
or U6808 (N_6808,N_5735,N_4479);
and U6809 (N_6809,N_4348,N_5892);
nand U6810 (N_6810,N_5618,N_4717);
nand U6811 (N_6811,N_4080,N_4950);
nor U6812 (N_6812,N_4410,N_4029);
nand U6813 (N_6813,N_5149,N_5255);
nand U6814 (N_6814,N_4867,N_4364);
nor U6815 (N_6815,N_5200,N_5730);
or U6816 (N_6816,N_4811,N_5784);
nand U6817 (N_6817,N_5817,N_5403);
nor U6818 (N_6818,N_5656,N_5736);
nand U6819 (N_6819,N_4564,N_5760);
or U6820 (N_6820,N_4818,N_5565);
or U6821 (N_6821,N_5186,N_5777);
and U6822 (N_6822,N_5153,N_4510);
and U6823 (N_6823,N_4577,N_5146);
and U6824 (N_6824,N_4291,N_5770);
nor U6825 (N_6825,N_4907,N_4098);
nand U6826 (N_6826,N_5194,N_4520);
and U6827 (N_6827,N_4971,N_5890);
or U6828 (N_6828,N_5420,N_4037);
nand U6829 (N_6829,N_5635,N_5811);
nand U6830 (N_6830,N_5016,N_4611);
nand U6831 (N_6831,N_4414,N_4470);
and U6832 (N_6832,N_4628,N_5540);
or U6833 (N_6833,N_4449,N_5404);
xor U6834 (N_6834,N_5229,N_4854);
and U6835 (N_6835,N_5514,N_4456);
or U6836 (N_6836,N_4544,N_4231);
or U6837 (N_6837,N_5495,N_4312);
nor U6838 (N_6838,N_4069,N_5183);
and U6839 (N_6839,N_5526,N_4690);
and U6840 (N_6840,N_4678,N_4284);
and U6841 (N_6841,N_5174,N_4799);
xnor U6842 (N_6842,N_5935,N_4779);
or U6843 (N_6843,N_5373,N_5214);
or U6844 (N_6844,N_5767,N_4596);
and U6845 (N_6845,N_5014,N_4266);
and U6846 (N_6846,N_5664,N_5804);
nor U6847 (N_6847,N_4338,N_4575);
nand U6848 (N_6848,N_5449,N_5205);
nand U6849 (N_6849,N_5467,N_4258);
nand U6850 (N_6850,N_4543,N_4055);
nand U6851 (N_6851,N_5075,N_5924);
and U6852 (N_6852,N_5998,N_5673);
or U6853 (N_6853,N_4376,N_4540);
nor U6854 (N_6854,N_5966,N_5652);
nor U6855 (N_6855,N_4089,N_4917);
nand U6856 (N_6856,N_4923,N_5880);
nor U6857 (N_6857,N_4182,N_4221);
and U6858 (N_6858,N_4972,N_4350);
or U6859 (N_6859,N_4127,N_4174);
and U6860 (N_6860,N_5724,N_5701);
or U6861 (N_6861,N_5458,N_5871);
and U6862 (N_6862,N_4073,N_4893);
and U6863 (N_6863,N_4363,N_5422);
and U6864 (N_6864,N_5025,N_5351);
nor U6865 (N_6865,N_4654,N_4111);
nand U6866 (N_6866,N_5226,N_4351);
nor U6867 (N_6867,N_5451,N_4466);
and U6868 (N_6868,N_5927,N_4774);
nor U6869 (N_6869,N_5137,N_5035);
or U6870 (N_6870,N_5533,N_4095);
and U6871 (N_6871,N_5589,N_5104);
or U6872 (N_6872,N_4384,N_5721);
nand U6873 (N_6873,N_5801,N_5556);
and U6874 (N_6874,N_5487,N_5043);
or U6875 (N_6875,N_4800,N_5191);
nor U6876 (N_6876,N_5606,N_5666);
nor U6877 (N_6877,N_5172,N_4724);
nor U6878 (N_6878,N_4286,N_4754);
nor U6879 (N_6879,N_5437,N_4049);
nor U6880 (N_6880,N_4944,N_4926);
or U6881 (N_6881,N_4597,N_4443);
nand U6882 (N_6882,N_4166,N_5711);
and U6883 (N_6883,N_5089,N_5732);
nand U6884 (N_6884,N_5047,N_4458);
nor U6885 (N_6885,N_5587,N_5501);
nand U6886 (N_6886,N_5671,N_4232);
and U6887 (N_6887,N_5270,N_4626);
or U6888 (N_6888,N_4633,N_4805);
nor U6889 (N_6889,N_5729,N_5366);
nor U6890 (N_6890,N_4594,N_5262);
and U6891 (N_6891,N_5218,N_4878);
and U6892 (N_6892,N_5869,N_4145);
nand U6893 (N_6893,N_5222,N_4032);
nand U6894 (N_6894,N_4528,N_5256);
and U6895 (N_6895,N_4691,N_4297);
nand U6896 (N_6896,N_4096,N_5152);
nor U6897 (N_6897,N_4023,N_4316);
or U6898 (N_6898,N_4140,N_5008);
nand U6899 (N_6899,N_4868,N_5778);
or U6900 (N_6900,N_4728,N_4965);
nand U6901 (N_6901,N_5432,N_5042);
nor U6902 (N_6902,N_4580,N_5631);
or U6903 (N_6903,N_4431,N_5265);
or U6904 (N_6904,N_5867,N_5827);
nor U6905 (N_6905,N_4078,N_5504);
nand U6906 (N_6906,N_5335,N_4100);
and U6907 (N_6907,N_4736,N_4315);
and U6908 (N_6908,N_5710,N_4910);
and U6909 (N_6909,N_5605,N_4821);
nand U6910 (N_6910,N_4228,N_5597);
or U6911 (N_6911,N_4509,N_4124);
or U6912 (N_6912,N_4588,N_5855);
or U6913 (N_6913,N_4102,N_4646);
and U6914 (N_6914,N_4413,N_4146);
and U6915 (N_6915,N_5011,N_4780);
or U6916 (N_6916,N_4886,N_5246);
or U6917 (N_6917,N_5090,N_5455);
nand U6918 (N_6918,N_5276,N_5374);
nor U6919 (N_6919,N_5443,N_5980);
and U6920 (N_6920,N_5323,N_4106);
nand U6921 (N_6921,N_4322,N_4876);
or U6922 (N_6922,N_4420,N_5552);
nor U6923 (N_6923,N_4574,N_4957);
and U6924 (N_6924,N_5883,N_5755);
and U6925 (N_6925,N_4268,N_5835);
nand U6926 (N_6926,N_5017,N_5337);
nor U6927 (N_6927,N_4604,N_4434);
nand U6928 (N_6928,N_4308,N_5698);
nand U6929 (N_6929,N_5002,N_5020);
and U6930 (N_6930,N_4177,N_4942);
or U6931 (N_6931,N_5690,N_4656);
or U6932 (N_6932,N_5284,N_5530);
nor U6933 (N_6933,N_4525,N_4719);
and U6934 (N_6934,N_4841,N_4371);
nor U6935 (N_6935,N_4770,N_4053);
or U6936 (N_6936,N_5028,N_5637);
or U6937 (N_6937,N_4005,N_4058);
and U6938 (N_6938,N_4623,N_5080);
or U6939 (N_6939,N_4552,N_4844);
xor U6940 (N_6940,N_4618,N_5968);
nor U6941 (N_6941,N_5239,N_4052);
nand U6942 (N_6942,N_4245,N_4403);
nor U6943 (N_6943,N_4164,N_4184);
nor U6944 (N_6944,N_5293,N_4343);
nor U6945 (N_6945,N_5251,N_5056);
nor U6946 (N_6946,N_5304,N_5716);
nand U6947 (N_6947,N_5427,N_5763);
nor U6948 (N_6948,N_5692,N_4857);
or U6949 (N_6949,N_5987,N_5672);
nand U6950 (N_6950,N_4021,N_4463);
or U6951 (N_6951,N_4827,N_4064);
and U6952 (N_6952,N_4968,N_4300);
or U6953 (N_6953,N_5377,N_5594);
and U6954 (N_6954,N_4900,N_4270);
and U6955 (N_6955,N_4980,N_4872);
nor U6956 (N_6956,N_5534,N_5515);
nand U6957 (N_6957,N_4459,N_5010);
or U6958 (N_6958,N_5786,N_5371);
nor U6959 (N_6959,N_5833,N_5865);
nand U6960 (N_6960,N_4936,N_5491);
and U6961 (N_6961,N_5163,N_4729);
and U6962 (N_6962,N_5644,N_4415);
or U6963 (N_6963,N_5470,N_5541);
nor U6964 (N_6964,N_5921,N_5120);
nor U6965 (N_6965,N_4446,N_5704);
or U6966 (N_6966,N_4747,N_5965);
or U6967 (N_6967,N_5902,N_5988);
or U6968 (N_6968,N_4209,N_4966);
or U6969 (N_6969,N_5242,N_4642);
nor U6970 (N_6970,N_5563,N_4390);
and U6971 (N_6971,N_5925,N_5065);
and U6972 (N_6972,N_4712,N_5640);
nand U6973 (N_6973,N_5461,N_4094);
nand U6974 (N_6974,N_5102,N_4426);
and U6975 (N_6975,N_5614,N_5788);
and U6976 (N_6976,N_4680,N_4812);
nor U6977 (N_6977,N_4155,N_4493);
or U6978 (N_6978,N_5523,N_4303);
or U6979 (N_6979,N_5821,N_4001);
nor U6980 (N_6980,N_5658,N_5574);
and U6981 (N_6981,N_4850,N_5375);
or U6982 (N_6982,N_5310,N_4485);
and U6983 (N_6983,N_4861,N_4859);
or U6984 (N_6984,N_4020,N_5874);
and U6985 (N_6985,N_4902,N_4809);
nor U6986 (N_6986,N_5668,N_4700);
or U6987 (N_6987,N_4707,N_5122);
and U6988 (N_6988,N_4172,N_4281);
nand U6989 (N_6989,N_4919,N_4630);
and U6990 (N_6990,N_5499,N_4394);
nand U6991 (N_6991,N_4549,N_4863);
nand U6992 (N_6992,N_5211,N_4605);
nor U6993 (N_6993,N_5520,N_4275);
and U6994 (N_6994,N_4189,N_5842);
nor U6995 (N_6995,N_4356,N_5894);
or U6996 (N_6996,N_4296,N_5857);
or U6997 (N_6997,N_5321,N_4051);
or U6998 (N_6998,N_4283,N_4582);
or U6999 (N_6999,N_4030,N_5204);
and U7000 (N_7000,N_4765,N_5584);
or U7001 (N_7001,N_5751,N_4892);
nor U7002 (N_7002,N_5230,N_5035);
or U7003 (N_7003,N_5132,N_4838);
or U7004 (N_7004,N_4478,N_4229);
nand U7005 (N_7005,N_5187,N_4011);
and U7006 (N_7006,N_5057,N_5807);
and U7007 (N_7007,N_5206,N_5804);
and U7008 (N_7008,N_5455,N_5317);
nor U7009 (N_7009,N_5133,N_4873);
nor U7010 (N_7010,N_5847,N_4289);
nand U7011 (N_7011,N_4696,N_5782);
or U7012 (N_7012,N_4023,N_5936);
nor U7013 (N_7013,N_5687,N_4333);
and U7014 (N_7014,N_5636,N_4876);
nand U7015 (N_7015,N_4174,N_5536);
nor U7016 (N_7016,N_5815,N_5031);
nand U7017 (N_7017,N_5866,N_4445);
or U7018 (N_7018,N_4266,N_5535);
nor U7019 (N_7019,N_5712,N_5273);
and U7020 (N_7020,N_4386,N_4960);
or U7021 (N_7021,N_4344,N_4906);
and U7022 (N_7022,N_5207,N_5213);
or U7023 (N_7023,N_4593,N_4829);
and U7024 (N_7024,N_5780,N_5066);
nor U7025 (N_7025,N_4345,N_4335);
or U7026 (N_7026,N_5502,N_5859);
or U7027 (N_7027,N_4352,N_5491);
nand U7028 (N_7028,N_5266,N_5752);
nor U7029 (N_7029,N_4492,N_5171);
nand U7030 (N_7030,N_4949,N_5100);
or U7031 (N_7031,N_5445,N_5621);
or U7032 (N_7032,N_4004,N_5105);
and U7033 (N_7033,N_4922,N_5202);
and U7034 (N_7034,N_5789,N_5351);
and U7035 (N_7035,N_4981,N_5671);
and U7036 (N_7036,N_4858,N_5033);
nand U7037 (N_7037,N_4771,N_5382);
nor U7038 (N_7038,N_5770,N_5309);
and U7039 (N_7039,N_4858,N_4720);
nand U7040 (N_7040,N_4220,N_4928);
nor U7041 (N_7041,N_5891,N_5473);
nand U7042 (N_7042,N_5305,N_4373);
nor U7043 (N_7043,N_4299,N_5341);
or U7044 (N_7044,N_5676,N_4557);
or U7045 (N_7045,N_4635,N_4992);
or U7046 (N_7046,N_5086,N_4471);
nand U7047 (N_7047,N_4707,N_5226);
nand U7048 (N_7048,N_5701,N_4112);
xnor U7049 (N_7049,N_5500,N_5064);
and U7050 (N_7050,N_5351,N_5217);
nand U7051 (N_7051,N_4176,N_5437);
or U7052 (N_7052,N_5075,N_4251);
nand U7053 (N_7053,N_4226,N_5582);
nand U7054 (N_7054,N_5522,N_4492);
nand U7055 (N_7055,N_4122,N_5722);
and U7056 (N_7056,N_5050,N_5240);
nor U7057 (N_7057,N_5009,N_5574);
nor U7058 (N_7058,N_5267,N_4196);
or U7059 (N_7059,N_4853,N_4293);
nand U7060 (N_7060,N_5003,N_5198);
nor U7061 (N_7061,N_5328,N_4753);
and U7062 (N_7062,N_4014,N_5969);
nand U7063 (N_7063,N_4238,N_4204);
nand U7064 (N_7064,N_5859,N_5597);
nor U7065 (N_7065,N_5757,N_5081);
nor U7066 (N_7066,N_5775,N_5801);
xnor U7067 (N_7067,N_5015,N_5609);
or U7068 (N_7068,N_4237,N_5179);
or U7069 (N_7069,N_4077,N_5942);
xor U7070 (N_7070,N_5076,N_4979);
nand U7071 (N_7071,N_4932,N_5477);
nand U7072 (N_7072,N_5506,N_5314);
nor U7073 (N_7073,N_5817,N_5093);
nand U7074 (N_7074,N_4079,N_4483);
or U7075 (N_7075,N_5106,N_4429);
or U7076 (N_7076,N_5766,N_4287);
and U7077 (N_7077,N_4593,N_4308);
nor U7078 (N_7078,N_4694,N_4156);
or U7079 (N_7079,N_4956,N_4864);
or U7080 (N_7080,N_4804,N_5916);
or U7081 (N_7081,N_4695,N_5452);
or U7082 (N_7082,N_4319,N_4680);
nor U7083 (N_7083,N_5286,N_4830);
nand U7084 (N_7084,N_4454,N_5590);
or U7085 (N_7085,N_4765,N_5306);
nand U7086 (N_7086,N_4043,N_5277);
and U7087 (N_7087,N_5641,N_5263);
nand U7088 (N_7088,N_5164,N_4486);
nand U7089 (N_7089,N_4079,N_5869);
nor U7090 (N_7090,N_5780,N_5189);
and U7091 (N_7091,N_4116,N_4874);
or U7092 (N_7092,N_5666,N_4536);
and U7093 (N_7093,N_5767,N_5017);
nand U7094 (N_7094,N_4748,N_5073);
nor U7095 (N_7095,N_4481,N_5012);
or U7096 (N_7096,N_5374,N_4493);
and U7097 (N_7097,N_5445,N_4827);
or U7098 (N_7098,N_4166,N_5105);
nand U7099 (N_7099,N_5280,N_4620);
or U7100 (N_7100,N_4640,N_5678);
nand U7101 (N_7101,N_5370,N_5130);
or U7102 (N_7102,N_4308,N_5191);
nor U7103 (N_7103,N_5776,N_5311);
and U7104 (N_7104,N_5483,N_4163);
and U7105 (N_7105,N_5188,N_4235);
or U7106 (N_7106,N_5968,N_4432);
nand U7107 (N_7107,N_4053,N_4152);
or U7108 (N_7108,N_4802,N_5627);
and U7109 (N_7109,N_4744,N_5102);
nor U7110 (N_7110,N_5332,N_5159);
or U7111 (N_7111,N_5616,N_5149);
nand U7112 (N_7112,N_5249,N_4881);
nor U7113 (N_7113,N_4740,N_4710);
or U7114 (N_7114,N_5386,N_4972);
nand U7115 (N_7115,N_5043,N_5007);
nor U7116 (N_7116,N_4977,N_5249);
and U7117 (N_7117,N_5732,N_5498);
nor U7118 (N_7118,N_4628,N_4456);
or U7119 (N_7119,N_5608,N_4637);
and U7120 (N_7120,N_4147,N_4331);
and U7121 (N_7121,N_5306,N_4651);
or U7122 (N_7122,N_5576,N_5916);
nand U7123 (N_7123,N_5522,N_5213);
nand U7124 (N_7124,N_5925,N_5049);
or U7125 (N_7125,N_5955,N_4505);
nand U7126 (N_7126,N_5859,N_4747);
nand U7127 (N_7127,N_4530,N_5683);
nor U7128 (N_7128,N_4277,N_4575);
nand U7129 (N_7129,N_4084,N_4285);
nand U7130 (N_7130,N_5829,N_5051);
or U7131 (N_7131,N_4421,N_4810);
and U7132 (N_7132,N_4025,N_4810);
and U7133 (N_7133,N_4560,N_4687);
and U7134 (N_7134,N_4974,N_4146);
or U7135 (N_7135,N_5474,N_4048);
or U7136 (N_7136,N_4975,N_5470);
nor U7137 (N_7137,N_5810,N_5997);
or U7138 (N_7138,N_5765,N_4185);
nor U7139 (N_7139,N_5191,N_5797);
or U7140 (N_7140,N_5282,N_5491);
nor U7141 (N_7141,N_4253,N_4484);
nor U7142 (N_7142,N_4555,N_5230);
nand U7143 (N_7143,N_5751,N_5802);
nand U7144 (N_7144,N_5395,N_4820);
or U7145 (N_7145,N_5385,N_4865);
or U7146 (N_7146,N_4328,N_4243);
nor U7147 (N_7147,N_4798,N_4042);
nor U7148 (N_7148,N_4963,N_4086);
and U7149 (N_7149,N_5889,N_5805);
or U7150 (N_7150,N_5100,N_4309);
nor U7151 (N_7151,N_4107,N_5012);
nand U7152 (N_7152,N_4797,N_5241);
nor U7153 (N_7153,N_5704,N_4376);
and U7154 (N_7154,N_4452,N_4650);
nand U7155 (N_7155,N_4484,N_4338);
and U7156 (N_7156,N_5742,N_5891);
nand U7157 (N_7157,N_4287,N_4402);
nor U7158 (N_7158,N_4495,N_5511);
nor U7159 (N_7159,N_4893,N_4147);
nand U7160 (N_7160,N_4473,N_5022);
or U7161 (N_7161,N_5272,N_4242);
nand U7162 (N_7162,N_5444,N_5788);
nor U7163 (N_7163,N_5141,N_5416);
and U7164 (N_7164,N_5932,N_4214);
or U7165 (N_7165,N_4529,N_5730);
nor U7166 (N_7166,N_4973,N_5034);
and U7167 (N_7167,N_5879,N_5158);
nor U7168 (N_7168,N_5939,N_4679);
nand U7169 (N_7169,N_5609,N_5179);
nor U7170 (N_7170,N_5020,N_4596);
and U7171 (N_7171,N_4686,N_4794);
and U7172 (N_7172,N_4009,N_4832);
xor U7173 (N_7173,N_5750,N_4145);
nor U7174 (N_7174,N_5063,N_4189);
or U7175 (N_7175,N_4559,N_5733);
and U7176 (N_7176,N_4143,N_5956);
or U7177 (N_7177,N_4090,N_5762);
or U7178 (N_7178,N_4146,N_5549);
and U7179 (N_7179,N_5795,N_4992);
or U7180 (N_7180,N_5911,N_4271);
or U7181 (N_7181,N_5931,N_5655);
nand U7182 (N_7182,N_5263,N_4942);
nand U7183 (N_7183,N_4173,N_4607);
or U7184 (N_7184,N_5260,N_4935);
and U7185 (N_7185,N_5035,N_5239);
or U7186 (N_7186,N_5746,N_5510);
or U7187 (N_7187,N_5918,N_4666);
nor U7188 (N_7188,N_5085,N_5578);
and U7189 (N_7189,N_5143,N_4558);
and U7190 (N_7190,N_5305,N_4996);
or U7191 (N_7191,N_5357,N_5018);
and U7192 (N_7192,N_4823,N_5371);
or U7193 (N_7193,N_4357,N_5595);
or U7194 (N_7194,N_5586,N_5722);
and U7195 (N_7195,N_5619,N_4441);
and U7196 (N_7196,N_5154,N_5984);
and U7197 (N_7197,N_4627,N_4636);
nor U7198 (N_7198,N_5350,N_5667);
nor U7199 (N_7199,N_4711,N_4772);
and U7200 (N_7200,N_4705,N_4103);
nand U7201 (N_7201,N_4044,N_5844);
nor U7202 (N_7202,N_5264,N_5761);
or U7203 (N_7203,N_4936,N_4154);
or U7204 (N_7204,N_5471,N_4150);
or U7205 (N_7205,N_5111,N_4129);
and U7206 (N_7206,N_4383,N_5236);
or U7207 (N_7207,N_4016,N_4435);
or U7208 (N_7208,N_4740,N_4964);
and U7209 (N_7209,N_4531,N_4478);
nor U7210 (N_7210,N_5557,N_4794);
nand U7211 (N_7211,N_5430,N_5812);
or U7212 (N_7212,N_4871,N_5860);
and U7213 (N_7213,N_5082,N_5651);
nor U7214 (N_7214,N_4036,N_5326);
nand U7215 (N_7215,N_5554,N_5136);
nand U7216 (N_7216,N_4843,N_5821);
nor U7217 (N_7217,N_4506,N_5970);
nand U7218 (N_7218,N_4610,N_5642);
nor U7219 (N_7219,N_4020,N_4956);
nand U7220 (N_7220,N_4844,N_5683);
nand U7221 (N_7221,N_5767,N_5943);
nor U7222 (N_7222,N_4907,N_5061);
nor U7223 (N_7223,N_4362,N_5023);
and U7224 (N_7224,N_5174,N_4728);
nand U7225 (N_7225,N_5256,N_5165);
nor U7226 (N_7226,N_5385,N_4586);
nand U7227 (N_7227,N_4615,N_5551);
and U7228 (N_7228,N_5747,N_4606);
nand U7229 (N_7229,N_5898,N_4658);
or U7230 (N_7230,N_4063,N_4104);
or U7231 (N_7231,N_4495,N_4216);
nor U7232 (N_7232,N_4426,N_4451);
and U7233 (N_7233,N_5691,N_4385);
nand U7234 (N_7234,N_5570,N_4269);
or U7235 (N_7235,N_5273,N_5749);
or U7236 (N_7236,N_4366,N_4521);
or U7237 (N_7237,N_4876,N_5331);
nor U7238 (N_7238,N_4971,N_5132);
nand U7239 (N_7239,N_5048,N_4076);
nor U7240 (N_7240,N_5749,N_5852);
nor U7241 (N_7241,N_5166,N_4456);
or U7242 (N_7242,N_4528,N_5249);
nor U7243 (N_7243,N_4988,N_4456);
nor U7244 (N_7244,N_4958,N_4203);
and U7245 (N_7245,N_4872,N_5141);
or U7246 (N_7246,N_4773,N_4562);
and U7247 (N_7247,N_5087,N_5055);
or U7248 (N_7248,N_4986,N_5989);
nand U7249 (N_7249,N_5950,N_5816);
and U7250 (N_7250,N_4962,N_4679);
or U7251 (N_7251,N_5154,N_4082);
xor U7252 (N_7252,N_5202,N_5005);
and U7253 (N_7253,N_5167,N_5489);
or U7254 (N_7254,N_5590,N_4168);
nand U7255 (N_7255,N_5725,N_5511);
or U7256 (N_7256,N_5859,N_5870);
nand U7257 (N_7257,N_5385,N_5960);
nand U7258 (N_7258,N_4585,N_5846);
nand U7259 (N_7259,N_4381,N_5689);
nor U7260 (N_7260,N_4636,N_5117);
nor U7261 (N_7261,N_4990,N_5830);
or U7262 (N_7262,N_5784,N_4906);
nor U7263 (N_7263,N_4761,N_5906);
nor U7264 (N_7264,N_5175,N_4794);
nand U7265 (N_7265,N_4061,N_5292);
or U7266 (N_7266,N_5625,N_5196);
or U7267 (N_7267,N_5847,N_5502);
and U7268 (N_7268,N_5396,N_4299);
nand U7269 (N_7269,N_4088,N_5887);
nand U7270 (N_7270,N_5935,N_4943);
or U7271 (N_7271,N_4958,N_5158);
or U7272 (N_7272,N_4300,N_5662);
nor U7273 (N_7273,N_5591,N_4678);
nor U7274 (N_7274,N_5322,N_5541);
or U7275 (N_7275,N_4751,N_4922);
nor U7276 (N_7276,N_5760,N_5296);
nor U7277 (N_7277,N_5839,N_4428);
or U7278 (N_7278,N_4558,N_5551);
and U7279 (N_7279,N_4712,N_5284);
nor U7280 (N_7280,N_5357,N_5233);
and U7281 (N_7281,N_4017,N_4037);
or U7282 (N_7282,N_5517,N_5336);
nor U7283 (N_7283,N_4241,N_4743);
and U7284 (N_7284,N_4617,N_5200);
nor U7285 (N_7285,N_5003,N_4486);
nand U7286 (N_7286,N_5869,N_5777);
and U7287 (N_7287,N_5636,N_5962);
or U7288 (N_7288,N_5617,N_5470);
and U7289 (N_7289,N_5373,N_5080);
nand U7290 (N_7290,N_4119,N_4256);
or U7291 (N_7291,N_4882,N_5944);
nor U7292 (N_7292,N_4516,N_4780);
nor U7293 (N_7293,N_4155,N_5705);
or U7294 (N_7294,N_5305,N_4082);
nand U7295 (N_7295,N_5626,N_4212);
or U7296 (N_7296,N_4308,N_5573);
nor U7297 (N_7297,N_5893,N_4235);
nand U7298 (N_7298,N_5696,N_5900);
and U7299 (N_7299,N_5176,N_4302);
nand U7300 (N_7300,N_5018,N_4431);
and U7301 (N_7301,N_5303,N_5147);
or U7302 (N_7302,N_4737,N_5056);
nor U7303 (N_7303,N_4300,N_5380);
nor U7304 (N_7304,N_4498,N_4291);
or U7305 (N_7305,N_5146,N_4932);
or U7306 (N_7306,N_4366,N_5226);
and U7307 (N_7307,N_4886,N_5723);
nand U7308 (N_7308,N_4841,N_4763);
or U7309 (N_7309,N_5923,N_4644);
nand U7310 (N_7310,N_4866,N_5481);
nor U7311 (N_7311,N_5759,N_5424);
nor U7312 (N_7312,N_4443,N_4718);
nand U7313 (N_7313,N_4847,N_5567);
nand U7314 (N_7314,N_4192,N_5642);
nor U7315 (N_7315,N_4104,N_4266);
and U7316 (N_7316,N_5821,N_5205);
or U7317 (N_7317,N_4321,N_5015);
or U7318 (N_7318,N_4334,N_4387);
nand U7319 (N_7319,N_4392,N_5105);
and U7320 (N_7320,N_4204,N_4228);
and U7321 (N_7321,N_5755,N_4285);
nand U7322 (N_7322,N_5066,N_5243);
or U7323 (N_7323,N_4357,N_5338);
nand U7324 (N_7324,N_5939,N_4295);
nand U7325 (N_7325,N_5515,N_4811);
and U7326 (N_7326,N_4325,N_4544);
and U7327 (N_7327,N_4438,N_4390);
nor U7328 (N_7328,N_5369,N_5427);
nor U7329 (N_7329,N_4987,N_5008);
nor U7330 (N_7330,N_4016,N_5676);
nand U7331 (N_7331,N_4600,N_5623);
nand U7332 (N_7332,N_5194,N_5009);
nor U7333 (N_7333,N_4073,N_4415);
nand U7334 (N_7334,N_4609,N_5470);
or U7335 (N_7335,N_4600,N_5346);
nor U7336 (N_7336,N_5891,N_4323);
and U7337 (N_7337,N_4923,N_5280);
xor U7338 (N_7338,N_4054,N_5361);
and U7339 (N_7339,N_4533,N_5160);
or U7340 (N_7340,N_5929,N_4863);
and U7341 (N_7341,N_4490,N_4244);
and U7342 (N_7342,N_5930,N_4788);
or U7343 (N_7343,N_5817,N_4236);
nor U7344 (N_7344,N_5017,N_5394);
or U7345 (N_7345,N_4210,N_4657);
nand U7346 (N_7346,N_4214,N_5702);
and U7347 (N_7347,N_4643,N_4371);
and U7348 (N_7348,N_5683,N_5078);
nor U7349 (N_7349,N_5561,N_4115);
nor U7350 (N_7350,N_5626,N_4343);
nand U7351 (N_7351,N_4394,N_5475);
nor U7352 (N_7352,N_5113,N_4058);
and U7353 (N_7353,N_5293,N_5056);
nand U7354 (N_7354,N_4212,N_5132);
and U7355 (N_7355,N_4720,N_5763);
or U7356 (N_7356,N_5606,N_4594);
nor U7357 (N_7357,N_5037,N_5781);
nor U7358 (N_7358,N_5790,N_5413);
nand U7359 (N_7359,N_4916,N_4187);
and U7360 (N_7360,N_4874,N_5069);
nand U7361 (N_7361,N_5353,N_4903);
nor U7362 (N_7362,N_4785,N_5424);
and U7363 (N_7363,N_5311,N_5271);
nand U7364 (N_7364,N_5722,N_5562);
nand U7365 (N_7365,N_4600,N_5923);
or U7366 (N_7366,N_4071,N_4326);
and U7367 (N_7367,N_5384,N_4332);
or U7368 (N_7368,N_5470,N_4410);
or U7369 (N_7369,N_4419,N_4643);
nand U7370 (N_7370,N_4767,N_4762);
and U7371 (N_7371,N_4329,N_5873);
nand U7372 (N_7372,N_5284,N_4841);
nand U7373 (N_7373,N_4114,N_4963);
nor U7374 (N_7374,N_4353,N_5638);
and U7375 (N_7375,N_5788,N_4524);
or U7376 (N_7376,N_5208,N_5149);
and U7377 (N_7377,N_4345,N_4892);
nand U7378 (N_7378,N_4063,N_5816);
and U7379 (N_7379,N_5896,N_4838);
and U7380 (N_7380,N_5367,N_4372);
nor U7381 (N_7381,N_5092,N_5576);
or U7382 (N_7382,N_5209,N_5083);
and U7383 (N_7383,N_4069,N_4973);
and U7384 (N_7384,N_5026,N_5043);
nand U7385 (N_7385,N_5862,N_4791);
or U7386 (N_7386,N_4610,N_4224);
or U7387 (N_7387,N_4215,N_5694);
nor U7388 (N_7388,N_4070,N_4169);
or U7389 (N_7389,N_5942,N_4804);
or U7390 (N_7390,N_5037,N_5520);
and U7391 (N_7391,N_5734,N_4882);
and U7392 (N_7392,N_4343,N_4467);
and U7393 (N_7393,N_4875,N_4821);
or U7394 (N_7394,N_5172,N_4384);
and U7395 (N_7395,N_4253,N_5592);
nand U7396 (N_7396,N_4283,N_5277);
and U7397 (N_7397,N_5976,N_4555);
and U7398 (N_7398,N_4784,N_5255);
and U7399 (N_7399,N_4977,N_4664);
and U7400 (N_7400,N_4582,N_4456);
and U7401 (N_7401,N_4090,N_4151);
or U7402 (N_7402,N_5976,N_5210);
and U7403 (N_7403,N_4806,N_4446);
or U7404 (N_7404,N_4363,N_5547);
and U7405 (N_7405,N_4275,N_5920);
or U7406 (N_7406,N_4440,N_5010);
or U7407 (N_7407,N_5853,N_5119);
nor U7408 (N_7408,N_4517,N_5971);
nand U7409 (N_7409,N_4419,N_4008);
nand U7410 (N_7410,N_4444,N_5714);
and U7411 (N_7411,N_5713,N_5814);
or U7412 (N_7412,N_4750,N_4495);
nor U7413 (N_7413,N_4727,N_5741);
xor U7414 (N_7414,N_5366,N_5343);
or U7415 (N_7415,N_4079,N_4427);
or U7416 (N_7416,N_4562,N_4116);
and U7417 (N_7417,N_4452,N_5722);
nand U7418 (N_7418,N_4369,N_5715);
nand U7419 (N_7419,N_5568,N_4280);
nand U7420 (N_7420,N_5858,N_4215);
nand U7421 (N_7421,N_4271,N_4573);
or U7422 (N_7422,N_5899,N_5688);
and U7423 (N_7423,N_5408,N_4071);
or U7424 (N_7424,N_4398,N_5525);
and U7425 (N_7425,N_5420,N_4414);
nor U7426 (N_7426,N_5244,N_5439);
nand U7427 (N_7427,N_5654,N_5480);
nand U7428 (N_7428,N_5914,N_5031);
nand U7429 (N_7429,N_4783,N_4454);
or U7430 (N_7430,N_5764,N_4742);
or U7431 (N_7431,N_4467,N_5596);
nand U7432 (N_7432,N_4490,N_4420);
and U7433 (N_7433,N_4864,N_4159);
and U7434 (N_7434,N_5542,N_4451);
nor U7435 (N_7435,N_4357,N_4081);
nand U7436 (N_7436,N_5184,N_5896);
nor U7437 (N_7437,N_5923,N_4236);
or U7438 (N_7438,N_5665,N_5399);
and U7439 (N_7439,N_4379,N_5788);
xor U7440 (N_7440,N_5711,N_4018);
and U7441 (N_7441,N_4465,N_5272);
and U7442 (N_7442,N_5074,N_4334);
or U7443 (N_7443,N_5547,N_4101);
and U7444 (N_7444,N_5328,N_4229);
or U7445 (N_7445,N_5575,N_4512);
or U7446 (N_7446,N_4956,N_5793);
nand U7447 (N_7447,N_4522,N_4807);
nand U7448 (N_7448,N_4315,N_5162);
nand U7449 (N_7449,N_5236,N_4282);
nor U7450 (N_7450,N_5579,N_5195);
or U7451 (N_7451,N_5827,N_5300);
nor U7452 (N_7452,N_5832,N_5414);
and U7453 (N_7453,N_5629,N_5498);
nand U7454 (N_7454,N_5586,N_4971);
nor U7455 (N_7455,N_5129,N_4546);
and U7456 (N_7456,N_4822,N_5720);
nand U7457 (N_7457,N_5825,N_5508);
nor U7458 (N_7458,N_4760,N_5309);
and U7459 (N_7459,N_4941,N_4137);
nor U7460 (N_7460,N_5540,N_5312);
nor U7461 (N_7461,N_4499,N_5356);
nor U7462 (N_7462,N_5018,N_5039);
and U7463 (N_7463,N_4045,N_4876);
nor U7464 (N_7464,N_5742,N_5500);
or U7465 (N_7465,N_5741,N_5615);
nand U7466 (N_7466,N_4609,N_5413);
nor U7467 (N_7467,N_5401,N_5451);
nand U7468 (N_7468,N_5338,N_5126);
nor U7469 (N_7469,N_4552,N_4567);
and U7470 (N_7470,N_4787,N_5545);
nand U7471 (N_7471,N_5689,N_5531);
nor U7472 (N_7472,N_5095,N_4672);
nor U7473 (N_7473,N_4403,N_5702);
or U7474 (N_7474,N_4232,N_5281);
xor U7475 (N_7475,N_4617,N_5726);
and U7476 (N_7476,N_4137,N_5288);
or U7477 (N_7477,N_4426,N_4636);
nor U7478 (N_7478,N_5290,N_4712);
nand U7479 (N_7479,N_4158,N_5398);
and U7480 (N_7480,N_5037,N_5317);
or U7481 (N_7481,N_5935,N_5633);
or U7482 (N_7482,N_5412,N_5541);
nand U7483 (N_7483,N_5536,N_5535);
nor U7484 (N_7484,N_4886,N_4571);
nor U7485 (N_7485,N_4101,N_4622);
nand U7486 (N_7486,N_4707,N_4577);
and U7487 (N_7487,N_5901,N_4864);
or U7488 (N_7488,N_4614,N_5488);
nor U7489 (N_7489,N_4931,N_5849);
and U7490 (N_7490,N_4283,N_4113);
nand U7491 (N_7491,N_4246,N_5782);
and U7492 (N_7492,N_4200,N_4481);
nand U7493 (N_7493,N_4062,N_4688);
or U7494 (N_7494,N_4057,N_4151);
nor U7495 (N_7495,N_5430,N_5876);
or U7496 (N_7496,N_4941,N_5523);
or U7497 (N_7497,N_5386,N_4462);
and U7498 (N_7498,N_4514,N_5479);
nand U7499 (N_7499,N_4812,N_5600);
or U7500 (N_7500,N_4552,N_5625);
nand U7501 (N_7501,N_5851,N_4881);
and U7502 (N_7502,N_4691,N_4500);
and U7503 (N_7503,N_5603,N_4446);
nand U7504 (N_7504,N_5707,N_5097);
nand U7505 (N_7505,N_4297,N_4721);
and U7506 (N_7506,N_5966,N_4847);
and U7507 (N_7507,N_4626,N_5996);
and U7508 (N_7508,N_4786,N_5143);
nand U7509 (N_7509,N_4803,N_4036);
or U7510 (N_7510,N_5563,N_4037);
or U7511 (N_7511,N_4507,N_5825);
nand U7512 (N_7512,N_4025,N_5168);
or U7513 (N_7513,N_4265,N_4831);
nor U7514 (N_7514,N_5712,N_5288);
nor U7515 (N_7515,N_5838,N_5223);
nand U7516 (N_7516,N_5228,N_5852);
nand U7517 (N_7517,N_4487,N_4272);
or U7518 (N_7518,N_4767,N_4442);
nand U7519 (N_7519,N_5505,N_4631);
nand U7520 (N_7520,N_4137,N_5226);
or U7521 (N_7521,N_4021,N_5144);
nand U7522 (N_7522,N_4927,N_4037);
nand U7523 (N_7523,N_5536,N_5115);
and U7524 (N_7524,N_5974,N_4528);
nand U7525 (N_7525,N_4598,N_5198);
or U7526 (N_7526,N_5092,N_4359);
nand U7527 (N_7527,N_5920,N_4619);
or U7528 (N_7528,N_4872,N_4726);
or U7529 (N_7529,N_4825,N_5963);
and U7530 (N_7530,N_5868,N_4126);
or U7531 (N_7531,N_4560,N_5189);
and U7532 (N_7532,N_4873,N_4176);
and U7533 (N_7533,N_5451,N_4290);
and U7534 (N_7534,N_4694,N_5267);
or U7535 (N_7535,N_5127,N_5102);
nor U7536 (N_7536,N_5478,N_5700);
or U7537 (N_7537,N_5439,N_4608);
and U7538 (N_7538,N_5396,N_4852);
and U7539 (N_7539,N_4569,N_4911);
nand U7540 (N_7540,N_5311,N_5662);
nor U7541 (N_7541,N_5142,N_5725);
or U7542 (N_7542,N_5921,N_4817);
nand U7543 (N_7543,N_4380,N_5125);
or U7544 (N_7544,N_4604,N_4986);
or U7545 (N_7545,N_5328,N_4954);
and U7546 (N_7546,N_4118,N_4099);
and U7547 (N_7547,N_4695,N_5300);
and U7548 (N_7548,N_5189,N_5260);
nor U7549 (N_7549,N_5809,N_4096);
and U7550 (N_7550,N_4061,N_4625);
nor U7551 (N_7551,N_4977,N_5595);
xnor U7552 (N_7552,N_5267,N_4391);
nand U7553 (N_7553,N_4010,N_5977);
nand U7554 (N_7554,N_4386,N_5804);
xor U7555 (N_7555,N_4689,N_4658);
nand U7556 (N_7556,N_4027,N_4579);
nor U7557 (N_7557,N_4649,N_4681);
nand U7558 (N_7558,N_4460,N_5917);
nand U7559 (N_7559,N_5538,N_5759);
nor U7560 (N_7560,N_4272,N_5548);
nand U7561 (N_7561,N_4735,N_4960);
or U7562 (N_7562,N_5588,N_4481);
nand U7563 (N_7563,N_4419,N_5949);
nand U7564 (N_7564,N_5154,N_4563);
or U7565 (N_7565,N_5073,N_5812);
nor U7566 (N_7566,N_4830,N_5982);
nor U7567 (N_7567,N_4322,N_4839);
nand U7568 (N_7568,N_4819,N_4902);
nand U7569 (N_7569,N_5518,N_5217);
or U7570 (N_7570,N_4932,N_4277);
nor U7571 (N_7571,N_4469,N_5723);
nor U7572 (N_7572,N_5352,N_4984);
nor U7573 (N_7573,N_5595,N_4194);
or U7574 (N_7574,N_4179,N_4332);
nand U7575 (N_7575,N_5723,N_4780);
or U7576 (N_7576,N_4487,N_4175);
and U7577 (N_7577,N_5033,N_5894);
nor U7578 (N_7578,N_5013,N_5825);
nand U7579 (N_7579,N_4660,N_5948);
nand U7580 (N_7580,N_5788,N_4766);
nor U7581 (N_7581,N_5142,N_4790);
nand U7582 (N_7582,N_4455,N_4883);
or U7583 (N_7583,N_5024,N_5558);
or U7584 (N_7584,N_4550,N_5879);
nand U7585 (N_7585,N_4593,N_5153);
and U7586 (N_7586,N_4773,N_4356);
or U7587 (N_7587,N_4609,N_4159);
or U7588 (N_7588,N_4707,N_4068);
nand U7589 (N_7589,N_5935,N_5024);
and U7590 (N_7590,N_5411,N_5799);
nor U7591 (N_7591,N_5476,N_4361);
or U7592 (N_7592,N_4745,N_5657);
nor U7593 (N_7593,N_5206,N_4740);
nor U7594 (N_7594,N_5792,N_4182);
nor U7595 (N_7595,N_5041,N_4957);
and U7596 (N_7596,N_4202,N_4891);
or U7597 (N_7597,N_4940,N_5467);
nand U7598 (N_7598,N_5301,N_5622);
and U7599 (N_7599,N_4600,N_4829);
or U7600 (N_7600,N_4186,N_4785);
nand U7601 (N_7601,N_4134,N_4442);
nand U7602 (N_7602,N_4652,N_4964);
or U7603 (N_7603,N_4518,N_5309);
nand U7604 (N_7604,N_5191,N_5990);
nand U7605 (N_7605,N_4443,N_4018);
or U7606 (N_7606,N_4531,N_4311);
or U7607 (N_7607,N_4645,N_4542);
nand U7608 (N_7608,N_4814,N_5971);
nand U7609 (N_7609,N_4762,N_5980);
nor U7610 (N_7610,N_4008,N_5788);
nand U7611 (N_7611,N_5819,N_5192);
or U7612 (N_7612,N_5230,N_5731);
nor U7613 (N_7613,N_4796,N_4514);
nor U7614 (N_7614,N_4595,N_4440);
or U7615 (N_7615,N_5468,N_5849);
nor U7616 (N_7616,N_5912,N_4218);
nand U7617 (N_7617,N_4698,N_5304);
and U7618 (N_7618,N_5191,N_5704);
and U7619 (N_7619,N_4447,N_4913);
nand U7620 (N_7620,N_4923,N_5169);
nor U7621 (N_7621,N_5538,N_5854);
or U7622 (N_7622,N_5755,N_4838);
nor U7623 (N_7623,N_4279,N_5122);
nor U7624 (N_7624,N_4949,N_5920);
or U7625 (N_7625,N_5597,N_4645);
or U7626 (N_7626,N_5217,N_4426);
nor U7627 (N_7627,N_5180,N_5030);
nor U7628 (N_7628,N_4911,N_4030);
xor U7629 (N_7629,N_4760,N_5678);
nor U7630 (N_7630,N_4401,N_5835);
or U7631 (N_7631,N_5845,N_4224);
nand U7632 (N_7632,N_4907,N_5583);
nand U7633 (N_7633,N_5093,N_4513);
and U7634 (N_7634,N_4541,N_4991);
and U7635 (N_7635,N_5287,N_5187);
or U7636 (N_7636,N_5827,N_5548);
nor U7637 (N_7637,N_5884,N_5019);
nand U7638 (N_7638,N_4979,N_5680);
nor U7639 (N_7639,N_5396,N_5642);
and U7640 (N_7640,N_5354,N_4938);
nand U7641 (N_7641,N_5358,N_5913);
nor U7642 (N_7642,N_4202,N_4878);
nand U7643 (N_7643,N_5838,N_5619);
or U7644 (N_7644,N_5084,N_4835);
nand U7645 (N_7645,N_5976,N_5694);
nand U7646 (N_7646,N_5820,N_5157);
xnor U7647 (N_7647,N_5721,N_5321);
nor U7648 (N_7648,N_4075,N_4407);
nand U7649 (N_7649,N_5816,N_5546);
and U7650 (N_7650,N_5526,N_5393);
nor U7651 (N_7651,N_5329,N_5721);
or U7652 (N_7652,N_4917,N_5137);
and U7653 (N_7653,N_4451,N_4628);
or U7654 (N_7654,N_4459,N_4130);
or U7655 (N_7655,N_5612,N_4398);
nor U7656 (N_7656,N_5539,N_4870);
nor U7657 (N_7657,N_5282,N_4872);
and U7658 (N_7658,N_5671,N_4367);
nand U7659 (N_7659,N_5618,N_4947);
nand U7660 (N_7660,N_5587,N_5957);
and U7661 (N_7661,N_5590,N_4196);
or U7662 (N_7662,N_5501,N_5371);
and U7663 (N_7663,N_4741,N_5762);
nand U7664 (N_7664,N_4088,N_5861);
nor U7665 (N_7665,N_4648,N_5531);
or U7666 (N_7666,N_5194,N_5874);
nand U7667 (N_7667,N_5121,N_5823);
nor U7668 (N_7668,N_5795,N_4569);
or U7669 (N_7669,N_4921,N_5281);
nand U7670 (N_7670,N_5377,N_5342);
nor U7671 (N_7671,N_4057,N_4277);
and U7672 (N_7672,N_4805,N_4573);
nand U7673 (N_7673,N_5318,N_4549);
or U7674 (N_7674,N_5059,N_4486);
nor U7675 (N_7675,N_4302,N_5440);
nor U7676 (N_7676,N_5380,N_5487);
nand U7677 (N_7677,N_4400,N_5424);
and U7678 (N_7678,N_5349,N_5895);
nand U7679 (N_7679,N_4303,N_4731);
and U7680 (N_7680,N_4699,N_5978);
and U7681 (N_7681,N_4575,N_5079);
nor U7682 (N_7682,N_4994,N_5692);
and U7683 (N_7683,N_4658,N_5679);
nand U7684 (N_7684,N_4792,N_4951);
nand U7685 (N_7685,N_5292,N_4842);
and U7686 (N_7686,N_5047,N_4535);
and U7687 (N_7687,N_4467,N_5039);
nor U7688 (N_7688,N_4086,N_4989);
or U7689 (N_7689,N_5875,N_5550);
or U7690 (N_7690,N_5579,N_4620);
nor U7691 (N_7691,N_4634,N_5142);
or U7692 (N_7692,N_5549,N_4624);
or U7693 (N_7693,N_4178,N_4535);
and U7694 (N_7694,N_4452,N_4028);
and U7695 (N_7695,N_4426,N_5239);
nor U7696 (N_7696,N_5156,N_5020);
or U7697 (N_7697,N_5463,N_4239);
or U7698 (N_7698,N_4882,N_4373);
nand U7699 (N_7699,N_4182,N_4269);
nand U7700 (N_7700,N_5732,N_4199);
or U7701 (N_7701,N_5902,N_4797);
nor U7702 (N_7702,N_5014,N_4173);
and U7703 (N_7703,N_4394,N_4221);
or U7704 (N_7704,N_4495,N_5831);
and U7705 (N_7705,N_4038,N_4031);
or U7706 (N_7706,N_4047,N_4767);
nand U7707 (N_7707,N_4256,N_5314);
or U7708 (N_7708,N_4343,N_4340);
nand U7709 (N_7709,N_4913,N_5970);
nor U7710 (N_7710,N_5626,N_5422);
nand U7711 (N_7711,N_4577,N_4649);
or U7712 (N_7712,N_4130,N_4953);
or U7713 (N_7713,N_5135,N_4752);
or U7714 (N_7714,N_5290,N_4643);
nand U7715 (N_7715,N_4016,N_5699);
xor U7716 (N_7716,N_5921,N_4432);
nor U7717 (N_7717,N_4357,N_4116);
nor U7718 (N_7718,N_5443,N_4650);
or U7719 (N_7719,N_4589,N_4245);
and U7720 (N_7720,N_4163,N_5967);
nand U7721 (N_7721,N_5027,N_4555);
or U7722 (N_7722,N_4640,N_5471);
and U7723 (N_7723,N_5880,N_4422);
nand U7724 (N_7724,N_5132,N_5692);
nor U7725 (N_7725,N_5627,N_4804);
or U7726 (N_7726,N_5649,N_5000);
or U7727 (N_7727,N_4434,N_5505);
and U7728 (N_7728,N_5904,N_5249);
nor U7729 (N_7729,N_4643,N_4980);
nor U7730 (N_7730,N_4918,N_4980);
nor U7731 (N_7731,N_5594,N_4569);
nand U7732 (N_7732,N_5376,N_5358);
and U7733 (N_7733,N_5045,N_5648);
or U7734 (N_7734,N_5541,N_4625);
and U7735 (N_7735,N_4664,N_4068);
and U7736 (N_7736,N_5390,N_4049);
and U7737 (N_7737,N_4874,N_4811);
nor U7738 (N_7738,N_4666,N_5258);
nand U7739 (N_7739,N_5559,N_5533);
nand U7740 (N_7740,N_5163,N_4546);
and U7741 (N_7741,N_4505,N_5275);
nor U7742 (N_7742,N_4678,N_4114);
nand U7743 (N_7743,N_4369,N_5788);
or U7744 (N_7744,N_4539,N_4652);
nor U7745 (N_7745,N_4611,N_5414);
nor U7746 (N_7746,N_5761,N_5007);
nor U7747 (N_7747,N_5208,N_4455);
nor U7748 (N_7748,N_5598,N_4969);
nand U7749 (N_7749,N_4834,N_5230);
and U7750 (N_7750,N_4617,N_5781);
nor U7751 (N_7751,N_4227,N_5353);
or U7752 (N_7752,N_5414,N_4369);
and U7753 (N_7753,N_4868,N_4885);
or U7754 (N_7754,N_5727,N_4725);
and U7755 (N_7755,N_4994,N_5691);
nor U7756 (N_7756,N_4225,N_4554);
and U7757 (N_7757,N_4663,N_4738);
nand U7758 (N_7758,N_4638,N_4405);
or U7759 (N_7759,N_4119,N_4731);
or U7760 (N_7760,N_5213,N_4564);
and U7761 (N_7761,N_5481,N_5671);
or U7762 (N_7762,N_4841,N_5715);
nand U7763 (N_7763,N_4882,N_4595);
and U7764 (N_7764,N_5984,N_5146);
or U7765 (N_7765,N_4869,N_5357);
nor U7766 (N_7766,N_5430,N_4118);
or U7767 (N_7767,N_4404,N_4594);
nor U7768 (N_7768,N_4795,N_4612);
or U7769 (N_7769,N_5521,N_4812);
nor U7770 (N_7770,N_5179,N_5182);
nand U7771 (N_7771,N_4068,N_4485);
nor U7772 (N_7772,N_4018,N_5809);
or U7773 (N_7773,N_5635,N_5237);
or U7774 (N_7774,N_4498,N_4959);
and U7775 (N_7775,N_5490,N_5752);
and U7776 (N_7776,N_5491,N_4485);
and U7777 (N_7777,N_5298,N_5996);
nor U7778 (N_7778,N_4849,N_4046);
nand U7779 (N_7779,N_4941,N_5151);
nor U7780 (N_7780,N_5939,N_5335);
nor U7781 (N_7781,N_5983,N_5637);
nor U7782 (N_7782,N_4979,N_5729);
nand U7783 (N_7783,N_5141,N_5927);
and U7784 (N_7784,N_5723,N_5149);
or U7785 (N_7785,N_5751,N_5658);
and U7786 (N_7786,N_4582,N_4558);
nor U7787 (N_7787,N_5211,N_4865);
or U7788 (N_7788,N_4522,N_5750);
or U7789 (N_7789,N_5117,N_4467);
xnor U7790 (N_7790,N_4447,N_5343);
and U7791 (N_7791,N_5927,N_4746);
nand U7792 (N_7792,N_4934,N_5995);
nor U7793 (N_7793,N_5638,N_5159);
nand U7794 (N_7794,N_5371,N_4205);
nor U7795 (N_7795,N_4555,N_4706);
or U7796 (N_7796,N_4077,N_5334);
nor U7797 (N_7797,N_5944,N_4958);
and U7798 (N_7798,N_4808,N_4799);
or U7799 (N_7799,N_4020,N_4279);
nor U7800 (N_7800,N_5110,N_5142);
and U7801 (N_7801,N_4332,N_5579);
nand U7802 (N_7802,N_4120,N_4668);
or U7803 (N_7803,N_5103,N_4414);
or U7804 (N_7804,N_5374,N_4792);
and U7805 (N_7805,N_4058,N_4117);
and U7806 (N_7806,N_4908,N_5178);
nand U7807 (N_7807,N_5855,N_5283);
nor U7808 (N_7808,N_4420,N_4574);
nor U7809 (N_7809,N_5264,N_4193);
nand U7810 (N_7810,N_4210,N_5461);
and U7811 (N_7811,N_4352,N_5828);
and U7812 (N_7812,N_5405,N_5192);
and U7813 (N_7813,N_4884,N_5132);
or U7814 (N_7814,N_4921,N_5938);
nor U7815 (N_7815,N_4628,N_4522);
and U7816 (N_7816,N_5964,N_4205);
and U7817 (N_7817,N_4619,N_4208);
or U7818 (N_7818,N_4418,N_5944);
nand U7819 (N_7819,N_4241,N_5802);
nand U7820 (N_7820,N_5384,N_5633);
and U7821 (N_7821,N_5002,N_5084);
xor U7822 (N_7822,N_4252,N_4480);
or U7823 (N_7823,N_5406,N_4394);
nand U7824 (N_7824,N_4570,N_4191);
and U7825 (N_7825,N_4646,N_5488);
and U7826 (N_7826,N_5867,N_4461);
or U7827 (N_7827,N_5045,N_4344);
and U7828 (N_7828,N_5431,N_4953);
and U7829 (N_7829,N_5210,N_5637);
nor U7830 (N_7830,N_4147,N_4269);
nand U7831 (N_7831,N_5741,N_4213);
nor U7832 (N_7832,N_4545,N_4820);
nand U7833 (N_7833,N_4635,N_5782);
xor U7834 (N_7834,N_5499,N_4999);
or U7835 (N_7835,N_4635,N_4387);
nand U7836 (N_7836,N_4970,N_5547);
nand U7837 (N_7837,N_5576,N_4008);
nor U7838 (N_7838,N_5680,N_5920);
or U7839 (N_7839,N_4148,N_5721);
nor U7840 (N_7840,N_5441,N_4157);
and U7841 (N_7841,N_4092,N_4714);
nor U7842 (N_7842,N_5826,N_5253);
nand U7843 (N_7843,N_4809,N_5532);
nor U7844 (N_7844,N_4122,N_4117);
nor U7845 (N_7845,N_4376,N_5892);
nand U7846 (N_7846,N_5864,N_4938);
nand U7847 (N_7847,N_5362,N_5843);
and U7848 (N_7848,N_5701,N_5411);
nor U7849 (N_7849,N_5944,N_5458);
nor U7850 (N_7850,N_5260,N_4222);
nor U7851 (N_7851,N_5945,N_4080);
and U7852 (N_7852,N_5457,N_4561);
and U7853 (N_7853,N_4990,N_5965);
and U7854 (N_7854,N_4678,N_5565);
nand U7855 (N_7855,N_4417,N_5766);
and U7856 (N_7856,N_4086,N_5408);
or U7857 (N_7857,N_5962,N_5193);
and U7858 (N_7858,N_4068,N_4924);
and U7859 (N_7859,N_5594,N_5794);
nor U7860 (N_7860,N_4239,N_4991);
or U7861 (N_7861,N_4155,N_5094);
and U7862 (N_7862,N_4041,N_4599);
nand U7863 (N_7863,N_5785,N_4416);
or U7864 (N_7864,N_4985,N_4609);
nand U7865 (N_7865,N_4011,N_5455);
nor U7866 (N_7866,N_5132,N_4059);
nand U7867 (N_7867,N_4767,N_4082);
or U7868 (N_7868,N_5073,N_4885);
nor U7869 (N_7869,N_5349,N_4534);
or U7870 (N_7870,N_5933,N_4755);
and U7871 (N_7871,N_4771,N_5293);
nor U7872 (N_7872,N_5346,N_4228);
nor U7873 (N_7873,N_4163,N_4389);
nand U7874 (N_7874,N_5402,N_4451);
nor U7875 (N_7875,N_5282,N_4135);
or U7876 (N_7876,N_4126,N_5125);
nor U7877 (N_7877,N_4738,N_5040);
nor U7878 (N_7878,N_4216,N_5486);
nand U7879 (N_7879,N_4681,N_5121);
or U7880 (N_7880,N_5841,N_5851);
and U7881 (N_7881,N_4487,N_5386);
nor U7882 (N_7882,N_5502,N_5914);
and U7883 (N_7883,N_5737,N_4215);
nor U7884 (N_7884,N_4739,N_5286);
and U7885 (N_7885,N_4749,N_4332);
nand U7886 (N_7886,N_4522,N_4979);
nor U7887 (N_7887,N_5702,N_4559);
and U7888 (N_7888,N_5081,N_4761);
or U7889 (N_7889,N_4544,N_5874);
and U7890 (N_7890,N_5843,N_4684);
and U7891 (N_7891,N_4002,N_5456);
nor U7892 (N_7892,N_5511,N_4283);
nand U7893 (N_7893,N_4120,N_4789);
or U7894 (N_7894,N_4286,N_4543);
nor U7895 (N_7895,N_4029,N_4247);
nor U7896 (N_7896,N_4067,N_5818);
or U7897 (N_7897,N_4122,N_5967);
nand U7898 (N_7898,N_4621,N_5084);
or U7899 (N_7899,N_4243,N_4483);
and U7900 (N_7900,N_5127,N_5386);
or U7901 (N_7901,N_4202,N_4227);
nand U7902 (N_7902,N_4116,N_4935);
or U7903 (N_7903,N_4579,N_4947);
or U7904 (N_7904,N_5410,N_5901);
nor U7905 (N_7905,N_5376,N_5540);
or U7906 (N_7906,N_4807,N_4551);
and U7907 (N_7907,N_5820,N_5752);
nor U7908 (N_7908,N_5809,N_4110);
and U7909 (N_7909,N_5601,N_5874);
and U7910 (N_7910,N_4121,N_5450);
and U7911 (N_7911,N_4209,N_4205);
nor U7912 (N_7912,N_5779,N_5224);
nand U7913 (N_7913,N_4614,N_4365);
nand U7914 (N_7914,N_4169,N_5519);
and U7915 (N_7915,N_4983,N_4467);
nand U7916 (N_7916,N_5691,N_5277);
and U7917 (N_7917,N_5536,N_5747);
nand U7918 (N_7918,N_4344,N_4842);
or U7919 (N_7919,N_5542,N_4271);
nor U7920 (N_7920,N_5957,N_5390);
nor U7921 (N_7921,N_5326,N_4515);
or U7922 (N_7922,N_4488,N_5215);
and U7923 (N_7923,N_5419,N_5729);
nand U7924 (N_7924,N_5233,N_4001);
nand U7925 (N_7925,N_4249,N_4552);
nor U7926 (N_7926,N_5182,N_4742);
nor U7927 (N_7927,N_4462,N_5349);
nand U7928 (N_7928,N_4975,N_5222);
nor U7929 (N_7929,N_5985,N_4950);
nor U7930 (N_7930,N_4401,N_5750);
or U7931 (N_7931,N_4185,N_4485);
nor U7932 (N_7932,N_4156,N_5127);
nor U7933 (N_7933,N_4147,N_5305);
and U7934 (N_7934,N_5030,N_5632);
or U7935 (N_7935,N_4617,N_4612);
nand U7936 (N_7936,N_5810,N_4813);
nor U7937 (N_7937,N_5187,N_4735);
or U7938 (N_7938,N_4429,N_4370);
and U7939 (N_7939,N_4293,N_5000);
and U7940 (N_7940,N_4545,N_4745);
and U7941 (N_7941,N_4863,N_4790);
and U7942 (N_7942,N_4851,N_4481);
nand U7943 (N_7943,N_5105,N_4549);
or U7944 (N_7944,N_5087,N_4190);
nor U7945 (N_7945,N_4246,N_4005);
and U7946 (N_7946,N_5596,N_5265);
or U7947 (N_7947,N_4439,N_4859);
or U7948 (N_7948,N_4451,N_4853);
nor U7949 (N_7949,N_5852,N_4274);
or U7950 (N_7950,N_5043,N_4926);
nand U7951 (N_7951,N_5503,N_5959);
nand U7952 (N_7952,N_4487,N_4810);
nor U7953 (N_7953,N_5027,N_4471);
and U7954 (N_7954,N_5735,N_4010);
or U7955 (N_7955,N_5025,N_5879);
nand U7956 (N_7956,N_4025,N_5463);
nand U7957 (N_7957,N_4177,N_4633);
nand U7958 (N_7958,N_4961,N_4385);
or U7959 (N_7959,N_5080,N_5008);
and U7960 (N_7960,N_4645,N_4094);
nand U7961 (N_7961,N_4700,N_5025);
nand U7962 (N_7962,N_4931,N_4816);
and U7963 (N_7963,N_5809,N_5921);
and U7964 (N_7964,N_4659,N_4241);
nand U7965 (N_7965,N_4551,N_4358);
and U7966 (N_7966,N_4910,N_4063);
nand U7967 (N_7967,N_5561,N_5785);
xor U7968 (N_7968,N_4786,N_4021);
and U7969 (N_7969,N_5219,N_4182);
nand U7970 (N_7970,N_4539,N_5358);
nand U7971 (N_7971,N_5687,N_5737);
and U7972 (N_7972,N_4581,N_5578);
or U7973 (N_7973,N_5060,N_5473);
nand U7974 (N_7974,N_5728,N_5146);
nor U7975 (N_7975,N_4562,N_4405);
and U7976 (N_7976,N_5921,N_5917);
nand U7977 (N_7977,N_5582,N_5680);
or U7978 (N_7978,N_4638,N_4043);
and U7979 (N_7979,N_5228,N_4863);
xnor U7980 (N_7980,N_5103,N_5549);
nor U7981 (N_7981,N_4341,N_5566);
or U7982 (N_7982,N_4779,N_4962);
nor U7983 (N_7983,N_4002,N_4166);
or U7984 (N_7984,N_4913,N_5265);
or U7985 (N_7985,N_4576,N_5444);
nor U7986 (N_7986,N_5597,N_4396);
nor U7987 (N_7987,N_4742,N_4351);
or U7988 (N_7988,N_4731,N_5976);
nor U7989 (N_7989,N_5858,N_5083);
or U7990 (N_7990,N_4591,N_5867);
or U7991 (N_7991,N_4417,N_4002);
nand U7992 (N_7992,N_4809,N_5719);
xnor U7993 (N_7993,N_5154,N_4949);
nand U7994 (N_7994,N_5185,N_5081);
or U7995 (N_7995,N_4315,N_5316);
nor U7996 (N_7996,N_5483,N_4543);
or U7997 (N_7997,N_5405,N_5689);
nor U7998 (N_7998,N_5864,N_5390);
nand U7999 (N_7999,N_4605,N_5507);
nand U8000 (N_8000,N_6446,N_7123);
nand U8001 (N_8001,N_6548,N_7110);
or U8002 (N_8002,N_7332,N_7209);
or U8003 (N_8003,N_7634,N_7826);
and U8004 (N_8004,N_7410,N_7360);
and U8005 (N_8005,N_7927,N_7248);
nor U8006 (N_8006,N_6623,N_7664);
nand U8007 (N_8007,N_6852,N_7379);
nor U8008 (N_8008,N_6785,N_7338);
or U8009 (N_8009,N_7330,N_7294);
nand U8010 (N_8010,N_7255,N_7496);
or U8011 (N_8011,N_7234,N_6168);
nor U8012 (N_8012,N_7336,N_6713);
or U8013 (N_8013,N_6604,N_6320);
nand U8014 (N_8014,N_7731,N_6230);
nor U8015 (N_8015,N_6349,N_7484);
and U8016 (N_8016,N_7468,N_6676);
nor U8017 (N_8017,N_6626,N_6301);
nand U8018 (N_8018,N_7708,N_6120);
and U8019 (N_8019,N_7710,N_6053);
nand U8020 (N_8020,N_7241,N_7808);
nor U8021 (N_8021,N_6654,N_7010);
and U8022 (N_8022,N_6355,N_7450);
nor U8023 (N_8023,N_7992,N_7632);
or U8024 (N_8024,N_6140,N_7202);
nand U8025 (N_8025,N_6228,N_7122);
and U8026 (N_8026,N_7852,N_6402);
and U8027 (N_8027,N_7188,N_7836);
or U8028 (N_8028,N_6924,N_7069);
or U8029 (N_8029,N_6501,N_6240);
nand U8030 (N_8030,N_7888,N_7427);
nand U8031 (N_8031,N_7896,N_7617);
nor U8032 (N_8032,N_6507,N_7506);
nand U8033 (N_8033,N_7637,N_6559);
nand U8034 (N_8034,N_6553,N_7872);
nor U8035 (N_8035,N_7090,N_7426);
or U8036 (N_8036,N_6717,N_7325);
nor U8037 (N_8037,N_7959,N_7044);
or U8038 (N_8038,N_7551,N_7193);
nor U8039 (N_8039,N_6188,N_6844);
and U8040 (N_8040,N_6211,N_6768);
nand U8041 (N_8041,N_6444,N_6272);
nand U8042 (N_8042,N_7037,N_7579);
nand U8043 (N_8043,N_7622,N_7062);
and U8044 (N_8044,N_6975,N_7536);
nand U8045 (N_8045,N_7507,N_7340);
nand U8046 (N_8046,N_6739,N_6652);
nand U8047 (N_8047,N_6024,N_7827);
nand U8048 (N_8048,N_7096,N_7750);
nor U8049 (N_8049,N_7543,N_7635);
nor U8050 (N_8050,N_6586,N_6085);
or U8051 (N_8051,N_7077,N_6822);
nand U8052 (N_8052,N_7985,N_6389);
nand U8053 (N_8053,N_7965,N_7283);
nand U8054 (N_8054,N_6690,N_6712);
or U8055 (N_8055,N_6260,N_7716);
nor U8056 (N_8056,N_7799,N_6049);
and U8057 (N_8057,N_7412,N_7464);
nor U8058 (N_8058,N_7855,N_6394);
or U8059 (N_8059,N_6421,N_7017);
nor U8060 (N_8060,N_6890,N_7995);
nor U8061 (N_8061,N_7859,N_7968);
or U8062 (N_8062,N_6647,N_7016);
nand U8063 (N_8063,N_6476,N_6467);
nand U8064 (N_8064,N_7268,N_6487);
or U8065 (N_8065,N_7133,N_7073);
nand U8066 (N_8066,N_7386,N_7803);
nand U8067 (N_8067,N_7944,N_7973);
nand U8068 (N_8068,N_6640,N_6758);
and U8069 (N_8069,N_7366,N_6418);
nor U8070 (N_8070,N_6895,N_6527);
nand U8071 (N_8071,N_6959,N_7436);
and U8072 (N_8072,N_7142,N_7671);
nor U8073 (N_8073,N_7215,N_7478);
nand U8074 (N_8074,N_6919,N_6189);
or U8075 (N_8075,N_7726,N_7686);
or U8076 (N_8076,N_6773,N_7790);
nor U8077 (N_8077,N_7626,N_7175);
and U8078 (N_8078,N_7287,N_6082);
xnor U8079 (N_8079,N_6458,N_7694);
nand U8080 (N_8080,N_7982,N_6019);
nor U8081 (N_8081,N_7994,N_6858);
nor U8082 (N_8082,N_7176,N_6535);
and U8083 (N_8083,N_6839,N_7627);
and U8084 (N_8084,N_6315,N_6601);
nand U8085 (N_8085,N_7546,N_6457);
and U8086 (N_8086,N_7805,N_6770);
nor U8087 (N_8087,N_6625,N_6245);
nor U8088 (N_8088,N_6000,N_7333);
nand U8089 (N_8089,N_6552,N_7561);
nor U8090 (N_8090,N_6789,N_6144);
nand U8091 (N_8091,N_6434,N_7920);
and U8092 (N_8092,N_7935,N_6371);
nor U8093 (N_8093,N_7831,N_6563);
nand U8094 (N_8094,N_6236,N_6400);
nand U8095 (N_8095,N_6877,N_7232);
nand U8096 (N_8096,N_7095,N_7934);
xnor U8097 (N_8097,N_6414,N_7440);
and U8098 (N_8098,N_7754,N_7302);
nor U8099 (N_8099,N_6622,N_6021);
nor U8100 (N_8100,N_7993,N_6513);
and U8101 (N_8101,N_6738,N_7243);
and U8102 (N_8102,N_7448,N_7608);
nor U8103 (N_8103,N_6939,N_7857);
and U8104 (N_8104,N_6727,N_7313);
nor U8105 (N_8105,N_7022,N_7873);
nand U8106 (N_8106,N_7199,N_6537);
and U8107 (N_8107,N_6607,N_6209);
nand U8108 (N_8108,N_7931,N_6533);
and U8109 (N_8109,N_6169,N_6463);
nor U8110 (N_8110,N_7030,N_7134);
or U8111 (N_8111,N_7988,N_6792);
or U8112 (N_8112,N_6433,N_7348);
nor U8113 (N_8113,N_7769,N_6945);
or U8114 (N_8114,N_7548,N_7054);
and U8115 (N_8115,N_7117,N_7876);
nand U8116 (N_8116,N_6908,N_7963);
or U8117 (N_8117,N_6608,N_6088);
or U8118 (N_8118,N_6733,N_7584);
nand U8119 (N_8119,N_7497,N_7401);
nand U8120 (N_8120,N_7958,N_6497);
nor U8121 (N_8121,N_7829,N_6590);
or U8122 (N_8122,N_7862,N_6706);
nand U8123 (N_8123,N_6749,N_7774);
and U8124 (N_8124,N_6688,N_6368);
or U8125 (N_8125,N_6341,N_7303);
or U8126 (N_8126,N_7717,N_7703);
nor U8127 (N_8127,N_7508,N_6461);
and U8128 (N_8128,N_6139,N_7361);
nand U8129 (N_8129,N_6160,N_6635);
and U8130 (N_8130,N_7770,N_6293);
or U8131 (N_8131,N_7793,N_7670);
nand U8132 (N_8132,N_7537,N_7003);
nor U8133 (N_8133,N_7527,N_6557);
nand U8134 (N_8134,N_6011,N_6041);
or U8135 (N_8135,N_7056,N_7319);
nor U8136 (N_8136,N_6947,N_6070);
or U8137 (N_8137,N_7388,N_6427);
or U8138 (N_8138,N_7522,N_6828);
nor U8139 (N_8139,N_6439,N_7495);
and U8140 (N_8140,N_7221,N_7633);
or U8141 (N_8141,N_7345,N_7048);
nor U8142 (N_8142,N_7893,N_6985);
nand U8143 (N_8143,N_7154,N_7012);
nand U8144 (N_8144,N_6353,N_6473);
nand U8145 (N_8145,N_7911,N_6202);
or U8146 (N_8146,N_7130,N_7595);
and U8147 (N_8147,N_7918,N_6281);
and U8148 (N_8148,N_7699,N_6724);
or U8149 (N_8149,N_7639,N_7374);
nand U8150 (N_8150,N_6916,N_7141);
nand U8151 (N_8151,N_6014,N_6982);
nand U8152 (N_8152,N_6835,N_6996);
nor U8153 (N_8153,N_6471,N_7079);
or U8154 (N_8154,N_6883,N_7138);
and U8155 (N_8155,N_6171,N_7515);
and U8156 (N_8156,N_6380,N_6905);
nand U8157 (N_8157,N_6386,N_7192);
or U8158 (N_8158,N_7800,N_6767);
and U8159 (N_8159,N_6932,N_7493);
nand U8160 (N_8160,N_7815,N_7779);
and U8161 (N_8161,N_6793,N_7155);
nand U8162 (N_8162,N_6269,N_7324);
or U8163 (N_8163,N_7660,N_7086);
or U8164 (N_8164,N_7885,N_7528);
and U8165 (N_8165,N_6752,N_7292);
and U8166 (N_8166,N_6665,N_6574);
or U8167 (N_8167,N_6798,N_7083);
and U8168 (N_8168,N_7165,N_7486);
nor U8169 (N_8169,N_7001,N_6498);
nand U8170 (N_8170,N_6783,N_7736);
nand U8171 (N_8171,N_6338,N_6317);
and U8172 (N_8172,N_7572,N_6613);
or U8173 (N_8173,N_7682,N_7359);
or U8174 (N_8174,N_7169,N_7631);
nor U8175 (N_8175,N_6016,N_7843);
and U8176 (N_8176,N_6063,N_7033);
and U8177 (N_8177,N_7877,N_7695);
or U8178 (N_8178,N_6263,N_6830);
or U8179 (N_8179,N_6600,N_6555);
nor U8180 (N_8180,N_6304,N_7005);
nor U8181 (N_8181,N_6186,N_6725);
nor U8182 (N_8182,N_6915,N_6278);
nand U8183 (N_8183,N_6728,N_7414);
or U8184 (N_8184,N_6478,N_6679);
nand U8185 (N_8185,N_7351,N_7317);
nand U8186 (N_8186,N_7451,N_7197);
nor U8187 (N_8187,N_6350,N_7700);
nor U8188 (N_8188,N_6755,N_6510);
nand U8189 (N_8189,N_6210,N_7163);
or U8190 (N_8190,N_7422,N_7218);
nand U8191 (N_8191,N_6261,N_7646);
nor U8192 (N_8192,N_7838,N_6382);
nor U8193 (N_8193,N_7137,N_6565);
or U8194 (N_8194,N_7534,N_6383);
or U8195 (N_8195,N_6333,N_7740);
nor U8196 (N_8196,N_6403,N_6157);
and U8197 (N_8197,N_6373,N_6115);
and U8198 (N_8198,N_7737,N_6656);
and U8199 (N_8199,N_6208,N_6855);
or U8200 (N_8200,N_6201,N_6080);
and U8201 (N_8201,N_7288,N_6631);
nor U8202 (N_8202,N_6732,N_6106);
nor U8203 (N_8203,N_7198,N_6399);
nor U8204 (N_8204,N_7061,N_7544);
nor U8205 (N_8205,N_7747,N_7961);
nand U8206 (N_8206,N_6076,N_7156);
nor U8207 (N_8207,N_6370,N_7798);
and U8208 (N_8208,N_7604,N_7773);
and U8209 (N_8209,N_6824,N_6584);
and U8210 (N_8210,N_7880,N_7323);
or U8211 (N_8211,N_6853,N_7078);
nand U8212 (N_8212,N_7066,N_7605);
nand U8213 (N_8213,N_6112,N_6721);
or U8214 (N_8214,N_6992,N_6215);
nor U8215 (N_8215,N_7214,N_6187);
nand U8216 (N_8216,N_6372,N_6432);
nor U8217 (N_8217,N_7295,N_6413);
and U8218 (N_8218,N_7228,N_6454);
and U8219 (N_8219,N_6522,N_7794);
nand U8220 (N_8220,N_7084,N_6314);
nor U8221 (N_8221,N_6166,N_6815);
nand U8222 (N_8222,N_6217,N_6582);
nand U8223 (N_8223,N_6838,N_7190);
or U8224 (N_8224,N_6954,N_6766);
or U8225 (N_8225,N_7203,N_6920);
nor U8226 (N_8226,N_6764,N_7185);
nor U8227 (N_8227,N_7607,N_7247);
or U8228 (N_8228,N_7786,N_6084);
and U8229 (N_8229,N_6790,N_7310);
nor U8230 (N_8230,N_7580,N_7820);
or U8231 (N_8231,N_6784,N_6391);
nand U8232 (N_8232,N_6328,N_7854);
nand U8233 (N_8233,N_6401,N_6643);
nor U8234 (N_8234,N_6059,N_7170);
and U8235 (N_8235,N_6089,N_6181);
nor U8236 (N_8236,N_6807,N_6980);
nor U8237 (N_8237,N_6788,N_6193);
or U8238 (N_8238,N_6816,N_6662);
or U8239 (N_8239,N_7870,N_6312);
or U8240 (N_8240,N_7306,N_6158);
nand U8241 (N_8241,N_6927,N_6868);
and U8242 (N_8242,N_6462,N_6722);
nand U8243 (N_8243,N_6252,N_7796);
or U8244 (N_8244,N_6067,N_6221);
nor U8245 (N_8245,N_7712,N_6957);
and U8246 (N_8246,N_6289,N_7613);
or U8247 (N_8247,N_7269,N_6499);
and U8248 (N_8248,N_6012,N_7264);
nor U8249 (N_8249,N_7246,N_7356);
nor U8250 (N_8250,N_7969,N_7498);
nand U8251 (N_8251,N_7733,N_7739);
and U8252 (N_8252,N_7656,N_6031);
nor U8253 (N_8253,N_6633,N_6197);
nor U8254 (N_8254,N_6036,N_6104);
nor U8255 (N_8255,N_7430,N_7471);
nand U8256 (N_8256,N_7952,N_7948);
or U8257 (N_8257,N_7727,N_6406);
nand U8258 (N_8258,N_7663,N_7477);
nand U8259 (N_8259,N_7600,N_6695);
nor U8260 (N_8260,N_6040,N_7897);
and U8261 (N_8261,N_7625,N_7178);
nor U8262 (N_8262,N_6431,N_7589);
nor U8263 (N_8263,N_7363,N_7970);
or U8264 (N_8264,N_7933,N_6464);
or U8265 (N_8265,N_6701,N_7026);
and U8266 (N_8266,N_7512,N_7676);
or U8267 (N_8267,N_7819,N_6101);
nor U8268 (N_8268,N_6550,N_6359);
nor U8269 (N_8269,N_6829,N_6337);
and U8270 (N_8270,N_6532,N_7575);
nand U8271 (N_8271,N_6653,N_6025);
nand U8272 (N_8272,N_7305,N_7402);
nand U8273 (N_8273,N_7946,N_7435);
nor U8274 (N_8274,N_6365,N_7068);
nand U8275 (N_8275,N_7641,N_6943);
nand U8276 (N_8276,N_6229,N_6650);
and U8277 (N_8277,N_7749,N_6762);
nor U8278 (N_8278,N_6010,N_7370);
and U8279 (N_8279,N_6700,N_6265);
and U8280 (N_8280,N_7023,N_7977);
or U8281 (N_8281,N_6592,N_7258);
nor U8282 (N_8282,N_6319,N_6672);
nand U8283 (N_8283,N_6154,N_6897);
nor U8284 (N_8284,N_6955,N_7494);
nand U8285 (N_8285,N_7709,N_7687);
or U8286 (N_8286,N_6285,N_7669);
nand U8287 (N_8287,N_6124,N_7902);
and U8288 (N_8288,N_7906,N_6405);
and U8289 (N_8289,N_7164,N_7092);
nand U8290 (N_8290,N_7021,N_7955);
or U8291 (N_8291,N_6857,N_7148);
and U8292 (N_8292,N_7167,N_6671);
nor U8293 (N_8293,N_7334,N_7168);
nand U8294 (N_8294,N_6743,N_6420);
or U8295 (N_8295,N_6558,N_6133);
or U8296 (N_8296,N_7581,N_7525);
and U8297 (N_8297,N_7114,N_6551);
and U8298 (N_8298,N_7636,N_7446);
or U8299 (N_8299,N_7504,N_7685);
nor U8300 (N_8300,N_6356,N_6912);
nand U8301 (N_8301,N_6944,N_6212);
and U8302 (N_8302,N_6375,N_6628);
or U8303 (N_8303,N_7009,N_7256);
and U8304 (N_8304,N_6846,N_7213);
nand U8305 (N_8305,N_6691,N_6914);
nor U8306 (N_8306,N_7301,N_7445);
and U8307 (N_8307,N_7681,N_6437);
nor U8308 (N_8308,N_6184,N_7943);
and U8309 (N_8309,N_7704,N_7488);
nand U8310 (N_8310,N_6925,N_7316);
and U8311 (N_8311,N_7298,N_7368);
nor U8312 (N_8312,N_7889,N_6495);
nor U8313 (N_8313,N_7652,N_7623);
and U8314 (N_8314,N_6668,N_7558);
or U8315 (N_8315,N_7075,N_6449);
and U8316 (N_8316,N_6595,N_7592);
and U8317 (N_8317,N_7153,N_6251);
nand U8318 (N_8318,N_6504,N_6342);
nand U8319 (N_8319,N_7449,N_6569);
and U8320 (N_8320,N_6587,N_7385);
nand U8321 (N_8321,N_7491,N_7204);
and U8322 (N_8322,N_6491,N_7586);
or U8323 (N_8323,N_7742,N_6456);
nand U8324 (N_8324,N_7150,N_6322);
and U8325 (N_8325,N_6493,N_7028);
and U8326 (N_8326,N_7706,N_7014);
nand U8327 (N_8327,N_7285,N_6442);
nand U8328 (N_8328,N_6893,N_6620);
or U8329 (N_8329,N_6207,N_6441);
nor U8330 (N_8330,N_6506,N_7915);
nor U8331 (N_8331,N_7470,N_7485);
and U8332 (N_8332,N_6159,N_7015);
and U8333 (N_8333,N_7908,N_7618);
or U8334 (N_8334,N_7042,N_6074);
and U8335 (N_8335,N_6429,N_7398);
and U8336 (N_8336,N_7650,N_6440);
nand U8337 (N_8337,N_7904,N_6981);
nand U8338 (N_8338,N_6681,N_7252);
nand U8339 (N_8339,N_7104,N_7503);
nor U8340 (N_8340,N_6489,N_6685);
or U8341 (N_8341,N_6316,N_6630);
and U8342 (N_8342,N_6071,N_7335);
nand U8343 (N_8343,N_7487,N_7738);
or U8344 (N_8344,N_7901,N_7281);
nor U8345 (N_8345,N_6697,N_7802);
and U8346 (N_8346,N_6863,N_7018);
and U8347 (N_8347,N_6572,N_7538);
or U8348 (N_8348,N_6664,N_6997);
and U8349 (N_8349,N_7828,N_6205);
or U8350 (N_8350,N_6987,N_6416);
or U8351 (N_8351,N_6198,N_7382);
and U8352 (N_8352,N_7049,N_6398);
or U8353 (N_8353,N_6292,N_6745);
or U8354 (N_8354,N_6942,N_7147);
nand U8355 (N_8355,N_6488,N_7437);
and U8356 (N_8356,N_7384,N_7320);
nor U8357 (N_8357,N_7358,N_6938);
nand U8358 (N_8358,N_6984,N_7299);
or U8359 (N_8359,N_7936,N_6087);
and U8360 (N_8360,N_6117,N_7986);
and U8361 (N_8361,N_7611,N_6347);
nor U8362 (N_8362,N_7787,N_7315);
nand U8363 (N_8363,N_7980,N_6183);
nor U8364 (N_8364,N_7705,N_7217);
nor U8365 (N_8365,N_7041,N_6095);
nor U8366 (N_8366,N_6810,N_6485);
and U8367 (N_8367,N_6109,N_7046);
and U8368 (N_8368,N_6837,N_6191);
nand U8369 (N_8369,N_7883,N_7780);
or U8370 (N_8370,N_6042,N_7628);
or U8371 (N_8371,N_6564,N_7296);
and U8372 (N_8372,N_6926,N_6377);
nand U8373 (N_8373,N_7085,N_6075);
and U8374 (N_8374,N_6177,N_7851);
nor U8375 (N_8375,N_6744,N_6026);
nand U8376 (N_8376,N_6268,N_6541);
or U8377 (N_8377,N_6151,N_7957);
nand U8378 (N_8378,N_7945,N_6588);
and U8379 (N_8379,N_6906,N_7131);
or U8380 (N_8380,N_7250,N_7289);
nand U8381 (N_8381,N_7677,N_7173);
and U8382 (N_8382,N_6936,N_7443);
nand U8383 (N_8383,N_7542,N_7020);
nand U8384 (N_8384,N_6161,N_7499);
or U8385 (N_8385,N_7554,N_7718);
nand U8386 (N_8386,N_6083,N_6703);
nand U8387 (N_8387,N_7643,N_6450);
nand U8388 (N_8388,N_6203,N_6978);
and U8389 (N_8389,N_7757,N_6616);
and U8390 (N_8390,N_7956,N_6866);
nor U8391 (N_8391,N_7954,N_6256);
nand U8392 (N_8392,N_7984,N_6683);
nand U8393 (N_8393,N_6156,N_6466);
or U8394 (N_8394,N_7849,N_7523);
nand U8395 (N_8395,N_6332,N_6892);
nor U8396 (N_8396,N_6173,N_7035);
nand U8397 (N_8397,N_7112,N_7050);
or U8398 (N_8398,N_7040,N_7569);
and U8399 (N_8399,N_6060,N_7121);
and U8400 (N_8400,N_7601,N_7549);
nor U8401 (N_8401,N_7689,N_6424);
nand U8402 (N_8402,N_7594,N_7300);
or U8403 (N_8403,N_6052,N_6940);
or U8404 (N_8404,N_7365,N_7032);
nor U8405 (N_8405,N_7932,N_7233);
or U8406 (N_8406,N_7157,N_7051);
or U8407 (N_8407,N_7352,N_6220);
and U8408 (N_8408,N_6583,N_6481);
nor U8409 (N_8409,N_6967,N_7866);
nor U8410 (N_8410,N_7762,N_7698);
or U8411 (N_8411,N_7070,N_7951);
and U8412 (N_8412,N_7830,N_7093);
nand U8413 (N_8413,N_6232,N_6775);
nor U8414 (N_8414,N_6632,N_6748);
nand U8415 (N_8415,N_6966,N_6518);
or U8416 (N_8416,N_6663,N_7417);
nand U8417 (N_8417,N_6577,N_6093);
nor U8418 (N_8418,N_6058,N_6061);
nand U8419 (N_8419,N_7433,N_6235);
and U8420 (N_8420,N_7272,N_6266);
nor U8421 (N_8421,N_6288,N_6561);
xnor U8422 (N_8422,N_6192,N_7349);
and U8423 (N_8423,N_6619,N_6667);
nor U8424 (N_8424,N_6470,N_7219);
nand U8425 (N_8425,N_7166,N_7612);
nor U8426 (N_8426,N_6327,N_6308);
nor U8427 (N_8427,N_6958,N_6410);
or U8428 (N_8428,N_6390,N_6219);
nand U8429 (N_8429,N_6834,N_7967);
nand U8430 (N_8430,N_7647,N_6425);
or U8431 (N_8431,N_6833,N_6545);
nor U8432 (N_8432,N_7072,N_6129);
or U8433 (N_8433,N_6477,N_7583);
or U8434 (N_8434,N_7439,N_7892);
nand U8435 (N_8435,N_7823,N_6995);
or U8436 (N_8436,N_7149,N_6296);
and U8437 (N_8437,N_7262,N_7875);
nand U8438 (N_8438,N_6249,N_6880);
nor U8439 (N_8439,N_6069,N_7128);
nand U8440 (N_8440,N_6199,N_7890);
or U8441 (N_8441,N_7690,N_7684);
or U8442 (N_8442,N_6763,N_7222);
or U8443 (N_8443,N_7413,N_7432);
or U8444 (N_8444,N_6702,N_6153);
and U8445 (N_8445,N_6731,N_7107);
or U8446 (N_8446,N_7778,N_6843);
and U8447 (N_8447,N_6149,N_7377);
and U8448 (N_8448,N_7720,N_7210);
and U8449 (N_8449,N_6262,N_6005);
nor U8450 (N_8450,N_7587,N_7242);
and U8451 (N_8451,N_6546,N_6796);
or U8452 (N_8452,N_7223,N_7251);
nand U8453 (N_8453,N_7059,N_7910);
and U8454 (N_8454,N_7949,N_7891);
nor U8455 (N_8455,N_7763,N_7545);
and U8456 (N_8456,N_7753,N_7314);
nor U8457 (N_8457,N_7597,N_7161);
nand U8458 (N_8458,N_7732,N_7614);
nor U8459 (N_8459,N_6962,N_6742);
and U8460 (N_8460,N_6689,N_6412);
nor U8461 (N_8461,N_7991,N_6132);
nor U8462 (N_8462,N_6436,N_6407);
nand U8463 (N_8463,N_7509,N_6801);
nand U8464 (N_8464,N_7566,N_7002);
nor U8465 (N_8465,N_7089,N_6605);
and U8466 (N_8466,N_7111,N_6960);
nand U8467 (N_8467,N_7758,N_7282);
nand U8468 (N_8468,N_7346,N_6544);
or U8469 (N_8469,N_7329,N_6970);
and U8470 (N_8470,N_7881,N_7620);
nand U8471 (N_8471,N_6264,N_7714);
nor U8472 (N_8472,N_6279,N_7972);
or U8473 (N_8473,N_7942,N_7856);
nand U8474 (N_8474,N_6043,N_7804);
and U8475 (N_8475,N_6769,N_6017);
or U8476 (N_8476,N_6331,N_7833);
nor U8477 (N_8477,N_6455,N_7372);
and U8478 (N_8478,N_7088,N_7781);
nand U8479 (N_8479,N_7362,N_6324);
or U8480 (N_8480,N_6649,N_6351);
and U8481 (N_8481,N_6879,N_6213);
or U8482 (N_8482,N_6358,N_7277);
nor U8483 (N_8483,N_6542,N_7118);
or U8484 (N_8484,N_6469,N_7521);
nor U8485 (N_8485,N_7013,N_6660);
nand U8486 (N_8486,N_7615,N_7730);
and U8487 (N_8487,N_6345,N_7886);
nor U8488 (N_8488,N_7469,N_6659);
and U8489 (N_8489,N_6699,N_7869);
and U8490 (N_8490,N_6718,N_7532);
nand U8491 (N_8491,N_7582,N_6873);
or U8492 (N_8492,N_7693,N_7816);
nor U8493 (N_8493,N_6517,N_6979);
and U8494 (N_8494,N_7841,N_7102);
and U8495 (N_8495,N_6735,N_6859);
nor U8496 (N_8496,N_6538,N_7999);
nor U8497 (N_8497,N_6512,N_7474);
or U8498 (N_8498,N_6986,N_6468);
nor U8499 (N_8499,N_7339,N_7159);
nand U8500 (N_8500,N_6539,N_7925);
or U8501 (N_8501,N_7903,N_7309);
and U8502 (N_8502,N_6170,N_6804);
nand U8503 (N_8503,N_7567,N_6490);
nand U8504 (N_8504,N_7539,N_7785);
and U8505 (N_8505,N_6524,N_7293);
or U8506 (N_8506,N_6057,N_6903);
and U8507 (N_8507,N_6831,N_7321);
nor U8508 (N_8508,N_7530,N_7179);
nor U8509 (N_8509,N_7394,N_7201);
or U8510 (N_8510,N_6854,N_6484);
and U8511 (N_8511,N_7236,N_6566);
nor U8512 (N_8512,N_7842,N_7113);
nand U8513 (N_8513,N_7513,N_7492);
and U8514 (N_8514,N_7053,N_6645);
nor U8515 (N_8515,N_6241,N_6677);
nand U8516 (N_8516,N_6795,N_7821);
and U8517 (N_8517,N_6684,N_7490);
or U8518 (N_8518,N_6127,N_6864);
nand U8519 (N_8519,N_6448,N_6870);
nand U8520 (N_8520,N_7297,N_6786);
nand U8521 (N_8521,N_6746,N_7074);
nor U8522 (N_8522,N_6802,N_7404);
nand U8523 (N_8523,N_6756,N_6806);
nor U8524 (N_8524,N_6282,N_7208);
and U8525 (N_8525,N_7206,N_7578);
or U8526 (N_8526,N_6185,N_6778);
nor U8527 (N_8527,N_7563,N_7375);
nand U8528 (N_8528,N_6030,N_6861);
or U8529 (N_8529,N_6573,N_7364);
nor U8530 (N_8530,N_6990,N_6675);
nand U8531 (N_8531,N_6765,N_6494);
and U8532 (N_8532,N_7189,N_6443);
or U8533 (N_8533,N_7744,N_6298);
and U8534 (N_8534,N_7171,N_6845);
nand U8535 (N_8535,N_7226,N_7678);
and U8536 (N_8536,N_6730,N_7752);
and U8537 (N_8537,N_7560,N_6921);
nor U8538 (N_8538,N_7280,N_7237);
and U8539 (N_8539,N_6847,N_6963);
nor U8540 (N_8540,N_6226,N_6385);
nor U8541 (N_8541,N_6658,N_6352);
and U8542 (N_8542,N_6163,N_7183);
nand U8543 (N_8543,N_7541,N_6318);
nor U8544 (N_8544,N_7265,N_6135);
and U8545 (N_8545,N_6387,N_6591);
nand U8546 (N_8546,N_6287,N_6255);
or U8547 (N_8547,N_6715,N_6362);
nand U8548 (N_8548,N_6842,N_7570);
and U8549 (N_8549,N_7143,N_6521);
or U8550 (N_8550,N_6611,N_6344);
nor U8551 (N_8551,N_7253,N_7279);
or U8552 (N_8552,N_6369,N_7884);
and U8553 (N_8553,N_7132,N_6378);
nor U8554 (N_8554,N_7200,N_7393);
nand U8555 (N_8555,N_6760,N_6710);
nand U8556 (N_8556,N_6445,N_7813);
nand U8557 (N_8557,N_7459,N_6409);
and U8558 (N_8558,N_6881,N_6239);
nor U8559 (N_8559,N_6593,N_7181);
nand U8560 (N_8560,N_7225,N_7395);
and U8561 (N_8561,N_7502,N_7034);
or U8562 (N_8562,N_7724,N_6624);
xnor U8563 (N_8563,N_7483,N_6634);
and U8564 (N_8564,N_6146,N_6502);
nor U8565 (N_8565,N_7576,N_7921);
and U8566 (N_8566,N_7501,N_7308);
nand U8567 (N_8567,N_6736,N_6346);
or U8568 (N_8568,N_6291,N_6651);
xor U8569 (N_8569,N_7761,N_6805);
nand U8570 (N_8570,N_6142,N_6460);
and U8571 (N_8571,N_7930,N_6354);
or U8572 (N_8572,N_7844,N_6267);
or U8573 (N_8573,N_7688,N_7659);
nor U8574 (N_8574,N_7928,N_6038);
and U8575 (N_8575,N_6780,N_6560);
and U8576 (N_8576,N_6361,N_7658);
nor U8577 (N_8577,N_6162,N_6617);
nand U8578 (N_8578,N_7397,N_7811);
and U8579 (N_8579,N_6180,N_6428);
nand U8580 (N_8580,N_6013,N_6747);
or U8581 (N_8581,N_6705,N_6008);
nor U8582 (N_8582,N_6422,N_7376);
and U8583 (N_8583,N_7619,N_7832);
nor U8584 (N_8584,N_7505,N_7254);
or U8585 (N_8585,N_7400,N_7467);
nor U8586 (N_8586,N_6761,N_6872);
and U8587 (N_8587,N_7853,N_6270);
or U8588 (N_8588,N_6003,N_7212);
or U8589 (N_8589,N_7116,N_7697);
nand U8590 (N_8590,N_7326,N_6172);
nor U8591 (N_8591,N_7568,N_6734);
nor U8592 (N_8592,N_7529,N_6134);
and U8593 (N_8593,N_6941,N_6430);
or U8594 (N_8594,N_6708,N_6379);
nor U8595 (N_8595,N_7644,N_7909);
and U8596 (N_8596,N_7249,N_7008);
nand U8597 (N_8597,N_6898,N_6274);
nand U8598 (N_8598,N_6817,N_7180);
or U8599 (N_8599,N_7602,N_6048);
nand U8600 (N_8600,N_6147,N_6964);
and U8601 (N_8601,N_6899,N_7460);
and U8602 (N_8602,N_7719,N_7692);
nand U8603 (N_8603,N_6143,N_6107);
or U8604 (N_8604,N_6204,N_7438);
or U8605 (N_8605,N_6257,N_6678);
nor U8606 (N_8606,N_6492,N_6900);
and U8607 (N_8607,N_6929,N_7158);
nand U8608 (N_8608,N_6636,N_7369);
or U8609 (N_8609,N_7144,N_7599);
and U8610 (N_8610,N_6034,N_7735);
or U8611 (N_8611,N_6108,N_6259);
nand U8612 (N_8612,N_7186,N_7441);
or U8613 (N_8613,N_7146,N_6931);
or U8614 (N_8614,N_7343,N_6972);
and U8615 (N_8615,N_6004,N_6599);
or U8616 (N_8616,N_7331,N_7184);
nor U8617 (N_8617,N_7598,N_7978);
or U8618 (N_8618,N_6687,N_6556);
or U8619 (N_8619,N_6580,N_6097);
and U8620 (N_8620,N_6612,N_6233);
nor U8621 (N_8621,N_7416,N_6100);
nand U8622 (N_8622,N_6214,N_6503);
and U8623 (N_8623,N_7825,N_6295);
nand U8624 (N_8624,N_7937,N_6195);
xnor U8625 (N_8625,N_7473,N_7998);
or U8626 (N_8626,N_6820,N_6055);
nor U8627 (N_8627,N_6105,N_6099);
and U8628 (N_8628,N_6224,N_6145);
or U8629 (N_8629,N_7748,N_6875);
nor U8630 (N_8630,N_6886,N_6928);
nor U8631 (N_8631,N_6799,N_7429);
nor U8632 (N_8632,N_6917,N_7286);
or U8633 (N_8633,N_6751,N_6125);
nor U8634 (N_8634,N_6937,N_7461);
xnor U8635 (N_8635,N_7520,N_6549);
nand U8636 (N_8636,N_6871,N_6062);
and U8637 (N_8637,N_7462,N_6111);
and U8638 (N_8638,N_6505,N_7983);
and U8639 (N_8639,N_6519,N_7220);
or U8640 (N_8640,N_6392,N_7812);
or U8641 (N_8641,N_7367,N_7043);
nor U8642 (N_8642,N_6737,N_6130);
and U8643 (N_8643,N_6950,N_6138);
and U8644 (N_8644,N_6782,N_6977);
or U8645 (N_8645,N_6306,N_6222);
or U8646 (N_8646,N_6137,N_7454);
or U8647 (N_8647,N_6238,N_6543);
or U8648 (N_8648,N_7792,N_6234);
nand U8649 (N_8649,N_6136,N_7373);
or U8650 (N_8650,N_6426,N_6661);
nand U8651 (N_8651,N_7729,N_7728);
nor U8652 (N_8652,N_6032,N_6299);
and U8653 (N_8653,N_6196,N_7058);
and U8654 (N_8654,N_7244,N_6244);
or U8655 (N_8655,N_7661,N_7564);
or U8656 (N_8656,N_7177,N_6913);
and U8657 (N_8657,N_6772,N_7899);
nor U8658 (N_8658,N_7807,N_6534);
or U8659 (N_8659,N_7741,N_7482);
or U8660 (N_8660,N_7447,N_6885);
or U8661 (N_8661,N_7809,N_7725);
nand U8662 (N_8662,N_7355,N_7481);
or U8663 (N_8663,N_6453,N_6302);
and U8664 (N_8664,N_6646,N_7105);
nand U8665 (N_8665,N_6823,N_6825);
nor U8666 (N_8666,N_6567,N_6237);
nor U8667 (N_8667,N_7434,N_6121);
nor U8668 (N_8668,N_6891,N_7344);
nor U8669 (N_8669,N_7610,N_7775);
nor U8670 (N_8670,N_7953,N_7907);
or U8671 (N_8671,N_6020,N_7000);
nor U8672 (N_8672,N_7848,N_6998);
and U8673 (N_8673,N_7860,N_7257);
nand U8674 (N_8674,N_6575,N_7997);
nor U8675 (N_8675,N_7751,N_6849);
nor U8676 (N_8676,N_7390,N_6629);
or U8677 (N_8677,N_7913,N_6714);
nor U8678 (N_8678,N_7235,N_7555);
nor U8679 (N_8679,N_7871,N_6094);
nor U8680 (N_8680,N_7666,N_6723);
nor U8681 (N_8681,N_6388,N_7011);
nor U8682 (N_8682,N_7711,N_6808);
nand U8683 (N_8683,N_7874,N_7347);
and U8684 (N_8684,N_6343,N_6225);
or U8685 (N_8685,N_7103,N_7065);
nand U8686 (N_8686,N_7900,N_7100);
and U8687 (N_8687,N_7878,N_7019);
nand U8688 (N_8688,N_7514,N_7964);
nor U8689 (N_8689,N_7472,N_6247);
or U8690 (N_8690,N_6141,N_7428);
nor U8691 (N_8691,N_6206,N_6174);
nor U8692 (N_8692,N_6283,N_6800);
nand U8693 (N_8693,N_7950,N_6297);
nor U8694 (N_8694,N_6709,N_7817);
nand U8695 (N_8695,N_6482,N_6415);
and U8696 (N_8696,N_7453,N_6596);
and U8697 (N_8697,N_6531,N_7526);
nand U8698 (N_8698,N_6644,N_6176);
or U8699 (N_8699,N_6848,N_6576);
nand U8700 (N_8700,N_6911,N_7824);
nor U8701 (N_8701,N_6971,N_7174);
nand U8702 (N_8702,N_6419,N_7195);
nand U8703 (N_8703,N_6047,N_6809);
nor U8704 (N_8704,N_6079,N_7229);
and U8705 (N_8705,N_6757,N_7571);
nor U8706 (N_8706,N_7245,N_6719);
and U8707 (N_8707,N_7962,N_6515);
nand U8708 (N_8708,N_6882,N_7409);
and U8709 (N_8709,N_7721,N_7354);
nor U8710 (N_8710,N_6113,N_7052);
or U8711 (N_8711,N_7063,N_6528);
or U8712 (N_8712,N_6585,N_7091);
nor U8713 (N_8713,N_6812,N_7621);
or U8714 (N_8714,N_7031,N_6103);
nor U8715 (N_8715,N_7696,N_6194);
and U8716 (N_8716,N_7519,N_7259);
nor U8717 (N_8717,N_6329,N_6155);
and U8718 (N_8718,N_7124,N_7408);
nor U8719 (N_8719,N_7552,N_6568);
nor U8720 (N_8720,N_7760,N_6330);
or U8721 (N_8721,N_6716,N_6867);
and U8722 (N_8722,N_7989,N_6547);
nor U8723 (N_8723,N_6821,N_6178);
nor U8724 (N_8724,N_6618,N_7590);
nor U8725 (N_8725,N_6035,N_6459);
nor U8726 (N_8726,N_7172,N_6918);
and U8727 (N_8727,N_6357,N_7645);
nor U8728 (N_8728,N_7867,N_6175);
nor U8729 (N_8729,N_7834,N_6803);
or U8730 (N_8730,N_7160,N_6781);
nor U8731 (N_8731,N_7887,N_7789);
or U8732 (N_8732,N_6704,N_6248);
nor U8733 (N_8733,N_6081,N_6680);
and U8734 (N_8734,N_7327,N_6759);
nor U8735 (N_8735,N_7938,N_7912);
nor U8736 (N_8736,N_7667,N_6988);
nand U8737 (N_8737,N_7455,N_7196);
and U8738 (N_8738,N_7328,N_6693);
nand U8739 (N_8739,N_7947,N_6486);
nand U8740 (N_8740,N_7387,N_7765);
nand U8741 (N_8741,N_7318,N_7060);
and U8742 (N_8742,N_6218,N_6581);
nor U8743 (N_8743,N_6152,N_6707);
and U8744 (N_8744,N_7839,N_7127);
and U8745 (N_8745,N_7638,N_7510);
or U8746 (N_8746,N_6500,N_6974);
or U8747 (N_8747,N_6423,N_7357);
nand U8748 (N_8748,N_6114,N_6325);
or U8749 (N_8749,N_6033,N_7759);
nor U8750 (N_8750,N_7668,N_6741);
or U8751 (N_8751,N_7341,N_7120);
nand U8752 (N_8752,N_7458,N_7518);
or U8753 (N_8753,N_7271,N_6674);
nand U8754 (N_8754,N_6814,N_6102);
and U8755 (N_8755,N_7797,N_7981);
or U8756 (N_8756,N_7624,N_6227);
nand U8757 (N_8757,N_6148,N_6949);
nor U8758 (N_8758,N_7067,N_6190);
nand U8759 (N_8759,N_7879,N_6028);
and U8760 (N_8760,N_7094,N_7630);
nor U8761 (N_8761,N_6638,N_6948);
and U8762 (N_8762,N_7261,N_6290);
or U8763 (N_8763,N_7940,N_6452);
nor U8764 (N_8764,N_6313,N_6711);
or U8765 (N_8765,N_6754,N_7457);
nand U8766 (N_8766,N_7553,N_7378);
nand U8767 (N_8767,N_6860,N_7311);
or U8768 (N_8768,N_7916,N_6673);
nand U8769 (N_8769,N_7036,N_7152);
or U8770 (N_8770,N_7511,N_6131);
nor U8771 (N_8771,N_6334,N_7898);
or U8772 (N_8772,N_7865,N_6642);
nor U8773 (N_8773,N_6696,N_7755);
and U8774 (N_8774,N_6836,N_6050);
and U8775 (N_8775,N_6694,N_7480);
xor U8776 (N_8776,N_7603,N_6254);
or U8777 (N_8777,N_7847,N_7276);
or U8778 (N_8778,N_6827,N_6326);
nand U8779 (N_8779,N_6669,N_6054);
nor U8780 (N_8780,N_7591,N_7990);
nor U8781 (N_8781,N_6408,N_6096);
and U8782 (N_8782,N_6068,N_6091);
nand U8783 (N_8783,N_6077,N_7284);
nand U8784 (N_8784,N_7227,N_7776);
nand U8785 (N_8785,N_6526,N_7230);
or U8786 (N_8786,N_6018,N_7126);
nor U8787 (N_8787,N_7108,N_6774);
nand U8788 (N_8788,N_6909,N_6300);
nor U8789 (N_8789,N_6064,N_7456);
or U8790 (N_8790,N_6273,N_6946);
nor U8791 (N_8791,N_7322,N_6280);
nor U8792 (N_8792,N_7837,N_7444);
and U8793 (N_8793,N_7562,N_7917);
nand U8794 (N_8794,N_6993,N_6923);
or U8795 (N_8795,N_6360,N_6999);
or U8796 (N_8796,N_7976,N_7266);
nor U8797 (N_8797,N_6046,N_7672);
or U8798 (N_8798,N_6002,N_6397);
nand U8799 (N_8799,N_7411,N_7371);
and U8800 (N_8800,N_7960,N_6475);
or U8801 (N_8801,N_7691,N_6367);
or U8802 (N_8802,N_6323,N_6904);
and U8803 (N_8803,N_6856,N_6983);
and U8804 (N_8804,N_7971,N_7743);
and U8805 (N_8805,N_7533,N_6110);
nor U8806 (N_8806,N_6045,N_7784);
or U8807 (N_8807,N_7047,N_7822);
nor U8808 (N_8808,N_7679,N_6065);
or U8809 (N_8809,N_6396,N_7500);
or U8810 (N_8810,N_6182,N_7675);
nand U8811 (N_8811,N_7766,N_7996);
or U8812 (N_8812,N_6310,N_6787);
nand U8813 (N_8813,N_6973,N_7895);
or U8814 (N_8814,N_7924,N_7715);
or U8815 (N_8815,N_6540,N_7115);
nor U8816 (N_8816,N_6627,N_6878);
or U8817 (N_8817,N_6150,N_6570);
nor U8818 (N_8818,N_7596,N_6348);
or U8819 (N_8819,N_6001,N_7777);
nand U8820 (N_8820,N_6771,N_6794);
or U8821 (N_8821,N_7466,N_6023);
nand U8822 (N_8822,N_7756,N_6511);
nor U8823 (N_8823,N_7649,N_7651);
nand U8824 (N_8824,N_6006,N_7723);
or U8825 (N_8825,N_7629,N_7383);
and U8826 (N_8826,N_7405,N_6606);
nand U8827 (N_8827,N_7923,N_7864);
nor U8828 (N_8828,N_7606,N_7380);
or U8829 (N_8829,N_6670,N_7136);
or U8830 (N_8830,N_6393,N_6078);
and U8831 (N_8831,N_6682,N_7260);
nor U8832 (N_8832,N_6976,N_7099);
or U8833 (N_8833,N_6216,N_6366);
nand U8834 (N_8834,N_6305,N_6086);
and U8835 (N_8835,N_6339,N_7151);
nand U8836 (N_8836,N_7722,N_6516);
or U8837 (N_8837,N_6951,N_7039);
and U8838 (N_8838,N_6483,N_6092);
or U8839 (N_8839,N_6364,N_7129);
or U8840 (N_8840,N_7391,N_7588);
nand U8841 (N_8841,N_6435,N_6777);
nand U8842 (N_8842,N_6404,N_7791);
and U8843 (N_8843,N_7939,N_6603);
nand U8844 (N_8844,N_7673,N_7680);
xor U8845 (N_8845,N_7531,N_6307);
and U8846 (N_8846,N_6119,N_6164);
nand U8847 (N_8847,N_7653,N_7746);
or U8848 (N_8848,N_7304,N_7403);
nand U8849 (N_8849,N_7642,N_7004);
or U8850 (N_8850,N_7609,N_7767);
or U8851 (N_8851,N_6753,N_6294);
or U8852 (N_8852,N_7291,N_7846);
and U8853 (N_8853,N_7045,N_6200);
and U8854 (N_8854,N_6965,N_6051);
and U8855 (N_8855,N_6411,N_7038);
nand U8856 (N_8856,N_6884,N_7423);
or U8857 (N_8857,N_6797,N_6363);
nand U8858 (N_8858,N_6271,N_6729);
and U8859 (N_8859,N_7547,N_7055);
and U8860 (N_8860,N_7353,N_7406);
xnor U8861 (N_8861,N_6284,N_6989);
nand U8862 (N_8862,N_7524,N_7655);
or U8863 (N_8863,N_6123,N_6509);
nor U8864 (N_8864,N_7463,N_7922);
nand U8865 (N_8865,N_7974,N_7810);
nand U8866 (N_8866,N_6641,N_6258);
and U8867 (N_8867,N_7109,N_6242);
nor U8868 (N_8868,N_7987,N_6098);
nand U8869 (N_8869,N_6956,N_6374);
or U8870 (N_8870,N_7654,N_6637);
or U8871 (N_8871,N_6465,N_7006);
nand U8872 (N_8872,N_6750,N_6116);
nor U8873 (N_8873,N_6009,N_7024);
or U8874 (N_8874,N_7941,N_6508);
and U8875 (N_8875,N_6029,N_6529);
and U8876 (N_8876,N_7389,N_7187);
nor U8877 (N_8877,N_7914,N_7162);
nor U8878 (N_8878,N_6571,N_7135);
nor U8879 (N_8879,N_7119,N_7662);
and U8880 (N_8880,N_6165,N_7064);
nand U8881 (N_8881,N_7707,N_6819);
nor U8882 (N_8882,N_7392,N_7419);
nor U8883 (N_8883,N_6930,N_6027);
or U8884 (N_8884,N_7840,N_6907);
nor U8885 (N_8885,N_7516,N_7431);
and U8886 (N_8886,N_7489,N_6776);
nor U8887 (N_8887,N_6536,N_7835);
nand U8888 (N_8888,N_6952,N_6874);
or U8889 (N_8889,N_7081,N_7905);
nand U8890 (N_8890,N_7224,N_7979);
nand U8891 (N_8891,N_6961,N_6610);
nand U8892 (N_8892,N_6639,N_7350);
and U8893 (N_8893,N_6813,N_7674);
and U8894 (N_8894,N_6523,N_7290);
xor U8895 (N_8895,N_7850,N_6417);
nor U8896 (N_8896,N_6935,N_6791);
or U8897 (N_8897,N_7145,N_6231);
and U8898 (N_8898,N_6179,N_7025);
nand U8899 (N_8899,N_6384,N_7087);
and U8900 (N_8900,N_6876,N_6826);
or U8901 (N_8901,N_7557,N_6602);
nand U8902 (N_8902,N_6869,N_6335);
and U8903 (N_8903,N_6594,N_6862);
or U8904 (N_8904,N_6128,N_6520);
or U8905 (N_8905,N_7071,N_6655);
or U8906 (N_8906,N_7337,N_6562);
or U8907 (N_8907,N_7097,N_7745);
nand U8908 (N_8908,N_6614,N_7407);
and U8909 (N_8909,N_6496,N_7101);
or U8910 (N_8910,N_6968,N_6579);
or U8911 (N_8911,N_6910,N_7795);
or U8912 (N_8912,N_6250,N_7080);
or U8913 (N_8913,N_6922,N_7442);
nor U8914 (N_8914,N_6126,N_6015);
nand U8915 (N_8915,N_6615,N_7182);
nor U8916 (N_8916,N_6726,N_6597);
nand U8917 (N_8917,N_7929,N_7845);
and U8918 (N_8918,N_7771,N_7540);
or U8919 (N_8919,N_7307,N_7858);
or U8920 (N_8920,N_6276,N_6275);
nand U8921 (N_8921,N_6303,N_6686);
nor U8922 (N_8922,N_7275,N_7342);
nand U8923 (N_8923,N_6395,N_7772);
and U8924 (N_8924,N_6321,N_6451);
or U8925 (N_8925,N_7782,N_7274);
or U8926 (N_8926,N_7421,N_7535);
nor U8927 (N_8927,N_6698,N_6851);
nor U8928 (N_8928,N_7205,N_7139);
and U8929 (N_8929,N_6589,N_6648);
nand U8930 (N_8930,N_6832,N_6525);
and U8931 (N_8931,N_7863,N_6969);
nand U8932 (N_8932,N_6902,N_6953);
or U8933 (N_8933,N_6167,N_6072);
or U8934 (N_8934,N_7593,N_6666);
and U8935 (N_8935,N_6376,N_7418);
nor U8936 (N_8936,N_7550,N_6223);
nand U8937 (N_8937,N_7683,N_7399);
nand U8938 (N_8938,N_7027,N_7420);
nor U8939 (N_8939,N_6090,N_7194);
nor U8940 (N_8940,N_7734,N_6578);
and U8941 (N_8941,N_6621,N_7106);
nor U8942 (N_8942,N_6811,N_7263);
nor U8943 (N_8943,N_6309,N_7238);
and U8944 (N_8944,N_6479,N_6933);
and U8945 (N_8945,N_6066,N_7007);
nand U8946 (N_8946,N_7207,N_7894);
nand U8947 (N_8947,N_7585,N_6530);
nand U8948 (N_8948,N_7616,N_7517);
or U8949 (N_8949,N_6657,N_7806);
or U8950 (N_8950,N_7312,N_6381);
nand U8951 (N_8951,N_7191,N_7814);
nand U8952 (N_8952,N_6598,N_7919);
and U8953 (N_8953,N_6447,N_6894);
nor U8954 (N_8954,N_7239,N_6991);
nand U8955 (N_8955,N_6896,N_7057);
and U8956 (N_8956,N_7768,N_7125);
nand U8957 (N_8957,N_7465,N_7966);
or U8958 (N_8958,N_7882,N_7783);
and U8959 (N_8959,N_7098,N_6994);
and U8960 (N_8960,N_7425,N_7975);
nand U8961 (N_8961,N_7240,N_6056);
nor U8962 (N_8962,N_6311,N_6073);
nand U8963 (N_8963,N_7475,N_6720);
and U8964 (N_8964,N_6901,N_7216);
and U8965 (N_8965,N_6286,N_7926);
or U8966 (N_8966,N_7788,N_6865);
nand U8967 (N_8967,N_6740,N_6514);
nor U8968 (N_8968,N_7665,N_6609);
nand U8969 (N_8969,N_6438,N_6480);
nor U8970 (N_8970,N_7396,N_6118);
and U8971 (N_8971,N_6841,N_6692);
and U8972 (N_8972,N_7270,N_6277);
nor U8973 (N_8973,N_7424,N_6039);
or U8974 (N_8974,N_6243,N_7211);
xor U8975 (N_8975,N_7565,N_6122);
or U8976 (N_8976,N_7076,N_7231);
nand U8977 (N_8977,N_6850,N_7764);
or U8978 (N_8978,N_6336,N_7577);
or U8979 (N_8979,N_6888,N_6934);
or U8980 (N_8980,N_7861,N_7082);
nor U8981 (N_8981,N_7801,N_6007);
or U8982 (N_8982,N_6044,N_7648);
or U8983 (N_8983,N_7559,N_7140);
and U8984 (N_8984,N_7574,N_6887);
nor U8985 (N_8985,N_7273,N_7818);
nand U8986 (N_8986,N_7556,N_7868);
or U8987 (N_8987,N_6246,N_6554);
nand U8988 (N_8988,N_7476,N_7381);
nor U8989 (N_8989,N_7267,N_6253);
nand U8990 (N_8990,N_6779,N_7278);
nand U8991 (N_8991,N_6022,N_7479);
nor U8992 (N_8992,N_7713,N_7701);
nand U8993 (N_8993,N_7029,N_7657);
and U8994 (N_8994,N_6340,N_6472);
nand U8995 (N_8995,N_6037,N_6474);
nor U8996 (N_8996,N_6889,N_6818);
nand U8997 (N_8997,N_7640,N_7573);
and U8998 (N_8998,N_7415,N_7702);
or U8999 (N_8999,N_6840,N_7452);
nand U9000 (N_9000,N_7760,N_6590);
nor U9001 (N_9001,N_7373,N_6037);
and U9002 (N_9002,N_6239,N_6633);
and U9003 (N_9003,N_7400,N_6929);
nor U9004 (N_9004,N_7161,N_6282);
or U9005 (N_9005,N_7536,N_7047);
or U9006 (N_9006,N_6657,N_7300);
nor U9007 (N_9007,N_6570,N_6067);
nor U9008 (N_9008,N_7686,N_7693);
and U9009 (N_9009,N_7744,N_6915);
and U9010 (N_9010,N_7501,N_7326);
and U9011 (N_9011,N_6176,N_7791);
nand U9012 (N_9012,N_7277,N_7266);
and U9013 (N_9013,N_6765,N_7424);
nand U9014 (N_9014,N_7073,N_7539);
nor U9015 (N_9015,N_6982,N_6635);
nor U9016 (N_9016,N_7726,N_7524);
or U9017 (N_9017,N_6949,N_6487);
and U9018 (N_9018,N_7137,N_7296);
or U9019 (N_9019,N_6401,N_6995);
nor U9020 (N_9020,N_6577,N_6203);
or U9021 (N_9021,N_6236,N_6690);
or U9022 (N_9022,N_6446,N_6610);
nor U9023 (N_9023,N_6458,N_6735);
and U9024 (N_9024,N_6442,N_6721);
nor U9025 (N_9025,N_6019,N_6632);
and U9026 (N_9026,N_6967,N_6244);
or U9027 (N_9027,N_7811,N_6537);
and U9028 (N_9028,N_7133,N_7807);
and U9029 (N_9029,N_7747,N_6075);
and U9030 (N_9030,N_7470,N_7531);
or U9031 (N_9031,N_6072,N_6221);
or U9032 (N_9032,N_6792,N_6782);
nor U9033 (N_9033,N_7956,N_7377);
and U9034 (N_9034,N_7930,N_7457);
nand U9035 (N_9035,N_7456,N_6661);
and U9036 (N_9036,N_6160,N_6759);
nand U9037 (N_9037,N_6972,N_6264);
nand U9038 (N_9038,N_7472,N_6520);
nand U9039 (N_9039,N_7940,N_7392);
or U9040 (N_9040,N_6154,N_7760);
nor U9041 (N_9041,N_7958,N_6135);
or U9042 (N_9042,N_6564,N_7671);
or U9043 (N_9043,N_6908,N_7516);
nand U9044 (N_9044,N_6253,N_6787);
and U9045 (N_9045,N_6137,N_7250);
nor U9046 (N_9046,N_7879,N_6829);
nor U9047 (N_9047,N_7200,N_7955);
and U9048 (N_9048,N_7990,N_7878);
nor U9049 (N_9049,N_7674,N_6591);
nor U9050 (N_9050,N_6140,N_7275);
or U9051 (N_9051,N_6275,N_7555);
or U9052 (N_9052,N_7364,N_6302);
nor U9053 (N_9053,N_7536,N_6016);
nand U9054 (N_9054,N_6752,N_6692);
nand U9055 (N_9055,N_7065,N_7963);
nor U9056 (N_9056,N_7923,N_7011);
nand U9057 (N_9057,N_6338,N_6888);
or U9058 (N_9058,N_6543,N_7585);
nor U9059 (N_9059,N_6812,N_6169);
nand U9060 (N_9060,N_6707,N_6698);
and U9061 (N_9061,N_7700,N_6164);
nand U9062 (N_9062,N_7210,N_7832);
xnor U9063 (N_9063,N_6436,N_7041);
nor U9064 (N_9064,N_6658,N_7175);
and U9065 (N_9065,N_6335,N_7667);
nor U9066 (N_9066,N_7274,N_6788);
nor U9067 (N_9067,N_7756,N_7181);
and U9068 (N_9068,N_7164,N_6790);
nor U9069 (N_9069,N_6930,N_7712);
nor U9070 (N_9070,N_6283,N_6545);
and U9071 (N_9071,N_6692,N_7362);
or U9072 (N_9072,N_7109,N_7592);
or U9073 (N_9073,N_6208,N_7521);
nor U9074 (N_9074,N_7717,N_7670);
nor U9075 (N_9075,N_6877,N_7271);
nand U9076 (N_9076,N_7062,N_6879);
and U9077 (N_9077,N_6433,N_6841);
nor U9078 (N_9078,N_7759,N_6343);
nand U9079 (N_9079,N_7818,N_7624);
or U9080 (N_9080,N_6516,N_7453);
nor U9081 (N_9081,N_6342,N_6574);
or U9082 (N_9082,N_7625,N_6818);
and U9083 (N_9083,N_7027,N_7709);
nor U9084 (N_9084,N_6009,N_7500);
and U9085 (N_9085,N_6645,N_7059);
nor U9086 (N_9086,N_6269,N_6092);
nor U9087 (N_9087,N_7860,N_6084);
nor U9088 (N_9088,N_6542,N_7379);
nor U9089 (N_9089,N_7579,N_7254);
and U9090 (N_9090,N_6478,N_7512);
or U9091 (N_9091,N_7020,N_7425);
nand U9092 (N_9092,N_7205,N_6772);
nand U9093 (N_9093,N_6915,N_7986);
nor U9094 (N_9094,N_7072,N_7818);
or U9095 (N_9095,N_7289,N_7129);
nor U9096 (N_9096,N_6117,N_7669);
and U9097 (N_9097,N_6404,N_7677);
xor U9098 (N_9098,N_6759,N_6452);
and U9099 (N_9099,N_7563,N_7650);
nand U9100 (N_9100,N_7709,N_7804);
nor U9101 (N_9101,N_6684,N_7198);
nand U9102 (N_9102,N_7961,N_7548);
nand U9103 (N_9103,N_7349,N_7408);
or U9104 (N_9104,N_6932,N_7074);
nand U9105 (N_9105,N_6092,N_7828);
nor U9106 (N_9106,N_7085,N_7982);
nand U9107 (N_9107,N_7884,N_7227);
nand U9108 (N_9108,N_7891,N_6081);
xor U9109 (N_9109,N_7032,N_6299);
and U9110 (N_9110,N_6232,N_6250);
and U9111 (N_9111,N_6768,N_7605);
and U9112 (N_9112,N_6362,N_7933);
or U9113 (N_9113,N_7827,N_7304);
nand U9114 (N_9114,N_7426,N_7842);
or U9115 (N_9115,N_7714,N_7551);
and U9116 (N_9116,N_7149,N_7509);
nand U9117 (N_9117,N_6781,N_7061);
nor U9118 (N_9118,N_6736,N_7973);
and U9119 (N_9119,N_6766,N_7956);
and U9120 (N_9120,N_6883,N_7311);
nand U9121 (N_9121,N_7347,N_6896);
nor U9122 (N_9122,N_6959,N_7842);
nand U9123 (N_9123,N_6553,N_7652);
or U9124 (N_9124,N_7296,N_6465);
nand U9125 (N_9125,N_6422,N_7634);
or U9126 (N_9126,N_6495,N_7579);
nor U9127 (N_9127,N_6019,N_7023);
or U9128 (N_9128,N_7495,N_6655);
nor U9129 (N_9129,N_7270,N_6748);
nand U9130 (N_9130,N_7274,N_6687);
nor U9131 (N_9131,N_7401,N_6981);
nand U9132 (N_9132,N_6097,N_7537);
nor U9133 (N_9133,N_6956,N_6111);
nor U9134 (N_9134,N_7151,N_6205);
nor U9135 (N_9135,N_7329,N_7855);
or U9136 (N_9136,N_6027,N_7602);
nor U9137 (N_9137,N_6103,N_7878);
or U9138 (N_9138,N_6397,N_6275);
and U9139 (N_9139,N_7001,N_7883);
nor U9140 (N_9140,N_6786,N_6500);
nand U9141 (N_9141,N_6744,N_7769);
and U9142 (N_9142,N_7274,N_7292);
and U9143 (N_9143,N_7874,N_7836);
or U9144 (N_9144,N_7576,N_7488);
nor U9145 (N_9145,N_7613,N_6517);
nand U9146 (N_9146,N_6355,N_7689);
xnor U9147 (N_9147,N_7720,N_7053);
and U9148 (N_9148,N_6375,N_7101);
nand U9149 (N_9149,N_7559,N_7907);
and U9150 (N_9150,N_7449,N_6508);
nor U9151 (N_9151,N_7002,N_7433);
or U9152 (N_9152,N_7244,N_7597);
and U9153 (N_9153,N_7910,N_6383);
or U9154 (N_9154,N_7155,N_6620);
nand U9155 (N_9155,N_6301,N_6817);
nor U9156 (N_9156,N_7670,N_6448);
and U9157 (N_9157,N_6239,N_6953);
nand U9158 (N_9158,N_6714,N_6212);
nor U9159 (N_9159,N_7702,N_7058);
nor U9160 (N_9160,N_6707,N_7736);
or U9161 (N_9161,N_6398,N_7548);
and U9162 (N_9162,N_6699,N_6848);
or U9163 (N_9163,N_6776,N_6533);
nor U9164 (N_9164,N_6545,N_7722);
nand U9165 (N_9165,N_7784,N_6558);
nand U9166 (N_9166,N_6306,N_7637);
nand U9167 (N_9167,N_7686,N_7617);
nor U9168 (N_9168,N_7654,N_6900);
and U9169 (N_9169,N_6723,N_6248);
nand U9170 (N_9170,N_7265,N_7703);
nand U9171 (N_9171,N_6096,N_7527);
or U9172 (N_9172,N_7084,N_6401);
or U9173 (N_9173,N_6086,N_6735);
or U9174 (N_9174,N_6161,N_7662);
nor U9175 (N_9175,N_7823,N_7061);
or U9176 (N_9176,N_6869,N_6029);
and U9177 (N_9177,N_7434,N_6578);
nor U9178 (N_9178,N_6466,N_7327);
and U9179 (N_9179,N_7323,N_7271);
nand U9180 (N_9180,N_6391,N_6181);
nand U9181 (N_9181,N_6658,N_7193);
xor U9182 (N_9182,N_7711,N_7655);
and U9183 (N_9183,N_7810,N_6623);
nand U9184 (N_9184,N_7235,N_7782);
nand U9185 (N_9185,N_6186,N_7227);
or U9186 (N_9186,N_7688,N_7547);
or U9187 (N_9187,N_6949,N_6691);
nor U9188 (N_9188,N_6906,N_7004);
and U9189 (N_9189,N_7562,N_6750);
and U9190 (N_9190,N_6448,N_6882);
nand U9191 (N_9191,N_7271,N_6436);
nand U9192 (N_9192,N_6437,N_6338);
or U9193 (N_9193,N_7807,N_6018);
and U9194 (N_9194,N_6025,N_6751);
or U9195 (N_9195,N_7086,N_7565);
xor U9196 (N_9196,N_6229,N_6244);
nor U9197 (N_9197,N_7382,N_6348);
nor U9198 (N_9198,N_6029,N_7017);
or U9199 (N_9199,N_6734,N_7577);
or U9200 (N_9200,N_7328,N_7001);
nand U9201 (N_9201,N_6458,N_6456);
nand U9202 (N_9202,N_7081,N_7538);
or U9203 (N_9203,N_7988,N_6269);
and U9204 (N_9204,N_7774,N_7265);
and U9205 (N_9205,N_6517,N_6016);
or U9206 (N_9206,N_7514,N_7609);
and U9207 (N_9207,N_7966,N_7177);
and U9208 (N_9208,N_7081,N_6182);
or U9209 (N_9209,N_7208,N_7921);
nor U9210 (N_9210,N_6669,N_7636);
and U9211 (N_9211,N_6130,N_7589);
and U9212 (N_9212,N_7656,N_6957);
nor U9213 (N_9213,N_7376,N_6821);
nand U9214 (N_9214,N_6212,N_6167);
nor U9215 (N_9215,N_6055,N_6998);
or U9216 (N_9216,N_7646,N_6027);
nor U9217 (N_9217,N_6685,N_7866);
nor U9218 (N_9218,N_7542,N_7162);
nand U9219 (N_9219,N_6156,N_6068);
or U9220 (N_9220,N_7805,N_6566);
and U9221 (N_9221,N_6134,N_7053);
and U9222 (N_9222,N_6036,N_7339);
or U9223 (N_9223,N_6603,N_7576);
nand U9224 (N_9224,N_7356,N_6216);
nand U9225 (N_9225,N_6659,N_7754);
nand U9226 (N_9226,N_7806,N_6854);
nor U9227 (N_9227,N_6803,N_7776);
and U9228 (N_9228,N_6832,N_6454);
or U9229 (N_9229,N_6005,N_6163);
and U9230 (N_9230,N_6446,N_7588);
and U9231 (N_9231,N_7891,N_7213);
nand U9232 (N_9232,N_6845,N_6475);
and U9233 (N_9233,N_7664,N_7651);
nor U9234 (N_9234,N_7157,N_6825);
nor U9235 (N_9235,N_7268,N_6766);
nand U9236 (N_9236,N_6965,N_6916);
nand U9237 (N_9237,N_7697,N_6249);
nor U9238 (N_9238,N_7418,N_7813);
nand U9239 (N_9239,N_6320,N_6298);
and U9240 (N_9240,N_7221,N_6349);
and U9241 (N_9241,N_7004,N_6994);
and U9242 (N_9242,N_7300,N_7735);
nand U9243 (N_9243,N_7060,N_7114);
nor U9244 (N_9244,N_6847,N_7871);
nand U9245 (N_9245,N_7743,N_6874);
nand U9246 (N_9246,N_6893,N_6523);
nand U9247 (N_9247,N_7898,N_7221);
and U9248 (N_9248,N_6542,N_7080);
nor U9249 (N_9249,N_7928,N_7559);
and U9250 (N_9250,N_7139,N_6977);
or U9251 (N_9251,N_6020,N_6718);
and U9252 (N_9252,N_6005,N_7450);
or U9253 (N_9253,N_6566,N_7521);
or U9254 (N_9254,N_6647,N_6419);
nand U9255 (N_9255,N_6800,N_6648);
nand U9256 (N_9256,N_7071,N_7851);
or U9257 (N_9257,N_7566,N_7580);
and U9258 (N_9258,N_6931,N_7823);
and U9259 (N_9259,N_7613,N_6721);
and U9260 (N_9260,N_7441,N_7998);
nor U9261 (N_9261,N_6846,N_6382);
and U9262 (N_9262,N_6301,N_7662);
or U9263 (N_9263,N_6379,N_7411);
xor U9264 (N_9264,N_6427,N_7986);
or U9265 (N_9265,N_6161,N_7812);
or U9266 (N_9266,N_6994,N_7274);
and U9267 (N_9267,N_6373,N_7183);
nor U9268 (N_9268,N_6789,N_7212);
nand U9269 (N_9269,N_7261,N_6488);
nor U9270 (N_9270,N_7256,N_7024);
nor U9271 (N_9271,N_6927,N_7803);
and U9272 (N_9272,N_7347,N_7251);
nand U9273 (N_9273,N_7333,N_7067);
or U9274 (N_9274,N_7682,N_6258);
and U9275 (N_9275,N_6419,N_7605);
xnor U9276 (N_9276,N_7536,N_7115);
nand U9277 (N_9277,N_7260,N_7734);
nand U9278 (N_9278,N_7123,N_6543);
and U9279 (N_9279,N_7817,N_6531);
and U9280 (N_9280,N_7734,N_6330);
and U9281 (N_9281,N_7550,N_7816);
nor U9282 (N_9282,N_7332,N_7120);
and U9283 (N_9283,N_7048,N_7261);
nand U9284 (N_9284,N_6448,N_7960);
nor U9285 (N_9285,N_6988,N_7528);
xnor U9286 (N_9286,N_6344,N_6994);
nor U9287 (N_9287,N_7266,N_6058);
or U9288 (N_9288,N_6746,N_6902);
nor U9289 (N_9289,N_7876,N_6768);
nand U9290 (N_9290,N_7352,N_7539);
nand U9291 (N_9291,N_7939,N_6132);
and U9292 (N_9292,N_6266,N_6887);
nor U9293 (N_9293,N_6474,N_7921);
nor U9294 (N_9294,N_6597,N_6928);
or U9295 (N_9295,N_6584,N_6778);
or U9296 (N_9296,N_6395,N_6127);
nor U9297 (N_9297,N_6859,N_6427);
nand U9298 (N_9298,N_6219,N_6006);
nand U9299 (N_9299,N_6283,N_7829);
and U9300 (N_9300,N_6855,N_7149);
nor U9301 (N_9301,N_7914,N_7275);
and U9302 (N_9302,N_7870,N_6713);
or U9303 (N_9303,N_6640,N_7850);
nand U9304 (N_9304,N_6077,N_7099);
nor U9305 (N_9305,N_7572,N_6446);
nand U9306 (N_9306,N_7069,N_6831);
nand U9307 (N_9307,N_6074,N_7275);
nand U9308 (N_9308,N_7973,N_7592);
nand U9309 (N_9309,N_6442,N_7154);
or U9310 (N_9310,N_6636,N_7827);
or U9311 (N_9311,N_6400,N_7601);
and U9312 (N_9312,N_7187,N_7213);
nand U9313 (N_9313,N_7620,N_6097);
or U9314 (N_9314,N_7385,N_7635);
or U9315 (N_9315,N_6369,N_6688);
nand U9316 (N_9316,N_7159,N_7203);
nand U9317 (N_9317,N_7786,N_7414);
nand U9318 (N_9318,N_7360,N_6341);
nor U9319 (N_9319,N_6921,N_7150);
or U9320 (N_9320,N_6473,N_6241);
nor U9321 (N_9321,N_7493,N_6335);
or U9322 (N_9322,N_6057,N_7937);
nor U9323 (N_9323,N_7241,N_7167);
nor U9324 (N_9324,N_7653,N_6119);
and U9325 (N_9325,N_7410,N_7925);
nand U9326 (N_9326,N_7466,N_7064);
nor U9327 (N_9327,N_6603,N_7078);
nor U9328 (N_9328,N_7487,N_6631);
nor U9329 (N_9329,N_6460,N_7659);
or U9330 (N_9330,N_6609,N_6250);
and U9331 (N_9331,N_7760,N_7287);
nor U9332 (N_9332,N_6233,N_6138);
and U9333 (N_9333,N_6728,N_6225);
and U9334 (N_9334,N_7134,N_7817);
nand U9335 (N_9335,N_7547,N_7723);
nand U9336 (N_9336,N_6424,N_7893);
and U9337 (N_9337,N_7494,N_6275);
nand U9338 (N_9338,N_7940,N_6877);
and U9339 (N_9339,N_6944,N_7539);
nand U9340 (N_9340,N_7197,N_7126);
or U9341 (N_9341,N_6619,N_6647);
nand U9342 (N_9342,N_7218,N_6200);
or U9343 (N_9343,N_6260,N_6222);
nand U9344 (N_9344,N_7574,N_6713);
or U9345 (N_9345,N_7693,N_6387);
nor U9346 (N_9346,N_6000,N_7688);
nor U9347 (N_9347,N_6879,N_6066);
nand U9348 (N_9348,N_7105,N_7647);
nand U9349 (N_9349,N_7329,N_6489);
nor U9350 (N_9350,N_7492,N_6741);
nor U9351 (N_9351,N_7697,N_7616);
or U9352 (N_9352,N_7701,N_7092);
and U9353 (N_9353,N_6760,N_7274);
and U9354 (N_9354,N_6387,N_6104);
or U9355 (N_9355,N_6037,N_6888);
and U9356 (N_9356,N_6134,N_7396);
nor U9357 (N_9357,N_7875,N_6718);
and U9358 (N_9358,N_6903,N_7542);
nor U9359 (N_9359,N_6211,N_7619);
or U9360 (N_9360,N_6712,N_6151);
nand U9361 (N_9361,N_6529,N_7318);
nor U9362 (N_9362,N_6095,N_6652);
nand U9363 (N_9363,N_6741,N_7321);
nand U9364 (N_9364,N_7519,N_7657);
and U9365 (N_9365,N_7972,N_6721);
and U9366 (N_9366,N_7747,N_6630);
or U9367 (N_9367,N_6306,N_6538);
nand U9368 (N_9368,N_7921,N_7552);
and U9369 (N_9369,N_7475,N_6800);
nand U9370 (N_9370,N_7586,N_7196);
nor U9371 (N_9371,N_7043,N_6771);
and U9372 (N_9372,N_6669,N_6765);
and U9373 (N_9373,N_7593,N_6714);
nor U9374 (N_9374,N_6304,N_7698);
nor U9375 (N_9375,N_7226,N_7556);
nand U9376 (N_9376,N_6796,N_6704);
nor U9377 (N_9377,N_6197,N_7611);
nand U9378 (N_9378,N_6492,N_7742);
nand U9379 (N_9379,N_6460,N_6214);
or U9380 (N_9380,N_6898,N_7024);
or U9381 (N_9381,N_6664,N_6121);
nand U9382 (N_9382,N_7647,N_6140);
nand U9383 (N_9383,N_7788,N_6752);
nor U9384 (N_9384,N_6533,N_6365);
and U9385 (N_9385,N_6150,N_7841);
nand U9386 (N_9386,N_7433,N_7769);
or U9387 (N_9387,N_6942,N_6338);
nor U9388 (N_9388,N_7380,N_6000);
or U9389 (N_9389,N_6522,N_7828);
and U9390 (N_9390,N_6971,N_6688);
nor U9391 (N_9391,N_7981,N_7672);
nand U9392 (N_9392,N_7801,N_6016);
nor U9393 (N_9393,N_6693,N_6142);
nand U9394 (N_9394,N_6526,N_6109);
or U9395 (N_9395,N_7874,N_6105);
nand U9396 (N_9396,N_7120,N_6643);
or U9397 (N_9397,N_6368,N_6355);
nor U9398 (N_9398,N_6463,N_6818);
and U9399 (N_9399,N_7440,N_6154);
or U9400 (N_9400,N_6869,N_7352);
or U9401 (N_9401,N_7454,N_6918);
and U9402 (N_9402,N_7395,N_7385);
or U9403 (N_9403,N_6637,N_6748);
or U9404 (N_9404,N_7002,N_7631);
nor U9405 (N_9405,N_7435,N_6779);
nor U9406 (N_9406,N_6955,N_7070);
and U9407 (N_9407,N_7363,N_6404);
nor U9408 (N_9408,N_7686,N_7325);
nand U9409 (N_9409,N_7079,N_6412);
nand U9410 (N_9410,N_7481,N_7924);
or U9411 (N_9411,N_6653,N_6717);
and U9412 (N_9412,N_7158,N_6573);
or U9413 (N_9413,N_7930,N_6102);
nor U9414 (N_9414,N_6332,N_6398);
nor U9415 (N_9415,N_6303,N_7813);
or U9416 (N_9416,N_6365,N_7657);
or U9417 (N_9417,N_7677,N_7445);
and U9418 (N_9418,N_6100,N_6269);
nand U9419 (N_9419,N_6452,N_7463);
or U9420 (N_9420,N_7584,N_7301);
nand U9421 (N_9421,N_7413,N_7864);
and U9422 (N_9422,N_7618,N_7332);
or U9423 (N_9423,N_6298,N_6958);
and U9424 (N_9424,N_7524,N_6199);
nor U9425 (N_9425,N_6676,N_6493);
or U9426 (N_9426,N_6500,N_6255);
and U9427 (N_9427,N_6474,N_7423);
and U9428 (N_9428,N_6628,N_6484);
nand U9429 (N_9429,N_6317,N_7227);
nor U9430 (N_9430,N_7034,N_6963);
nand U9431 (N_9431,N_6164,N_6522);
and U9432 (N_9432,N_7063,N_7431);
or U9433 (N_9433,N_6240,N_6605);
nand U9434 (N_9434,N_7007,N_6005);
or U9435 (N_9435,N_7755,N_6642);
and U9436 (N_9436,N_7450,N_6086);
and U9437 (N_9437,N_6429,N_6762);
or U9438 (N_9438,N_6942,N_7114);
and U9439 (N_9439,N_6006,N_7296);
nand U9440 (N_9440,N_7632,N_7588);
nand U9441 (N_9441,N_6214,N_6176);
and U9442 (N_9442,N_6786,N_7905);
nor U9443 (N_9443,N_7219,N_7360);
nor U9444 (N_9444,N_7573,N_6888);
nor U9445 (N_9445,N_7967,N_6330);
or U9446 (N_9446,N_6524,N_7421);
and U9447 (N_9447,N_6569,N_7089);
nand U9448 (N_9448,N_6232,N_6629);
and U9449 (N_9449,N_6713,N_7275);
or U9450 (N_9450,N_6882,N_7464);
or U9451 (N_9451,N_6977,N_6863);
nor U9452 (N_9452,N_7241,N_6270);
and U9453 (N_9453,N_7234,N_6133);
or U9454 (N_9454,N_7446,N_7666);
nor U9455 (N_9455,N_7657,N_7992);
and U9456 (N_9456,N_7084,N_7270);
or U9457 (N_9457,N_6015,N_7128);
nor U9458 (N_9458,N_7799,N_6728);
or U9459 (N_9459,N_6158,N_7211);
or U9460 (N_9460,N_6821,N_6706);
or U9461 (N_9461,N_6476,N_7976);
nand U9462 (N_9462,N_6104,N_7977);
nand U9463 (N_9463,N_7062,N_6741);
nand U9464 (N_9464,N_7035,N_7015);
or U9465 (N_9465,N_7143,N_6982);
nor U9466 (N_9466,N_6640,N_7457);
and U9467 (N_9467,N_6945,N_7145);
and U9468 (N_9468,N_6869,N_7006);
nor U9469 (N_9469,N_6196,N_7281);
nand U9470 (N_9470,N_7386,N_7086);
nor U9471 (N_9471,N_7443,N_6220);
or U9472 (N_9472,N_6788,N_6645);
or U9473 (N_9473,N_6235,N_7021);
and U9474 (N_9474,N_6419,N_6214);
and U9475 (N_9475,N_7673,N_6115);
and U9476 (N_9476,N_7676,N_7984);
nand U9477 (N_9477,N_7193,N_6551);
nand U9478 (N_9478,N_6684,N_7460);
nor U9479 (N_9479,N_6616,N_7184);
and U9480 (N_9480,N_6773,N_7053);
nor U9481 (N_9481,N_7450,N_7498);
nand U9482 (N_9482,N_6550,N_6708);
nor U9483 (N_9483,N_6504,N_6063);
nand U9484 (N_9484,N_7200,N_6243);
and U9485 (N_9485,N_6605,N_6809);
or U9486 (N_9486,N_6157,N_6930);
and U9487 (N_9487,N_6366,N_7967);
nand U9488 (N_9488,N_7998,N_6021);
nor U9489 (N_9489,N_6693,N_6023);
nor U9490 (N_9490,N_6303,N_6698);
and U9491 (N_9491,N_7510,N_7407);
nor U9492 (N_9492,N_6483,N_6435);
nand U9493 (N_9493,N_6272,N_6803);
and U9494 (N_9494,N_6952,N_6912);
or U9495 (N_9495,N_6483,N_7987);
nand U9496 (N_9496,N_7222,N_6812);
xor U9497 (N_9497,N_6417,N_6920);
or U9498 (N_9498,N_6047,N_7533);
or U9499 (N_9499,N_6463,N_7222);
nand U9500 (N_9500,N_6819,N_6589);
nor U9501 (N_9501,N_6424,N_6399);
nor U9502 (N_9502,N_7158,N_7819);
or U9503 (N_9503,N_7429,N_6997);
xor U9504 (N_9504,N_6041,N_7880);
and U9505 (N_9505,N_6303,N_7935);
nand U9506 (N_9506,N_6100,N_6646);
nor U9507 (N_9507,N_6175,N_6336);
xnor U9508 (N_9508,N_7896,N_7269);
or U9509 (N_9509,N_7146,N_7198);
and U9510 (N_9510,N_6349,N_7522);
nand U9511 (N_9511,N_6329,N_6679);
nor U9512 (N_9512,N_7387,N_6559);
and U9513 (N_9513,N_7084,N_7954);
nor U9514 (N_9514,N_7554,N_7698);
or U9515 (N_9515,N_6104,N_7006);
nand U9516 (N_9516,N_6178,N_6942);
nor U9517 (N_9517,N_7623,N_7640);
nor U9518 (N_9518,N_7078,N_6229);
or U9519 (N_9519,N_6501,N_7498);
and U9520 (N_9520,N_7319,N_7271);
and U9521 (N_9521,N_7241,N_6414);
nor U9522 (N_9522,N_6231,N_6602);
nor U9523 (N_9523,N_6353,N_6064);
nand U9524 (N_9524,N_7512,N_7591);
nor U9525 (N_9525,N_7081,N_7053);
and U9526 (N_9526,N_6873,N_6810);
or U9527 (N_9527,N_7784,N_7252);
or U9528 (N_9528,N_7555,N_6522);
and U9529 (N_9529,N_7236,N_7090);
and U9530 (N_9530,N_6372,N_6879);
or U9531 (N_9531,N_6464,N_6634);
and U9532 (N_9532,N_6289,N_7300);
or U9533 (N_9533,N_7612,N_6087);
nand U9534 (N_9534,N_7426,N_6553);
and U9535 (N_9535,N_7628,N_7954);
nand U9536 (N_9536,N_6838,N_7399);
and U9537 (N_9537,N_6659,N_6142);
nor U9538 (N_9538,N_7962,N_6115);
xnor U9539 (N_9539,N_6218,N_6947);
or U9540 (N_9540,N_7445,N_6782);
or U9541 (N_9541,N_7899,N_6823);
and U9542 (N_9542,N_6070,N_6231);
or U9543 (N_9543,N_7291,N_6753);
nand U9544 (N_9544,N_6128,N_7406);
and U9545 (N_9545,N_7298,N_6087);
xnor U9546 (N_9546,N_7196,N_6064);
nor U9547 (N_9547,N_6206,N_6916);
or U9548 (N_9548,N_7055,N_7083);
nor U9549 (N_9549,N_6921,N_7148);
nor U9550 (N_9550,N_6629,N_6890);
or U9551 (N_9551,N_7508,N_6350);
nor U9552 (N_9552,N_7678,N_7749);
or U9553 (N_9553,N_6922,N_7137);
nor U9554 (N_9554,N_6917,N_7364);
nor U9555 (N_9555,N_6114,N_6291);
nand U9556 (N_9556,N_6236,N_6637);
nand U9557 (N_9557,N_7186,N_6192);
nor U9558 (N_9558,N_7585,N_7721);
and U9559 (N_9559,N_7162,N_7194);
and U9560 (N_9560,N_7748,N_7184);
nor U9561 (N_9561,N_6859,N_6071);
and U9562 (N_9562,N_7133,N_7328);
nor U9563 (N_9563,N_7961,N_6453);
nand U9564 (N_9564,N_7637,N_6639);
and U9565 (N_9565,N_6366,N_6378);
nor U9566 (N_9566,N_6623,N_6573);
and U9567 (N_9567,N_6067,N_7077);
and U9568 (N_9568,N_7899,N_7228);
nor U9569 (N_9569,N_7865,N_7133);
and U9570 (N_9570,N_6401,N_7666);
nand U9571 (N_9571,N_7504,N_6488);
nor U9572 (N_9572,N_7377,N_6467);
nor U9573 (N_9573,N_6079,N_7005);
and U9574 (N_9574,N_7109,N_7886);
and U9575 (N_9575,N_6341,N_6109);
nand U9576 (N_9576,N_7114,N_6715);
and U9577 (N_9577,N_6858,N_7271);
or U9578 (N_9578,N_7195,N_7375);
nand U9579 (N_9579,N_7078,N_7602);
nand U9580 (N_9580,N_6624,N_6611);
xnor U9581 (N_9581,N_7877,N_6008);
and U9582 (N_9582,N_6549,N_7943);
or U9583 (N_9583,N_7286,N_6689);
and U9584 (N_9584,N_7234,N_7324);
nor U9585 (N_9585,N_7244,N_7639);
nand U9586 (N_9586,N_6885,N_6829);
nand U9587 (N_9587,N_6056,N_7610);
nand U9588 (N_9588,N_7296,N_7014);
nor U9589 (N_9589,N_7550,N_6226);
nand U9590 (N_9590,N_6973,N_6171);
and U9591 (N_9591,N_6218,N_6729);
and U9592 (N_9592,N_7485,N_6911);
and U9593 (N_9593,N_7557,N_6158);
nor U9594 (N_9594,N_7510,N_6959);
nor U9595 (N_9595,N_6235,N_6657);
nor U9596 (N_9596,N_7392,N_7655);
nand U9597 (N_9597,N_6038,N_6288);
and U9598 (N_9598,N_7520,N_6893);
and U9599 (N_9599,N_6005,N_7409);
and U9600 (N_9600,N_6725,N_7739);
and U9601 (N_9601,N_7896,N_6237);
and U9602 (N_9602,N_6450,N_6748);
and U9603 (N_9603,N_6575,N_7507);
and U9604 (N_9604,N_7811,N_6359);
or U9605 (N_9605,N_6581,N_6456);
or U9606 (N_9606,N_6305,N_7347);
nor U9607 (N_9607,N_7502,N_7248);
and U9608 (N_9608,N_6029,N_7753);
nand U9609 (N_9609,N_7789,N_7832);
nand U9610 (N_9610,N_7164,N_6713);
xor U9611 (N_9611,N_6511,N_7559);
nor U9612 (N_9612,N_7668,N_7432);
or U9613 (N_9613,N_7291,N_6673);
nor U9614 (N_9614,N_6260,N_7711);
or U9615 (N_9615,N_7245,N_7364);
nand U9616 (N_9616,N_6490,N_6777);
nand U9617 (N_9617,N_7556,N_7745);
or U9618 (N_9618,N_7931,N_7150);
or U9619 (N_9619,N_7593,N_6605);
or U9620 (N_9620,N_7388,N_7111);
or U9621 (N_9621,N_6800,N_7705);
and U9622 (N_9622,N_7673,N_6941);
or U9623 (N_9623,N_6854,N_6348);
nor U9624 (N_9624,N_7407,N_7789);
nand U9625 (N_9625,N_6015,N_6655);
and U9626 (N_9626,N_6912,N_7981);
or U9627 (N_9627,N_7734,N_6546);
or U9628 (N_9628,N_7852,N_6028);
nor U9629 (N_9629,N_7380,N_6563);
and U9630 (N_9630,N_6621,N_7318);
or U9631 (N_9631,N_6706,N_7285);
nand U9632 (N_9632,N_6804,N_7315);
or U9633 (N_9633,N_7017,N_7506);
or U9634 (N_9634,N_7413,N_6757);
and U9635 (N_9635,N_7843,N_7268);
nor U9636 (N_9636,N_6219,N_7713);
and U9637 (N_9637,N_7775,N_7833);
nand U9638 (N_9638,N_6063,N_7952);
or U9639 (N_9639,N_7743,N_7089);
nand U9640 (N_9640,N_6263,N_7704);
xnor U9641 (N_9641,N_7082,N_6810);
nor U9642 (N_9642,N_6432,N_7743);
nand U9643 (N_9643,N_7896,N_6045);
nand U9644 (N_9644,N_7954,N_7273);
or U9645 (N_9645,N_6170,N_7361);
nor U9646 (N_9646,N_7850,N_7682);
nand U9647 (N_9647,N_7272,N_6079);
nand U9648 (N_9648,N_7048,N_7672);
nand U9649 (N_9649,N_6025,N_6269);
nor U9650 (N_9650,N_6509,N_6991);
and U9651 (N_9651,N_6305,N_6440);
nand U9652 (N_9652,N_6271,N_7593);
nand U9653 (N_9653,N_7331,N_7633);
nand U9654 (N_9654,N_7370,N_7033);
nand U9655 (N_9655,N_6249,N_6380);
or U9656 (N_9656,N_6393,N_7409);
and U9657 (N_9657,N_7964,N_7706);
or U9658 (N_9658,N_7671,N_7775);
or U9659 (N_9659,N_6379,N_7044);
or U9660 (N_9660,N_7220,N_6746);
or U9661 (N_9661,N_6109,N_7998);
and U9662 (N_9662,N_7960,N_7570);
nor U9663 (N_9663,N_6939,N_6085);
or U9664 (N_9664,N_6875,N_6655);
nor U9665 (N_9665,N_6478,N_6967);
nor U9666 (N_9666,N_6041,N_7953);
nand U9667 (N_9667,N_7246,N_7140);
and U9668 (N_9668,N_7414,N_7958);
nand U9669 (N_9669,N_6597,N_7451);
nor U9670 (N_9670,N_6539,N_7568);
nor U9671 (N_9671,N_6157,N_7862);
or U9672 (N_9672,N_7560,N_6243);
nand U9673 (N_9673,N_7819,N_6375);
nand U9674 (N_9674,N_6158,N_7131);
nor U9675 (N_9675,N_7617,N_7826);
nand U9676 (N_9676,N_6265,N_7375);
or U9677 (N_9677,N_7612,N_7353);
and U9678 (N_9678,N_7371,N_6286);
nor U9679 (N_9679,N_7580,N_7329);
and U9680 (N_9680,N_7934,N_6778);
and U9681 (N_9681,N_7774,N_7294);
nor U9682 (N_9682,N_6736,N_6748);
nand U9683 (N_9683,N_6569,N_6578);
nand U9684 (N_9684,N_7783,N_7759);
and U9685 (N_9685,N_7433,N_7797);
or U9686 (N_9686,N_6090,N_6244);
and U9687 (N_9687,N_6679,N_7711);
or U9688 (N_9688,N_7246,N_6028);
and U9689 (N_9689,N_7760,N_6486);
and U9690 (N_9690,N_6420,N_7086);
or U9691 (N_9691,N_6892,N_6525);
nand U9692 (N_9692,N_7386,N_7664);
or U9693 (N_9693,N_6121,N_7559);
nor U9694 (N_9694,N_7946,N_6284);
nand U9695 (N_9695,N_7480,N_7856);
nor U9696 (N_9696,N_7697,N_7820);
or U9697 (N_9697,N_7818,N_7898);
nor U9698 (N_9698,N_7998,N_6362);
and U9699 (N_9699,N_7974,N_6045);
nand U9700 (N_9700,N_7274,N_7820);
and U9701 (N_9701,N_7844,N_6035);
or U9702 (N_9702,N_6496,N_7511);
or U9703 (N_9703,N_6890,N_6624);
and U9704 (N_9704,N_7602,N_7763);
nand U9705 (N_9705,N_6919,N_7510);
and U9706 (N_9706,N_7265,N_6979);
nand U9707 (N_9707,N_6524,N_6207);
nor U9708 (N_9708,N_6656,N_6572);
nor U9709 (N_9709,N_6786,N_6891);
and U9710 (N_9710,N_7428,N_6156);
and U9711 (N_9711,N_7710,N_6415);
or U9712 (N_9712,N_7043,N_7053);
or U9713 (N_9713,N_6049,N_7129);
nand U9714 (N_9714,N_6179,N_7553);
nand U9715 (N_9715,N_6044,N_7146);
and U9716 (N_9716,N_6509,N_7068);
and U9717 (N_9717,N_7392,N_6921);
nand U9718 (N_9718,N_6669,N_7294);
or U9719 (N_9719,N_7130,N_7415);
and U9720 (N_9720,N_6768,N_7451);
and U9721 (N_9721,N_6007,N_7142);
and U9722 (N_9722,N_7885,N_7431);
and U9723 (N_9723,N_6136,N_7056);
and U9724 (N_9724,N_6638,N_7768);
xnor U9725 (N_9725,N_6392,N_7992);
nor U9726 (N_9726,N_6158,N_7406);
or U9727 (N_9727,N_7188,N_7654);
or U9728 (N_9728,N_6407,N_7918);
or U9729 (N_9729,N_7228,N_7698);
and U9730 (N_9730,N_7268,N_6430);
nor U9731 (N_9731,N_7757,N_7309);
nand U9732 (N_9732,N_6381,N_6710);
nor U9733 (N_9733,N_7069,N_7415);
nor U9734 (N_9734,N_7672,N_7025);
and U9735 (N_9735,N_7966,N_7769);
nand U9736 (N_9736,N_7254,N_7695);
or U9737 (N_9737,N_7874,N_6201);
and U9738 (N_9738,N_6362,N_7387);
or U9739 (N_9739,N_6892,N_7835);
or U9740 (N_9740,N_7676,N_7594);
nor U9741 (N_9741,N_6492,N_7464);
and U9742 (N_9742,N_7967,N_7877);
nor U9743 (N_9743,N_7773,N_7187);
nor U9744 (N_9744,N_6740,N_7401);
or U9745 (N_9745,N_6948,N_6223);
and U9746 (N_9746,N_6416,N_7290);
nor U9747 (N_9747,N_7559,N_6180);
nor U9748 (N_9748,N_7005,N_7536);
nor U9749 (N_9749,N_7044,N_7585);
or U9750 (N_9750,N_6505,N_7093);
nor U9751 (N_9751,N_6472,N_7969);
nand U9752 (N_9752,N_7646,N_7721);
or U9753 (N_9753,N_7362,N_7349);
nand U9754 (N_9754,N_6950,N_7437);
nor U9755 (N_9755,N_7327,N_6669);
nor U9756 (N_9756,N_6909,N_7306);
or U9757 (N_9757,N_7312,N_6361);
nor U9758 (N_9758,N_6226,N_6586);
nand U9759 (N_9759,N_6489,N_6111);
nor U9760 (N_9760,N_7943,N_7080);
nor U9761 (N_9761,N_6447,N_6510);
or U9762 (N_9762,N_7344,N_6593);
nor U9763 (N_9763,N_7086,N_6230);
nor U9764 (N_9764,N_6957,N_7388);
nand U9765 (N_9765,N_6995,N_7918);
or U9766 (N_9766,N_7319,N_6516);
nor U9767 (N_9767,N_6640,N_7250);
and U9768 (N_9768,N_7492,N_7598);
or U9769 (N_9769,N_7511,N_7780);
nor U9770 (N_9770,N_7487,N_7785);
nor U9771 (N_9771,N_7826,N_7598);
nand U9772 (N_9772,N_6282,N_6716);
nor U9773 (N_9773,N_6056,N_7112);
or U9774 (N_9774,N_6006,N_6103);
nor U9775 (N_9775,N_6520,N_7793);
or U9776 (N_9776,N_6440,N_7701);
and U9777 (N_9777,N_7810,N_6749);
nor U9778 (N_9778,N_7488,N_6244);
nand U9779 (N_9779,N_6587,N_6362);
nor U9780 (N_9780,N_7238,N_6751);
and U9781 (N_9781,N_7324,N_6180);
and U9782 (N_9782,N_7386,N_6632);
or U9783 (N_9783,N_6635,N_6317);
or U9784 (N_9784,N_6221,N_6602);
nor U9785 (N_9785,N_7383,N_6948);
and U9786 (N_9786,N_6360,N_6274);
nand U9787 (N_9787,N_6846,N_6013);
xor U9788 (N_9788,N_7232,N_7261);
nand U9789 (N_9789,N_6131,N_6778);
nor U9790 (N_9790,N_7617,N_6608);
or U9791 (N_9791,N_7869,N_6416);
nand U9792 (N_9792,N_7584,N_7409);
nor U9793 (N_9793,N_6888,N_6769);
and U9794 (N_9794,N_7686,N_7954);
nand U9795 (N_9795,N_7006,N_6497);
nand U9796 (N_9796,N_7226,N_6943);
xnor U9797 (N_9797,N_6260,N_6530);
and U9798 (N_9798,N_7964,N_6614);
or U9799 (N_9799,N_7212,N_7035);
nor U9800 (N_9800,N_6798,N_7116);
nor U9801 (N_9801,N_7275,N_7204);
nor U9802 (N_9802,N_7969,N_7002);
nor U9803 (N_9803,N_7234,N_7568);
and U9804 (N_9804,N_6202,N_6895);
or U9805 (N_9805,N_7742,N_6979);
nor U9806 (N_9806,N_7764,N_6154);
or U9807 (N_9807,N_6950,N_7409);
or U9808 (N_9808,N_7653,N_7599);
nand U9809 (N_9809,N_7130,N_7121);
or U9810 (N_9810,N_7400,N_7473);
nor U9811 (N_9811,N_6508,N_7577);
nand U9812 (N_9812,N_7459,N_6270);
or U9813 (N_9813,N_7517,N_7709);
nand U9814 (N_9814,N_7033,N_6946);
nand U9815 (N_9815,N_7913,N_6616);
and U9816 (N_9816,N_6917,N_6149);
and U9817 (N_9817,N_6413,N_7183);
or U9818 (N_9818,N_7486,N_6976);
nand U9819 (N_9819,N_7007,N_7477);
nand U9820 (N_9820,N_7318,N_6784);
or U9821 (N_9821,N_7988,N_6866);
or U9822 (N_9822,N_7110,N_6543);
and U9823 (N_9823,N_7947,N_7294);
and U9824 (N_9824,N_6888,N_6422);
nor U9825 (N_9825,N_7568,N_7724);
nand U9826 (N_9826,N_6419,N_7709);
nor U9827 (N_9827,N_6234,N_7929);
nor U9828 (N_9828,N_7034,N_7925);
or U9829 (N_9829,N_6068,N_7619);
nor U9830 (N_9830,N_6783,N_7871);
nand U9831 (N_9831,N_6475,N_6408);
nand U9832 (N_9832,N_7891,N_6313);
and U9833 (N_9833,N_7987,N_7464);
nor U9834 (N_9834,N_7821,N_7583);
or U9835 (N_9835,N_7190,N_7741);
and U9836 (N_9836,N_6466,N_7509);
and U9837 (N_9837,N_6323,N_6414);
or U9838 (N_9838,N_6050,N_6489);
nor U9839 (N_9839,N_6875,N_6890);
and U9840 (N_9840,N_6308,N_7308);
or U9841 (N_9841,N_7659,N_6608);
nand U9842 (N_9842,N_7512,N_7633);
nor U9843 (N_9843,N_7017,N_6795);
and U9844 (N_9844,N_7158,N_6554);
or U9845 (N_9845,N_6699,N_6750);
or U9846 (N_9846,N_6343,N_6444);
nor U9847 (N_9847,N_6286,N_7927);
nand U9848 (N_9848,N_7411,N_7684);
nand U9849 (N_9849,N_7083,N_6205);
nand U9850 (N_9850,N_6208,N_7754);
or U9851 (N_9851,N_6964,N_7804);
nor U9852 (N_9852,N_7372,N_7607);
and U9853 (N_9853,N_7084,N_6749);
nand U9854 (N_9854,N_6834,N_6235);
nand U9855 (N_9855,N_7029,N_7032);
and U9856 (N_9856,N_6930,N_7601);
nand U9857 (N_9857,N_7241,N_6545);
and U9858 (N_9858,N_6173,N_7843);
or U9859 (N_9859,N_7371,N_6166);
nand U9860 (N_9860,N_7164,N_6083);
nor U9861 (N_9861,N_6516,N_7113);
nor U9862 (N_9862,N_7358,N_6176);
nor U9863 (N_9863,N_7074,N_6857);
or U9864 (N_9864,N_6442,N_6285);
nand U9865 (N_9865,N_6071,N_6438);
nand U9866 (N_9866,N_6121,N_6148);
nor U9867 (N_9867,N_7785,N_7815);
or U9868 (N_9868,N_6425,N_7295);
or U9869 (N_9869,N_6356,N_7278);
and U9870 (N_9870,N_6185,N_7565);
or U9871 (N_9871,N_6199,N_6497);
nand U9872 (N_9872,N_7039,N_7932);
nand U9873 (N_9873,N_7162,N_7254);
nor U9874 (N_9874,N_6173,N_6245);
nor U9875 (N_9875,N_7728,N_7606);
and U9876 (N_9876,N_6986,N_6940);
nor U9877 (N_9877,N_6273,N_7830);
nor U9878 (N_9878,N_6350,N_7113);
nor U9879 (N_9879,N_6900,N_6618);
or U9880 (N_9880,N_7693,N_6933);
nand U9881 (N_9881,N_6049,N_7240);
nor U9882 (N_9882,N_6966,N_6209);
nand U9883 (N_9883,N_6089,N_7677);
nand U9884 (N_9884,N_7527,N_6036);
or U9885 (N_9885,N_7516,N_6127);
nand U9886 (N_9886,N_6854,N_6655);
nand U9887 (N_9887,N_6402,N_6138);
nor U9888 (N_9888,N_6042,N_6473);
and U9889 (N_9889,N_6440,N_7169);
and U9890 (N_9890,N_7903,N_6420);
or U9891 (N_9891,N_7961,N_7702);
nand U9892 (N_9892,N_6264,N_6247);
and U9893 (N_9893,N_6860,N_6543);
nor U9894 (N_9894,N_7556,N_7490);
nand U9895 (N_9895,N_7309,N_7966);
or U9896 (N_9896,N_7159,N_6072);
and U9897 (N_9897,N_6231,N_6965);
or U9898 (N_9898,N_7247,N_6750);
nor U9899 (N_9899,N_7337,N_7593);
and U9900 (N_9900,N_6128,N_6310);
nand U9901 (N_9901,N_7285,N_7776);
nor U9902 (N_9902,N_7465,N_7972);
and U9903 (N_9903,N_6939,N_6560);
nor U9904 (N_9904,N_6027,N_6625);
xnor U9905 (N_9905,N_7381,N_7354);
or U9906 (N_9906,N_6004,N_6723);
or U9907 (N_9907,N_7777,N_7599);
nor U9908 (N_9908,N_6406,N_7677);
and U9909 (N_9909,N_6936,N_7936);
or U9910 (N_9910,N_7779,N_7840);
nand U9911 (N_9911,N_7401,N_7560);
or U9912 (N_9912,N_6408,N_6923);
nand U9913 (N_9913,N_6547,N_7760);
or U9914 (N_9914,N_7506,N_7276);
nand U9915 (N_9915,N_7185,N_7181);
nand U9916 (N_9916,N_6329,N_7343);
nor U9917 (N_9917,N_7526,N_7171);
nor U9918 (N_9918,N_7243,N_6364);
or U9919 (N_9919,N_7783,N_6089);
nand U9920 (N_9920,N_6598,N_6756);
nor U9921 (N_9921,N_6139,N_7329);
or U9922 (N_9922,N_6250,N_6331);
nor U9923 (N_9923,N_7806,N_7724);
or U9924 (N_9924,N_6442,N_6429);
nand U9925 (N_9925,N_7096,N_7410);
or U9926 (N_9926,N_7918,N_7278);
nand U9927 (N_9927,N_7965,N_7735);
or U9928 (N_9928,N_6581,N_6162);
nand U9929 (N_9929,N_6431,N_6022);
or U9930 (N_9930,N_7210,N_7760);
nand U9931 (N_9931,N_6726,N_6202);
nand U9932 (N_9932,N_7389,N_7120);
nand U9933 (N_9933,N_6638,N_7178);
and U9934 (N_9934,N_6554,N_7411);
nand U9935 (N_9935,N_7746,N_6225);
or U9936 (N_9936,N_7377,N_6703);
or U9937 (N_9937,N_7712,N_6314);
or U9938 (N_9938,N_7815,N_7055);
xor U9939 (N_9939,N_7574,N_7886);
nand U9940 (N_9940,N_7959,N_6632);
nor U9941 (N_9941,N_7381,N_7102);
nand U9942 (N_9942,N_6786,N_7042);
or U9943 (N_9943,N_7557,N_7103);
or U9944 (N_9944,N_6275,N_7022);
and U9945 (N_9945,N_6614,N_6490);
or U9946 (N_9946,N_7557,N_7496);
xnor U9947 (N_9947,N_6948,N_7570);
nand U9948 (N_9948,N_6843,N_6525);
nor U9949 (N_9949,N_6001,N_6387);
and U9950 (N_9950,N_6159,N_6970);
and U9951 (N_9951,N_7501,N_7766);
or U9952 (N_9952,N_6465,N_7983);
nand U9953 (N_9953,N_7133,N_6138);
or U9954 (N_9954,N_6452,N_6429);
or U9955 (N_9955,N_7072,N_7466);
nand U9956 (N_9956,N_6406,N_6491);
nand U9957 (N_9957,N_6807,N_7080);
and U9958 (N_9958,N_7220,N_7143);
or U9959 (N_9959,N_7905,N_6417);
or U9960 (N_9960,N_6120,N_7589);
nor U9961 (N_9961,N_7124,N_6684);
or U9962 (N_9962,N_7664,N_7000);
nand U9963 (N_9963,N_6366,N_6033);
nor U9964 (N_9964,N_6712,N_6204);
or U9965 (N_9965,N_6559,N_7261);
nand U9966 (N_9966,N_6049,N_6995);
and U9967 (N_9967,N_7940,N_7296);
nand U9968 (N_9968,N_7230,N_7741);
or U9969 (N_9969,N_7021,N_6055);
or U9970 (N_9970,N_6038,N_6827);
and U9971 (N_9971,N_7238,N_6890);
nand U9972 (N_9972,N_6421,N_6001);
nor U9973 (N_9973,N_7836,N_6469);
nand U9974 (N_9974,N_7635,N_6510);
or U9975 (N_9975,N_7936,N_7528);
and U9976 (N_9976,N_6932,N_6090);
or U9977 (N_9977,N_7758,N_7288);
or U9978 (N_9978,N_7180,N_6940);
nor U9979 (N_9979,N_6514,N_7102);
and U9980 (N_9980,N_7201,N_6197);
and U9981 (N_9981,N_7785,N_7598);
nor U9982 (N_9982,N_6323,N_6160);
or U9983 (N_9983,N_6783,N_7269);
nor U9984 (N_9984,N_7968,N_7956);
or U9985 (N_9985,N_7334,N_6151);
or U9986 (N_9986,N_7390,N_7443);
nor U9987 (N_9987,N_7238,N_6799);
nor U9988 (N_9988,N_7925,N_7880);
and U9989 (N_9989,N_7390,N_6877);
or U9990 (N_9990,N_6397,N_7989);
and U9991 (N_9991,N_7841,N_6261);
nor U9992 (N_9992,N_7127,N_6468);
nor U9993 (N_9993,N_7206,N_6563);
or U9994 (N_9994,N_7056,N_7875);
nand U9995 (N_9995,N_7913,N_7779);
nor U9996 (N_9996,N_6336,N_7343);
and U9997 (N_9997,N_7644,N_7246);
nand U9998 (N_9998,N_7350,N_6844);
and U9999 (N_9999,N_6353,N_7060);
and UO_0 (O_0,N_8421,N_9948);
and UO_1 (O_1,N_9819,N_9576);
nand UO_2 (O_2,N_8576,N_9324);
or UO_3 (O_3,N_9409,N_9730);
or UO_4 (O_4,N_8072,N_8363);
and UO_5 (O_5,N_8760,N_8737);
and UO_6 (O_6,N_8508,N_8387);
and UO_7 (O_7,N_8346,N_9037);
and UO_8 (O_8,N_9935,N_9284);
or UO_9 (O_9,N_9374,N_9673);
nand UO_10 (O_10,N_8726,N_9241);
nand UO_11 (O_11,N_9139,N_9053);
nand UO_12 (O_12,N_8846,N_8173);
nor UO_13 (O_13,N_8769,N_9990);
and UO_14 (O_14,N_9516,N_9445);
and UO_15 (O_15,N_9890,N_8970);
nor UO_16 (O_16,N_8233,N_8168);
or UO_17 (O_17,N_8990,N_9155);
or UO_18 (O_18,N_9862,N_9809);
or UO_19 (O_19,N_9810,N_8376);
nand UO_20 (O_20,N_8322,N_9893);
nor UO_21 (O_21,N_8592,N_9301);
or UO_22 (O_22,N_9785,N_8195);
or UO_23 (O_23,N_8086,N_9589);
or UO_24 (O_24,N_9916,N_9071);
nand UO_25 (O_25,N_9114,N_8248);
nand UO_26 (O_26,N_8748,N_8965);
nor UO_27 (O_27,N_8039,N_8773);
nor UO_28 (O_28,N_9822,N_9408);
and UO_29 (O_29,N_8669,N_9024);
and UO_30 (O_30,N_9010,N_9419);
nor UO_31 (O_31,N_8134,N_8901);
or UO_32 (O_32,N_9683,N_8619);
nor UO_33 (O_33,N_9630,N_8936);
nor UO_34 (O_34,N_9404,N_8133);
or UO_35 (O_35,N_9422,N_8780);
or UO_36 (O_36,N_9080,N_8277);
or UO_37 (O_37,N_8019,N_9031);
or UO_38 (O_38,N_9616,N_9216);
nor UO_39 (O_39,N_8577,N_8758);
and UO_40 (O_40,N_8526,N_8336);
nand UO_41 (O_41,N_9447,N_9738);
nand UO_42 (O_42,N_8550,N_8488);
and UO_43 (O_43,N_8152,N_8274);
nand UO_44 (O_44,N_9805,N_8136);
nor UO_45 (O_45,N_8492,N_8319);
nand UO_46 (O_46,N_9760,N_9944);
nor UO_47 (O_47,N_9966,N_9192);
and UO_48 (O_48,N_8715,N_8880);
nand UO_49 (O_49,N_9619,N_8243);
nand UO_50 (O_50,N_8507,N_8854);
and UO_51 (O_51,N_8660,N_9364);
or UO_52 (O_52,N_9190,N_8190);
nor UO_53 (O_53,N_8255,N_9503);
nor UO_54 (O_54,N_8128,N_8124);
or UO_55 (O_55,N_9588,N_9380);
or UO_56 (O_56,N_8501,N_9107);
and UO_57 (O_57,N_8077,N_8158);
and UO_58 (O_58,N_9117,N_9686);
or UO_59 (O_59,N_9163,N_8711);
or UO_60 (O_60,N_8410,N_8432);
and UO_61 (O_61,N_8025,N_8462);
nand UO_62 (O_62,N_9631,N_8858);
and UO_63 (O_63,N_8043,N_8533);
nor UO_64 (O_64,N_8397,N_8700);
nand UO_65 (O_65,N_8349,N_9270);
and UO_66 (O_66,N_8296,N_9933);
nand UO_67 (O_67,N_9199,N_9759);
and UO_68 (O_68,N_8157,N_9495);
or UO_69 (O_69,N_9230,N_8044);
nand UO_70 (O_70,N_9474,N_8101);
nand UO_71 (O_71,N_9318,N_9959);
or UO_72 (O_72,N_8824,N_9291);
and UO_73 (O_73,N_9109,N_9883);
and UO_74 (O_74,N_8581,N_8777);
and UO_75 (O_75,N_8436,N_9140);
nor UO_76 (O_76,N_8759,N_9855);
or UO_77 (O_77,N_9020,N_9484);
nand UO_78 (O_78,N_9652,N_8112);
nor UO_79 (O_79,N_9193,N_8254);
or UO_80 (O_80,N_9922,N_9558);
nor UO_81 (O_81,N_8151,N_9072);
and UO_82 (O_82,N_8862,N_9965);
and UO_83 (O_83,N_9793,N_9919);
nor UO_84 (O_84,N_9086,N_9650);
or UO_85 (O_85,N_9598,N_8093);
nand UO_86 (O_86,N_9055,N_8515);
xnor UO_87 (O_87,N_9359,N_8722);
nor UO_88 (O_88,N_9989,N_9223);
or UO_89 (O_89,N_9001,N_9747);
nand UO_90 (O_90,N_8915,N_9787);
or UO_91 (O_91,N_9036,N_9283);
or UO_92 (O_92,N_8107,N_8871);
and UO_93 (O_93,N_8645,N_9699);
nand UO_94 (O_94,N_9361,N_9549);
nand UO_95 (O_95,N_8247,N_8616);
or UO_96 (O_96,N_8092,N_8371);
and UO_97 (O_97,N_8536,N_8041);
nor UO_98 (O_98,N_8976,N_8940);
and UO_99 (O_99,N_8188,N_9614);
and UO_100 (O_100,N_8539,N_8182);
and UO_101 (O_101,N_8518,N_9562);
nor UO_102 (O_102,N_8042,N_8315);
nor UO_103 (O_103,N_9913,N_8078);
nand UO_104 (O_104,N_8847,N_8806);
or UO_105 (O_105,N_8015,N_9632);
nor UO_106 (O_106,N_9387,N_8008);
nand UO_107 (O_107,N_8307,N_9543);
nand UO_108 (O_108,N_9112,N_8359);
or UO_109 (O_109,N_9256,N_9519);
and UO_110 (O_110,N_9566,N_8207);
and UO_111 (O_111,N_9337,N_9836);
or UO_112 (O_112,N_9574,N_8183);
or UO_113 (O_113,N_8330,N_9911);
or UO_114 (O_114,N_9426,N_9479);
xor UO_115 (O_115,N_8540,N_9290);
nor UO_116 (O_116,N_8196,N_9537);
nor UO_117 (O_117,N_8289,N_8565);
nor UO_118 (O_118,N_9006,N_8732);
or UO_119 (O_119,N_8206,N_9377);
nand UO_120 (O_120,N_9626,N_8252);
nand UO_121 (O_121,N_9781,N_9110);
nand UO_122 (O_122,N_8447,N_8429);
or UO_123 (O_123,N_9670,N_8974);
nand UO_124 (O_124,N_8301,N_9817);
and UO_125 (O_125,N_8543,N_9949);
nor UO_126 (O_126,N_8786,N_8293);
nor UO_127 (O_127,N_8024,N_9187);
or UO_128 (O_128,N_9532,N_8351);
and UO_129 (O_129,N_8099,N_8426);
nor UO_130 (O_130,N_9804,N_8352);
or UO_131 (O_131,N_8521,N_8941);
and UO_132 (O_132,N_9698,N_9154);
nor UO_133 (O_133,N_8882,N_9127);
or UO_134 (O_134,N_8561,N_8889);
or UO_135 (O_135,N_9253,N_9400);
and UO_136 (O_136,N_8756,N_8181);
or UO_137 (O_137,N_8689,N_9635);
and UO_138 (O_138,N_8912,N_9803);
and UO_139 (O_139,N_8930,N_8412);
and UO_140 (O_140,N_8624,N_9617);
or UO_141 (O_141,N_8563,N_9482);
and UO_142 (O_142,N_8353,N_8598);
and UO_143 (O_143,N_8529,N_9688);
and UO_144 (O_144,N_8789,N_9229);
and UO_145 (O_145,N_8910,N_9525);
or UO_146 (O_146,N_8163,N_8708);
or UO_147 (O_147,N_8609,N_8762);
and UO_148 (O_148,N_8027,N_8479);
nor UO_149 (O_149,N_8291,N_9000);
nand UO_150 (O_150,N_9251,N_9884);
nand UO_151 (O_151,N_9074,N_8822);
and UO_152 (O_152,N_8164,N_8143);
or UO_153 (O_153,N_8870,N_8791);
or UO_154 (O_154,N_8551,N_8063);
nand UO_155 (O_155,N_9233,N_9603);
nor UO_156 (O_156,N_8203,N_8498);
nand UO_157 (O_157,N_8323,N_9937);
nor UO_158 (O_158,N_8810,N_9368);
nand UO_159 (O_159,N_8853,N_8053);
nor UO_160 (O_160,N_8674,N_9834);
nor UO_161 (O_161,N_8900,N_9593);
xnor UO_162 (O_162,N_8094,N_8408);
nand UO_163 (O_163,N_9932,N_9719);
nand UO_164 (O_164,N_9015,N_8909);
or UO_165 (O_165,N_9946,N_9880);
nor UO_166 (O_166,N_8931,N_8145);
xnor UO_167 (O_167,N_8682,N_8456);
nand UO_168 (O_168,N_9713,N_9395);
nand UO_169 (O_169,N_9385,N_8154);
and UO_170 (O_170,N_9048,N_9848);
and UO_171 (O_171,N_9153,N_9449);
and UO_172 (O_172,N_8090,N_8913);
nand UO_173 (O_173,N_9958,N_9552);
or UO_174 (O_174,N_8194,N_9840);
or UO_175 (O_175,N_9066,N_8985);
nand UO_176 (O_176,N_8069,N_8765);
or UO_177 (O_177,N_9026,N_8714);
nand UO_178 (O_178,N_9041,N_9999);
or UO_179 (O_179,N_9069,N_8681);
nor UO_180 (O_180,N_9583,N_8127);
nor UO_181 (O_181,N_9750,N_8055);
and UO_182 (O_182,N_9649,N_8073);
nor UO_183 (O_183,N_9797,N_8830);
nand UO_184 (O_184,N_8317,N_9826);
nor UO_185 (O_185,N_8868,N_9434);
nor UO_186 (O_186,N_9628,N_9182);
nand UO_187 (O_187,N_9300,N_9876);
or UO_188 (O_188,N_8391,N_9352);
nor UO_189 (O_189,N_8415,N_9950);
or UO_190 (O_190,N_8833,N_8744);
and UO_191 (O_191,N_8832,N_8097);
nor UO_192 (O_192,N_8013,N_9287);
nor UO_193 (O_193,N_8999,N_8485);
and UO_194 (O_194,N_9746,N_8713);
or UO_195 (O_195,N_8630,N_8360);
or UO_196 (O_196,N_9691,N_8369);
nor UO_197 (O_197,N_8724,N_8358);
nor UO_198 (O_198,N_9108,N_9396);
nor UO_199 (O_199,N_9962,N_9097);
or UO_200 (O_200,N_9240,N_9902);
or UO_201 (O_201,N_9220,N_8811);
nor UO_202 (O_202,N_9178,N_9601);
nor UO_203 (O_203,N_9172,N_9130);
and UO_204 (O_204,N_9266,N_9070);
and UO_205 (O_205,N_8819,N_9047);
nand UO_206 (O_206,N_9013,N_8220);
nor UO_207 (O_207,N_9551,N_9706);
or UO_208 (O_208,N_9701,N_9844);
nor UO_209 (O_209,N_9068,N_8299);
nor UO_210 (O_210,N_9101,N_8570);
nor UO_211 (O_211,N_8656,N_9972);
nor UO_212 (O_212,N_9378,N_8440);
or UO_213 (O_213,N_8401,N_8155);
or UO_214 (O_214,N_9038,N_9757);
and UO_215 (O_215,N_9818,N_9046);
or UO_216 (O_216,N_9025,N_9498);
or UO_217 (O_217,N_8723,N_9742);
nand UO_218 (O_218,N_8345,N_8794);
nor UO_219 (O_219,N_9232,N_9800);
nor UO_220 (O_220,N_8951,N_8281);
nand UO_221 (O_221,N_9620,N_9360);
nand UO_222 (O_222,N_9436,N_8392);
xnor UO_223 (O_223,N_9612,N_9079);
or UO_224 (O_224,N_9145,N_9005);
or UO_225 (O_225,N_8750,N_8860);
nor UO_226 (O_226,N_8694,N_9656);
and UO_227 (O_227,N_8249,N_8489);
nor UO_228 (O_228,N_8787,N_9205);
or UO_229 (O_229,N_9597,N_8100);
nand UO_230 (O_230,N_9606,N_8738);
or UO_231 (O_231,N_8239,N_8678);
or UO_232 (O_232,N_9481,N_8422);
nor UO_233 (O_233,N_8608,N_9580);
nor UO_234 (O_234,N_9162,N_8741);
and UO_235 (O_235,N_8208,N_8535);
and UO_236 (O_236,N_9263,N_8405);
and UO_237 (O_237,N_9149,N_8165);
nand UO_238 (O_238,N_8348,N_9639);
or UO_239 (O_239,N_8467,N_9638);
nor UO_240 (O_240,N_8211,N_8788);
nand UO_241 (O_241,N_9444,N_8890);
nand UO_242 (O_242,N_9823,N_8251);
nor UO_243 (O_243,N_8720,N_8218);
nor UO_244 (O_244,N_9424,N_8375);
nand UO_245 (O_245,N_8482,N_9769);
nand UO_246 (O_246,N_9717,N_8403);
or UO_247 (O_247,N_9741,N_9556);
or UO_248 (O_248,N_9973,N_9869);
or UO_249 (O_249,N_9177,N_8423);
and UO_250 (O_250,N_8464,N_9982);
nor UO_251 (O_251,N_8085,N_9390);
or UO_252 (O_252,N_8704,N_8395);
nand UO_253 (O_253,N_9100,N_8439);
and UO_254 (O_254,N_8776,N_8227);
nand UO_255 (O_255,N_8861,N_8178);
nand UO_256 (O_256,N_9217,N_8054);
or UO_257 (O_257,N_8877,N_9564);
nand UO_258 (O_258,N_9943,N_9280);
and UO_259 (O_259,N_9956,N_8059);
or UO_260 (O_260,N_8799,N_9665);
or UO_261 (O_261,N_8021,N_8591);
or UO_262 (O_262,N_8804,N_9915);
and UO_263 (O_263,N_8443,N_9347);
nand UO_264 (O_264,N_8823,N_8216);
or UO_265 (O_265,N_9329,N_9505);
and UO_266 (O_266,N_9753,N_8625);
and UO_267 (O_267,N_9144,N_9767);
nor UO_268 (O_268,N_8753,N_8751);
nand UO_269 (O_269,N_9856,N_8244);
or UO_270 (O_270,N_9092,N_8803);
and UO_271 (O_271,N_9465,N_8567);
or UO_272 (O_272,N_8434,N_8851);
and UO_273 (O_273,N_8106,N_9555);
or UO_274 (O_274,N_8884,N_9493);
and UO_275 (O_275,N_8525,N_8463);
nand UO_276 (O_276,N_9322,N_8778);
and UO_277 (O_277,N_8368,N_9923);
and UO_278 (O_278,N_8197,N_9511);
xor UO_279 (O_279,N_9295,N_8454);
or UO_280 (O_280,N_8082,N_8473);
nand UO_281 (O_281,N_8600,N_8981);
or UO_282 (O_282,N_8548,N_8933);
nand UO_283 (O_283,N_9243,N_9033);
nand UO_284 (O_284,N_9427,N_8259);
and UO_285 (O_285,N_9708,N_8691);
nor UO_286 (O_286,N_9064,N_9211);
or UO_287 (O_287,N_8643,N_9294);
and UO_288 (O_288,N_9341,N_9311);
nand UO_289 (O_289,N_8826,N_8172);
nand UO_290 (O_290,N_9860,N_9816);
nand UO_291 (O_291,N_9488,N_8506);
and UO_292 (O_292,N_8784,N_9658);
nand UO_293 (O_293,N_9039,N_8932);
or UO_294 (O_294,N_9731,N_8728);
and UO_295 (O_295,N_8505,N_9740);
nand UO_296 (O_296,N_8098,N_8111);
nor UO_297 (O_297,N_9842,N_9023);
nor UO_298 (O_298,N_9843,N_9342);
nor UO_299 (O_299,N_9866,N_9718);
nand UO_300 (O_300,N_8010,N_8657);
nand UO_301 (O_301,N_9472,N_9147);
and UO_302 (O_302,N_8560,N_8167);
nor UO_303 (O_303,N_9931,N_9248);
nor UO_304 (O_304,N_8963,N_9030);
and UO_305 (O_305,N_9567,N_8279);
nand UO_306 (O_306,N_8170,N_8272);
and UO_307 (O_307,N_8613,N_8471);
nor UO_308 (O_308,N_9271,N_9681);
or UO_309 (O_309,N_9435,N_8303);
nand UO_310 (O_310,N_9968,N_9363);
nor UO_311 (O_311,N_9514,N_9260);
or UO_312 (O_312,N_8047,N_9174);
nor UO_313 (O_313,N_8649,N_8148);
nand UO_314 (O_314,N_9779,N_8962);
or UO_315 (O_315,N_8849,N_9858);
and UO_316 (O_316,N_8316,N_9554);
nor UO_317 (O_317,N_8209,N_9573);
nand UO_318 (O_318,N_8399,N_9274);
nor UO_319 (O_319,N_9084,N_8324);
nand UO_320 (O_320,N_9045,N_9729);
and UO_321 (O_321,N_8772,N_9778);
and UO_322 (O_322,N_8215,N_9338);
and UO_323 (O_323,N_8103,N_9040);
nor UO_324 (O_324,N_9032,N_8448);
nand UO_325 (O_325,N_9736,N_8005);
or UO_326 (O_326,N_8374,N_8874);
nor UO_327 (O_327,N_9788,N_9831);
and UO_328 (O_328,N_9689,N_8400);
nand UO_329 (O_329,N_9541,N_9640);
nor UO_330 (O_330,N_9315,N_9406);
nor UO_331 (O_331,N_8840,N_9508);
nand UO_332 (O_332,N_8838,N_8364);
nor UO_333 (O_333,N_9204,N_9975);
nor UO_334 (O_334,N_9735,N_8524);
nand UO_335 (O_335,N_9924,N_8574);
nor UO_336 (O_336,N_9090,N_8528);
nor UO_337 (O_337,N_8716,N_8568);
and UO_338 (O_338,N_9119,N_9825);
nand UO_339 (O_339,N_8650,N_9325);
or UO_340 (O_340,N_9375,N_9995);
nand UO_341 (O_341,N_9540,N_8821);
or UO_342 (O_342,N_9486,N_9367);
xnor UO_343 (O_343,N_9456,N_9702);
nand UO_344 (O_344,N_8727,N_9997);
nand UO_345 (O_345,N_8084,N_9986);
or UO_346 (O_346,N_9722,N_9507);
or UO_347 (O_347,N_8096,N_9796);
nor UO_348 (O_348,N_9952,N_8622);
nor UO_349 (O_349,N_9448,N_9320);
nor UO_350 (O_350,N_9129,N_9158);
or UO_351 (O_351,N_9083,N_8420);
or UO_352 (O_352,N_8928,N_9442);
nand UO_353 (O_353,N_8068,N_9016);
or UO_354 (O_354,N_8557,N_8357);
and UO_355 (O_355,N_9469,N_8334);
nor UO_356 (O_356,N_8491,N_9586);
and UO_357 (O_357,N_8721,N_9725);
nor UO_358 (O_358,N_8888,N_8265);
or UO_359 (O_359,N_9553,N_8531);
nand UO_360 (O_360,N_8937,N_9401);
nand UO_361 (O_361,N_8636,N_9776);
nor UO_362 (O_362,N_9500,N_9238);
nor UO_363 (O_363,N_9113,N_9168);
nor UO_364 (O_364,N_9141,N_8418);
xnor UO_365 (O_365,N_8232,N_9506);
and UO_366 (O_366,N_9716,N_8419);
and UO_367 (O_367,N_8333,N_9176);
nor UO_368 (O_368,N_9389,N_8843);
or UO_369 (O_369,N_9712,N_8618);
xnor UO_370 (O_370,N_9941,N_8137);
or UO_371 (O_371,N_9350,N_8594);
nor UO_372 (O_372,N_9179,N_9415);
nor UO_373 (O_373,N_9684,N_9607);
nor UO_374 (O_374,N_8952,N_9279);
nor UO_375 (O_375,N_9136,N_9641);
nor UO_376 (O_376,N_8051,N_9700);
nand UO_377 (O_377,N_8764,N_8825);
and UO_378 (O_378,N_9403,N_8470);
or UO_379 (O_379,N_9462,N_8000);
and UO_380 (O_380,N_8327,N_8534);
nand UO_381 (O_381,N_9675,N_9160);
nand UO_382 (O_382,N_8511,N_8997);
and UO_383 (O_383,N_8661,N_9927);
and UO_384 (O_384,N_9526,N_8193);
and UO_385 (O_385,N_9061,N_9226);
or UO_386 (O_386,N_9476,N_9587);
nand UO_387 (O_387,N_9595,N_8729);
nand UO_388 (O_388,N_8413,N_9898);
and UO_389 (O_389,N_8706,N_8673);
or UO_390 (O_390,N_9653,N_9407);
and UO_391 (O_391,N_9734,N_8564);
and UO_392 (O_392,N_9200,N_8130);
and UO_393 (O_393,N_9191,N_8542);
nor UO_394 (O_394,N_9981,N_8245);
nor UO_395 (O_395,N_9739,N_9570);
or UO_396 (O_396,N_9296,N_9466);
nor UO_397 (O_397,N_8311,N_8883);
and UO_398 (O_398,N_9221,N_8646);
and UO_399 (O_399,N_8587,N_9382);
nand UO_400 (O_400,N_9875,N_8876);
or UO_401 (O_401,N_9373,N_9164);
nand UO_402 (O_402,N_8222,N_8958);
nor UO_403 (O_403,N_9728,N_9314);
or UO_404 (O_404,N_9920,N_8018);
or UO_405 (O_405,N_9116,N_8431);
nand UO_406 (O_406,N_8031,N_9930);
nor UO_407 (O_407,N_9925,N_9124);
or UO_408 (O_408,N_9726,N_9611);
nand UO_409 (O_409,N_8050,N_8983);
nand UO_410 (O_410,N_8246,N_9323);
or UO_411 (O_411,N_9398,N_9622);
or UO_412 (O_412,N_8261,N_8174);
nor UO_413 (O_413,N_9581,N_9985);
nand UO_414 (O_414,N_8497,N_8407);
and UO_415 (O_415,N_9687,N_9386);
and UO_416 (O_416,N_9335,N_9664);
nor UO_417 (O_417,N_9346,N_8873);
or UO_418 (O_418,N_9604,N_8921);
nor UO_419 (O_419,N_9544,N_9678);
and UO_420 (O_420,N_8615,N_8670);
or UO_421 (O_421,N_9692,N_9228);
nand UO_422 (O_422,N_9798,N_8703);
or UO_423 (O_423,N_9410,N_8665);
or UO_424 (O_424,N_8960,N_8852);
xor UO_425 (O_425,N_8588,N_8905);
nor UO_426 (O_426,N_8627,N_9065);
nor UO_427 (O_427,N_8026,N_8156);
nand UO_428 (O_428,N_9413,N_9623);
nand UO_429 (O_429,N_8584,N_8520);
and UO_430 (O_430,N_9646,N_8070);
xor UO_431 (O_431,N_8386,N_8979);
nand UO_432 (O_432,N_8198,N_9633);
or UO_433 (O_433,N_8309,N_8503);
and UO_434 (O_434,N_8549,N_8731);
or UO_435 (O_435,N_9710,N_9870);
nand UO_436 (O_436,N_9629,N_8035);
nor UO_437 (O_437,N_8552,N_9478);
or UO_438 (O_438,N_9018,N_8580);
and UO_439 (O_439,N_9169,N_9845);
and UO_440 (O_440,N_9402,N_9808);
nor UO_441 (O_441,N_8798,N_8828);
nor UO_442 (O_442,N_9872,N_8679);
nand UO_443 (O_443,N_9494,N_9605);
nand UO_444 (O_444,N_9326,N_8238);
or UO_445 (O_445,N_9480,N_9264);
nand UO_446 (O_446,N_9304,N_9830);
nor UO_447 (O_447,N_8064,N_8438);
nand UO_448 (O_448,N_9269,N_9207);
nand UO_449 (O_449,N_8453,N_8487);
and UO_450 (O_450,N_8340,N_8815);
nand UO_451 (O_451,N_8586,N_8801);
or UO_452 (O_452,N_8425,N_8892);
or UO_453 (O_453,N_9417,N_8867);
and UO_454 (O_454,N_8617,N_9585);
nand UO_455 (O_455,N_8411,N_9067);
nand UO_456 (O_456,N_8290,N_8257);
nor UO_457 (O_457,N_9208,N_9391);
or UO_458 (O_458,N_9874,N_8667);
nand UO_459 (O_459,N_9235,N_9520);
nand UO_460 (O_460,N_8109,N_9912);
nand UO_461 (O_461,N_8747,N_9655);
or UO_462 (O_462,N_9578,N_8445);
nor UO_463 (O_463,N_8201,N_9278);
nand UO_464 (O_464,N_9093,N_9272);
and UO_465 (O_465,N_8538,N_9381);
or UO_466 (O_466,N_8339,N_8320);
and UO_467 (O_467,N_8893,N_9019);
xnor UO_468 (O_468,N_8949,N_9483);
nand UO_469 (O_469,N_9369,N_9414);
nor UO_470 (O_470,N_8541,N_9887);
nor UO_471 (O_471,N_8475,N_9947);
nand UO_472 (O_472,N_9547,N_9321);
nor UO_473 (O_473,N_9420,N_9051);
or UO_474 (O_474,N_8335,N_8469);
and UO_475 (O_475,N_8709,N_9327);
and UO_476 (O_476,N_8262,N_8509);
nor UO_477 (O_477,N_8337,N_8476);
and UO_478 (O_478,N_8396,N_8012);
and UO_479 (O_479,N_8441,N_9859);
nand UO_480 (O_480,N_9522,N_9259);
nand UO_481 (O_481,N_9418,N_9098);
nand UO_482 (O_482,N_8088,N_9261);
and UO_483 (O_483,N_9945,N_9529);
or UO_484 (O_484,N_9237,N_8685);
nor UO_485 (O_485,N_8306,N_9076);
and UO_486 (O_486,N_8341,N_8125);
nand UO_487 (O_487,N_9954,N_9345);
nor UO_488 (O_488,N_9215,N_8023);
xor UO_489 (O_489,N_8002,N_9955);
nand UO_490 (O_490,N_9978,N_8486);
nand UO_491 (O_491,N_8342,N_9286);
and UO_492 (O_492,N_9977,N_9773);
nand UO_493 (O_493,N_9302,N_8424);
nand UO_494 (O_494,N_8835,N_9209);
and UO_495 (O_495,N_9245,N_8663);
nor UO_496 (O_496,N_8954,N_8972);
or UO_497 (O_497,N_8677,N_9443);
nand UO_498 (O_498,N_8601,N_8959);
or UO_499 (O_499,N_8260,N_8995);
or UO_500 (O_500,N_8699,N_8350);
nand UO_501 (O_501,N_9584,N_8739);
nand UO_502 (O_502,N_8554,N_9042);
nand UO_503 (O_503,N_8036,N_9732);
nand UO_504 (O_504,N_9143,N_8131);
nor UO_505 (O_505,N_8973,N_8149);
and UO_506 (O_506,N_9662,N_9636);
nor UO_507 (O_507,N_9146,N_8775);
or UO_508 (O_508,N_8304,N_9851);
and UO_509 (O_509,N_9257,N_9685);
nand UO_510 (O_510,N_8907,N_9050);
or UO_511 (O_511,N_8210,N_8820);
nor UO_512 (O_512,N_8943,N_8914);
nor UO_513 (O_513,N_8014,N_9971);
nand UO_514 (O_514,N_9907,N_8046);
or UO_515 (O_515,N_8161,N_9850);
or UO_516 (O_516,N_8944,N_9596);
nand UO_517 (O_517,N_9452,N_9827);
nor UO_518 (O_518,N_8553,N_8326);
nor UO_519 (O_519,N_9976,N_8717);
nand UO_520 (O_520,N_8675,N_8079);
or UO_521 (O_521,N_8460,N_9561);
nor UO_522 (O_522,N_9438,N_9120);
or UO_523 (O_523,N_8920,N_8795);
nor UO_524 (O_524,N_8159,N_8062);
or UO_525 (O_525,N_8637,N_9756);
nand UO_526 (O_526,N_8621,N_8466);
and UO_527 (O_527,N_8171,N_9499);
or UO_528 (O_528,N_8639,N_9060);
nand UO_529 (O_529,N_8141,N_8373);
nand UO_530 (O_530,N_9057,N_9697);
nor UO_531 (O_531,N_8771,N_8573);
and UO_532 (O_532,N_9743,N_8620);
nor UO_533 (O_533,N_9864,N_8652);
nor UO_534 (O_534,N_9458,N_9942);
or UO_535 (O_535,N_9453,N_9059);
nor UO_536 (O_536,N_8468,N_8075);
or UO_537 (O_537,N_8782,N_8927);
xor UO_538 (O_538,N_8842,N_9905);
xor UO_539 (O_539,N_8555,N_9889);
nor UO_540 (O_540,N_8225,N_8437);
nor UO_541 (O_541,N_9592,N_9393);
or UO_542 (O_542,N_9682,N_8904);
nand UO_543 (O_543,N_8923,N_9807);
nand UO_544 (O_544,N_8433,N_9674);
or UO_545 (O_545,N_9002,N_9824);
nor UO_546 (O_546,N_9085,N_8305);
nor UO_547 (O_547,N_9988,N_9334);
or UO_548 (O_548,N_9671,N_9908);
and UO_549 (O_549,N_8638,N_9461);
and UO_550 (O_550,N_8474,N_9089);
nor UO_551 (O_551,N_8066,N_8430);
and UO_552 (O_552,N_8916,N_9313);
nand UO_553 (O_553,N_8452,N_8297);
nand UO_554 (O_554,N_8402,N_9298);
and UO_555 (O_555,N_8752,N_8185);
and UO_556 (O_556,N_9470,N_9695);
nand UO_557 (O_557,N_9014,N_8120);
and UO_558 (O_558,N_9694,N_8235);
nand UO_559 (O_559,N_9195,N_9744);
or UO_560 (O_560,N_8966,N_9303);
nand UO_561 (O_561,N_8427,N_8530);
or UO_562 (O_562,N_8294,N_9276);
xnor UO_563 (O_563,N_9104,N_9615);
nor UO_564 (O_564,N_8104,N_8362);
nor UO_565 (O_565,N_8022,N_8903);
or UO_566 (O_566,N_9992,N_9600);
or UO_567 (O_567,N_8523,N_9610);
and UO_568 (O_568,N_8740,N_9096);
nor UO_569 (O_569,N_8147,N_8918);
and UO_570 (O_570,N_8734,N_9513);
and UO_571 (O_571,N_8153,N_9548);
and UO_572 (O_572,N_9571,N_8366);
nor UO_573 (O_573,N_9839,N_9181);
or UO_574 (O_574,N_9125,N_9812);
and UO_575 (O_575,N_9963,N_8857);
nand UO_576 (O_576,N_8696,N_9648);
or UO_577 (O_577,N_8271,N_8599);
or UO_578 (O_578,N_9714,N_9863);
and UO_579 (O_579,N_9349,N_8200);
nor UO_580 (O_580,N_8404,N_9009);
nand UO_581 (O_581,N_8455,N_8977);
or UO_582 (O_582,N_9878,N_8606);
nor UO_583 (O_583,N_8117,N_9703);
or UO_584 (O_584,N_8370,N_8605);
and UO_585 (O_585,N_8219,N_8545);
xor UO_586 (O_586,N_9250,N_9293);
and UO_587 (O_587,N_9669,N_8229);
nand UO_588 (O_588,N_9774,N_8325);
and UO_589 (O_589,N_8276,N_9464);
and UO_590 (O_590,N_9142,N_9316);
nor UO_591 (O_591,N_9613,N_8205);
and UO_592 (O_592,N_9161,N_8829);
nor UO_593 (O_593,N_9886,N_8917);
or UO_594 (O_594,N_9277,N_8634);
nor UO_595 (O_595,N_9721,N_8083);
and UO_596 (O_596,N_8991,N_9171);
or UO_597 (O_597,N_8633,N_8865);
or UO_598 (O_598,N_9225,N_8998);
and UO_599 (O_599,N_8268,N_9467);
or UO_600 (O_600,N_8742,N_9926);
or UO_601 (O_601,N_8283,N_8644);
nor UO_602 (O_602,N_8113,N_9151);
or UO_603 (O_603,N_8504,N_8061);
nand UO_604 (O_604,N_9213,N_8267);
and UO_605 (O_605,N_9106,N_8558);
or UO_606 (O_606,N_9940,N_8175);
or UO_607 (O_607,N_8994,N_8409);
nor UO_608 (O_608,N_9197,N_8956);
or UO_609 (O_609,N_8514,N_9659);
and UO_610 (O_610,N_8308,N_9340);
nand UO_611 (O_611,N_8365,N_9806);
nand UO_612 (O_612,N_8033,N_8802);
and UO_613 (O_613,N_9951,N_8115);
or UO_614 (O_614,N_8926,N_9813);
nor UO_615 (O_615,N_8519,N_8761);
or UO_616 (O_616,N_8595,N_9412);
or UO_617 (O_617,N_9429,N_9914);
nor UO_618 (O_618,N_8589,N_8969);
xnor UO_619 (O_619,N_9376,N_8242);
nor UO_620 (O_620,N_8382,N_9696);
or UO_621 (O_621,N_8126,N_8878);
or UO_622 (O_622,N_8692,N_9421);
nor UO_623 (O_623,N_8234,N_9786);
and UO_624 (O_624,N_8108,N_9095);
nor UO_625 (O_625,N_9579,N_8793);
nand UO_626 (O_626,N_9761,N_8680);
nor UO_627 (O_627,N_8478,N_8048);
or UO_628 (O_628,N_9255,N_8465);
or UO_629 (O_629,N_8813,N_9835);
and UO_630 (O_630,N_8338,N_9288);
or UO_631 (O_631,N_9267,N_8935);
or UO_632 (O_632,N_8416,N_9967);
nor UO_633 (O_633,N_8745,N_8578);
and UO_634 (O_634,N_9173,N_8603);
nand UO_635 (O_635,N_9425,N_8672);
nor UO_636 (O_636,N_8783,N_9437);
or UO_637 (O_637,N_8017,N_8122);
or UO_638 (O_638,N_9939,N_9964);
or UO_639 (O_639,N_8459,N_9765);
nand UO_640 (O_640,N_8864,N_8483);
and UO_641 (O_641,N_9333,N_9471);
nand UO_642 (O_642,N_8698,N_9838);
nand UO_643 (O_643,N_9910,N_8629);
and UO_644 (O_644,N_9088,N_8733);
nand UO_645 (O_645,N_9577,N_8314);
and UO_646 (O_646,N_9899,N_9441);
or UO_647 (O_647,N_8848,N_9468);
xor UO_648 (O_648,N_8458,N_8067);
nand UO_649 (O_649,N_8768,N_9133);
and UO_650 (O_650,N_8948,N_9078);
and UO_651 (O_651,N_8361,N_9974);
nand UO_652 (O_652,N_8547,N_9996);
or UO_653 (O_653,N_8354,N_8356);
nand UO_654 (O_654,N_9405,N_9432);
nor UO_655 (O_655,N_8502,N_9103);
nand UO_656 (O_656,N_8393,N_9196);
or UO_657 (O_657,N_9258,N_8179);
nand UO_658 (O_658,N_9077,N_8950);
and UO_659 (O_659,N_8398,N_9917);
and UO_660 (O_660,N_8032,N_8284);
or UO_661 (O_661,N_9938,N_8658);
nor UO_662 (O_662,N_8996,N_8797);
or UO_663 (O_663,N_8902,N_9569);
nand UO_664 (O_664,N_8390,N_8280);
and UO_665 (O_665,N_9249,N_9693);
nor UO_666 (O_666,N_8135,N_8355);
nand UO_667 (O_667,N_8705,N_8377);
or UO_668 (O_668,N_9560,N_8612);
and UO_669 (O_669,N_9820,N_9709);
nand UO_670 (O_670,N_8057,N_9663);
nand UO_671 (O_671,N_8556,N_8695);
and UO_672 (O_672,N_8500,N_9370);
nand UO_673 (O_673,N_8499,N_8767);
nor UO_674 (O_674,N_8385,N_8142);
nor UO_675 (O_675,N_9704,N_9450);
and UO_676 (O_676,N_9762,N_8648);
nand UO_677 (O_677,N_9877,N_9530);
nor UO_678 (O_678,N_8102,N_9099);
nand UO_679 (O_679,N_8004,N_8987);
nor UO_680 (O_680,N_9170,N_8285);
nor UO_681 (O_681,N_9081,N_9440);
nor UO_682 (O_682,N_9236,N_8081);
nor UO_683 (O_683,N_9459,N_9512);
or UO_684 (O_684,N_9022,N_9102);
nor UO_685 (O_685,N_8986,N_8451);
nand UO_686 (O_686,N_8110,N_8980);
and UO_687 (O_687,N_9189,N_8192);
nor UO_688 (O_688,N_8911,N_9957);
or UO_689 (O_689,N_8671,N_9501);
nor UO_690 (O_690,N_8065,N_9837);
nand UO_691 (O_691,N_9029,N_9594);
or UO_692 (O_692,N_8449,N_9156);
nand UO_693 (O_693,N_8056,N_9582);
and UO_694 (O_694,N_8632,N_9307);
nor UO_695 (O_695,N_8253,N_9539);
nor UO_696 (O_696,N_8331,N_8329);
or UO_697 (O_697,N_8831,N_9305);
nor UO_698 (O_698,N_9821,N_8312);
or UO_699 (O_699,N_9677,N_9814);
or UO_700 (O_700,N_9657,N_8095);
nor UO_701 (O_701,N_8953,N_9752);
or UO_702 (O_702,N_8076,N_9473);
nor UO_703 (O_703,N_9201,N_9904);
nor UO_704 (O_704,N_9194,N_9993);
or UO_705 (O_705,N_9536,N_8189);
or UO_706 (O_706,N_9292,N_9980);
or UO_707 (O_707,N_9772,N_9921);
or UO_708 (O_708,N_9672,N_9521);
and UO_709 (O_709,N_9185,N_8697);
and UO_710 (O_710,N_9091,N_8146);
and UO_711 (O_711,N_9841,N_8809);
nand UO_712 (O_712,N_8446,N_9004);
or UO_713 (O_713,N_8169,N_9477);
or UO_714 (O_714,N_8011,N_9538);
and UO_715 (O_715,N_9075,N_8604);
or UO_716 (O_716,N_9165,N_9795);
nor UO_717 (O_717,N_9531,N_8763);
nand UO_718 (O_718,N_8114,N_8712);
nor UO_719 (O_719,N_8805,N_9868);
or UO_720 (O_720,N_8662,N_9642);
or UO_721 (O_721,N_8684,N_8481);
nor UO_722 (O_722,N_9527,N_8544);
nand UO_723 (O_723,N_8906,N_9524);
or UO_724 (O_724,N_9897,N_9517);
and UO_725 (O_725,N_9763,N_9011);
and UO_726 (O_726,N_8480,N_9599);
nand UO_727 (O_727,N_8725,N_8812);
and UO_728 (O_728,N_9775,N_9128);
or UO_729 (O_729,N_8582,N_8919);
nand UO_730 (O_730,N_9297,N_9052);
nand UO_731 (O_731,N_8975,N_8579);
and UO_732 (O_732,N_8121,N_9126);
and UO_733 (O_733,N_8105,N_8484);
xor UO_734 (O_734,N_9043,N_8707);
nor UO_735 (O_735,N_9994,N_9309);
nor UO_736 (O_736,N_9766,N_8808);
nand UO_737 (O_737,N_8757,N_8264);
nand UO_738 (O_738,N_9265,N_8383);
nor UO_739 (O_739,N_9987,N_9854);
nand UO_740 (O_740,N_8237,N_9789);
nand UO_741 (O_741,N_8571,N_9791);
and UO_742 (O_742,N_8642,N_9273);
and UO_743 (O_743,N_8298,N_9792);
nor UO_744 (O_744,N_8001,N_9882);
nor UO_745 (O_745,N_8367,N_8347);
and UO_746 (O_746,N_8635,N_8651);
or UO_747 (O_747,N_9439,N_9829);
nor UO_748 (O_748,N_9523,N_9847);
and UO_749 (O_749,N_9206,N_9132);
and UO_750 (O_750,N_9222,N_9777);
or UO_751 (O_751,N_8258,N_9308);
or UO_752 (O_752,N_9634,N_8343);
xor UO_753 (O_753,N_8654,N_8736);
and UO_754 (O_754,N_9861,N_8160);
or UO_755 (O_755,N_8187,N_9332);
or UO_756 (O_756,N_9397,N_8749);
nand UO_757 (O_757,N_9627,N_9111);
and UO_758 (O_758,N_8886,N_8144);
nand UO_759 (O_759,N_8743,N_9184);
or UO_760 (O_760,N_9563,N_8754);
nor UO_761 (O_761,N_8686,N_9219);
nand UO_762 (O_762,N_9832,N_8814);
nor UO_763 (O_763,N_9984,N_8850);
and UO_764 (O_764,N_8040,N_9203);
nor UO_765 (O_765,N_9454,N_9485);
nand UO_766 (O_766,N_9903,N_8278);
nor UO_767 (O_767,N_9455,N_8746);
nand UO_768 (O_768,N_8428,N_9463);
nand UO_769 (O_769,N_8007,N_9063);
or UO_770 (O_770,N_9247,N_9310);
nand UO_771 (O_771,N_9644,N_8372);
and UO_772 (O_772,N_8655,N_9348);
nand UO_773 (O_773,N_9319,N_8957);
nand UO_774 (O_774,N_9159,N_9550);
nor UO_775 (O_775,N_9970,N_9661);
nor UO_776 (O_776,N_9509,N_9654);
and UO_777 (O_777,N_8701,N_9504);
or UO_778 (O_778,N_8118,N_9384);
or UO_779 (O_779,N_9007,N_8310);
or UO_780 (O_780,N_9979,N_8946);
nor UO_781 (O_781,N_9900,N_8532);
and UO_782 (O_782,N_9572,N_9166);
and UO_783 (O_783,N_8875,N_8295);
nor UO_784 (O_784,N_8461,N_9998);
or UO_785 (O_785,N_8947,N_9609);
nand UO_786 (O_786,N_9328,N_9188);
nor UO_787 (O_787,N_8908,N_8982);
nand UO_788 (O_788,N_9366,N_9515);
and UO_789 (O_789,N_9846,N_9928);
or UO_790 (O_790,N_8388,N_9351);
or UO_791 (O_791,N_8510,N_8176);
xor UO_792 (O_792,N_9833,N_9667);
or UO_793 (O_793,N_9724,N_9645);
nor UO_794 (O_794,N_8989,N_8702);
nor UO_795 (O_795,N_9991,N_9118);
or UO_796 (O_796,N_9138,N_9715);
nand UO_797 (O_797,N_8978,N_8213);
or UO_798 (O_798,N_9857,N_8730);
nand UO_799 (O_799,N_8925,N_9720);
nand UO_800 (O_800,N_9901,N_9723);
and UO_801 (O_801,N_9546,N_9637);
and UO_802 (O_802,N_8841,N_9647);
and UO_803 (O_803,N_8231,N_9799);
and UO_804 (O_804,N_9198,N_9282);
nor UO_805 (O_805,N_8770,N_9231);
or UO_806 (O_806,N_9428,N_9244);
nand UO_807 (O_807,N_8881,N_8869);
nand UO_808 (O_808,N_8597,N_9815);
or UO_809 (O_809,N_9344,N_9888);
and UO_810 (O_810,N_9285,N_8866);
nor UO_811 (O_811,N_8993,N_9497);
nor UO_812 (O_812,N_8968,N_9423);
or UO_813 (O_813,N_8191,N_9510);
and UO_814 (O_814,N_9383,N_8060);
nand UO_815 (O_815,N_9969,N_9012);
nand UO_816 (O_816,N_8300,N_8186);
and UO_817 (O_817,N_8522,N_8955);
or UO_818 (O_818,N_8517,N_8228);
or UO_819 (O_819,N_8263,N_8585);
nand UO_820 (O_820,N_8961,N_8087);
nor UO_821 (O_821,N_8045,N_8575);
nor UO_822 (O_822,N_8938,N_8816);
or UO_823 (O_823,N_9121,N_9242);
nand UO_824 (O_824,N_8929,N_9475);
nor UO_825 (O_825,N_9867,N_8282);
or UO_826 (O_826,N_8781,N_9559);
or UO_827 (O_827,N_9306,N_9056);
or UO_828 (O_828,N_9496,N_9122);
or UO_829 (O_829,N_9918,N_9749);
and UO_830 (O_830,N_9707,N_8177);
nand UO_831 (O_831,N_9894,N_8074);
or UO_832 (O_832,N_9115,N_8256);
nand UO_833 (O_833,N_9852,N_8834);
nor UO_834 (O_834,N_8344,N_9533);
and UO_835 (O_835,N_8394,N_8855);
or UO_836 (O_836,N_8332,N_8224);
or UO_837 (O_837,N_8537,N_9254);
and UO_838 (O_838,N_9355,N_8379);
or UO_839 (O_839,N_8562,N_9343);
or UO_840 (O_840,N_8049,N_8016);
and UO_841 (O_841,N_9771,N_8328);
and UO_842 (O_842,N_8626,N_9227);
nor UO_843 (O_843,N_8071,N_9105);
or UO_844 (O_844,N_9802,N_8653);
nand UO_845 (O_845,N_8596,N_8718);
and UO_846 (O_846,N_8792,N_9357);
xnor UO_847 (O_847,N_9565,N_9542);
nand UO_848 (O_848,N_8693,N_9224);
nand UO_849 (O_849,N_8292,N_8735);
nor UO_850 (O_850,N_8988,N_8992);
nor UO_851 (O_851,N_8898,N_8318);
nand UO_852 (O_852,N_9094,N_8513);
nand UO_853 (O_853,N_9021,N_9214);
or UO_854 (O_854,N_9365,N_8058);
nand UO_855 (O_855,N_9934,N_9953);
xor UO_856 (O_856,N_8647,N_8688);
nor UO_857 (O_857,N_9733,N_9281);
and UO_858 (O_858,N_9618,N_8450);
nor UO_859 (O_859,N_8559,N_8477);
nand UO_860 (O_860,N_9262,N_9073);
nand UO_861 (O_861,N_9602,N_9234);
and UO_862 (O_862,N_8683,N_8240);
nand UO_863 (O_863,N_8006,N_9148);
and UO_864 (O_864,N_9960,N_9489);
nand UO_865 (O_865,N_8628,N_9895);
or UO_866 (O_866,N_9679,N_8607);
or UO_867 (O_867,N_9909,N_8894);
or UO_868 (O_868,N_9457,N_8199);
nor UO_869 (O_869,N_8774,N_9008);
xor UO_870 (O_870,N_9252,N_9399);
and UO_871 (O_871,N_9983,N_8800);
nand UO_872 (O_872,N_8038,N_9754);
nand UO_873 (O_873,N_9885,N_9502);
or UO_874 (O_874,N_9782,N_8321);
nor UO_875 (O_875,N_8029,N_8899);
or UO_876 (O_876,N_8236,N_8659);
nor UO_877 (O_877,N_8807,N_9062);
nor UO_878 (O_878,N_8241,N_9394);
nand UO_879 (O_879,N_9534,N_9379);
nand UO_880 (O_880,N_8139,N_9054);
or UO_881 (O_881,N_9246,N_8891);
nand UO_882 (O_882,N_9210,N_8879);
and UO_883 (O_883,N_9058,N_9783);
nand UO_884 (O_884,N_9017,N_8934);
or UO_885 (O_885,N_8384,N_9331);
or UO_886 (O_886,N_8223,N_8212);
nor UO_887 (O_887,N_8273,N_8286);
nand UO_888 (O_888,N_9299,N_8872);
nand UO_889 (O_889,N_8924,N_8269);
and UO_890 (O_890,N_8818,N_9748);
and UO_891 (O_891,N_9487,N_8527);
nor UO_892 (O_892,N_8668,N_8859);
nand UO_893 (O_893,N_9590,N_9034);
and UO_894 (O_894,N_9680,N_8406);
nor UO_895 (O_895,N_8472,N_9545);
nand UO_896 (O_896,N_9768,N_9892);
xor UO_897 (O_897,N_9218,N_8710);
nand UO_898 (O_898,N_8945,N_8984);
or UO_899 (O_899,N_9660,N_9289);
nand UO_900 (O_900,N_9666,N_9676);
nand UO_901 (O_901,N_9764,N_9035);
nor UO_902 (O_902,N_9751,N_8964);
and UO_903 (O_903,N_8184,N_9575);
nor UO_904 (O_904,N_8381,N_9643);
nand UO_905 (O_905,N_8089,N_9134);
and UO_906 (O_906,N_8034,N_9568);
nand UO_907 (O_907,N_9705,N_8493);
nand UO_908 (O_908,N_8516,N_9811);
nor UO_909 (O_909,N_8414,N_9853);
and UO_910 (O_910,N_8221,N_9790);
nor UO_911 (O_911,N_9801,N_9727);
or UO_912 (O_912,N_8140,N_9131);
nor UO_913 (O_913,N_8313,N_9491);
or UO_914 (O_914,N_9336,N_9755);
nand UO_915 (O_915,N_8288,N_9906);
nand UO_916 (O_916,N_9625,N_8442);
and UO_917 (O_917,N_8610,N_8495);
or UO_918 (O_918,N_8836,N_9371);
and UO_919 (O_919,N_9873,N_9770);
and UO_920 (O_920,N_8270,N_9135);
nor UO_921 (O_921,N_9745,N_8435);
and UO_922 (O_922,N_8566,N_9608);
nand UO_923 (O_923,N_8676,N_8569);
or UO_924 (O_924,N_8895,N_9362);
or UO_925 (O_925,N_9651,N_8226);
and UO_926 (O_926,N_8942,N_9268);
and UO_927 (O_927,N_8116,N_8755);
or UO_928 (O_928,N_9896,N_9411);
nand UO_929 (O_929,N_9737,N_9891);
and UO_930 (O_930,N_9275,N_8593);
or UO_931 (O_931,N_8839,N_9150);
nand UO_932 (O_932,N_8687,N_9202);
nand UO_933 (O_933,N_8897,N_8132);
and UO_934 (O_934,N_8666,N_8150);
nor UO_935 (O_935,N_8380,N_9621);
or UO_936 (O_936,N_9431,N_8028);
or UO_937 (O_937,N_9879,N_8020);
nor UO_938 (O_938,N_9183,N_9137);
nand UO_939 (O_939,N_8827,N_8922);
and UO_940 (O_940,N_9784,N_9528);
and UO_941 (O_941,N_9317,N_9049);
or UO_942 (O_942,N_9087,N_8719);
and UO_943 (O_943,N_8631,N_8602);
nand UO_944 (O_944,N_8287,N_8546);
or UO_945 (O_945,N_8275,N_8180);
nor UO_946 (O_946,N_8572,N_8583);
or UO_947 (O_947,N_8611,N_8496);
and UO_948 (O_948,N_8845,N_9339);
nand UO_949 (O_949,N_8230,N_8266);
nand UO_950 (O_950,N_8250,N_9044);
and UO_951 (O_951,N_8214,N_9591);
or UO_952 (O_952,N_9356,N_8494);
and UO_953 (O_953,N_9849,N_8138);
and UO_954 (O_954,N_9828,N_9388);
or UO_955 (O_955,N_8785,N_9082);
and UO_956 (O_956,N_9690,N_9936);
nor UO_957 (O_957,N_9028,N_9557);
nor UO_958 (O_958,N_8030,N_8457);
nand UO_959 (O_959,N_8129,N_8166);
and UO_960 (O_960,N_8091,N_9535);
or UO_961 (O_961,N_8490,N_9392);
nor UO_962 (O_962,N_9758,N_8417);
or UO_963 (O_963,N_8590,N_9372);
or UO_964 (O_964,N_8837,N_9354);
or UO_965 (O_965,N_9518,N_9451);
nor UO_966 (O_966,N_9212,N_8389);
or UO_967 (O_967,N_9490,N_8887);
nor UO_968 (O_968,N_8119,N_9312);
and UO_969 (O_969,N_9167,N_8378);
or UO_970 (O_970,N_8885,N_8217);
nand UO_971 (O_971,N_8971,N_9492);
nand UO_972 (O_972,N_8967,N_8664);
nand UO_973 (O_973,N_8009,N_9003);
or UO_974 (O_974,N_8302,N_8512);
nand UO_975 (O_975,N_9780,N_9929);
or UO_976 (O_976,N_8844,N_8444);
nor UO_977 (O_977,N_8052,N_8939);
nand UO_978 (O_978,N_8896,N_9416);
nor UO_979 (O_979,N_8779,N_9668);
or UO_980 (O_980,N_9711,N_9353);
and UO_981 (O_981,N_8162,N_8003);
or UO_982 (O_982,N_9624,N_8796);
nor UO_983 (O_983,N_9358,N_8204);
or UO_984 (O_984,N_9180,N_8790);
or UO_985 (O_985,N_8640,N_9881);
nor UO_986 (O_986,N_9460,N_8123);
nand UO_987 (O_987,N_9871,N_9175);
or UO_988 (O_988,N_8766,N_8690);
nand UO_989 (O_989,N_9239,N_9152);
nand UO_990 (O_990,N_9186,N_9961);
nor UO_991 (O_991,N_8037,N_8856);
or UO_992 (O_992,N_9330,N_8623);
nor UO_993 (O_993,N_9433,N_8863);
nor UO_994 (O_994,N_8080,N_8202);
or UO_995 (O_995,N_8641,N_9430);
nand UO_996 (O_996,N_9027,N_9865);
and UO_997 (O_997,N_9123,N_9446);
nand UO_998 (O_998,N_8614,N_8817);
xor UO_999 (O_999,N_9157,N_9794);
and UO_1000 (O_1000,N_8582,N_9692);
or UO_1001 (O_1001,N_9860,N_9113);
nand UO_1002 (O_1002,N_8571,N_8268);
and UO_1003 (O_1003,N_8700,N_9643);
nor UO_1004 (O_1004,N_8956,N_8955);
or UO_1005 (O_1005,N_8551,N_9513);
or UO_1006 (O_1006,N_8323,N_9237);
nand UO_1007 (O_1007,N_8783,N_9860);
and UO_1008 (O_1008,N_8983,N_9533);
or UO_1009 (O_1009,N_9006,N_9777);
and UO_1010 (O_1010,N_8402,N_9460);
or UO_1011 (O_1011,N_8065,N_9113);
and UO_1012 (O_1012,N_8612,N_8668);
or UO_1013 (O_1013,N_9315,N_9410);
nand UO_1014 (O_1014,N_9153,N_9610);
and UO_1015 (O_1015,N_8014,N_9822);
and UO_1016 (O_1016,N_8084,N_9373);
xnor UO_1017 (O_1017,N_8485,N_9948);
and UO_1018 (O_1018,N_8611,N_9570);
nor UO_1019 (O_1019,N_8502,N_9437);
and UO_1020 (O_1020,N_9623,N_9198);
nand UO_1021 (O_1021,N_9252,N_9018);
nor UO_1022 (O_1022,N_9628,N_9712);
and UO_1023 (O_1023,N_8585,N_9868);
or UO_1024 (O_1024,N_8950,N_8672);
and UO_1025 (O_1025,N_8050,N_9670);
nand UO_1026 (O_1026,N_9379,N_8801);
nor UO_1027 (O_1027,N_9214,N_8781);
nand UO_1028 (O_1028,N_9918,N_9078);
nor UO_1029 (O_1029,N_9175,N_9196);
and UO_1030 (O_1030,N_9292,N_8130);
or UO_1031 (O_1031,N_8658,N_8186);
and UO_1032 (O_1032,N_8512,N_9964);
and UO_1033 (O_1033,N_9833,N_9463);
nor UO_1034 (O_1034,N_9434,N_8343);
and UO_1035 (O_1035,N_8782,N_8745);
nand UO_1036 (O_1036,N_9876,N_8915);
nand UO_1037 (O_1037,N_9211,N_8939);
nand UO_1038 (O_1038,N_9893,N_8181);
and UO_1039 (O_1039,N_9910,N_8932);
or UO_1040 (O_1040,N_8464,N_9777);
and UO_1041 (O_1041,N_8499,N_8501);
or UO_1042 (O_1042,N_9704,N_9057);
or UO_1043 (O_1043,N_9182,N_9611);
nand UO_1044 (O_1044,N_8858,N_9869);
or UO_1045 (O_1045,N_9145,N_9526);
or UO_1046 (O_1046,N_9974,N_8086);
and UO_1047 (O_1047,N_9495,N_9377);
or UO_1048 (O_1048,N_9909,N_9567);
xor UO_1049 (O_1049,N_9226,N_9491);
and UO_1050 (O_1050,N_8309,N_8949);
or UO_1051 (O_1051,N_8797,N_8605);
nand UO_1052 (O_1052,N_8613,N_9724);
nor UO_1053 (O_1053,N_8311,N_9794);
and UO_1054 (O_1054,N_9782,N_8017);
nand UO_1055 (O_1055,N_9608,N_8839);
nor UO_1056 (O_1056,N_9218,N_9969);
and UO_1057 (O_1057,N_9282,N_8241);
nor UO_1058 (O_1058,N_8043,N_9173);
or UO_1059 (O_1059,N_8473,N_9602);
nand UO_1060 (O_1060,N_9440,N_9907);
nor UO_1061 (O_1061,N_8073,N_9464);
or UO_1062 (O_1062,N_8945,N_8861);
nor UO_1063 (O_1063,N_9114,N_9025);
and UO_1064 (O_1064,N_9213,N_9816);
nand UO_1065 (O_1065,N_8972,N_8546);
nor UO_1066 (O_1066,N_9430,N_9189);
nor UO_1067 (O_1067,N_9023,N_8275);
nor UO_1068 (O_1068,N_9741,N_8473);
nor UO_1069 (O_1069,N_9586,N_8033);
nor UO_1070 (O_1070,N_9747,N_8812);
or UO_1071 (O_1071,N_9888,N_8229);
nor UO_1072 (O_1072,N_8896,N_8763);
nor UO_1073 (O_1073,N_8322,N_9434);
nand UO_1074 (O_1074,N_9578,N_8291);
nor UO_1075 (O_1075,N_8799,N_8669);
nand UO_1076 (O_1076,N_9514,N_8323);
or UO_1077 (O_1077,N_8154,N_9390);
nand UO_1078 (O_1078,N_8954,N_8401);
and UO_1079 (O_1079,N_8496,N_8770);
nand UO_1080 (O_1080,N_8697,N_8485);
or UO_1081 (O_1081,N_8232,N_8631);
nor UO_1082 (O_1082,N_9287,N_9106);
nand UO_1083 (O_1083,N_8968,N_9537);
nand UO_1084 (O_1084,N_9099,N_8157);
nor UO_1085 (O_1085,N_8385,N_9074);
and UO_1086 (O_1086,N_9734,N_8284);
or UO_1087 (O_1087,N_8369,N_9087);
nor UO_1088 (O_1088,N_8393,N_8857);
and UO_1089 (O_1089,N_8058,N_9230);
nor UO_1090 (O_1090,N_8614,N_9206);
or UO_1091 (O_1091,N_8060,N_8370);
nand UO_1092 (O_1092,N_9781,N_9840);
or UO_1093 (O_1093,N_8654,N_8953);
and UO_1094 (O_1094,N_8589,N_9144);
nand UO_1095 (O_1095,N_9369,N_8648);
nor UO_1096 (O_1096,N_8142,N_8397);
and UO_1097 (O_1097,N_8187,N_8431);
nand UO_1098 (O_1098,N_8214,N_9189);
or UO_1099 (O_1099,N_9523,N_9041);
nand UO_1100 (O_1100,N_8004,N_9030);
or UO_1101 (O_1101,N_8834,N_9238);
nand UO_1102 (O_1102,N_9992,N_8085);
or UO_1103 (O_1103,N_8925,N_8328);
nor UO_1104 (O_1104,N_9471,N_8132);
nor UO_1105 (O_1105,N_9434,N_9409);
and UO_1106 (O_1106,N_8477,N_8049);
or UO_1107 (O_1107,N_9568,N_8209);
or UO_1108 (O_1108,N_8066,N_9761);
and UO_1109 (O_1109,N_9538,N_9686);
nand UO_1110 (O_1110,N_9239,N_8165);
nand UO_1111 (O_1111,N_9046,N_9492);
or UO_1112 (O_1112,N_8295,N_9939);
nor UO_1113 (O_1113,N_8695,N_9713);
nor UO_1114 (O_1114,N_8317,N_8573);
nand UO_1115 (O_1115,N_8963,N_9675);
and UO_1116 (O_1116,N_8449,N_8272);
and UO_1117 (O_1117,N_8455,N_8373);
nor UO_1118 (O_1118,N_8470,N_8942);
nor UO_1119 (O_1119,N_9496,N_9943);
nand UO_1120 (O_1120,N_8684,N_8926);
or UO_1121 (O_1121,N_8710,N_9655);
nand UO_1122 (O_1122,N_8364,N_9713);
nor UO_1123 (O_1123,N_8061,N_8685);
or UO_1124 (O_1124,N_9918,N_8918);
nand UO_1125 (O_1125,N_9930,N_9791);
and UO_1126 (O_1126,N_8661,N_8910);
or UO_1127 (O_1127,N_8515,N_8815);
nor UO_1128 (O_1128,N_9069,N_9177);
and UO_1129 (O_1129,N_9065,N_8267);
or UO_1130 (O_1130,N_9204,N_8299);
and UO_1131 (O_1131,N_9333,N_8539);
nor UO_1132 (O_1132,N_9591,N_9012);
or UO_1133 (O_1133,N_9513,N_9958);
nor UO_1134 (O_1134,N_8925,N_8784);
and UO_1135 (O_1135,N_9206,N_9627);
xor UO_1136 (O_1136,N_8295,N_8856);
nand UO_1137 (O_1137,N_8132,N_9722);
nor UO_1138 (O_1138,N_9312,N_8191);
and UO_1139 (O_1139,N_9791,N_9504);
or UO_1140 (O_1140,N_9221,N_9441);
nand UO_1141 (O_1141,N_8584,N_9268);
nand UO_1142 (O_1142,N_9753,N_8584);
or UO_1143 (O_1143,N_9733,N_9561);
nor UO_1144 (O_1144,N_8801,N_8456);
nand UO_1145 (O_1145,N_9044,N_9088);
nand UO_1146 (O_1146,N_9223,N_9440);
nor UO_1147 (O_1147,N_8900,N_8640);
and UO_1148 (O_1148,N_9383,N_8065);
nor UO_1149 (O_1149,N_8634,N_9699);
nand UO_1150 (O_1150,N_9574,N_8265);
or UO_1151 (O_1151,N_8033,N_8567);
nand UO_1152 (O_1152,N_8500,N_8533);
and UO_1153 (O_1153,N_9472,N_8575);
and UO_1154 (O_1154,N_8117,N_8474);
nor UO_1155 (O_1155,N_8114,N_8009);
nor UO_1156 (O_1156,N_8419,N_9065);
nor UO_1157 (O_1157,N_8094,N_8169);
nor UO_1158 (O_1158,N_8356,N_8206);
and UO_1159 (O_1159,N_8192,N_8845);
and UO_1160 (O_1160,N_9101,N_8594);
or UO_1161 (O_1161,N_8661,N_8938);
nand UO_1162 (O_1162,N_8647,N_8016);
nand UO_1163 (O_1163,N_9789,N_9536);
and UO_1164 (O_1164,N_9654,N_9140);
and UO_1165 (O_1165,N_8471,N_9653);
and UO_1166 (O_1166,N_8291,N_8536);
or UO_1167 (O_1167,N_8548,N_8750);
nor UO_1168 (O_1168,N_8049,N_8612);
and UO_1169 (O_1169,N_9086,N_9497);
nor UO_1170 (O_1170,N_8246,N_8068);
and UO_1171 (O_1171,N_9361,N_9158);
and UO_1172 (O_1172,N_8304,N_9711);
or UO_1173 (O_1173,N_9736,N_9961);
nor UO_1174 (O_1174,N_9466,N_9681);
nor UO_1175 (O_1175,N_8553,N_9831);
and UO_1176 (O_1176,N_8570,N_8098);
nor UO_1177 (O_1177,N_9283,N_8749);
nor UO_1178 (O_1178,N_9673,N_8596);
and UO_1179 (O_1179,N_9826,N_8190);
nand UO_1180 (O_1180,N_8323,N_8361);
and UO_1181 (O_1181,N_8106,N_9276);
and UO_1182 (O_1182,N_9692,N_9488);
nand UO_1183 (O_1183,N_8535,N_9620);
and UO_1184 (O_1184,N_8102,N_9432);
nor UO_1185 (O_1185,N_9127,N_8385);
nor UO_1186 (O_1186,N_9498,N_9345);
and UO_1187 (O_1187,N_9016,N_9460);
or UO_1188 (O_1188,N_8436,N_8653);
or UO_1189 (O_1189,N_8249,N_8748);
or UO_1190 (O_1190,N_8817,N_8407);
nand UO_1191 (O_1191,N_9449,N_8834);
and UO_1192 (O_1192,N_8237,N_9654);
nor UO_1193 (O_1193,N_9677,N_8450);
nand UO_1194 (O_1194,N_8259,N_9649);
nor UO_1195 (O_1195,N_8136,N_9943);
and UO_1196 (O_1196,N_9452,N_8377);
nand UO_1197 (O_1197,N_8184,N_8189);
and UO_1198 (O_1198,N_8392,N_8124);
nand UO_1199 (O_1199,N_9126,N_8215);
and UO_1200 (O_1200,N_8978,N_9364);
nor UO_1201 (O_1201,N_9643,N_9457);
nand UO_1202 (O_1202,N_8228,N_9596);
and UO_1203 (O_1203,N_9192,N_9654);
or UO_1204 (O_1204,N_8283,N_8561);
nand UO_1205 (O_1205,N_8125,N_8485);
or UO_1206 (O_1206,N_9316,N_9238);
nor UO_1207 (O_1207,N_9798,N_8489);
xnor UO_1208 (O_1208,N_9938,N_8673);
and UO_1209 (O_1209,N_9515,N_9011);
and UO_1210 (O_1210,N_8935,N_8862);
and UO_1211 (O_1211,N_8997,N_8916);
nor UO_1212 (O_1212,N_9753,N_8977);
nand UO_1213 (O_1213,N_9077,N_8261);
and UO_1214 (O_1214,N_8074,N_9647);
and UO_1215 (O_1215,N_8696,N_8413);
or UO_1216 (O_1216,N_8687,N_9195);
or UO_1217 (O_1217,N_8266,N_9790);
or UO_1218 (O_1218,N_8771,N_9626);
nor UO_1219 (O_1219,N_8913,N_9306);
nand UO_1220 (O_1220,N_9647,N_9989);
nor UO_1221 (O_1221,N_9949,N_9994);
nand UO_1222 (O_1222,N_9856,N_9967);
or UO_1223 (O_1223,N_9351,N_9452);
or UO_1224 (O_1224,N_9142,N_8866);
nor UO_1225 (O_1225,N_9833,N_8437);
nand UO_1226 (O_1226,N_8979,N_8036);
and UO_1227 (O_1227,N_8380,N_9264);
nor UO_1228 (O_1228,N_8597,N_8543);
and UO_1229 (O_1229,N_8887,N_8424);
and UO_1230 (O_1230,N_9555,N_9118);
and UO_1231 (O_1231,N_9483,N_8953);
nor UO_1232 (O_1232,N_8215,N_9269);
or UO_1233 (O_1233,N_9439,N_9489);
nor UO_1234 (O_1234,N_9250,N_9964);
and UO_1235 (O_1235,N_9690,N_9938);
nor UO_1236 (O_1236,N_9472,N_8161);
and UO_1237 (O_1237,N_9490,N_9200);
or UO_1238 (O_1238,N_8428,N_8341);
nand UO_1239 (O_1239,N_9205,N_8641);
or UO_1240 (O_1240,N_9609,N_9424);
nor UO_1241 (O_1241,N_9968,N_9052);
nand UO_1242 (O_1242,N_8710,N_8381);
nand UO_1243 (O_1243,N_9940,N_9533);
or UO_1244 (O_1244,N_9911,N_9037);
or UO_1245 (O_1245,N_9263,N_8240);
and UO_1246 (O_1246,N_9091,N_9739);
nor UO_1247 (O_1247,N_8937,N_9853);
nand UO_1248 (O_1248,N_9452,N_8461);
nor UO_1249 (O_1249,N_9436,N_8406);
or UO_1250 (O_1250,N_8612,N_8116);
nand UO_1251 (O_1251,N_9209,N_9949);
or UO_1252 (O_1252,N_8408,N_8537);
nor UO_1253 (O_1253,N_8195,N_8525);
nor UO_1254 (O_1254,N_9056,N_8331);
nand UO_1255 (O_1255,N_9178,N_9237);
nor UO_1256 (O_1256,N_9462,N_9253);
nand UO_1257 (O_1257,N_8899,N_9279);
or UO_1258 (O_1258,N_9504,N_9203);
or UO_1259 (O_1259,N_9635,N_8358);
nor UO_1260 (O_1260,N_9841,N_8461);
nand UO_1261 (O_1261,N_8471,N_9827);
and UO_1262 (O_1262,N_8241,N_9387);
nand UO_1263 (O_1263,N_8021,N_9956);
nor UO_1264 (O_1264,N_8445,N_9177);
or UO_1265 (O_1265,N_9786,N_9802);
and UO_1266 (O_1266,N_8986,N_9240);
nor UO_1267 (O_1267,N_8324,N_8338);
nand UO_1268 (O_1268,N_9829,N_8040);
nor UO_1269 (O_1269,N_8487,N_8031);
nand UO_1270 (O_1270,N_9628,N_8940);
nor UO_1271 (O_1271,N_8764,N_9426);
nor UO_1272 (O_1272,N_9841,N_8351);
xnor UO_1273 (O_1273,N_8842,N_9778);
nand UO_1274 (O_1274,N_9335,N_8438);
or UO_1275 (O_1275,N_9451,N_9334);
and UO_1276 (O_1276,N_9355,N_9611);
nor UO_1277 (O_1277,N_9840,N_9237);
and UO_1278 (O_1278,N_8686,N_9741);
or UO_1279 (O_1279,N_8521,N_9306);
and UO_1280 (O_1280,N_9300,N_8028);
nor UO_1281 (O_1281,N_9716,N_9448);
and UO_1282 (O_1282,N_9517,N_9815);
nor UO_1283 (O_1283,N_8179,N_8030);
nand UO_1284 (O_1284,N_9400,N_8402);
nand UO_1285 (O_1285,N_9806,N_9921);
nand UO_1286 (O_1286,N_8154,N_8676);
or UO_1287 (O_1287,N_9284,N_8977);
or UO_1288 (O_1288,N_8914,N_9880);
and UO_1289 (O_1289,N_8596,N_9257);
or UO_1290 (O_1290,N_8929,N_8260);
nor UO_1291 (O_1291,N_8082,N_9419);
nand UO_1292 (O_1292,N_8934,N_8825);
nand UO_1293 (O_1293,N_9443,N_8652);
nor UO_1294 (O_1294,N_9861,N_9411);
nor UO_1295 (O_1295,N_9229,N_8111);
nor UO_1296 (O_1296,N_8370,N_9358);
or UO_1297 (O_1297,N_9976,N_8928);
nand UO_1298 (O_1298,N_8161,N_9964);
and UO_1299 (O_1299,N_8050,N_8910);
and UO_1300 (O_1300,N_8127,N_9281);
and UO_1301 (O_1301,N_9112,N_9491);
or UO_1302 (O_1302,N_9854,N_9781);
xnor UO_1303 (O_1303,N_9193,N_8297);
or UO_1304 (O_1304,N_9775,N_9898);
and UO_1305 (O_1305,N_9300,N_9405);
nor UO_1306 (O_1306,N_9703,N_8178);
nand UO_1307 (O_1307,N_8635,N_9919);
nand UO_1308 (O_1308,N_9797,N_9862);
nand UO_1309 (O_1309,N_8950,N_8215);
and UO_1310 (O_1310,N_9934,N_8688);
nor UO_1311 (O_1311,N_8405,N_8647);
and UO_1312 (O_1312,N_9862,N_9159);
nor UO_1313 (O_1313,N_8683,N_8603);
or UO_1314 (O_1314,N_9197,N_9206);
or UO_1315 (O_1315,N_9770,N_8778);
and UO_1316 (O_1316,N_9745,N_8416);
and UO_1317 (O_1317,N_8388,N_8315);
or UO_1318 (O_1318,N_8153,N_9775);
and UO_1319 (O_1319,N_8120,N_8845);
or UO_1320 (O_1320,N_8480,N_8046);
and UO_1321 (O_1321,N_8671,N_9968);
nor UO_1322 (O_1322,N_9244,N_9113);
and UO_1323 (O_1323,N_9925,N_9400);
and UO_1324 (O_1324,N_9936,N_8688);
and UO_1325 (O_1325,N_8577,N_8957);
or UO_1326 (O_1326,N_9896,N_8047);
nor UO_1327 (O_1327,N_9173,N_8110);
and UO_1328 (O_1328,N_9277,N_8524);
or UO_1329 (O_1329,N_8401,N_9884);
and UO_1330 (O_1330,N_9015,N_8445);
and UO_1331 (O_1331,N_9883,N_8986);
and UO_1332 (O_1332,N_8448,N_8959);
and UO_1333 (O_1333,N_8145,N_9120);
and UO_1334 (O_1334,N_9568,N_9329);
nand UO_1335 (O_1335,N_8389,N_9038);
nor UO_1336 (O_1336,N_8727,N_9215);
and UO_1337 (O_1337,N_8328,N_8408);
or UO_1338 (O_1338,N_8856,N_9471);
nand UO_1339 (O_1339,N_8600,N_9433);
nor UO_1340 (O_1340,N_8340,N_8950);
or UO_1341 (O_1341,N_8055,N_8504);
or UO_1342 (O_1342,N_9274,N_9408);
nor UO_1343 (O_1343,N_9263,N_8385);
and UO_1344 (O_1344,N_8639,N_8193);
and UO_1345 (O_1345,N_9610,N_9133);
nand UO_1346 (O_1346,N_9070,N_9075);
and UO_1347 (O_1347,N_9503,N_9006);
and UO_1348 (O_1348,N_8226,N_8383);
nand UO_1349 (O_1349,N_9947,N_8876);
or UO_1350 (O_1350,N_8109,N_9149);
nor UO_1351 (O_1351,N_9773,N_9212);
nor UO_1352 (O_1352,N_8108,N_9147);
nor UO_1353 (O_1353,N_8929,N_8371);
or UO_1354 (O_1354,N_8141,N_9158);
nand UO_1355 (O_1355,N_8193,N_8435);
nor UO_1356 (O_1356,N_9390,N_8203);
nand UO_1357 (O_1357,N_8267,N_9936);
or UO_1358 (O_1358,N_9613,N_9668);
nor UO_1359 (O_1359,N_9645,N_9846);
or UO_1360 (O_1360,N_8780,N_8344);
nor UO_1361 (O_1361,N_9454,N_9143);
or UO_1362 (O_1362,N_9188,N_8553);
or UO_1363 (O_1363,N_9549,N_9770);
nand UO_1364 (O_1364,N_9445,N_9596);
and UO_1365 (O_1365,N_8246,N_9358);
or UO_1366 (O_1366,N_9369,N_8773);
nor UO_1367 (O_1367,N_9322,N_8411);
and UO_1368 (O_1368,N_9401,N_9866);
or UO_1369 (O_1369,N_9687,N_9397);
and UO_1370 (O_1370,N_8590,N_9987);
and UO_1371 (O_1371,N_9888,N_9025);
nor UO_1372 (O_1372,N_9115,N_9183);
and UO_1373 (O_1373,N_8769,N_9750);
or UO_1374 (O_1374,N_9751,N_9299);
nand UO_1375 (O_1375,N_8505,N_8412);
or UO_1376 (O_1376,N_9342,N_9117);
nor UO_1377 (O_1377,N_8443,N_8168);
and UO_1378 (O_1378,N_8771,N_9561);
nand UO_1379 (O_1379,N_9841,N_9314);
nand UO_1380 (O_1380,N_8949,N_9871);
nor UO_1381 (O_1381,N_8022,N_9815);
nand UO_1382 (O_1382,N_8905,N_9845);
nor UO_1383 (O_1383,N_8562,N_9185);
or UO_1384 (O_1384,N_9990,N_8028);
nand UO_1385 (O_1385,N_9354,N_9932);
or UO_1386 (O_1386,N_8411,N_9169);
nand UO_1387 (O_1387,N_9912,N_8009);
nor UO_1388 (O_1388,N_9197,N_9802);
nand UO_1389 (O_1389,N_8657,N_8421);
and UO_1390 (O_1390,N_9620,N_9098);
and UO_1391 (O_1391,N_8371,N_9212);
nor UO_1392 (O_1392,N_9863,N_8139);
nand UO_1393 (O_1393,N_8721,N_9890);
nor UO_1394 (O_1394,N_8875,N_9220);
and UO_1395 (O_1395,N_8586,N_8998);
or UO_1396 (O_1396,N_8158,N_8421);
and UO_1397 (O_1397,N_8524,N_8311);
or UO_1398 (O_1398,N_9938,N_9748);
and UO_1399 (O_1399,N_8748,N_9287);
or UO_1400 (O_1400,N_9650,N_8032);
nor UO_1401 (O_1401,N_9019,N_8007);
nor UO_1402 (O_1402,N_8016,N_8525);
nand UO_1403 (O_1403,N_9234,N_8726);
and UO_1404 (O_1404,N_8174,N_8094);
or UO_1405 (O_1405,N_9685,N_8190);
nor UO_1406 (O_1406,N_8134,N_9128);
and UO_1407 (O_1407,N_8760,N_9505);
or UO_1408 (O_1408,N_8782,N_9408);
nand UO_1409 (O_1409,N_9194,N_8647);
or UO_1410 (O_1410,N_8781,N_9710);
and UO_1411 (O_1411,N_9536,N_9147);
or UO_1412 (O_1412,N_8672,N_8970);
nand UO_1413 (O_1413,N_8376,N_8878);
nor UO_1414 (O_1414,N_9702,N_9148);
or UO_1415 (O_1415,N_9167,N_8391);
nor UO_1416 (O_1416,N_9189,N_9536);
nor UO_1417 (O_1417,N_8163,N_8646);
nand UO_1418 (O_1418,N_8537,N_9865);
and UO_1419 (O_1419,N_9788,N_8966);
nor UO_1420 (O_1420,N_8646,N_8144);
nand UO_1421 (O_1421,N_9773,N_8296);
nand UO_1422 (O_1422,N_9967,N_8827);
nor UO_1423 (O_1423,N_9242,N_9231);
nor UO_1424 (O_1424,N_8757,N_9782);
or UO_1425 (O_1425,N_8859,N_8903);
nor UO_1426 (O_1426,N_8449,N_8722);
nor UO_1427 (O_1427,N_9344,N_9458);
and UO_1428 (O_1428,N_8424,N_9156);
or UO_1429 (O_1429,N_9482,N_9057);
and UO_1430 (O_1430,N_8144,N_8770);
nand UO_1431 (O_1431,N_9959,N_8547);
or UO_1432 (O_1432,N_8383,N_9563);
nor UO_1433 (O_1433,N_8055,N_9551);
nand UO_1434 (O_1434,N_8132,N_8367);
nor UO_1435 (O_1435,N_9642,N_9826);
and UO_1436 (O_1436,N_8097,N_8635);
and UO_1437 (O_1437,N_8194,N_8559);
nor UO_1438 (O_1438,N_8196,N_8280);
or UO_1439 (O_1439,N_9340,N_8196);
nand UO_1440 (O_1440,N_9137,N_8653);
and UO_1441 (O_1441,N_8770,N_8482);
or UO_1442 (O_1442,N_9796,N_8856);
or UO_1443 (O_1443,N_9389,N_8159);
or UO_1444 (O_1444,N_9621,N_9439);
or UO_1445 (O_1445,N_9807,N_9816);
or UO_1446 (O_1446,N_8405,N_8691);
and UO_1447 (O_1447,N_9749,N_9278);
and UO_1448 (O_1448,N_9571,N_8868);
and UO_1449 (O_1449,N_8794,N_8968);
nor UO_1450 (O_1450,N_8204,N_8665);
and UO_1451 (O_1451,N_9784,N_8296);
and UO_1452 (O_1452,N_8564,N_8871);
and UO_1453 (O_1453,N_9846,N_8087);
nor UO_1454 (O_1454,N_9685,N_9135);
nor UO_1455 (O_1455,N_9910,N_9967);
nand UO_1456 (O_1456,N_9315,N_8380);
or UO_1457 (O_1457,N_9613,N_9940);
nor UO_1458 (O_1458,N_9873,N_9312);
and UO_1459 (O_1459,N_8530,N_9107);
or UO_1460 (O_1460,N_9822,N_8252);
nor UO_1461 (O_1461,N_8856,N_9122);
and UO_1462 (O_1462,N_8027,N_8341);
and UO_1463 (O_1463,N_8924,N_9360);
or UO_1464 (O_1464,N_8230,N_9662);
and UO_1465 (O_1465,N_8159,N_8775);
nand UO_1466 (O_1466,N_8231,N_8809);
nand UO_1467 (O_1467,N_9214,N_9089);
nand UO_1468 (O_1468,N_9478,N_8485);
and UO_1469 (O_1469,N_8421,N_9928);
nor UO_1470 (O_1470,N_9089,N_8091);
xnor UO_1471 (O_1471,N_8674,N_9238);
nor UO_1472 (O_1472,N_9428,N_8586);
and UO_1473 (O_1473,N_9966,N_8630);
nand UO_1474 (O_1474,N_9990,N_9049);
nand UO_1475 (O_1475,N_8890,N_9162);
nand UO_1476 (O_1476,N_9638,N_9191);
and UO_1477 (O_1477,N_8834,N_9873);
or UO_1478 (O_1478,N_9596,N_9729);
nor UO_1479 (O_1479,N_8188,N_9098);
and UO_1480 (O_1480,N_8115,N_8686);
or UO_1481 (O_1481,N_8964,N_8455);
nand UO_1482 (O_1482,N_9626,N_9273);
or UO_1483 (O_1483,N_9138,N_9043);
or UO_1484 (O_1484,N_9180,N_9124);
nor UO_1485 (O_1485,N_9810,N_8933);
nor UO_1486 (O_1486,N_8440,N_8517);
nand UO_1487 (O_1487,N_8001,N_9096);
or UO_1488 (O_1488,N_8797,N_9137);
and UO_1489 (O_1489,N_8182,N_9014);
or UO_1490 (O_1490,N_9362,N_8796);
or UO_1491 (O_1491,N_8533,N_8536);
nor UO_1492 (O_1492,N_8925,N_8368);
nor UO_1493 (O_1493,N_9928,N_8574);
or UO_1494 (O_1494,N_9182,N_8038);
nor UO_1495 (O_1495,N_9819,N_8230);
nor UO_1496 (O_1496,N_9234,N_9389);
and UO_1497 (O_1497,N_8988,N_8982);
nor UO_1498 (O_1498,N_9309,N_9549);
nor UO_1499 (O_1499,N_8557,N_9641);
endmodule