module basic_1000_10000_1500_20_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_146,In_740);
nor U1 (N_1,In_711,In_344);
nor U2 (N_2,In_935,In_123);
xnor U3 (N_3,In_939,In_14);
nand U4 (N_4,In_167,In_696);
nor U5 (N_5,In_235,In_495);
and U6 (N_6,In_483,In_591);
nand U7 (N_7,In_117,In_868);
nor U8 (N_8,In_583,In_21);
or U9 (N_9,In_330,In_38);
nand U10 (N_10,In_76,In_16);
xnor U11 (N_11,In_357,In_378);
nand U12 (N_12,In_527,In_165);
and U13 (N_13,In_744,In_534);
nor U14 (N_14,In_305,In_862);
and U15 (N_15,In_962,In_452);
or U16 (N_16,In_30,In_810);
nor U17 (N_17,In_215,In_408);
or U18 (N_18,In_951,In_808);
or U19 (N_19,In_660,In_647);
and U20 (N_20,In_365,In_645);
or U21 (N_21,In_875,In_648);
xnor U22 (N_22,In_861,In_331);
xnor U23 (N_23,In_888,In_263);
nand U24 (N_24,In_33,In_23);
nor U25 (N_25,In_960,In_796);
xnor U26 (N_26,In_34,In_335);
and U27 (N_27,In_746,In_289);
nor U28 (N_28,In_61,In_688);
or U29 (N_29,In_659,In_946);
or U30 (N_30,In_689,In_639);
nor U31 (N_31,In_731,In_652);
nor U32 (N_32,In_972,In_109);
xnor U33 (N_33,In_158,In_499);
and U34 (N_34,In_20,In_773);
and U35 (N_35,In_572,In_280);
and U36 (N_36,In_870,In_363);
xor U37 (N_37,In_260,In_716);
or U38 (N_38,In_551,In_249);
or U39 (N_39,In_36,In_269);
xor U40 (N_40,In_677,In_785);
nand U41 (N_41,In_928,In_427);
and U42 (N_42,In_826,In_850);
or U43 (N_43,In_374,In_518);
and U44 (N_44,In_292,In_623);
nor U45 (N_45,In_754,In_206);
and U46 (N_46,In_39,In_461);
and U47 (N_47,In_113,In_291);
nor U48 (N_48,In_863,In_601);
xnor U49 (N_49,In_224,In_899);
xor U50 (N_50,In_787,In_662);
nand U51 (N_51,In_341,In_661);
and U52 (N_52,In_979,In_144);
or U53 (N_53,In_790,In_306);
and U54 (N_54,In_467,In_223);
nor U55 (N_55,In_838,In_369);
nor U56 (N_56,In_135,In_811);
nor U57 (N_57,In_548,In_698);
nand U58 (N_58,In_4,In_122);
or U59 (N_59,In_567,In_610);
nor U60 (N_60,In_388,In_431);
and U61 (N_61,In_99,In_470);
or U62 (N_62,In_926,In_320);
or U63 (N_63,In_493,In_697);
and U64 (N_64,In_90,In_817);
and U65 (N_65,In_471,In_839);
or U66 (N_66,In_624,In_103);
nand U67 (N_67,In_575,In_799);
and U68 (N_68,In_65,In_613);
nor U69 (N_69,In_789,In_555);
xnor U70 (N_70,In_699,In_145);
and U71 (N_71,In_425,In_856);
nand U72 (N_72,In_830,In_89);
nor U73 (N_73,In_924,In_867);
and U74 (N_74,In_56,In_426);
nand U75 (N_75,In_469,In_98);
nand U76 (N_76,In_506,In_675);
nand U77 (N_77,In_514,In_152);
nand U78 (N_78,In_190,In_18);
xor U79 (N_79,In_543,In_642);
nor U80 (N_80,In_195,In_929);
and U81 (N_81,In_170,In_42);
and U82 (N_82,In_406,In_321);
nor U83 (N_83,In_756,In_748);
and U84 (N_84,In_893,In_304);
xor U85 (N_85,In_142,In_912);
nor U86 (N_86,In_442,In_398);
nand U87 (N_87,In_214,In_156);
nor U88 (N_88,In_614,In_159);
or U89 (N_89,In_164,In_261);
nor U90 (N_90,In_553,In_405);
nand U91 (N_91,In_456,In_719);
and U92 (N_92,In_539,In_582);
nor U93 (N_93,In_668,In_718);
nor U94 (N_94,In_255,In_332);
or U95 (N_95,In_735,In_457);
or U96 (N_96,In_940,In_581);
and U97 (N_97,In_869,In_997);
nand U98 (N_98,In_161,In_995);
or U99 (N_99,In_941,In_47);
nand U100 (N_100,In_307,In_294);
or U101 (N_101,In_737,In_447);
or U102 (N_102,In_881,In_965);
nor U103 (N_103,In_745,In_252);
xor U104 (N_104,In_732,In_903);
and U105 (N_105,In_368,In_410);
xnor U106 (N_106,In_636,In_397);
xnor U107 (N_107,In_72,In_772);
and U108 (N_108,In_890,In_829);
and U109 (N_109,In_742,In_999);
and U110 (N_110,In_638,In_905);
and U111 (N_111,In_723,In_356);
nand U112 (N_112,In_919,In_713);
nand U113 (N_113,In_379,In_312);
or U114 (N_114,In_600,In_88);
nor U115 (N_115,In_812,In_706);
nand U116 (N_116,In_664,In_492);
nand U117 (N_117,In_372,In_24);
nand U118 (N_118,In_414,In_532);
or U119 (N_119,In_181,In_377);
and U120 (N_120,In_651,In_632);
or U121 (N_121,In_12,In_542);
nor U122 (N_122,In_262,In_690);
nor U123 (N_123,In_464,In_107);
nand U124 (N_124,In_878,In_104);
and U125 (N_125,In_818,In_900);
or U126 (N_126,In_857,In_412);
and U127 (N_127,In_348,In_409);
or U128 (N_128,In_315,In_340);
xnor U129 (N_129,In_91,In_174);
or U130 (N_130,In_399,In_526);
or U131 (N_131,In_157,In_546);
and U132 (N_132,In_803,In_679);
nand U133 (N_133,In_653,In_561);
and U134 (N_134,In_512,In_820);
nor U135 (N_135,In_445,In_239);
or U136 (N_136,In_982,In_694);
or U137 (N_137,In_43,In_212);
and U138 (N_138,In_242,In_956);
or U139 (N_139,In_80,In_10);
xor U140 (N_140,In_500,In_26);
nand U141 (N_141,In_57,In_504);
nand U142 (N_142,In_448,In_992);
xor U143 (N_143,In_937,In_271);
xor U144 (N_144,In_84,In_957);
nor U145 (N_145,In_488,In_188);
and U146 (N_146,In_859,In_436);
nand U147 (N_147,In_138,In_895);
and U148 (N_148,In_333,In_686);
or U149 (N_149,In_665,In_392);
or U150 (N_150,In_337,In_288);
xnor U151 (N_151,In_743,In_133);
nand U152 (N_152,In_360,In_684);
or U153 (N_153,In_120,In_715);
nand U154 (N_154,In_259,In_631);
nor U155 (N_155,In_886,In_316);
and U156 (N_156,In_703,In_116);
and U157 (N_157,In_906,In_173);
xor U158 (N_158,In_130,In_588);
and U159 (N_159,In_32,In_955);
nor U160 (N_160,In_83,In_626);
and U161 (N_161,In_513,In_967);
nand U162 (N_162,In_359,In_840);
nand U163 (N_163,In_299,In_343);
nor U164 (N_164,In_5,In_871);
or U165 (N_165,In_481,In_205);
and U166 (N_166,In_666,In_761);
nor U167 (N_167,In_282,In_550);
nor U168 (N_168,In_669,In_184);
xnor U169 (N_169,In_336,In_44);
or U170 (N_170,In_792,In_250);
nand U171 (N_171,In_615,In_275);
nand U172 (N_172,In_231,In_667);
xor U173 (N_173,In_189,In_437);
or U174 (N_174,In_3,In_247);
nor U175 (N_175,In_177,In_202);
nor U176 (N_176,In_420,In_396);
xnor U177 (N_177,In_450,In_355);
and U178 (N_178,In_914,In_149);
or U179 (N_179,In_938,In_864);
and U180 (N_180,In_927,In_185);
nand U181 (N_181,In_986,In_930);
xor U182 (N_182,In_63,In_860);
or U183 (N_183,In_465,In_423);
or U184 (N_184,In_272,In_303);
and U185 (N_185,In_768,In_961);
or U186 (N_186,In_137,In_942);
xnor U187 (N_187,In_324,In_503);
nor U188 (N_188,In_1,In_809);
nor U189 (N_189,In_484,In_650);
nor U190 (N_190,In_97,In_166);
or U191 (N_191,In_455,In_563);
and U192 (N_192,In_644,In_987);
nand U193 (N_193,In_580,In_883);
xnor U194 (N_194,In_985,In_367);
or U195 (N_195,In_314,In_449);
or U196 (N_196,In_676,In_201);
nand U197 (N_197,In_576,In_920);
nor U198 (N_198,In_150,In_602);
and U199 (N_199,In_317,In_0);
nor U200 (N_200,In_53,In_558);
nand U201 (N_201,In_27,In_508);
nor U202 (N_202,In_106,In_620);
or U203 (N_203,In_727,In_918);
or U204 (N_204,In_48,In_805);
and U205 (N_205,In_371,In_521);
nor U206 (N_206,In_384,In_963);
nand U207 (N_207,In_435,In_362);
nor U208 (N_208,In_110,In_973);
and U209 (N_209,In_901,In_898);
nor U210 (N_210,In_326,In_778);
or U211 (N_211,In_954,In_519);
nand U212 (N_212,In_605,In_846);
and U213 (N_213,In_510,In_277);
or U214 (N_214,In_329,In_169);
nor U215 (N_215,In_621,In_788);
nand U216 (N_216,In_739,In_976);
nand U217 (N_217,In_441,In_760);
or U218 (N_218,In_25,In_627);
nor U219 (N_219,In_628,In_227);
and U220 (N_220,In_276,In_108);
nor U221 (N_221,In_222,In_385);
or U222 (N_222,In_708,In_656);
or U223 (N_223,In_6,In_832);
or U224 (N_224,In_172,In_411);
nor U225 (N_225,In_487,In_700);
nor U226 (N_226,In_351,In_168);
nand U227 (N_227,In_894,In_253);
and U228 (N_228,In_234,In_729);
nand U229 (N_229,In_619,In_295);
nand U230 (N_230,In_264,In_124);
and U231 (N_231,In_948,In_78);
and U232 (N_232,In_328,In_489);
or U233 (N_233,In_641,In_528);
and U234 (N_234,In_118,In_153);
nand U235 (N_235,In_834,In_682);
nand U236 (N_236,In_203,In_180);
nor U237 (N_237,In_350,In_643);
or U238 (N_238,In_854,In_775);
and U239 (N_239,In_238,In_257);
nor U240 (N_240,In_889,In_390);
nand U241 (N_241,In_964,In_474);
and U242 (N_242,In_759,In_815);
and U243 (N_243,In_556,In_485);
or U244 (N_244,In_183,In_453);
or U245 (N_245,In_70,In_523);
or U246 (N_246,In_244,In_728);
xor U247 (N_247,In_907,In_592);
or U248 (N_248,In_625,In_687);
nand U249 (N_249,In_611,In_609);
xor U250 (N_250,In_278,In_428);
and U251 (N_251,In_251,In_128);
nor U252 (N_252,In_313,In_767);
nor U253 (N_253,In_95,In_801);
or U254 (N_254,In_421,In_240);
nand U255 (N_255,In_115,In_349);
nor U256 (N_256,In_7,In_584);
nand U257 (N_257,In_463,In_755);
nor U258 (N_258,In_52,In_389);
or U259 (N_259,In_917,In_670);
and U260 (N_260,In_454,In_836);
nor U261 (N_261,In_717,In_994);
nor U262 (N_262,In_593,In_217);
nand U263 (N_263,In_931,In_400);
nor U264 (N_264,In_87,In_594);
nand U265 (N_265,In_496,In_245);
or U266 (N_266,In_419,In_640);
nand U267 (N_267,In_66,In_13);
and U268 (N_268,In_798,In_874);
or U269 (N_269,In_258,In_909);
nand U270 (N_270,In_568,In_701);
nor U271 (N_271,In_725,In_286);
xnor U272 (N_272,In_816,In_629);
and U273 (N_273,In_978,In_139);
nand U274 (N_274,In_129,In_191);
or U275 (N_275,In_779,In_8);
and U276 (N_276,In_843,In_923);
nand U277 (N_277,In_771,In_204);
and U278 (N_278,In_475,In_800);
nand U279 (N_279,In_327,In_765);
nand U280 (N_280,In_570,In_422);
and U281 (N_281,In_111,In_85);
or U282 (N_282,In_193,In_216);
nand U283 (N_283,In_179,In_134);
and U284 (N_284,In_9,In_733);
nor U285 (N_285,In_589,In_402);
nor U286 (N_286,In_762,In_678);
nand U287 (N_287,In_19,In_763);
and U288 (N_288,In_552,In_199);
or U289 (N_289,In_969,In_37);
nor U290 (N_290,In_444,In_777);
or U291 (N_291,In_221,In_430);
or U292 (N_292,In_352,In_807);
or U293 (N_293,In_683,In_579);
xor U294 (N_294,In_908,In_380);
nor U295 (N_295,In_608,In_657);
and U296 (N_296,In_387,In_462);
nand U297 (N_297,In_71,In_910);
xor U298 (N_298,In_571,In_975);
nand U299 (N_299,In_925,In_171);
or U300 (N_300,In_322,In_607);
nand U301 (N_301,In_947,In_491);
or U302 (N_302,In_62,In_822);
nand U303 (N_303,In_695,In_301);
or U304 (N_304,In_383,In_58);
nand U305 (N_305,In_366,In_538);
and U306 (N_306,In_218,In_851);
and U307 (N_307,In_712,In_902);
nor U308 (N_308,In_49,In_692);
and U309 (N_309,In_738,In_270);
or U310 (N_310,In_966,In_891);
nor U311 (N_311,In_557,In_952);
nor U312 (N_312,In_599,In_560);
or U313 (N_313,In_848,In_604);
and U314 (N_314,In_782,In_182);
or U315 (N_315,In_776,In_780);
or U316 (N_316,In_793,In_46);
and U317 (N_317,In_502,In_681);
and U318 (N_318,In_101,In_287);
and U319 (N_319,In_254,In_934);
or U320 (N_320,In_824,In_382);
or U321 (N_321,In_691,In_443);
nand U322 (N_322,In_75,In_418);
xnor U323 (N_323,In_598,In_198);
or U324 (N_324,In_59,In_364);
nor U325 (N_325,In_279,In_154);
nand U326 (N_326,In_766,In_77);
nor U327 (N_327,In_837,In_845);
nand U328 (N_328,In_415,In_79);
or U329 (N_329,In_17,In_35);
and U330 (N_330,In_451,In_882);
nor U331 (N_331,In_825,In_424);
nor U332 (N_332,In_509,In_459);
xor U333 (N_333,In_578,In_268);
nand U334 (N_334,In_724,In_704);
and U335 (N_335,In_232,In_119);
or U336 (N_336,In_64,In_554);
nand U337 (N_337,In_143,In_220);
nand U338 (N_338,In_308,In_273);
xnor U339 (N_339,In_597,In_998);
nand U340 (N_340,In_403,In_633);
nand U341 (N_341,In_354,In_866);
or U342 (N_342,In_841,In_347);
nor U343 (N_343,In_786,In_750);
nand U344 (N_344,In_769,In_884);
nor U345 (N_345,In_617,In_281);
nand U346 (N_346,In_540,In_702);
and U347 (N_347,In_865,In_847);
and U348 (N_348,In_635,In_827);
nor U349 (N_349,In_873,In_968);
nand U350 (N_350,In_243,In_515);
nand U351 (N_351,In_720,In_933);
or U352 (N_352,In_256,In_194);
nor U353 (N_353,In_595,In_187);
or U354 (N_354,In_603,In_311);
or U355 (N_355,In_705,In_783);
nand U356 (N_356,In_569,In_285);
xor U357 (N_357,In_877,In_213);
or U358 (N_358,In_516,In_823);
and U359 (N_359,In_974,In_15);
and U360 (N_360,In_69,In_86);
or U361 (N_361,In_94,In_752);
xnor U362 (N_362,In_634,In_842);
nand U363 (N_363,In_93,In_674);
nor U364 (N_364,In_784,In_274);
and U365 (N_365,In_228,In_693);
and U366 (N_366,In_490,In_28);
or U367 (N_367,In_612,In_980);
nand U368 (N_368,In_114,In_233);
or U369 (N_369,In_585,In_429);
and U370 (N_370,In_524,In_334);
nand U371 (N_371,In_105,In_791);
nand U372 (N_372,In_844,In_208);
nor U373 (N_373,In_297,In_781);
nand U374 (N_374,In_916,In_804);
nand U375 (N_375,In_440,In_741);
nand U376 (N_376,In_92,In_872);
and U377 (N_377,In_479,In_544);
nor U378 (N_378,In_573,In_988);
or U379 (N_379,In_685,In_977);
xor U380 (N_380,In_125,In_186);
nor U381 (N_381,In_525,In_658);
and U382 (N_382,In_749,In_813);
or U383 (N_383,In_22,In_541);
and U384 (N_384,In_505,In_432);
or U385 (N_385,In_932,In_310);
xor U386 (N_386,In_229,In_112);
and U387 (N_387,In_394,In_82);
and U388 (N_388,In_753,In_672);
and U389 (N_389,In_529,In_821);
xnor U390 (N_390,In_226,In_849);
or U391 (N_391,In_913,In_858);
and U392 (N_392,In_950,In_473);
and U393 (N_393,In_345,In_880);
nor U394 (N_394,In_757,In_852);
xnor U395 (N_395,In_989,In_879);
nand U396 (N_396,In_819,In_163);
nand U397 (N_397,In_339,In_943);
or U398 (N_398,In_81,In_559);
or U399 (N_399,In_802,In_407);
and U400 (N_400,In_160,In_68);
xnor U401 (N_401,In_774,In_530);
nand U402 (N_402,In_707,In_155);
nor U403 (N_403,In_806,In_438);
or U404 (N_404,In_478,In_547);
nand U405 (N_405,In_885,In_209);
and U406 (N_406,In_971,In_549);
nand U407 (N_407,In_795,In_897);
or U408 (N_408,In_637,In_751);
nand U409 (N_409,In_562,In_590);
nor U410 (N_410,In_480,In_51);
and U411 (N_411,In_248,In_486);
nor U412 (N_412,In_545,In_892);
nand U413 (N_413,In_655,In_266);
nand U414 (N_414,In_2,In_853);
nor U415 (N_415,In_358,In_482);
nand U416 (N_416,In_855,In_439);
xnor U417 (N_417,In_325,In_574);
xor U418 (N_418,In_293,In_833);
nor U419 (N_419,In_680,In_141);
or U420 (N_420,In_835,In_498);
and U421 (N_421,In_586,In_446);
nor U422 (N_422,In_646,In_671);
nor U423 (N_423,In_323,In_507);
or U424 (N_424,In_45,In_953);
nand U425 (N_425,In_151,In_225);
nand U426 (N_426,In_472,In_136);
or U427 (N_427,In_981,In_814);
and U428 (N_428,In_54,In_60);
and U429 (N_429,In_577,In_494);
or U430 (N_430,In_346,In_433);
nor U431 (N_431,In_606,In_132);
nand U432 (N_432,In_921,In_175);
nand U433 (N_433,In_40,In_797);
xnor U434 (N_434,In_196,In_984);
nand U435 (N_435,In_758,In_126);
or U436 (N_436,In_460,In_393);
nand U437 (N_437,In_537,In_596);
nand U438 (N_438,In_404,In_714);
nor U439 (N_439,In_533,In_649);
or U440 (N_440,In_219,In_991);
or U441 (N_441,In_73,In_29);
nand U442 (N_442,In_722,In_501);
and U443 (N_443,In_50,In_236);
or U444 (N_444,In_401,In_74);
nor U445 (N_445,In_993,In_361);
nor U446 (N_446,In_721,In_230);
or U447 (N_447,In_381,In_710);
and U448 (N_448,In_100,In_990);
and U449 (N_449,In_434,In_131);
nand U450 (N_450,In_945,In_983);
or U451 (N_451,In_416,In_267);
or U452 (N_452,In_318,In_477);
and U453 (N_453,In_915,In_734);
and U454 (N_454,In_284,In_876);
xor U455 (N_455,In_709,In_375);
nor U456 (N_456,In_831,In_726);
and U457 (N_457,In_319,In_342);
nand U458 (N_458,In_148,In_970);
nand U459 (N_459,In_517,In_162);
and U460 (N_460,In_370,In_298);
nand U461 (N_461,In_911,In_564);
nor U462 (N_462,In_497,In_468);
nand U463 (N_463,In_207,In_41);
nand U464 (N_464,In_353,In_296);
and U465 (N_465,In_476,In_904);
or U466 (N_466,In_949,In_654);
and U467 (N_467,In_376,In_794);
or U468 (N_468,In_140,In_200);
nor U469 (N_469,In_673,In_55);
nor U470 (N_470,In_616,In_197);
or U471 (N_471,In_466,In_730);
or U472 (N_472,In_958,In_511);
and U473 (N_473,In_265,In_622);
nor U474 (N_474,In_31,In_67);
nand U475 (N_475,In_211,In_192);
and U476 (N_476,In_922,In_531);
nand U477 (N_477,In_386,In_127);
or U478 (N_478,In_373,In_887);
nand U479 (N_479,In_944,In_241);
nand U480 (N_480,In_828,In_618);
nand U481 (N_481,In_290,In_102);
xor U482 (N_482,In_176,In_565);
nand U483 (N_483,In_338,In_309);
or U484 (N_484,In_747,In_11);
nor U485 (N_485,In_413,In_630);
and U486 (N_486,In_96,In_246);
nand U487 (N_487,In_522,In_210);
nor U488 (N_488,In_959,In_566);
or U489 (N_489,In_896,In_395);
or U490 (N_490,In_520,In_587);
or U491 (N_491,In_283,In_770);
nand U492 (N_492,In_764,In_237);
and U493 (N_493,In_936,In_147);
nor U494 (N_494,In_391,In_535);
nor U495 (N_495,In_302,In_121);
or U496 (N_496,In_300,In_736);
or U497 (N_497,In_996,In_417);
xnor U498 (N_498,In_458,In_663);
and U499 (N_499,In_178,In_536);
nand U500 (N_500,N_493,N_110);
xnor U501 (N_501,N_166,N_448);
nand U502 (N_502,N_286,N_93);
or U503 (N_503,N_60,N_413);
and U504 (N_504,N_442,N_131);
or U505 (N_505,N_328,N_36);
nor U506 (N_506,N_171,N_485);
or U507 (N_507,N_28,N_265);
nor U508 (N_508,N_400,N_1);
or U509 (N_509,N_221,N_133);
nand U510 (N_510,N_406,N_169);
and U511 (N_511,N_360,N_106);
or U512 (N_512,N_25,N_48);
nor U513 (N_513,N_42,N_372);
and U514 (N_514,N_317,N_252);
nor U515 (N_515,N_52,N_426);
nor U516 (N_516,N_301,N_95);
and U517 (N_517,N_346,N_75);
nor U518 (N_518,N_136,N_473);
or U519 (N_519,N_441,N_460);
nor U520 (N_520,N_68,N_316);
or U521 (N_521,N_300,N_429);
nand U522 (N_522,N_283,N_471);
nand U523 (N_523,N_233,N_148);
nor U524 (N_524,N_210,N_90);
or U525 (N_525,N_211,N_386);
or U526 (N_526,N_38,N_65);
and U527 (N_527,N_497,N_320);
nand U528 (N_528,N_76,N_54);
nand U529 (N_529,N_405,N_327);
nor U530 (N_530,N_355,N_79);
nor U531 (N_531,N_50,N_127);
and U532 (N_532,N_86,N_198);
xnor U533 (N_533,N_183,N_103);
or U534 (N_534,N_91,N_230);
nor U535 (N_535,N_226,N_15);
and U536 (N_536,N_14,N_396);
nor U537 (N_537,N_255,N_475);
or U538 (N_538,N_321,N_308);
nor U539 (N_539,N_185,N_200);
nor U540 (N_540,N_254,N_378);
nor U541 (N_541,N_403,N_481);
or U542 (N_542,N_495,N_44);
xor U543 (N_543,N_145,N_137);
nand U544 (N_544,N_425,N_21);
or U545 (N_545,N_279,N_375);
nand U546 (N_546,N_268,N_351);
xor U547 (N_547,N_61,N_175);
or U548 (N_548,N_26,N_109);
nand U549 (N_549,N_488,N_203);
or U550 (N_550,N_8,N_276);
nand U551 (N_551,N_179,N_438);
nand U552 (N_552,N_0,N_58);
nand U553 (N_553,N_353,N_339);
or U554 (N_554,N_369,N_247);
and U555 (N_555,N_77,N_359);
or U556 (N_556,N_384,N_462);
and U557 (N_557,N_157,N_242);
and U558 (N_558,N_6,N_22);
or U559 (N_559,N_88,N_204);
nand U560 (N_560,N_260,N_105);
nand U561 (N_561,N_187,N_241);
nor U562 (N_562,N_326,N_464);
xnor U563 (N_563,N_463,N_323);
xnor U564 (N_564,N_153,N_285);
nand U565 (N_565,N_57,N_2);
nand U566 (N_566,N_487,N_7);
or U567 (N_567,N_251,N_370);
and U568 (N_568,N_262,N_480);
nand U569 (N_569,N_420,N_214);
or U570 (N_570,N_232,N_31);
nand U571 (N_571,N_150,N_12);
nor U572 (N_572,N_291,N_461);
nand U573 (N_573,N_223,N_212);
nand U574 (N_574,N_423,N_134);
nor U575 (N_575,N_97,N_410);
nand U576 (N_576,N_394,N_416);
nand U577 (N_577,N_310,N_253);
nor U578 (N_578,N_250,N_45);
or U579 (N_579,N_334,N_120);
and U580 (N_580,N_4,N_20);
nor U581 (N_581,N_284,N_78);
nor U582 (N_582,N_368,N_296);
and U583 (N_583,N_486,N_427);
xor U584 (N_584,N_82,N_468);
nand U585 (N_585,N_193,N_382);
nor U586 (N_586,N_318,N_305);
or U587 (N_587,N_62,N_356);
nor U588 (N_588,N_287,N_195);
nor U589 (N_589,N_391,N_408);
nor U590 (N_590,N_274,N_99);
nand U591 (N_591,N_39,N_281);
nor U592 (N_592,N_104,N_272);
or U593 (N_593,N_118,N_451);
or U594 (N_594,N_174,N_436);
and U595 (N_595,N_432,N_398);
nand U596 (N_596,N_474,N_182);
and U597 (N_597,N_155,N_213);
or U598 (N_598,N_392,N_123);
or U599 (N_599,N_139,N_458);
nand U600 (N_600,N_362,N_361);
and U601 (N_601,N_496,N_498);
nand U602 (N_602,N_83,N_409);
nand U603 (N_603,N_350,N_302);
nand U604 (N_604,N_132,N_490);
or U605 (N_605,N_470,N_388);
and U606 (N_606,N_494,N_47);
xnor U607 (N_607,N_231,N_112);
nor U608 (N_608,N_377,N_341);
xnor U609 (N_609,N_261,N_266);
and U610 (N_610,N_271,N_435);
nor U611 (N_611,N_417,N_189);
nand U612 (N_612,N_440,N_428);
nand U613 (N_613,N_437,N_84);
or U614 (N_614,N_69,N_217);
nand U615 (N_615,N_479,N_239);
or U616 (N_616,N_349,N_202);
nand U617 (N_617,N_224,N_176);
or U618 (N_618,N_344,N_383);
nor U619 (N_619,N_122,N_72);
or U620 (N_620,N_35,N_264);
or U621 (N_621,N_414,N_331);
or U622 (N_622,N_121,N_173);
and U623 (N_623,N_13,N_24);
nor U624 (N_624,N_222,N_484);
nor U625 (N_625,N_191,N_46);
nor U626 (N_626,N_395,N_228);
nand U627 (N_627,N_135,N_333);
and U628 (N_628,N_366,N_269);
and U629 (N_629,N_162,N_55);
or U630 (N_630,N_172,N_444);
nor U631 (N_631,N_161,N_259);
xnor U632 (N_632,N_111,N_290);
nand U633 (N_633,N_483,N_219);
xor U634 (N_634,N_186,N_263);
nor U635 (N_635,N_130,N_141);
nor U636 (N_636,N_335,N_100);
and U637 (N_637,N_245,N_70);
nand U638 (N_638,N_126,N_304);
nand U639 (N_639,N_455,N_297);
and U640 (N_640,N_390,N_397);
xnor U641 (N_641,N_348,N_142);
and U642 (N_642,N_312,N_41);
xor U643 (N_643,N_220,N_146);
nand U644 (N_644,N_453,N_342);
and U645 (N_645,N_154,N_240);
nor U646 (N_646,N_190,N_404);
and U647 (N_647,N_332,N_168);
nor U648 (N_648,N_450,N_11);
or U649 (N_649,N_337,N_147);
xor U650 (N_650,N_180,N_401);
nand U651 (N_651,N_129,N_439);
or U652 (N_652,N_199,N_299);
or U653 (N_653,N_376,N_81);
or U654 (N_654,N_143,N_116);
nor U655 (N_655,N_466,N_352);
and U656 (N_656,N_215,N_277);
nand U657 (N_657,N_295,N_354);
nor U658 (N_658,N_107,N_364);
nand U659 (N_659,N_373,N_30);
or U660 (N_660,N_492,N_419);
and U661 (N_661,N_119,N_443);
nor U662 (N_662,N_125,N_282);
nor U663 (N_663,N_138,N_298);
xnor U664 (N_664,N_381,N_114);
nor U665 (N_665,N_365,N_445);
or U666 (N_666,N_10,N_206);
or U667 (N_667,N_152,N_23);
nor U668 (N_668,N_74,N_34);
and U669 (N_669,N_9,N_209);
or U670 (N_670,N_482,N_258);
and U671 (N_671,N_37,N_67);
and U672 (N_672,N_201,N_307);
or U673 (N_673,N_216,N_73);
xor U674 (N_674,N_345,N_280);
nor U675 (N_675,N_17,N_66);
and U676 (N_676,N_367,N_399);
xor U677 (N_677,N_159,N_273);
nor U678 (N_678,N_32,N_165);
nor U679 (N_679,N_256,N_207);
and U680 (N_680,N_319,N_446);
xnor U681 (N_681,N_467,N_140);
nand U682 (N_682,N_192,N_177);
and U683 (N_683,N_108,N_156);
or U684 (N_684,N_340,N_387);
nand U685 (N_685,N_489,N_336);
and U686 (N_686,N_433,N_246);
nor U687 (N_687,N_53,N_87);
nand U688 (N_688,N_56,N_347);
nor U689 (N_689,N_469,N_456);
xor U690 (N_690,N_343,N_160);
nand U691 (N_691,N_96,N_306);
xor U692 (N_692,N_208,N_178);
and U693 (N_693,N_324,N_236);
and U694 (N_694,N_314,N_64);
or U695 (N_695,N_267,N_477);
nand U696 (N_696,N_115,N_371);
or U697 (N_697,N_167,N_457);
or U698 (N_698,N_275,N_430);
xnor U699 (N_699,N_311,N_447);
and U700 (N_700,N_412,N_329);
nand U701 (N_701,N_94,N_421);
and U702 (N_702,N_170,N_205);
nand U703 (N_703,N_51,N_393);
xor U704 (N_704,N_144,N_128);
nand U705 (N_705,N_196,N_227);
nor U706 (N_706,N_124,N_248);
nand U707 (N_707,N_49,N_472);
nand U708 (N_708,N_293,N_101);
and U709 (N_709,N_424,N_292);
or U710 (N_710,N_163,N_243);
nor U711 (N_711,N_235,N_452);
or U712 (N_712,N_3,N_402);
nor U713 (N_713,N_43,N_257);
nor U714 (N_714,N_465,N_71);
or U715 (N_715,N_313,N_309);
xnor U716 (N_716,N_113,N_27);
nand U717 (N_717,N_63,N_92);
nand U718 (N_718,N_181,N_237);
and U719 (N_719,N_449,N_270);
or U720 (N_720,N_415,N_434);
nor U721 (N_721,N_151,N_379);
nor U722 (N_722,N_229,N_19);
xnor U723 (N_723,N_98,N_459);
or U724 (N_724,N_5,N_374);
nor U725 (N_725,N_225,N_330);
xor U726 (N_726,N_40,N_218);
nand U727 (N_727,N_238,N_476);
nand U728 (N_728,N_158,N_249);
nor U729 (N_729,N_244,N_149);
or U730 (N_730,N_325,N_278);
and U731 (N_731,N_407,N_363);
nand U732 (N_732,N_303,N_288);
and U733 (N_733,N_380,N_322);
or U734 (N_734,N_358,N_389);
and U735 (N_735,N_18,N_422);
nor U736 (N_736,N_188,N_499);
nor U737 (N_737,N_315,N_85);
and U738 (N_738,N_184,N_418);
xnor U739 (N_739,N_194,N_16);
or U740 (N_740,N_385,N_89);
and U741 (N_741,N_357,N_491);
nand U742 (N_742,N_234,N_117);
or U743 (N_743,N_478,N_431);
nor U744 (N_744,N_454,N_411);
nand U745 (N_745,N_29,N_338);
nand U746 (N_746,N_294,N_80);
or U747 (N_747,N_33,N_164);
nor U748 (N_748,N_289,N_102);
or U749 (N_749,N_59,N_197);
nand U750 (N_750,N_408,N_33);
xor U751 (N_751,N_150,N_391);
and U752 (N_752,N_392,N_224);
nor U753 (N_753,N_271,N_48);
and U754 (N_754,N_301,N_440);
nor U755 (N_755,N_467,N_300);
nand U756 (N_756,N_366,N_157);
and U757 (N_757,N_347,N_82);
nor U758 (N_758,N_195,N_126);
and U759 (N_759,N_214,N_136);
nor U760 (N_760,N_402,N_217);
and U761 (N_761,N_242,N_307);
xor U762 (N_762,N_231,N_105);
nor U763 (N_763,N_373,N_108);
nand U764 (N_764,N_61,N_67);
nand U765 (N_765,N_399,N_156);
or U766 (N_766,N_295,N_483);
and U767 (N_767,N_415,N_325);
or U768 (N_768,N_373,N_185);
nor U769 (N_769,N_66,N_198);
nor U770 (N_770,N_452,N_445);
and U771 (N_771,N_100,N_278);
and U772 (N_772,N_183,N_123);
xor U773 (N_773,N_5,N_204);
nand U774 (N_774,N_50,N_158);
nor U775 (N_775,N_47,N_428);
nor U776 (N_776,N_249,N_122);
or U777 (N_777,N_270,N_198);
nand U778 (N_778,N_291,N_426);
xor U779 (N_779,N_403,N_383);
and U780 (N_780,N_489,N_313);
nand U781 (N_781,N_464,N_404);
nor U782 (N_782,N_25,N_279);
nand U783 (N_783,N_386,N_420);
or U784 (N_784,N_43,N_211);
nand U785 (N_785,N_80,N_421);
nor U786 (N_786,N_54,N_439);
and U787 (N_787,N_458,N_110);
nor U788 (N_788,N_430,N_494);
and U789 (N_789,N_220,N_304);
nand U790 (N_790,N_353,N_300);
nor U791 (N_791,N_211,N_27);
nor U792 (N_792,N_302,N_430);
nor U793 (N_793,N_488,N_379);
xor U794 (N_794,N_287,N_350);
nor U795 (N_795,N_161,N_169);
and U796 (N_796,N_13,N_408);
or U797 (N_797,N_268,N_408);
nand U798 (N_798,N_362,N_249);
and U799 (N_799,N_159,N_374);
nor U800 (N_800,N_3,N_229);
or U801 (N_801,N_122,N_44);
nand U802 (N_802,N_481,N_320);
nor U803 (N_803,N_190,N_158);
nor U804 (N_804,N_453,N_364);
or U805 (N_805,N_211,N_13);
nand U806 (N_806,N_230,N_297);
nor U807 (N_807,N_78,N_354);
nand U808 (N_808,N_487,N_339);
and U809 (N_809,N_54,N_120);
xor U810 (N_810,N_459,N_238);
and U811 (N_811,N_246,N_144);
and U812 (N_812,N_12,N_389);
or U813 (N_813,N_341,N_1);
nand U814 (N_814,N_417,N_331);
or U815 (N_815,N_173,N_48);
or U816 (N_816,N_65,N_429);
nand U817 (N_817,N_280,N_305);
nand U818 (N_818,N_0,N_226);
or U819 (N_819,N_273,N_45);
and U820 (N_820,N_452,N_213);
xnor U821 (N_821,N_258,N_350);
nand U822 (N_822,N_118,N_162);
nor U823 (N_823,N_290,N_115);
or U824 (N_824,N_274,N_74);
and U825 (N_825,N_403,N_264);
or U826 (N_826,N_13,N_200);
and U827 (N_827,N_293,N_177);
and U828 (N_828,N_290,N_82);
or U829 (N_829,N_218,N_168);
xor U830 (N_830,N_387,N_326);
and U831 (N_831,N_91,N_316);
xor U832 (N_832,N_465,N_182);
or U833 (N_833,N_44,N_270);
or U834 (N_834,N_458,N_331);
and U835 (N_835,N_33,N_332);
nor U836 (N_836,N_337,N_421);
nand U837 (N_837,N_351,N_77);
and U838 (N_838,N_389,N_208);
or U839 (N_839,N_341,N_69);
or U840 (N_840,N_378,N_69);
nor U841 (N_841,N_363,N_419);
nand U842 (N_842,N_87,N_151);
xor U843 (N_843,N_25,N_28);
and U844 (N_844,N_283,N_160);
or U845 (N_845,N_361,N_444);
and U846 (N_846,N_144,N_268);
nand U847 (N_847,N_423,N_259);
nand U848 (N_848,N_12,N_44);
or U849 (N_849,N_96,N_2);
and U850 (N_850,N_256,N_295);
nor U851 (N_851,N_377,N_58);
nor U852 (N_852,N_66,N_60);
and U853 (N_853,N_161,N_404);
or U854 (N_854,N_238,N_295);
or U855 (N_855,N_429,N_74);
xor U856 (N_856,N_276,N_236);
or U857 (N_857,N_434,N_253);
and U858 (N_858,N_143,N_145);
and U859 (N_859,N_109,N_276);
nand U860 (N_860,N_355,N_83);
and U861 (N_861,N_233,N_394);
or U862 (N_862,N_309,N_101);
and U863 (N_863,N_39,N_59);
nor U864 (N_864,N_138,N_432);
and U865 (N_865,N_207,N_171);
xnor U866 (N_866,N_399,N_441);
or U867 (N_867,N_430,N_412);
or U868 (N_868,N_217,N_290);
and U869 (N_869,N_379,N_17);
and U870 (N_870,N_118,N_415);
or U871 (N_871,N_334,N_48);
xnor U872 (N_872,N_91,N_268);
and U873 (N_873,N_439,N_452);
and U874 (N_874,N_206,N_360);
nor U875 (N_875,N_363,N_357);
nor U876 (N_876,N_247,N_39);
or U877 (N_877,N_27,N_21);
nor U878 (N_878,N_399,N_255);
nand U879 (N_879,N_82,N_495);
nand U880 (N_880,N_209,N_282);
nor U881 (N_881,N_28,N_168);
nand U882 (N_882,N_236,N_30);
and U883 (N_883,N_57,N_281);
nor U884 (N_884,N_449,N_257);
nor U885 (N_885,N_174,N_370);
or U886 (N_886,N_25,N_439);
and U887 (N_887,N_328,N_218);
nand U888 (N_888,N_489,N_206);
nor U889 (N_889,N_174,N_385);
and U890 (N_890,N_276,N_358);
or U891 (N_891,N_191,N_318);
nor U892 (N_892,N_376,N_262);
nor U893 (N_893,N_244,N_96);
nor U894 (N_894,N_408,N_76);
nand U895 (N_895,N_96,N_171);
nor U896 (N_896,N_346,N_408);
nor U897 (N_897,N_247,N_183);
xor U898 (N_898,N_411,N_247);
nand U899 (N_899,N_494,N_141);
or U900 (N_900,N_470,N_453);
nor U901 (N_901,N_241,N_352);
xnor U902 (N_902,N_68,N_347);
and U903 (N_903,N_65,N_26);
nand U904 (N_904,N_173,N_6);
nand U905 (N_905,N_105,N_45);
or U906 (N_906,N_134,N_102);
and U907 (N_907,N_130,N_159);
and U908 (N_908,N_262,N_406);
and U909 (N_909,N_461,N_330);
xnor U910 (N_910,N_37,N_287);
or U911 (N_911,N_300,N_394);
nor U912 (N_912,N_234,N_226);
and U913 (N_913,N_190,N_11);
nor U914 (N_914,N_42,N_313);
nand U915 (N_915,N_290,N_221);
nor U916 (N_916,N_443,N_422);
and U917 (N_917,N_383,N_12);
or U918 (N_918,N_360,N_8);
xor U919 (N_919,N_75,N_87);
and U920 (N_920,N_353,N_157);
and U921 (N_921,N_304,N_150);
nand U922 (N_922,N_121,N_311);
nand U923 (N_923,N_9,N_203);
nor U924 (N_924,N_427,N_455);
or U925 (N_925,N_209,N_140);
and U926 (N_926,N_96,N_282);
and U927 (N_927,N_130,N_51);
nor U928 (N_928,N_176,N_183);
or U929 (N_929,N_496,N_5);
nor U930 (N_930,N_297,N_351);
or U931 (N_931,N_465,N_48);
xnor U932 (N_932,N_411,N_319);
nor U933 (N_933,N_101,N_474);
or U934 (N_934,N_246,N_37);
nor U935 (N_935,N_137,N_367);
and U936 (N_936,N_421,N_333);
or U937 (N_937,N_238,N_87);
nand U938 (N_938,N_147,N_41);
xor U939 (N_939,N_253,N_307);
xor U940 (N_940,N_319,N_167);
nor U941 (N_941,N_188,N_31);
or U942 (N_942,N_351,N_197);
nor U943 (N_943,N_340,N_214);
xnor U944 (N_944,N_358,N_386);
nor U945 (N_945,N_375,N_288);
and U946 (N_946,N_355,N_117);
xor U947 (N_947,N_394,N_492);
nor U948 (N_948,N_139,N_331);
or U949 (N_949,N_399,N_467);
xor U950 (N_950,N_63,N_97);
xor U951 (N_951,N_346,N_51);
or U952 (N_952,N_53,N_461);
nand U953 (N_953,N_374,N_40);
nor U954 (N_954,N_236,N_306);
nand U955 (N_955,N_352,N_469);
nand U956 (N_956,N_144,N_245);
and U957 (N_957,N_269,N_125);
nand U958 (N_958,N_463,N_453);
nand U959 (N_959,N_94,N_349);
or U960 (N_960,N_229,N_74);
xor U961 (N_961,N_324,N_125);
or U962 (N_962,N_215,N_278);
nor U963 (N_963,N_28,N_151);
or U964 (N_964,N_26,N_449);
nor U965 (N_965,N_130,N_264);
and U966 (N_966,N_419,N_83);
nor U967 (N_967,N_322,N_111);
nand U968 (N_968,N_364,N_376);
nor U969 (N_969,N_123,N_339);
or U970 (N_970,N_15,N_254);
nor U971 (N_971,N_253,N_69);
nand U972 (N_972,N_87,N_107);
or U973 (N_973,N_303,N_405);
nand U974 (N_974,N_134,N_482);
and U975 (N_975,N_339,N_78);
nor U976 (N_976,N_344,N_453);
or U977 (N_977,N_306,N_149);
and U978 (N_978,N_142,N_20);
nand U979 (N_979,N_10,N_24);
nor U980 (N_980,N_221,N_391);
and U981 (N_981,N_8,N_66);
or U982 (N_982,N_430,N_393);
nor U983 (N_983,N_267,N_193);
and U984 (N_984,N_322,N_210);
nand U985 (N_985,N_19,N_231);
nand U986 (N_986,N_91,N_59);
or U987 (N_987,N_358,N_273);
or U988 (N_988,N_496,N_161);
or U989 (N_989,N_131,N_470);
xnor U990 (N_990,N_395,N_488);
or U991 (N_991,N_255,N_458);
nor U992 (N_992,N_460,N_53);
nor U993 (N_993,N_241,N_266);
or U994 (N_994,N_76,N_149);
xor U995 (N_995,N_376,N_218);
nor U996 (N_996,N_417,N_487);
nand U997 (N_997,N_114,N_29);
or U998 (N_998,N_185,N_23);
nor U999 (N_999,N_396,N_207);
and U1000 (N_1000,N_612,N_954);
and U1001 (N_1001,N_682,N_753);
nor U1002 (N_1002,N_801,N_807);
xor U1003 (N_1003,N_935,N_722);
or U1004 (N_1004,N_571,N_538);
nand U1005 (N_1005,N_604,N_570);
nand U1006 (N_1006,N_528,N_669);
and U1007 (N_1007,N_728,N_852);
and U1008 (N_1008,N_664,N_884);
and U1009 (N_1009,N_972,N_760);
or U1010 (N_1010,N_556,N_514);
or U1011 (N_1011,N_955,N_877);
xnor U1012 (N_1012,N_867,N_687);
and U1013 (N_1013,N_762,N_983);
nand U1014 (N_1014,N_993,N_778);
or U1015 (N_1015,N_500,N_841);
or U1016 (N_1016,N_531,N_900);
or U1017 (N_1017,N_584,N_675);
nor U1018 (N_1018,N_859,N_748);
and U1019 (N_1019,N_743,N_880);
and U1020 (N_1020,N_836,N_525);
and U1021 (N_1021,N_513,N_712);
and U1022 (N_1022,N_716,N_700);
xor U1023 (N_1023,N_517,N_910);
and U1024 (N_1024,N_978,N_749);
and U1025 (N_1025,N_765,N_860);
nand U1026 (N_1026,N_816,N_620);
nor U1027 (N_1027,N_793,N_740);
or U1028 (N_1028,N_624,N_789);
nand U1029 (N_1029,N_565,N_835);
or U1030 (N_1030,N_638,N_804);
or U1031 (N_1031,N_694,N_651);
nand U1032 (N_1032,N_674,N_924);
nor U1033 (N_1033,N_999,N_876);
and U1034 (N_1034,N_666,N_803);
nand U1035 (N_1035,N_794,N_779);
nand U1036 (N_1036,N_643,N_961);
and U1037 (N_1037,N_908,N_710);
and U1038 (N_1038,N_781,N_815);
nand U1039 (N_1039,N_695,N_953);
or U1040 (N_1040,N_809,N_882);
nor U1041 (N_1041,N_990,N_599);
nand U1042 (N_1042,N_614,N_906);
or U1043 (N_1043,N_977,N_527);
nand U1044 (N_1044,N_826,N_667);
nand U1045 (N_1045,N_504,N_865);
nand U1046 (N_1046,N_697,N_621);
nor U1047 (N_1047,N_799,N_692);
and U1048 (N_1048,N_555,N_560);
and U1049 (N_1049,N_640,N_970);
nand U1050 (N_1050,N_656,N_505);
or U1051 (N_1051,N_639,N_855);
and U1052 (N_1052,N_548,N_995);
and U1053 (N_1053,N_521,N_573);
nor U1054 (N_1054,N_768,N_685);
nand U1055 (N_1055,N_863,N_683);
nand U1056 (N_1056,N_788,N_557);
or U1057 (N_1057,N_524,N_979);
nand U1058 (N_1058,N_702,N_535);
nor U1059 (N_1059,N_838,N_719);
nand U1060 (N_1060,N_818,N_647);
nor U1061 (N_1061,N_546,N_750);
nor U1062 (N_1062,N_948,N_917);
nor U1063 (N_1063,N_795,N_580);
or U1064 (N_1064,N_627,N_926);
and U1065 (N_1065,N_597,N_886);
nor U1066 (N_1066,N_777,N_958);
or U1067 (N_1067,N_976,N_537);
nor U1068 (N_1068,N_622,N_704);
nand U1069 (N_1069,N_520,N_610);
nor U1070 (N_1070,N_997,N_629);
nor U1071 (N_1071,N_774,N_840);
nor U1072 (N_1072,N_893,N_844);
nor U1073 (N_1073,N_864,N_897);
nand U1074 (N_1074,N_982,N_888);
and U1075 (N_1075,N_681,N_628);
or U1076 (N_1076,N_644,N_892);
or U1077 (N_1077,N_652,N_601);
and U1078 (N_1078,N_988,N_737);
nor U1079 (N_1079,N_655,N_654);
nand U1080 (N_1080,N_941,N_733);
xnor U1081 (N_1081,N_657,N_909);
or U1082 (N_1082,N_649,N_585);
or U1083 (N_1083,N_755,N_945);
nor U1084 (N_1084,N_709,N_767);
or U1085 (N_1085,N_751,N_928);
nand U1086 (N_1086,N_678,N_530);
nor U1087 (N_1087,N_872,N_870);
nand U1088 (N_1088,N_746,N_745);
and U1089 (N_1089,N_756,N_559);
nand U1090 (N_1090,N_632,N_889);
nor U1091 (N_1091,N_819,N_980);
nand U1092 (N_1092,N_831,N_786);
and U1093 (N_1093,N_849,N_853);
or U1094 (N_1094,N_944,N_741);
nor U1095 (N_1095,N_551,N_890);
nand U1096 (N_1096,N_938,N_785);
and U1097 (N_1097,N_994,N_532);
or U1098 (N_1098,N_858,N_856);
nand U1099 (N_1099,N_752,N_519);
nand U1100 (N_1100,N_846,N_761);
xor U1101 (N_1101,N_706,N_964);
xor U1102 (N_1102,N_773,N_792);
xor U1103 (N_1103,N_518,N_625);
or U1104 (N_1104,N_626,N_763);
nand U1105 (N_1105,N_642,N_526);
or U1106 (N_1106,N_608,N_996);
nor U1107 (N_1107,N_800,N_633);
and U1108 (N_1108,N_775,N_830);
nand U1109 (N_1109,N_617,N_729);
and U1110 (N_1110,N_688,N_973);
or U1111 (N_1111,N_757,N_873);
nor U1112 (N_1112,N_934,N_673);
nand U1113 (N_1113,N_501,N_575);
xor U1114 (N_1114,N_658,N_850);
or U1115 (N_1115,N_588,N_966);
and U1116 (N_1116,N_554,N_820);
and U1117 (N_1117,N_933,N_582);
and U1118 (N_1118,N_506,N_904);
or U1119 (N_1119,N_663,N_529);
and U1120 (N_1120,N_827,N_959);
nand U1121 (N_1121,N_613,N_914);
and U1122 (N_1122,N_566,N_572);
and U1123 (N_1123,N_833,N_805);
nand U1124 (N_1124,N_808,N_583);
xor U1125 (N_1125,N_713,N_828);
nor U1126 (N_1126,N_915,N_821);
nor U1127 (N_1127,N_851,N_593);
and U1128 (N_1128,N_829,N_698);
nand U1129 (N_1129,N_711,N_534);
or U1130 (N_1130,N_616,N_545);
nand U1131 (N_1131,N_871,N_736);
or U1132 (N_1132,N_881,N_854);
or U1133 (N_1133,N_516,N_609);
xnor U1134 (N_1134,N_540,N_986);
or U1135 (N_1135,N_596,N_603);
nor U1136 (N_1136,N_802,N_747);
or U1137 (N_1137,N_732,N_600);
or U1138 (N_1138,N_734,N_962);
xnor U1139 (N_1139,N_590,N_998);
xnor U1140 (N_1140,N_512,N_949);
nand U1141 (N_1141,N_776,N_672);
and U1142 (N_1142,N_842,N_707);
xnor U1143 (N_1143,N_739,N_845);
nand U1144 (N_1144,N_696,N_641);
or U1145 (N_1145,N_984,N_561);
or U1146 (N_1146,N_951,N_940);
xor U1147 (N_1147,N_701,N_987);
nor U1148 (N_1148,N_703,N_857);
or U1149 (N_1149,N_536,N_634);
or U1150 (N_1150,N_916,N_677);
and U1151 (N_1151,N_731,N_907);
nor U1152 (N_1152,N_630,N_797);
nand U1153 (N_1153,N_509,N_637);
or U1154 (N_1154,N_541,N_960);
xnor U1155 (N_1155,N_563,N_885);
nand U1156 (N_1156,N_587,N_725);
nand U1157 (N_1157,N_783,N_971);
or U1158 (N_1158,N_502,N_868);
xor U1159 (N_1159,N_550,N_942);
or U1160 (N_1160,N_533,N_861);
nor U1161 (N_1161,N_898,N_635);
xor U1162 (N_1162,N_595,N_772);
or U1163 (N_1163,N_931,N_661);
or U1164 (N_1164,N_592,N_539);
and U1165 (N_1165,N_887,N_963);
nand U1166 (N_1166,N_899,N_562);
nor U1167 (N_1167,N_759,N_847);
or U1168 (N_1168,N_992,N_659);
and U1169 (N_1169,N_932,N_866);
and U1170 (N_1170,N_782,N_766);
nand U1171 (N_1171,N_567,N_883);
nor U1172 (N_1172,N_686,N_758);
or U1173 (N_1173,N_579,N_730);
or U1174 (N_1174,N_586,N_947);
nand U1175 (N_1175,N_848,N_552);
nor U1176 (N_1176,N_645,N_558);
or U1177 (N_1177,N_939,N_665);
xnor U1178 (N_1178,N_771,N_875);
and U1179 (N_1179,N_508,N_679);
nand U1180 (N_1180,N_879,N_822);
xor U1181 (N_1181,N_929,N_581);
nor U1182 (N_1182,N_544,N_901);
nor U1183 (N_1183,N_589,N_985);
or U1184 (N_1184,N_738,N_650);
nand U1185 (N_1185,N_812,N_720);
or U1186 (N_1186,N_598,N_619);
nor U1187 (N_1187,N_576,N_891);
and U1188 (N_1188,N_918,N_974);
and U1189 (N_1189,N_930,N_648);
or U1190 (N_1190,N_925,N_811);
or U1191 (N_1191,N_618,N_832);
or U1192 (N_1192,N_594,N_549);
or U1193 (N_1193,N_726,N_507);
or U1194 (N_1194,N_723,N_834);
and U1195 (N_1195,N_814,N_724);
or U1196 (N_1196,N_912,N_668);
nor U1197 (N_1197,N_965,N_670);
or U1198 (N_1198,N_913,N_956);
nand U1199 (N_1199,N_744,N_991);
nor U1200 (N_1200,N_862,N_511);
and U1201 (N_1201,N_605,N_896);
nand U1202 (N_1202,N_680,N_510);
nor U1203 (N_1203,N_611,N_981);
nor U1204 (N_1204,N_869,N_791);
or U1205 (N_1205,N_523,N_784);
nor U1206 (N_1206,N_577,N_717);
and U1207 (N_1207,N_905,N_967);
and U1208 (N_1208,N_787,N_894);
nand U1209 (N_1209,N_754,N_542);
nor U1210 (N_1210,N_553,N_543);
or U1211 (N_1211,N_950,N_568);
nand U1212 (N_1212,N_503,N_969);
nor U1213 (N_1213,N_769,N_721);
nor U1214 (N_1214,N_689,N_602);
nor U1215 (N_1215,N_684,N_813);
or U1216 (N_1216,N_957,N_823);
nor U1217 (N_1217,N_690,N_569);
or U1218 (N_1218,N_607,N_646);
nor U1219 (N_1219,N_718,N_825);
or U1220 (N_1220,N_631,N_671);
or U1221 (N_1221,N_839,N_764);
xnor U1222 (N_1222,N_919,N_727);
or U1223 (N_1223,N_923,N_662);
or U1224 (N_1224,N_975,N_615);
nand U1225 (N_1225,N_927,N_699);
nor U1226 (N_1226,N_946,N_903);
xor U1227 (N_1227,N_660,N_653);
nand U1228 (N_1228,N_522,N_606);
and U1229 (N_1229,N_564,N_943);
and U1230 (N_1230,N_798,N_591);
and U1231 (N_1231,N_810,N_806);
nor U1232 (N_1232,N_817,N_952);
nor U1233 (N_1233,N_902,N_936);
xnor U1234 (N_1234,N_878,N_989);
nand U1235 (N_1235,N_796,N_636);
nor U1236 (N_1236,N_735,N_742);
or U1237 (N_1237,N_715,N_547);
and U1238 (N_1238,N_824,N_895);
or U1239 (N_1239,N_911,N_920);
nor U1240 (N_1240,N_837,N_623);
nand U1241 (N_1241,N_968,N_578);
or U1242 (N_1242,N_770,N_708);
xnor U1243 (N_1243,N_921,N_676);
nand U1244 (N_1244,N_780,N_790);
and U1245 (N_1245,N_705,N_874);
and U1246 (N_1246,N_515,N_691);
nor U1247 (N_1247,N_937,N_574);
nor U1248 (N_1248,N_714,N_693);
nor U1249 (N_1249,N_922,N_843);
or U1250 (N_1250,N_602,N_984);
and U1251 (N_1251,N_741,N_896);
and U1252 (N_1252,N_796,N_704);
nand U1253 (N_1253,N_757,N_912);
nor U1254 (N_1254,N_882,N_682);
nand U1255 (N_1255,N_943,N_707);
nor U1256 (N_1256,N_542,N_606);
nand U1257 (N_1257,N_831,N_626);
xnor U1258 (N_1258,N_598,N_786);
and U1259 (N_1259,N_958,N_837);
nor U1260 (N_1260,N_863,N_617);
nand U1261 (N_1261,N_676,N_527);
or U1262 (N_1262,N_599,N_950);
or U1263 (N_1263,N_793,N_831);
or U1264 (N_1264,N_856,N_754);
and U1265 (N_1265,N_596,N_812);
and U1266 (N_1266,N_791,N_862);
or U1267 (N_1267,N_523,N_862);
and U1268 (N_1268,N_845,N_575);
and U1269 (N_1269,N_695,N_757);
xnor U1270 (N_1270,N_899,N_705);
or U1271 (N_1271,N_897,N_965);
nand U1272 (N_1272,N_850,N_665);
or U1273 (N_1273,N_697,N_699);
and U1274 (N_1274,N_516,N_669);
xnor U1275 (N_1275,N_969,N_629);
nor U1276 (N_1276,N_719,N_670);
or U1277 (N_1277,N_509,N_918);
and U1278 (N_1278,N_793,N_561);
nand U1279 (N_1279,N_761,N_688);
or U1280 (N_1280,N_634,N_985);
or U1281 (N_1281,N_805,N_664);
xor U1282 (N_1282,N_672,N_798);
nand U1283 (N_1283,N_706,N_612);
nor U1284 (N_1284,N_820,N_599);
xor U1285 (N_1285,N_558,N_965);
and U1286 (N_1286,N_992,N_804);
nand U1287 (N_1287,N_803,N_948);
nand U1288 (N_1288,N_550,N_526);
or U1289 (N_1289,N_609,N_591);
nand U1290 (N_1290,N_571,N_629);
nand U1291 (N_1291,N_646,N_715);
nand U1292 (N_1292,N_577,N_684);
nand U1293 (N_1293,N_898,N_568);
or U1294 (N_1294,N_567,N_972);
nand U1295 (N_1295,N_585,N_627);
nand U1296 (N_1296,N_685,N_993);
and U1297 (N_1297,N_778,N_675);
and U1298 (N_1298,N_751,N_873);
and U1299 (N_1299,N_756,N_881);
nor U1300 (N_1300,N_971,N_953);
nor U1301 (N_1301,N_705,N_853);
nor U1302 (N_1302,N_680,N_686);
nand U1303 (N_1303,N_546,N_986);
nor U1304 (N_1304,N_832,N_681);
nand U1305 (N_1305,N_522,N_843);
nand U1306 (N_1306,N_550,N_935);
or U1307 (N_1307,N_614,N_806);
nor U1308 (N_1308,N_801,N_924);
or U1309 (N_1309,N_695,N_927);
or U1310 (N_1310,N_688,N_694);
and U1311 (N_1311,N_530,N_639);
nor U1312 (N_1312,N_608,N_880);
and U1313 (N_1313,N_731,N_871);
xnor U1314 (N_1314,N_865,N_749);
xor U1315 (N_1315,N_515,N_598);
and U1316 (N_1316,N_713,N_575);
and U1317 (N_1317,N_974,N_926);
or U1318 (N_1318,N_737,N_613);
and U1319 (N_1319,N_534,N_563);
and U1320 (N_1320,N_647,N_600);
nor U1321 (N_1321,N_587,N_942);
nor U1322 (N_1322,N_710,N_954);
nor U1323 (N_1323,N_843,N_641);
nor U1324 (N_1324,N_697,N_591);
nor U1325 (N_1325,N_566,N_567);
nor U1326 (N_1326,N_618,N_547);
or U1327 (N_1327,N_670,N_638);
and U1328 (N_1328,N_567,N_672);
nor U1329 (N_1329,N_615,N_681);
xor U1330 (N_1330,N_921,N_810);
nand U1331 (N_1331,N_505,N_696);
or U1332 (N_1332,N_673,N_721);
and U1333 (N_1333,N_701,N_920);
nor U1334 (N_1334,N_527,N_819);
and U1335 (N_1335,N_729,N_543);
nand U1336 (N_1336,N_762,N_654);
nor U1337 (N_1337,N_684,N_788);
and U1338 (N_1338,N_519,N_745);
nor U1339 (N_1339,N_932,N_916);
nor U1340 (N_1340,N_971,N_912);
and U1341 (N_1341,N_676,N_829);
nand U1342 (N_1342,N_635,N_685);
or U1343 (N_1343,N_976,N_525);
and U1344 (N_1344,N_557,N_927);
nor U1345 (N_1345,N_709,N_877);
nor U1346 (N_1346,N_867,N_905);
nor U1347 (N_1347,N_715,N_929);
nor U1348 (N_1348,N_569,N_870);
xnor U1349 (N_1349,N_784,N_754);
nor U1350 (N_1350,N_989,N_705);
nand U1351 (N_1351,N_980,N_744);
and U1352 (N_1352,N_517,N_737);
or U1353 (N_1353,N_925,N_552);
and U1354 (N_1354,N_914,N_569);
and U1355 (N_1355,N_786,N_617);
nand U1356 (N_1356,N_953,N_877);
and U1357 (N_1357,N_747,N_657);
or U1358 (N_1358,N_521,N_871);
xor U1359 (N_1359,N_501,N_519);
or U1360 (N_1360,N_551,N_883);
nand U1361 (N_1361,N_842,N_612);
nor U1362 (N_1362,N_702,N_622);
nand U1363 (N_1363,N_993,N_553);
xnor U1364 (N_1364,N_808,N_753);
and U1365 (N_1365,N_930,N_816);
or U1366 (N_1366,N_807,N_632);
nand U1367 (N_1367,N_639,N_563);
nand U1368 (N_1368,N_933,N_814);
or U1369 (N_1369,N_966,N_803);
or U1370 (N_1370,N_671,N_836);
nor U1371 (N_1371,N_936,N_801);
nor U1372 (N_1372,N_657,N_939);
nand U1373 (N_1373,N_760,N_743);
and U1374 (N_1374,N_513,N_950);
nor U1375 (N_1375,N_831,N_658);
xor U1376 (N_1376,N_960,N_556);
nor U1377 (N_1377,N_672,N_565);
and U1378 (N_1378,N_994,N_550);
nor U1379 (N_1379,N_635,N_615);
or U1380 (N_1380,N_862,N_858);
nand U1381 (N_1381,N_581,N_686);
or U1382 (N_1382,N_906,N_873);
and U1383 (N_1383,N_927,N_996);
and U1384 (N_1384,N_862,N_639);
nand U1385 (N_1385,N_955,N_832);
xnor U1386 (N_1386,N_876,N_918);
or U1387 (N_1387,N_780,N_775);
and U1388 (N_1388,N_540,N_744);
and U1389 (N_1389,N_748,N_803);
and U1390 (N_1390,N_787,N_603);
and U1391 (N_1391,N_689,N_921);
and U1392 (N_1392,N_522,N_831);
and U1393 (N_1393,N_535,N_775);
nor U1394 (N_1394,N_752,N_832);
nor U1395 (N_1395,N_670,N_633);
nand U1396 (N_1396,N_630,N_911);
or U1397 (N_1397,N_767,N_719);
or U1398 (N_1398,N_664,N_899);
nand U1399 (N_1399,N_830,N_809);
or U1400 (N_1400,N_680,N_862);
and U1401 (N_1401,N_814,N_799);
nor U1402 (N_1402,N_901,N_545);
or U1403 (N_1403,N_700,N_702);
nand U1404 (N_1404,N_730,N_940);
nand U1405 (N_1405,N_857,N_563);
nand U1406 (N_1406,N_797,N_825);
nand U1407 (N_1407,N_987,N_553);
or U1408 (N_1408,N_724,N_997);
nand U1409 (N_1409,N_995,N_534);
nand U1410 (N_1410,N_523,N_873);
nand U1411 (N_1411,N_579,N_919);
xor U1412 (N_1412,N_984,N_728);
or U1413 (N_1413,N_910,N_779);
xnor U1414 (N_1414,N_500,N_988);
nand U1415 (N_1415,N_774,N_898);
nand U1416 (N_1416,N_973,N_868);
and U1417 (N_1417,N_943,N_629);
xor U1418 (N_1418,N_967,N_848);
and U1419 (N_1419,N_811,N_622);
or U1420 (N_1420,N_987,N_669);
and U1421 (N_1421,N_654,N_689);
nor U1422 (N_1422,N_723,N_606);
nor U1423 (N_1423,N_653,N_989);
xor U1424 (N_1424,N_533,N_855);
nand U1425 (N_1425,N_523,N_766);
nand U1426 (N_1426,N_813,N_844);
nor U1427 (N_1427,N_808,N_743);
and U1428 (N_1428,N_798,N_500);
or U1429 (N_1429,N_685,N_948);
nor U1430 (N_1430,N_678,N_693);
xnor U1431 (N_1431,N_515,N_730);
nand U1432 (N_1432,N_781,N_836);
nand U1433 (N_1433,N_659,N_618);
and U1434 (N_1434,N_906,N_589);
or U1435 (N_1435,N_767,N_617);
or U1436 (N_1436,N_660,N_806);
xnor U1437 (N_1437,N_654,N_817);
nand U1438 (N_1438,N_708,N_795);
and U1439 (N_1439,N_936,N_770);
nand U1440 (N_1440,N_627,N_952);
nand U1441 (N_1441,N_746,N_817);
or U1442 (N_1442,N_688,N_825);
or U1443 (N_1443,N_738,N_523);
nand U1444 (N_1444,N_677,N_852);
nor U1445 (N_1445,N_666,N_921);
and U1446 (N_1446,N_654,N_831);
xor U1447 (N_1447,N_513,N_894);
and U1448 (N_1448,N_616,N_560);
and U1449 (N_1449,N_959,N_517);
or U1450 (N_1450,N_508,N_722);
or U1451 (N_1451,N_979,N_543);
xor U1452 (N_1452,N_793,N_699);
xnor U1453 (N_1453,N_788,N_940);
nand U1454 (N_1454,N_656,N_578);
nor U1455 (N_1455,N_988,N_716);
xor U1456 (N_1456,N_870,N_841);
nor U1457 (N_1457,N_593,N_758);
nor U1458 (N_1458,N_685,N_658);
and U1459 (N_1459,N_601,N_742);
nor U1460 (N_1460,N_829,N_969);
and U1461 (N_1461,N_865,N_996);
nor U1462 (N_1462,N_723,N_513);
nand U1463 (N_1463,N_821,N_653);
or U1464 (N_1464,N_671,N_627);
nor U1465 (N_1465,N_684,N_973);
xnor U1466 (N_1466,N_651,N_671);
and U1467 (N_1467,N_838,N_816);
xnor U1468 (N_1468,N_818,N_878);
nor U1469 (N_1469,N_912,N_900);
nand U1470 (N_1470,N_953,N_542);
nor U1471 (N_1471,N_780,N_592);
or U1472 (N_1472,N_581,N_803);
and U1473 (N_1473,N_695,N_818);
or U1474 (N_1474,N_984,N_704);
and U1475 (N_1475,N_614,N_749);
nor U1476 (N_1476,N_574,N_532);
nor U1477 (N_1477,N_747,N_865);
and U1478 (N_1478,N_875,N_528);
and U1479 (N_1479,N_970,N_811);
nor U1480 (N_1480,N_750,N_657);
and U1481 (N_1481,N_947,N_604);
nand U1482 (N_1482,N_673,N_564);
nor U1483 (N_1483,N_703,N_630);
and U1484 (N_1484,N_624,N_947);
or U1485 (N_1485,N_862,N_670);
nand U1486 (N_1486,N_833,N_868);
nand U1487 (N_1487,N_923,N_702);
nand U1488 (N_1488,N_878,N_565);
or U1489 (N_1489,N_756,N_693);
nand U1490 (N_1490,N_636,N_540);
and U1491 (N_1491,N_697,N_650);
or U1492 (N_1492,N_758,N_664);
nand U1493 (N_1493,N_970,N_726);
nor U1494 (N_1494,N_956,N_738);
nand U1495 (N_1495,N_852,N_708);
and U1496 (N_1496,N_998,N_612);
nand U1497 (N_1497,N_532,N_570);
or U1498 (N_1498,N_533,N_650);
nand U1499 (N_1499,N_504,N_983);
or U1500 (N_1500,N_1342,N_1158);
and U1501 (N_1501,N_1003,N_1248);
or U1502 (N_1502,N_1262,N_1284);
nor U1503 (N_1503,N_1013,N_1153);
nand U1504 (N_1504,N_1217,N_1310);
nand U1505 (N_1505,N_1047,N_1415);
nand U1506 (N_1506,N_1497,N_1211);
nand U1507 (N_1507,N_1133,N_1467);
nand U1508 (N_1508,N_1352,N_1054);
xnor U1509 (N_1509,N_1406,N_1106);
nand U1510 (N_1510,N_1495,N_1006);
or U1511 (N_1511,N_1143,N_1256);
and U1512 (N_1512,N_1268,N_1345);
xnor U1513 (N_1513,N_1329,N_1382);
nand U1514 (N_1514,N_1420,N_1025);
or U1515 (N_1515,N_1241,N_1332);
nand U1516 (N_1516,N_1434,N_1376);
nand U1517 (N_1517,N_1028,N_1242);
or U1518 (N_1518,N_1177,N_1088);
nand U1519 (N_1519,N_1138,N_1353);
nor U1520 (N_1520,N_1094,N_1036);
nor U1521 (N_1521,N_1271,N_1404);
xor U1522 (N_1522,N_1338,N_1354);
or U1523 (N_1523,N_1289,N_1044);
nor U1524 (N_1524,N_1032,N_1431);
nand U1525 (N_1525,N_1040,N_1341);
nand U1526 (N_1526,N_1269,N_1100);
nand U1527 (N_1527,N_1232,N_1317);
or U1528 (N_1528,N_1369,N_1294);
nor U1529 (N_1529,N_1444,N_1492);
nand U1530 (N_1530,N_1461,N_1438);
nor U1531 (N_1531,N_1179,N_1280);
and U1532 (N_1532,N_1049,N_1257);
and U1533 (N_1533,N_1162,N_1334);
nor U1534 (N_1534,N_1087,N_1261);
or U1535 (N_1535,N_1286,N_1251);
nor U1536 (N_1536,N_1199,N_1163);
and U1537 (N_1537,N_1250,N_1347);
nor U1538 (N_1538,N_1074,N_1193);
nand U1539 (N_1539,N_1400,N_1195);
and U1540 (N_1540,N_1039,N_1290);
and U1541 (N_1541,N_1442,N_1010);
nand U1542 (N_1542,N_1270,N_1385);
nor U1543 (N_1543,N_1459,N_1229);
nor U1544 (N_1544,N_1455,N_1101);
nor U1545 (N_1545,N_1117,N_1204);
nor U1546 (N_1546,N_1408,N_1424);
nand U1547 (N_1547,N_1356,N_1086);
and U1548 (N_1548,N_1129,N_1246);
xnor U1549 (N_1549,N_1393,N_1165);
and U1550 (N_1550,N_1171,N_1285);
and U1551 (N_1551,N_1399,N_1125);
or U1552 (N_1552,N_1365,N_1348);
or U1553 (N_1553,N_1279,N_1389);
nor U1554 (N_1554,N_1140,N_1202);
and U1555 (N_1555,N_1330,N_1145);
or U1556 (N_1556,N_1429,N_1273);
nand U1557 (N_1557,N_1196,N_1239);
nor U1558 (N_1558,N_1346,N_1056);
and U1559 (N_1559,N_1447,N_1466);
nor U1560 (N_1560,N_1453,N_1070);
and U1561 (N_1561,N_1107,N_1333);
nor U1562 (N_1562,N_1212,N_1092);
and U1563 (N_1563,N_1157,N_1083);
or U1564 (N_1564,N_1377,N_1035);
or U1565 (N_1565,N_1433,N_1128);
nand U1566 (N_1566,N_1200,N_1343);
and U1567 (N_1567,N_1395,N_1033);
or U1568 (N_1568,N_1267,N_1413);
and U1569 (N_1569,N_1038,N_1243);
or U1570 (N_1570,N_1244,N_1476);
nand U1571 (N_1571,N_1458,N_1090);
nand U1572 (N_1572,N_1253,N_1226);
or U1573 (N_1573,N_1339,N_1115);
nand U1574 (N_1574,N_1148,N_1237);
nand U1575 (N_1575,N_1197,N_1421);
nor U1576 (N_1576,N_1015,N_1063);
xnor U1577 (N_1577,N_1309,N_1266);
nand U1578 (N_1578,N_1072,N_1020);
nand U1579 (N_1579,N_1483,N_1487);
xnor U1580 (N_1580,N_1029,N_1331);
nor U1581 (N_1581,N_1122,N_1474);
or U1582 (N_1582,N_1287,N_1045);
nor U1583 (N_1583,N_1478,N_1378);
and U1584 (N_1584,N_1323,N_1154);
xnor U1585 (N_1585,N_1223,N_1062);
nand U1586 (N_1586,N_1439,N_1392);
and U1587 (N_1587,N_1225,N_1452);
xnor U1588 (N_1588,N_1412,N_1149);
nand U1589 (N_1589,N_1141,N_1189);
nand U1590 (N_1590,N_1471,N_1077);
and U1591 (N_1591,N_1233,N_1097);
and U1592 (N_1592,N_1203,N_1186);
and U1593 (N_1593,N_1313,N_1336);
or U1594 (N_1594,N_1379,N_1367);
nand U1595 (N_1595,N_1301,N_1252);
and U1596 (N_1596,N_1238,N_1282);
nand U1597 (N_1597,N_1000,N_1052);
nor U1598 (N_1598,N_1084,N_1218);
nand U1599 (N_1599,N_1110,N_1017);
and U1600 (N_1600,N_1457,N_1118);
xor U1601 (N_1601,N_1103,N_1208);
nor U1602 (N_1602,N_1247,N_1078);
and U1603 (N_1603,N_1411,N_1430);
and U1604 (N_1604,N_1037,N_1178);
nand U1605 (N_1605,N_1009,N_1391);
or U1606 (N_1606,N_1014,N_1007);
nor U1607 (N_1607,N_1123,N_1401);
or U1608 (N_1608,N_1181,N_1245);
nor U1609 (N_1609,N_1479,N_1277);
nor U1610 (N_1610,N_1335,N_1222);
nand U1611 (N_1611,N_1394,N_1234);
or U1612 (N_1612,N_1135,N_1325);
or U1613 (N_1613,N_1364,N_1350);
or U1614 (N_1614,N_1470,N_1386);
nor U1615 (N_1615,N_1390,N_1099);
nor U1616 (N_1616,N_1283,N_1221);
or U1617 (N_1617,N_1180,N_1058);
nor U1618 (N_1618,N_1296,N_1319);
or U1619 (N_1619,N_1405,N_1236);
or U1620 (N_1620,N_1355,N_1164);
and U1621 (N_1621,N_1494,N_1201);
or U1622 (N_1622,N_1215,N_1308);
or U1623 (N_1623,N_1098,N_1051);
nand U1624 (N_1624,N_1361,N_1278);
nor U1625 (N_1625,N_1224,N_1272);
nand U1626 (N_1626,N_1344,N_1275);
nor U1627 (N_1627,N_1079,N_1360);
and U1628 (N_1628,N_1050,N_1081);
nor U1629 (N_1629,N_1060,N_1220);
and U1630 (N_1630,N_1209,N_1126);
nand U1631 (N_1631,N_1298,N_1034);
and U1632 (N_1632,N_1432,N_1303);
or U1633 (N_1633,N_1191,N_1048);
xor U1634 (N_1634,N_1291,N_1004);
or U1635 (N_1635,N_1327,N_1446);
or U1636 (N_1636,N_1228,N_1023);
nand U1637 (N_1637,N_1016,N_1198);
xnor U1638 (N_1638,N_1167,N_1407);
or U1639 (N_1639,N_1320,N_1134);
and U1640 (N_1640,N_1485,N_1136);
nand U1641 (N_1641,N_1067,N_1076);
xor U1642 (N_1642,N_1489,N_1300);
or U1643 (N_1643,N_1064,N_1417);
nor U1644 (N_1644,N_1210,N_1384);
xnor U1645 (N_1645,N_1440,N_1418);
nand U1646 (N_1646,N_1019,N_1041);
nor U1647 (N_1647,N_1147,N_1130);
nand U1648 (N_1648,N_1073,N_1185);
nand U1649 (N_1649,N_1264,N_1473);
or U1650 (N_1650,N_1441,N_1046);
nand U1651 (N_1651,N_1426,N_1435);
nor U1652 (N_1652,N_1449,N_1175);
nor U1653 (N_1653,N_1340,N_1161);
nand U1654 (N_1654,N_1091,N_1219);
nor U1655 (N_1655,N_1012,N_1055);
or U1656 (N_1656,N_1005,N_1383);
and U1657 (N_1657,N_1295,N_1159);
nand U1658 (N_1658,N_1119,N_1468);
and U1659 (N_1659,N_1469,N_1030);
nor U1660 (N_1660,N_1281,N_1465);
xor U1661 (N_1661,N_1190,N_1358);
xnor U1662 (N_1662,N_1302,N_1160);
nand U1663 (N_1663,N_1372,N_1057);
nor U1664 (N_1664,N_1463,N_1373);
xor U1665 (N_1665,N_1443,N_1374);
or U1666 (N_1666,N_1001,N_1150);
nand U1667 (N_1667,N_1416,N_1230);
nand U1668 (N_1668,N_1397,N_1318);
nor U1669 (N_1669,N_1305,N_1255);
nand U1670 (N_1670,N_1089,N_1486);
nand U1671 (N_1671,N_1113,N_1192);
and U1672 (N_1672,N_1328,N_1460);
nor U1673 (N_1673,N_1182,N_1349);
or U1674 (N_1674,N_1075,N_1065);
xnor U1675 (N_1675,N_1082,N_1357);
nor U1676 (N_1676,N_1214,N_1425);
nor U1677 (N_1677,N_1121,N_1152);
nor U1678 (N_1678,N_1370,N_1423);
nand U1679 (N_1679,N_1464,N_1388);
nand U1680 (N_1680,N_1368,N_1324);
or U1681 (N_1681,N_1096,N_1022);
nand U1682 (N_1682,N_1205,N_1381);
and U1683 (N_1683,N_1026,N_1169);
or U1684 (N_1684,N_1496,N_1166);
nor U1685 (N_1685,N_1151,N_1396);
and U1686 (N_1686,N_1366,N_1254);
nor U1687 (N_1687,N_1482,N_1448);
xnor U1688 (N_1688,N_1375,N_1297);
nand U1689 (N_1689,N_1231,N_1306);
or U1690 (N_1690,N_1174,N_1498);
nand U1691 (N_1691,N_1351,N_1337);
nor U1692 (N_1692,N_1315,N_1168);
or U1693 (N_1693,N_1428,N_1265);
and U1694 (N_1694,N_1488,N_1419);
or U1695 (N_1695,N_1027,N_1363);
xor U1696 (N_1696,N_1227,N_1112);
xor U1697 (N_1697,N_1093,N_1146);
and U1698 (N_1698,N_1484,N_1475);
nand U1699 (N_1699,N_1116,N_1131);
nand U1700 (N_1700,N_1207,N_1276);
or U1701 (N_1701,N_1462,N_1480);
nand U1702 (N_1702,N_1206,N_1491);
nor U1703 (N_1703,N_1316,N_1002);
or U1704 (N_1704,N_1059,N_1410);
and U1705 (N_1705,N_1042,N_1304);
nor U1706 (N_1706,N_1021,N_1155);
or U1707 (N_1707,N_1362,N_1326);
or U1708 (N_1708,N_1144,N_1111);
nor U1709 (N_1709,N_1031,N_1445);
nor U1710 (N_1710,N_1371,N_1490);
nor U1711 (N_1711,N_1477,N_1137);
nand U1712 (N_1712,N_1071,N_1322);
nor U1713 (N_1713,N_1437,N_1321);
nand U1714 (N_1714,N_1293,N_1085);
and U1715 (N_1715,N_1108,N_1259);
nor U1716 (N_1716,N_1450,N_1194);
or U1717 (N_1717,N_1249,N_1176);
and U1718 (N_1718,N_1080,N_1314);
xor U1719 (N_1719,N_1139,N_1102);
nand U1720 (N_1720,N_1451,N_1008);
or U1721 (N_1721,N_1359,N_1053);
or U1722 (N_1722,N_1061,N_1312);
and U1723 (N_1723,N_1018,N_1311);
and U1724 (N_1724,N_1120,N_1114);
nor U1725 (N_1725,N_1456,N_1307);
nand U1726 (N_1726,N_1235,N_1170);
xnor U1727 (N_1727,N_1403,N_1499);
nand U1728 (N_1728,N_1240,N_1024);
nand U1729 (N_1729,N_1402,N_1213);
nand U1730 (N_1730,N_1493,N_1066);
nand U1731 (N_1731,N_1260,N_1188);
nand U1732 (N_1732,N_1069,N_1292);
or U1733 (N_1733,N_1187,N_1068);
and U1734 (N_1734,N_1409,N_1109);
or U1735 (N_1735,N_1216,N_1184);
and U1736 (N_1736,N_1436,N_1454);
xor U1737 (N_1737,N_1258,N_1472);
and U1738 (N_1738,N_1481,N_1299);
nor U1739 (N_1739,N_1263,N_1043);
nor U1740 (N_1740,N_1127,N_1142);
nand U1741 (N_1741,N_1172,N_1274);
and U1742 (N_1742,N_1173,N_1422);
nor U1743 (N_1743,N_1183,N_1132);
nor U1744 (N_1744,N_1380,N_1011);
and U1745 (N_1745,N_1387,N_1124);
nand U1746 (N_1746,N_1104,N_1414);
and U1747 (N_1747,N_1095,N_1288);
nand U1748 (N_1748,N_1398,N_1427);
and U1749 (N_1749,N_1105,N_1156);
nor U1750 (N_1750,N_1226,N_1012);
nand U1751 (N_1751,N_1251,N_1182);
nor U1752 (N_1752,N_1343,N_1494);
and U1753 (N_1753,N_1400,N_1138);
or U1754 (N_1754,N_1207,N_1099);
or U1755 (N_1755,N_1480,N_1119);
nor U1756 (N_1756,N_1357,N_1094);
or U1757 (N_1757,N_1067,N_1246);
nor U1758 (N_1758,N_1255,N_1245);
nand U1759 (N_1759,N_1132,N_1362);
and U1760 (N_1760,N_1026,N_1433);
and U1761 (N_1761,N_1347,N_1096);
xor U1762 (N_1762,N_1269,N_1258);
nand U1763 (N_1763,N_1083,N_1127);
or U1764 (N_1764,N_1211,N_1251);
xor U1765 (N_1765,N_1126,N_1098);
nand U1766 (N_1766,N_1192,N_1067);
or U1767 (N_1767,N_1487,N_1204);
nor U1768 (N_1768,N_1014,N_1179);
nor U1769 (N_1769,N_1157,N_1338);
nor U1770 (N_1770,N_1157,N_1006);
xor U1771 (N_1771,N_1263,N_1226);
or U1772 (N_1772,N_1339,N_1045);
nor U1773 (N_1773,N_1107,N_1351);
or U1774 (N_1774,N_1445,N_1165);
or U1775 (N_1775,N_1212,N_1221);
nor U1776 (N_1776,N_1054,N_1034);
nand U1777 (N_1777,N_1406,N_1313);
or U1778 (N_1778,N_1405,N_1259);
nand U1779 (N_1779,N_1010,N_1454);
or U1780 (N_1780,N_1268,N_1184);
xnor U1781 (N_1781,N_1261,N_1329);
nor U1782 (N_1782,N_1462,N_1042);
or U1783 (N_1783,N_1378,N_1131);
nand U1784 (N_1784,N_1156,N_1255);
or U1785 (N_1785,N_1368,N_1439);
xor U1786 (N_1786,N_1056,N_1044);
nor U1787 (N_1787,N_1345,N_1065);
and U1788 (N_1788,N_1290,N_1303);
or U1789 (N_1789,N_1344,N_1400);
and U1790 (N_1790,N_1169,N_1293);
nand U1791 (N_1791,N_1235,N_1429);
nand U1792 (N_1792,N_1334,N_1399);
nand U1793 (N_1793,N_1473,N_1005);
or U1794 (N_1794,N_1196,N_1435);
nor U1795 (N_1795,N_1070,N_1032);
nor U1796 (N_1796,N_1340,N_1279);
and U1797 (N_1797,N_1061,N_1492);
or U1798 (N_1798,N_1353,N_1197);
and U1799 (N_1799,N_1403,N_1250);
nand U1800 (N_1800,N_1324,N_1058);
nor U1801 (N_1801,N_1372,N_1454);
xor U1802 (N_1802,N_1411,N_1109);
nand U1803 (N_1803,N_1401,N_1211);
or U1804 (N_1804,N_1276,N_1432);
or U1805 (N_1805,N_1332,N_1046);
or U1806 (N_1806,N_1406,N_1155);
nor U1807 (N_1807,N_1018,N_1325);
nor U1808 (N_1808,N_1069,N_1071);
and U1809 (N_1809,N_1387,N_1430);
and U1810 (N_1810,N_1276,N_1314);
and U1811 (N_1811,N_1268,N_1258);
nor U1812 (N_1812,N_1045,N_1241);
nand U1813 (N_1813,N_1188,N_1386);
xor U1814 (N_1814,N_1421,N_1067);
nand U1815 (N_1815,N_1440,N_1067);
or U1816 (N_1816,N_1281,N_1106);
or U1817 (N_1817,N_1040,N_1398);
or U1818 (N_1818,N_1411,N_1205);
and U1819 (N_1819,N_1195,N_1333);
and U1820 (N_1820,N_1070,N_1100);
nand U1821 (N_1821,N_1474,N_1453);
nand U1822 (N_1822,N_1390,N_1027);
or U1823 (N_1823,N_1268,N_1419);
xor U1824 (N_1824,N_1151,N_1315);
xnor U1825 (N_1825,N_1135,N_1446);
nor U1826 (N_1826,N_1120,N_1122);
nand U1827 (N_1827,N_1089,N_1293);
nand U1828 (N_1828,N_1104,N_1120);
nor U1829 (N_1829,N_1467,N_1366);
nand U1830 (N_1830,N_1132,N_1486);
or U1831 (N_1831,N_1213,N_1154);
or U1832 (N_1832,N_1464,N_1417);
or U1833 (N_1833,N_1306,N_1114);
nor U1834 (N_1834,N_1322,N_1424);
xnor U1835 (N_1835,N_1060,N_1294);
nor U1836 (N_1836,N_1092,N_1140);
or U1837 (N_1837,N_1190,N_1285);
or U1838 (N_1838,N_1281,N_1080);
xor U1839 (N_1839,N_1038,N_1335);
nor U1840 (N_1840,N_1341,N_1073);
and U1841 (N_1841,N_1439,N_1300);
nand U1842 (N_1842,N_1273,N_1115);
or U1843 (N_1843,N_1423,N_1337);
or U1844 (N_1844,N_1003,N_1193);
or U1845 (N_1845,N_1325,N_1118);
and U1846 (N_1846,N_1458,N_1183);
nor U1847 (N_1847,N_1367,N_1084);
nand U1848 (N_1848,N_1029,N_1483);
nand U1849 (N_1849,N_1229,N_1058);
and U1850 (N_1850,N_1483,N_1424);
or U1851 (N_1851,N_1179,N_1438);
or U1852 (N_1852,N_1260,N_1066);
and U1853 (N_1853,N_1136,N_1034);
and U1854 (N_1854,N_1489,N_1461);
nor U1855 (N_1855,N_1235,N_1182);
nor U1856 (N_1856,N_1000,N_1207);
nand U1857 (N_1857,N_1249,N_1017);
nor U1858 (N_1858,N_1034,N_1177);
nor U1859 (N_1859,N_1153,N_1028);
xnor U1860 (N_1860,N_1111,N_1310);
xor U1861 (N_1861,N_1117,N_1055);
nand U1862 (N_1862,N_1248,N_1165);
nor U1863 (N_1863,N_1181,N_1016);
and U1864 (N_1864,N_1215,N_1460);
and U1865 (N_1865,N_1467,N_1443);
nand U1866 (N_1866,N_1090,N_1188);
and U1867 (N_1867,N_1218,N_1311);
and U1868 (N_1868,N_1212,N_1466);
and U1869 (N_1869,N_1048,N_1482);
or U1870 (N_1870,N_1059,N_1320);
or U1871 (N_1871,N_1144,N_1397);
and U1872 (N_1872,N_1045,N_1407);
or U1873 (N_1873,N_1031,N_1122);
and U1874 (N_1874,N_1019,N_1451);
xnor U1875 (N_1875,N_1172,N_1324);
and U1876 (N_1876,N_1213,N_1167);
and U1877 (N_1877,N_1250,N_1342);
xor U1878 (N_1878,N_1267,N_1339);
nand U1879 (N_1879,N_1149,N_1188);
nor U1880 (N_1880,N_1074,N_1087);
nor U1881 (N_1881,N_1295,N_1206);
xor U1882 (N_1882,N_1383,N_1361);
nand U1883 (N_1883,N_1450,N_1039);
nand U1884 (N_1884,N_1224,N_1411);
or U1885 (N_1885,N_1155,N_1482);
or U1886 (N_1886,N_1492,N_1385);
nor U1887 (N_1887,N_1386,N_1116);
nand U1888 (N_1888,N_1371,N_1480);
and U1889 (N_1889,N_1171,N_1265);
xnor U1890 (N_1890,N_1240,N_1006);
nor U1891 (N_1891,N_1230,N_1478);
and U1892 (N_1892,N_1157,N_1206);
and U1893 (N_1893,N_1356,N_1352);
nor U1894 (N_1894,N_1307,N_1118);
or U1895 (N_1895,N_1143,N_1271);
and U1896 (N_1896,N_1495,N_1183);
nand U1897 (N_1897,N_1318,N_1051);
or U1898 (N_1898,N_1084,N_1119);
nand U1899 (N_1899,N_1389,N_1305);
nand U1900 (N_1900,N_1454,N_1398);
nand U1901 (N_1901,N_1101,N_1235);
xor U1902 (N_1902,N_1077,N_1090);
or U1903 (N_1903,N_1031,N_1141);
nor U1904 (N_1904,N_1121,N_1352);
nand U1905 (N_1905,N_1299,N_1490);
or U1906 (N_1906,N_1255,N_1486);
nand U1907 (N_1907,N_1074,N_1222);
or U1908 (N_1908,N_1206,N_1253);
or U1909 (N_1909,N_1058,N_1221);
nand U1910 (N_1910,N_1453,N_1144);
nor U1911 (N_1911,N_1063,N_1085);
nand U1912 (N_1912,N_1045,N_1208);
or U1913 (N_1913,N_1225,N_1203);
nand U1914 (N_1914,N_1392,N_1243);
nor U1915 (N_1915,N_1304,N_1164);
and U1916 (N_1916,N_1257,N_1182);
xnor U1917 (N_1917,N_1436,N_1066);
nor U1918 (N_1918,N_1137,N_1144);
nor U1919 (N_1919,N_1004,N_1471);
nand U1920 (N_1920,N_1120,N_1280);
nor U1921 (N_1921,N_1385,N_1366);
nand U1922 (N_1922,N_1399,N_1017);
or U1923 (N_1923,N_1060,N_1466);
or U1924 (N_1924,N_1353,N_1214);
and U1925 (N_1925,N_1231,N_1193);
nand U1926 (N_1926,N_1399,N_1251);
nand U1927 (N_1927,N_1002,N_1200);
nor U1928 (N_1928,N_1306,N_1442);
nand U1929 (N_1929,N_1051,N_1192);
nand U1930 (N_1930,N_1399,N_1295);
or U1931 (N_1931,N_1414,N_1357);
or U1932 (N_1932,N_1376,N_1370);
or U1933 (N_1933,N_1037,N_1089);
and U1934 (N_1934,N_1439,N_1183);
or U1935 (N_1935,N_1058,N_1371);
nand U1936 (N_1936,N_1454,N_1452);
nor U1937 (N_1937,N_1161,N_1327);
or U1938 (N_1938,N_1378,N_1046);
nor U1939 (N_1939,N_1044,N_1450);
nand U1940 (N_1940,N_1321,N_1252);
or U1941 (N_1941,N_1277,N_1148);
and U1942 (N_1942,N_1119,N_1435);
nor U1943 (N_1943,N_1076,N_1294);
or U1944 (N_1944,N_1481,N_1028);
xnor U1945 (N_1945,N_1347,N_1310);
nor U1946 (N_1946,N_1471,N_1407);
nand U1947 (N_1947,N_1116,N_1073);
xnor U1948 (N_1948,N_1330,N_1430);
nor U1949 (N_1949,N_1163,N_1017);
and U1950 (N_1950,N_1469,N_1395);
nor U1951 (N_1951,N_1229,N_1131);
nor U1952 (N_1952,N_1071,N_1045);
or U1953 (N_1953,N_1126,N_1393);
xor U1954 (N_1954,N_1384,N_1073);
nand U1955 (N_1955,N_1166,N_1362);
nand U1956 (N_1956,N_1128,N_1077);
nand U1957 (N_1957,N_1130,N_1048);
nand U1958 (N_1958,N_1484,N_1364);
xnor U1959 (N_1959,N_1214,N_1343);
and U1960 (N_1960,N_1394,N_1404);
or U1961 (N_1961,N_1222,N_1220);
nand U1962 (N_1962,N_1318,N_1439);
or U1963 (N_1963,N_1234,N_1157);
nand U1964 (N_1964,N_1432,N_1127);
or U1965 (N_1965,N_1043,N_1380);
nand U1966 (N_1966,N_1012,N_1299);
or U1967 (N_1967,N_1159,N_1184);
nor U1968 (N_1968,N_1042,N_1433);
or U1969 (N_1969,N_1483,N_1167);
nor U1970 (N_1970,N_1464,N_1493);
nand U1971 (N_1971,N_1362,N_1047);
or U1972 (N_1972,N_1350,N_1132);
and U1973 (N_1973,N_1321,N_1494);
nor U1974 (N_1974,N_1295,N_1042);
nor U1975 (N_1975,N_1160,N_1457);
or U1976 (N_1976,N_1055,N_1053);
nand U1977 (N_1977,N_1239,N_1306);
nand U1978 (N_1978,N_1330,N_1065);
or U1979 (N_1979,N_1190,N_1101);
nand U1980 (N_1980,N_1275,N_1326);
nor U1981 (N_1981,N_1296,N_1250);
and U1982 (N_1982,N_1023,N_1229);
nor U1983 (N_1983,N_1396,N_1487);
and U1984 (N_1984,N_1176,N_1032);
nand U1985 (N_1985,N_1382,N_1126);
and U1986 (N_1986,N_1331,N_1262);
nand U1987 (N_1987,N_1078,N_1197);
nand U1988 (N_1988,N_1016,N_1089);
nor U1989 (N_1989,N_1482,N_1435);
xor U1990 (N_1990,N_1014,N_1068);
and U1991 (N_1991,N_1041,N_1247);
nand U1992 (N_1992,N_1157,N_1023);
nand U1993 (N_1993,N_1397,N_1082);
nand U1994 (N_1994,N_1288,N_1000);
and U1995 (N_1995,N_1152,N_1353);
nand U1996 (N_1996,N_1125,N_1227);
and U1997 (N_1997,N_1066,N_1267);
nand U1998 (N_1998,N_1098,N_1023);
or U1999 (N_1999,N_1267,N_1376);
xor U2000 (N_2000,N_1684,N_1624);
nor U2001 (N_2001,N_1846,N_1770);
nand U2002 (N_2002,N_1735,N_1821);
nand U2003 (N_2003,N_1849,N_1960);
xor U2004 (N_2004,N_1566,N_1513);
and U2005 (N_2005,N_1810,N_1549);
or U2006 (N_2006,N_1812,N_1948);
xor U2007 (N_2007,N_1608,N_1522);
and U2008 (N_2008,N_1905,N_1583);
and U2009 (N_2009,N_1701,N_1896);
nor U2010 (N_2010,N_1628,N_1559);
nor U2011 (N_2011,N_1553,N_1520);
or U2012 (N_2012,N_1723,N_1973);
or U2013 (N_2013,N_1502,N_1994);
and U2014 (N_2014,N_1571,N_1681);
nor U2015 (N_2015,N_1825,N_1858);
or U2016 (N_2016,N_1534,N_1861);
nor U2017 (N_2017,N_1878,N_1646);
and U2018 (N_2018,N_1840,N_1610);
nor U2019 (N_2019,N_1658,N_1511);
nor U2020 (N_2020,N_1990,N_1563);
nand U2021 (N_2021,N_1989,N_1816);
and U2022 (N_2022,N_1867,N_1524);
or U2023 (N_2023,N_1761,N_1817);
and U2024 (N_2024,N_1804,N_1565);
nor U2025 (N_2025,N_1737,N_1977);
or U2026 (N_2026,N_1712,N_1556);
nor U2027 (N_2027,N_1783,N_1983);
nand U2028 (N_2028,N_1743,N_1791);
nor U2029 (N_2029,N_1668,N_1677);
and U2030 (N_2030,N_1719,N_1865);
nor U2031 (N_2031,N_1580,N_1777);
nor U2032 (N_2032,N_1708,N_1975);
nand U2033 (N_2033,N_1922,N_1870);
nand U2034 (N_2034,N_1699,N_1730);
and U2035 (N_2035,N_1531,N_1798);
nand U2036 (N_2036,N_1614,N_1832);
or U2037 (N_2037,N_1823,N_1724);
xnor U2038 (N_2038,N_1954,N_1796);
nand U2039 (N_2039,N_1753,N_1733);
or U2040 (N_2040,N_1956,N_1911);
and U2041 (N_2041,N_1898,N_1696);
and U2042 (N_2042,N_1551,N_1751);
nand U2043 (N_2043,N_1933,N_1567);
and U2044 (N_2044,N_1711,N_1670);
nor U2045 (N_2045,N_1820,N_1797);
nor U2046 (N_2046,N_1931,N_1962);
and U2047 (N_2047,N_1585,N_1609);
and U2048 (N_2048,N_1885,N_1899);
nor U2049 (N_2049,N_1757,N_1533);
or U2050 (N_2050,N_1717,N_1809);
nor U2051 (N_2051,N_1795,N_1833);
nand U2052 (N_2052,N_1845,N_1987);
nor U2053 (N_2053,N_1946,N_1768);
or U2054 (N_2054,N_1552,N_1572);
nor U2055 (N_2055,N_1710,N_1790);
nor U2056 (N_2056,N_1625,N_1961);
nand U2057 (N_2057,N_1864,N_1852);
nor U2058 (N_2058,N_1607,N_1755);
and U2059 (N_2059,N_1574,N_1792);
nor U2060 (N_2060,N_1655,N_1665);
nor U2061 (N_2061,N_1857,N_1603);
nand U2062 (N_2062,N_1651,N_1635);
and U2063 (N_2063,N_1758,N_1843);
nand U2064 (N_2064,N_1570,N_1813);
and U2065 (N_2065,N_1507,N_1588);
and U2066 (N_2066,N_1561,N_1965);
nor U2067 (N_2067,N_1675,N_1526);
nor U2068 (N_2068,N_1891,N_1660);
nand U2069 (N_2069,N_1537,N_1914);
xnor U2070 (N_2070,N_1974,N_1606);
and U2071 (N_2071,N_1872,N_1506);
xor U2072 (N_2072,N_1985,N_1998);
nand U2073 (N_2073,N_1692,N_1540);
xnor U2074 (N_2074,N_1923,N_1634);
xnor U2075 (N_2075,N_1640,N_1890);
nor U2076 (N_2076,N_1579,N_1638);
nand U2077 (N_2077,N_1765,N_1767);
and U2078 (N_2078,N_1969,N_1562);
nor U2079 (N_2079,N_1793,N_1676);
and U2080 (N_2080,N_1882,N_1532);
nor U2081 (N_2081,N_1869,N_1672);
or U2082 (N_2082,N_1970,N_1953);
and U2083 (N_2083,N_1913,N_1966);
nor U2084 (N_2084,N_1955,N_1822);
or U2085 (N_2085,N_1764,N_1666);
and U2086 (N_2086,N_1678,N_1824);
and U2087 (N_2087,N_1976,N_1988);
nand U2088 (N_2088,N_1694,N_1829);
nand U2089 (N_2089,N_1863,N_1859);
and U2090 (N_2090,N_1721,N_1952);
and U2091 (N_2091,N_1695,N_1643);
or U2092 (N_2092,N_1892,N_1661);
or U2093 (N_2093,N_1957,N_1926);
or U2094 (N_2094,N_1741,N_1541);
nor U2095 (N_2095,N_1932,N_1999);
or U2096 (N_2096,N_1910,N_1577);
nor U2097 (N_2097,N_1853,N_1897);
or U2098 (N_2098,N_1831,N_1727);
nand U2099 (N_2099,N_1828,N_1653);
or U2100 (N_2100,N_1802,N_1544);
and U2101 (N_2101,N_1584,N_1545);
nand U2102 (N_2102,N_1862,N_1629);
and U2103 (N_2103,N_1698,N_1763);
nor U2104 (N_2104,N_1980,N_1877);
or U2105 (N_2105,N_1903,N_1729);
or U2106 (N_2106,N_1842,N_1601);
or U2107 (N_2107,N_1978,N_1801);
and U2108 (N_2108,N_1972,N_1787);
and U2109 (N_2109,N_1568,N_1742);
nand U2110 (N_2110,N_1554,N_1641);
and U2111 (N_2111,N_1928,N_1659);
xor U2112 (N_2112,N_1766,N_1748);
or U2113 (N_2113,N_1871,N_1731);
nor U2114 (N_2114,N_1626,N_1738);
nand U2115 (N_2115,N_1967,N_1535);
or U2116 (N_2116,N_1819,N_1868);
nand U2117 (N_2117,N_1652,N_1908);
nor U2118 (N_2118,N_1774,N_1686);
xnor U2119 (N_2119,N_1647,N_1521);
and U2120 (N_2120,N_1781,N_1935);
or U2121 (N_2121,N_1620,N_1664);
and U2122 (N_2122,N_1945,N_1778);
or U2123 (N_2123,N_1762,N_1706);
and U2124 (N_2124,N_1780,N_1599);
or U2125 (N_2125,N_1744,N_1505);
and U2126 (N_2126,N_1848,N_1503);
or U2127 (N_2127,N_1662,N_1622);
and U2128 (N_2128,N_1683,N_1939);
nor U2129 (N_2129,N_1907,N_1916);
or U2130 (N_2130,N_1573,N_1514);
nand U2131 (N_2131,N_1516,N_1656);
or U2132 (N_2132,N_1979,N_1673);
or U2133 (N_2133,N_1631,N_1538);
nor U2134 (N_2134,N_1720,N_1806);
and U2135 (N_2135,N_1648,N_1779);
or U2136 (N_2136,N_1611,N_1587);
nor U2137 (N_2137,N_1536,N_1927);
xor U2138 (N_2138,N_1800,N_1598);
nor U2139 (N_2139,N_1938,N_1918);
nand U2140 (N_2140,N_1834,N_1886);
nand U2141 (N_2141,N_1616,N_1942);
and U2142 (N_2142,N_1995,N_1936);
or U2143 (N_2143,N_1997,N_1924);
and U2144 (N_2144,N_1700,N_1900);
or U2145 (N_2145,N_1595,N_1504);
nor U2146 (N_2146,N_1881,N_1794);
xnor U2147 (N_2147,N_1838,N_1725);
nor U2148 (N_2148,N_1591,N_1688);
nor U2149 (N_2149,N_1645,N_1959);
nor U2150 (N_2150,N_1940,N_1887);
xnor U2151 (N_2151,N_1736,N_1600);
nand U2152 (N_2152,N_1732,N_1826);
nand U2153 (N_2153,N_1917,N_1811);
nor U2154 (N_2154,N_1746,N_1951);
and U2155 (N_2155,N_1803,N_1623);
or U2156 (N_2156,N_1508,N_1921);
nand U2157 (N_2157,N_1636,N_1697);
or U2158 (N_2158,N_1747,N_1775);
nor U2159 (N_2159,N_1714,N_1884);
xnor U2160 (N_2160,N_1739,N_1654);
and U2161 (N_2161,N_1944,N_1612);
xnor U2162 (N_2162,N_1934,N_1754);
nand U2163 (N_2163,N_1740,N_1937);
or U2164 (N_2164,N_1771,N_1992);
nor U2165 (N_2165,N_1749,N_1847);
and U2166 (N_2166,N_1875,N_1509);
nor U2167 (N_2167,N_1642,N_1958);
and U2168 (N_2168,N_1830,N_1663);
and U2169 (N_2169,N_1680,N_1617);
or U2170 (N_2170,N_1690,N_1582);
nor U2171 (N_2171,N_1964,N_1734);
or U2172 (N_2172,N_1947,N_1703);
or U2173 (N_2173,N_1873,N_1557);
nand U2174 (N_2174,N_1715,N_1895);
or U2175 (N_2175,N_1827,N_1605);
and U2176 (N_2176,N_1968,N_1604);
nand U2177 (N_2177,N_1630,N_1915);
xor U2178 (N_2178,N_1799,N_1518);
nor U2179 (N_2179,N_1836,N_1860);
nand U2180 (N_2180,N_1888,N_1685);
nor U2181 (N_2181,N_1594,N_1578);
nand U2182 (N_2182,N_1618,N_1613);
or U2183 (N_2183,N_1707,N_1632);
nor U2184 (N_2184,N_1991,N_1909);
or U2185 (N_2185,N_1805,N_1726);
xnor U2186 (N_2186,N_1691,N_1602);
nor U2187 (N_2187,N_1519,N_1550);
nand U2188 (N_2188,N_1621,N_1713);
xnor U2189 (N_2189,N_1906,N_1704);
xor U2190 (N_2190,N_1589,N_1784);
nand U2191 (N_2191,N_1528,N_1530);
nand U2192 (N_2192,N_1889,N_1527);
nor U2193 (N_2193,N_1639,N_1785);
and U2194 (N_2194,N_1709,N_1716);
nand U2195 (N_2195,N_1941,N_1650);
nand U2196 (N_2196,N_1543,N_1950);
or U2197 (N_2197,N_1517,N_1593);
and U2198 (N_2198,N_1649,N_1548);
and U2199 (N_2199,N_1856,N_1682);
nor U2200 (N_2200,N_1515,N_1745);
and U2201 (N_2201,N_1510,N_1689);
nor U2202 (N_2202,N_1525,N_1949);
nand U2203 (N_2203,N_1564,N_1679);
or U2204 (N_2204,N_1523,N_1883);
xor U2205 (N_2205,N_1808,N_1818);
nor U2206 (N_2206,N_1841,N_1837);
or U2207 (N_2207,N_1560,N_1788);
nor U2208 (N_2208,N_1904,N_1993);
and U2209 (N_2209,N_1986,N_1971);
nand U2210 (N_2210,N_1912,N_1529);
nor U2211 (N_2211,N_1996,N_1773);
nand U2212 (N_2212,N_1547,N_1671);
and U2213 (N_2213,N_1718,N_1592);
and U2214 (N_2214,N_1637,N_1512);
and U2215 (N_2215,N_1558,N_1876);
nand U2216 (N_2216,N_1728,N_1919);
or U2217 (N_2217,N_1880,N_1879);
nand U2218 (N_2218,N_1929,N_1644);
nand U2219 (N_2219,N_1866,N_1657);
nor U2220 (N_2220,N_1586,N_1615);
or U2221 (N_2221,N_1501,N_1555);
nand U2222 (N_2222,N_1569,N_1815);
and U2223 (N_2223,N_1542,N_1575);
xor U2224 (N_2224,N_1669,N_1789);
nand U2225 (N_2225,N_1854,N_1590);
nor U2226 (N_2226,N_1851,N_1687);
xor U2227 (N_2227,N_1667,N_1920);
nor U2228 (N_2228,N_1839,N_1925);
and U2229 (N_2229,N_1814,N_1981);
nand U2230 (N_2230,N_1752,N_1894);
and U2231 (N_2231,N_1769,N_1930);
and U2232 (N_2232,N_1943,N_1902);
xnor U2233 (N_2233,N_1850,N_1756);
nor U2234 (N_2234,N_1705,N_1893);
nand U2235 (N_2235,N_1901,N_1807);
and U2236 (N_2236,N_1627,N_1772);
and U2237 (N_2237,N_1874,N_1855);
nor U2238 (N_2238,N_1633,N_1702);
nand U2239 (N_2239,N_1546,N_1782);
or U2240 (N_2240,N_1500,N_1759);
nand U2241 (N_2241,N_1619,N_1576);
xor U2242 (N_2242,N_1776,N_1596);
and U2243 (N_2243,N_1835,N_1539);
xnor U2244 (N_2244,N_1963,N_1722);
nand U2245 (N_2245,N_1984,N_1750);
nand U2246 (N_2246,N_1844,N_1693);
and U2247 (N_2247,N_1597,N_1982);
and U2248 (N_2248,N_1674,N_1581);
and U2249 (N_2249,N_1760,N_1786);
nand U2250 (N_2250,N_1701,N_1686);
nand U2251 (N_2251,N_1965,N_1550);
and U2252 (N_2252,N_1604,N_1986);
nand U2253 (N_2253,N_1952,N_1648);
nand U2254 (N_2254,N_1626,N_1574);
or U2255 (N_2255,N_1674,N_1609);
nor U2256 (N_2256,N_1828,N_1701);
and U2257 (N_2257,N_1986,N_1610);
nand U2258 (N_2258,N_1652,N_1854);
nor U2259 (N_2259,N_1547,N_1827);
and U2260 (N_2260,N_1940,N_1584);
or U2261 (N_2261,N_1974,N_1815);
or U2262 (N_2262,N_1743,N_1723);
nand U2263 (N_2263,N_1802,N_1906);
nand U2264 (N_2264,N_1534,N_1662);
and U2265 (N_2265,N_1700,N_1539);
nor U2266 (N_2266,N_1573,N_1740);
xnor U2267 (N_2267,N_1523,N_1970);
xnor U2268 (N_2268,N_1729,N_1782);
or U2269 (N_2269,N_1570,N_1999);
and U2270 (N_2270,N_1911,N_1670);
nor U2271 (N_2271,N_1602,N_1913);
nor U2272 (N_2272,N_1936,N_1700);
nand U2273 (N_2273,N_1800,N_1734);
and U2274 (N_2274,N_1616,N_1945);
or U2275 (N_2275,N_1940,N_1872);
nor U2276 (N_2276,N_1943,N_1649);
or U2277 (N_2277,N_1571,N_1741);
nor U2278 (N_2278,N_1555,N_1533);
nor U2279 (N_2279,N_1712,N_1951);
nand U2280 (N_2280,N_1538,N_1548);
nand U2281 (N_2281,N_1820,N_1823);
and U2282 (N_2282,N_1708,N_1510);
and U2283 (N_2283,N_1558,N_1864);
or U2284 (N_2284,N_1605,N_1996);
nand U2285 (N_2285,N_1570,N_1600);
nor U2286 (N_2286,N_1715,N_1827);
or U2287 (N_2287,N_1660,N_1541);
nor U2288 (N_2288,N_1576,N_1590);
and U2289 (N_2289,N_1615,N_1578);
and U2290 (N_2290,N_1594,N_1882);
and U2291 (N_2291,N_1982,N_1989);
nor U2292 (N_2292,N_1564,N_1723);
nor U2293 (N_2293,N_1813,N_1801);
or U2294 (N_2294,N_1599,N_1637);
nor U2295 (N_2295,N_1910,N_1786);
nand U2296 (N_2296,N_1789,N_1684);
and U2297 (N_2297,N_1804,N_1781);
nor U2298 (N_2298,N_1897,N_1726);
and U2299 (N_2299,N_1723,N_1557);
and U2300 (N_2300,N_1867,N_1560);
nand U2301 (N_2301,N_1684,N_1753);
and U2302 (N_2302,N_1750,N_1841);
nand U2303 (N_2303,N_1769,N_1895);
nor U2304 (N_2304,N_1514,N_1689);
nand U2305 (N_2305,N_1796,N_1792);
nand U2306 (N_2306,N_1672,N_1681);
nand U2307 (N_2307,N_1919,N_1842);
or U2308 (N_2308,N_1560,N_1759);
and U2309 (N_2309,N_1535,N_1998);
nor U2310 (N_2310,N_1826,N_1718);
nor U2311 (N_2311,N_1543,N_1629);
and U2312 (N_2312,N_1957,N_1614);
or U2313 (N_2313,N_1791,N_1704);
or U2314 (N_2314,N_1718,N_1635);
nor U2315 (N_2315,N_1986,N_1724);
or U2316 (N_2316,N_1842,N_1612);
nand U2317 (N_2317,N_1869,N_1668);
nand U2318 (N_2318,N_1839,N_1711);
and U2319 (N_2319,N_1797,N_1913);
and U2320 (N_2320,N_1830,N_1870);
nand U2321 (N_2321,N_1756,N_1705);
nor U2322 (N_2322,N_1890,N_1528);
and U2323 (N_2323,N_1702,N_1801);
nor U2324 (N_2324,N_1841,N_1730);
nor U2325 (N_2325,N_1596,N_1950);
and U2326 (N_2326,N_1933,N_1947);
xor U2327 (N_2327,N_1524,N_1573);
and U2328 (N_2328,N_1864,N_1715);
or U2329 (N_2329,N_1961,N_1602);
and U2330 (N_2330,N_1897,N_1995);
or U2331 (N_2331,N_1634,N_1515);
nand U2332 (N_2332,N_1595,N_1521);
and U2333 (N_2333,N_1657,N_1841);
nand U2334 (N_2334,N_1736,N_1717);
nand U2335 (N_2335,N_1645,N_1797);
and U2336 (N_2336,N_1943,N_1508);
nand U2337 (N_2337,N_1873,N_1765);
nor U2338 (N_2338,N_1828,N_1967);
or U2339 (N_2339,N_1902,N_1950);
and U2340 (N_2340,N_1877,N_1679);
or U2341 (N_2341,N_1624,N_1930);
and U2342 (N_2342,N_1556,N_1611);
nand U2343 (N_2343,N_1736,N_1761);
or U2344 (N_2344,N_1763,N_1886);
and U2345 (N_2345,N_1929,N_1721);
and U2346 (N_2346,N_1674,N_1729);
and U2347 (N_2347,N_1513,N_1577);
and U2348 (N_2348,N_1981,N_1534);
nand U2349 (N_2349,N_1666,N_1911);
or U2350 (N_2350,N_1636,N_1535);
and U2351 (N_2351,N_1904,N_1776);
and U2352 (N_2352,N_1756,N_1626);
nand U2353 (N_2353,N_1681,N_1581);
nor U2354 (N_2354,N_1505,N_1518);
xnor U2355 (N_2355,N_1776,N_1885);
nand U2356 (N_2356,N_1854,N_1529);
nor U2357 (N_2357,N_1613,N_1932);
xnor U2358 (N_2358,N_1826,N_1815);
nor U2359 (N_2359,N_1981,N_1550);
and U2360 (N_2360,N_1723,N_1844);
nor U2361 (N_2361,N_1868,N_1906);
xnor U2362 (N_2362,N_1601,N_1660);
nand U2363 (N_2363,N_1956,N_1707);
xnor U2364 (N_2364,N_1517,N_1926);
nand U2365 (N_2365,N_1649,N_1505);
and U2366 (N_2366,N_1941,N_1501);
and U2367 (N_2367,N_1891,N_1940);
or U2368 (N_2368,N_1877,N_1864);
or U2369 (N_2369,N_1853,N_1607);
nand U2370 (N_2370,N_1845,N_1639);
and U2371 (N_2371,N_1997,N_1798);
nand U2372 (N_2372,N_1722,N_1609);
and U2373 (N_2373,N_1893,N_1920);
or U2374 (N_2374,N_1791,N_1735);
or U2375 (N_2375,N_1508,N_1657);
nor U2376 (N_2376,N_1537,N_1807);
nor U2377 (N_2377,N_1848,N_1828);
nand U2378 (N_2378,N_1805,N_1627);
and U2379 (N_2379,N_1586,N_1885);
or U2380 (N_2380,N_1927,N_1520);
xor U2381 (N_2381,N_1508,N_1827);
xnor U2382 (N_2382,N_1857,N_1504);
nand U2383 (N_2383,N_1822,N_1937);
or U2384 (N_2384,N_1818,N_1964);
and U2385 (N_2385,N_1608,N_1842);
xor U2386 (N_2386,N_1938,N_1851);
nand U2387 (N_2387,N_1961,N_1832);
nand U2388 (N_2388,N_1786,N_1715);
nor U2389 (N_2389,N_1832,N_1843);
nand U2390 (N_2390,N_1745,N_1959);
or U2391 (N_2391,N_1856,N_1621);
and U2392 (N_2392,N_1522,N_1912);
and U2393 (N_2393,N_1688,N_1824);
or U2394 (N_2394,N_1977,N_1667);
nand U2395 (N_2395,N_1600,N_1630);
nand U2396 (N_2396,N_1724,N_1744);
nor U2397 (N_2397,N_1946,N_1739);
and U2398 (N_2398,N_1680,N_1660);
xor U2399 (N_2399,N_1718,N_1569);
or U2400 (N_2400,N_1916,N_1720);
nand U2401 (N_2401,N_1546,N_1884);
nor U2402 (N_2402,N_1559,N_1578);
nand U2403 (N_2403,N_1826,N_1673);
and U2404 (N_2404,N_1579,N_1863);
or U2405 (N_2405,N_1716,N_1854);
and U2406 (N_2406,N_1614,N_1661);
or U2407 (N_2407,N_1992,N_1510);
nor U2408 (N_2408,N_1624,N_1655);
and U2409 (N_2409,N_1570,N_1894);
nor U2410 (N_2410,N_1990,N_1708);
nand U2411 (N_2411,N_1838,N_1706);
and U2412 (N_2412,N_1809,N_1506);
nand U2413 (N_2413,N_1707,N_1904);
or U2414 (N_2414,N_1693,N_1757);
and U2415 (N_2415,N_1728,N_1726);
nand U2416 (N_2416,N_1848,N_1586);
or U2417 (N_2417,N_1711,N_1827);
and U2418 (N_2418,N_1892,N_1516);
nor U2419 (N_2419,N_1885,N_1861);
or U2420 (N_2420,N_1778,N_1704);
nand U2421 (N_2421,N_1515,N_1672);
nor U2422 (N_2422,N_1552,N_1798);
nor U2423 (N_2423,N_1679,N_1962);
or U2424 (N_2424,N_1952,N_1761);
or U2425 (N_2425,N_1637,N_1650);
nor U2426 (N_2426,N_1793,N_1972);
nand U2427 (N_2427,N_1704,N_1598);
xor U2428 (N_2428,N_1714,N_1625);
and U2429 (N_2429,N_1512,N_1994);
or U2430 (N_2430,N_1895,N_1644);
nand U2431 (N_2431,N_1912,N_1634);
and U2432 (N_2432,N_1889,N_1503);
or U2433 (N_2433,N_1531,N_1564);
or U2434 (N_2434,N_1852,N_1749);
nand U2435 (N_2435,N_1845,N_1668);
nand U2436 (N_2436,N_1536,N_1601);
and U2437 (N_2437,N_1584,N_1553);
or U2438 (N_2438,N_1872,N_1889);
and U2439 (N_2439,N_1715,N_1537);
or U2440 (N_2440,N_1607,N_1680);
and U2441 (N_2441,N_1551,N_1734);
or U2442 (N_2442,N_1849,N_1577);
or U2443 (N_2443,N_1737,N_1734);
and U2444 (N_2444,N_1870,N_1951);
and U2445 (N_2445,N_1541,N_1594);
nor U2446 (N_2446,N_1621,N_1983);
nor U2447 (N_2447,N_1783,N_1722);
xor U2448 (N_2448,N_1879,N_1634);
nand U2449 (N_2449,N_1799,N_1854);
or U2450 (N_2450,N_1932,N_1694);
nand U2451 (N_2451,N_1509,N_1872);
nor U2452 (N_2452,N_1886,N_1600);
and U2453 (N_2453,N_1805,N_1634);
or U2454 (N_2454,N_1980,N_1708);
and U2455 (N_2455,N_1550,N_1697);
nand U2456 (N_2456,N_1549,N_1936);
or U2457 (N_2457,N_1725,N_1679);
and U2458 (N_2458,N_1700,N_1717);
and U2459 (N_2459,N_1893,N_1822);
nor U2460 (N_2460,N_1724,N_1807);
nand U2461 (N_2461,N_1818,N_1519);
nand U2462 (N_2462,N_1615,N_1539);
nand U2463 (N_2463,N_1643,N_1605);
nor U2464 (N_2464,N_1901,N_1953);
or U2465 (N_2465,N_1510,N_1623);
or U2466 (N_2466,N_1501,N_1657);
nand U2467 (N_2467,N_1655,N_1790);
and U2468 (N_2468,N_1638,N_1751);
and U2469 (N_2469,N_1828,N_1876);
and U2470 (N_2470,N_1968,N_1605);
nand U2471 (N_2471,N_1528,N_1510);
or U2472 (N_2472,N_1680,N_1608);
nor U2473 (N_2473,N_1954,N_1842);
nand U2474 (N_2474,N_1799,N_1679);
or U2475 (N_2475,N_1710,N_1786);
nand U2476 (N_2476,N_1796,N_1820);
nand U2477 (N_2477,N_1933,N_1685);
and U2478 (N_2478,N_1784,N_1550);
nor U2479 (N_2479,N_1847,N_1681);
nand U2480 (N_2480,N_1591,N_1516);
and U2481 (N_2481,N_1596,N_1734);
or U2482 (N_2482,N_1855,N_1507);
nand U2483 (N_2483,N_1697,N_1690);
nor U2484 (N_2484,N_1730,N_1698);
or U2485 (N_2485,N_1541,N_1592);
or U2486 (N_2486,N_1930,N_1864);
nor U2487 (N_2487,N_1810,N_1630);
or U2488 (N_2488,N_1955,N_1874);
nand U2489 (N_2489,N_1620,N_1523);
nand U2490 (N_2490,N_1919,N_1888);
xnor U2491 (N_2491,N_1793,N_1613);
nand U2492 (N_2492,N_1996,N_1575);
nor U2493 (N_2493,N_1913,N_1759);
nand U2494 (N_2494,N_1606,N_1737);
nor U2495 (N_2495,N_1886,N_1819);
or U2496 (N_2496,N_1746,N_1782);
or U2497 (N_2497,N_1753,N_1996);
nor U2498 (N_2498,N_1656,N_1775);
nor U2499 (N_2499,N_1877,N_1869);
nand U2500 (N_2500,N_2059,N_2005);
nand U2501 (N_2501,N_2485,N_2247);
nor U2502 (N_2502,N_2383,N_2011);
and U2503 (N_2503,N_2231,N_2331);
nor U2504 (N_2504,N_2474,N_2230);
xor U2505 (N_2505,N_2152,N_2174);
or U2506 (N_2506,N_2309,N_2394);
and U2507 (N_2507,N_2036,N_2143);
or U2508 (N_2508,N_2387,N_2255);
nand U2509 (N_2509,N_2377,N_2042);
nand U2510 (N_2510,N_2419,N_2115);
and U2511 (N_2511,N_2364,N_2168);
nand U2512 (N_2512,N_2139,N_2121);
xnor U2513 (N_2513,N_2234,N_2291);
and U2514 (N_2514,N_2102,N_2459);
nor U2515 (N_2515,N_2164,N_2223);
or U2516 (N_2516,N_2030,N_2211);
nand U2517 (N_2517,N_2285,N_2456);
nand U2518 (N_2518,N_2431,N_2018);
nand U2519 (N_2519,N_2055,N_2292);
nand U2520 (N_2520,N_2172,N_2490);
or U2521 (N_2521,N_2409,N_2111);
nand U2522 (N_2522,N_2410,N_2159);
nor U2523 (N_2523,N_2357,N_2279);
nor U2524 (N_2524,N_2250,N_2060);
nand U2525 (N_2525,N_2420,N_2026);
xnor U2526 (N_2526,N_2338,N_2393);
nand U2527 (N_2527,N_2244,N_2216);
nor U2528 (N_2528,N_2316,N_2296);
nand U2529 (N_2529,N_2155,N_2430);
nor U2530 (N_2530,N_2432,N_2233);
nor U2531 (N_2531,N_2403,N_2421);
nor U2532 (N_2532,N_2088,N_2012);
and U2533 (N_2533,N_2219,N_2069);
or U2534 (N_2534,N_2039,N_2087);
nand U2535 (N_2535,N_2356,N_2232);
or U2536 (N_2536,N_2192,N_2082);
and U2537 (N_2537,N_2312,N_2074);
or U2538 (N_2538,N_2463,N_2146);
and U2539 (N_2539,N_2161,N_2273);
and U2540 (N_2540,N_2217,N_2493);
nand U2541 (N_2541,N_2347,N_2045);
nor U2542 (N_2542,N_2204,N_2130);
or U2543 (N_2543,N_2259,N_2201);
nor U2544 (N_2544,N_2141,N_2458);
or U2545 (N_2545,N_2299,N_2272);
or U2546 (N_2546,N_2317,N_2099);
xor U2547 (N_2547,N_2149,N_2196);
or U2548 (N_2548,N_2344,N_2160);
or U2549 (N_2549,N_2235,N_2365);
and U2550 (N_2550,N_2491,N_2202);
nor U2551 (N_2551,N_2209,N_2107);
nor U2552 (N_2552,N_2256,N_2276);
nor U2553 (N_2553,N_2411,N_2423);
or U2554 (N_2554,N_2443,N_2437);
or U2555 (N_2555,N_2479,N_2402);
nand U2556 (N_2556,N_2305,N_2451);
nand U2557 (N_2557,N_2078,N_2123);
and U2558 (N_2558,N_2213,N_2212);
or U2559 (N_2559,N_2040,N_2448);
or U2560 (N_2560,N_2147,N_2390);
xor U2561 (N_2561,N_2095,N_2108);
or U2562 (N_2562,N_2298,N_2190);
nor U2563 (N_2563,N_2089,N_2466);
or U2564 (N_2564,N_2475,N_2484);
xor U2565 (N_2565,N_2348,N_2068);
nand U2566 (N_2566,N_2156,N_2416);
or U2567 (N_2567,N_2001,N_2341);
nand U2568 (N_2568,N_2206,N_2371);
nand U2569 (N_2569,N_2199,N_2311);
nand U2570 (N_2570,N_2313,N_2268);
and U2571 (N_2571,N_2062,N_2444);
nor U2572 (N_2572,N_2125,N_2414);
nand U2573 (N_2573,N_2142,N_2406);
nor U2574 (N_2574,N_2461,N_2304);
nor U2575 (N_2575,N_2081,N_2440);
or U2576 (N_2576,N_2265,N_2310);
nand U2577 (N_2577,N_2359,N_2385);
nand U2578 (N_2578,N_2085,N_2252);
nor U2579 (N_2579,N_2464,N_2072);
nor U2580 (N_2580,N_2200,N_2243);
nand U2581 (N_2581,N_2038,N_2119);
nor U2582 (N_2582,N_2096,N_2483);
nand U2583 (N_2583,N_2395,N_2236);
and U2584 (N_2584,N_2028,N_2024);
and U2585 (N_2585,N_2091,N_2127);
and U2586 (N_2586,N_2282,N_2425);
and U2587 (N_2587,N_2009,N_2242);
or U2588 (N_2588,N_2408,N_2381);
nor U2589 (N_2589,N_2225,N_2157);
xor U2590 (N_2590,N_2071,N_2436);
xor U2591 (N_2591,N_2048,N_2013);
nand U2592 (N_2592,N_2092,N_2194);
or U2593 (N_2593,N_2162,N_2433);
nand U2594 (N_2594,N_2375,N_2270);
nor U2595 (N_2595,N_2056,N_2495);
and U2596 (N_2596,N_2446,N_2195);
xnor U2597 (N_2597,N_2128,N_2413);
and U2598 (N_2598,N_2000,N_2277);
nand U2599 (N_2599,N_2379,N_2301);
xor U2600 (N_2600,N_2294,N_2037);
nor U2601 (N_2601,N_2333,N_2358);
nor U2602 (N_2602,N_2049,N_2083);
and U2603 (N_2603,N_2441,N_2284);
and U2604 (N_2604,N_2281,N_2260);
or U2605 (N_2605,N_2271,N_2468);
or U2606 (N_2606,N_2065,N_2266);
xor U2607 (N_2607,N_2224,N_2227);
nand U2608 (N_2608,N_2245,N_2480);
nor U2609 (N_2609,N_2166,N_2114);
and U2610 (N_2610,N_2469,N_2335);
nand U2611 (N_2611,N_2498,N_2171);
or U2612 (N_2612,N_2486,N_2424);
or U2613 (N_2613,N_2354,N_2120);
nand U2614 (N_2614,N_2417,N_2322);
or U2615 (N_2615,N_2315,N_2360);
or U2616 (N_2616,N_2006,N_2035);
and U2617 (N_2617,N_2499,N_2457);
nand U2618 (N_2618,N_2496,N_2138);
or U2619 (N_2619,N_2452,N_2189);
and U2620 (N_2620,N_2439,N_2080);
nand U2621 (N_2621,N_2004,N_2382);
and U2622 (N_2622,N_2366,N_2465);
nand U2623 (N_2623,N_2163,N_2497);
xor U2624 (N_2624,N_2349,N_2133);
xor U2625 (N_2625,N_2239,N_2057);
nand U2626 (N_2626,N_2346,N_2186);
nand U2627 (N_2627,N_2388,N_2391);
xnor U2628 (N_2628,N_2117,N_2257);
nor U2629 (N_2629,N_2422,N_2113);
or U2630 (N_2630,N_2492,N_2396);
and U2631 (N_2631,N_2207,N_2473);
nand U2632 (N_2632,N_2470,N_2210);
and U2633 (N_2633,N_2105,N_2428);
and U2634 (N_2634,N_2010,N_2263);
xor U2635 (N_2635,N_2150,N_2450);
nor U2636 (N_2636,N_2106,N_2022);
xor U2637 (N_2637,N_2077,N_2286);
or U2638 (N_2638,N_2218,N_2144);
nor U2639 (N_2639,N_2253,N_2453);
or U2640 (N_2640,N_2140,N_2280);
and U2641 (N_2641,N_2302,N_2215);
or U2642 (N_2642,N_2398,N_2368);
nor U2643 (N_2643,N_2399,N_2367);
nand U2644 (N_2644,N_2454,N_2021);
nand U2645 (N_2645,N_2400,N_2460);
or U2646 (N_2646,N_2203,N_2182);
or U2647 (N_2647,N_2476,N_2249);
nand U2648 (N_2648,N_2044,N_2169);
nor U2649 (N_2649,N_2261,N_2293);
and U2650 (N_2650,N_2027,N_2307);
nor U2651 (N_2651,N_2337,N_2240);
or U2652 (N_2652,N_2401,N_2447);
or U2653 (N_2653,N_2445,N_2122);
nand U2654 (N_2654,N_2325,N_2154);
and U2655 (N_2655,N_2179,N_2061);
and U2656 (N_2656,N_2334,N_2058);
nor U2657 (N_2657,N_2165,N_2041);
and U2658 (N_2658,N_2407,N_2370);
or U2659 (N_2659,N_2003,N_2369);
nor U2660 (N_2660,N_2258,N_2241);
xnor U2661 (N_2661,N_2124,N_2101);
nand U2662 (N_2662,N_2449,N_2007);
or U2663 (N_2663,N_2067,N_2129);
or U2664 (N_2664,N_2295,N_2073);
nand U2665 (N_2665,N_2326,N_2118);
or U2666 (N_2666,N_2328,N_2153);
or U2667 (N_2667,N_2220,N_2208);
or U2668 (N_2668,N_2148,N_2246);
and U2669 (N_2669,N_2084,N_2254);
nand U2670 (N_2670,N_2467,N_2314);
and U2671 (N_2671,N_2187,N_2051);
or U2672 (N_2672,N_2435,N_2462);
nor U2673 (N_2673,N_2086,N_2248);
nand U2674 (N_2674,N_2029,N_2306);
nor U2675 (N_2675,N_2177,N_2237);
or U2676 (N_2676,N_2361,N_2329);
nor U2677 (N_2677,N_2287,N_2050);
or U2678 (N_2678,N_2275,N_2472);
nand U2679 (N_2679,N_2471,N_2308);
or U2680 (N_2680,N_2031,N_2226);
or U2681 (N_2681,N_2418,N_2412);
nor U2682 (N_2682,N_2350,N_2415);
or U2683 (N_2683,N_2170,N_2053);
or U2684 (N_2684,N_2264,N_2158);
nand U2685 (N_2685,N_2070,N_2145);
and U2686 (N_2686,N_2289,N_2278);
nor U2687 (N_2687,N_2362,N_2318);
and U2688 (N_2688,N_2345,N_2290);
nor U2689 (N_2689,N_2340,N_2426);
or U2690 (N_2690,N_2336,N_2100);
xor U2691 (N_2691,N_2327,N_2376);
and U2692 (N_2692,N_2098,N_2109);
and U2693 (N_2693,N_2330,N_2181);
and U2694 (N_2694,N_2269,N_2112);
nor U2695 (N_2695,N_2324,N_2303);
or U2696 (N_2696,N_2488,N_2339);
or U2697 (N_2697,N_2052,N_2191);
nand U2698 (N_2698,N_2380,N_2262);
and U2699 (N_2699,N_2297,N_2300);
nand U2700 (N_2700,N_2442,N_2015);
xor U2701 (N_2701,N_2033,N_2283);
or U2702 (N_2702,N_2481,N_2188);
or U2703 (N_2703,N_2228,N_2017);
and U2704 (N_2704,N_2126,N_2288);
or U2705 (N_2705,N_2372,N_2034);
and U2706 (N_2706,N_2222,N_2176);
or U2707 (N_2707,N_2332,N_2032);
nor U2708 (N_2708,N_2093,N_2386);
nand U2709 (N_2709,N_2355,N_2205);
xnor U2710 (N_2710,N_2405,N_2131);
nand U2711 (N_2711,N_2135,N_2097);
or U2712 (N_2712,N_2198,N_2267);
and U2713 (N_2713,N_2343,N_2494);
and U2714 (N_2714,N_2016,N_2487);
nor U2715 (N_2715,N_2229,N_2184);
nand U2716 (N_2716,N_2178,N_2238);
nor U2717 (N_2717,N_2116,N_2183);
and U2718 (N_2718,N_2353,N_2274);
and U2719 (N_2719,N_2389,N_2342);
and U2720 (N_2720,N_2478,N_2455);
or U2721 (N_2721,N_2134,N_2193);
or U2722 (N_2722,N_2063,N_2075);
and U2723 (N_2723,N_2167,N_2373);
nor U2724 (N_2724,N_2429,N_2173);
nand U2725 (N_2725,N_2221,N_2046);
nor U2726 (N_2726,N_2094,N_2137);
nand U2727 (N_2727,N_2090,N_2019);
or U2728 (N_2728,N_2008,N_2482);
nor U2729 (N_2729,N_2066,N_2002);
or U2730 (N_2730,N_2320,N_2438);
or U2731 (N_2731,N_2047,N_2014);
nand U2732 (N_2732,N_2104,N_2180);
nand U2733 (N_2733,N_2103,N_2374);
and U2734 (N_2734,N_2434,N_2185);
or U2735 (N_2735,N_2378,N_2392);
nand U2736 (N_2736,N_2025,N_2064);
or U2737 (N_2737,N_2427,N_2323);
nand U2738 (N_2738,N_2023,N_2020);
or U2739 (N_2739,N_2110,N_2214);
or U2740 (N_2740,N_2397,N_2352);
nand U2741 (N_2741,N_2404,N_2321);
xor U2742 (N_2742,N_2132,N_2351);
or U2743 (N_2743,N_2054,N_2251);
nor U2744 (N_2744,N_2175,N_2079);
nor U2745 (N_2745,N_2076,N_2151);
or U2746 (N_2746,N_2384,N_2363);
or U2747 (N_2747,N_2197,N_2489);
and U2748 (N_2748,N_2136,N_2477);
or U2749 (N_2749,N_2319,N_2043);
xnor U2750 (N_2750,N_2031,N_2007);
or U2751 (N_2751,N_2124,N_2293);
and U2752 (N_2752,N_2070,N_2139);
or U2753 (N_2753,N_2012,N_2289);
xnor U2754 (N_2754,N_2038,N_2021);
and U2755 (N_2755,N_2495,N_2182);
nand U2756 (N_2756,N_2273,N_2280);
nand U2757 (N_2757,N_2009,N_2063);
xor U2758 (N_2758,N_2363,N_2200);
nor U2759 (N_2759,N_2227,N_2196);
nor U2760 (N_2760,N_2233,N_2262);
nand U2761 (N_2761,N_2040,N_2014);
and U2762 (N_2762,N_2249,N_2430);
nor U2763 (N_2763,N_2137,N_2215);
or U2764 (N_2764,N_2005,N_2440);
and U2765 (N_2765,N_2213,N_2478);
or U2766 (N_2766,N_2018,N_2082);
and U2767 (N_2767,N_2235,N_2383);
xor U2768 (N_2768,N_2459,N_2464);
or U2769 (N_2769,N_2057,N_2041);
and U2770 (N_2770,N_2411,N_2206);
nand U2771 (N_2771,N_2292,N_2404);
xor U2772 (N_2772,N_2155,N_2340);
and U2773 (N_2773,N_2001,N_2316);
or U2774 (N_2774,N_2098,N_2447);
and U2775 (N_2775,N_2076,N_2484);
and U2776 (N_2776,N_2282,N_2102);
and U2777 (N_2777,N_2124,N_2490);
or U2778 (N_2778,N_2378,N_2341);
nor U2779 (N_2779,N_2311,N_2386);
nand U2780 (N_2780,N_2175,N_2200);
and U2781 (N_2781,N_2410,N_2241);
xor U2782 (N_2782,N_2424,N_2092);
nand U2783 (N_2783,N_2242,N_2005);
and U2784 (N_2784,N_2126,N_2108);
nand U2785 (N_2785,N_2105,N_2071);
or U2786 (N_2786,N_2328,N_2255);
and U2787 (N_2787,N_2499,N_2420);
or U2788 (N_2788,N_2173,N_2433);
nor U2789 (N_2789,N_2304,N_2336);
nand U2790 (N_2790,N_2196,N_2374);
nand U2791 (N_2791,N_2484,N_2101);
nor U2792 (N_2792,N_2285,N_2126);
xnor U2793 (N_2793,N_2273,N_2267);
nor U2794 (N_2794,N_2256,N_2477);
or U2795 (N_2795,N_2443,N_2380);
or U2796 (N_2796,N_2052,N_2226);
or U2797 (N_2797,N_2161,N_2057);
nand U2798 (N_2798,N_2359,N_2084);
or U2799 (N_2799,N_2325,N_2375);
or U2800 (N_2800,N_2045,N_2158);
or U2801 (N_2801,N_2010,N_2145);
or U2802 (N_2802,N_2047,N_2493);
nor U2803 (N_2803,N_2139,N_2476);
and U2804 (N_2804,N_2259,N_2234);
nand U2805 (N_2805,N_2218,N_2107);
nand U2806 (N_2806,N_2348,N_2142);
nor U2807 (N_2807,N_2114,N_2426);
nand U2808 (N_2808,N_2111,N_2269);
nor U2809 (N_2809,N_2110,N_2220);
or U2810 (N_2810,N_2288,N_2263);
nor U2811 (N_2811,N_2248,N_2048);
nand U2812 (N_2812,N_2141,N_2293);
nand U2813 (N_2813,N_2362,N_2377);
and U2814 (N_2814,N_2339,N_2491);
or U2815 (N_2815,N_2023,N_2145);
nor U2816 (N_2816,N_2060,N_2297);
or U2817 (N_2817,N_2112,N_2470);
or U2818 (N_2818,N_2474,N_2259);
nand U2819 (N_2819,N_2364,N_2259);
nand U2820 (N_2820,N_2028,N_2265);
and U2821 (N_2821,N_2107,N_2106);
nor U2822 (N_2822,N_2074,N_2226);
and U2823 (N_2823,N_2358,N_2350);
and U2824 (N_2824,N_2476,N_2090);
xnor U2825 (N_2825,N_2394,N_2079);
and U2826 (N_2826,N_2313,N_2000);
nand U2827 (N_2827,N_2207,N_2391);
and U2828 (N_2828,N_2410,N_2374);
nand U2829 (N_2829,N_2243,N_2146);
and U2830 (N_2830,N_2442,N_2204);
nand U2831 (N_2831,N_2175,N_2351);
or U2832 (N_2832,N_2259,N_2379);
nor U2833 (N_2833,N_2474,N_2264);
nand U2834 (N_2834,N_2193,N_2168);
or U2835 (N_2835,N_2118,N_2383);
nor U2836 (N_2836,N_2235,N_2310);
xor U2837 (N_2837,N_2395,N_2029);
nand U2838 (N_2838,N_2125,N_2473);
nand U2839 (N_2839,N_2154,N_2000);
nand U2840 (N_2840,N_2378,N_2139);
nor U2841 (N_2841,N_2311,N_2383);
and U2842 (N_2842,N_2170,N_2255);
or U2843 (N_2843,N_2115,N_2157);
nand U2844 (N_2844,N_2001,N_2013);
nand U2845 (N_2845,N_2226,N_2097);
and U2846 (N_2846,N_2492,N_2082);
nor U2847 (N_2847,N_2026,N_2193);
and U2848 (N_2848,N_2201,N_2293);
or U2849 (N_2849,N_2228,N_2332);
nor U2850 (N_2850,N_2467,N_2335);
nand U2851 (N_2851,N_2270,N_2480);
nor U2852 (N_2852,N_2472,N_2484);
and U2853 (N_2853,N_2404,N_2374);
nand U2854 (N_2854,N_2073,N_2003);
or U2855 (N_2855,N_2464,N_2011);
xor U2856 (N_2856,N_2462,N_2031);
and U2857 (N_2857,N_2353,N_2002);
nand U2858 (N_2858,N_2184,N_2329);
or U2859 (N_2859,N_2378,N_2049);
xor U2860 (N_2860,N_2156,N_2355);
and U2861 (N_2861,N_2190,N_2433);
xnor U2862 (N_2862,N_2300,N_2072);
or U2863 (N_2863,N_2259,N_2151);
or U2864 (N_2864,N_2182,N_2325);
nand U2865 (N_2865,N_2316,N_2162);
or U2866 (N_2866,N_2353,N_2409);
nand U2867 (N_2867,N_2359,N_2146);
or U2868 (N_2868,N_2349,N_2461);
and U2869 (N_2869,N_2212,N_2409);
nor U2870 (N_2870,N_2129,N_2463);
nand U2871 (N_2871,N_2020,N_2175);
nor U2872 (N_2872,N_2430,N_2055);
xor U2873 (N_2873,N_2450,N_2308);
or U2874 (N_2874,N_2141,N_2038);
and U2875 (N_2875,N_2193,N_2013);
nand U2876 (N_2876,N_2211,N_2249);
nand U2877 (N_2877,N_2032,N_2230);
and U2878 (N_2878,N_2034,N_2124);
nor U2879 (N_2879,N_2410,N_2455);
or U2880 (N_2880,N_2307,N_2280);
and U2881 (N_2881,N_2033,N_2022);
and U2882 (N_2882,N_2082,N_2357);
or U2883 (N_2883,N_2497,N_2467);
nand U2884 (N_2884,N_2496,N_2393);
nand U2885 (N_2885,N_2281,N_2371);
nand U2886 (N_2886,N_2445,N_2106);
and U2887 (N_2887,N_2032,N_2167);
xnor U2888 (N_2888,N_2419,N_2281);
xnor U2889 (N_2889,N_2378,N_2275);
and U2890 (N_2890,N_2100,N_2272);
or U2891 (N_2891,N_2333,N_2195);
or U2892 (N_2892,N_2013,N_2386);
nand U2893 (N_2893,N_2166,N_2182);
or U2894 (N_2894,N_2363,N_2007);
nor U2895 (N_2895,N_2178,N_2098);
nand U2896 (N_2896,N_2075,N_2313);
and U2897 (N_2897,N_2012,N_2025);
and U2898 (N_2898,N_2298,N_2031);
nand U2899 (N_2899,N_2130,N_2299);
nor U2900 (N_2900,N_2212,N_2252);
or U2901 (N_2901,N_2419,N_2239);
and U2902 (N_2902,N_2481,N_2205);
nor U2903 (N_2903,N_2373,N_2182);
nor U2904 (N_2904,N_2439,N_2486);
nand U2905 (N_2905,N_2179,N_2439);
and U2906 (N_2906,N_2327,N_2222);
nor U2907 (N_2907,N_2448,N_2490);
nand U2908 (N_2908,N_2323,N_2345);
nand U2909 (N_2909,N_2251,N_2204);
nand U2910 (N_2910,N_2021,N_2190);
and U2911 (N_2911,N_2399,N_2363);
or U2912 (N_2912,N_2131,N_2426);
and U2913 (N_2913,N_2081,N_2406);
and U2914 (N_2914,N_2203,N_2485);
or U2915 (N_2915,N_2405,N_2214);
or U2916 (N_2916,N_2308,N_2008);
nor U2917 (N_2917,N_2009,N_2466);
nand U2918 (N_2918,N_2025,N_2315);
nand U2919 (N_2919,N_2146,N_2158);
or U2920 (N_2920,N_2092,N_2160);
nor U2921 (N_2921,N_2073,N_2145);
xnor U2922 (N_2922,N_2012,N_2208);
or U2923 (N_2923,N_2135,N_2037);
xor U2924 (N_2924,N_2176,N_2021);
or U2925 (N_2925,N_2437,N_2189);
or U2926 (N_2926,N_2156,N_2415);
xor U2927 (N_2927,N_2328,N_2232);
or U2928 (N_2928,N_2034,N_2256);
and U2929 (N_2929,N_2095,N_2169);
nor U2930 (N_2930,N_2388,N_2397);
nand U2931 (N_2931,N_2096,N_2344);
and U2932 (N_2932,N_2185,N_2192);
nor U2933 (N_2933,N_2439,N_2079);
and U2934 (N_2934,N_2183,N_2266);
nand U2935 (N_2935,N_2278,N_2426);
or U2936 (N_2936,N_2476,N_2224);
or U2937 (N_2937,N_2363,N_2184);
or U2938 (N_2938,N_2480,N_2412);
nor U2939 (N_2939,N_2093,N_2229);
nor U2940 (N_2940,N_2067,N_2089);
nand U2941 (N_2941,N_2038,N_2363);
nand U2942 (N_2942,N_2278,N_2001);
and U2943 (N_2943,N_2482,N_2362);
nand U2944 (N_2944,N_2015,N_2036);
nand U2945 (N_2945,N_2103,N_2428);
nor U2946 (N_2946,N_2260,N_2136);
or U2947 (N_2947,N_2260,N_2231);
nand U2948 (N_2948,N_2055,N_2261);
or U2949 (N_2949,N_2054,N_2319);
or U2950 (N_2950,N_2342,N_2058);
xnor U2951 (N_2951,N_2277,N_2496);
and U2952 (N_2952,N_2288,N_2069);
and U2953 (N_2953,N_2449,N_2298);
nor U2954 (N_2954,N_2426,N_2241);
and U2955 (N_2955,N_2450,N_2013);
or U2956 (N_2956,N_2414,N_2362);
xnor U2957 (N_2957,N_2263,N_2334);
or U2958 (N_2958,N_2045,N_2130);
nand U2959 (N_2959,N_2145,N_2071);
xor U2960 (N_2960,N_2303,N_2459);
nand U2961 (N_2961,N_2208,N_2249);
or U2962 (N_2962,N_2266,N_2399);
or U2963 (N_2963,N_2402,N_2162);
and U2964 (N_2964,N_2407,N_2251);
xor U2965 (N_2965,N_2298,N_2324);
nor U2966 (N_2966,N_2402,N_2335);
and U2967 (N_2967,N_2267,N_2328);
nand U2968 (N_2968,N_2422,N_2362);
or U2969 (N_2969,N_2319,N_2092);
xnor U2970 (N_2970,N_2473,N_2161);
nand U2971 (N_2971,N_2042,N_2037);
and U2972 (N_2972,N_2118,N_2224);
nor U2973 (N_2973,N_2077,N_2427);
or U2974 (N_2974,N_2015,N_2016);
xor U2975 (N_2975,N_2122,N_2135);
nor U2976 (N_2976,N_2470,N_2339);
nand U2977 (N_2977,N_2444,N_2026);
nor U2978 (N_2978,N_2173,N_2382);
and U2979 (N_2979,N_2269,N_2299);
and U2980 (N_2980,N_2090,N_2279);
and U2981 (N_2981,N_2334,N_2371);
and U2982 (N_2982,N_2322,N_2111);
nor U2983 (N_2983,N_2052,N_2324);
and U2984 (N_2984,N_2001,N_2138);
and U2985 (N_2985,N_2123,N_2160);
and U2986 (N_2986,N_2052,N_2308);
and U2987 (N_2987,N_2232,N_2485);
or U2988 (N_2988,N_2345,N_2384);
nor U2989 (N_2989,N_2220,N_2250);
or U2990 (N_2990,N_2042,N_2263);
nor U2991 (N_2991,N_2368,N_2204);
or U2992 (N_2992,N_2449,N_2253);
or U2993 (N_2993,N_2487,N_2461);
nand U2994 (N_2994,N_2338,N_2359);
or U2995 (N_2995,N_2396,N_2266);
nand U2996 (N_2996,N_2069,N_2157);
nand U2997 (N_2997,N_2157,N_2260);
and U2998 (N_2998,N_2486,N_2303);
nand U2999 (N_2999,N_2297,N_2193);
nand U3000 (N_3000,N_2705,N_2620);
xor U3001 (N_3001,N_2501,N_2921);
nor U3002 (N_3002,N_2823,N_2808);
and U3003 (N_3003,N_2630,N_2642);
and U3004 (N_3004,N_2811,N_2662);
and U3005 (N_3005,N_2694,N_2856);
or U3006 (N_3006,N_2843,N_2989);
and U3007 (N_3007,N_2699,N_2708);
and U3008 (N_3008,N_2883,N_2554);
and U3009 (N_3009,N_2924,N_2665);
or U3010 (N_3010,N_2608,N_2936);
nor U3011 (N_3011,N_2701,N_2769);
and U3012 (N_3012,N_2686,N_2561);
xnor U3013 (N_3013,N_2857,N_2899);
nand U3014 (N_3014,N_2802,N_2616);
xnor U3015 (N_3015,N_2793,N_2969);
and U3016 (N_3016,N_2589,N_2884);
or U3017 (N_3017,N_2707,N_2555);
and U3018 (N_3018,N_2632,N_2988);
or U3019 (N_3019,N_2733,N_2613);
or U3020 (N_3020,N_2865,N_2978);
or U3021 (N_3021,N_2687,N_2901);
nand U3022 (N_3022,N_2556,N_2749);
or U3023 (N_3023,N_2890,N_2631);
nor U3024 (N_3024,N_2621,N_2680);
or U3025 (N_3025,N_2704,N_2675);
nor U3026 (N_3026,N_2731,N_2787);
nand U3027 (N_3027,N_2940,N_2738);
or U3028 (N_3028,N_2594,N_2909);
nor U3029 (N_3029,N_2752,N_2540);
nand U3030 (N_3030,N_2892,N_2805);
nand U3031 (N_3031,N_2814,N_2848);
nand U3032 (N_3032,N_2548,N_2502);
nand U3033 (N_3033,N_2746,N_2963);
nor U3034 (N_3034,N_2618,N_2813);
and U3035 (N_3035,N_2654,N_2640);
nor U3036 (N_3036,N_2624,N_2755);
and U3037 (N_3037,N_2717,N_2550);
and U3038 (N_3038,N_2923,N_2954);
nand U3039 (N_3039,N_2649,N_2816);
xnor U3040 (N_3040,N_2774,N_2584);
or U3041 (N_3041,N_2847,N_2653);
and U3042 (N_3042,N_2551,N_2801);
or U3043 (N_3043,N_2879,N_2671);
nand U3044 (N_3044,N_2937,N_2505);
nor U3045 (N_3045,N_2919,N_2971);
and U3046 (N_3046,N_2754,N_2711);
and U3047 (N_3047,N_2809,N_2543);
and U3048 (N_3048,N_2734,N_2677);
and U3049 (N_3049,N_2944,N_2688);
nand U3050 (N_3050,N_2840,N_2775);
xor U3051 (N_3051,N_2852,N_2743);
and U3052 (N_3052,N_2633,N_2927);
nand U3053 (N_3053,N_2986,N_2600);
nand U3054 (N_3054,N_2881,N_2693);
nand U3055 (N_3055,N_2770,N_2957);
nor U3056 (N_3056,N_2850,N_2966);
nand U3057 (N_3057,N_2634,N_2602);
or U3058 (N_3058,N_2635,N_2724);
nor U3059 (N_3059,N_2636,N_2612);
xor U3060 (N_3060,N_2532,N_2508);
and U3061 (N_3061,N_2511,N_2663);
or U3062 (N_3062,N_2762,N_2827);
nand U3063 (N_3063,N_2539,N_2896);
and U3064 (N_3064,N_2519,N_2860);
nand U3065 (N_3065,N_2619,N_2975);
and U3066 (N_3066,N_2776,N_2789);
or U3067 (N_3067,N_2666,N_2715);
nor U3068 (N_3068,N_2629,N_2567);
or U3069 (N_3069,N_2737,N_2898);
nor U3070 (N_3070,N_2744,N_2646);
and U3071 (N_3071,N_2572,N_2930);
and U3072 (N_3072,N_2784,N_2991);
xor U3073 (N_3073,N_2709,N_2796);
nor U3074 (N_3074,N_2875,N_2753);
xnor U3075 (N_3075,N_2974,N_2534);
and U3076 (N_3076,N_2798,N_2582);
xnor U3077 (N_3077,N_2997,N_2985);
or U3078 (N_3078,N_2571,N_2580);
nor U3079 (N_3079,N_2895,N_2723);
nor U3080 (N_3080,N_2617,N_2506);
nor U3081 (N_3081,N_2660,N_2751);
nor U3082 (N_3082,N_2569,N_2657);
and U3083 (N_3083,N_2515,N_2943);
nor U3084 (N_3084,N_2728,N_2845);
and U3085 (N_3085,N_2696,N_2512);
nor U3086 (N_3086,N_2670,N_2570);
and U3087 (N_3087,N_2907,N_2651);
and U3088 (N_3088,N_2968,N_2729);
nor U3089 (N_3089,N_2503,N_2839);
nor U3090 (N_3090,N_2819,N_2983);
nor U3091 (N_3091,N_2524,N_2804);
xor U3092 (N_3092,N_2607,N_2626);
nand U3093 (N_3093,N_2535,N_2574);
xnor U3094 (N_3094,N_2588,N_2960);
and U3095 (N_3095,N_2664,N_2722);
xnor U3096 (N_3096,N_2807,N_2911);
nor U3097 (N_3097,N_2702,N_2851);
nor U3098 (N_3098,N_2598,N_2609);
and U3099 (N_3099,N_2586,N_2868);
and U3100 (N_3100,N_2961,N_2538);
nor U3101 (N_3101,N_2964,N_2672);
and U3102 (N_3102,N_2806,N_2623);
xor U3103 (N_3103,N_2523,N_2591);
nor U3104 (N_3104,N_2973,N_2577);
nor U3105 (N_3105,N_2541,N_2563);
or U3106 (N_3106,N_2956,N_2810);
nor U3107 (N_3107,N_2815,N_2922);
xor U3108 (N_3108,N_2976,N_2597);
xnor U3109 (N_3109,N_2903,N_2934);
or U3110 (N_3110,N_2627,N_2500);
nor U3111 (N_3111,N_2926,N_2880);
and U3112 (N_3112,N_2557,N_2844);
xnor U3113 (N_3113,N_2996,N_2596);
nor U3114 (N_3114,N_2849,N_2732);
or U3115 (N_3115,N_2977,N_2526);
nor U3116 (N_3116,N_2866,N_2656);
and U3117 (N_3117,N_2716,N_2763);
and U3118 (N_3118,N_2610,N_2833);
or U3119 (N_3119,N_2533,N_2575);
nand U3120 (N_3120,N_2887,N_2999);
or U3121 (N_3121,N_2862,N_2949);
nor U3122 (N_3122,N_2611,N_2683);
nand U3123 (N_3123,N_2894,N_2792);
nand U3124 (N_3124,N_2908,N_2703);
nor U3125 (N_3125,N_2528,N_2652);
nor U3126 (N_3126,N_2928,N_2948);
nand U3127 (N_3127,N_2982,N_2786);
xor U3128 (N_3128,N_2552,N_2527);
or U3129 (N_3129,N_2993,N_2720);
or U3130 (N_3130,N_2842,N_2767);
nand U3131 (N_3131,N_2760,N_2546);
nand U3132 (N_3132,N_2648,N_2782);
nor U3133 (N_3133,N_2891,N_2537);
or U3134 (N_3134,N_2521,N_2593);
nand U3135 (N_3135,N_2525,N_2689);
or U3136 (N_3136,N_2685,N_2727);
nor U3137 (N_3137,N_2622,N_2573);
or U3138 (N_3138,N_2545,N_2773);
or U3139 (N_3139,N_2859,N_2544);
and U3140 (N_3140,N_2529,N_2886);
nor U3141 (N_3141,N_2872,N_2513);
xor U3142 (N_3142,N_2914,N_2951);
or U3143 (N_3143,N_2658,N_2765);
or U3144 (N_3144,N_2564,N_2542);
nand U3145 (N_3145,N_2910,N_2669);
or U3146 (N_3146,N_2935,N_2992);
and U3147 (N_3147,N_2504,N_2674);
or U3148 (N_3148,N_2742,N_2710);
nand U3149 (N_3149,N_2931,N_2592);
xnor U3150 (N_3150,N_2771,N_2583);
nand U3151 (N_3151,N_2897,N_2825);
nand U3152 (N_3152,N_2870,N_2605);
nor U3153 (N_3153,N_2599,N_2863);
nand U3154 (N_3154,N_2867,N_2614);
nor U3155 (N_3155,N_2695,N_2873);
and U3156 (N_3156,N_2604,N_2691);
xor U3157 (N_3157,N_2920,N_2871);
and U3158 (N_3158,N_2861,N_2576);
nand U3159 (N_3159,N_2668,N_2667);
nor U3160 (N_3160,N_2950,N_2522);
or U3161 (N_3161,N_2877,N_2779);
nand U3162 (N_3162,N_2566,N_2579);
nor U3163 (N_3163,N_2967,N_2706);
nand U3164 (N_3164,N_2509,N_2641);
nor U3165 (N_3165,N_2970,N_2780);
and U3166 (N_3166,N_2718,N_2628);
nand U3167 (N_3167,N_2719,N_2778);
nand U3168 (N_3168,N_2739,N_2854);
nor U3169 (N_3169,N_2955,N_2747);
or U3170 (N_3170,N_2888,N_2925);
or U3171 (N_3171,N_2748,N_2531);
or U3172 (N_3172,N_2998,N_2714);
nand U3173 (N_3173,N_2741,N_2726);
nand U3174 (N_3174,N_2637,N_2692);
and U3175 (N_3175,N_2581,N_2824);
nand U3176 (N_3176,N_2536,N_2794);
and U3177 (N_3177,N_2939,N_2791);
nand U3178 (N_3178,N_2812,N_2834);
and U3179 (N_3179,N_2800,N_2979);
or U3180 (N_3180,N_2638,N_2797);
nor U3181 (N_3181,N_2777,N_2684);
or U3182 (N_3182,N_2725,N_2981);
or U3183 (N_3183,N_2595,N_2952);
or U3184 (N_3184,N_2846,N_2915);
or U3185 (N_3185,N_2517,N_2962);
and U3186 (N_3186,N_2995,N_2678);
nand U3187 (N_3187,N_2945,N_2822);
nor U3188 (N_3188,N_2874,N_2905);
nand U3189 (N_3189,N_2958,N_2980);
nor U3190 (N_3190,N_2878,N_2549);
and U3191 (N_3191,N_2818,N_2757);
and U3192 (N_3192,N_2510,N_2941);
or U3193 (N_3193,N_2547,N_2606);
nor U3194 (N_3194,N_2698,N_2601);
nand U3195 (N_3195,N_2946,N_2768);
or U3196 (N_3196,N_2838,N_2918);
nor U3197 (N_3197,N_2644,N_2953);
or U3198 (N_3198,N_2697,N_2837);
nor U3199 (N_3199,N_2929,N_2507);
or U3200 (N_3200,N_2565,N_2713);
xnor U3201 (N_3201,N_2984,N_2916);
and U3202 (N_3202,N_2766,N_2917);
xor U3203 (N_3203,N_2906,N_2959);
and U3204 (N_3204,N_2817,N_2730);
or U3205 (N_3205,N_2876,N_2785);
or U3206 (N_3206,N_2942,N_2759);
nand U3207 (N_3207,N_2869,N_2700);
xnor U3208 (N_3208,N_2965,N_2756);
or U3209 (N_3209,N_2758,N_2832);
and U3210 (N_3210,N_2795,N_2821);
nor U3211 (N_3211,N_2740,N_2885);
nor U3212 (N_3212,N_2639,N_2994);
and U3213 (N_3213,N_2650,N_2659);
nor U3214 (N_3214,N_2553,N_2820);
nand U3215 (N_3215,N_2585,N_2900);
or U3216 (N_3216,N_2882,N_2745);
nand U3217 (N_3217,N_2790,N_2655);
nand U3218 (N_3218,N_2625,N_2736);
or U3219 (N_3219,N_2735,N_2645);
nand U3220 (N_3220,N_2712,N_2841);
or U3221 (N_3221,N_2562,N_2750);
and U3222 (N_3222,N_2568,N_2858);
or U3223 (N_3223,N_2912,N_2514);
xor U3224 (N_3224,N_2830,N_2615);
nor U3225 (N_3225,N_2853,N_2772);
and U3226 (N_3226,N_2836,N_2972);
nand U3227 (N_3227,N_2690,N_2520);
or U3228 (N_3228,N_2893,N_2803);
nor U3229 (N_3229,N_2516,N_2987);
or U3230 (N_3230,N_2682,N_2558);
xnor U3231 (N_3231,N_2643,N_2559);
or U3232 (N_3232,N_2933,N_2938);
or U3233 (N_3233,N_2902,N_2947);
and U3234 (N_3234,N_2826,N_2799);
and U3235 (N_3235,N_2788,N_2855);
and U3236 (N_3236,N_2530,N_2764);
nand U3237 (N_3237,N_2990,N_2676);
and U3238 (N_3238,N_2647,N_2889);
or U3239 (N_3239,N_2679,N_2761);
nand U3240 (N_3240,N_2828,N_2518);
or U3241 (N_3241,N_2673,N_2603);
nor U3242 (N_3242,N_2587,N_2829);
nand U3243 (N_3243,N_2681,N_2560);
nor U3244 (N_3244,N_2932,N_2831);
nand U3245 (N_3245,N_2578,N_2783);
nor U3246 (N_3246,N_2721,N_2835);
nand U3247 (N_3247,N_2781,N_2904);
or U3248 (N_3248,N_2913,N_2590);
nor U3249 (N_3249,N_2864,N_2661);
nand U3250 (N_3250,N_2666,N_2855);
and U3251 (N_3251,N_2578,N_2987);
nor U3252 (N_3252,N_2937,N_2646);
or U3253 (N_3253,N_2942,N_2717);
xnor U3254 (N_3254,N_2541,N_2704);
or U3255 (N_3255,N_2942,N_2965);
nand U3256 (N_3256,N_2651,N_2894);
and U3257 (N_3257,N_2571,N_2733);
nor U3258 (N_3258,N_2697,N_2787);
or U3259 (N_3259,N_2942,N_2730);
or U3260 (N_3260,N_2996,N_2983);
nand U3261 (N_3261,N_2660,N_2803);
nand U3262 (N_3262,N_2844,N_2556);
nand U3263 (N_3263,N_2650,N_2522);
nor U3264 (N_3264,N_2970,N_2935);
or U3265 (N_3265,N_2989,N_2561);
or U3266 (N_3266,N_2638,N_2555);
xor U3267 (N_3267,N_2886,N_2965);
nand U3268 (N_3268,N_2773,N_2711);
and U3269 (N_3269,N_2700,N_2800);
nand U3270 (N_3270,N_2676,N_2516);
or U3271 (N_3271,N_2903,N_2841);
or U3272 (N_3272,N_2993,N_2930);
nor U3273 (N_3273,N_2626,N_2690);
or U3274 (N_3274,N_2938,N_2737);
or U3275 (N_3275,N_2804,N_2880);
nor U3276 (N_3276,N_2701,N_2502);
nand U3277 (N_3277,N_2672,N_2601);
xnor U3278 (N_3278,N_2585,N_2609);
nor U3279 (N_3279,N_2988,N_2647);
or U3280 (N_3280,N_2819,N_2746);
nor U3281 (N_3281,N_2542,N_2904);
nor U3282 (N_3282,N_2832,N_2987);
nor U3283 (N_3283,N_2666,N_2507);
nand U3284 (N_3284,N_2729,N_2590);
and U3285 (N_3285,N_2548,N_2667);
xnor U3286 (N_3286,N_2881,N_2721);
and U3287 (N_3287,N_2658,N_2551);
and U3288 (N_3288,N_2786,N_2632);
or U3289 (N_3289,N_2921,N_2519);
nor U3290 (N_3290,N_2758,N_2650);
or U3291 (N_3291,N_2532,N_2945);
nor U3292 (N_3292,N_2673,N_2648);
nor U3293 (N_3293,N_2921,N_2626);
nor U3294 (N_3294,N_2786,N_2767);
nand U3295 (N_3295,N_2562,N_2860);
and U3296 (N_3296,N_2590,N_2851);
nand U3297 (N_3297,N_2966,N_2924);
xnor U3298 (N_3298,N_2819,N_2948);
xnor U3299 (N_3299,N_2829,N_2763);
nor U3300 (N_3300,N_2845,N_2843);
and U3301 (N_3301,N_2991,N_2546);
and U3302 (N_3302,N_2873,N_2646);
xnor U3303 (N_3303,N_2686,N_2972);
and U3304 (N_3304,N_2789,N_2558);
nand U3305 (N_3305,N_2596,N_2553);
nand U3306 (N_3306,N_2682,N_2566);
or U3307 (N_3307,N_2651,N_2963);
or U3308 (N_3308,N_2529,N_2513);
nor U3309 (N_3309,N_2967,N_2745);
or U3310 (N_3310,N_2849,N_2799);
nor U3311 (N_3311,N_2696,N_2599);
or U3312 (N_3312,N_2793,N_2994);
nand U3313 (N_3313,N_2509,N_2664);
or U3314 (N_3314,N_2601,N_2793);
nor U3315 (N_3315,N_2921,N_2974);
nor U3316 (N_3316,N_2685,N_2572);
or U3317 (N_3317,N_2893,N_2620);
nor U3318 (N_3318,N_2758,N_2655);
or U3319 (N_3319,N_2717,N_2962);
or U3320 (N_3320,N_2646,N_2644);
or U3321 (N_3321,N_2796,N_2961);
nor U3322 (N_3322,N_2953,N_2578);
nor U3323 (N_3323,N_2776,N_2931);
or U3324 (N_3324,N_2995,N_2599);
and U3325 (N_3325,N_2827,N_2765);
and U3326 (N_3326,N_2849,N_2991);
nand U3327 (N_3327,N_2665,N_2974);
and U3328 (N_3328,N_2758,N_2678);
xnor U3329 (N_3329,N_2792,N_2948);
or U3330 (N_3330,N_2650,N_2623);
and U3331 (N_3331,N_2520,N_2607);
or U3332 (N_3332,N_2910,N_2698);
nor U3333 (N_3333,N_2778,N_2968);
nand U3334 (N_3334,N_2778,N_2980);
nor U3335 (N_3335,N_2726,N_2949);
nand U3336 (N_3336,N_2572,N_2618);
nor U3337 (N_3337,N_2731,N_2907);
xnor U3338 (N_3338,N_2762,N_2773);
nor U3339 (N_3339,N_2689,N_2644);
and U3340 (N_3340,N_2900,N_2930);
xor U3341 (N_3341,N_2958,N_2928);
nor U3342 (N_3342,N_2595,N_2703);
xnor U3343 (N_3343,N_2910,N_2957);
nor U3344 (N_3344,N_2735,N_2517);
and U3345 (N_3345,N_2726,N_2844);
and U3346 (N_3346,N_2640,N_2562);
nand U3347 (N_3347,N_2707,N_2828);
or U3348 (N_3348,N_2832,N_2784);
nand U3349 (N_3349,N_2752,N_2647);
nand U3350 (N_3350,N_2756,N_2859);
or U3351 (N_3351,N_2781,N_2889);
or U3352 (N_3352,N_2569,N_2557);
or U3353 (N_3353,N_2988,N_2602);
or U3354 (N_3354,N_2733,N_2752);
nand U3355 (N_3355,N_2544,N_2725);
and U3356 (N_3356,N_2997,N_2766);
or U3357 (N_3357,N_2806,N_2894);
xnor U3358 (N_3358,N_2709,N_2805);
nor U3359 (N_3359,N_2689,N_2622);
nand U3360 (N_3360,N_2937,N_2721);
or U3361 (N_3361,N_2723,N_2514);
and U3362 (N_3362,N_2881,N_2772);
nor U3363 (N_3363,N_2806,N_2834);
or U3364 (N_3364,N_2638,N_2857);
nand U3365 (N_3365,N_2518,N_2587);
and U3366 (N_3366,N_2533,N_2933);
xnor U3367 (N_3367,N_2605,N_2561);
xnor U3368 (N_3368,N_2611,N_2892);
nor U3369 (N_3369,N_2900,N_2654);
nand U3370 (N_3370,N_2637,N_2987);
or U3371 (N_3371,N_2998,N_2694);
or U3372 (N_3372,N_2545,N_2606);
and U3373 (N_3373,N_2504,N_2613);
nor U3374 (N_3374,N_2756,N_2600);
or U3375 (N_3375,N_2743,N_2523);
xnor U3376 (N_3376,N_2734,N_2621);
nor U3377 (N_3377,N_2862,N_2547);
or U3378 (N_3378,N_2883,N_2572);
and U3379 (N_3379,N_2989,N_2667);
and U3380 (N_3380,N_2862,N_2850);
xor U3381 (N_3381,N_2851,N_2969);
xnor U3382 (N_3382,N_2555,N_2502);
nor U3383 (N_3383,N_2502,N_2710);
and U3384 (N_3384,N_2641,N_2721);
nand U3385 (N_3385,N_2516,N_2937);
nor U3386 (N_3386,N_2890,N_2996);
and U3387 (N_3387,N_2626,N_2817);
nor U3388 (N_3388,N_2841,N_2943);
or U3389 (N_3389,N_2789,N_2767);
nand U3390 (N_3390,N_2949,N_2867);
or U3391 (N_3391,N_2998,N_2970);
xor U3392 (N_3392,N_2880,N_2941);
or U3393 (N_3393,N_2997,N_2968);
and U3394 (N_3394,N_2562,N_2991);
nand U3395 (N_3395,N_2668,N_2965);
nor U3396 (N_3396,N_2850,N_2665);
nand U3397 (N_3397,N_2525,N_2955);
xor U3398 (N_3398,N_2944,N_2640);
and U3399 (N_3399,N_2869,N_2879);
nand U3400 (N_3400,N_2779,N_2573);
nor U3401 (N_3401,N_2722,N_2755);
nor U3402 (N_3402,N_2589,N_2597);
nor U3403 (N_3403,N_2695,N_2835);
or U3404 (N_3404,N_2761,N_2947);
or U3405 (N_3405,N_2667,N_2962);
or U3406 (N_3406,N_2841,N_2649);
nor U3407 (N_3407,N_2622,N_2546);
nor U3408 (N_3408,N_2879,N_2826);
xnor U3409 (N_3409,N_2829,N_2834);
xor U3410 (N_3410,N_2679,N_2869);
or U3411 (N_3411,N_2762,N_2930);
and U3412 (N_3412,N_2795,N_2878);
nand U3413 (N_3413,N_2998,N_2739);
nand U3414 (N_3414,N_2617,N_2762);
and U3415 (N_3415,N_2733,N_2945);
and U3416 (N_3416,N_2826,N_2956);
or U3417 (N_3417,N_2660,N_2839);
and U3418 (N_3418,N_2599,N_2855);
and U3419 (N_3419,N_2676,N_2622);
and U3420 (N_3420,N_2895,N_2623);
and U3421 (N_3421,N_2781,N_2721);
nor U3422 (N_3422,N_2769,N_2742);
nor U3423 (N_3423,N_2741,N_2665);
and U3424 (N_3424,N_2837,N_2640);
xnor U3425 (N_3425,N_2865,N_2736);
or U3426 (N_3426,N_2652,N_2660);
and U3427 (N_3427,N_2529,N_2878);
nand U3428 (N_3428,N_2781,N_2583);
or U3429 (N_3429,N_2827,N_2634);
and U3430 (N_3430,N_2569,N_2977);
or U3431 (N_3431,N_2822,N_2510);
nand U3432 (N_3432,N_2874,N_2833);
and U3433 (N_3433,N_2723,N_2992);
xnor U3434 (N_3434,N_2850,N_2868);
nand U3435 (N_3435,N_2637,N_2808);
or U3436 (N_3436,N_2507,N_2804);
nand U3437 (N_3437,N_2731,N_2819);
xnor U3438 (N_3438,N_2677,N_2595);
and U3439 (N_3439,N_2831,N_2502);
nor U3440 (N_3440,N_2763,N_2953);
and U3441 (N_3441,N_2808,N_2660);
nor U3442 (N_3442,N_2709,N_2663);
or U3443 (N_3443,N_2914,N_2941);
nand U3444 (N_3444,N_2544,N_2652);
xor U3445 (N_3445,N_2857,N_2604);
nor U3446 (N_3446,N_2787,N_2990);
nor U3447 (N_3447,N_2836,N_2578);
nand U3448 (N_3448,N_2745,N_2878);
and U3449 (N_3449,N_2892,N_2946);
nand U3450 (N_3450,N_2663,N_2573);
nand U3451 (N_3451,N_2775,N_2510);
and U3452 (N_3452,N_2699,N_2582);
xor U3453 (N_3453,N_2697,N_2581);
or U3454 (N_3454,N_2975,N_2817);
and U3455 (N_3455,N_2913,N_2818);
nor U3456 (N_3456,N_2757,N_2867);
or U3457 (N_3457,N_2854,N_2926);
or U3458 (N_3458,N_2860,N_2964);
nand U3459 (N_3459,N_2921,N_2751);
or U3460 (N_3460,N_2733,N_2843);
nor U3461 (N_3461,N_2518,N_2965);
nand U3462 (N_3462,N_2730,N_2835);
nand U3463 (N_3463,N_2673,N_2533);
or U3464 (N_3464,N_2781,N_2996);
or U3465 (N_3465,N_2817,N_2890);
and U3466 (N_3466,N_2774,N_2725);
nor U3467 (N_3467,N_2936,N_2934);
nand U3468 (N_3468,N_2528,N_2593);
nand U3469 (N_3469,N_2933,N_2708);
and U3470 (N_3470,N_2677,N_2729);
nor U3471 (N_3471,N_2645,N_2884);
nand U3472 (N_3472,N_2675,N_2637);
or U3473 (N_3473,N_2800,N_2743);
nor U3474 (N_3474,N_2711,N_2916);
and U3475 (N_3475,N_2533,N_2779);
nor U3476 (N_3476,N_2542,N_2643);
and U3477 (N_3477,N_2652,N_2816);
and U3478 (N_3478,N_2964,N_2554);
or U3479 (N_3479,N_2767,N_2892);
and U3480 (N_3480,N_2758,N_2772);
nand U3481 (N_3481,N_2753,N_2682);
nor U3482 (N_3482,N_2852,N_2991);
nor U3483 (N_3483,N_2593,N_2840);
and U3484 (N_3484,N_2867,N_2880);
and U3485 (N_3485,N_2942,N_2666);
nor U3486 (N_3486,N_2521,N_2836);
and U3487 (N_3487,N_2821,N_2729);
or U3488 (N_3488,N_2654,N_2651);
nor U3489 (N_3489,N_2645,N_2978);
and U3490 (N_3490,N_2629,N_2647);
and U3491 (N_3491,N_2689,N_2901);
xor U3492 (N_3492,N_2694,N_2938);
and U3493 (N_3493,N_2640,N_2901);
nor U3494 (N_3494,N_2686,N_2746);
and U3495 (N_3495,N_2972,N_2623);
or U3496 (N_3496,N_2882,N_2795);
and U3497 (N_3497,N_2744,N_2813);
and U3498 (N_3498,N_2509,N_2517);
nand U3499 (N_3499,N_2863,N_2742);
and U3500 (N_3500,N_3157,N_3192);
nand U3501 (N_3501,N_3073,N_3079);
nand U3502 (N_3502,N_3323,N_3200);
nor U3503 (N_3503,N_3242,N_3400);
or U3504 (N_3504,N_3089,N_3003);
nand U3505 (N_3505,N_3229,N_3091);
xnor U3506 (N_3506,N_3189,N_3288);
nand U3507 (N_3507,N_3343,N_3130);
nand U3508 (N_3508,N_3397,N_3252);
nand U3509 (N_3509,N_3456,N_3396);
nand U3510 (N_3510,N_3218,N_3096);
nand U3511 (N_3511,N_3086,N_3271);
nand U3512 (N_3512,N_3162,N_3384);
or U3513 (N_3513,N_3365,N_3195);
nor U3514 (N_3514,N_3301,N_3366);
nor U3515 (N_3515,N_3125,N_3029);
nor U3516 (N_3516,N_3101,N_3220);
nor U3517 (N_3517,N_3449,N_3175);
and U3518 (N_3518,N_3196,N_3420);
nand U3519 (N_3519,N_3442,N_3163);
and U3520 (N_3520,N_3121,N_3497);
nor U3521 (N_3521,N_3124,N_3139);
nor U3522 (N_3522,N_3174,N_3466);
nand U3523 (N_3523,N_3487,N_3117);
or U3524 (N_3524,N_3319,N_3007);
or U3525 (N_3525,N_3006,N_3374);
nor U3526 (N_3526,N_3053,N_3055);
nand U3527 (N_3527,N_3338,N_3309);
nand U3528 (N_3528,N_3041,N_3186);
or U3529 (N_3529,N_3226,N_3092);
and U3530 (N_3530,N_3077,N_3326);
nor U3531 (N_3531,N_3132,N_3317);
nor U3532 (N_3532,N_3280,N_3316);
and U3533 (N_3533,N_3274,N_3215);
nand U3534 (N_3534,N_3263,N_3257);
nor U3535 (N_3535,N_3310,N_3403);
nand U3536 (N_3536,N_3122,N_3388);
and U3537 (N_3537,N_3005,N_3234);
nor U3538 (N_3538,N_3232,N_3045);
or U3539 (N_3539,N_3284,N_3430);
nor U3540 (N_3540,N_3297,N_3399);
and U3541 (N_3541,N_3455,N_3467);
and U3542 (N_3542,N_3231,N_3290);
and U3543 (N_3543,N_3225,N_3152);
nor U3544 (N_3544,N_3415,N_3219);
nor U3545 (N_3545,N_3034,N_3390);
or U3546 (N_3546,N_3472,N_3193);
or U3547 (N_3547,N_3134,N_3318);
xor U3548 (N_3548,N_3459,N_3008);
nor U3549 (N_3549,N_3105,N_3362);
and U3550 (N_3550,N_3372,N_3253);
nand U3551 (N_3551,N_3462,N_3227);
or U3552 (N_3552,N_3141,N_3037);
or U3553 (N_3553,N_3367,N_3416);
and U3554 (N_3554,N_3019,N_3381);
or U3555 (N_3555,N_3216,N_3081);
nor U3556 (N_3556,N_3346,N_3294);
nor U3557 (N_3557,N_3247,N_3431);
and U3558 (N_3558,N_3061,N_3350);
nand U3559 (N_3559,N_3046,N_3114);
nor U3560 (N_3560,N_3417,N_3217);
or U3561 (N_3561,N_3022,N_3410);
or U3562 (N_3562,N_3481,N_3230);
xor U3563 (N_3563,N_3123,N_3491);
nand U3564 (N_3564,N_3389,N_3460);
nand U3565 (N_3565,N_3398,N_3426);
nor U3566 (N_3566,N_3382,N_3475);
nand U3567 (N_3567,N_3210,N_3349);
and U3568 (N_3568,N_3048,N_3205);
xor U3569 (N_3569,N_3348,N_3411);
nand U3570 (N_3570,N_3289,N_3413);
and U3571 (N_3571,N_3213,N_3333);
nand U3572 (N_3572,N_3379,N_3102);
nor U3573 (N_3573,N_3276,N_3080);
xnor U3574 (N_3574,N_3255,N_3357);
xor U3575 (N_3575,N_3119,N_3039);
xor U3576 (N_3576,N_3261,N_3451);
or U3577 (N_3577,N_3228,N_3441);
and U3578 (N_3578,N_3116,N_3058);
nand U3579 (N_3579,N_3070,N_3407);
and U3580 (N_3580,N_3044,N_3111);
nand U3581 (N_3581,N_3243,N_3069);
nand U3582 (N_3582,N_3260,N_3206);
or U3583 (N_3583,N_3386,N_3298);
nand U3584 (N_3584,N_3265,N_3304);
and U3585 (N_3585,N_3408,N_3394);
nor U3586 (N_3586,N_3401,N_3015);
and U3587 (N_3587,N_3203,N_3207);
or U3588 (N_3588,N_3340,N_3402);
nand U3589 (N_3589,N_3282,N_3308);
nor U3590 (N_3590,N_3075,N_3158);
and U3591 (N_3591,N_3036,N_3393);
or U3592 (N_3592,N_3392,N_3178);
nand U3593 (N_3593,N_3352,N_3236);
and U3594 (N_3594,N_3454,N_3358);
nand U3595 (N_3595,N_3090,N_3306);
nor U3596 (N_3596,N_3469,N_3238);
and U3597 (N_3597,N_3001,N_3468);
xnor U3598 (N_3598,N_3115,N_3097);
nand U3599 (N_3599,N_3272,N_3251);
or U3600 (N_3600,N_3083,N_3273);
or U3601 (N_3601,N_3427,N_3136);
nand U3602 (N_3602,N_3143,N_3355);
nor U3603 (N_3603,N_3214,N_3336);
nor U3604 (N_3604,N_3328,N_3364);
nor U3605 (N_3605,N_3423,N_3324);
nor U3606 (N_3606,N_3153,N_3464);
nand U3607 (N_3607,N_3470,N_3342);
nand U3608 (N_3608,N_3054,N_3100);
nand U3609 (N_3609,N_3445,N_3154);
and U3610 (N_3610,N_3293,N_3063);
and U3611 (N_3611,N_3068,N_3444);
and U3612 (N_3612,N_3223,N_3076);
or U3613 (N_3613,N_3176,N_3188);
nand U3614 (N_3614,N_3118,N_3295);
nor U3615 (N_3615,N_3438,N_3126);
xnor U3616 (N_3616,N_3237,N_3275);
and U3617 (N_3617,N_3485,N_3099);
and U3618 (N_3618,N_3002,N_3179);
and U3619 (N_3619,N_3133,N_3016);
and U3620 (N_3620,N_3110,N_3313);
nand U3621 (N_3621,N_3248,N_3047);
nor U3622 (N_3622,N_3279,N_3359);
and U3623 (N_3623,N_3199,N_3221);
or U3624 (N_3624,N_3440,N_3000);
or U3625 (N_3625,N_3320,N_3138);
and U3626 (N_3626,N_3190,N_3373);
nand U3627 (N_3627,N_3021,N_3361);
nand U3628 (N_3628,N_3249,N_3033);
and U3629 (N_3629,N_3065,N_3254);
and U3630 (N_3630,N_3183,N_3377);
or U3631 (N_3631,N_3109,N_3267);
and U3632 (N_3632,N_3287,N_3406);
or U3633 (N_3633,N_3233,N_3281);
or U3634 (N_3634,N_3093,N_3378);
nand U3635 (N_3635,N_3160,N_3197);
and U3636 (N_3636,N_3159,N_3018);
or U3637 (N_3637,N_3329,N_3014);
and U3638 (N_3638,N_3347,N_3030);
nand U3639 (N_3639,N_3250,N_3494);
nor U3640 (N_3640,N_3339,N_3478);
and U3641 (N_3641,N_3314,N_3270);
or U3642 (N_3642,N_3443,N_3151);
and U3643 (N_3643,N_3480,N_3296);
or U3644 (N_3644,N_3148,N_3269);
and U3645 (N_3645,N_3483,N_3439);
nand U3646 (N_3646,N_3020,N_3062);
and U3647 (N_3647,N_3170,N_3173);
nor U3648 (N_3648,N_3064,N_3165);
nand U3649 (N_3649,N_3049,N_3038);
and U3650 (N_3650,N_3493,N_3421);
xor U3651 (N_3651,N_3057,N_3259);
nand U3652 (N_3652,N_3245,N_3424);
nand U3653 (N_3653,N_3476,N_3147);
or U3654 (N_3654,N_3428,N_3127);
or U3655 (N_3655,N_3448,N_3375);
nor U3656 (N_3656,N_3258,N_3180);
or U3657 (N_3657,N_3129,N_3322);
and U3658 (N_3658,N_3344,N_3409);
nand U3659 (N_3659,N_3369,N_3161);
nand U3660 (N_3660,N_3286,N_3164);
xnor U3661 (N_3661,N_3325,N_3351);
nor U3662 (N_3662,N_3473,N_3465);
nand U3663 (N_3663,N_3050,N_3332);
nor U3664 (N_3664,N_3078,N_3060);
xnor U3665 (N_3665,N_3471,N_3435);
and U3666 (N_3666,N_3177,N_3071);
or U3667 (N_3667,N_3376,N_3458);
nor U3668 (N_3668,N_3484,N_3302);
or U3669 (N_3669,N_3330,N_3026);
and U3670 (N_3670,N_3490,N_3385);
and U3671 (N_3671,N_3149,N_3321);
nor U3672 (N_3672,N_3202,N_3447);
and U3673 (N_3673,N_3285,N_3433);
nand U3674 (N_3674,N_3204,N_3341);
and U3675 (N_3675,N_3169,N_3354);
nor U3676 (N_3676,N_3266,N_3425);
xnor U3677 (N_3677,N_3395,N_3477);
or U3678 (N_3678,N_3434,N_3488);
and U3679 (N_3679,N_3419,N_3268);
nor U3680 (N_3680,N_3040,N_3499);
or U3681 (N_3681,N_3144,N_3067);
nor U3682 (N_3682,N_3235,N_3299);
nand U3683 (N_3683,N_3224,N_3017);
xor U3684 (N_3684,N_3042,N_3140);
nor U3685 (N_3685,N_3283,N_3131);
nor U3686 (N_3686,N_3305,N_3356);
nand U3687 (N_3687,N_3201,N_3031);
nand U3688 (N_3688,N_3412,N_3166);
xnor U3689 (N_3689,N_3052,N_3422);
xnor U3690 (N_3690,N_3498,N_3262);
xor U3691 (N_3691,N_3155,N_3387);
or U3692 (N_3692,N_3292,N_3012);
nor U3693 (N_3693,N_3404,N_3185);
xor U3694 (N_3694,N_3345,N_3461);
nand U3695 (N_3695,N_3380,N_3331);
nand U3696 (N_3696,N_3011,N_3450);
nor U3697 (N_3697,N_3150,N_3327);
xor U3698 (N_3698,N_3437,N_3209);
nor U3699 (N_3699,N_3056,N_3107);
or U3700 (N_3700,N_3277,N_3264);
nand U3701 (N_3701,N_3194,N_3446);
nor U3702 (N_3702,N_3168,N_3010);
nand U3703 (N_3703,N_3212,N_3146);
nor U3704 (N_3704,N_3051,N_3391);
nand U3705 (N_3705,N_3240,N_3241);
nor U3706 (N_3706,N_3479,N_3486);
nor U3707 (N_3707,N_3104,N_3337);
nand U3708 (N_3708,N_3072,N_3429);
and U3709 (N_3709,N_3106,N_3187);
and U3710 (N_3710,N_3082,N_3436);
nand U3711 (N_3711,N_3315,N_3004);
nor U3712 (N_3712,N_3098,N_3360);
or U3713 (N_3713,N_3208,N_3492);
xor U3714 (N_3714,N_3135,N_3156);
xor U3715 (N_3715,N_3244,N_3085);
or U3716 (N_3716,N_3495,N_3463);
nor U3717 (N_3717,N_3088,N_3432);
nand U3718 (N_3718,N_3094,N_3043);
nand U3719 (N_3719,N_3084,N_3167);
nor U3720 (N_3720,N_3027,N_3311);
nand U3721 (N_3721,N_3383,N_3137);
or U3722 (N_3722,N_3103,N_3452);
or U3723 (N_3723,N_3108,N_3182);
nor U3724 (N_3724,N_3095,N_3489);
or U3725 (N_3725,N_3278,N_3353);
and U3726 (N_3726,N_3307,N_3457);
nor U3727 (N_3727,N_3112,N_3246);
nor U3728 (N_3728,N_3368,N_3184);
or U3729 (N_3729,N_3172,N_3145);
nor U3730 (N_3730,N_3303,N_3113);
nand U3731 (N_3731,N_3418,N_3474);
nor U3732 (N_3732,N_3066,N_3256);
and U3733 (N_3733,N_3059,N_3171);
and U3734 (N_3734,N_3370,N_3291);
nand U3735 (N_3735,N_3198,N_3363);
nor U3736 (N_3736,N_3414,N_3142);
nor U3737 (N_3737,N_3087,N_3032);
xor U3738 (N_3738,N_3024,N_3334);
nor U3739 (N_3739,N_3312,N_3023);
and U3740 (N_3740,N_3028,N_3035);
or U3741 (N_3741,N_3496,N_3025);
and U3742 (N_3742,N_3191,N_3181);
nand U3743 (N_3743,N_3222,N_3335);
or U3744 (N_3744,N_3013,N_3074);
and U3745 (N_3745,N_3211,N_3009);
nand U3746 (N_3746,N_3120,N_3128);
nor U3747 (N_3747,N_3482,N_3300);
or U3748 (N_3748,N_3405,N_3371);
nand U3749 (N_3749,N_3453,N_3239);
or U3750 (N_3750,N_3028,N_3139);
nor U3751 (N_3751,N_3184,N_3277);
xnor U3752 (N_3752,N_3447,N_3398);
or U3753 (N_3753,N_3270,N_3039);
or U3754 (N_3754,N_3264,N_3117);
and U3755 (N_3755,N_3369,N_3397);
or U3756 (N_3756,N_3120,N_3156);
nand U3757 (N_3757,N_3290,N_3173);
nand U3758 (N_3758,N_3285,N_3219);
xnor U3759 (N_3759,N_3059,N_3498);
or U3760 (N_3760,N_3283,N_3282);
nand U3761 (N_3761,N_3098,N_3122);
and U3762 (N_3762,N_3388,N_3029);
and U3763 (N_3763,N_3064,N_3292);
or U3764 (N_3764,N_3493,N_3123);
nor U3765 (N_3765,N_3306,N_3202);
nand U3766 (N_3766,N_3051,N_3246);
nand U3767 (N_3767,N_3060,N_3432);
or U3768 (N_3768,N_3191,N_3119);
or U3769 (N_3769,N_3302,N_3102);
and U3770 (N_3770,N_3321,N_3315);
and U3771 (N_3771,N_3140,N_3432);
nor U3772 (N_3772,N_3081,N_3143);
or U3773 (N_3773,N_3368,N_3342);
nor U3774 (N_3774,N_3044,N_3025);
nor U3775 (N_3775,N_3242,N_3226);
or U3776 (N_3776,N_3151,N_3357);
or U3777 (N_3777,N_3159,N_3394);
and U3778 (N_3778,N_3183,N_3462);
and U3779 (N_3779,N_3379,N_3192);
and U3780 (N_3780,N_3292,N_3203);
and U3781 (N_3781,N_3347,N_3412);
and U3782 (N_3782,N_3488,N_3451);
xnor U3783 (N_3783,N_3450,N_3352);
xnor U3784 (N_3784,N_3324,N_3178);
or U3785 (N_3785,N_3045,N_3473);
or U3786 (N_3786,N_3144,N_3213);
and U3787 (N_3787,N_3360,N_3170);
xnor U3788 (N_3788,N_3012,N_3186);
nand U3789 (N_3789,N_3397,N_3498);
xnor U3790 (N_3790,N_3233,N_3237);
nand U3791 (N_3791,N_3190,N_3179);
or U3792 (N_3792,N_3134,N_3282);
nand U3793 (N_3793,N_3433,N_3280);
and U3794 (N_3794,N_3498,N_3179);
and U3795 (N_3795,N_3237,N_3301);
or U3796 (N_3796,N_3467,N_3286);
or U3797 (N_3797,N_3283,N_3018);
nor U3798 (N_3798,N_3223,N_3194);
or U3799 (N_3799,N_3017,N_3210);
nand U3800 (N_3800,N_3408,N_3113);
xor U3801 (N_3801,N_3250,N_3459);
nand U3802 (N_3802,N_3485,N_3408);
xor U3803 (N_3803,N_3365,N_3164);
xor U3804 (N_3804,N_3033,N_3225);
and U3805 (N_3805,N_3303,N_3252);
and U3806 (N_3806,N_3419,N_3302);
and U3807 (N_3807,N_3437,N_3277);
or U3808 (N_3808,N_3126,N_3055);
or U3809 (N_3809,N_3051,N_3133);
xnor U3810 (N_3810,N_3300,N_3264);
and U3811 (N_3811,N_3212,N_3455);
xnor U3812 (N_3812,N_3269,N_3211);
and U3813 (N_3813,N_3042,N_3309);
nor U3814 (N_3814,N_3249,N_3288);
nor U3815 (N_3815,N_3057,N_3476);
nand U3816 (N_3816,N_3235,N_3081);
nor U3817 (N_3817,N_3144,N_3282);
nand U3818 (N_3818,N_3109,N_3151);
or U3819 (N_3819,N_3477,N_3126);
nor U3820 (N_3820,N_3395,N_3167);
and U3821 (N_3821,N_3246,N_3459);
or U3822 (N_3822,N_3118,N_3094);
or U3823 (N_3823,N_3411,N_3093);
and U3824 (N_3824,N_3100,N_3146);
nor U3825 (N_3825,N_3112,N_3262);
or U3826 (N_3826,N_3141,N_3051);
nand U3827 (N_3827,N_3461,N_3177);
and U3828 (N_3828,N_3486,N_3499);
nand U3829 (N_3829,N_3399,N_3043);
and U3830 (N_3830,N_3115,N_3161);
nand U3831 (N_3831,N_3090,N_3289);
or U3832 (N_3832,N_3484,N_3392);
and U3833 (N_3833,N_3447,N_3112);
and U3834 (N_3834,N_3318,N_3026);
nor U3835 (N_3835,N_3137,N_3284);
nor U3836 (N_3836,N_3044,N_3328);
and U3837 (N_3837,N_3353,N_3005);
nor U3838 (N_3838,N_3357,N_3285);
or U3839 (N_3839,N_3161,N_3450);
nand U3840 (N_3840,N_3018,N_3180);
and U3841 (N_3841,N_3478,N_3326);
nor U3842 (N_3842,N_3125,N_3242);
nor U3843 (N_3843,N_3021,N_3144);
nand U3844 (N_3844,N_3091,N_3297);
xor U3845 (N_3845,N_3256,N_3058);
or U3846 (N_3846,N_3325,N_3134);
nor U3847 (N_3847,N_3475,N_3446);
or U3848 (N_3848,N_3208,N_3100);
nand U3849 (N_3849,N_3104,N_3239);
nor U3850 (N_3850,N_3216,N_3326);
nand U3851 (N_3851,N_3015,N_3086);
or U3852 (N_3852,N_3187,N_3173);
and U3853 (N_3853,N_3212,N_3274);
and U3854 (N_3854,N_3219,N_3160);
xor U3855 (N_3855,N_3319,N_3281);
nor U3856 (N_3856,N_3088,N_3209);
nor U3857 (N_3857,N_3013,N_3120);
nand U3858 (N_3858,N_3315,N_3207);
or U3859 (N_3859,N_3230,N_3462);
nand U3860 (N_3860,N_3095,N_3025);
nand U3861 (N_3861,N_3338,N_3132);
and U3862 (N_3862,N_3244,N_3106);
or U3863 (N_3863,N_3434,N_3326);
nand U3864 (N_3864,N_3115,N_3118);
or U3865 (N_3865,N_3410,N_3475);
nand U3866 (N_3866,N_3285,N_3027);
and U3867 (N_3867,N_3044,N_3193);
nor U3868 (N_3868,N_3173,N_3440);
or U3869 (N_3869,N_3450,N_3375);
nand U3870 (N_3870,N_3230,N_3092);
nand U3871 (N_3871,N_3082,N_3220);
or U3872 (N_3872,N_3444,N_3497);
or U3873 (N_3873,N_3455,N_3318);
nor U3874 (N_3874,N_3244,N_3435);
or U3875 (N_3875,N_3269,N_3005);
or U3876 (N_3876,N_3242,N_3464);
and U3877 (N_3877,N_3075,N_3377);
and U3878 (N_3878,N_3270,N_3048);
nor U3879 (N_3879,N_3347,N_3363);
nand U3880 (N_3880,N_3043,N_3198);
or U3881 (N_3881,N_3364,N_3061);
nor U3882 (N_3882,N_3164,N_3027);
nand U3883 (N_3883,N_3165,N_3336);
nor U3884 (N_3884,N_3191,N_3324);
nand U3885 (N_3885,N_3400,N_3208);
and U3886 (N_3886,N_3286,N_3144);
and U3887 (N_3887,N_3432,N_3351);
nor U3888 (N_3888,N_3398,N_3042);
or U3889 (N_3889,N_3103,N_3322);
nor U3890 (N_3890,N_3340,N_3308);
and U3891 (N_3891,N_3278,N_3129);
nand U3892 (N_3892,N_3366,N_3150);
and U3893 (N_3893,N_3070,N_3092);
nor U3894 (N_3894,N_3101,N_3407);
and U3895 (N_3895,N_3356,N_3383);
or U3896 (N_3896,N_3010,N_3242);
nand U3897 (N_3897,N_3173,N_3073);
or U3898 (N_3898,N_3108,N_3398);
or U3899 (N_3899,N_3475,N_3224);
and U3900 (N_3900,N_3307,N_3343);
nor U3901 (N_3901,N_3077,N_3255);
or U3902 (N_3902,N_3359,N_3167);
nor U3903 (N_3903,N_3228,N_3429);
nor U3904 (N_3904,N_3157,N_3087);
or U3905 (N_3905,N_3466,N_3464);
nor U3906 (N_3906,N_3335,N_3084);
xnor U3907 (N_3907,N_3324,N_3041);
and U3908 (N_3908,N_3406,N_3054);
and U3909 (N_3909,N_3424,N_3350);
or U3910 (N_3910,N_3181,N_3144);
nor U3911 (N_3911,N_3478,N_3388);
nor U3912 (N_3912,N_3358,N_3202);
and U3913 (N_3913,N_3111,N_3330);
nand U3914 (N_3914,N_3028,N_3099);
or U3915 (N_3915,N_3313,N_3493);
nand U3916 (N_3916,N_3003,N_3197);
xnor U3917 (N_3917,N_3097,N_3118);
or U3918 (N_3918,N_3498,N_3169);
nor U3919 (N_3919,N_3165,N_3470);
nor U3920 (N_3920,N_3146,N_3009);
and U3921 (N_3921,N_3063,N_3294);
nor U3922 (N_3922,N_3479,N_3402);
nor U3923 (N_3923,N_3165,N_3071);
or U3924 (N_3924,N_3358,N_3147);
xnor U3925 (N_3925,N_3033,N_3270);
nand U3926 (N_3926,N_3337,N_3287);
or U3927 (N_3927,N_3397,N_3233);
nand U3928 (N_3928,N_3456,N_3112);
nand U3929 (N_3929,N_3349,N_3247);
nand U3930 (N_3930,N_3255,N_3101);
and U3931 (N_3931,N_3471,N_3016);
nand U3932 (N_3932,N_3487,N_3399);
and U3933 (N_3933,N_3048,N_3466);
nand U3934 (N_3934,N_3038,N_3285);
nor U3935 (N_3935,N_3110,N_3153);
nand U3936 (N_3936,N_3181,N_3054);
nand U3937 (N_3937,N_3146,N_3399);
nand U3938 (N_3938,N_3480,N_3014);
nand U3939 (N_3939,N_3430,N_3385);
or U3940 (N_3940,N_3339,N_3452);
nand U3941 (N_3941,N_3258,N_3344);
or U3942 (N_3942,N_3436,N_3453);
nand U3943 (N_3943,N_3430,N_3471);
nand U3944 (N_3944,N_3076,N_3322);
xor U3945 (N_3945,N_3238,N_3437);
xor U3946 (N_3946,N_3156,N_3112);
xor U3947 (N_3947,N_3355,N_3480);
and U3948 (N_3948,N_3075,N_3488);
nor U3949 (N_3949,N_3195,N_3070);
xnor U3950 (N_3950,N_3405,N_3159);
nand U3951 (N_3951,N_3468,N_3347);
and U3952 (N_3952,N_3206,N_3042);
nor U3953 (N_3953,N_3468,N_3279);
or U3954 (N_3954,N_3009,N_3036);
nand U3955 (N_3955,N_3186,N_3471);
nor U3956 (N_3956,N_3459,N_3035);
and U3957 (N_3957,N_3459,N_3225);
nor U3958 (N_3958,N_3032,N_3119);
nor U3959 (N_3959,N_3470,N_3390);
nand U3960 (N_3960,N_3182,N_3131);
and U3961 (N_3961,N_3426,N_3177);
nand U3962 (N_3962,N_3088,N_3285);
and U3963 (N_3963,N_3371,N_3246);
nor U3964 (N_3964,N_3334,N_3439);
or U3965 (N_3965,N_3398,N_3262);
nor U3966 (N_3966,N_3193,N_3182);
or U3967 (N_3967,N_3487,N_3381);
xor U3968 (N_3968,N_3233,N_3474);
or U3969 (N_3969,N_3191,N_3078);
nor U3970 (N_3970,N_3218,N_3280);
or U3971 (N_3971,N_3366,N_3225);
nand U3972 (N_3972,N_3436,N_3402);
nor U3973 (N_3973,N_3079,N_3056);
and U3974 (N_3974,N_3472,N_3264);
and U3975 (N_3975,N_3377,N_3378);
or U3976 (N_3976,N_3288,N_3280);
and U3977 (N_3977,N_3120,N_3359);
nand U3978 (N_3978,N_3498,N_3304);
nand U3979 (N_3979,N_3297,N_3229);
nor U3980 (N_3980,N_3432,N_3446);
xor U3981 (N_3981,N_3102,N_3064);
and U3982 (N_3982,N_3217,N_3199);
or U3983 (N_3983,N_3207,N_3233);
and U3984 (N_3984,N_3434,N_3037);
nor U3985 (N_3985,N_3378,N_3031);
and U3986 (N_3986,N_3430,N_3398);
nor U3987 (N_3987,N_3357,N_3332);
nor U3988 (N_3988,N_3269,N_3184);
xor U3989 (N_3989,N_3379,N_3163);
nand U3990 (N_3990,N_3196,N_3211);
nand U3991 (N_3991,N_3165,N_3024);
and U3992 (N_3992,N_3069,N_3242);
nor U3993 (N_3993,N_3400,N_3130);
nor U3994 (N_3994,N_3392,N_3285);
nor U3995 (N_3995,N_3092,N_3239);
and U3996 (N_3996,N_3034,N_3366);
or U3997 (N_3997,N_3126,N_3086);
and U3998 (N_3998,N_3074,N_3213);
or U3999 (N_3999,N_3105,N_3021);
nand U4000 (N_4000,N_3634,N_3520);
or U4001 (N_4001,N_3991,N_3593);
or U4002 (N_4002,N_3856,N_3512);
or U4003 (N_4003,N_3891,N_3502);
xor U4004 (N_4004,N_3691,N_3849);
and U4005 (N_4005,N_3610,N_3730);
or U4006 (N_4006,N_3548,N_3619);
nand U4007 (N_4007,N_3846,N_3763);
nor U4008 (N_4008,N_3901,N_3716);
xor U4009 (N_4009,N_3889,N_3776);
nor U4010 (N_4010,N_3981,N_3818);
and U4011 (N_4011,N_3959,N_3808);
nand U4012 (N_4012,N_3890,N_3822);
nand U4013 (N_4013,N_3695,N_3706);
nand U4014 (N_4014,N_3598,N_3838);
or U4015 (N_4015,N_3579,N_3554);
nor U4016 (N_4016,N_3774,N_3560);
nor U4017 (N_4017,N_3814,N_3577);
and U4018 (N_4018,N_3642,N_3592);
or U4019 (N_4019,N_3793,N_3865);
nand U4020 (N_4020,N_3601,N_3907);
xnor U4021 (N_4021,N_3905,N_3727);
nand U4022 (N_4022,N_3582,N_3569);
xnor U4023 (N_4023,N_3513,N_3875);
or U4024 (N_4024,N_3982,N_3500);
nand U4025 (N_4025,N_3783,N_3717);
nor U4026 (N_4026,N_3650,N_3511);
xnor U4027 (N_4027,N_3723,N_3769);
nand U4028 (N_4028,N_3969,N_3620);
nand U4029 (N_4029,N_3622,N_3536);
or U4030 (N_4030,N_3702,N_3629);
nand U4031 (N_4031,N_3874,N_3694);
and U4032 (N_4032,N_3683,N_3742);
or U4033 (N_4033,N_3927,N_3603);
nor U4034 (N_4034,N_3854,N_3938);
nand U4035 (N_4035,N_3953,N_3992);
and U4036 (N_4036,N_3597,N_3934);
and U4037 (N_4037,N_3555,N_3613);
or U4038 (N_4038,N_3624,N_3819);
nand U4039 (N_4039,N_3962,N_3711);
and U4040 (N_4040,N_3677,N_3882);
nand U4041 (N_4041,N_3957,N_3584);
xnor U4042 (N_4042,N_3626,N_3858);
nand U4043 (N_4043,N_3954,N_3583);
or U4044 (N_4044,N_3766,N_3750);
nor U4045 (N_4045,N_3964,N_3839);
and U4046 (N_4046,N_3514,N_3649);
xnor U4047 (N_4047,N_3551,N_3754);
and U4048 (N_4048,N_3881,N_3549);
nor U4049 (N_4049,N_3509,N_3698);
nor U4050 (N_4050,N_3563,N_3998);
xnor U4051 (N_4051,N_3581,N_3547);
xnor U4052 (N_4052,N_3524,N_3707);
and U4053 (N_4053,N_3893,N_3987);
nand U4054 (N_4054,N_3872,N_3848);
or U4055 (N_4055,N_3796,N_3712);
and U4056 (N_4056,N_3955,N_3761);
or U4057 (N_4057,N_3956,N_3894);
nor U4058 (N_4058,N_3572,N_3735);
and U4059 (N_4059,N_3724,N_3945);
nor U4060 (N_4060,N_3916,N_3663);
or U4061 (N_4061,N_3672,N_3923);
or U4062 (N_4062,N_3784,N_3625);
and U4063 (N_4063,N_3896,N_3937);
nand U4064 (N_4064,N_3741,N_3713);
nand U4065 (N_4065,N_3952,N_3946);
and U4066 (N_4066,N_3647,N_3505);
nor U4067 (N_4067,N_3725,N_3869);
nor U4068 (N_4068,N_3518,N_3556);
nor U4069 (N_4069,N_3749,N_3704);
and U4070 (N_4070,N_3773,N_3508);
xnor U4071 (N_4071,N_3553,N_3720);
or U4072 (N_4072,N_3503,N_3861);
nor U4073 (N_4073,N_3764,N_3811);
nand U4074 (N_4074,N_3574,N_3616);
nor U4075 (N_4075,N_3633,N_3585);
and U4076 (N_4076,N_3543,N_3950);
nand U4077 (N_4077,N_3900,N_3758);
or U4078 (N_4078,N_3545,N_3636);
nand U4079 (N_4079,N_3605,N_3990);
and U4080 (N_4080,N_3841,N_3664);
and U4081 (N_4081,N_3803,N_3989);
xnor U4082 (N_4082,N_3929,N_3681);
or U4083 (N_4083,N_3604,N_3851);
and U4084 (N_4084,N_3523,N_3996);
nor U4085 (N_4085,N_3732,N_3618);
and U4086 (N_4086,N_3963,N_3570);
or U4087 (N_4087,N_3798,N_3747);
and U4088 (N_4088,N_3842,N_3718);
or U4089 (N_4089,N_3745,N_3837);
and U4090 (N_4090,N_3997,N_3826);
nor U4091 (N_4091,N_3590,N_3654);
or U4092 (N_4092,N_3971,N_3655);
xnor U4093 (N_4093,N_3641,N_3639);
and U4094 (N_4094,N_3596,N_3738);
nor U4095 (N_4095,N_3611,N_3644);
nor U4096 (N_4096,N_3886,N_3740);
nor U4097 (N_4097,N_3544,N_3667);
or U4098 (N_4098,N_3968,N_3507);
and U4099 (N_4099,N_3948,N_3657);
nor U4100 (N_4100,N_3501,N_3831);
or U4101 (N_4101,N_3699,N_3904);
and U4102 (N_4102,N_3791,N_3786);
and U4103 (N_4103,N_3802,N_3692);
xnor U4104 (N_4104,N_3844,N_3974);
or U4105 (N_4105,N_3933,N_3941);
and U4106 (N_4106,N_3534,N_3679);
nand U4107 (N_4107,N_3733,N_3995);
nand U4108 (N_4108,N_3922,N_3794);
and U4109 (N_4109,N_3888,N_3531);
nand U4110 (N_4110,N_3805,N_3777);
and U4111 (N_4111,N_3859,N_3746);
nand U4112 (N_4112,N_3812,N_3669);
nand U4113 (N_4113,N_3748,N_3607);
and U4114 (N_4114,N_3515,N_3873);
and U4115 (N_4115,N_3671,N_3685);
and U4116 (N_4116,N_3516,N_3751);
and U4117 (N_4117,N_3753,N_3744);
and U4118 (N_4118,N_3600,N_3780);
nor U4119 (N_4119,N_3526,N_3715);
or U4120 (N_4120,N_3689,N_3850);
nand U4121 (N_4121,N_3867,N_3845);
nand U4122 (N_4122,N_3662,N_3521);
and U4123 (N_4123,N_3658,N_3883);
and U4124 (N_4124,N_3797,N_3835);
and U4125 (N_4125,N_3862,N_3853);
nor U4126 (N_4126,N_3973,N_3958);
and U4127 (N_4127,N_3972,N_3813);
and U4128 (N_4128,N_3876,N_3529);
and U4129 (N_4129,N_3721,N_3911);
xnor U4130 (N_4130,N_3504,N_3880);
nand U4131 (N_4131,N_3985,N_3586);
nand U4132 (N_4132,N_3756,N_3977);
or U4133 (N_4133,N_3827,N_3980);
nand U4134 (N_4134,N_3631,N_3621);
or U4135 (N_4135,N_3871,N_3617);
or U4136 (N_4136,N_3921,N_3926);
xor U4137 (N_4137,N_3775,N_3860);
xnor U4138 (N_4138,N_3594,N_3628);
and U4139 (N_4139,N_3696,N_3656);
or U4140 (N_4140,N_3868,N_3675);
or U4141 (N_4141,N_3676,N_3944);
and U4142 (N_4142,N_3807,N_3771);
and U4143 (N_4143,N_3895,N_3847);
or U4144 (N_4144,N_3834,N_3668);
xor U4145 (N_4145,N_3726,N_3762);
nand U4146 (N_4146,N_3903,N_3734);
nand U4147 (N_4147,N_3897,N_3918);
or U4148 (N_4148,N_3648,N_3612);
and U4149 (N_4149,N_3510,N_3986);
and U4150 (N_4150,N_3825,N_3552);
nor U4151 (N_4151,N_3930,N_3589);
nand U4152 (N_4152,N_3627,N_3877);
and U4153 (N_4153,N_3866,N_3943);
nor U4154 (N_4154,N_3759,N_3653);
nor U4155 (N_4155,N_3539,N_3722);
nand U4156 (N_4156,N_3898,N_3770);
and U4157 (N_4157,N_3660,N_3737);
nor U4158 (N_4158,N_3863,N_3565);
nand U4159 (N_4159,N_3884,N_3568);
or U4160 (N_4160,N_3994,N_3908);
nor U4161 (N_4161,N_3984,N_3645);
or U4162 (N_4162,N_3815,N_3821);
xnor U4163 (N_4163,N_3525,N_3806);
or U4164 (N_4164,N_3789,N_3787);
or U4165 (N_4165,N_3820,N_3975);
or U4166 (N_4166,N_3540,N_3928);
or U4167 (N_4167,N_3940,N_3580);
nor U4168 (N_4168,N_3527,N_3533);
or U4169 (N_4169,N_3652,N_3832);
and U4170 (N_4170,N_3804,N_3729);
or U4171 (N_4171,N_3799,N_3566);
and U4172 (N_4172,N_3708,N_3693);
xnor U4173 (N_4173,N_3546,N_3537);
and U4174 (N_4174,N_3947,N_3768);
and U4175 (N_4175,N_3782,N_3522);
and U4176 (N_4176,N_3710,N_3714);
and U4177 (N_4177,N_3519,N_3591);
and U4178 (N_4178,N_3638,N_3541);
and U4179 (N_4179,N_3765,N_3942);
or U4180 (N_4180,N_3700,N_3795);
or U4181 (N_4181,N_3678,N_3557);
nand U4182 (N_4182,N_3752,N_3951);
and U4183 (N_4183,N_3912,N_3965);
and U4184 (N_4184,N_3779,N_3673);
and U4185 (N_4185,N_3575,N_3778);
xor U4186 (N_4186,N_3506,N_3757);
and U4187 (N_4187,N_3816,N_3935);
and U4188 (N_4188,N_3760,N_3587);
nand U4189 (N_4189,N_3615,N_3792);
and U4190 (N_4190,N_3767,N_3573);
nand U4191 (N_4191,N_3665,N_3830);
nor U4192 (N_4192,N_3606,N_3632);
and U4193 (N_4193,N_3931,N_3697);
and U4194 (N_4194,N_3785,N_3824);
nor U4195 (N_4195,N_3670,N_3906);
nor U4196 (N_4196,N_3970,N_3801);
nand U4197 (N_4197,N_3703,N_3550);
nand U4198 (N_4198,N_3719,N_3578);
nand U4199 (N_4199,N_3736,N_3640);
or U4200 (N_4200,N_3651,N_3559);
nand U4201 (N_4201,N_3909,N_3978);
or U4202 (N_4202,N_3879,N_3567);
nand U4203 (N_4203,N_3614,N_3686);
xor U4204 (N_4204,N_3637,N_3674);
and U4205 (N_4205,N_3885,N_3661);
nor U4206 (N_4206,N_3932,N_3781);
nand U4207 (N_4207,N_3528,N_3961);
nand U4208 (N_4208,N_3772,N_3680);
nor U4209 (N_4209,N_3562,N_3530);
or U4210 (N_4210,N_3852,N_3517);
xor U4211 (N_4211,N_3983,N_3829);
and U4212 (N_4212,N_3728,N_3608);
nand U4213 (N_4213,N_3659,N_3870);
or U4214 (N_4214,N_3701,N_3892);
or U4215 (N_4215,N_3855,N_3966);
or U4216 (N_4216,N_3690,N_3902);
nor U4217 (N_4217,N_3688,N_3915);
xor U4218 (N_4218,N_3684,N_3833);
xnor U4219 (N_4219,N_3999,N_3817);
or U4220 (N_4220,N_3810,N_3857);
nand U4221 (N_4221,N_3755,N_3682);
and U4222 (N_4222,N_3790,N_3936);
nor U4223 (N_4223,N_3609,N_3705);
or U4224 (N_4224,N_3571,N_3564);
nand U4225 (N_4225,N_3828,N_3635);
nand U4226 (N_4226,N_3843,N_3993);
nand U4227 (N_4227,N_3910,N_3630);
nand U4228 (N_4228,N_3836,N_3920);
or U4229 (N_4229,N_3823,N_3914);
and U4230 (N_4230,N_3887,N_3960);
and U4231 (N_4231,N_3709,N_3576);
nor U4232 (N_4232,N_3939,N_3623);
xor U4233 (N_4233,N_3687,N_3538);
nor U4234 (N_4234,N_3643,N_3602);
or U4235 (N_4235,N_3809,N_3967);
and U4236 (N_4236,N_3917,N_3558);
or U4237 (N_4237,N_3532,N_3595);
and U4238 (N_4238,N_3599,N_3561);
or U4239 (N_4239,N_3743,N_3949);
nor U4240 (N_4240,N_3788,N_3588);
nand U4241 (N_4241,N_3913,N_3864);
and U4242 (N_4242,N_3924,N_3976);
and U4243 (N_4243,N_3535,N_3979);
xnor U4244 (N_4244,N_3988,N_3731);
nor U4245 (N_4245,N_3878,N_3925);
nor U4246 (N_4246,N_3800,N_3739);
nor U4247 (N_4247,N_3646,N_3840);
nor U4248 (N_4248,N_3666,N_3919);
nor U4249 (N_4249,N_3542,N_3899);
xor U4250 (N_4250,N_3602,N_3763);
or U4251 (N_4251,N_3657,N_3867);
and U4252 (N_4252,N_3809,N_3533);
nand U4253 (N_4253,N_3519,N_3532);
and U4254 (N_4254,N_3702,N_3947);
and U4255 (N_4255,N_3788,N_3903);
xor U4256 (N_4256,N_3935,N_3901);
nor U4257 (N_4257,N_3825,N_3679);
nor U4258 (N_4258,N_3631,N_3524);
and U4259 (N_4259,N_3584,N_3691);
nor U4260 (N_4260,N_3506,N_3639);
nor U4261 (N_4261,N_3890,N_3748);
and U4262 (N_4262,N_3992,N_3723);
and U4263 (N_4263,N_3595,N_3742);
and U4264 (N_4264,N_3656,N_3681);
and U4265 (N_4265,N_3609,N_3949);
or U4266 (N_4266,N_3590,N_3548);
and U4267 (N_4267,N_3848,N_3679);
nand U4268 (N_4268,N_3961,N_3873);
nand U4269 (N_4269,N_3851,N_3924);
nand U4270 (N_4270,N_3616,N_3615);
or U4271 (N_4271,N_3604,N_3861);
or U4272 (N_4272,N_3610,N_3708);
xnor U4273 (N_4273,N_3970,N_3699);
nand U4274 (N_4274,N_3513,N_3737);
nand U4275 (N_4275,N_3938,N_3598);
or U4276 (N_4276,N_3669,N_3962);
and U4277 (N_4277,N_3724,N_3791);
and U4278 (N_4278,N_3653,N_3790);
xnor U4279 (N_4279,N_3972,N_3560);
and U4280 (N_4280,N_3902,N_3629);
nand U4281 (N_4281,N_3712,N_3831);
nand U4282 (N_4282,N_3611,N_3539);
and U4283 (N_4283,N_3997,N_3647);
and U4284 (N_4284,N_3670,N_3824);
xnor U4285 (N_4285,N_3846,N_3791);
or U4286 (N_4286,N_3720,N_3802);
nor U4287 (N_4287,N_3869,N_3923);
nor U4288 (N_4288,N_3667,N_3554);
nor U4289 (N_4289,N_3528,N_3545);
xor U4290 (N_4290,N_3692,N_3840);
and U4291 (N_4291,N_3719,N_3900);
or U4292 (N_4292,N_3661,N_3596);
nand U4293 (N_4293,N_3992,N_3729);
nand U4294 (N_4294,N_3992,N_3731);
or U4295 (N_4295,N_3742,N_3902);
xor U4296 (N_4296,N_3977,N_3922);
nand U4297 (N_4297,N_3957,N_3987);
or U4298 (N_4298,N_3675,N_3895);
or U4299 (N_4299,N_3848,N_3879);
nor U4300 (N_4300,N_3700,N_3631);
and U4301 (N_4301,N_3686,N_3814);
nor U4302 (N_4302,N_3761,N_3789);
and U4303 (N_4303,N_3657,N_3597);
nor U4304 (N_4304,N_3715,N_3875);
or U4305 (N_4305,N_3833,N_3687);
nor U4306 (N_4306,N_3904,N_3510);
nand U4307 (N_4307,N_3957,N_3518);
xnor U4308 (N_4308,N_3890,N_3593);
and U4309 (N_4309,N_3892,N_3565);
and U4310 (N_4310,N_3750,N_3736);
nand U4311 (N_4311,N_3915,N_3518);
nor U4312 (N_4312,N_3653,N_3522);
or U4313 (N_4313,N_3664,N_3772);
or U4314 (N_4314,N_3882,N_3809);
and U4315 (N_4315,N_3867,N_3795);
and U4316 (N_4316,N_3680,N_3930);
nor U4317 (N_4317,N_3576,N_3938);
or U4318 (N_4318,N_3500,N_3752);
xor U4319 (N_4319,N_3837,N_3857);
nand U4320 (N_4320,N_3787,N_3519);
nor U4321 (N_4321,N_3790,N_3796);
nor U4322 (N_4322,N_3917,N_3523);
and U4323 (N_4323,N_3741,N_3898);
xor U4324 (N_4324,N_3997,N_3580);
nor U4325 (N_4325,N_3615,N_3597);
and U4326 (N_4326,N_3855,N_3560);
xnor U4327 (N_4327,N_3585,N_3582);
nand U4328 (N_4328,N_3861,N_3844);
nand U4329 (N_4329,N_3789,N_3732);
nand U4330 (N_4330,N_3762,N_3921);
xor U4331 (N_4331,N_3914,N_3642);
nor U4332 (N_4332,N_3738,N_3726);
nand U4333 (N_4333,N_3856,N_3574);
nand U4334 (N_4334,N_3770,N_3673);
xnor U4335 (N_4335,N_3753,N_3772);
or U4336 (N_4336,N_3835,N_3823);
nor U4337 (N_4337,N_3777,N_3946);
nor U4338 (N_4338,N_3502,N_3582);
or U4339 (N_4339,N_3592,N_3784);
xnor U4340 (N_4340,N_3515,N_3724);
nand U4341 (N_4341,N_3781,N_3887);
or U4342 (N_4342,N_3722,N_3696);
or U4343 (N_4343,N_3875,N_3648);
nor U4344 (N_4344,N_3936,N_3726);
and U4345 (N_4345,N_3582,N_3522);
or U4346 (N_4346,N_3998,N_3579);
and U4347 (N_4347,N_3643,N_3778);
and U4348 (N_4348,N_3751,N_3986);
and U4349 (N_4349,N_3628,N_3793);
nor U4350 (N_4350,N_3550,N_3575);
nand U4351 (N_4351,N_3987,N_3750);
xnor U4352 (N_4352,N_3928,N_3748);
and U4353 (N_4353,N_3747,N_3970);
or U4354 (N_4354,N_3817,N_3907);
nor U4355 (N_4355,N_3535,N_3677);
or U4356 (N_4356,N_3530,N_3750);
nor U4357 (N_4357,N_3682,N_3547);
or U4358 (N_4358,N_3952,N_3587);
and U4359 (N_4359,N_3761,N_3961);
nor U4360 (N_4360,N_3816,N_3603);
nand U4361 (N_4361,N_3994,N_3940);
nand U4362 (N_4362,N_3578,N_3583);
xor U4363 (N_4363,N_3783,N_3813);
and U4364 (N_4364,N_3877,N_3551);
and U4365 (N_4365,N_3807,N_3926);
nor U4366 (N_4366,N_3924,N_3986);
nor U4367 (N_4367,N_3844,N_3809);
and U4368 (N_4368,N_3695,N_3628);
xor U4369 (N_4369,N_3742,N_3867);
or U4370 (N_4370,N_3926,N_3788);
nand U4371 (N_4371,N_3517,N_3574);
and U4372 (N_4372,N_3747,N_3715);
nand U4373 (N_4373,N_3649,N_3768);
and U4374 (N_4374,N_3828,N_3839);
or U4375 (N_4375,N_3717,N_3933);
and U4376 (N_4376,N_3741,N_3641);
and U4377 (N_4377,N_3800,N_3726);
nand U4378 (N_4378,N_3815,N_3876);
and U4379 (N_4379,N_3837,N_3777);
nand U4380 (N_4380,N_3903,N_3820);
or U4381 (N_4381,N_3936,N_3695);
or U4382 (N_4382,N_3958,N_3708);
xor U4383 (N_4383,N_3976,N_3502);
or U4384 (N_4384,N_3668,N_3657);
and U4385 (N_4385,N_3556,N_3558);
and U4386 (N_4386,N_3918,N_3841);
and U4387 (N_4387,N_3815,N_3635);
nor U4388 (N_4388,N_3872,N_3650);
nor U4389 (N_4389,N_3954,N_3992);
or U4390 (N_4390,N_3998,N_3799);
or U4391 (N_4391,N_3570,N_3815);
nand U4392 (N_4392,N_3570,N_3942);
nand U4393 (N_4393,N_3786,N_3505);
or U4394 (N_4394,N_3964,N_3644);
xor U4395 (N_4395,N_3710,N_3911);
and U4396 (N_4396,N_3621,N_3636);
nand U4397 (N_4397,N_3738,N_3995);
or U4398 (N_4398,N_3880,N_3592);
or U4399 (N_4399,N_3775,N_3590);
or U4400 (N_4400,N_3598,N_3574);
or U4401 (N_4401,N_3834,N_3872);
nand U4402 (N_4402,N_3587,N_3840);
nand U4403 (N_4403,N_3904,N_3591);
and U4404 (N_4404,N_3742,N_3790);
and U4405 (N_4405,N_3956,N_3962);
nand U4406 (N_4406,N_3929,N_3933);
nor U4407 (N_4407,N_3936,N_3802);
nand U4408 (N_4408,N_3760,N_3651);
nand U4409 (N_4409,N_3721,N_3995);
and U4410 (N_4410,N_3597,N_3603);
nand U4411 (N_4411,N_3644,N_3888);
nor U4412 (N_4412,N_3579,N_3739);
and U4413 (N_4413,N_3680,N_3532);
and U4414 (N_4414,N_3692,N_3838);
or U4415 (N_4415,N_3752,N_3638);
nor U4416 (N_4416,N_3689,N_3724);
nand U4417 (N_4417,N_3638,N_3768);
nand U4418 (N_4418,N_3862,N_3579);
or U4419 (N_4419,N_3703,N_3893);
nand U4420 (N_4420,N_3644,N_3557);
or U4421 (N_4421,N_3914,N_3916);
and U4422 (N_4422,N_3532,N_3749);
nor U4423 (N_4423,N_3654,N_3532);
xor U4424 (N_4424,N_3797,N_3781);
xnor U4425 (N_4425,N_3521,N_3740);
and U4426 (N_4426,N_3709,N_3984);
or U4427 (N_4427,N_3749,N_3869);
nand U4428 (N_4428,N_3595,N_3576);
nor U4429 (N_4429,N_3508,N_3939);
nand U4430 (N_4430,N_3946,N_3607);
and U4431 (N_4431,N_3540,N_3651);
and U4432 (N_4432,N_3538,N_3703);
or U4433 (N_4433,N_3759,N_3824);
nand U4434 (N_4434,N_3813,N_3715);
and U4435 (N_4435,N_3638,N_3598);
nand U4436 (N_4436,N_3833,N_3700);
or U4437 (N_4437,N_3589,N_3591);
xnor U4438 (N_4438,N_3763,N_3634);
or U4439 (N_4439,N_3770,N_3558);
and U4440 (N_4440,N_3579,N_3562);
xor U4441 (N_4441,N_3881,N_3768);
and U4442 (N_4442,N_3953,N_3896);
or U4443 (N_4443,N_3768,N_3583);
nand U4444 (N_4444,N_3842,N_3777);
nor U4445 (N_4445,N_3815,N_3752);
or U4446 (N_4446,N_3836,N_3925);
and U4447 (N_4447,N_3960,N_3996);
or U4448 (N_4448,N_3591,N_3980);
or U4449 (N_4449,N_3609,N_3698);
and U4450 (N_4450,N_3800,N_3805);
xnor U4451 (N_4451,N_3615,N_3847);
and U4452 (N_4452,N_3950,N_3732);
nand U4453 (N_4453,N_3673,N_3679);
or U4454 (N_4454,N_3904,N_3704);
and U4455 (N_4455,N_3598,N_3953);
nor U4456 (N_4456,N_3811,N_3624);
or U4457 (N_4457,N_3796,N_3734);
and U4458 (N_4458,N_3964,N_3749);
nor U4459 (N_4459,N_3640,N_3707);
nand U4460 (N_4460,N_3613,N_3577);
and U4461 (N_4461,N_3844,N_3897);
or U4462 (N_4462,N_3949,N_3646);
nand U4463 (N_4463,N_3566,N_3506);
nand U4464 (N_4464,N_3609,N_3636);
and U4465 (N_4465,N_3776,N_3862);
nor U4466 (N_4466,N_3989,N_3946);
and U4467 (N_4467,N_3766,N_3976);
nor U4468 (N_4468,N_3602,N_3521);
xor U4469 (N_4469,N_3871,N_3905);
nor U4470 (N_4470,N_3536,N_3799);
nand U4471 (N_4471,N_3986,N_3987);
and U4472 (N_4472,N_3953,N_3647);
or U4473 (N_4473,N_3954,N_3629);
and U4474 (N_4474,N_3767,N_3615);
xnor U4475 (N_4475,N_3823,N_3546);
nor U4476 (N_4476,N_3809,N_3872);
nor U4477 (N_4477,N_3928,N_3575);
or U4478 (N_4478,N_3991,N_3669);
and U4479 (N_4479,N_3892,N_3831);
and U4480 (N_4480,N_3807,N_3970);
nor U4481 (N_4481,N_3784,N_3672);
or U4482 (N_4482,N_3881,N_3871);
nand U4483 (N_4483,N_3999,N_3648);
nand U4484 (N_4484,N_3551,N_3524);
or U4485 (N_4485,N_3541,N_3652);
nor U4486 (N_4486,N_3832,N_3574);
nor U4487 (N_4487,N_3595,N_3593);
nand U4488 (N_4488,N_3540,N_3701);
or U4489 (N_4489,N_3730,N_3836);
nor U4490 (N_4490,N_3653,N_3948);
or U4491 (N_4491,N_3751,N_3984);
nor U4492 (N_4492,N_3972,N_3786);
and U4493 (N_4493,N_3609,N_3932);
or U4494 (N_4494,N_3833,N_3842);
xnor U4495 (N_4495,N_3750,N_3899);
or U4496 (N_4496,N_3706,N_3900);
nor U4497 (N_4497,N_3958,N_3563);
or U4498 (N_4498,N_3592,N_3831);
nand U4499 (N_4499,N_3936,N_3716);
and U4500 (N_4500,N_4216,N_4440);
or U4501 (N_4501,N_4226,N_4311);
or U4502 (N_4502,N_4132,N_4228);
or U4503 (N_4503,N_4140,N_4383);
and U4504 (N_4504,N_4125,N_4048);
and U4505 (N_4505,N_4336,N_4263);
nand U4506 (N_4506,N_4200,N_4395);
and U4507 (N_4507,N_4161,N_4445);
and U4508 (N_4508,N_4441,N_4066);
nor U4509 (N_4509,N_4266,N_4317);
or U4510 (N_4510,N_4436,N_4334);
xor U4511 (N_4511,N_4407,N_4337);
nand U4512 (N_4512,N_4284,N_4054);
xor U4513 (N_4513,N_4032,N_4053);
and U4514 (N_4514,N_4398,N_4123);
nor U4515 (N_4515,N_4479,N_4056);
nand U4516 (N_4516,N_4184,N_4260);
or U4517 (N_4517,N_4478,N_4202);
and U4518 (N_4518,N_4307,N_4212);
or U4519 (N_4519,N_4039,N_4232);
nand U4520 (N_4520,N_4370,N_4380);
or U4521 (N_4521,N_4245,N_4325);
nor U4522 (N_4522,N_4406,N_4084);
or U4523 (N_4523,N_4244,N_4328);
nand U4524 (N_4524,N_4483,N_4196);
and U4525 (N_4525,N_4008,N_4168);
and U4526 (N_4526,N_4120,N_4428);
or U4527 (N_4527,N_4220,N_4405);
nor U4528 (N_4528,N_4322,N_4074);
and U4529 (N_4529,N_4018,N_4486);
and U4530 (N_4530,N_4448,N_4189);
nand U4531 (N_4531,N_4111,N_4493);
or U4532 (N_4532,N_4213,N_4136);
nor U4533 (N_4533,N_4484,N_4449);
and U4534 (N_4534,N_4366,N_4078);
or U4535 (N_4535,N_4464,N_4210);
xor U4536 (N_4536,N_4057,N_4319);
and U4537 (N_4537,N_4207,N_4432);
and U4538 (N_4538,N_4062,N_4287);
or U4539 (N_4539,N_4482,N_4270);
and U4540 (N_4540,N_4434,N_4242);
nand U4541 (N_4541,N_4169,N_4102);
nand U4542 (N_4542,N_4218,N_4147);
nor U4543 (N_4543,N_4138,N_4190);
xor U4544 (N_4544,N_4480,N_4193);
nor U4545 (N_4545,N_4352,N_4149);
or U4546 (N_4546,N_4496,N_4064);
nor U4547 (N_4547,N_4122,N_4162);
xnor U4548 (N_4548,N_4238,N_4070);
nor U4549 (N_4549,N_4022,N_4058);
or U4550 (N_4550,N_4429,N_4192);
and U4551 (N_4551,N_4014,N_4153);
and U4552 (N_4552,N_4324,N_4378);
nand U4553 (N_4553,N_4283,N_4485);
or U4554 (N_4554,N_4261,N_4376);
or U4555 (N_4555,N_4451,N_4470);
and U4556 (N_4556,N_4129,N_4180);
nor U4557 (N_4557,N_4155,N_4320);
and U4558 (N_4558,N_4257,N_4060);
nor U4559 (N_4559,N_4049,N_4494);
nor U4560 (N_4560,N_4357,N_4194);
xor U4561 (N_4561,N_4385,N_4025);
and U4562 (N_4562,N_4239,N_4217);
xnor U4563 (N_4563,N_4331,N_4061);
and U4564 (N_4564,N_4401,N_4412);
nand U4565 (N_4565,N_4003,N_4314);
xor U4566 (N_4566,N_4017,N_4041);
or U4567 (N_4567,N_4349,N_4249);
or U4568 (N_4568,N_4291,N_4077);
and U4569 (N_4569,N_4335,N_4312);
nand U4570 (N_4570,N_4420,N_4112);
nor U4571 (N_4571,N_4214,N_4033);
xor U4572 (N_4572,N_4492,N_4069);
nand U4573 (N_4573,N_4150,N_4497);
nand U4574 (N_4574,N_4046,N_4076);
or U4575 (N_4575,N_4124,N_4143);
nor U4576 (N_4576,N_4409,N_4045);
xor U4577 (N_4577,N_4113,N_4297);
and U4578 (N_4578,N_4499,N_4175);
nor U4579 (N_4579,N_4198,N_4354);
nand U4580 (N_4580,N_4462,N_4410);
xor U4581 (N_4581,N_4103,N_4174);
nand U4582 (N_4582,N_4256,N_4002);
xor U4583 (N_4583,N_4438,N_4293);
nand U4584 (N_4584,N_4304,N_4313);
nand U4585 (N_4585,N_4463,N_4182);
nor U4586 (N_4586,N_4344,N_4345);
and U4587 (N_4587,N_4030,N_4443);
nand U4588 (N_4588,N_4197,N_4298);
or U4589 (N_4589,N_4423,N_4036);
and U4590 (N_4590,N_4130,N_4421);
or U4591 (N_4591,N_4170,N_4294);
xor U4592 (N_4592,N_4148,N_4157);
or U4593 (N_4593,N_4404,N_4342);
nor U4594 (N_4594,N_4005,N_4301);
nand U4595 (N_4595,N_4396,N_4173);
and U4596 (N_4596,N_4458,N_4387);
and U4597 (N_4597,N_4021,N_4278);
nor U4598 (N_4598,N_4333,N_4326);
and U4599 (N_4599,N_4348,N_4350);
nand U4600 (N_4600,N_4075,N_4374);
nand U4601 (N_4601,N_4452,N_4177);
xnor U4602 (N_4602,N_4286,N_4364);
and U4603 (N_4603,N_4188,N_4139);
or U4604 (N_4604,N_4063,N_4471);
nand U4605 (N_4605,N_4165,N_4164);
and U4606 (N_4606,N_4183,N_4179);
xnor U4607 (N_4607,N_4158,N_4388);
nand U4608 (N_4608,N_4085,N_4013);
or U4609 (N_4609,N_4365,N_4347);
nor U4610 (N_4610,N_4251,N_4465);
and U4611 (N_4611,N_4230,N_4371);
nand U4612 (N_4612,N_4050,N_4023);
nor U4613 (N_4613,N_4391,N_4394);
nand U4614 (N_4614,N_4431,N_4386);
xor U4615 (N_4615,N_4031,N_4418);
nor U4616 (N_4616,N_4040,N_4456);
or U4617 (N_4617,N_4302,N_4204);
or U4618 (N_4618,N_4327,N_4255);
nand U4619 (N_4619,N_4323,N_4106);
nand U4620 (N_4620,N_4424,N_4426);
nor U4621 (N_4621,N_4108,N_4340);
nor U4622 (N_4622,N_4459,N_4476);
nor U4623 (N_4623,N_4247,N_4289);
nand U4624 (N_4624,N_4231,N_4495);
or U4625 (N_4625,N_4097,N_4309);
and U4626 (N_4626,N_4355,N_4248);
and U4627 (N_4627,N_4167,N_4027);
nand U4628 (N_4628,N_4467,N_4274);
nor U4629 (N_4629,N_4279,N_4093);
or U4630 (N_4630,N_4305,N_4332);
or U4631 (N_4631,N_4363,N_4346);
or U4632 (N_4632,N_4088,N_4315);
nand U4633 (N_4633,N_4159,N_4430);
or U4634 (N_4634,N_4071,N_4016);
or U4635 (N_4635,N_4110,N_4145);
nand U4636 (N_4636,N_4012,N_4107);
and U4637 (N_4637,N_4259,N_4367);
nor U4638 (N_4638,N_4072,N_4382);
xnor U4639 (N_4639,N_4215,N_4425);
and U4640 (N_4640,N_4083,N_4098);
nand U4641 (N_4641,N_4393,N_4273);
nor U4642 (N_4642,N_4392,N_4359);
and U4643 (N_4643,N_4466,N_4191);
and U4644 (N_4644,N_4019,N_4267);
xor U4645 (N_4645,N_4390,N_4474);
nor U4646 (N_4646,N_4099,N_4253);
xnor U4647 (N_4647,N_4038,N_4341);
nand U4648 (N_4648,N_4362,N_4460);
or U4649 (N_4649,N_4498,N_4490);
and U4650 (N_4650,N_4221,N_4330);
and U4651 (N_4651,N_4300,N_4372);
xor U4652 (N_4652,N_4000,N_4379);
and U4653 (N_4653,N_4422,N_4353);
nor U4654 (N_4654,N_4186,N_4360);
or U4655 (N_4655,N_4181,N_4203);
or U4656 (N_4656,N_4416,N_4176);
or U4657 (N_4657,N_4389,N_4417);
and U4658 (N_4658,N_4455,N_4358);
and U4659 (N_4659,N_4236,N_4115);
or U4660 (N_4660,N_4450,N_4100);
and U4661 (N_4661,N_4272,N_4473);
nor U4662 (N_4662,N_4092,N_4199);
nor U4663 (N_4663,N_4152,N_4067);
nand U4664 (N_4664,N_4368,N_4400);
nor U4665 (N_4665,N_4280,N_4243);
nor U4666 (N_4666,N_4006,N_4338);
and U4667 (N_4667,N_4044,N_4310);
and U4668 (N_4668,N_4276,N_4185);
nand U4669 (N_4669,N_4361,N_4381);
or U4670 (N_4670,N_4223,N_4369);
nor U4671 (N_4671,N_4117,N_4234);
nor U4672 (N_4672,N_4010,N_4321);
xnor U4673 (N_4673,N_4413,N_4308);
or U4674 (N_4674,N_4195,N_4246);
nand U4675 (N_4675,N_4096,N_4264);
or U4676 (N_4676,N_4042,N_4079);
and U4677 (N_4677,N_4468,N_4026);
nand U4678 (N_4678,N_4487,N_4166);
and U4679 (N_4679,N_4375,N_4240);
and U4680 (N_4680,N_4094,N_4402);
xnor U4681 (N_4681,N_4211,N_4051);
or U4682 (N_4682,N_4403,N_4227);
nor U4683 (N_4683,N_4219,N_4271);
and U4684 (N_4684,N_4101,N_4029);
and U4685 (N_4685,N_4109,N_4068);
nand U4686 (N_4686,N_4082,N_4275);
nand U4687 (N_4687,N_4035,N_4472);
xnor U4688 (N_4688,N_4089,N_4292);
or U4689 (N_4689,N_4126,N_4475);
nand U4690 (N_4690,N_4172,N_4206);
nand U4691 (N_4691,N_4343,N_4268);
and U4692 (N_4692,N_4454,N_4020);
nor U4693 (N_4693,N_4116,N_4281);
or U4694 (N_4694,N_4090,N_4299);
or U4695 (N_4695,N_4446,N_4160);
or U4696 (N_4696,N_4269,N_4444);
or U4697 (N_4697,N_4151,N_4419);
nand U4698 (N_4698,N_4144,N_4034);
or U4699 (N_4699,N_4373,N_4081);
or U4700 (N_4700,N_4303,N_4316);
or U4701 (N_4701,N_4131,N_4224);
nand U4702 (N_4702,N_4397,N_4439);
nor U4703 (N_4703,N_4222,N_4241);
or U4704 (N_4704,N_4119,N_4235);
and U4705 (N_4705,N_4156,N_4262);
and U4706 (N_4706,N_4285,N_4427);
xnor U4707 (N_4707,N_4233,N_4001);
or U4708 (N_4708,N_4043,N_4250);
nand U4709 (N_4709,N_4351,N_4229);
and U4710 (N_4710,N_4171,N_4055);
nor U4711 (N_4711,N_4208,N_4146);
or U4712 (N_4712,N_4329,N_4073);
xor U4713 (N_4713,N_4415,N_4118);
and U4714 (N_4714,N_4178,N_4209);
nor U4715 (N_4715,N_4258,N_4137);
and U4716 (N_4716,N_4356,N_4225);
and U4717 (N_4717,N_4414,N_4133);
xor U4718 (N_4718,N_4141,N_4254);
nand U4719 (N_4719,N_4295,N_4059);
nor U4720 (N_4720,N_4469,N_4205);
nor U4721 (N_4721,N_4411,N_4104);
and U4722 (N_4722,N_4288,N_4134);
and U4723 (N_4723,N_4457,N_4052);
and U4724 (N_4724,N_4489,N_4007);
nor U4725 (N_4725,N_4009,N_4399);
and U4726 (N_4726,N_4318,N_4154);
nor U4727 (N_4727,N_4437,N_4065);
nor U4728 (N_4728,N_4028,N_4237);
or U4729 (N_4729,N_4114,N_4477);
nand U4730 (N_4730,N_4091,N_4265);
and U4731 (N_4731,N_4252,N_4087);
nor U4732 (N_4732,N_4290,N_4105);
nor U4733 (N_4733,N_4481,N_4037);
nor U4734 (N_4734,N_4142,N_4187);
and U4735 (N_4735,N_4442,N_4491);
or U4736 (N_4736,N_4282,N_4024);
xor U4737 (N_4737,N_4453,N_4201);
and U4738 (N_4738,N_4086,N_4339);
nand U4739 (N_4739,N_4433,N_4095);
or U4740 (N_4740,N_4047,N_4447);
or U4741 (N_4741,N_4015,N_4121);
nor U4742 (N_4742,N_4488,N_4384);
and U4743 (N_4743,N_4461,N_4306);
or U4744 (N_4744,N_4277,N_4435);
nand U4745 (N_4745,N_4135,N_4163);
and U4746 (N_4746,N_4011,N_4004);
nor U4747 (N_4747,N_4296,N_4377);
or U4748 (N_4748,N_4408,N_4127);
or U4749 (N_4749,N_4128,N_4080);
nand U4750 (N_4750,N_4007,N_4114);
nor U4751 (N_4751,N_4421,N_4489);
xnor U4752 (N_4752,N_4083,N_4075);
nand U4753 (N_4753,N_4227,N_4429);
or U4754 (N_4754,N_4203,N_4160);
or U4755 (N_4755,N_4150,N_4052);
xnor U4756 (N_4756,N_4362,N_4405);
or U4757 (N_4757,N_4097,N_4110);
and U4758 (N_4758,N_4057,N_4468);
nor U4759 (N_4759,N_4445,N_4191);
or U4760 (N_4760,N_4100,N_4072);
nand U4761 (N_4761,N_4072,N_4289);
or U4762 (N_4762,N_4054,N_4281);
and U4763 (N_4763,N_4125,N_4061);
and U4764 (N_4764,N_4465,N_4298);
and U4765 (N_4765,N_4069,N_4163);
nand U4766 (N_4766,N_4338,N_4305);
nor U4767 (N_4767,N_4088,N_4094);
and U4768 (N_4768,N_4451,N_4358);
nor U4769 (N_4769,N_4331,N_4162);
nor U4770 (N_4770,N_4256,N_4348);
nand U4771 (N_4771,N_4126,N_4450);
nand U4772 (N_4772,N_4252,N_4260);
nor U4773 (N_4773,N_4335,N_4253);
or U4774 (N_4774,N_4113,N_4145);
nor U4775 (N_4775,N_4256,N_4205);
and U4776 (N_4776,N_4261,N_4016);
or U4777 (N_4777,N_4144,N_4278);
and U4778 (N_4778,N_4173,N_4127);
and U4779 (N_4779,N_4164,N_4293);
and U4780 (N_4780,N_4497,N_4165);
or U4781 (N_4781,N_4151,N_4184);
nand U4782 (N_4782,N_4473,N_4315);
nor U4783 (N_4783,N_4182,N_4140);
nand U4784 (N_4784,N_4452,N_4357);
nor U4785 (N_4785,N_4385,N_4396);
or U4786 (N_4786,N_4293,N_4046);
or U4787 (N_4787,N_4358,N_4045);
xnor U4788 (N_4788,N_4419,N_4202);
nor U4789 (N_4789,N_4029,N_4420);
nor U4790 (N_4790,N_4134,N_4173);
or U4791 (N_4791,N_4233,N_4029);
xnor U4792 (N_4792,N_4165,N_4235);
nand U4793 (N_4793,N_4351,N_4437);
and U4794 (N_4794,N_4010,N_4107);
nor U4795 (N_4795,N_4119,N_4150);
or U4796 (N_4796,N_4342,N_4298);
nor U4797 (N_4797,N_4045,N_4297);
or U4798 (N_4798,N_4083,N_4031);
or U4799 (N_4799,N_4264,N_4294);
nand U4800 (N_4800,N_4289,N_4357);
nand U4801 (N_4801,N_4173,N_4477);
and U4802 (N_4802,N_4419,N_4111);
nand U4803 (N_4803,N_4428,N_4327);
xor U4804 (N_4804,N_4136,N_4304);
and U4805 (N_4805,N_4321,N_4057);
xor U4806 (N_4806,N_4316,N_4024);
and U4807 (N_4807,N_4344,N_4375);
nand U4808 (N_4808,N_4145,N_4336);
and U4809 (N_4809,N_4472,N_4253);
nor U4810 (N_4810,N_4203,N_4271);
or U4811 (N_4811,N_4062,N_4257);
nor U4812 (N_4812,N_4237,N_4329);
nor U4813 (N_4813,N_4359,N_4366);
or U4814 (N_4814,N_4444,N_4227);
or U4815 (N_4815,N_4298,N_4300);
and U4816 (N_4816,N_4061,N_4299);
and U4817 (N_4817,N_4265,N_4067);
nor U4818 (N_4818,N_4446,N_4010);
nor U4819 (N_4819,N_4085,N_4326);
nand U4820 (N_4820,N_4286,N_4351);
nand U4821 (N_4821,N_4130,N_4172);
nand U4822 (N_4822,N_4310,N_4164);
or U4823 (N_4823,N_4343,N_4163);
or U4824 (N_4824,N_4355,N_4030);
and U4825 (N_4825,N_4234,N_4113);
and U4826 (N_4826,N_4036,N_4172);
or U4827 (N_4827,N_4248,N_4440);
or U4828 (N_4828,N_4485,N_4097);
xnor U4829 (N_4829,N_4022,N_4103);
and U4830 (N_4830,N_4350,N_4148);
nor U4831 (N_4831,N_4424,N_4454);
or U4832 (N_4832,N_4201,N_4109);
or U4833 (N_4833,N_4042,N_4394);
or U4834 (N_4834,N_4362,N_4366);
xnor U4835 (N_4835,N_4423,N_4091);
and U4836 (N_4836,N_4385,N_4268);
nand U4837 (N_4837,N_4225,N_4234);
xor U4838 (N_4838,N_4132,N_4171);
and U4839 (N_4839,N_4498,N_4441);
or U4840 (N_4840,N_4200,N_4439);
nand U4841 (N_4841,N_4001,N_4377);
nand U4842 (N_4842,N_4201,N_4358);
and U4843 (N_4843,N_4269,N_4487);
nand U4844 (N_4844,N_4084,N_4019);
nor U4845 (N_4845,N_4110,N_4236);
or U4846 (N_4846,N_4321,N_4319);
and U4847 (N_4847,N_4057,N_4357);
and U4848 (N_4848,N_4153,N_4269);
and U4849 (N_4849,N_4064,N_4097);
and U4850 (N_4850,N_4100,N_4345);
xnor U4851 (N_4851,N_4170,N_4496);
or U4852 (N_4852,N_4065,N_4483);
and U4853 (N_4853,N_4239,N_4134);
nand U4854 (N_4854,N_4439,N_4294);
and U4855 (N_4855,N_4239,N_4065);
nand U4856 (N_4856,N_4234,N_4278);
nor U4857 (N_4857,N_4311,N_4196);
xnor U4858 (N_4858,N_4311,N_4131);
nor U4859 (N_4859,N_4451,N_4379);
nor U4860 (N_4860,N_4416,N_4139);
and U4861 (N_4861,N_4163,N_4057);
nand U4862 (N_4862,N_4454,N_4358);
or U4863 (N_4863,N_4211,N_4490);
and U4864 (N_4864,N_4082,N_4030);
nor U4865 (N_4865,N_4034,N_4197);
and U4866 (N_4866,N_4174,N_4360);
or U4867 (N_4867,N_4403,N_4050);
or U4868 (N_4868,N_4170,N_4442);
nand U4869 (N_4869,N_4425,N_4213);
or U4870 (N_4870,N_4100,N_4465);
or U4871 (N_4871,N_4366,N_4086);
xnor U4872 (N_4872,N_4386,N_4145);
nor U4873 (N_4873,N_4417,N_4465);
or U4874 (N_4874,N_4006,N_4027);
nand U4875 (N_4875,N_4057,N_4150);
nand U4876 (N_4876,N_4184,N_4446);
nand U4877 (N_4877,N_4197,N_4249);
nor U4878 (N_4878,N_4279,N_4260);
xnor U4879 (N_4879,N_4124,N_4487);
or U4880 (N_4880,N_4024,N_4289);
or U4881 (N_4881,N_4387,N_4247);
nand U4882 (N_4882,N_4249,N_4168);
nand U4883 (N_4883,N_4008,N_4432);
and U4884 (N_4884,N_4142,N_4340);
nor U4885 (N_4885,N_4174,N_4096);
or U4886 (N_4886,N_4142,N_4366);
and U4887 (N_4887,N_4286,N_4292);
xnor U4888 (N_4888,N_4278,N_4050);
or U4889 (N_4889,N_4476,N_4160);
and U4890 (N_4890,N_4098,N_4200);
nor U4891 (N_4891,N_4499,N_4087);
and U4892 (N_4892,N_4051,N_4141);
and U4893 (N_4893,N_4157,N_4248);
and U4894 (N_4894,N_4282,N_4109);
nor U4895 (N_4895,N_4161,N_4457);
or U4896 (N_4896,N_4147,N_4069);
nor U4897 (N_4897,N_4355,N_4338);
nor U4898 (N_4898,N_4442,N_4212);
nand U4899 (N_4899,N_4255,N_4190);
nor U4900 (N_4900,N_4273,N_4191);
xnor U4901 (N_4901,N_4113,N_4142);
and U4902 (N_4902,N_4000,N_4082);
or U4903 (N_4903,N_4028,N_4097);
or U4904 (N_4904,N_4041,N_4310);
nand U4905 (N_4905,N_4155,N_4211);
nor U4906 (N_4906,N_4226,N_4198);
or U4907 (N_4907,N_4472,N_4034);
or U4908 (N_4908,N_4146,N_4075);
and U4909 (N_4909,N_4059,N_4266);
or U4910 (N_4910,N_4152,N_4063);
xnor U4911 (N_4911,N_4460,N_4221);
and U4912 (N_4912,N_4485,N_4297);
or U4913 (N_4913,N_4049,N_4477);
nand U4914 (N_4914,N_4031,N_4466);
nor U4915 (N_4915,N_4092,N_4088);
nor U4916 (N_4916,N_4156,N_4471);
and U4917 (N_4917,N_4365,N_4018);
nor U4918 (N_4918,N_4251,N_4174);
nand U4919 (N_4919,N_4351,N_4340);
nor U4920 (N_4920,N_4098,N_4108);
nor U4921 (N_4921,N_4051,N_4025);
and U4922 (N_4922,N_4082,N_4167);
and U4923 (N_4923,N_4437,N_4128);
xor U4924 (N_4924,N_4260,N_4144);
or U4925 (N_4925,N_4143,N_4043);
or U4926 (N_4926,N_4472,N_4146);
or U4927 (N_4927,N_4223,N_4323);
nand U4928 (N_4928,N_4037,N_4237);
nor U4929 (N_4929,N_4100,N_4294);
or U4930 (N_4930,N_4413,N_4206);
nor U4931 (N_4931,N_4055,N_4095);
and U4932 (N_4932,N_4077,N_4363);
nand U4933 (N_4933,N_4245,N_4120);
nor U4934 (N_4934,N_4111,N_4431);
nand U4935 (N_4935,N_4133,N_4365);
and U4936 (N_4936,N_4057,N_4452);
nand U4937 (N_4937,N_4015,N_4475);
nand U4938 (N_4938,N_4041,N_4446);
nand U4939 (N_4939,N_4459,N_4153);
nand U4940 (N_4940,N_4219,N_4016);
nor U4941 (N_4941,N_4261,N_4482);
nor U4942 (N_4942,N_4063,N_4089);
and U4943 (N_4943,N_4198,N_4070);
nand U4944 (N_4944,N_4413,N_4496);
nand U4945 (N_4945,N_4207,N_4260);
and U4946 (N_4946,N_4152,N_4078);
or U4947 (N_4947,N_4305,N_4493);
or U4948 (N_4948,N_4324,N_4483);
nand U4949 (N_4949,N_4258,N_4064);
nand U4950 (N_4950,N_4287,N_4156);
nor U4951 (N_4951,N_4152,N_4449);
and U4952 (N_4952,N_4335,N_4409);
nor U4953 (N_4953,N_4264,N_4017);
and U4954 (N_4954,N_4078,N_4262);
xor U4955 (N_4955,N_4490,N_4492);
and U4956 (N_4956,N_4159,N_4443);
nor U4957 (N_4957,N_4392,N_4279);
nor U4958 (N_4958,N_4440,N_4095);
nor U4959 (N_4959,N_4206,N_4400);
nor U4960 (N_4960,N_4102,N_4096);
xnor U4961 (N_4961,N_4326,N_4088);
nand U4962 (N_4962,N_4165,N_4290);
nand U4963 (N_4963,N_4203,N_4432);
or U4964 (N_4964,N_4484,N_4006);
nor U4965 (N_4965,N_4016,N_4278);
or U4966 (N_4966,N_4306,N_4333);
nand U4967 (N_4967,N_4366,N_4239);
and U4968 (N_4968,N_4480,N_4400);
or U4969 (N_4969,N_4384,N_4207);
and U4970 (N_4970,N_4182,N_4442);
nand U4971 (N_4971,N_4217,N_4286);
nand U4972 (N_4972,N_4112,N_4402);
and U4973 (N_4973,N_4022,N_4237);
and U4974 (N_4974,N_4283,N_4203);
nand U4975 (N_4975,N_4455,N_4074);
xnor U4976 (N_4976,N_4250,N_4408);
or U4977 (N_4977,N_4385,N_4236);
or U4978 (N_4978,N_4311,N_4222);
nand U4979 (N_4979,N_4193,N_4078);
or U4980 (N_4980,N_4163,N_4488);
nand U4981 (N_4981,N_4303,N_4291);
or U4982 (N_4982,N_4308,N_4442);
nor U4983 (N_4983,N_4028,N_4321);
nand U4984 (N_4984,N_4483,N_4209);
nand U4985 (N_4985,N_4085,N_4285);
nor U4986 (N_4986,N_4418,N_4119);
and U4987 (N_4987,N_4235,N_4238);
and U4988 (N_4988,N_4039,N_4432);
nor U4989 (N_4989,N_4179,N_4039);
and U4990 (N_4990,N_4361,N_4215);
or U4991 (N_4991,N_4353,N_4000);
or U4992 (N_4992,N_4002,N_4291);
or U4993 (N_4993,N_4476,N_4217);
nor U4994 (N_4994,N_4245,N_4055);
nand U4995 (N_4995,N_4374,N_4043);
nand U4996 (N_4996,N_4413,N_4236);
or U4997 (N_4997,N_4243,N_4246);
nor U4998 (N_4998,N_4104,N_4210);
nor U4999 (N_4999,N_4035,N_4439);
or U5000 (N_5000,N_4926,N_4930);
or U5001 (N_5001,N_4935,N_4957);
nand U5002 (N_5002,N_4985,N_4651);
or U5003 (N_5003,N_4510,N_4916);
nor U5004 (N_5004,N_4839,N_4641);
or U5005 (N_5005,N_4553,N_4749);
xnor U5006 (N_5006,N_4689,N_4673);
nor U5007 (N_5007,N_4722,N_4789);
or U5008 (N_5008,N_4794,N_4950);
xor U5009 (N_5009,N_4921,N_4909);
nand U5010 (N_5010,N_4569,N_4831);
nand U5011 (N_5011,N_4773,N_4680);
or U5012 (N_5012,N_4638,N_4948);
and U5013 (N_5013,N_4523,N_4843);
nor U5014 (N_5014,N_4715,N_4650);
or U5015 (N_5015,N_4645,N_4898);
or U5016 (N_5016,N_4941,N_4819);
xor U5017 (N_5017,N_4601,N_4859);
xnor U5018 (N_5018,N_4772,N_4817);
and U5019 (N_5019,N_4706,N_4575);
xor U5020 (N_5020,N_4590,N_4549);
or U5021 (N_5021,N_4894,N_4571);
or U5022 (N_5022,N_4633,N_4765);
nor U5023 (N_5023,N_4559,N_4649);
and U5024 (N_5024,N_4798,N_4602);
and U5025 (N_5025,N_4723,N_4864);
nor U5026 (N_5026,N_4812,N_4613);
and U5027 (N_5027,N_4937,N_4530);
xor U5028 (N_5028,N_4529,N_4932);
nand U5029 (N_5029,N_4825,N_4534);
and U5030 (N_5030,N_4628,N_4768);
or U5031 (N_5031,N_4755,N_4629);
nor U5032 (N_5032,N_4631,N_4929);
nor U5033 (N_5033,N_4877,N_4588);
nand U5034 (N_5034,N_4848,N_4987);
xnor U5035 (N_5035,N_4992,N_4885);
or U5036 (N_5036,N_4933,N_4584);
nor U5037 (N_5037,N_4993,N_4668);
xor U5038 (N_5038,N_4873,N_4657);
or U5039 (N_5039,N_4835,N_4964);
nand U5040 (N_5040,N_4671,N_4536);
xor U5041 (N_5041,N_4805,N_4740);
nor U5042 (N_5042,N_4544,N_4648);
nand U5043 (N_5043,N_4676,N_4797);
or U5044 (N_5044,N_4558,N_4607);
nor U5045 (N_5045,N_4672,N_4999);
nand U5046 (N_5046,N_4736,N_4770);
or U5047 (N_5047,N_4745,N_4983);
and U5048 (N_5048,N_4900,N_4524);
and U5049 (N_5049,N_4617,N_4512);
or U5050 (N_5050,N_4750,N_4681);
nand U5051 (N_5051,N_4783,N_4764);
or U5052 (N_5052,N_4686,N_4568);
nand U5053 (N_5053,N_4838,N_4832);
nand U5054 (N_5054,N_4920,N_4962);
or U5055 (N_5055,N_4662,N_4517);
nand U5056 (N_5056,N_4531,N_4579);
or U5057 (N_5057,N_4971,N_4827);
nand U5058 (N_5058,N_4989,N_4542);
nand U5059 (N_5059,N_4868,N_4829);
nand U5060 (N_5060,N_4847,N_4753);
or U5061 (N_5061,N_4997,N_4806);
and U5062 (N_5062,N_4842,N_4702);
nand U5063 (N_5063,N_4612,N_4578);
and U5064 (N_5064,N_4924,N_4786);
xnor U5065 (N_5065,N_4796,N_4952);
nand U5066 (N_5066,N_4851,N_4775);
and U5067 (N_5067,N_4860,N_4988);
or U5068 (N_5068,N_4659,N_4562);
or U5069 (N_5069,N_4748,N_4514);
nor U5070 (N_5070,N_4508,N_4743);
nand U5071 (N_5071,N_4866,N_4876);
and U5072 (N_5072,N_4897,N_4756);
nor U5073 (N_5073,N_4778,N_4721);
nand U5074 (N_5074,N_4608,N_4734);
xor U5075 (N_5075,N_4513,N_4966);
and U5076 (N_5076,N_4521,N_4511);
nand U5077 (N_5077,N_4582,N_4986);
nor U5078 (N_5078,N_4587,N_4803);
or U5079 (N_5079,N_4954,N_4888);
nor U5080 (N_5080,N_4914,N_4967);
nor U5081 (N_5081,N_4846,N_4718);
xor U5082 (N_5082,N_4507,N_4527);
xnor U5083 (N_5083,N_4733,N_4807);
nor U5084 (N_5084,N_4515,N_4732);
and U5085 (N_5085,N_4639,N_4901);
and U5086 (N_5086,N_4543,N_4801);
nand U5087 (N_5087,N_4624,N_4746);
nor U5088 (N_5088,N_4593,N_4737);
or U5089 (N_5089,N_4946,N_4960);
nor U5090 (N_5090,N_4959,N_4574);
xor U5091 (N_5091,N_4698,N_4991);
or U5092 (N_5092,N_4965,N_4632);
nand U5093 (N_5093,N_4580,N_4961);
and U5094 (N_5094,N_4573,N_4713);
and U5095 (N_5095,N_4699,N_4912);
or U5096 (N_5096,N_4939,N_4881);
and U5097 (N_5097,N_4707,N_4548);
nor U5098 (N_5098,N_4928,N_4841);
nand U5099 (N_5099,N_4795,N_4857);
and U5100 (N_5100,N_4940,N_4661);
xnor U5101 (N_5101,N_4793,N_4776);
xor U5102 (N_5102,N_4627,N_4654);
and U5103 (N_5103,N_4620,N_4904);
and U5104 (N_5104,N_4518,N_4554);
or U5105 (N_5105,N_4594,N_4758);
nor U5106 (N_5106,N_4762,N_4844);
nor U5107 (N_5107,N_4665,N_4906);
nor U5108 (N_5108,N_4836,N_4705);
xor U5109 (N_5109,N_4856,N_4977);
and U5110 (N_5110,N_4953,N_4934);
nand U5111 (N_5111,N_4799,N_4688);
nor U5112 (N_5112,N_4871,N_4730);
and U5113 (N_5113,N_4763,N_4727);
xnor U5114 (N_5114,N_4902,N_4643);
or U5115 (N_5115,N_4696,N_4863);
and U5116 (N_5116,N_4526,N_4927);
xnor U5117 (N_5117,N_4821,N_4867);
nor U5118 (N_5118,N_4609,N_4958);
or U5119 (N_5119,N_4996,N_4604);
nand U5120 (N_5120,N_4744,N_4973);
nor U5121 (N_5121,N_4576,N_4591);
or U5122 (N_5122,N_4923,N_4809);
or U5123 (N_5123,N_4760,N_4545);
nand U5124 (N_5124,N_4739,N_4840);
nor U5125 (N_5125,N_4896,N_4567);
nand U5126 (N_5126,N_4975,N_4931);
xor U5127 (N_5127,N_4815,N_4625);
xnor U5128 (N_5128,N_4982,N_4899);
or U5129 (N_5129,N_4994,N_4541);
or U5130 (N_5130,N_4626,N_4800);
nor U5131 (N_5131,N_4810,N_4656);
nor U5132 (N_5132,N_4535,N_4502);
xor U5133 (N_5133,N_4981,N_4879);
and U5134 (N_5134,N_4572,N_4826);
and U5135 (N_5135,N_4501,N_4943);
nand U5136 (N_5136,N_4540,N_4777);
nor U5137 (N_5137,N_4949,N_4837);
and U5138 (N_5138,N_4849,N_4589);
nand U5139 (N_5139,N_4915,N_4684);
nor U5140 (N_5140,N_4751,N_4556);
or U5141 (N_5141,N_4884,N_4664);
and U5142 (N_5142,N_4725,N_4972);
or U5143 (N_5143,N_4566,N_4917);
or U5144 (N_5144,N_4675,N_4710);
or U5145 (N_5145,N_4890,N_4603);
or U5146 (N_5146,N_4887,N_4979);
xnor U5147 (N_5147,N_4595,N_4895);
nand U5148 (N_5148,N_4854,N_4586);
nand U5149 (N_5149,N_4791,N_4822);
nand U5150 (N_5150,N_4532,N_4616);
nand U5151 (N_5151,N_4855,N_4630);
nand U5152 (N_5152,N_4984,N_4550);
and U5153 (N_5153,N_4944,N_4919);
nand U5154 (N_5154,N_4766,N_4911);
and U5155 (N_5155,N_4802,N_4634);
and U5156 (N_5156,N_4677,N_4581);
and U5157 (N_5157,N_4720,N_4500);
nor U5158 (N_5158,N_4539,N_4947);
and U5159 (N_5159,N_4889,N_4708);
and U5160 (N_5160,N_4853,N_4754);
nand U5161 (N_5161,N_4875,N_4956);
and U5162 (N_5162,N_4598,N_4828);
nor U5163 (N_5163,N_4728,N_4522);
nand U5164 (N_5164,N_4623,N_4907);
or U5165 (N_5165,N_4910,N_4606);
nand U5166 (N_5166,N_4731,N_4703);
or U5167 (N_5167,N_4872,N_4564);
or U5168 (N_5168,N_4874,N_4978);
nand U5169 (N_5169,N_4711,N_4729);
or U5170 (N_5170,N_4820,N_4850);
nand U5171 (N_5171,N_4998,N_4615);
and U5172 (N_5172,N_4974,N_4913);
nor U5173 (N_5173,N_4903,N_4714);
nor U5174 (N_5174,N_4716,N_4771);
and U5175 (N_5175,N_4834,N_4596);
and U5176 (N_5176,N_4642,N_4968);
or U5177 (N_5177,N_4779,N_4516);
nand U5178 (N_5178,N_4788,N_4726);
or U5179 (N_5179,N_4865,N_4666);
nand U5180 (N_5180,N_4878,N_4891);
nand U5181 (N_5181,N_4883,N_4787);
or U5182 (N_5182,N_4611,N_4552);
or U5183 (N_5183,N_4519,N_4683);
and U5184 (N_5184,N_4719,N_4570);
and U5185 (N_5185,N_4976,N_4538);
or U5186 (N_5186,N_4520,N_4690);
nor U5187 (N_5187,N_4980,N_4561);
or U5188 (N_5188,N_4674,N_4813);
nor U5189 (N_5189,N_4824,N_4785);
or U5190 (N_5190,N_4741,N_4942);
nand U5191 (N_5191,N_4685,N_4555);
or U5192 (N_5192,N_4970,N_4862);
and U5193 (N_5193,N_4660,N_4951);
nor U5194 (N_5194,N_4990,N_4945);
nand U5195 (N_5195,N_4635,N_4767);
nor U5196 (N_5196,N_4557,N_4599);
nand U5197 (N_5197,N_4742,N_4687);
and U5198 (N_5198,N_4506,N_4533);
nor U5199 (N_5199,N_4963,N_4780);
and U5200 (N_5200,N_4709,N_4636);
nor U5201 (N_5201,N_4852,N_4647);
xnor U5202 (N_5202,N_4644,N_4525);
xor U5203 (N_5203,N_4610,N_4892);
and U5204 (N_5204,N_4790,N_4908);
or U5205 (N_5205,N_4692,N_4869);
nand U5206 (N_5206,N_4936,N_4995);
and U5207 (N_5207,N_4693,N_4861);
nand U5208 (N_5208,N_4577,N_4547);
nand U5209 (N_5209,N_4747,N_4761);
nor U5210 (N_5210,N_4759,N_4667);
nand U5211 (N_5211,N_4804,N_4583);
and U5212 (N_5212,N_4505,N_4646);
and U5213 (N_5213,N_4735,N_4619);
nor U5214 (N_5214,N_4823,N_4653);
and U5215 (N_5215,N_4504,N_4528);
and U5216 (N_5216,N_4697,N_4622);
or U5217 (N_5217,N_4682,N_4774);
and U5218 (N_5218,N_4700,N_4605);
and U5219 (N_5219,N_4955,N_4679);
or U5220 (N_5220,N_4757,N_4565);
nand U5221 (N_5221,N_4925,N_4652);
nor U5222 (N_5222,N_4882,N_4585);
and U5223 (N_5223,N_4724,N_4814);
or U5224 (N_5224,N_4669,N_4922);
nor U5225 (N_5225,N_4870,N_4658);
or U5226 (N_5226,N_4738,N_4663);
nand U5227 (N_5227,N_4695,N_4551);
or U5228 (N_5228,N_4614,N_4691);
and U5229 (N_5229,N_4600,N_4592);
and U5230 (N_5230,N_4503,N_4655);
xnor U5231 (N_5231,N_4563,N_4969);
and U5232 (N_5232,N_4792,N_4537);
nor U5233 (N_5233,N_4811,N_4782);
nor U5234 (N_5234,N_4717,N_4712);
nor U5235 (N_5235,N_4678,N_4818);
or U5236 (N_5236,N_4905,N_4781);
or U5237 (N_5237,N_4784,N_4637);
xnor U5238 (N_5238,N_4880,N_4618);
and U5239 (N_5239,N_4816,N_4509);
and U5240 (N_5240,N_4858,N_4546);
or U5241 (N_5241,N_4830,N_4701);
or U5242 (N_5242,N_4808,N_4886);
nand U5243 (N_5243,N_4704,N_4597);
nand U5244 (N_5244,N_4752,N_4769);
or U5245 (N_5245,N_4845,N_4833);
and U5246 (N_5246,N_4918,N_4560);
and U5247 (N_5247,N_4640,N_4621);
nor U5248 (N_5248,N_4938,N_4694);
or U5249 (N_5249,N_4670,N_4893);
or U5250 (N_5250,N_4597,N_4817);
nor U5251 (N_5251,N_4654,N_4651);
or U5252 (N_5252,N_4593,N_4949);
and U5253 (N_5253,N_4628,N_4979);
or U5254 (N_5254,N_4753,N_4824);
xor U5255 (N_5255,N_4597,N_4554);
nand U5256 (N_5256,N_4980,N_4793);
or U5257 (N_5257,N_4896,N_4800);
nand U5258 (N_5258,N_4866,N_4661);
nor U5259 (N_5259,N_4526,N_4539);
nand U5260 (N_5260,N_4753,N_4965);
nor U5261 (N_5261,N_4906,N_4910);
nor U5262 (N_5262,N_4887,N_4834);
or U5263 (N_5263,N_4670,N_4963);
and U5264 (N_5264,N_4652,N_4521);
nor U5265 (N_5265,N_4750,N_4668);
and U5266 (N_5266,N_4868,N_4787);
nand U5267 (N_5267,N_4993,N_4780);
and U5268 (N_5268,N_4950,N_4585);
nor U5269 (N_5269,N_4659,N_4959);
or U5270 (N_5270,N_4813,N_4971);
or U5271 (N_5271,N_4791,N_4730);
or U5272 (N_5272,N_4765,N_4882);
nand U5273 (N_5273,N_4686,N_4779);
and U5274 (N_5274,N_4925,N_4976);
nor U5275 (N_5275,N_4992,N_4715);
nand U5276 (N_5276,N_4962,N_4793);
nand U5277 (N_5277,N_4778,N_4600);
nand U5278 (N_5278,N_4933,N_4958);
nor U5279 (N_5279,N_4804,N_4976);
nor U5280 (N_5280,N_4746,N_4627);
nor U5281 (N_5281,N_4515,N_4772);
nand U5282 (N_5282,N_4657,N_4668);
or U5283 (N_5283,N_4716,N_4815);
nand U5284 (N_5284,N_4642,N_4501);
nor U5285 (N_5285,N_4550,N_4533);
nand U5286 (N_5286,N_4973,N_4809);
xnor U5287 (N_5287,N_4846,N_4793);
or U5288 (N_5288,N_4719,N_4765);
nand U5289 (N_5289,N_4955,N_4534);
nand U5290 (N_5290,N_4979,N_4592);
nand U5291 (N_5291,N_4808,N_4983);
or U5292 (N_5292,N_4571,N_4759);
nor U5293 (N_5293,N_4554,N_4574);
nand U5294 (N_5294,N_4914,N_4658);
and U5295 (N_5295,N_4623,N_4994);
or U5296 (N_5296,N_4831,N_4554);
xor U5297 (N_5297,N_4836,N_4942);
or U5298 (N_5298,N_4723,N_4790);
xnor U5299 (N_5299,N_4927,N_4727);
or U5300 (N_5300,N_4895,N_4760);
nand U5301 (N_5301,N_4641,N_4506);
and U5302 (N_5302,N_4988,N_4508);
xnor U5303 (N_5303,N_4878,N_4651);
nand U5304 (N_5304,N_4921,N_4542);
and U5305 (N_5305,N_4695,N_4553);
xor U5306 (N_5306,N_4877,N_4712);
nand U5307 (N_5307,N_4680,N_4753);
or U5308 (N_5308,N_4642,N_4940);
or U5309 (N_5309,N_4546,N_4932);
nor U5310 (N_5310,N_4850,N_4846);
nand U5311 (N_5311,N_4543,N_4937);
and U5312 (N_5312,N_4824,N_4716);
or U5313 (N_5313,N_4939,N_4608);
nor U5314 (N_5314,N_4746,N_4893);
nor U5315 (N_5315,N_4996,N_4866);
nor U5316 (N_5316,N_4510,N_4695);
or U5317 (N_5317,N_4771,N_4974);
or U5318 (N_5318,N_4888,N_4774);
or U5319 (N_5319,N_4964,N_4597);
or U5320 (N_5320,N_4554,N_4887);
nand U5321 (N_5321,N_4742,N_4559);
nor U5322 (N_5322,N_4972,N_4621);
or U5323 (N_5323,N_4947,N_4508);
nand U5324 (N_5324,N_4601,N_4633);
nor U5325 (N_5325,N_4800,N_4560);
and U5326 (N_5326,N_4848,N_4893);
nor U5327 (N_5327,N_4746,N_4546);
nand U5328 (N_5328,N_4603,N_4820);
nand U5329 (N_5329,N_4589,N_4579);
and U5330 (N_5330,N_4582,N_4623);
nand U5331 (N_5331,N_4505,N_4556);
nor U5332 (N_5332,N_4619,N_4818);
and U5333 (N_5333,N_4572,N_4803);
or U5334 (N_5334,N_4975,N_4838);
nor U5335 (N_5335,N_4643,N_4548);
nor U5336 (N_5336,N_4801,N_4833);
nor U5337 (N_5337,N_4784,N_4653);
and U5338 (N_5338,N_4729,N_4587);
or U5339 (N_5339,N_4935,N_4894);
nor U5340 (N_5340,N_4842,N_4902);
nor U5341 (N_5341,N_4950,N_4686);
or U5342 (N_5342,N_4951,N_4917);
nor U5343 (N_5343,N_4741,N_4912);
nor U5344 (N_5344,N_4775,N_4652);
or U5345 (N_5345,N_4761,N_4568);
nand U5346 (N_5346,N_4757,N_4533);
and U5347 (N_5347,N_4598,N_4895);
or U5348 (N_5348,N_4948,N_4938);
nand U5349 (N_5349,N_4935,N_4999);
nand U5350 (N_5350,N_4609,N_4736);
nor U5351 (N_5351,N_4784,N_4699);
nor U5352 (N_5352,N_4719,N_4860);
and U5353 (N_5353,N_4557,N_4756);
or U5354 (N_5354,N_4641,N_4791);
nand U5355 (N_5355,N_4521,N_4504);
nor U5356 (N_5356,N_4724,N_4928);
nor U5357 (N_5357,N_4955,N_4969);
xor U5358 (N_5358,N_4913,N_4643);
nor U5359 (N_5359,N_4700,N_4735);
or U5360 (N_5360,N_4702,N_4528);
or U5361 (N_5361,N_4525,N_4970);
and U5362 (N_5362,N_4641,N_4920);
or U5363 (N_5363,N_4693,N_4515);
nand U5364 (N_5364,N_4618,N_4826);
nand U5365 (N_5365,N_4912,N_4725);
nor U5366 (N_5366,N_4980,N_4643);
and U5367 (N_5367,N_4856,N_4894);
nor U5368 (N_5368,N_4992,N_4520);
xnor U5369 (N_5369,N_4717,N_4510);
xor U5370 (N_5370,N_4529,N_4691);
nand U5371 (N_5371,N_4734,N_4622);
or U5372 (N_5372,N_4983,N_4684);
and U5373 (N_5373,N_4637,N_4529);
or U5374 (N_5374,N_4978,N_4838);
nand U5375 (N_5375,N_4587,N_4555);
nand U5376 (N_5376,N_4677,N_4560);
or U5377 (N_5377,N_4813,N_4810);
or U5378 (N_5378,N_4932,N_4708);
and U5379 (N_5379,N_4753,N_4895);
or U5380 (N_5380,N_4750,N_4954);
and U5381 (N_5381,N_4531,N_4944);
or U5382 (N_5382,N_4843,N_4562);
nand U5383 (N_5383,N_4568,N_4730);
nor U5384 (N_5384,N_4626,N_4873);
or U5385 (N_5385,N_4792,N_4947);
nand U5386 (N_5386,N_4529,N_4976);
and U5387 (N_5387,N_4700,N_4964);
nor U5388 (N_5388,N_4952,N_4784);
and U5389 (N_5389,N_4533,N_4728);
xor U5390 (N_5390,N_4846,N_4773);
nor U5391 (N_5391,N_4923,N_4893);
or U5392 (N_5392,N_4639,N_4969);
nor U5393 (N_5393,N_4588,N_4993);
nor U5394 (N_5394,N_4720,N_4734);
nand U5395 (N_5395,N_4841,N_4929);
or U5396 (N_5396,N_4758,N_4831);
or U5397 (N_5397,N_4693,N_4632);
and U5398 (N_5398,N_4637,N_4717);
nor U5399 (N_5399,N_4925,N_4759);
xor U5400 (N_5400,N_4888,N_4628);
xor U5401 (N_5401,N_4942,N_4689);
or U5402 (N_5402,N_4825,N_4565);
and U5403 (N_5403,N_4800,N_4961);
or U5404 (N_5404,N_4975,N_4938);
and U5405 (N_5405,N_4968,N_4897);
nand U5406 (N_5406,N_4882,N_4847);
or U5407 (N_5407,N_4571,N_4732);
or U5408 (N_5408,N_4589,N_4732);
or U5409 (N_5409,N_4786,N_4990);
or U5410 (N_5410,N_4588,N_4733);
nand U5411 (N_5411,N_4833,N_4977);
nor U5412 (N_5412,N_4964,N_4963);
or U5413 (N_5413,N_4795,N_4906);
nor U5414 (N_5414,N_4892,N_4947);
or U5415 (N_5415,N_4636,N_4997);
or U5416 (N_5416,N_4733,N_4821);
nand U5417 (N_5417,N_4872,N_4688);
and U5418 (N_5418,N_4683,N_4902);
nand U5419 (N_5419,N_4630,N_4632);
nor U5420 (N_5420,N_4724,N_4613);
and U5421 (N_5421,N_4657,N_4792);
nor U5422 (N_5422,N_4660,N_4866);
and U5423 (N_5423,N_4578,N_4609);
and U5424 (N_5424,N_4936,N_4958);
and U5425 (N_5425,N_4578,N_4981);
nand U5426 (N_5426,N_4971,N_4733);
and U5427 (N_5427,N_4583,N_4523);
or U5428 (N_5428,N_4753,N_4897);
nand U5429 (N_5429,N_4691,N_4829);
and U5430 (N_5430,N_4994,N_4883);
or U5431 (N_5431,N_4859,N_4584);
nand U5432 (N_5432,N_4929,N_4963);
nor U5433 (N_5433,N_4505,N_4753);
nand U5434 (N_5434,N_4882,N_4551);
and U5435 (N_5435,N_4920,N_4931);
nor U5436 (N_5436,N_4839,N_4562);
nor U5437 (N_5437,N_4547,N_4764);
nor U5438 (N_5438,N_4749,N_4614);
and U5439 (N_5439,N_4551,N_4766);
nand U5440 (N_5440,N_4500,N_4659);
and U5441 (N_5441,N_4694,N_4611);
nor U5442 (N_5442,N_4764,N_4817);
nor U5443 (N_5443,N_4713,N_4917);
and U5444 (N_5444,N_4671,N_4795);
nor U5445 (N_5445,N_4778,N_4801);
nor U5446 (N_5446,N_4957,N_4692);
or U5447 (N_5447,N_4651,N_4871);
or U5448 (N_5448,N_4890,N_4651);
or U5449 (N_5449,N_4821,N_4916);
and U5450 (N_5450,N_4640,N_4677);
nand U5451 (N_5451,N_4518,N_4534);
nand U5452 (N_5452,N_4673,N_4979);
nor U5453 (N_5453,N_4505,N_4954);
and U5454 (N_5454,N_4714,N_4958);
or U5455 (N_5455,N_4963,N_4507);
nor U5456 (N_5456,N_4594,N_4626);
nor U5457 (N_5457,N_4579,N_4841);
or U5458 (N_5458,N_4866,N_4513);
or U5459 (N_5459,N_4990,N_4804);
nand U5460 (N_5460,N_4550,N_4514);
and U5461 (N_5461,N_4612,N_4964);
nor U5462 (N_5462,N_4779,N_4604);
nor U5463 (N_5463,N_4799,N_4919);
nand U5464 (N_5464,N_4711,N_4772);
and U5465 (N_5465,N_4899,N_4782);
or U5466 (N_5466,N_4575,N_4778);
or U5467 (N_5467,N_4561,N_4602);
and U5468 (N_5468,N_4656,N_4860);
or U5469 (N_5469,N_4713,N_4843);
or U5470 (N_5470,N_4792,N_4963);
xor U5471 (N_5471,N_4567,N_4947);
xor U5472 (N_5472,N_4523,N_4891);
nor U5473 (N_5473,N_4547,N_4826);
xor U5474 (N_5474,N_4999,N_4864);
and U5475 (N_5475,N_4706,N_4642);
nand U5476 (N_5476,N_4745,N_4696);
nor U5477 (N_5477,N_4684,N_4862);
xor U5478 (N_5478,N_4618,N_4789);
or U5479 (N_5479,N_4882,N_4947);
nand U5480 (N_5480,N_4850,N_4771);
and U5481 (N_5481,N_4807,N_4567);
nand U5482 (N_5482,N_4531,N_4898);
nor U5483 (N_5483,N_4970,N_4588);
nand U5484 (N_5484,N_4824,N_4673);
nand U5485 (N_5485,N_4863,N_4551);
or U5486 (N_5486,N_4799,N_4983);
nand U5487 (N_5487,N_4721,N_4801);
nor U5488 (N_5488,N_4995,N_4767);
and U5489 (N_5489,N_4993,N_4829);
nor U5490 (N_5490,N_4748,N_4897);
or U5491 (N_5491,N_4951,N_4676);
nor U5492 (N_5492,N_4649,N_4524);
or U5493 (N_5493,N_4868,N_4959);
and U5494 (N_5494,N_4635,N_4736);
and U5495 (N_5495,N_4964,N_4836);
xor U5496 (N_5496,N_4916,N_4524);
and U5497 (N_5497,N_4931,N_4576);
and U5498 (N_5498,N_4930,N_4864);
and U5499 (N_5499,N_4584,N_4583);
nor U5500 (N_5500,N_5421,N_5474);
or U5501 (N_5501,N_5483,N_5326);
and U5502 (N_5502,N_5296,N_5202);
nand U5503 (N_5503,N_5079,N_5220);
nand U5504 (N_5504,N_5117,N_5283);
xnor U5505 (N_5505,N_5178,N_5052);
and U5506 (N_5506,N_5103,N_5418);
nor U5507 (N_5507,N_5351,N_5349);
nand U5508 (N_5508,N_5286,N_5200);
or U5509 (N_5509,N_5437,N_5243);
nor U5510 (N_5510,N_5392,N_5261);
and U5511 (N_5511,N_5191,N_5016);
and U5512 (N_5512,N_5284,N_5354);
and U5513 (N_5513,N_5025,N_5409);
xor U5514 (N_5514,N_5106,N_5299);
or U5515 (N_5515,N_5438,N_5030);
or U5516 (N_5516,N_5318,N_5381);
nand U5517 (N_5517,N_5213,N_5441);
xor U5518 (N_5518,N_5021,N_5221);
nor U5519 (N_5519,N_5132,N_5336);
nand U5520 (N_5520,N_5301,N_5471);
nand U5521 (N_5521,N_5176,N_5477);
and U5522 (N_5522,N_5434,N_5164);
nand U5523 (N_5523,N_5264,N_5179);
nor U5524 (N_5524,N_5001,N_5169);
or U5525 (N_5525,N_5153,N_5435);
or U5526 (N_5526,N_5156,N_5250);
or U5527 (N_5527,N_5259,N_5494);
or U5528 (N_5528,N_5073,N_5090);
or U5529 (N_5529,N_5372,N_5230);
xnor U5530 (N_5530,N_5212,N_5334);
nor U5531 (N_5531,N_5249,N_5024);
or U5532 (N_5532,N_5088,N_5094);
nor U5533 (N_5533,N_5187,N_5246);
nand U5534 (N_5534,N_5029,N_5274);
and U5535 (N_5535,N_5379,N_5214);
or U5536 (N_5536,N_5330,N_5129);
nor U5537 (N_5537,N_5462,N_5035);
or U5538 (N_5538,N_5444,N_5498);
xnor U5539 (N_5539,N_5255,N_5127);
xor U5540 (N_5540,N_5415,N_5161);
nand U5541 (N_5541,N_5452,N_5321);
xor U5542 (N_5542,N_5171,N_5057);
nand U5543 (N_5543,N_5064,N_5124);
nor U5544 (N_5544,N_5279,N_5219);
nor U5545 (N_5545,N_5263,N_5428);
or U5546 (N_5546,N_5065,N_5130);
and U5547 (N_5547,N_5458,N_5207);
xor U5548 (N_5548,N_5196,N_5155);
nor U5549 (N_5549,N_5235,N_5059);
and U5550 (N_5550,N_5363,N_5037);
and U5551 (N_5551,N_5137,N_5185);
or U5552 (N_5552,N_5201,N_5232);
nand U5553 (N_5553,N_5039,N_5451);
xnor U5554 (N_5554,N_5180,N_5484);
and U5555 (N_5555,N_5173,N_5231);
or U5556 (N_5556,N_5136,N_5463);
and U5557 (N_5557,N_5256,N_5044);
or U5558 (N_5558,N_5273,N_5206);
or U5559 (N_5559,N_5152,N_5100);
nor U5560 (N_5560,N_5416,N_5112);
nor U5561 (N_5561,N_5125,N_5291);
or U5562 (N_5562,N_5399,N_5011);
xor U5563 (N_5563,N_5266,N_5116);
xnor U5564 (N_5564,N_5072,N_5108);
and U5565 (N_5565,N_5373,N_5377);
xor U5566 (N_5566,N_5087,N_5069);
nand U5567 (N_5567,N_5407,N_5455);
and U5568 (N_5568,N_5461,N_5186);
or U5569 (N_5569,N_5468,N_5002);
nor U5570 (N_5570,N_5209,N_5017);
nand U5571 (N_5571,N_5048,N_5181);
and U5572 (N_5572,N_5348,N_5226);
or U5573 (N_5573,N_5095,N_5329);
and U5574 (N_5574,N_5205,N_5384);
or U5575 (N_5575,N_5028,N_5085);
nand U5576 (N_5576,N_5303,N_5380);
nand U5577 (N_5577,N_5216,N_5271);
nand U5578 (N_5578,N_5092,N_5242);
and U5579 (N_5579,N_5429,N_5008);
xor U5580 (N_5580,N_5022,N_5140);
or U5581 (N_5581,N_5473,N_5055);
nand U5582 (N_5582,N_5158,N_5188);
nor U5583 (N_5583,N_5375,N_5281);
nand U5584 (N_5584,N_5332,N_5390);
and U5585 (N_5585,N_5010,N_5149);
xor U5586 (N_5586,N_5410,N_5223);
nand U5587 (N_5587,N_5472,N_5436);
nand U5588 (N_5588,N_5075,N_5298);
nor U5589 (N_5589,N_5033,N_5497);
xnor U5590 (N_5590,N_5282,N_5275);
and U5591 (N_5591,N_5224,N_5113);
xnor U5592 (N_5592,N_5424,N_5306);
nor U5593 (N_5593,N_5066,N_5105);
nand U5594 (N_5594,N_5370,N_5210);
and U5595 (N_5595,N_5096,N_5386);
nor U5596 (N_5596,N_5005,N_5107);
xnor U5597 (N_5597,N_5225,N_5228);
nor U5598 (N_5598,N_5238,N_5162);
nor U5599 (N_5599,N_5115,N_5371);
xor U5600 (N_5600,N_5426,N_5431);
or U5601 (N_5601,N_5151,N_5218);
nand U5602 (N_5602,N_5450,N_5419);
or U5603 (N_5603,N_5333,N_5111);
or U5604 (N_5604,N_5475,N_5167);
xnor U5605 (N_5605,N_5109,N_5466);
nand U5606 (N_5606,N_5395,N_5104);
nand U5607 (N_5607,N_5402,N_5182);
or U5608 (N_5608,N_5358,N_5018);
xnor U5609 (N_5609,N_5406,N_5076);
or U5610 (N_5610,N_5383,N_5070);
nand U5611 (N_5611,N_5063,N_5311);
nor U5612 (N_5612,N_5364,N_5396);
and U5613 (N_5613,N_5175,N_5004);
nor U5614 (N_5614,N_5040,N_5194);
or U5615 (N_5615,N_5270,N_5049);
nor U5616 (N_5616,N_5252,N_5482);
nand U5617 (N_5617,N_5053,N_5014);
and U5618 (N_5618,N_5289,N_5486);
or U5619 (N_5619,N_5082,N_5074);
nor U5620 (N_5620,N_5367,N_5313);
or U5621 (N_5621,N_5229,N_5138);
or U5622 (N_5622,N_5071,N_5346);
xnor U5623 (N_5623,N_5335,N_5480);
nand U5624 (N_5624,N_5099,N_5496);
or U5625 (N_5625,N_5160,N_5293);
nand U5626 (N_5626,N_5304,N_5265);
nor U5627 (N_5627,N_5062,N_5203);
xnor U5628 (N_5628,N_5453,N_5404);
and U5629 (N_5629,N_5045,N_5081);
nor U5630 (N_5630,N_5278,N_5183);
or U5631 (N_5631,N_5401,N_5403);
and U5632 (N_5632,N_5012,N_5459);
nand U5633 (N_5633,N_5067,N_5485);
or U5634 (N_5634,N_5487,N_5248);
nor U5635 (N_5635,N_5476,N_5262);
xnor U5636 (N_5636,N_5433,N_5470);
nand U5637 (N_5637,N_5241,N_5341);
nor U5638 (N_5638,N_5397,N_5222);
or U5639 (N_5639,N_5050,N_5312);
nor U5640 (N_5640,N_5456,N_5280);
nand U5641 (N_5641,N_5056,N_5009);
and U5642 (N_5642,N_5240,N_5051);
nor U5643 (N_5643,N_5172,N_5000);
nor U5644 (N_5644,N_5378,N_5123);
nand U5645 (N_5645,N_5208,N_5089);
nand U5646 (N_5646,N_5192,N_5247);
nor U5647 (N_5647,N_5369,N_5454);
nor U5648 (N_5648,N_5412,N_5362);
xnor U5649 (N_5649,N_5032,N_5297);
nor U5650 (N_5650,N_5327,N_5350);
nand U5651 (N_5651,N_5091,N_5041);
or U5652 (N_5652,N_5078,N_5315);
nor U5653 (N_5653,N_5337,N_5325);
nand U5654 (N_5654,N_5295,N_5143);
nand U5655 (N_5655,N_5144,N_5423);
and U5656 (N_5656,N_5083,N_5310);
nor U5657 (N_5657,N_5184,N_5440);
and U5658 (N_5658,N_5495,N_5142);
and U5659 (N_5659,N_5054,N_5465);
xor U5660 (N_5660,N_5170,N_5294);
or U5661 (N_5661,N_5368,N_5417);
and U5662 (N_5662,N_5093,N_5150);
xor U5663 (N_5663,N_5260,N_5128);
or U5664 (N_5664,N_5199,N_5215);
xnor U5665 (N_5665,N_5493,N_5323);
and U5666 (N_5666,N_5338,N_5133);
and U5667 (N_5667,N_5147,N_5491);
nand U5668 (N_5668,N_5126,N_5359);
xnor U5669 (N_5669,N_5003,N_5422);
nor U5670 (N_5670,N_5393,N_5139);
nor U5671 (N_5671,N_5007,N_5269);
nand U5672 (N_5672,N_5239,N_5253);
or U5673 (N_5673,N_5445,N_5068);
xor U5674 (N_5674,N_5447,N_5177);
nor U5675 (N_5675,N_5145,N_5305);
or U5676 (N_5676,N_5394,N_5258);
and U5677 (N_5677,N_5425,N_5020);
or U5678 (N_5678,N_5322,N_5101);
or U5679 (N_5679,N_5060,N_5148);
nand U5680 (N_5680,N_5227,N_5233);
and U5681 (N_5681,N_5388,N_5342);
or U5682 (N_5682,N_5097,N_5361);
or U5683 (N_5683,N_5135,N_5080);
or U5684 (N_5684,N_5360,N_5340);
or U5685 (N_5685,N_5339,N_5174);
and U5686 (N_5686,N_5355,N_5254);
nor U5687 (N_5687,N_5319,N_5442);
nand U5688 (N_5688,N_5443,N_5490);
nor U5689 (N_5689,N_5168,N_5120);
or U5690 (N_5690,N_5257,N_5036);
or U5691 (N_5691,N_5084,N_5457);
or U5692 (N_5692,N_5328,N_5098);
and U5693 (N_5693,N_5157,N_5027);
or U5694 (N_5694,N_5408,N_5046);
and U5695 (N_5695,N_5119,N_5043);
nand U5696 (N_5696,N_5251,N_5287);
nand U5697 (N_5697,N_5244,N_5376);
or U5698 (N_5698,N_5405,N_5331);
nor U5699 (N_5699,N_5420,N_5195);
xor U5700 (N_5700,N_5122,N_5234);
or U5701 (N_5701,N_5460,N_5288);
or U5702 (N_5702,N_5204,N_5047);
xor U5703 (N_5703,N_5488,N_5019);
or U5704 (N_5704,N_5324,N_5439);
or U5705 (N_5705,N_5352,N_5110);
and U5706 (N_5706,N_5481,N_5290);
or U5707 (N_5707,N_5141,N_5277);
nand U5708 (N_5708,N_5307,N_5146);
and U5709 (N_5709,N_5374,N_5314);
nand U5710 (N_5710,N_5382,N_5006);
nor U5711 (N_5711,N_5357,N_5013);
and U5712 (N_5712,N_5479,N_5285);
and U5713 (N_5713,N_5058,N_5302);
nand U5714 (N_5714,N_5189,N_5347);
nand U5715 (N_5715,N_5427,N_5414);
or U5716 (N_5716,N_5446,N_5038);
or U5717 (N_5717,N_5316,N_5356);
and U5718 (N_5718,N_5366,N_5398);
and U5719 (N_5719,N_5118,N_5077);
nor U5720 (N_5720,N_5114,N_5217);
nand U5721 (N_5721,N_5190,N_5292);
and U5722 (N_5722,N_5385,N_5023);
nand U5723 (N_5723,N_5272,N_5245);
nand U5724 (N_5724,N_5309,N_5086);
nand U5725 (N_5725,N_5163,N_5134);
and U5726 (N_5726,N_5197,N_5131);
or U5727 (N_5727,N_5489,N_5268);
xor U5728 (N_5728,N_5353,N_5198);
nand U5729 (N_5729,N_5267,N_5300);
or U5730 (N_5730,N_5430,N_5061);
or U5731 (N_5731,N_5121,N_5469);
or U5732 (N_5732,N_5344,N_5448);
xnor U5733 (N_5733,N_5387,N_5236);
and U5734 (N_5734,N_5042,N_5276);
and U5735 (N_5735,N_5413,N_5343);
nor U5736 (N_5736,N_5193,N_5432);
nor U5737 (N_5737,N_5389,N_5345);
and U5738 (N_5738,N_5308,N_5166);
nand U5739 (N_5739,N_5492,N_5317);
nand U5740 (N_5740,N_5159,N_5391);
nand U5741 (N_5741,N_5237,N_5464);
or U5742 (N_5742,N_5449,N_5499);
nand U5743 (N_5743,N_5478,N_5015);
xnor U5744 (N_5744,N_5154,N_5034);
nand U5745 (N_5745,N_5365,N_5320);
xor U5746 (N_5746,N_5026,N_5031);
nand U5747 (N_5747,N_5467,N_5411);
xor U5748 (N_5748,N_5400,N_5165);
or U5749 (N_5749,N_5211,N_5102);
xor U5750 (N_5750,N_5326,N_5181);
and U5751 (N_5751,N_5239,N_5497);
and U5752 (N_5752,N_5475,N_5498);
nand U5753 (N_5753,N_5435,N_5133);
and U5754 (N_5754,N_5460,N_5236);
nor U5755 (N_5755,N_5384,N_5028);
and U5756 (N_5756,N_5384,N_5269);
nand U5757 (N_5757,N_5056,N_5299);
and U5758 (N_5758,N_5197,N_5114);
and U5759 (N_5759,N_5054,N_5372);
or U5760 (N_5760,N_5151,N_5442);
or U5761 (N_5761,N_5272,N_5487);
nor U5762 (N_5762,N_5170,N_5375);
xor U5763 (N_5763,N_5326,N_5319);
or U5764 (N_5764,N_5349,N_5360);
nand U5765 (N_5765,N_5254,N_5443);
nor U5766 (N_5766,N_5232,N_5121);
and U5767 (N_5767,N_5142,N_5060);
and U5768 (N_5768,N_5235,N_5408);
nor U5769 (N_5769,N_5395,N_5473);
nor U5770 (N_5770,N_5140,N_5123);
xnor U5771 (N_5771,N_5166,N_5186);
and U5772 (N_5772,N_5388,N_5428);
xnor U5773 (N_5773,N_5064,N_5032);
nand U5774 (N_5774,N_5270,N_5390);
nor U5775 (N_5775,N_5157,N_5097);
nor U5776 (N_5776,N_5359,N_5404);
nor U5777 (N_5777,N_5435,N_5432);
or U5778 (N_5778,N_5170,N_5309);
xnor U5779 (N_5779,N_5492,N_5281);
or U5780 (N_5780,N_5484,N_5316);
xor U5781 (N_5781,N_5460,N_5421);
and U5782 (N_5782,N_5029,N_5273);
or U5783 (N_5783,N_5131,N_5296);
and U5784 (N_5784,N_5325,N_5031);
xor U5785 (N_5785,N_5324,N_5187);
or U5786 (N_5786,N_5493,N_5349);
nand U5787 (N_5787,N_5290,N_5212);
and U5788 (N_5788,N_5288,N_5312);
nor U5789 (N_5789,N_5369,N_5139);
nor U5790 (N_5790,N_5202,N_5262);
nand U5791 (N_5791,N_5381,N_5488);
and U5792 (N_5792,N_5194,N_5429);
nor U5793 (N_5793,N_5284,N_5156);
nand U5794 (N_5794,N_5217,N_5136);
or U5795 (N_5795,N_5181,N_5083);
nor U5796 (N_5796,N_5273,N_5319);
nor U5797 (N_5797,N_5134,N_5411);
nand U5798 (N_5798,N_5379,N_5156);
nand U5799 (N_5799,N_5400,N_5079);
or U5800 (N_5800,N_5379,N_5012);
nor U5801 (N_5801,N_5389,N_5150);
xnor U5802 (N_5802,N_5121,N_5324);
xnor U5803 (N_5803,N_5009,N_5439);
nand U5804 (N_5804,N_5307,N_5218);
and U5805 (N_5805,N_5474,N_5161);
nor U5806 (N_5806,N_5471,N_5240);
and U5807 (N_5807,N_5374,N_5211);
nand U5808 (N_5808,N_5099,N_5498);
or U5809 (N_5809,N_5475,N_5155);
and U5810 (N_5810,N_5360,N_5147);
and U5811 (N_5811,N_5341,N_5457);
and U5812 (N_5812,N_5206,N_5172);
and U5813 (N_5813,N_5198,N_5376);
nand U5814 (N_5814,N_5372,N_5112);
nor U5815 (N_5815,N_5486,N_5483);
and U5816 (N_5816,N_5388,N_5393);
or U5817 (N_5817,N_5385,N_5029);
or U5818 (N_5818,N_5089,N_5154);
and U5819 (N_5819,N_5337,N_5051);
xnor U5820 (N_5820,N_5292,N_5008);
and U5821 (N_5821,N_5309,N_5440);
and U5822 (N_5822,N_5354,N_5415);
or U5823 (N_5823,N_5182,N_5338);
nand U5824 (N_5824,N_5214,N_5192);
nand U5825 (N_5825,N_5049,N_5245);
and U5826 (N_5826,N_5445,N_5412);
nand U5827 (N_5827,N_5261,N_5464);
nor U5828 (N_5828,N_5255,N_5294);
nand U5829 (N_5829,N_5100,N_5130);
nand U5830 (N_5830,N_5154,N_5167);
or U5831 (N_5831,N_5340,N_5090);
or U5832 (N_5832,N_5338,N_5140);
nor U5833 (N_5833,N_5313,N_5052);
nand U5834 (N_5834,N_5100,N_5263);
and U5835 (N_5835,N_5067,N_5075);
and U5836 (N_5836,N_5349,N_5133);
xnor U5837 (N_5837,N_5078,N_5246);
nor U5838 (N_5838,N_5447,N_5451);
xor U5839 (N_5839,N_5031,N_5461);
and U5840 (N_5840,N_5055,N_5233);
or U5841 (N_5841,N_5045,N_5228);
and U5842 (N_5842,N_5131,N_5165);
and U5843 (N_5843,N_5353,N_5105);
and U5844 (N_5844,N_5286,N_5372);
xor U5845 (N_5845,N_5316,N_5057);
and U5846 (N_5846,N_5126,N_5270);
and U5847 (N_5847,N_5162,N_5079);
nor U5848 (N_5848,N_5473,N_5171);
and U5849 (N_5849,N_5461,N_5093);
or U5850 (N_5850,N_5043,N_5102);
nor U5851 (N_5851,N_5024,N_5047);
or U5852 (N_5852,N_5329,N_5127);
and U5853 (N_5853,N_5176,N_5394);
nand U5854 (N_5854,N_5338,N_5128);
nand U5855 (N_5855,N_5053,N_5442);
and U5856 (N_5856,N_5056,N_5236);
nand U5857 (N_5857,N_5410,N_5259);
or U5858 (N_5858,N_5050,N_5336);
or U5859 (N_5859,N_5129,N_5114);
and U5860 (N_5860,N_5013,N_5349);
nor U5861 (N_5861,N_5494,N_5321);
and U5862 (N_5862,N_5487,N_5341);
nand U5863 (N_5863,N_5459,N_5437);
and U5864 (N_5864,N_5250,N_5301);
and U5865 (N_5865,N_5493,N_5364);
nand U5866 (N_5866,N_5349,N_5215);
nor U5867 (N_5867,N_5380,N_5108);
or U5868 (N_5868,N_5449,N_5183);
xor U5869 (N_5869,N_5238,N_5269);
nand U5870 (N_5870,N_5092,N_5181);
nor U5871 (N_5871,N_5338,N_5061);
or U5872 (N_5872,N_5495,N_5203);
and U5873 (N_5873,N_5426,N_5395);
nand U5874 (N_5874,N_5129,N_5051);
xnor U5875 (N_5875,N_5031,N_5484);
nand U5876 (N_5876,N_5006,N_5439);
nor U5877 (N_5877,N_5328,N_5225);
or U5878 (N_5878,N_5499,N_5108);
and U5879 (N_5879,N_5066,N_5188);
or U5880 (N_5880,N_5286,N_5429);
and U5881 (N_5881,N_5294,N_5103);
and U5882 (N_5882,N_5038,N_5479);
and U5883 (N_5883,N_5061,N_5251);
and U5884 (N_5884,N_5312,N_5134);
nand U5885 (N_5885,N_5438,N_5107);
nand U5886 (N_5886,N_5361,N_5201);
and U5887 (N_5887,N_5413,N_5055);
and U5888 (N_5888,N_5463,N_5237);
nand U5889 (N_5889,N_5265,N_5384);
nand U5890 (N_5890,N_5404,N_5021);
nor U5891 (N_5891,N_5371,N_5438);
and U5892 (N_5892,N_5250,N_5014);
nand U5893 (N_5893,N_5336,N_5358);
nand U5894 (N_5894,N_5175,N_5425);
nor U5895 (N_5895,N_5459,N_5216);
or U5896 (N_5896,N_5334,N_5191);
and U5897 (N_5897,N_5069,N_5413);
or U5898 (N_5898,N_5228,N_5361);
or U5899 (N_5899,N_5154,N_5010);
xnor U5900 (N_5900,N_5091,N_5390);
nand U5901 (N_5901,N_5030,N_5104);
nor U5902 (N_5902,N_5348,N_5165);
or U5903 (N_5903,N_5457,N_5362);
or U5904 (N_5904,N_5459,N_5424);
nor U5905 (N_5905,N_5371,N_5367);
nand U5906 (N_5906,N_5336,N_5414);
nor U5907 (N_5907,N_5042,N_5062);
nor U5908 (N_5908,N_5313,N_5291);
nor U5909 (N_5909,N_5009,N_5119);
nand U5910 (N_5910,N_5047,N_5430);
nor U5911 (N_5911,N_5296,N_5226);
nand U5912 (N_5912,N_5154,N_5164);
or U5913 (N_5913,N_5304,N_5354);
nor U5914 (N_5914,N_5386,N_5230);
nor U5915 (N_5915,N_5453,N_5240);
xor U5916 (N_5916,N_5205,N_5148);
nand U5917 (N_5917,N_5000,N_5343);
or U5918 (N_5918,N_5079,N_5422);
or U5919 (N_5919,N_5043,N_5492);
or U5920 (N_5920,N_5438,N_5040);
xor U5921 (N_5921,N_5229,N_5224);
or U5922 (N_5922,N_5238,N_5353);
xnor U5923 (N_5923,N_5450,N_5106);
nand U5924 (N_5924,N_5230,N_5010);
nand U5925 (N_5925,N_5037,N_5211);
and U5926 (N_5926,N_5170,N_5010);
nor U5927 (N_5927,N_5488,N_5435);
nor U5928 (N_5928,N_5131,N_5281);
nor U5929 (N_5929,N_5081,N_5437);
nor U5930 (N_5930,N_5429,N_5452);
nand U5931 (N_5931,N_5045,N_5365);
or U5932 (N_5932,N_5006,N_5147);
and U5933 (N_5933,N_5309,N_5132);
and U5934 (N_5934,N_5377,N_5309);
and U5935 (N_5935,N_5098,N_5060);
nor U5936 (N_5936,N_5107,N_5024);
and U5937 (N_5937,N_5294,N_5432);
nor U5938 (N_5938,N_5425,N_5172);
or U5939 (N_5939,N_5002,N_5136);
nand U5940 (N_5940,N_5459,N_5392);
nand U5941 (N_5941,N_5265,N_5144);
nand U5942 (N_5942,N_5155,N_5423);
and U5943 (N_5943,N_5062,N_5310);
nand U5944 (N_5944,N_5391,N_5153);
or U5945 (N_5945,N_5172,N_5412);
nor U5946 (N_5946,N_5097,N_5332);
xnor U5947 (N_5947,N_5248,N_5202);
and U5948 (N_5948,N_5282,N_5380);
xnor U5949 (N_5949,N_5437,N_5390);
nor U5950 (N_5950,N_5104,N_5231);
or U5951 (N_5951,N_5494,N_5133);
and U5952 (N_5952,N_5057,N_5249);
nor U5953 (N_5953,N_5282,N_5231);
nor U5954 (N_5954,N_5024,N_5103);
and U5955 (N_5955,N_5374,N_5175);
nand U5956 (N_5956,N_5466,N_5376);
or U5957 (N_5957,N_5152,N_5462);
nand U5958 (N_5958,N_5189,N_5142);
xnor U5959 (N_5959,N_5218,N_5231);
and U5960 (N_5960,N_5182,N_5245);
nor U5961 (N_5961,N_5038,N_5426);
xor U5962 (N_5962,N_5432,N_5288);
or U5963 (N_5963,N_5172,N_5153);
nand U5964 (N_5964,N_5211,N_5062);
and U5965 (N_5965,N_5255,N_5263);
nand U5966 (N_5966,N_5469,N_5230);
or U5967 (N_5967,N_5490,N_5339);
nor U5968 (N_5968,N_5236,N_5465);
or U5969 (N_5969,N_5352,N_5362);
xor U5970 (N_5970,N_5324,N_5434);
nor U5971 (N_5971,N_5410,N_5430);
nand U5972 (N_5972,N_5215,N_5031);
and U5973 (N_5973,N_5422,N_5050);
or U5974 (N_5974,N_5312,N_5235);
and U5975 (N_5975,N_5466,N_5044);
and U5976 (N_5976,N_5313,N_5144);
or U5977 (N_5977,N_5070,N_5457);
and U5978 (N_5978,N_5152,N_5472);
nand U5979 (N_5979,N_5288,N_5207);
or U5980 (N_5980,N_5237,N_5089);
and U5981 (N_5981,N_5218,N_5000);
nand U5982 (N_5982,N_5498,N_5081);
nand U5983 (N_5983,N_5466,N_5479);
xnor U5984 (N_5984,N_5076,N_5054);
nand U5985 (N_5985,N_5004,N_5368);
nor U5986 (N_5986,N_5320,N_5415);
or U5987 (N_5987,N_5049,N_5031);
and U5988 (N_5988,N_5117,N_5352);
or U5989 (N_5989,N_5227,N_5275);
xnor U5990 (N_5990,N_5123,N_5427);
or U5991 (N_5991,N_5158,N_5452);
nor U5992 (N_5992,N_5312,N_5148);
nor U5993 (N_5993,N_5288,N_5376);
and U5994 (N_5994,N_5145,N_5302);
and U5995 (N_5995,N_5044,N_5277);
nand U5996 (N_5996,N_5028,N_5414);
nand U5997 (N_5997,N_5282,N_5169);
and U5998 (N_5998,N_5320,N_5148);
nand U5999 (N_5999,N_5159,N_5265);
or U6000 (N_6000,N_5636,N_5901);
or U6001 (N_6001,N_5956,N_5593);
or U6002 (N_6002,N_5624,N_5869);
xnor U6003 (N_6003,N_5508,N_5530);
or U6004 (N_6004,N_5719,N_5726);
nand U6005 (N_6005,N_5724,N_5537);
nor U6006 (N_6006,N_5880,N_5543);
nand U6007 (N_6007,N_5617,N_5698);
nand U6008 (N_6008,N_5524,N_5737);
and U6009 (N_6009,N_5884,N_5587);
or U6010 (N_6010,N_5656,N_5538);
nand U6011 (N_6011,N_5977,N_5986);
and U6012 (N_6012,N_5984,N_5888);
and U6013 (N_6013,N_5818,N_5792);
or U6014 (N_6014,N_5753,N_5970);
xor U6015 (N_6015,N_5575,N_5758);
nand U6016 (N_6016,N_5500,N_5692);
and U6017 (N_6017,N_5722,N_5582);
and U6018 (N_6018,N_5931,N_5682);
and U6019 (N_6019,N_5921,N_5657);
or U6020 (N_6020,N_5772,N_5746);
xor U6021 (N_6021,N_5777,N_5728);
nand U6022 (N_6022,N_5563,N_5566);
nor U6023 (N_6023,N_5628,N_5664);
nand U6024 (N_6024,N_5847,N_5825);
nand U6025 (N_6025,N_5525,N_5509);
or U6026 (N_6026,N_5705,N_5642);
nand U6027 (N_6027,N_5765,N_5936);
nor U6028 (N_6028,N_5916,N_5735);
nand U6029 (N_6029,N_5954,N_5790);
or U6030 (N_6030,N_5793,N_5743);
and U6031 (N_6031,N_5996,N_5623);
and U6032 (N_6032,N_5748,N_5544);
nor U6033 (N_6033,N_5852,N_5565);
nand U6034 (N_6034,N_5967,N_5943);
nand U6035 (N_6035,N_5928,N_5640);
nor U6036 (N_6036,N_5918,N_5653);
and U6037 (N_6037,N_5620,N_5570);
nor U6038 (N_6038,N_5929,N_5590);
or U6039 (N_6039,N_5740,N_5502);
or U6040 (N_6040,N_5545,N_5529);
or U6041 (N_6041,N_5554,N_5690);
nand U6042 (N_6042,N_5896,N_5650);
nand U6043 (N_6043,N_5811,N_5742);
nor U6044 (N_6044,N_5823,N_5668);
and U6045 (N_6045,N_5798,N_5534);
or U6046 (N_6046,N_5787,N_5932);
or U6047 (N_6047,N_5683,N_5714);
nand U6048 (N_6048,N_5906,N_5859);
and U6049 (N_6049,N_5696,N_5820);
xor U6050 (N_6050,N_5540,N_5716);
nor U6051 (N_6051,N_5837,N_5908);
nor U6052 (N_6052,N_5618,N_5842);
nor U6053 (N_6053,N_5784,N_5843);
nor U6054 (N_6054,N_5872,N_5699);
or U6055 (N_6055,N_5754,N_5581);
or U6056 (N_6056,N_5942,N_5868);
nor U6057 (N_6057,N_5881,N_5681);
and U6058 (N_6058,N_5610,N_5514);
nor U6059 (N_6059,N_5971,N_5713);
nor U6060 (N_6060,N_5834,N_5652);
nor U6061 (N_6061,N_5505,N_5677);
or U6062 (N_6062,N_5518,N_5973);
nand U6063 (N_6063,N_5694,N_5938);
nand U6064 (N_6064,N_5531,N_5991);
nand U6065 (N_6065,N_5846,N_5645);
nand U6066 (N_6066,N_5701,N_5526);
nor U6067 (N_6067,N_5813,N_5771);
or U6068 (N_6068,N_5700,N_5957);
nand U6069 (N_6069,N_5584,N_5744);
or U6070 (N_6070,N_5638,N_5976);
nand U6071 (N_6071,N_5717,N_5999);
xnor U6072 (N_6072,N_5863,N_5568);
xor U6073 (N_6073,N_5604,N_5731);
and U6074 (N_6074,N_5785,N_5964);
xnor U6075 (N_6075,N_5870,N_5797);
nand U6076 (N_6076,N_5802,N_5925);
nand U6077 (N_6077,N_5806,N_5560);
nand U6078 (N_6078,N_5917,N_5639);
and U6079 (N_6079,N_5774,N_5800);
and U6080 (N_6080,N_5559,N_5648);
xnor U6081 (N_6081,N_5807,N_5920);
or U6082 (N_6082,N_5879,N_5861);
and U6083 (N_6083,N_5789,N_5952);
xor U6084 (N_6084,N_5539,N_5583);
xnor U6085 (N_6085,N_5609,N_5550);
and U6086 (N_6086,N_5835,N_5911);
xnor U6087 (N_6087,N_5962,N_5541);
or U6088 (N_6088,N_5643,N_5886);
and U6089 (N_6089,N_5922,N_5632);
nand U6090 (N_6090,N_5972,N_5569);
and U6091 (N_6091,N_5893,N_5527);
and U6092 (N_6092,N_5864,N_5989);
nor U6093 (N_6093,N_5902,N_5833);
nor U6094 (N_6094,N_5799,N_5738);
or U6095 (N_6095,N_5891,N_5909);
and U6096 (N_6096,N_5907,N_5979);
and U6097 (N_6097,N_5983,N_5990);
and U6098 (N_6098,N_5598,N_5619);
nand U6099 (N_6099,N_5821,N_5615);
or U6100 (N_6100,N_5873,N_5998);
or U6101 (N_6101,N_5899,N_5766);
nand U6102 (N_6102,N_5519,N_5764);
nand U6103 (N_6103,N_5750,N_5839);
and U6104 (N_6104,N_5840,N_5562);
nor U6105 (N_6105,N_5564,N_5555);
or U6106 (N_6106,N_5997,N_5558);
or U6107 (N_6107,N_5680,N_5588);
nand U6108 (N_6108,N_5781,N_5730);
nor U6109 (N_6109,N_5892,N_5702);
nand U6110 (N_6110,N_5578,N_5994);
and U6111 (N_6111,N_5723,N_5817);
nand U6112 (N_6112,N_5860,N_5599);
nor U6113 (N_6113,N_5670,N_5912);
nor U6114 (N_6114,N_5944,N_5549);
and U6115 (N_6115,N_5733,N_5732);
nand U6116 (N_6116,N_5595,N_5865);
or U6117 (N_6117,N_5987,N_5579);
nor U6118 (N_6118,N_5969,N_5646);
and U6119 (N_6119,N_5779,N_5915);
or U6120 (N_6120,N_5801,N_5946);
xnor U6121 (N_6121,N_5889,N_5858);
xor U6122 (N_6122,N_5651,N_5769);
xor U6123 (N_6123,N_5824,N_5649);
or U6124 (N_6124,N_5751,N_5535);
and U6125 (N_6125,N_5605,N_5795);
xnor U6126 (N_6126,N_5687,N_5745);
nand U6127 (N_6127,N_5673,N_5600);
nor U6128 (N_6128,N_5857,N_5506);
or U6129 (N_6129,N_5688,N_5819);
nor U6130 (N_6130,N_5803,N_5547);
and U6131 (N_6131,N_5783,N_5796);
or U6132 (N_6132,N_5725,N_5577);
and U6133 (N_6133,N_5591,N_5988);
and U6134 (N_6134,N_5704,N_5760);
xnor U6135 (N_6135,N_5992,N_5955);
and U6136 (N_6136,N_5883,N_5561);
or U6137 (N_6137,N_5721,N_5836);
nor U6138 (N_6138,N_5630,N_5845);
nand U6139 (N_6139,N_5691,N_5878);
or U6140 (N_6140,N_5631,N_5809);
nor U6141 (N_6141,N_5968,N_5685);
and U6142 (N_6142,N_5963,N_5671);
nand U6143 (N_6143,N_5965,N_5612);
nor U6144 (N_6144,N_5551,N_5904);
and U6145 (N_6145,N_5810,N_5930);
xnor U6146 (N_6146,N_5669,N_5940);
or U6147 (N_6147,N_5981,N_5676);
nor U6148 (N_6148,N_5849,N_5914);
nor U6149 (N_6149,N_5655,N_5910);
and U6150 (N_6150,N_5625,N_5718);
nand U6151 (N_6151,N_5934,N_5712);
or U6152 (N_6152,N_5993,N_5557);
or U6153 (N_6153,N_5603,N_5850);
or U6154 (N_6154,N_5975,N_5585);
nor U6155 (N_6155,N_5567,N_5596);
nor U6156 (N_6156,N_5814,N_5747);
nor U6157 (N_6157,N_5621,N_5919);
or U6158 (N_6158,N_5961,N_5887);
or U6159 (N_6159,N_5542,N_5895);
nand U6160 (N_6160,N_5877,N_5788);
or U6161 (N_6161,N_5660,N_5511);
nand U6162 (N_6162,N_5826,N_5903);
and U6163 (N_6163,N_5611,N_5851);
or U6164 (N_6164,N_5629,N_5951);
and U6165 (N_6165,N_5644,N_5770);
nor U6166 (N_6166,N_5586,N_5985);
nand U6167 (N_6167,N_5841,N_5900);
nor U6168 (N_6168,N_5815,N_5830);
nand U6169 (N_6169,N_5667,N_5672);
and U6170 (N_6170,N_5749,N_5866);
or U6171 (N_6171,N_5752,N_5601);
nor U6172 (N_6172,N_5768,N_5614);
nand U6173 (N_6173,N_5707,N_5710);
xnor U6174 (N_6174,N_5831,N_5945);
or U6175 (N_6175,N_5756,N_5695);
or U6176 (N_6176,N_5662,N_5854);
or U6177 (N_6177,N_5520,N_5924);
or U6178 (N_6178,N_5693,N_5533);
xnor U6179 (N_6179,N_5580,N_5727);
nand U6180 (N_6180,N_5678,N_5855);
nand U6181 (N_6181,N_5808,N_5980);
and U6182 (N_6182,N_5504,N_5926);
nand U6183 (N_6183,N_5947,N_5822);
xor U6184 (N_6184,N_5602,N_5510);
and U6185 (N_6185,N_5776,N_5734);
xnor U6186 (N_6186,N_5715,N_5927);
or U6187 (N_6187,N_5829,N_5757);
nor U6188 (N_6188,N_5546,N_5503);
or U6189 (N_6189,N_5665,N_5708);
nor U6190 (N_6190,N_5689,N_5606);
nand U6191 (N_6191,N_5923,N_5675);
and U6192 (N_6192,N_5939,N_5736);
nor U6193 (N_6193,N_5536,N_5882);
nor U6194 (N_6194,N_5515,N_5513);
or U6195 (N_6195,N_5607,N_5637);
nor U6196 (N_6196,N_5684,N_5523);
nor U6197 (N_6197,N_5871,N_5832);
nand U6198 (N_6198,N_5828,N_5633);
or U6199 (N_6199,N_5532,N_5661);
nor U6200 (N_6200,N_5626,N_5804);
nand U6201 (N_6201,N_5573,N_5780);
nor U6202 (N_6202,N_5791,N_5966);
or U6203 (N_6203,N_5805,N_5978);
or U6204 (N_6204,N_5572,N_5627);
nor U6205 (N_6205,N_5816,N_5674);
and U6206 (N_6206,N_5641,N_5666);
xnor U6207 (N_6207,N_5786,N_5827);
nor U6208 (N_6208,N_5521,N_5634);
nor U6209 (N_6209,N_5528,N_5720);
nor U6210 (N_6210,N_5773,N_5862);
or U6211 (N_6211,N_5594,N_5812);
and U6212 (N_6212,N_5876,N_5890);
xor U6213 (N_6213,N_5517,N_5686);
nand U6214 (N_6214,N_5767,N_5553);
nand U6215 (N_6215,N_5658,N_5763);
and U6216 (N_6216,N_5522,N_5755);
or U6217 (N_6217,N_5709,N_5574);
xor U6218 (N_6218,N_5654,N_5597);
nor U6219 (N_6219,N_5875,N_5608);
nand U6220 (N_6220,N_5759,N_5512);
or U6221 (N_6221,N_5838,N_5933);
nor U6222 (N_6222,N_5711,N_5706);
nand U6223 (N_6223,N_5663,N_5794);
or U6224 (N_6224,N_5741,N_5613);
nand U6225 (N_6225,N_5635,N_5935);
or U6226 (N_6226,N_5867,N_5897);
nor U6227 (N_6227,N_5697,N_5974);
and U6228 (N_6228,N_5552,N_5622);
nand U6229 (N_6229,N_5729,N_5950);
or U6230 (N_6230,N_5941,N_5995);
and U6231 (N_6231,N_5761,N_5856);
xor U6232 (N_6232,N_5576,N_5953);
nor U6233 (N_6233,N_5960,N_5616);
nand U6234 (N_6234,N_5982,N_5948);
nand U6235 (N_6235,N_5949,N_5958);
or U6236 (N_6236,N_5501,N_5679);
nand U6237 (N_6237,N_5905,N_5844);
or U6238 (N_6238,N_5592,N_5913);
xor U6239 (N_6239,N_5548,N_5659);
nor U6240 (N_6240,N_5778,N_5571);
nand U6241 (N_6241,N_5556,N_5589);
and U6242 (N_6242,N_5762,N_5894);
or U6243 (N_6243,N_5898,N_5516);
or U6244 (N_6244,N_5853,N_5782);
or U6245 (N_6245,N_5775,N_5885);
and U6246 (N_6246,N_5937,N_5848);
or U6247 (N_6247,N_5874,N_5703);
nand U6248 (N_6248,N_5647,N_5959);
or U6249 (N_6249,N_5739,N_5507);
nand U6250 (N_6250,N_5656,N_5976);
nor U6251 (N_6251,N_5706,N_5918);
and U6252 (N_6252,N_5674,N_5787);
xor U6253 (N_6253,N_5948,N_5542);
nor U6254 (N_6254,N_5747,N_5580);
and U6255 (N_6255,N_5570,N_5586);
nor U6256 (N_6256,N_5511,N_5954);
nand U6257 (N_6257,N_5505,N_5717);
or U6258 (N_6258,N_5584,N_5565);
nor U6259 (N_6259,N_5719,N_5909);
or U6260 (N_6260,N_5670,N_5913);
and U6261 (N_6261,N_5866,N_5932);
nor U6262 (N_6262,N_5639,N_5891);
xor U6263 (N_6263,N_5733,N_5607);
and U6264 (N_6264,N_5891,N_5587);
or U6265 (N_6265,N_5785,N_5887);
and U6266 (N_6266,N_5668,N_5783);
and U6267 (N_6267,N_5851,N_5582);
or U6268 (N_6268,N_5529,N_5719);
and U6269 (N_6269,N_5518,N_5910);
nand U6270 (N_6270,N_5984,N_5955);
nand U6271 (N_6271,N_5905,N_5653);
and U6272 (N_6272,N_5559,N_5565);
nand U6273 (N_6273,N_5768,N_5867);
nand U6274 (N_6274,N_5657,N_5990);
or U6275 (N_6275,N_5972,N_5998);
and U6276 (N_6276,N_5518,N_5557);
nand U6277 (N_6277,N_5911,N_5727);
and U6278 (N_6278,N_5719,N_5629);
or U6279 (N_6279,N_5713,N_5917);
xnor U6280 (N_6280,N_5732,N_5810);
nor U6281 (N_6281,N_5580,N_5558);
and U6282 (N_6282,N_5691,N_5546);
and U6283 (N_6283,N_5727,N_5707);
nor U6284 (N_6284,N_5915,N_5846);
or U6285 (N_6285,N_5766,N_5880);
and U6286 (N_6286,N_5921,N_5891);
or U6287 (N_6287,N_5901,N_5714);
nand U6288 (N_6288,N_5644,N_5659);
or U6289 (N_6289,N_5673,N_5902);
nor U6290 (N_6290,N_5912,N_5550);
nor U6291 (N_6291,N_5616,N_5948);
xor U6292 (N_6292,N_5668,N_5990);
and U6293 (N_6293,N_5705,N_5731);
xor U6294 (N_6294,N_5527,N_5946);
nand U6295 (N_6295,N_5986,N_5517);
nand U6296 (N_6296,N_5738,N_5867);
or U6297 (N_6297,N_5654,N_5744);
nor U6298 (N_6298,N_5646,N_5846);
nor U6299 (N_6299,N_5657,N_5905);
xnor U6300 (N_6300,N_5648,N_5563);
and U6301 (N_6301,N_5842,N_5744);
xnor U6302 (N_6302,N_5872,N_5900);
nand U6303 (N_6303,N_5813,N_5625);
nand U6304 (N_6304,N_5809,N_5873);
nand U6305 (N_6305,N_5839,N_5515);
nor U6306 (N_6306,N_5599,N_5788);
xnor U6307 (N_6307,N_5942,N_5908);
or U6308 (N_6308,N_5708,N_5938);
nand U6309 (N_6309,N_5597,N_5849);
and U6310 (N_6310,N_5954,N_5810);
or U6311 (N_6311,N_5898,N_5657);
and U6312 (N_6312,N_5634,N_5972);
and U6313 (N_6313,N_5747,N_5939);
nor U6314 (N_6314,N_5910,N_5839);
nor U6315 (N_6315,N_5612,N_5596);
nand U6316 (N_6316,N_5531,N_5784);
xor U6317 (N_6317,N_5860,N_5796);
nor U6318 (N_6318,N_5848,N_5880);
or U6319 (N_6319,N_5975,N_5782);
nor U6320 (N_6320,N_5833,N_5925);
or U6321 (N_6321,N_5955,N_5987);
nor U6322 (N_6322,N_5621,N_5568);
nand U6323 (N_6323,N_5718,N_5544);
and U6324 (N_6324,N_5835,N_5837);
nand U6325 (N_6325,N_5740,N_5840);
and U6326 (N_6326,N_5507,N_5949);
nand U6327 (N_6327,N_5779,N_5589);
or U6328 (N_6328,N_5998,N_5832);
nor U6329 (N_6329,N_5723,N_5764);
nor U6330 (N_6330,N_5888,N_5822);
nor U6331 (N_6331,N_5972,N_5598);
and U6332 (N_6332,N_5842,N_5616);
or U6333 (N_6333,N_5951,N_5585);
or U6334 (N_6334,N_5953,N_5843);
and U6335 (N_6335,N_5585,N_5518);
nor U6336 (N_6336,N_5706,N_5755);
xnor U6337 (N_6337,N_5693,N_5627);
or U6338 (N_6338,N_5684,N_5692);
or U6339 (N_6339,N_5614,N_5997);
xnor U6340 (N_6340,N_5764,N_5828);
nor U6341 (N_6341,N_5922,N_5771);
nor U6342 (N_6342,N_5628,N_5810);
nor U6343 (N_6343,N_5970,N_5712);
and U6344 (N_6344,N_5833,N_5559);
and U6345 (N_6345,N_5613,N_5688);
nor U6346 (N_6346,N_5869,N_5533);
nor U6347 (N_6347,N_5999,N_5912);
nand U6348 (N_6348,N_5555,N_5536);
nand U6349 (N_6349,N_5636,N_5725);
or U6350 (N_6350,N_5697,N_5949);
nand U6351 (N_6351,N_5843,N_5688);
and U6352 (N_6352,N_5713,N_5767);
nand U6353 (N_6353,N_5683,N_5915);
nand U6354 (N_6354,N_5762,N_5784);
nor U6355 (N_6355,N_5721,N_5699);
and U6356 (N_6356,N_5854,N_5806);
and U6357 (N_6357,N_5764,N_5870);
nor U6358 (N_6358,N_5658,N_5847);
nor U6359 (N_6359,N_5932,N_5784);
nand U6360 (N_6360,N_5717,N_5800);
or U6361 (N_6361,N_5861,N_5595);
nor U6362 (N_6362,N_5743,N_5944);
or U6363 (N_6363,N_5793,N_5609);
nor U6364 (N_6364,N_5734,N_5556);
xor U6365 (N_6365,N_5973,N_5754);
nand U6366 (N_6366,N_5804,N_5664);
nand U6367 (N_6367,N_5605,N_5533);
or U6368 (N_6368,N_5574,N_5640);
nand U6369 (N_6369,N_5569,N_5540);
and U6370 (N_6370,N_5916,N_5974);
nor U6371 (N_6371,N_5817,N_5533);
nand U6372 (N_6372,N_5806,N_5613);
nand U6373 (N_6373,N_5597,N_5818);
nor U6374 (N_6374,N_5954,N_5943);
or U6375 (N_6375,N_5766,N_5692);
nor U6376 (N_6376,N_5734,N_5879);
or U6377 (N_6377,N_5899,N_5583);
or U6378 (N_6378,N_5926,N_5867);
nor U6379 (N_6379,N_5983,N_5543);
nand U6380 (N_6380,N_5619,N_5879);
and U6381 (N_6381,N_5867,N_5504);
nor U6382 (N_6382,N_5514,N_5950);
or U6383 (N_6383,N_5820,N_5610);
nand U6384 (N_6384,N_5567,N_5819);
nor U6385 (N_6385,N_5934,N_5547);
nand U6386 (N_6386,N_5983,N_5851);
nand U6387 (N_6387,N_5512,N_5668);
or U6388 (N_6388,N_5735,N_5609);
or U6389 (N_6389,N_5983,N_5912);
xnor U6390 (N_6390,N_5954,N_5784);
nand U6391 (N_6391,N_5755,N_5619);
or U6392 (N_6392,N_5539,N_5943);
and U6393 (N_6393,N_5761,N_5816);
xor U6394 (N_6394,N_5926,N_5566);
and U6395 (N_6395,N_5508,N_5862);
xor U6396 (N_6396,N_5968,N_5740);
and U6397 (N_6397,N_5875,N_5800);
or U6398 (N_6398,N_5751,N_5513);
or U6399 (N_6399,N_5990,N_5754);
nand U6400 (N_6400,N_5768,N_5755);
xnor U6401 (N_6401,N_5796,N_5643);
nand U6402 (N_6402,N_5571,N_5956);
and U6403 (N_6403,N_5967,N_5936);
xnor U6404 (N_6404,N_5957,N_5897);
and U6405 (N_6405,N_5645,N_5606);
nand U6406 (N_6406,N_5945,N_5938);
nor U6407 (N_6407,N_5809,N_5523);
nor U6408 (N_6408,N_5717,N_5988);
nand U6409 (N_6409,N_5517,N_5821);
xnor U6410 (N_6410,N_5635,N_5911);
and U6411 (N_6411,N_5635,N_5548);
and U6412 (N_6412,N_5653,N_5575);
and U6413 (N_6413,N_5795,N_5933);
and U6414 (N_6414,N_5649,N_5538);
and U6415 (N_6415,N_5846,N_5961);
nor U6416 (N_6416,N_5781,N_5615);
nand U6417 (N_6417,N_5590,N_5570);
or U6418 (N_6418,N_5826,N_5896);
nand U6419 (N_6419,N_5740,N_5879);
or U6420 (N_6420,N_5765,N_5620);
nand U6421 (N_6421,N_5682,N_5750);
nand U6422 (N_6422,N_5738,N_5906);
or U6423 (N_6423,N_5639,N_5630);
nor U6424 (N_6424,N_5847,N_5937);
xor U6425 (N_6425,N_5816,N_5546);
nor U6426 (N_6426,N_5638,N_5762);
nor U6427 (N_6427,N_5785,N_5527);
and U6428 (N_6428,N_5881,N_5520);
and U6429 (N_6429,N_5763,N_5645);
nor U6430 (N_6430,N_5528,N_5777);
xor U6431 (N_6431,N_5555,N_5745);
and U6432 (N_6432,N_5987,N_5746);
nor U6433 (N_6433,N_5876,N_5575);
nand U6434 (N_6434,N_5632,N_5672);
nor U6435 (N_6435,N_5794,N_5725);
and U6436 (N_6436,N_5535,N_5903);
or U6437 (N_6437,N_5636,N_5639);
or U6438 (N_6438,N_5842,N_5832);
or U6439 (N_6439,N_5766,N_5907);
nor U6440 (N_6440,N_5740,N_5691);
nor U6441 (N_6441,N_5641,N_5865);
nor U6442 (N_6442,N_5964,N_5626);
nor U6443 (N_6443,N_5981,N_5709);
or U6444 (N_6444,N_5963,N_5988);
nand U6445 (N_6445,N_5971,N_5697);
and U6446 (N_6446,N_5510,N_5503);
or U6447 (N_6447,N_5639,N_5902);
nand U6448 (N_6448,N_5987,N_5928);
nand U6449 (N_6449,N_5654,N_5750);
nor U6450 (N_6450,N_5828,N_5513);
nor U6451 (N_6451,N_5627,N_5763);
or U6452 (N_6452,N_5581,N_5886);
xor U6453 (N_6453,N_5751,N_5571);
nand U6454 (N_6454,N_5984,N_5970);
nor U6455 (N_6455,N_5668,N_5989);
or U6456 (N_6456,N_5509,N_5752);
or U6457 (N_6457,N_5933,N_5843);
nor U6458 (N_6458,N_5914,N_5598);
nand U6459 (N_6459,N_5889,N_5707);
xnor U6460 (N_6460,N_5807,N_5719);
nor U6461 (N_6461,N_5746,N_5729);
or U6462 (N_6462,N_5513,N_5646);
nand U6463 (N_6463,N_5813,N_5832);
nor U6464 (N_6464,N_5809,N_5997);
nand U6465 (N_6465,N_5763,N_5966);
or U6466 (N_6466,N_5934,N_5721);
nand U6467 (N_6467,N_5652,N_5604);
or U6468 (N_6468,N_5625,N_5592);
nand U6469 (N_6469,N_5521,N_5982);
nand U6470 (N_6470,N_5851,N_5521);
nand U6471 (N_6471,N_5996,N_5909);
xor U6472 (N_6472,N_5623,N_5978);
nand U6473 (N_6473,N_5538,N_5880);
xnor U6474 (N_6474,N_5661,N_5677);
nor U6475 (N_6475,N_5627,N_5691);
nor U6476 (N_6476,N_5934,N_5562);
or U6477 (N_6477,N_5782,N_5524);
xnor U6478 (N_6478,N_5723,N_5933);
nand U6479 (N_6479,N_5691,N_5602);
and U6480 (N_6480,N_5660,N_5829);
nor U6481 (N_6481,N_5723,N_5640);
nor U6482 (N_6482,N_5976,N_5815);
or U6483 (N_6483,N_5706,N_5596);
or U6484 (N_6484,N_5763,N_5590);
and U6485 (N_6485,N_5613,N_5573);
nand U6486 (N_6486,N_5995,N_5622);
or U6487 (N_6487,N_5863,N_5903);
nor U6488 (N_6488,N_5894,N_5585);
nand U6489 (N_6489,N_5501,N_5582);
and U6490 (N_6490,N_5848,N_5734);
nor U6491 (N_6491,N_5559,N_5544);
and U6492 (N_6492,N_5987,N_5547);
or U6493 (N_6493,N_5992,N_5774);
nand U6494 (N_6494,N_5613,N_5558);
and U6495 (N_6495,N_5571,N_5883);
nand U6496 (N_6496,N_5717,N_5962);
nor U6497 (N_6497,N_5831,N_5545);
nor U6498 (N_6498,N_5937,N_5778);
or U6499 (N_6499,N_5824,N_5874);
nand U6500 (N_6500,N_6313,N_6186);
nand U6501 (N_6501,N_6085,N_6207);
nor U6502 (N_6502,N_6403,N_6081);
or U6503 (N_6503,N_6010,N_6420);
nor U6504 (N_6504,N_6386,N_6000);
nor U6505 (N_6505,N_6297,N_6099);
and U6506 (N_6506,N_6009,N_6361);
and U6507 (N_6507,N_6117,N_6499);
or U6508 (N_6508,N_6435,N_6131);
xor U6509 (N_6509,N_6123,N_6102);
or U6510 (N_6510,N_6409,N_6367);
and U6511 (N_6511,N_6395,N_6325);
nand U6512 (N_6512,N_6373,N_6048);
nand U6513 (N_6513,N_6265,N_6394);
nand U6514 (N_6514,N_6152,N_6227);
or U6515 (N_6515,N_6401,N_6416);
or U6516 (N_6516,N_6025,N_6114);
or U6517 (N_6517,N_6485,N_6143);
xor U6518 (N_6518,N_6302,N_6385);
or U6519 (N_6519,N_6321,N_6155);
nor U6520 (N_6520,N_6076,N_6380);
nand U6521 (N_6521,N_6262,N_6492);
and U6522 (N_6522,N_6029,N_6198);
and U6523 (N_6523,N_6182,N_6034);
and U6524 (N_6524,N_6032,N_6023);
and U6525 (N_6525,N_6204,N_6027);
xor U6526 (N_6526,N_6365,N_6467);
and U6527 (N_6527,N_6402,N_6413);
nor U6528 (N_6528,N_6101,N_6276);
nand U6529 (N_6529,N_6038,N_6135);
nand U6530 (N_6530,N_6478,N_6474);
nor U6531 (N_6531,N_6304,N_6178);
nor U6532 (N_6532,N_6372,N_6042);
or U6533 (N_6533,N_6315,N_6400);
or U6534 (N_6534,N_6011,N_6124);
or U6535 (N_6535,N_6169,N_6115);
or U6536 (N_6536,N_6342,N_6219);
and U6537 (N_6537,N_6410,N_6314);
and U6538 (N_6538,N_6352,N_6272);
nand U6539 (N_6539,N_6356,N_6377);
nor U6540 (N_6540,N_6061,N_6079);
nand U6541 (N_6541,N_6022,N_6484);
nor U6542 (N_6542,N_6285,N_6404);
and U6543 (N_6543,N_6220,N_6247);
xor U6544 (N_6544,N_6290,N_6370);
and U6545 (N_6545,N_6391,N_6133);
nand U6546 (N_6546,N_6084,N_6208);
and U6547 (N_6547,N_6466,N_6237);
and U6548 (N_6548,N_6390,N_6109);
or U6549 (N_6549,N_6344,N_6267);
or U6550 (N_6550,N_6147,N_6407);
or U6551 (N_6551,N_6206,N_6229);
or U6552 (N_6552,N_6111,N_6007);
or U6553 (N_6553,N_6482,N_6417);
and U6554 (N_6554,N_6296,N_6360);
or U6555 (N_6555,N_6008,N_6363);
and U6556 (N_6556,N_6187,N_6199);
nand U6557 (N_6557,N_6397,N_6246);
nand U6558 (N_6558,N_6288,N_6339);
or U6559 (N_6559,N_6145,N_6210);
and U6560 (N_6560,N_6298,N_6092);
nand U6561 (N_6561,N_6384,N_6211);
or U6562 (N_6562,N_6074,N_6281);
nor U6563 (N_6563,N_6450,N_6322);
or U6564 (N_6564,N_6162,N_6353);
and U6565 (N_6565,N_6129,N_6349);
or U6566 (N_6566,N_6055,N_6412);
and U6567 (N_6567,N_6013,N_6291);
nand U6568 (N_6568,N_6368,N_6461);
or U6569 (N_6569,N_6260,N_6170);
or U6570 (N_6570,N_6093,N_6088);
nor U6571 (N_6571,N_6414,N_6371);
or U6572 (N_6572,N_6355,N_6190);
nor U6573 (N_6573,N_6139,N_6427);
nand U6574 (N_6574,N_6137,N_6068);
nor U6575 (N_6575,N_6442,N_6446);
xnor U6576 (N_6576,N_6128,N_6497);
nand U6577 (N_6577,N_6158,N_6292);
or U6578 (N_6578,N_6398,N_6046);
nor U6579 (N_6579,N_6180,N_6421);
and U6580 (N_6580,N_6108,N_6036);
and U6581 (N_6581,N_6003,N_6033);
and U6582 (N_6582,N_6320,N_6345);
xnor U6583 (N_6583,N_6030,N_6477);
nand U6584 (N_6584,N_6144,N_6164);
or U6585 (N_6585,N_6358,N_6177);
or U6586 (N_6586,N_6159,N_6268);
and U6587 (N_6587,N_6346,N_6243);
and U6588 (N_6588,N_6455,N_6089);
nor U6589 (N_6589,N_6100,N_6098);
and U6590 (N_6590,N_6136,N_6459);
and U6591 (N_6591,N_6249,N_6294);
and U6592 (N_6592,N_6419,N_6406);
nand U6593 (N_6593,N_6496,N_6301);
or U6594 (N_6594,N_6264,N_6293);
xor U6595 (N_6595,N_6333,N_6426);
nand U6596 (N_6596,N_6295,N_6205);
nor U6597 (N_6597,N_6072,N_6222);
nand U6598 (N_6598,N_6437,N_6005);
nor U6599 (N_6599,N_6392,N_6388);
nand U6600 (N_6600,N_6095,N_6106);
and U6601 (N_6601,N_6443,N_6415);
nand U6602 (N_6602,N_6468,N_6430);
nand U6603 (N_6603,N_6319,N_6252);
and U6604 (N_6604,N_6266,N_6469);
nor U6605 (N_6605,N_6183,N_6122);
nand U6606 (N_6606,N_6004,N_6053);
nor U6607 (N_6607,N_6457,N_6052);
nor U6608 (N_6608,N_6423,N_6057);
nor U6609 (N_6609,N_6151,N_6141);
or U6610 (N_6610,N_6080,N_6375);
nand U6611 (N_6611,N_6006,N_6001);
nand U6612 (N_6612,N_6488,N_6357);
and U6613 (N_6613,N_6283,N_6056);
nor U6614 (N_6614,N_6432,N_6422);
and U6615 (N_6615,N_6203,N_6239);
nand U6616 (N_6616,N_6250,N_6326);
nand U6617 (N_6617,N_6238,N_6017);
or U6618 (N_6618,N_6387,N_6105);
or U6619 (N_6619,N_6480,N_6383);
xnor U6620 (N_6620,N_6411,N_6280);
nand U6621 (N_6621,N_6454,N_6335);
and U6622 (N_6622,N_6366,N_6282);
and U6623 (N_6623,N_6150,N_6261);
or U6624 (N_6624,N_6378,N_6334);
nand U6625 (N_6625,N_6138,N_6002);
and U6626 (N_6626,N_6494,N_6445);
nand U6627 (N_6627,N_6438,N_6031);
or U6628 (N_6628,N_6064,N_6347);
nand U6629 (N_6629,N_6316,N_6175);
and U6630 (N_6630,N_6495,N_6341);
xnor U6631 (N_6631,N_6194,N_6255);
nand U6632 (N_6632,N_6125,N_6493);
xnor U6633 (N_6633,N_6191,N_6224);
nor U6634 (N_6634,N_6132,N_6440);
or U6635 (N_6635,N_6018,N_6418);
nand U6636 (N_6636,N_6253,N_6309);
or U6637 (N_6637,N_6091,N_6331);
or U6638 (N_6638,N_6228,N_6082);
nor U6639 (N_6639,N_6118,N_6113);
and U6640 (N_6640,N_6110,N_6359);
and U6641 (N_6641,N_6305,N_6119);
nor U6642 (N_6642,N_6475,N_6241);
xor U6643 (N_6643,N_6498,N_6441);
nand U6644 (N_6644,N_6107,N_6157);
nand U6645 (N_6645,N_6188,N_6456);
or U6646 (N_6646,N_6160,N_6240);
or U6647 (N_6647,N_6037,N_6166);
nor U6648 (N_6648,N_6259,N_6234);
and U6649 (N_6649,N_6232,N_6436);
or U6650 (N_6650,N_6279,N_6086);
and U6651 (N_6651,N_6075,N_6287);
or U6652 (N_6652,N_6431,N_6306);
nand U6653 (N_6653,N_6213,N_6399);
or U6654 (N_6654,N_6311,N_6289);
nor U6655 (N_6655,N_6327,N_6214);
nor U6656 (N_6656,N_6172,N_6473);
or U6657 (N_6657,N_6070,N_6078);
and U6658 (N_6658,N_6449,N_6087);
nand U6659 (N_6659,N_6063,N_6263);
nand U6660 (N_6660,N_6116,N_6130);
xnor U6661 (N_6661,N_6323,N_6066);
or U6662 (N_6662,N_6458,N_6201);
nand U6663 (N_6663,N_6024,N_6140);
nor U6664 (N_6664,N_6434,N_6146);
and U6665 (N_6665,N_6196,N_6254);
nand U6666 (N_6666,N_6479,N_6049);
nor U6667 (N_6667,N_6258,N_6470);
nand U6668 (N_6668,N_6393,N_6065);
or U6669 (N_6669,N_6094,N_6257);
nand U6670 (N_6670,N_6168,N_6097);
or U6671 (N_6671,N_6154,N_6062);
nand U6672 (N_6672,N_6173,N_6134);
or U6673 (N_6673,N_6189,N_6483);
nand U6674 (N_6674,N_6215,N_6020);
or U6675 (N_6675,N_6424,N_6071);
nor U6676 (N_6676,N_6073,N_6083);
and U6677 (N_6677,N_6439,N_6405);
nand U6678 (N_6678,N_6184,N_6195);
and U6679 (N_6679,N_6197,N_6472);
and U6680 (N_6680,N_6307,N_6451);
xnor U6681 (N_6681,N_6340,N_6312);
nor U6682 (N_6682,N_6284,N_6120);
nand U6683 (N_6683,N_6021,N_6491);
nand U6684 (N_6684,N_6212,N_6428);
nand U6685 (N_6685,N_6389,N_6103);
nand U6686 (N_6686,N_6149,N_6269);
or U6687 (N_6687,N_6251,N_6028);
or U6688 (N_6688,N_6476,N_6332);
nor U6689 (N_6689,N_6058,N_6060);
nand U6690 (N_6690,N_6142,N_6047);
nand U6691 (N_6691,N_6487,N_6310);
xor U6692 (N_6692,N_6462,N_6444);
nor U6693 (N_6693,N_6045,N_6156);
or U6694 (N_6694,N_6354,N_6242);
nand U6695 (N_6695,N_6381,N_6303);
xnor U6696 (N_6696,N_6433,N_6223);
nand U6697 (N_6697,N_6221,N_6112);
or U6698 (N_6698,N_6054,N_6127);
and U6699 (N_6699,N_6216,N_6465);
nand U6700 (N_6700,N_6019,N_6270);
nor U6701 (N_6701,N_6273,N_6300);
nor U6702 (N_6702,N_6425,N_6176);
xor U6703 (N_6703,N_6464,N_6274);
and U6704 (N_6704,N_6012,N_6348);
nor U6705 (N_6705,N_6245,N_6362);
nor U6706 (N_6706,N_6096,N_6337);
nand U6707 (N_6707,N_6329,N_6452);
and U6708 (N_6708,N_6185,N_6278);
xnor U6709 (N_6709,N_6299,N_6148);
or U6710 (N_6710,N_6209,N_6364);
and U6711 (N_6711,N_6275,N_6244);
or U6712 (N_6712,N_6396,N_6126);
xor U6713 (N_6713,N_6351,N_6429);
xnor U6714 (N_6714,N_6202,N_6369);
xnor U6715 (N_6715,N_6104,N_6463);
nor U6716 (N_6716,N_6471,N_6059);
or U6717 (N_6717,N_6181,N_6489);
nor U6718 (N_6718,N_6350,N_6041);
nand U6719 (N_6719,N_6328,N_6448);
xnor U6720 (N_6720,N_6271,N_6040);
nor U6721 (N_6721,N_6077,N_6374);
nor U6722 (N_6722,N_6165,N_6051);
xor U6723 (N_6723,N_6050,N_6163);
nor U6724 (N_6724,N_6447,N_6330);
and U6725 (N_6725,N_6171,N_6343);
and U6726 (N_6726,N_6026,N_6039);
and U6727 (N_6727,N_6376,N_6067);
nor U6728 (N_6728,N_6200,N_6167);
nand U6729 (N_6729,N_6014,N_6460);
or U6730 (N_6730,N_6256,N_6486);
nor U6731 (N_6731,N_6379,N_6382);
nand U6732 (N_6732,N_6226,N_6192);
nand U6733 (N_6733,N_6016,N_6308);
and U6734 (N_6734,N_6336,N_6161);
and U6735 (N_6735,N_6217,N_6015);
or U6736 (N_6736,N_6453,N_6235);
or U6737 (N_6737,N_6248,N_6338);
nand U6738 (N_6738,N_6035,N_6090);
nand U6739 (N_6739,N_6193,N_6069);
and U6740 (N_6740,N_6231,N_6043);
nor U6741 (N_6741,N_6174,N_6318);
xor U6742 (N_6742,N_6324,N_6317);
nor U6743 (N_6743,N_6121,N_6481);
nor U6744 (N_6744,N_6233,N_6408);
or U6745 (N_6745,N_6218,N_6225);
or U6746 (N_6746,N_6277,N_6490);
nor U6747 (N_6747,N_6044,N_6236);
nor U6748 (N_6748,N_6286,N_6179);
nand U6749 (N_6749,N_6153,N_6230);
or U6750 (N_6750,N_6212,N_6117);
nand U6751 (N_6751,N_6240,N_6132);
xnor U6752 (N_6752,N_6456,N_6458);
or U6753 (N_6753,N_6056,N_6329);
and U6754 (N_6754,N_6253,N_6255);
nor U6755 (N_6755,N_6432,N_6146);
or U6756 (N_6756,N_6262,N_6007);
and U6757 (N_6757,N_6387,N_6441);
nor U6758 (N_6758,N_6296,N_6468);
nor U6759 (N_6759,N_6199,N_6336);
and U6760 (N_6760,N_6336,N_6408);
and U6761 (N_6761,N_6053,N_6173);
nand U6762 (N_6762,N_6480,N_6363);
nor U6763 (N_6763,N_6237,N_6343);
or U6764 (N_6764,N_6239,N_6327);
xnor U6765 (N_6765,N_6472,N_6468);
or U6766 (N_6766,N_6392,N_6325);
or U6767 (N_6767,N_6017,N_6130);
xor U6768 (N_6768,N_6169,N_6369);
nor U6769 (N_6769,N_6013,N_6418);
nor U6770 (N_6770,N_6364,N_6183);
nor U6771 (N_6771,N_6227,N_6146);
nand U6772 (N_6772,N_6333,N_6017);
or U6773 (N_6773,N_6049,N_6231);
nand U6774 (N_6774,N_6234,N_6232);
nand U6775 (N_6775,N_6036,N_6180);
nor U6776 (N_6776,N_6236,N_6027);
and U6777 (N_6777,N_6278,N_6368);
nand U6778 (N_6778,N_6331,N_6246);
nand U6779 (N_6779,N_6116,N_6170);
or U6780 (N_6780,N_6092,N_6295);
xor U6781 (N_6781,N_6245,N_6129);
nand U6782 (N_6782,N_6125,N_6007);
and U6783 (N_6783,N_6258,N_6118);
nor U6784 (N_6784,N_6145,N_6346);
or U6785 (N_6785,N_6160,N_6247);
xnor U6786 (N_6786,N_6440,N_6428);
and U6787 (N_6787,N_6236,N_6067);
nor U6788 (N_6788,N_6446,N_6454);
xnor U6789 (N_6789,N_6187,N_6242);
nor U6790 (N_6790,N_6305,N_6206);
and U6791 (N_6791,N_6143,N_6470);
nor U6792 (N_6792,N_6230,N_6111);
xor U6793 (N_6793,N_6430,N_6220);
or U6794 (N_6794,N_6353,N_6308);
nor U6795 (N_6795,N_6271,N_6416);
nor U6796 (N_6796,N_6482,N_6132);
xor U6797 (N_6797,N_6220,N_6134);
xor U6798 (N_6798,N_6262,N_6166);
or U6799 (N_6799,N_6146,N_6423);
and U6800 (N_6800,N_6488,N_6011);
nor U6801 (N_6801,N_6479,N_6474);
nand U6802 (N_6802,N_6377,N_6418);
or U6803 (N_6803,N_6383,N_6293);
or U6804 (N_6804,N_6318,N_6077);
and U6805 (N_6805,N_6224,N_6125);
or U6806 (N_6806,N_6023,N_6006);
xor U6807 (N_6807,N_6150,N_6137);
nor U6808 (N_6808,N_6471,N_6119);
nor U6809 (N_6809,N_6328,N_6187);
nand U6810 (N_6810,N_6237,N_6410);
or U6811 (N_6811,N_6263,N_6064);
and U6812 (N_6812,N_6061,N_6316);
and U6813 (N_6813,N_6066,N_6118);
nor U6814 (N_6814,N_6373,N_6236);
nor U6815 (N_6815,N_6080,N_6238);
nor U6816 (N_6816,N_6470,N_6006);
nand U6817 (N_6817,N_6465,N_6057);
nor U6818 (N_6818,N_6479,N_6473);
and U6819 (N_6819,N_6174,N_6235);
nor U6820 (N_6820,N_6176,N_6110);
nor U6821 (N_6821,N_6343,N_6215);
nand U6822 (N_6822,N_6405,N_6415);
or U6823 (N_6823,N_6231,N_6155);
nand U6824 (N_6824,N_6174,N_6425);
nand U6825 (N_6825,N_6008,N_6266);
and U6826 (N_6826,N_6470,N_6445);
nor U6827 (N_6827,N_6415,N_6212);
and U6828 (N_6828,N_6034,N_6149);
or U6829 (N_6829,N_6244,N_6455);
or U6830 (N_6830,N_6235,N_6068);
or U6831 (N_6831,N_6274,N_6045);
and U6832 (N_6832,N_6386,N_6403);
nor U6833 (N_6833,N_6242,N_6239);
and U6834 (N_6834,N_6127,N_6106);
or U6835 (N_6835,N_6205,N_6495);
nand U6836 (N_6836,N_6225,N_6418);
nor U6837 (N_6837,N_6212,N_6133);
and U6838 (N_6838,N_6066,N_6003);
or U6839 (N_6839,N_6424,N_6359);
nor U6840 (N_6840,N_6235,N_6058);
or U6841 (N_6841,N_6344,N_6144);
nand U6842 (N_6842,N_6379,N_6008);
and U6843 (N_6843,N_6329,N_6119);
nand U6844 (N_6844,N_6429,N_6026);
or U6845 (N_6845,N_6098,N_6012);
xnor U6846 (N_6846,N_6228,N_6459);
and U6847 (N_6847,N_6189,N_6224);
and U6848 (N_6848,N_6167,N_6041);
nand U6849 (N_6849,N_6337,N_6153);
nor U6850 (N_6850,N_6351,N_6049);
nand U6851 (N_6851,N_6273,N_6464);
or U6852 (N_6852,N_6380,N_6125);
or U6853 (N_6853,N_6138,N_6432);
and U6854 (N_6854,N_6159,N_6420);
or U6855 (N_6855,N_6344,N_6394);
and U6856 (N_6856,N_6372,N_6354);
nand U6857 (N_6857,N_6047,N_6242);
nor U6858 (N_6858,N_6310,N_6214);
nand U6859 (N_6859,N_6347,N_6221);
or U6860 (N_6860,N_6330,N_6060);
xnor U6861 (N_6861,N_6451,N_6170);
nor U6862 (N_6862,N_6417,N_6093);
or U6863 (N_6863,N_6105,N_6389);
and U6864 (N_6864,N_6272,N_6425);
or U6865 (N_6865,N_6340,N_6314);
xnor U6866 (N_6866,N_6193,N_6341);
or U6867 (N_6867,N_6053,N_6243);
or U6868 (N_6868,N_6274,N_6327);
and U6869 (N_6869,N_6373,N_6336);
nor U6870 (N_6870,N_6281,N_6080);
nor U6871 (N_6871,N_6049,N_6128);
or U6872 (N_6872,N_6334,N_6304);
or U6873 (N_6873,N_6360,N_6369);
nor U6874 (N_6874,N_6150,N_6423);
xnor U6875 (N_6875,N_6102,N_6359);
xnor U6876 (N_6876,N_6290,N_6244);
and U6877 (N_6877,N_6189,N_6277);
or U6878 (N_6878,N_6251,N_6103);
and U6879 (N_6879,N_6348,N_6191);
or U6880 (N_6880,N_6454,N_6171);
and U6881 (N_6881,N_6169,N_6477);
or U6882 (N_6882,N_6461,N_6024);
nor U6883 (N_6883,N_6380,N_6383);
or U6884 (N_6884,N_6053,N_6017);
and U6885 (N_6885,N_6306,N_6412);
nor U6886 (N_6886,N_6298,N_6398);
nor U6887 (N_6887,N_6349,N_6397);
or U6888 (N_6888,N_6040,N_6248);
and U6889 (N_6889,N_6059,N_6453);
nand U6890 (N_6890,N_6085,N_6477);
xnor U6891 (N_6891,N_6193,N_6469);
or U6892 (N_6892,N_6204,N_6104);
nor U6893 (N_6893,N_6235,N_6224);
or U6894 (N_6894,N_6282,N_6123);
xor U6895 (N_6895,N_6300,N_6412);
nor U6896 (N_6896,N_6214,N_6155);
nand U6897 (N_6897,N_6470,N_6127);
or U6898 (N_6898,N_6024,N_6243);
nand U6899 (N_6899,N_6371,N_6205);
nor U6900 (N_6900,N_6372,N_6355);
nor U6901 (N_6901,N_6160,N_6261);
nor U6902 (N_6902,N_6456,N_6300);
xnor U6903 (N_6903,N_6451,N_6014);
or U6904 (N_6904,N_6071,N_6034);
nor U6905 (N_6905,N_6337,N_6060);
nor U6906 (N_6906,N_6361,N_6111);
and U6907 (N_6907,N_6383,N_6017);
nand U6908 (N_6908,N_6417,N_6143);
nand U6909 (N_6909,N_6127,N_6323);
or U6910 (N_6910,N_6226,N_6104);
or U6911 (N_6911,N_6246,N_6423);
and U6912 (N_6912,N_6335,N_6314);
nand U6913 (N_6913,N_6113,N_6299);
nand U6914 (N_6914,N_6050,N_6329);
or U6915 (N_6915,N_6028,N_6447);
and U6916 (N_6916,N_6054,N_6107);
xnor U6917 (N_6917,N_6039,N_6351);
xnor U6918 (N_6918,N_6029,N_6373);
nor U6919 (N_6919,N_6401,N_6104);
and U6920 (N_6920,N_6421,N_6488);
or U6921 (N_6921,N_6271,N_6474);
and U6922 (N_6922,N_6379,N_6334);
and U6923 (N_6923,N_6450,N_6175);
and U6924 (N_6924,N_6348,N_6081);
nor U6925 (N_6925,N_6207,N_6032);
or U6926 (N_6926,N_6208,N_6157);
nand U6927 (N_6927,N_6263,N_6337);
nand U6928 (N_6928,N_6485,N_6021);
or U6929 (N_6929,N_6279,N_6139);
nand U6930 (N_6930,N_6227,N_6460);
nand U6931 (N_6931,N_6362,N_6178);
xnor U6932 (N_6932,N_6258,N_6011);
nand U6933 (N_6933,N_6381,N_6470);
or U6934 (N_6934,N_6113,N_6130);
nor U6935 (N_6935,N_6305,N_6098);
nor U6936 (N_6936,N_6138,N_6268);
nand U6937 (N_6937,N_6097,N_6184);
nor U6938 (N_6938,N_6096,N_6407);
nor U6939 (N_6939,N_6125,N_6212);
nand U6940 (N_6940,N_6476,N_6268);
or U6941 (N_6941,N_6077,N_6127);
nand U6942 (N_6942,N_6318,N_6410);
and U6943 (N_6943,N_6462,N_6233);
xnor U6944 (N_6944,N_6481,N_6415);
nor U6945 (N_6945,N_6112,N_6099);
nor U6946 (N_6946,N_6025,N_6441);
or U6947 (N_6947,N_6251,N_6273);
nand U6948 (N_6948,N_6348,N_6004);
or U6949 (N_6949,N_6479,N_6439);
nor U6950 (N_6950,N_6452,N_6201);
or U6951 (N_6951,N_6029,N_6015);
nor U6952 (N_6952,N_6208,N_6192);
and U6953 (N_6953,N_6022,N_6371);
and U6954 (N_6954,N_6491,N_6182);
nor U6955 (N_6955,N_6072,N_6299);
nor U6956 (N_6956,N_6265,N_6086);
and U6957 (N_6957,N_6174,N_6039);
or U6958 (N_6958,N_6442,N_6385);
nor U6959 (N_6959,N_6064,N_6429);
or U6960 (N_6960,N_6456,N_6393);
nor U6961 (N_6961,N_6422,N_6062);
or U6962 (N_6962,N_6289,N_6229);
nor U6963 (N_6963,N_6485,N_6324);
xor U6964 (N_6964,N_6206,N_6381);
xnor U6965 (N_6965,N_6458,N_6019);
and U6966 (N_6966,N_6083,N_6382);
nor U6967 (N_6967,N_6126,N_6136);
nand U6968 (N_6968,N_6134,N_6225);
nand U6969 (N_6969,N_6198,N_6339);
nor U6970 (N_6970,N_6336,N_6275);
nand U6971 (N_6971,N_6282,N_6410);
xor U6972 (N_6972,N_6064,N_6251);
or U6973 (N_6973,N_6140,N_6478);
and U6974 (N_6974,N_6224,N_6498);
and U6975 (N_6975,N_6227,N_6080);
nand U6976 (N_6976,N_6438,N_6489);
or U6977 (N_6977,N_6339,N_6079);
and U6978 (N_6978,N_6481,N_6227);
and U6979 (N_6979,N_6307,N_6265);
nand U6980 (N_6980,N_6248,N_6321);
xnor U6981 (N_6981,N_6057,N_6173);
and U6982 (N_6982,N_6351,N_6459);
and U6983 (N_6983,N_6254,N_6115);
nor U6984 (N_6984,N_6039,N_6321);
nand U6985 (N_6985,N_6023,N_6214);
or U6986 (N_6986,N_6142,N_6126);
and U6987 (N_6987,N_6348,N_6276);
xnor U6988 (N_6988,N_6031,N_6202);
nor U6989 (N_6989,N_6230,N_6090);
and U6990 (N_6990,N_6454,N_6247);
nor U6991 (N_6991,N_6007,N_6187);
or U6992 (N_6992,N_6105,N_6185);
xnor U6993 (N_6993,N_6058,N_6458);
or U6994 (N_6994,N_6318,N_6301);
nand U6995 (N_6995,N_6231,N_6055);
nor U6996 (N_6996,N_6074,N_6299);
and U6997 (N_6997,N_6246,N_6094);
and U6998 (N_6998,N_6471,N_6211);
xor U6999 (N_6999,N_6005,N_6393);
or U7000 (N_7000,N_6918,N_6664);
nand U7001 (N_7001,N_6609,N_6877);
xor U7002 (N_7002,N_6673,N_6981);
or U7003 (N_7003,N_6577,N_6778);
or U7004 (N_7004,N_6995,N_6527);
nor U7005 (N_7005,N_6945,N_6991);
nand U7006 (N_7006,N_6647,N_6696);
nor U7007 (N_7007,N_6815,N_6871);
and U7008 (N_7008,N_6912,N_6741);
and U7009 (N_7009,N_6579,N_6909);
and U7010 (N_7010,N_6888,N_6584);
or U7011 (N_7011,N_6729,N_6785);
nor U7012 (N_7012,N_6800,N_6545);
nand U7013 (N_7013,N_6866,N_6873);
nand U7014 (N_7014,N_6814,N_6801);
and U7015 (N_7015,N_6849,N_6992);
and U7016 (N_7016,N_6964,N_6663);
or U7017 (N_7017,N_6917,N_6575);
or U7018 (N_7018,N_6843,N_6959);
nor U7019 (N_7019,N_6797,N_6723);
nand U7020 (N_7020,N_6513,N_6533);
and U7021 (N_7021,N_6755,N_6896);
or U7022 (N_7022,N_6927,N_6675);
nand U7023 (N_7023,N_6689,N_6530);
nand U7024 (N_7024,N_6998,N_6955);
nand U7025 (N_7025,N_6605,N_6901);
nand U7026 (N_7026,N_6684,N_6744);
or U7027 (N_7027,N_6657,N_6963);
nor U7028 (N_7028,N_6953,N_6733);
and U7029 (N_7029,N_6668,N_6947);
nand U7030 (N_7030,N_6829,N_6523);
nor U7031 (N_7031,N_6769,N_6932);
xor U7032 (N_7032,N_6572,N_6886);
nand U7033 (N_7033,N_6655,N_6772);
and U7034 (N_7034,N_6891,N_6773);
and U7035 (N_7035,N_6948,N_6878);
and U7036 (N_7036,N_6565,N_6789);
nand U7037 (N_7037,N_6712,N_6905);
nor U7038 (N_7038,N_6511,N_6701);
and U7039 (N_7039,N_6682,N_6554);
nor U7040 (N_7040,N_6950,N_6933);
nand U7041 (N_7041,N_6857,N_6784);
and U7042 (N_7042,N_6922,N_6637);
nor U7043 (N_7043,N_6506,N_6699);
and U7044 (N_7044,N_6967,N_6844);
or U7045 (N_7045,N_6792,N_6855);
or U7046 (N_7046,N_6636,N_6706);
nor U7047 (N_7047,N_6553,N_6793);
and U7048 (N_7048,N_6568,N_6621);
nor U7049 (N_7049,N_6898,N_6547);
nand U7050 (N_7050,N_6686,N_6924);
nor U7051 (N_7051,N_6518,N_6975);
nor U7052 (N_7052,N_6560,N_6638);
or U7053 (N_7053,N_6854,N_6830);
or U7054 (N_7054,N_6630,N_6537);
and U7055 (N_7055,N_6810,N_6988);
and U7056 (N_7056,N_6875,N_6550);
or U7057 (N_7057,N_6714,N_6783);
or U7058 (N_7058,N_6786,N_6887);
nand U7059 (N_7059,N_6735,N_6587);
nand U7060 (N_7060,N_6957,N_6951);
xor U7061 (N_7061,N_6526,N_6811);
nor U7062 (N_7062,N_6805,N_6928);
or U7063 (N_7063,N_6987,N_6803);
or U7064 (N_7064,N_6790,N_6881);
nor U7065 (N_7065,N_6678,N_6507);
nand U7066 (N_7066,N_6517,N_6535);
nor U7067 (N_7067,N_6989,N_6916);
and U7068 (N_7068,N_6617,N_6958);
and U7069 (N_7069,N_6763,N_6727);
or U7070 (N_7070,N_6758,N_6962);
xor U7071 (N_7071,N_6685,N_6984);
nand U7072 (N_7072,N_6719,N_6923);
nand U7073 (N_7073,N_6616,N_6704);
nand U7074 (N_7074,N_6892,N_6563);
xnor U7075 (N_7075,N_6850,N_6960);
or U7076 (N_7076,N_6934,N_6653);
nor U7077 (N_7077,N_6721,N_6602);
nand U7078 (N_7078,N_6502,N_6585);
and U7079 (N_7079,N_6574,N_6580);
and U7080 (N_7080,N_6505,N_6831);
and U7081 (N_7081,N_6812,N_6884);
nand U7082 (N_7082,N_6827,N_6645);
and U7083 (N_7083,N_6973,N_6738);
nand U7084 (N_7084,N_6930,N_6557);
or U7085 (N_7085,N_6743,N_6718);
nand U7086 (N_7086,N_6816,N_6650);
nand U7087 (N_7087,N_6571,N_6641);
nor U7088 (N_7088,N_6648,N_6771);
xnor U7089 (N_7089,N_6532,N_6508);
or U7090 (N_7090,N_6819,N_6614);
nand U7091 (N_7091,N_6601,N_6567);
nand U7092 (N_7092,N_6556,N_6509);
and U7093 (N_7093,N_6809,N_6705);
nand U7094 (N_7094,N_6599,N_6749);
nand U7095 (N_7095,N_6525,N_6776);
and U7096 (N_7096,N_6952,N_6848);
nor U7097 (N_7097,N_6627,N_6868);
or U7098 (N_7098,N_6942,N_6745);
or U7099 (N_7099,N_6852,N_6795);
and U7100 (N_7100,N_6551,N_6845);
and U7101 (N_7101,N_6907,N_6536);
or U7102 (N_7102,N_6822,N_6885);
or U7103 (N_7103,N_6693,N_6549);
or U7104 (N_7104,N_6756,N_6658);
xnor U7105 (N_7105,N_6633,N_6543);
nand U7106 (N_7106,N_6608,N_6651);
and U7107 (N_7107,N_6842,N_6739);
nand U7108 (N_7108,N_6654,N_6634);
nand U7109 (N_7109,N_6774,N_6539);
xnor U7110 (N_7110,N_6558,N_6692);
nand U7111 (N_7111,N_6582,N_6826);
nand U7112 (N_7112,N_6725,N_6808);
xor U7113 (N_7113,N_6889,N_6751);
or U7114 (N_7114,N_6703,N_6799);
and U7115 (N_7115,N_6818,N_6902);
nor U7116 (N_7116,N_6593,N_6820);
or U7117 (N_7117,N_6944,N_6761);
and U7118 (N_7118,N_6978,N_6730);
nor U7119 (N_7119,N_6817,N_6644);
xor U7120 (N_7120,N_6669,N_6698);
nand U7121 (N_7121,N_6562,N_6913);
and U7122 (N_7122,N_6969,N_6976);
nand U7123 (N_7123,N_6980,N_6591);
and U7124 (N_7124,N_6846,N_6979);
or U7125 (N_7125,N_6764,N_6639);
nor U7126 (N_7126,N_6629,N_6880);
nor U7127 (N_7127,N_6695,N_6863);
or U7128 (N_7128,N_6697,N_6971);
xnor U7129 (N_7129,N_6643,N_6935);
or U7130 (N_7130,N_6919,N_6997);
nand U7131 (N_7131,N_6676,N_6966);
and U7132 (N_7132,N_6806,N_6956);
or U7133 (N_7133,N_6954,N_6836);
and U7134 (N_7134,N_6595,N_6985);
and U7135 (N_7135,N_6940,N_6710);
or U7136 (N_7136,N_6765,N_6752);
or U7137 (N_7137,N_6623,N_6894);
nand U7138 (N_7138,N_6564,N_6993);
xor U7139 (N_7139,N_6667,N_6807);
nor U7140 (N_7140,N_6740,N_6628);
and U7141 (N_7141,N_6748,N_6972);
and U7142 (N_7142,N_6529,N_6632);
or U7143 (N_7143,N_6690,N_6779);
nor U7144 (N_7144,N_6802,N_6631);
or U7145 (N_7145,N_6824,N_6670);
xor U7146 (N_7146,N_6711,N_6681);
nor U7147 (N_7147,N_6867,N_6770);
and U7148 (N_7148,N_6521,N_6897);
and U7149 (N_7149,N_6534,N_6589);
and U7150 (N_7150,N_6768,N_6757);
nand U7151 (N_7151,N_6840,N_6747);
and U7152 (N_7152,N_6861,N_6780);
nor U7153 (N_7153,N_6538,N_6870);
nor U7154 (N_7154,N_6825,N_6904);
nor U7155 (N_7155,N_6731,N_6833);
nor U7156 (N_7156,N_6970,N_6586);
xnor U7157 (N_7157,N_6679,N_6707);
nor U7158 (N_7158,N_6548,N_6626);
nor U7159 (N_7159,N_6869,N_6754);
and U7160 (N_7160,N_6835,N_6625);
nand U7161 (N_7161,N_6635,N_6804);
nor U7162 (N_7162,N_6569,N_6883);
or U7163 (N_7163,N_6566,N_6921);
and U7164 (N_7164,N_6708,N_6893);
nand U7165 (N_7165,N_6903,N_6908);
nand U7166 (N_7166,N_6618,N_6561);
nand U7167 (N_7167,N_6512,N_6974);
xnor U7168 (N_7168,N_6516,N_6760);
nor U7169 (N_7169,N_6936,N_6750);
nand U7170 (N_7170,N_6968,N_6859);
and U7171 (N_7171,N_6900,N_6914);
and U7172 (N_7172,N_6665,N_6541);
xnor U7173 (N_7173,N_6724,N_6937);
or U7174 (N_7174,N_6662,N_6920);
nand U7175 (N_7175,N_6581,N_6520);
nor U7176 (N_7176,N_6649,N_6990);
nor U7177 (N_7177,N_6911,N_6677);
nand U7178 (N_7178,N_6640,N_6734);
nand U7179 (N_7179,N_6736,N_6965);
or U7180 (N_7180,N_6544,N_6598);
nor U7181 (N_7181,N_6737,N_6588);
or U7182 (N_7182,N_6732,N_6624);
or U7183 (N_7183,N_6943,N_6528);
nor U7184 (N_7184,N_6838,N_6837);
or U7185 (N_7185,N_6746,N_6674);
nand U7186 (N_7186,N_6939,N_6890);
xor U7187 (N_7187,N_6832,N_6941);
or U7188 (N_7188,N_6726,N_6660);
xnor U7189 (N_7189,N_6700,N_6671);
nor U7190 (N_7190,N_6672,N_6879);
or U7191 (N_7191,N_6680,N_6798);
xor U7192 (N_7192,N_6860,N_6994);
xnor U7193 (N_7193,N_6977,N_6821);
or U7194 (N_7194,N_6646,N_6573);
or U7195 (N_7195,N_6504,N_6777);
or U7196 (N_7196,N_6656,N_6555);
and U7197 (N_7197,N_6787,N_6775);
and U7198 (N_7198,N_6552,N_6813);
and U7199 (N_7199,N_6851,N_6862);
and U7200 (N_7200,N_6659,N_6728);
and U7201 (N_7201,N_6753,N_6501);
nand U7202 (N_7202,N_6594,N_6619);
or U7203 (N_7203,N_6864,N_6986);
nor U7204 (N_7204,N_6856,N_6996);
nor U7205 (N_7205,N_6722,N_6620);
nand U7206 (N_7206,N_6666,N_6519);
and U7207 (N_7207,N_6613,N_6961);
nor U7208 (N_7208,N_6503,N_6983);
and U7209 (N_7209,N_6522,N_6874);
or U7210 (N_7210,N_6524,N_6949);
or U7211 (N_7211,N_6823,N_6915);
and U7212 (N_7212,N_6709,N_6578);
or U7213 (N_7213,N_6782,N_6702);
or U7214 (N_7214,N_6570,N_6542);
nand U7215 (N_7215,N_6611,N_6766);
and U7216 (N_7216,N_6759,N_6604);
nor U7217 (N_7217,N_6767,N_6999);
nand U7218 (N_7218,N_6590,N_6847);
nand U7219 (N_7219,N_6938,N_6615);
and U7220 (N_7220,N_6876,N_6683);
nand U7221 (N_7221,N_6694,N_6895);
xor U7222 (N_7222,N_6606,N_6510);
nand U7223 (N_7223,N_6600,N_6791);
nor U7224 (N_7224,N_6717,N_6781);
nand U7225 (N_7225,N_6926,N_6794);
and U7226 (N_7226,N_6853,N_6540);
and U7227 (N_7227,N_6713,N_6622);
nand U7228 (N_7228,N_6931,N_6882);
or U7229 (N_7229,N_6652,N_6906);
and U7230 (N_7230,N_6742,N_6546);
or U7231 (N_7231,N_6796,N_6531);
and U7232 (N_7232,N_6661,N_6607);
nor U7233 (N_7233,N_6910,N_6515);
nor U7234 (N_7234,N_6872,N_6642);
and U7235 (N_7235,N_6715,N_6828);
or U7236 (N_7236,N_6500,N_6982);
nor U7237 (N_7237,N_6946,N_6603);
nand U7238 (N_7238,N_6899,N_6839);
and U7239 (N_7239,N_6865,N_6610);
nand U7240 (N_7240,N_6858,N_6691);
or U7241 (N_7241,N_6612,N_6559);
nand U7242 (N_7242,N_6762,N_6925);
nand U7243 (N_7243,N_6597,N_6688);
or U7244 (N_7244,N_6929,N_6592);
or U7245 (N_7245,N_6514,N_6583);
and U7246 (N_7246,N_6841,N_6788);
nor U7247 (N_7247,N_6576,N_6716);
or U7248 (N_7248,N_6687,N_6720);
or U7249 (N_7249,N_6834,N_6596);
or U7250 (N_7250,N_6883,N_6624);
nor U7251 (N_7251,N_6836,N_6582);
and U7252 (N_7252,N_6665,N_6555);
and U7253 (N_7253,N_6559,N_6846);
and U7254 (N_7254,N_6894,N_6617);
and U7255 (N_7255,N_6753,N_6655);
or U7256 (N_7256,N_6565,N_6910);
or U7257 (N_7257,N_6768,N_6797);
nor U7258 (N_7258,N_6965,N_6501);
nand U7259 (N_7259,N_6710,N_6913);
and U7260 (N_7260,N_6622,N_6920);
or U7261 (N_7261,N_6902,N_6669);
or U7262 (N_7262,N_6666,N_6549);
and U7263 (N_7263,N_6621,N_6721);
xnor U7264 (N_7264,N_6759,N_6534);
nor U7265 (N_7265,N_6814,N_6772);
or U7266 (N_7266,N_6784,N_6854);
nor U7267 (N_7267,N_6898,N_6911);
nor U7268 (N_7268,N_6893,N_6522);
and U7269 (N_7269,N_6509,N_6668);
and U7270 (N_7270,N_6812,N_6757);
or U7271 (N_7271,N_6704,N_6580);
or U7272 (N_7272,N_6782,N_6745);
and U7273 (N_7273,N_6932,N_6981);
or U7274 (N_7274,N_6586,N_6593);
and U7275 (N_7275,N_6832,N_6577);
or U7276 (N_7276,N_6818,N_6850);
and U7277 (N_7277,N_6995,N_6560);
and U7278 (N_7278,N_6523,N_6895);
or U7279 (N_7279,N_6946,N_6767);
xnor U7280 (N_7280,N_6725,N_6718);
nand U7281 (N_7281,N_6889,N_6676);
nand U7282 (N_7282,N_6645,N_6610);
or U7283 (N_7283,N_6623,N_6858);
or U7284 (N_7284,N_6617,N_6756);
nor U7285 (N_7285,N_6531,N_6756);
nor U7286 (N_7286,N_6581,N_6500);
nand U7287 (N_7287,N_6547,N_6823);
nand U7288 (N_7288,N_6956,N_6795);
and U7289 (N_7289,N_6738,N_6525);
nand U7290 (N_7290,N_6719,N_6505);
and U7291 (N_7291,N_6573,N_6852);
nor U7292 (N_7292,N_6762,N_6988);
nor U7293 (N_7293,N_6710,N_6526);
nand U7294 (N_7294,N_6577,N_6895);
or U7295 (N_7295,N_6615,N_6869);
nand U7296 (N_7296,N_6688,N_6971);
or U7297 (N_7297,N_6552,N_6835);
and U7298 (N_7298,N_6801,N_6942);
or U7299 (N_7299,N_6887,N_6518);
and U7300 (N_7300,N_6752,N_6889);
and U7301 (N_7301,N_6574,N_6922);
or U7302 (N_7302,N_6616,N_6550);
and U7303 (N_7303,N_6589,N_6713);
nor U7304 (N_7304,N_6625,N_6753);
or U7305 (N_7305,N_6586,N_6790);
and U7306 (N_7306,N_6920,N_6957);
and U7307 (N_7307,N_6669,N_6768);
nand U7308 (N_7308,N_6694,N_6812);
nand U7309 (N_7309,N_6818,N_6782);
nand U7310 (N_7310,N_6729,N_6694);
nor U7311 (N_7311,N_6522,N_6617);
nand U7312 (N_7312,N_6756,N_6790);
xor U7313 (N_7313,N_6615,N_6647);
xnor U7314 (N_7314,N_6819,N_6659);
nand U7315 (N_7315,N_6669,N_6503);
or U7316 (N_7316,N_6518,N_6559);
nand U7317 (N_7317,N_6767,N_6894);
or U7318 (N_7318,N_6906,N_6896);
and U7319 (N_7319,N_6725,N_6783);
nand U7320 (N_7320,N_6889,N_6909);
and U7321 (N_7321,N_6668,N_6561);
xor U7322 (N_7322,N_6570,N_6654);
nor U7323 (N_7323,N_6542,N_6941);
or U7324 (N_7324,N_6705,N_6513);
nand U7325 (N_7325,N_6721,N_6941);
and U7326 (N_7326,N_6684,N_6971);
nor U7327 (N_7327,N_6744,N_6892);
and U7328 (N_7328,N_6872,N_6725);
and U7329 (N_7329,N_6504,N_6539);
nor U7330 (N_7330,N_6951,N_6853);
and U7331 (N_7331,N_6532,N_6901);
or U7332 (N_7332,N_6818,N_6726);
nand U7333 (N_7333,N_6660,N_6803);
nand U7334 (N_7334,N_6612,N_6760);
nand U7335 (N_7335,N_6638,N_6550);
xor U7336 (N_7336,N_6830,N_6727);
nor U7337 (N_7337,N_6533,N_6589);
nand U7338 (N_7338,N_6577,N_6730);
nor U7339 (N_7339,N_6938,N_6929);
nand U7340 (N_7340,N_6514,N_6794);
or U7341 (N_7341,N_6880,N_6525);
xnor U7342 (N_7342,N_6977,N_6877);
and U7343 (N_7343,N_6741,N_6680);
xnor U7344 (N_7344,N_6891,N_6840);
nor U7345 (N_7345,N_6739,N_6837);
nand U7346 (N_7346,N_6639,N_6931);
xor U7347 (N_7347,N_6856,N_6863);
nand U7348 (N_7348,N_6787,N_6500);
nand U7349 (N_7349,N_6791,N_6799);
or U7350 (N_7350,N_6853,N_6967);
nand U7351 (N_7351,N_6777,N_6920);
nor U7352 (N_7352,N_6600,N_6576);
and U7353 (N_7353,N_6881,N_6736);
or U7354 (N_7354,N_6538,N_6894);
nand U7355 (N_7355,N_6543,N_6876);
nand U7356 (N_7356,N_6601,N_6643);
nor U7357 (N_7357,N_6618,N_6623);
nor U7358 (N_7358,N_6604,N_6792);
and U7359 (N_7359,N_6983,N_6707);
nor U7360 (N_7360,N_6792,N_6645);
nand U7361 (N_7361,N_6838,N_6637);
and U7362 (N_7362,N_6726,N_6633);
nand U7363 (N_7363,N_6716,N_6981);
or U7364 (N_7364,N_6742,N_6782);
or U7365 (N_7365,N_6516,N_6868);
and U7366 (N_7366,N_6540,N_6709);
and U7367 (N_7367,N_6964,N_6565);
nor U7368 (N_7368,N_6956,N_6732);
nor U7369 (N_7369,N_6699,N_6630);
xor U7370 (N_7370,N_6792,N_6528);
nand U7371 (N_7371,N_6780,N_6881);
nor U7372 (N_7372,N_6673,N_6592);
or U7373 (N_7373,N_6683,N_6692);
and U7374 (N_7374,N_6539,N_6541);
and U7375 (N_7375,N_6632,N_6789);
nor U7376 (N_7376,N_6553,N_6614);
nand U7377 (N_7377,N_6726,N_6727);
and U7378 (N_7378,N_6517,N_6697);
nor U7379 (N_7379,N_6704,N_6971);
nor U7380 (N_7380,N_6692,N_6702);
nand U7381 (N_7381,N_6687,N_6721);
and U7382 (N_7382,N_6972,N_6909);
nand U7383 (N_7383,N_6845,N_6754);
xnor U7384 (N_7384,N_6856,N_6889);
nand U7385 (N_7385,N_6900,N_6799);
nand U7386 (N_7386,N_6580,N_6958);
or U7387 (N_7387,N_6503,N_6751);
nand U7388 (N_7388,N_6914,N_6593);
nor U7389 (N_7389,N_6722,N_6660);
nor U7390 (N_7390,N_6960,N_6841);
or U7391 (N_7391,N_6504,N_6523);
nor U7392 (N_7392,N_6922,N_6631);
nand U7393 (N_7393,N_6702,N_6913);
nand U7394 (N_7394,N_6654,N_6738);
nor U7395 (N_7395,N_6542,N_6668);
and U7396 (N_7396,N_6985,N_6716);
or U7397 (N_7397,N_6886,N_6520);
or U7398 (N_7398,N_6838,N_6684);
nand U7399 (N_7399,N_6960,N_6764);
xor U7400 (N_7400,N_6927,N_6924);
nor U7401 (N_7401,N_6884,N_6651);
nor U7402 (N_7402,N_6895,N_6801);
or U7403 (N_7403,N_6695,N_6631);
nor U7404 (N_7404,N_6659,N_6591);
and U7405 (N_7405,N_6756,N_6500);
or U7406 (N_7406,N_6708,N_6876);
xnor U7407 (N_7407,N_6670,N_6580);
or U7408 (N_7408,N_6570,N_6738);
and U7409 (N_7409,N_6503,N_6532);
and U7410 (N_7410,N_6648,N_6862);
nor U7411 (N_7411,N_6585,N_6867);
or U7412 (N_7412,N_6998,N_6898);
nand U7413 (N_7413,N_6663,N_6557);
and U7414 (N_7414,N_6989,N_6738);
or U7415 (N_7415,N_6502,N_6637);
nor U7416 (N_7416,N_6619,N_6521);
or U7417 (N_7417,N_6758,N_6743);
or U7418 (N_7418,N_6720,N_6678);
nand U7419 (N_7419,N_6794,N_6716);
nor U7420 (N_7420,N_6741,N_6746);
or U7421 (N_7421,N_6668,N_6886);
nand U7422 (N_7422,N_6531,N_6524);
and U7423 (N_7423,N_6952,N_6500);
nor U7424 (N_7424,N_6688,N_6980);
or U7425 (N_7425,N_6798,N_6756);
xor U7426 (N_7426,N_6726,N_6744);
xor U7427 (N_7427,N_6648,N_6715);
nor U7428 (N_7428,N_6969,N_6619);
nor U7429 (N_7429,N_6697,N_6655);
nand U7430 (N_7430,N_6975,N_6627);
or U7431 (N_7431,N_6745,N_6556);
nor U7432 (N_7432,N_6964,N_6584);
and U7433 (N_7433,N_6599,N_6787);
nand U7434 (N_7434,N_6799,N_6885);
nor U7435 (N_7435,N_6706,N_6619);
nor U7436 (N_7436,N_6959,N_6934);
or U7437 (N_7437,N_6799,N_6877);
nand U7438 (N_7438,N_6788,N_6755);
or U7439 (N_7439,N_6879,N_6614);
or U7440 (N_7440,N_6509,N_6792);
and U7441 (N_7441,N_6862,N_6545);
nand U7442 (N_7442,N_6971,N_6870);
and U7443 (N_7443,N_6515,N_6582);
nor U7444 (N_7444,N_6630,N_6719);
and U7445 (N_7445,N_6543,N_6975);
and U7446 (N_7446,N_6975,N_6644);
nand U7447 (N_7447,N_6883,N_6714);
or U7448 (N_7448,N_6896,N_6978);
nor U7449 (N_7449,N_6761,N_6914);
nor U7450 (N_7450,N_6624,N_6910);
or U7451 (N_7451,N_6681,N_6963);
nand U7452 (N_7452,N_6572,N_6540);
and U7453 (N_7453,N_6817,N_6776);
nand U7454 (N_7454,N_6948,N_6866);
nor U7455 (N_7455,N_6969,N_6985);
nor U7456 (N_7456,N_6671,N_6793);
or U7457 (N_7457,N_6931,N_6633);
nor U7458 (N_7458,N_6638,N_6644);
nor U7459 (N_7459,N_6512,N_6664);
nor U7460 (N_7460,N_6914,N_6920);
nor U7461 (N_7461,N_6980,N_6891);
nand U7462 (N_7462,N_6510,N_6523);
or U7463 (N_7463,N_6760,N_6733);
or U7464 (N_7464,N_6560,N_6958);
nand U7465 (N_7465,N_6685,N_6737);
nor U7466 (N_7466,N_6999,N_6826);
nand U7467 (N_7467,N_6967,N_6835);
or U7468 (N_7468,N_6860,N_6501);
xnor U7469 (N_7469,N_6999,N_6990);
nand U7470 (N_7470,N_6674,N_6657);
and U7471 (N_7471,N_6551,N_6780);
nor U7472 (N_7472,N_6658,N_6996);
and U7473 (N_7473,N_6577,N_6620);
or U7474 (N_7474,N_6583,N_6555);
nand U7475 (N_7475,N_6605,N_6681);
nor U7476 (N_7476,N_6877,N_6631);
nor U7477 (N_7477,N_6837,N_6806);
nor U7478 (N_7478,N_6988,N_6784);
xnor U7479 (N_7479,N_6849,N_6525);
xor U7480 (N_7480,N_6809,N_6982);
or U7481 (N_7481,N_6914,N_6510);
nor U7482 (N_7482,N_6832,N_6684);
nand U7483 (N_7483,N_6734,N_6511);
nor U7484 (N_7484,N_6563,N_6650);
nor U7485 (N_7485,N_6500,N_6623);
and U7486 (N_7486,N_6917,N_6748);
or U7487 (N_7487,N_6555,N_6823);
and U7488 (N_7488,N_6794,N_6924);
nor U7489 (N_7489,N_6626,N_6975);
xor U7490 (N_7490,N_6549,N_6877);
nand U7491 (N_7491,N_6711,N_6658);
or U7492 (N_7492,N_6870,N_6983);
nand U7493 (N_7493,N_6525,N_6500);
xor U7494 (N_7494,N_6968,N_6574);
and U7495 (N_7495,N_6827,N_6852);
nand U7496 (N_7496,N_6964,N_6875);
nand U7497 (N_7497,N_6572,N_6546);
or U7498 (N_7498,N_6702,N_6940);
nand U7499 (N_7499,N_6561,N_6514);
nand U7500 (N_7500,N_7219,N_7418);
and U7501 (N_7501,N_7319,N_7065);
or U7502 (N_7502,N_7133,N_7161);
and U7503 (N_7503,N_7461,N_7062);
or U7504 (N_7504,N_7046,N_7211);
or U7505 (N_7505,N_7198,N_7378);
nand U7506 (N_7506,N_7263,N_7075);
or U7507 (N_7507,N_7450,N_7489);
nor U7508 (N_7508,N_7283,N_7366);
nand U7509 (N_7509,N_7138,N_7428);
nor U7510 (N_7510,N_7475,N_7312);
and U7511 (N_7511,N_7324,N_7376);
or U7512 (N_7512,N_7496,N_7383);
and U7513 (N_7513,N_7302,N_7371);
nor U7514 (N_7514,N_7020,N_7479);
or U7515 (N_7515,N_7206,N_7273);
nor U7516 (N_7516,N_7003,N_7192);
nand U7517 (N_7517,N_7305,N_7044);
or U7518 (N_7518,N_7245,N_7420);
or U7519 (N_7519,N_7403,N_7149);
and U7520 (N_7520,N_7370,N_7117);
nand U7521 (N_7521,N_7226,N_7317);
nor U7522 (N_7522,N_7099,N_7181);
nand U7523 (N_7523,N_7431,N_7089);
nand U7524 (N_7524,N_7325,N_7369);
nor U7525 (N_7525,N_7147,N_7224);
or U7526 (N_7526,N_7018,N_7393);
xor U7527 (N_7527,N_7104,N_7172);
xnor U7528 (N_7528,N_7010,N_7021);
and U7529 (N_7529,N_7126,N_7222);
nand U7530 (N_7530,N_7372,N_7173);
and U7531 (N_7531,N_7063,N_7085);
and U7532 (N_7532,N_7377,N_7237);
or U7533 (N_7533,N_7308,N_7114);
or U7534 (N_7534,N_7110,N_7436);
nand U7535 (N_7535,N_7462,N_7073);
or U7536 (N_7536,N_7130,N_7470);
or U7537 (N_7537,N_7332,N_7122);
nand U7538 (N_7538,N_7105,N_7338);
and U7539 (N_7539,N_7427,N_7412);
or U7540 (N_7540,N_7129,N_7053);
and U7541 (N_7541,N_7035,N_7477);
or U7542 (N_7542,N_7030,N_7251);
nor U7543 (N_7543,N_7004,N_7002);
nand U7544 (N_7544,N_7280,N_7180);
nor U7545 (N_7545,N_7070,N_7025);
xnor U7546 (N_7546,N_7042,N_7109);
and U7547 (N_7547,N_7398,N_7112);
and U7548 (N_7548,N_7438,N_7026);
nand U7549 (N_7549,N_7357,N_7084);
nand U7550 (N_7550,N_7405,N_7417);
or U7551 (N_7551,N_7024,N_7353);
xor U7552 (N_7552,N_7032,N_7210);
nor U7553 (N_7553,N_7054,N_7297);
and U7554 (N_7554,N_7497,N_7118);
nor U7555 (N_7555,N_7277,N_7135);
nand U7556 (N_7556,N_7080,N_7086);
nor U7557 (N_7557,N_7387,N_7472);
or U7558 (N_7558,N_7242,N_7052);
nand U7559 (N_7559,N_7231,N_7166);
and U7560 (N_7560,N_7127,N_7334);
nand U7561 (N_7561,N_7270,N_7364);
nor U7562 (N_7562,N_7336,N_7047);
nor U7563 (N_7563,N_7131,N_7490);
and U7564 (N_7564,N_7139,N_7234);
nor U7565 (N_7565,N_7410,N_7184);
xnor U7566 (N_7566,N_7223,N_7300);
or U7567 (N_7567,N_7386,N_7485);
and U7568 (N_7568,N_7456,N_7159);
nor U7569 (N_7569,N_7352,N_7156);
nand U7570 (N_7570,N_7011,N_7392);
and U7571 (N_7571,N_7027,N_7136);
nor U7572 (N_7572,N_7401,N_7137);
nand U7573 (N_7573,N_7066,N_7097);
or U7574 (N_7574,N_7039,N_7186);
or U7575 (N_7575,N_7205,N_7426);
or U7576 (N_7576,N_7441,N_7487);
nand U7577 (N_7577,N_7228,N_7215);
and U7578 (N_7578,N_7279,N_7335);
nor U7579 (N_7579,N_7077,N_7200);
xnor U7580 (N_7580,N_7266,N_7028);
nand U7581 (N_7581,N_7278,N_7008);
or U7582 (N_7582,N_7061,N_7292);
nand U7583 (N_7583,N_7408,N_7390);
and U7584 (N_7584,N_7145,N_7082);
and U7585 (N_7585,N_7433,N_7079);
xor U7586 (N_7586,N_7007,N_7351);
nand U7587 (N_7587,N_7471,N_7113);
or U7588 (N_7588,N_7288,N_7177);
or U7589 (N_7589,N_7102,N_7217);
xnor U7590 (N_7590,N_7261,N_7255);
nor U7591 (N_7591,N_7074,N_7329);
nor U7592 (N_7592,N_7191,N_7321);
xnor U7593 (N_7593,N_7394,N_7482);
xor U7594 (N_7594,N_7264,N_7094);
and U7595 (N_7595,N_7157,N_7058);
or U7596 (N_7596,N_7246,N_7256);
xnor U7597 (N_7597,N_7252,N_7221);
and U7598 (N_7598,N_7388,N_7121);
nor U7599 (N_7599,N_7328,N_7214);
nand U7600 (N_7600,N_7488,N_7285);
xnor U7601 (N_7601,N_7259,N_7434);
nand U7602 (N_7602,N_7049,N_7313);
xnor U7603 (N_7603,N_7402,N_7385);
nor U7604 (N_7604,N_7171,N_7415);
or U7605 (N_7605,N_7142,N_7384);
nand U7606 (N_7606,N_7148,N_7009);
nand U7607 (N_7607,N_7204,N_7038);
nor U7608 (N_7608,N_7195,N_7268);
nor U7609 (N_7609,N_7060,N_7269);
xnor U7610 (N_7610,N_7474,N_7150);
nand U7611 (N_7611,N_7216,N_7006);
nand U7612 (N_7612,N_7484,N_7330);
and U7613 (N_7613,N_7048,N_7345);
and U7614 (N_7614,N_7340,N_7407);
or U7615 (N_7615,N_7001,N_7233);
nor U7616 (N_7616,N_7153,N_7416);
and U7617 (N_7617,N_7344,N_7301);
xor U7618 (N_7618,N_7187,N_7341);
or U7619 (N_7619,N_7454,N_7014);
nand U7620 (N_7620,N_7476,N_7435);
or U7621 (N_7621,N_7404,N_7017);
nand U7622 (N_7622,N_7419,N_7276);
or U7623 (N_7623,N_7493,N_7031);
nor U7624 (N_7624,N_7466,N_7023);
nand U7625 (N_7625,N_7355,N_7037);
or U7626 (N_7626,N_7169,N_7498);
nor U7627 (N_7627,N_7446,N_7125);
nand U7628 (N_7628,N_7499,N_7422);
and U7629 (N_7629,N_7076,N_7162);
nand U7630 (N_7630,N_7019,N_7381);
nor U7631 (N_7631,N_7087,N_7414);
nor U7632 (N_7632,N_7144,N_7347);
or U7633 (N_7633,N_7314,N_7421);
nand U7634 (N_7634,N_7111,N_7247);
and U7635 (N_7635,N_7123,N_7342);
and U7636 (N_7636,N_7323,N_7449);
and U7637 (N_7637,N_7391,N_7185);
and U7638 (N_7638,N_7348,N_7289);
nor U7639 (N_7639,N_7440,N_7235);
nand U7640 (N_7640,N_7067,N_7120);
nor U7641 (N_7641,N_7473,N_7178);
and U7642 (N_7642,N_7069,N_7349);
and U7643 (N_7643,N_7068,N_7430);
xor U7644 (N_7644,N_7107,N_7309);
nand U7645 (N_7645,N_7170,N_7101);
nor U7646 (N_7646,N_7453,N_7190);
and U7647 (N_7647,N_7005,N_7363);
or U7648 (N_7648,N_7424,N_7360);
nand U7649 (N_7649,N_7194,N_7400);
nand U7650 (N_7650,N_7163,N_7158);
or U7651 (N_7651,N_7483,N_7096);
nor U7652 (N_7652,N_7059,N_7298);
xnor U7653 (N_7653,N_7197,N_7250);
nand U7654 (N_7654,N_7088,N_7165);
or U7655 (N_7655,N_7304,N_7209);
nand U7656 (N_7656,N_7439,N_7128);
nor U7657 (N_7657,N_7100,N_7208);
xnor U7658 (N_7658,N_7152,N_7103);
and U7659 (N_7659,N_7199,N_7365);
and U7660 (N_7660,N_7327,N_7282);
nand U7661 (N_7661,N_7457,N_7480);
nor U7662 (N_7662,N_7290,N_7459);
nand U7663 (N_7663,N_7220,N_7106);
nor U7664 (N_7664,N_7124,N_7468);
xnor U7665 (N_7665,N_7154,N_7098);
and U7666 (N_7666,N_7310,N_7445);
nand U7667 (N_7667,N_7249,N_7262);
or U7668 (N_7668,N_7193,N_7202);
or U7669 (N_7669,N_7458,N_7492);
nor U7670 (N_7670,N_7116,N_7443);
nand U7671 (N_7671,N_7093,N_7397);
or U7672 (N_7672,N_7040,N_7429);
xnor U7673 (N_7673,N_7240,N_7322);
and U7674 (N_7674,N_7016,N_7326);
nand U7675 (N_7675,N_7375,N_7463);
and U7676 (N_7676,N_7295,N_7411);
nor U7677 (N_7677,N_7465,N_7146);
or U7678 (N_7678,N_7469,N_7333);
nor U7679 (N_7679,N_7346,N_7167);
or U7680 (N_7680,N_7361,N_7013);
and U7681 (N_7681,N_7367,N_7248);
and U7682 (N_7682,N_7423,N_7239);
nor U7683 (N_7683,N_7083,N_7207);
and U7684 (N_7684,N_7265,N_7291);
xor U7685 (N_7685,N_7115,N_7160);
xor U7686 (N_7686,N_7307,N_7274);
nor U7687 (N_7687,N_7303,N_7389);
nand U7688 (N_7688,N_7486,N_7442);
and U7689 (N_7689,N_7294,N_7331);
and U7690 (N_7690,N_7022,N_7119);
nor U7691 (N_7691,N_7225,N_7481);
nand U7692 (N_7692,N_7132,N_7081);
nand U7693 (N_7693,N_7232,N_7271);
nand U7694 (N_7694,N_7033,N_7241);
and U7695 (N_7695,N_7437,N_7238);
nor U7696 (N_7696,N_7293,N_7141);
nand U7697 (N_7697,N_7337,N_7164);
and U7698 (N_7698,N_7258,N_7350);
or U7699 (N_7699,N_7380,N_7451);
nor U7700 (N_7700,N_7374,N_7359);
nand U7701 (N_7701,N_7396,N_7034);
nand U7702 (N_7702,N_7196,N_7299);
and U7703 (N_7703,N_7409,N_7444);
nor U7704 (N_7704,N_7036,N_7368);
nor U7705 (N_7705,N_7108,N_7078);
and U7706 (N_7706,N_7236,N_7201);
or U7707 (N_7707,N_7212,N_7000);
nor U7708 (N_7708,N_7091,N_7316);
nand U7709 (N_7709,N_7494,N_7203);
or U7710 (N_7710,N_7179,N_7406);
and U7711 (N_7711,N_7092,N_7151);
or U7712 (N_7712,N_7296,N_7286);
or U7713 (N_7713,N_7029,N_7467);
nand U7714 (N_7714,N_7358,N_7315);
nor U7715 (N_7715,N_7455,N_7213);
or U7716 (N_7716,N_7399,N_7343);
and U7717 (N_7717,N_7218,N_7043);
nor U7718 (N_7718,N_7050,N_7311);
nor U7719 (N_7719,N_7071,N_7257);
nor U7720 (N_7720,N_7318,N_7460);
nor U7721 (N_7721,N_7055,N_7056);
or U7722 (N_7722,N_7281,N_7267);
and U7723 (N_7723,N_7495,N_7176);
and U7724 (N_7724,N_7095,N_7287);
nand U7725 (N_7725,N_7143,N_7064);
nand U7726 (N_7726,N_7373,N_7272);
xor U7727 (N_7727,N_7057,N_7432);
xnor U7728 (N_7728,N_7188,N_7354);
and U7729 (N_7729,N_7254,N_7362);
and U7730 (N_7730,N_7072,N_7452);
nor U7731 (N_7731,N_7413,N_7425);
or U7732 (N_7732,N_7379,N_7230);
or U7733 (N_7733,N_7491,N_7448);
nand U7734 (N_7734,N_7140,N_7041);
nand U7735 (N_7735,N_7183,N_7478);
nand U7736 (N_7736,N_7339,N_7244);
nand U7737 (N_7737,N_7447,N_7382);
and U7738 (N_7738,N_7284,N_7253);
xor U7739 (N_7739,N_7260,N_7174);
xor U7740 (N_7740,N_7015,N_7134);
or U7741 (N_7741,N_7182,N_7175);
and U7742 (N_7742,N_7395,N_7012);
nand U7743 (N_7743,N_7320,N_7356);
nor U7744 (N_7744,N_7090,N_7051);
nand U7745 (N_7745,N_7189,N_7275);
nor U7746 (N_7746,N_7229,N_7155);
and U7747 (N_7747,N_7168,N_7045);
nand U7748 (N_7748,N_7243,N_7227);
or U7749 (N_7749,N_7464,N_7306);
nand U7750 (N_7750,N_7455,N_7277);
and U7751 (N_7751,N_7074,N_7108);
or U7752 (N_7752,N_7309,N_7451);
nand U7753 (N_7753,N_7412,N_7174);
nand U7754 (N_7754,N_7336,N_7454);
and U7755 (N_7755,N_7487,N_7270);
nand U7756 (N_7756,N_7465,N_7162);
nor U7757 (N_7757,N_7053,N_7399);
or U7758 (N_7758,N_7335,N_7250);
and U7759 (N_7759,N_7499,N_7492);
and U7760 (N_7760,N_7255,N_7009);
or U7761 (N_7761,N_7294,N_7481);
nand U7762 (N_7762,N_7014,N_7330);
or U7763 (N_7763,N_7244,N_7478);
xnor U7764 (N_7764,N_7240,N_7375);
or U7765 (N_7765,N_7466,N_7490);
xor U7766 (N_7766,N_7296,N_7241);
or U7767 (N_7767,N_7039,N_7025);
nor U7768 (N_7768,N_7172,N_7206);
or U7769 (N_7769,N_7407,N_7006);
nor U7770 (N_7770,N_7328,N_7003);
or U7771 (N_7771,N_7087,N_7277);
and U7772 (N_7772,N_7471,N_7200);
and U7773 (N_7773,N_7437,N_7393);
nand U7774 (N_7774,N_7068,N_7186);
nor U7775 (N_7775,N_7000,N_7389);
nor U7776 (N_7776,N_7263,N_7459);
xnor U7777 (N_7777,N_7240,N_7074);
nor U7778 (N_7778,N_7049,N_7058);
nand U7779 (N_7779,N_7159,N_7119);
xor U7780 (N_7780,N_7245,N_7317);
nand U7781 (N_7781,N_7187,N_7116);
and U7782 (N_7782,N_7098,N_7081);
xnor U7783 (N_7783,N_7085,N_7067);
xor U7784 (N_7784,N_7238,N_7053);
xor U7785 (N_7785,N_7199,N_7247);
and U7786 (N_7786,N_7496,N_7446);
nand U7787 (N_7787,N_7244,N_7381);
nand U7788 (N_7788,N_7412,N_7342);
nand U7789 (N_7789,N_7386,N_7199);
nand U7790 (N_7790,N_7145,N_7383);
nand U7791 (N_7791,N_7394,N_7245);
and U7792 (N_7792,N_7131,N_7324);
or U7793 (N_7793,N_7310,N_7305);
nand U7794 (N_7794,N_7061,N_7100);
and U7795 (N_7795,N_7328,N_7261);
and U7796 (N_7796,N_7427,N_7325);
and U7797 (N_7797,N_7298,N_7282);
nor U7798 (N_7798,N_7123,N_7361);
and U7799 (N_7799,N_7094,N_7493);
and U7800 (N_7800,N_7108,N_7194);
xor U7801 (N_7801,N_7468,N_7157);
nand U7802 (N_7802,N_7129,N_7377);
and U7803 (N_7803,N_7038,N_7200);
and U7804 (N_7804,N_7086,N_7004);
or U7805 (N_7805,N_7155,N_7160);
and U7806 (N_7806,N_7140,N_7390);
nor U7807 (N_7807,N_7482,N_7222);
and U7808 (N_7808,N_7204,N_7375);
xnor U7809 (N_7809,N_7187,N_7195);
or U7810 (N_7810,N_7458,N_7228);
nand U7811 (N_7811,N_7024,N_7262);
nor U7812 (N_7812,N_7329,N_7058);
and U7813 (N_7813,N_7469,N_7252);
nand U7814 (N_7814,N_7080,N_7027);
xor U7815 (N_7815,N_7259,N_7457);
nor U7816 (N_7816,N_7370,N_7135);
or U7817 (N_7817,N_7433,N_7114);
and U7818 (N_7818,N_7063,N_7082);
and U7819 (N_7819,N_7291,N_7454);
nand U7820 (N_7820,N_7139,N_7059);
and U7821 (N_7821,N_7383,N_7297);
or U7822 (N_7822,N_7453,N_7441);
nand U7823 (N_7823,N_7025,N_7423);
nor U7824 (N_7824,N_7288,N_7312);
nand U7825 (N_7825,N_7274,N_7496);
nand U7826 (N_7826,N_7220,N_7041);
xor U7827 (N_7827,N_7228,N_7358);
nor U7828 (N_7828,N_7316,N_7202);
nand U7829 (N_7829,N_7097,N_7282);
nor U7830 (N_7830,N_7460,N_7436);
xnor U7831 (N_7831,N_7401,N_7158);
and U7832 (N_7832,N_7389,N_7235);
or U7833 (N_7833,N_7498,N_7335);
or U7834 (N_7834,N_7263,N_7006);
xnor U7835 (N_7835,N_7078,N_7321);
nor U7836 (N_7836,N_7056,N_7217);
nor U7837 (N_7837,N_7411,N_7182);
xor U7838 (N_7838,N_7320,N_7255);
xnor U7839 (N_7839,N_7269,N_7148);
and U7840 (N_7840,N_7131,N_7049);
or U7841 (N_7841,N_7391,N_7106);
xnor U7842 (N_7842,N_7223,N_7100);
and U7843 (N_7843,N_7423,N_7142);
nand U7844 (N_7844,N_7023,N_7055);
nand U7845 (N_7845,N_7314,N_7344);
nor U7846 (N_7846,N_7096,N_7412);
or U7847 (N_7847,N_7354,N_7056);
and U7848 (N_7848,N_7440,N_7483);
or U7849 (N_7849,N_7402,N_7031);
or U7850 (N_7850,N_7307,N_7293);
nand U7851 (N_7851,N_7305,N_7060);
xor U7852 (N_7852,N_7244,N_7136);
and U7853 (N_7853,N_7116,N_7036);
nor U7854 (N_7854,N_7108,N_7493);
nand U7855 (N_7855,N_7050,N_7256);
nor U7856 (N_7856,N_7049,N_7255);
and U7857 (N_7857,N_7001,N_7303);
nand U7858 (N_7858,N_7117,N_7129);
nor U7859 (N_7859,N_7363,N_7374);
and U7860 (N_7860,N_7203,N_7244);
nand U7861 (N_7861,N_7394,N_7363);
nand U7862 (N_7862,N_7417,N_7156);
nor U7863 (N_7863,N_7146,N_7088);
and U7864 (N_7864,N_7312,N_7317);
nor U7865 (N_7865,N_7454,N_7308);
or U7866 (N_7866,N_7052,N_7164);
or U7867 (N_7867,N_7102,N_7404);
nor U7868 (N_7868,N_7276,N_7359);
nor U7869 (N_7869,N_7431,N_7497);
nand U7870 (N_7870,N_7131,N_7214);
nand U7871 (N_7871,N_7115,N_7184);
and U7872 (N_7872,N_7018,N_7466);
or U7873 (N_7873,N_7408,N_7248);
nand U7874 (N_7874,N_7028,N_7093);
and U7875 (N_7875,N_7092,N_7432);
nand U7876 (N_7876,N_7085,N_7193);
and U7877 (N_7877,N_7419,N_7008);
xor U7878 (N_7878,N_7308,N_7222);
or U7879 (N_7879,N_7239,N_7262);
and U7880 (N_7880,N_7422,N_7384);
nor U7881 (N_7881,N_7215,N_7101);
or U7882 (N_7882,N_7484,N_7481);
and U7883 (N_7883,N_7394,N_7202);
nand U7884 (N_7884,N_7086,N_7304);
nand U7885 (N_7885,N_7051,N_7311);
nand U7886 (N_7886,N_7124,N_7316);
nand U7887 (N_7887,N_7441,N_7262);
and U7888 (N_7888,N_7066,N_7318);
or U7889 (N_7889,N_7416,N_7497);
xor U7890 (N_7890,N_7316,N_7397);
nor U7891 (N_7891,N_7165,N_7281);
xor U7892 (N_7892,N_7459,N_7180);
and U7893 (N_7893,N_7252,N_7149);
or U7894 (N_7894,N_7325,N_7399);
or U7895 (N_7895,N_7044,N_7200);
nand U7896 (N_7896,N_7416,N_7302);
or U7897 (N_7897,N_7428,N_7012);
or U7898 (N_7898,N_7316,N_7452);
xnor U7899 (N_7899,N_7383,N_7180);
nand U7900 (N_7900,N_7243,N_7314);
nand U7901 (N_7901,N_7473,N_7039);
nand U7902 (N_7902,N_7117,N_7029);
or U7903 (N_7903,N_7406,N_7084);
nand U7904 (N_7904,N_7087,N_7033);
nand U7905 (N_7905,N_7476,N_7373);
or U7906 (N_7906,N_7084,N_7089);
xnor U7907 (N_7907,N_7070,N_7403);
nand U7908 (N_7908,N_7099,N_7233);
and U7909 (N_7909,N_7339,N_7361);
nor U7910 (N_7910,N_7330,N_7256);
nor U7911 (N_7911,N_7414,N_7358);
nand U7912 (N_7912,N_7428,N_7290);
nor U7913 (N_7913,N_7337,N_7300);
and U7914 (N_7914,N_7154,N_7129);
xor U7915 (N_7915,N_7488,N_7408);
or U7916 (N_7916,N_7241,N_7092);
nor U7917 (N_7917,N_7343,N_7272);
and U7918 (N_7918,N_7464,N_7109);
nor U7919 (N_7919,N_7363,N_7316);
or U7920 (N_7920,N_7187,N_7356);
or U7921 (N_7921,N_7377,N_7227);
nor U7922 (N_7922,N_7048,N_7222);
nand U7923 (N_7923,N_7417,N_7127);
nand U7924 (N_7924,N_7058,N_7401);
or U7925 (N_7925,N_7443,N_7414);
or U7926 (N_7926,N_7275,N_7244);
or U7927 (N_7927,N_7394,N_7092);
and U7928 (N_7928,N_7402,N_7217);
and U7929 (N_7929,N_7201,N_7347);
xor U7930 (N_7930,N_7121,N_7074);
nor U7931 (N_7931,N_7112,N_7322);
or U7932 (N_7932,N_7245,N_7361);
nor U7933 (N_7933,N_7417,N_7318);
and U7934 (N_7934,N_7385,N_7082);
and U7935 (N_7935,N_7498,N_7324);
and U7936 (N_7936,N_7183,N_7493);
or U7937 (N_7937,N_7155,N_7370);
nand U7938 (N_7938,N_7424,N_7052);
nor U7939 (N_7939,N_7337,N_7364);
or U7940 (N_7940,N_7252,N_7196);
xnor U7941 (N_7941,N_7435,N_7304);
nor U7942 (N_7942,N_7220,N_7094);
or U7943 (N_7943,N_7108,N_7162);
nor U7944 (N_7944,N_7120,N_7011);
nand U7945 (N_7945,N_7064,N_7490);
and U7946 (N_7946,N_7442,N_7463);
nand U7947 (N_7947,N_7086,N_7063);
xnor U7948 (N_7948,N_7150,N_7172);
or U7949 (N_7949,N_7024,N_7043);
or U7950 (N_7950,N_7162,N_7286);
or U7951 (N_7951,N_7360,N_7290);
nand U7952 (N_7952,N_7421,N_7136);
nor U7953 (N_7953,N_7359,N_7207);
nor U7954 (N_7954,N_7338,N_7111);
xnor U7955 (N_7955,N_7038,N_7131);
nor U7956 (N_7956,N_7353,N_7364);
nor U7957 (N_7957,N_7485,N_7409);
xnor U7958 (N_7958,N_7031,N_7097);
nor U7959 (N_7959,N_7443,N_7311);
nor U7960 (N_7960,N_7149,N_7264);
nor U7961 (N_7961,N_7324,N_7074);
nand U7962 (N_7962,N_7418,N_7163);
xor U7963 (N_7963,N_7178,N_7072);
and U7964 (N_7964,N_7194,N_7079);
nor U7965 (N_7965,N_7196,N_7400);
nor U7966 (N_7966,N_7363,N_7182);
or U7967 (N_7967,N_7412,N_7470);
or U7968 (N_7968,N_7381,N_7332);
nand U7969 (N_7969,N_7108,N_7215);
and U7970 (N_7970,N_7248,N_7243);
nand U7971 (N_7971,N_7123,N_7487);
and U7972 (N_7972,N_7376,N_7272);
nand U7973 (N_7973,N_7462,N_7112);
xnor U7974 (N_7974,N_7391,N_7259);
nand U7975 (N_7975,N_7211,N_7166);
nor U7976 (N_7976,N_7002,N_7407);
nor U7977 (N_7977,N_7485,N_7287);
nand U7978 (N_7978,N_7451,N_7320);
and U7979 (N_7979,N_7286,N_7279);
or U7980 (N_7980,N_7445,N_7480);
nand U7981 (N_7981,N_7101,N_7192);
nor U7982 (N_7982,N_7127,N_7110);
or U7983 (N_7983,N_7311,N_7484);
nand U7984 (N_7984,N_7474,N_7329);
and U7985 (N_7985,N_7138,N_7406);
and U7986 (N_7986,N_7372,N_7116);
and U7987 (N_7987,N_7018,N_7115);
and U7988 (N_7988,N_7138,N_7236);
nor U7989 (N_7989,N_7087,N_7203);
nand U7990 (N_7990,N_7038,N_7203);
and U7991 (N_7991,N_7041,N_7435);
and U7992 (N_7992,N_7071,N_7042);
and U7993 (N_7993,N_7499,N_7322);
or U7994 (N_7994,N_7117,N_7368);
xor U7995 (N_7995,N_7275,N_7466);
nand U7996 (N_7996,N_7467,N_7425);
and U7997 (N_7997,N_7092,N_7497);
nand U7998 (N_7998,N_7438,N_7308);
or U7999 (N_7999,N_7253,N_7101);
or U8000 (N_8000,N_7882,N_7955);
or U8001 (N_8001,N_7585,N_7934);
nand U8002 (N_8002,N_7986,N_7869);
and U8003 (N_8003,N_7818,N_7687);
nand U8004 (N_8004,N_7633,N_7973);
nor U8005 (N_8005,N_7914,N_7651);
or U8006 (N_8006,N_7681,N_7948);
nor U8007 (N_8007,N_7971,N_7965);
or U8008 (N_8008,N_7957,N_7501);
and U8009 (N_8009,N_7755,N_7577);
nor U8010 (N_8010,N_7552,N_7580);
and U8011 (N_8011,N_7686,N_7921);
or U8012 (N_8012,N_7613,N_7677);
xor U8013 (N_8013,N_7944,N_7834);
xor U8014 (N_8014,N_7622,N_7930);
or U8015 (N_8015,N_7983,N_7823);
nor U8016 (N_8016,N_7674,N_7855);
and U8017 (N_8017,N_7516,N_7586);
xnor U8018 (N_8018,N_7806,N_7964);
nor U8019 (N_8019,N_7842,N_7984);
and U8020 (N_8020,N_7660,N_7940);
nand U8021 (N_8021,N_7993,N_7549);
nand U8022 (N_8022,N_7989,N_7551);
nand U8023 (N_8023,N_7545,N_7511);
nand U8024 (N_8024,N_7919,N_7562);
and U8025 (N_8025,N_7630,N_7859);
or U8026 (N_8026,N_7659,N_7889);
and U8027 (N_8027,N_7550,N_7891);
nand U8028 (N_8028,N_7902,N_7900);
and U8029 (N_8029,N_7694,N_7669);
and U8030 (N_8030,N_7915,N_7893);
and U8031 (N_8031,N_7932,N_7801);
and U8032 (N_8032,N_7715,N_7839);
and U8033 (N_8033,N_7627,N_7726);
or U8034 (N_8034,N_7979,N_7877);
nand U8035 (N_8035,N_7556,N_7961);
xnor U8036 (N_8036,N_7596,N_7739);
and U8037 (N_8037,N_7590,N_7904);
nor U8038 (N_8038,N_7609,N_7638);
nand U8039 (N_8039,N_7758,N_7886);
nor U8040 (N_8040,N_7679,N_7820);
or U8041 (N_8041,N_7935,N_7897);
xnor U8042 (N_8042,N_7720,N_7746);
and U8043 (N_8043,N_7636,N_7794);
nand U8044 (N_8044,N_7606,N_7525);
or U8045 (N_8045,N_7733,N_7647);
and U8046 (N_8046,N_7863,N_7532);
nand U8047 (N_8047,N_7872,N_7673);
nor U8048 (N_8048,N_7512,N_7728);
nand U8049 (N_8049,N_7905,N_7643);
nand U8050 (N_8050,N_7831,N_7527);
nand U8051 (N_8051,N_7724,N_7535);
nor U8052 (N_8052,N_7721,N_7587);
nand U8053 (N_8053,N_7712,N_7560);
or U8054 (N_8054,N_7765,N_7582);
or U8055 (N_8055,N_7785,N_7817);
nand U8056 (N_8056,N_7888,N_7798);
nand U8057 (N_8057,N_7608,N_7907);
nor U8058 (N_8058,N_7639,N_7812);
xor U8059 (N_8059,N_7774,N_7773);
xnor U8060 (N_8060,N_7941,N_7786);
nor U8061 (N_8061,N_7929,N_7602);
nor U8062 (N_8062,N_7953,N_7916);
xnor U8063 (N_8063,N_7998,N_7994);
or U8064 (N_8064,N_7912,N_7943);
or U8065 (N_8065,N_7578,N_7951);
and U8066 (N_8066,N_7620,N_7777);
or U8067 (N_8067,N_7665,N_7780);
or U8068 (N_8068,N_7672,N_7736);
xnor U8069 (N_8069,N_7753,N_7604);
nor U8070 (N_8070,N_7830,N_7650);
or U8071 (N_8071,N_7621,N_7561);
or U8072 (N_8072,N_7901,N_7959);
nor U8073 (N_8073,N_7533,N_7652);
nand U8074 (N_8074,N_7624,N_7862);
or U8075 (N_8075,N_7750,N_7937);
nor U8076 (N_8076,N_7866,N_7970);
nor U8077 (N_8077,N_7543,N_7908);
and U8078 (N_8078,N_7837,N_7748);
and U8079 (N_8079,N_7529,N_7641);
nor U8080 (N_8080,N_7827,N_7895);
or U8081 (N_8081,N_7565,N_7824);
nor U8082 (N_8082,N_7734,N_7988);
nor U8083 (N_8083,N_7534,N_7685);
nand U8084 (N_8084,N_7832,N_7506);
and U8085 (N_8085,N_7816,N_7729);
nand U8086 (N_8086,N_7992,N_7789);
nor U8087 (N_8087,N_7642,N_7693);
nand U8088 (N_8088,N_7595,N_7689);
nand U8089 (N_8089,N_7962,N_7514);
and U8090 (N_8090,N_7705,N_7795);
or U8091 (N_8091,N_7661,N_7709);
or U8092 (N_8092,N_7883,N_7942);
nor U8093 (N_8093,N_7803,N_7851);
nand U8094 (N_8094,N_7909,N_7711);
nand U8095 (N_8095,N_7960,N_7519);
or U8096 (N_8096,N_7749,N_7890);
and U8097 (N_8097,N_7509,N_7884);
xnor U8098 (N_8098,N_7618,N_7683);
and U8099 (N_8099,N_7635,N_7626);
and U8100 (N_8100,N_7822,N_7526);
or U8101 (N_8101,N_7975,N_7978);
and U8102 (N_8102,N_7906,N_7745);
and U8103 (N_8103,N_7579,N_7808);
nor U8104 (N_8104,N_7878,N_7564);
nand U8105 (N_8105,N_7787,N_7566);
or U8106 (N_8106,N_7881,N_7927);
xor U8107 (N_8107,N_7778,N_7852);
and U8108 (N_8108,N_7713,N_7903);
nand U8109 (N_8109,N_7697,N_7847);
or U8110 (N_8110,N_7860,N_7744);
and U8111 (N_8111,N_7968,N_7597);
and U8112 (N_8112,N_7856,N_7696);
or U8113 (N_8113,N_7528,N_7864);
nor U8114 (N_8114,N_7503,N_7548);
and U8115 (N_8115,N_7783,N_7771);
xnor U8116 (N_8116,N_7563,N_7536);
nand U8117 (N_8117,N_7699,N_7631);
and U8118 (N_8118,N_7688,N_7594);
and U8119 (N_8119,N_7751,N_7956);
xnor U8120 (N_8120,N_7767,N_7576);
or U8121 (N_8121,N_7896,N_7876);
or U8122 (N_8122,N_7592,N_7663);
nand U8123 (N_8123,N_7880,N_7752);
nand U8124 (N_8124,N_7658,N_7531);
or U8125 (N_8125,N_7518,N_7719);
and U8126 (N_8126,N_7938,N_7702);
or U8127 (N_8127,N_7589,N_7737);
nor U8128 (N_8128,N_7911,N_7857);
or U8129 (N_8129,N_7571,N_7504);
nand U8130 (N_8130,N_7850,N_7646);
nor U8131 (N_8131,N_7980,N_7985);
xor U8132 (N_8132,N_7871,N_7928);
or U8133 (N_8133,N_7873,N_7949);
nor U8134 (N_8134,N_7969,N_7678);
nand U8135 (N_8135,N_7568,N_7813);
nor U8136 (N_8136,N_7867,N_7990);
and U8137 (N_8137,N_7807,N_7861);
or U8138 (N_8138,N_7547,N_7800);
nand U8139 (N_8139,N_7792,N_7700);
xor U8140 (N_8140,N_7634,N_7917);
or U8141 (N_8141,N_7858,N_7649);
nand U8142 (N_8142,N_7682,N_7603);
and U8143 (N_8143,N_7828,N_7524);
and U8144 (N_8144,N_7797,N_7840);
xor U8145 (N_8145,N_7982,N_7553);
and U8146 (N_8146,N_7657,N_7763);
nand U8147 (N_8147,N_7821,N_7781);
nor U8148 (N_8148,N_7987,N_7799);
nor U8149 (N_8149,N_7588,N_7574);
and U8150 (N_8150,N_7698,N_7544);
nor U8151 (N_8151,N_7865,N_7796);
nor U8152 (N_8152,N_7950,N_7601);
or U8153 (N_8153,N_7567,N_7833);
and U8154 (N_8154,N_7841,N_7757);
nand U8155 (N_8155,N_7653,N_7887);
nor U8156 (N_8156,N_7760,N_7946);
nand U8157 (N_8157,N_7999,N_7868);
nand U8158 (N_8158,N_7676,N_7542);
nor U8159 (N_8159,N_7769,N_7605);
nand U8160 (N_8160,N_7584,N_7735);
nand U8161 (N_8161,N_7967,N_7540);
and U8162 (N_8162,N_7836,N_7617);
nand U8163 (N_8163,N_7684,N_7913);
nand U8164 (N_8164,N_7616,N_7637);
nor U8165 (N_8165,N_7575,N_7537);
xnor U8166 (N_8166,N_7559,N_7809);
or U8167 (N_8167,N_7510,N_7926);
or U8168 (N_8168,N_7591,N_7879);
nor U8169 (N_8169,N_7569,N_7522);
nor U8170 (N_8170,N_7885,N_7614);
nor U8171 (N_8171,N_7716,N_7838);
and U8172 (N_8172,N_7931,N_7936);
nor U8173 (N_8173,N_7875,N_7600);
or U8174 (N_8174,N_7958,N_7762);
and U8175 (N_8175,N_7654,N_7593);
nand U8176 (N_8176,N_7977,N_7554);
and U8177 (N_8177,N_7619,N_7668);
and U8178 (N_8178,N_7599,N_7991);
nor U8179 (N_8179,N_7640,N_7725);
xnor U8180 (N_8180,N_7732,N_7695);
nand U8181 (N_8181,N_7628,N_7632);
or U8182 (N_8182,N_7513,N_7692);
nor U8183 (N_8183,N_7925,N_7826);
or U8184 (N_8184,N_7764,N_7945);
or U8185 (N_8185,N_7517,N_7804);
and U8186 (N_8186,N_7558,N_7500);
nor U8187 (N_8187,N_7502,N_7741);
or U8188 (N_8188,N_7662,N_7811);
xor U8189 (N_8189,N_7790,N_7963);
nor U8190 (N_8190,N_7756,N_7680);
or U8191 (N_8191,N_7843,N_7974);
nand U8192 (N_8192,N_7788,N_7775);
and U8193 (N_8193,N_7910,N_7848);
xor U8194 (N_8194,N_7874,N_7920);
nor U8195 (N_8195,N_7710,N_7546);
nand U8196 (N_8196,N_7829,N_7976);
and U8197 (N_8197,N_7644,N_7555);
nand U8198 (N_8198,N_7708,N_7611);
nand U8199 (N_8199,N_7723,N_7899);
nand U8200 (N_8200,N_7924,N_7784);
or U8201 (N_8201,N_7623,N_7667);
nor U8202 (N_8202,N_7581,N_7718);
nor U8203 (N_8203,N_7598,N_7505);
nand U8204 (N_8204,N_7731,N_7759);
or U8205 (N_8205,N_7922,N_7791);
xor U8206 (N_8206,N_7814,N_7520);
and U8207 (N_8207,N_7738,N_7704);
or U8208 (N_8208,N_7761,N_7648);
nor U8209 (N_8209,N_7523,N_7810);
nor U8210 (N_8210,N_7918,N_7671);
nand U8211 (N_8211,N_7612,N_7703);
and U8212 (N_8212,N_7573,N_7655);
and U8213 (N_8213,N_7530,N_7538);
nand U8214 (N_8214,N_7894,N_7572);
nand U8215 (N_8215,N_7701,N_7779);
and U8216 (N_8216,N_7815,N_7892);
nand U8217 (N_8217,N_7666,N_7521);
nor U8218 (N_8218,N_7997,N_7583);
and U8219 (N_8219,N_7768,N_7947);
or U8220 (N_8220,N_7742,N_7670);
or U8221 (N_8221,N_7570,N_7766);
nor U8222 (N_8222,N_7727,N_7656);
nand U8223 (N_8223,N_7996,N_7966);
and U8224 (N_8224,N_7845,N_7747);
nand U8225 (N_8225,N_7690,N_7933);
nand U8226 (N_8226,N_7849,N_7691);
nor U8227 (N_8227,N_7972,N_7995);
xor U8228 (N_8228,N_7923,N_7870);
nand U8229 (N_8229,N_7557,N_7740);
nor U8230 (N_8230,N_7770,N_7782);
nand U8231 (N_8231,N_7898,N_7615);
nor U8232 (N_8232,N_7706,N_7776);
nand U8233 (N_8233,N_7853,N_7981);
and U8234 (N_8234,N_7664,N_7754);
or U8235 (N_8235,N_7707,N_7846);
nor U8236 (N_8236,N_7645,N_7629);
and U8237 (N_8237,N_7939,N_7772);
nor U8238 (N_8238,N_7625,N_7515);
and U8239 (N_8239,N_7730,N_7805);
or U8240 (N_8240,N_7835,N_7714);
nor U8241 (N_8241,N_7952,N_7541);
nor U8242 (N_8242,N_7743,N_7825);
nand U8243 (N_8243,N_7610,N_7722);
or U8244 (N_8244,N_7607,N_7954);
nand U8245 (N_8245,N_7854,N_7793);
nand U8246 (N_8246,N_7539,N_7717);
xor U8247 (N_8247,N_7508,N_7844);
or U8248 (N_8248,N_7819,N_7507);
nand U8249 (N_8249,N_7802,N_7675);
xor U8250 (N_8250,N_7941,N_7540);
nor U8251 (N_8251,N_7695,N_7767);
nor U8252 (N_8252,N_7687,N_7767);
nor U8253 (N_8253,N_7780,N_7845);
nor U8254 (N_8254,N_7883,N_7930);
or U8255 (N_8255,N_7649,N_7945);
and U8256 (N_8256,N_7810,N_7653);
and U8257 (N_8257,N_7881,N_7891);
nor U8258 (N_8258,N_7594,N_7957);
and U8259 (N_8259,N_7759,N_7954);
or U8260 (N_8260,N_7655,N_7895);
and U8261 (N_8261,N_7649,N_7902);
or U8262 (N_8262,N_7904,N_7960);
nand U8263 (N_8263,N_7922,N_7988);
and U8264 (N_8264,N_7755,N_7925);
xnor U8265 (N_8265,N_7955,N_7972);
xnor U8266 (N_8266,N_7784,N_7854);
nand U8267 (N_8267,N_7502,N_7656);
or U8268 (N_8268,N_7599,N_7704);
nor U8269 (N_8269,N_7699,N_7866);
nand U8270 (N_8270,N_7695,N_7821);
or U8271 (N_8271,N_7698,N_7594);
or U8272 (N_8272,N_7903,N_7902);
nand U8273 (N_8273,N_7996,N_7730);
and U8274 (N_8274,N_7773,N_7534);
nor U8275 (N_8275,N_7943,N_7748);
nand U8276 (N_8276,N_7504,N_7764);
nor U8277 (N_8277,N_7522,N_7533);
and U8278 (N_8278,N_7705,N_7728);
and U8279 (N_8279,N_7715,N_7597);
and U8280 (N_8280,N_7721,N_7507);
or U8281 (N_8281,N_7821,N_7571);
and U8282 (N_8282,N_7939,N_7849);
nand U8283 (N_8283,N_7712,N_7940);
and U8284 (N_8284,N_7808,N_7944);
and U8285 (N_8285,N_7750,N_7510);
nor U8286 (N_8286,N_7965,N_7813);
nor U8287 (N_8287,N_7514,N_7863);
or U8288 (N_8288,N_7667,N_7579);
or U8289 (N_8289,N_7603,N_7770);
nor U8290 (N_8290,N_7794,N_7779);
or U8291 (N_8291,N_7942,N_7652);
or U8292 (N_8292,N_7799,N_7755);
nand U8293 (N_8293,N_7850,N_7633);
or U8294 (N_8294,N_7793,N_7654);
nor U8295 (N_8295,N_7742,N_7949);
nor U8296 (N_8296,N_7742,N_7811);
and U8297 (N_8297,N_7974,N_7838);
or U8298 (N_8298,N_7888,N_7773);
and U8299 (N_8299,N_7808,N_7825);
nor U8300 (N_8300,N_7785,N_7917);
nor U8301 (N_8301,N_7934,N_7550);
nand U8302 (N_8302,N_7671,N_7628);
or U8303 (N_8303,N_7802,N_7889);
nand U8304 (N_8304,N_7547,N_7692);
nor U8305 (N_8305,N_7636,N_7873);
nor U8306 (N_8306,N_7579,N_7535);
xor U8307 (N_8307,N_7969,N_7535);
xor U8308 (N_8308,N_7894,N_7978);
nand U8309 (N_8309,N_7839,N_7759);
and U8310 (N_8310,N_7998,N_7640);
xnor U8311 (N_8311,N_7857,N_7873);
or U8312 (N_8312,N_7743,N_7786);
nand U8313 (N_8313,N_7894,N_7563);
nand U8314 (N_8314,N_7770,N_7999);
or U8315 (N_8315,N_7525,N_7727);
or U8316 (N_8316,N_7888,N_7538);
or U8317 (N_8317,N_7545,N_7746);
or U8318 (N_8318,N_7789,N_7760);
or U8319 (N_8319,N_7502,N_7568);
or U8320 (N_8320,N_7841,N_7531);
or U8321 (N_8321,N_7708,N_7675);
nand U8322 (N_8322,N_7670,N_7615);
xnor U8323 (N_8323,N_7679,N_7824);
and U8324 (N_8324,N_7632,N_7870);
nand U8325 (N_8325,N_7945,N_7765);
or U8326 (N_8326,N_7664,N_7899);
or U8327 (N_8327,N_7780,N_7835);
nor U8328 (N_8328,N_7702,N_7694);
xor U8329 (N_8329,N_7821,N_7635);
nor U8330 (N_8330,N_7925,N_7511);
nand U8331 (N_8331,N_7997,N_7983);
nor U8332 (N_8332,N_7901,N_7759);
nand U8333 (N_8333,N_7611,N_7770);
or U8334 (N_8334,N_7679,N_7507);
or U8335 (N_8335,N_7613,N_7521);
and U8336 (N_8336,N_7718,N_7549);
or U8337 (N_8337,N_7939,N_7639);
or U8338 (N_8338,N_7651,N_7622);
nand U8339 (N_8339,N_7768,N_7697);
xnor U8340 (N_8340,N_7796,N_7586);
or U8341 (N_8341,N_7824,N_7673);
or U8342 (N_8342,N_7779,N_7813);
and U8343 (N_8343,N_7691,N_7760);
and U8344 (N_8344,N_7613,N_7660);
nor U8345 (N_8345,N_7754,N_7717);
and U8346 (N_8346,N_7957,N_7504);
or U8347 (N_8347,N_7772,N_7944);
nand U8348 (N_8348,N_7594,N_7510);
or U8349 (N_8349,N_7605,N_7872);
or U8350 (N_8350,N_7575,N_7776);
nor U8351 (N_8351,N_7765,N_7612);
and U8352 (N_8352,N_7752,N_7911);
nor U8353 (N_8353,N_7933,N_7801);
xnor U8354 (N_8354,N_7558,N_7568);
xor U8355 (N_8355,N_7618,N_7847);
nor U8356 (N_8356,N_7648,N_7651);
xnor U8357 (N_8357,N_7963,N_7788);
nor U8358 (N_8358,N_7528,N_7712);
and U8359 (N_8359,N_7913,N_7826);
nand U8360 (N_8360,N_7690,N_7963);
and U8361 (N_8361,N_7585,N_7867);
and U8362 (N_8362,N_7689,N_7520);
nor U8363 (N_8363,N_7526,N_7624);
nand U8364 (N_8364,N_7991,N_7595);
nand U8365 (N_8365,N_7737,N_7684);
or U8366 (N_8366,N_7702,N_7557);
nor U8367 (N_8367,N_7633,N_7913);
or U8368 (N_8368,N_7576,N_7634);
and U8369 (N_8369,N_7622,N_7667);
or U8370 (N_8370,N_7856,N_7707);
nor U8371 (N_8371,N_7586,N_7513);
xnor U8372 (N_8372,N_7908,N_7707);
nor U8373 (N_8373,N_7739,N_7754);
nor U8374 (N_8374,N_7896,N_7905);
nor U8375 (N_8375,N_7631,N_7851);
and U8376 (N_8376,N_7610,N_7876);
and U8377 (N_8377,N_7583,N_7594);
nand U8378 (N_8378,N_7654,N_7649);
nand U8379 (N_8379,N_7515,N_7815);
or U8380 (N_8380,N_7622,N_7806);
xor U8381 (N_8381,N_7633,N_7793);
xnor U8382 (N_8382,N_7799,N_7566);
or U8383 (N_8383,N_7562,N_7913);
or U8384 (N_8384,N_7844,N_7522);
and U8385 (N_8385,N_7546,N_7972);
nor U8386 (N_8386,N_7677,N_7698);
xor U8387 (N_8387,N_7717,N_7948);
or U8388 (N_8388,N_7789,N_7896);
nand U8389 (N_8389,N_7777,N_7955);
or U8390 (N_8390,N_7675,N_7922);
nor U8391 (N_8391,N_7644,N_7508);
nor U8392 (N_8392,N_7743,N_7980);
xor U8393 (N_8393,N_7888,N_7792);
nand U8394 (N_8394,N_7879,N_7734);
nand U8395 (N_8395,N_7796,N_7760);
xor U8396 (N_8396,N_7613,N_7967);
xnor U8397 (N_8397,N_7928,N_7757);
nand U8398 (N_8398,N_7614,N_7552);
xnor U8399 (N_8399,N_7855,N_7996);
nor U8400 (N_8400,N_7857,N_7872);
nand U8401 (N_8401,N_7515,N_7611);
or U8402 (N_8402,N_7766,N_7614);
nand U8403 (N_8403,N_7597,N_7751);
nand U8404 (N_8404,N_7679,N_7626);
and U8405 (N_8405,N_7598,N_7576);
xnor U8406 (N_8406,N_7999,N_7605);
nand U8407 (N_8407,N_7857,N_7953);
or U8408 (N_8408,N_7744,N_7500);
nand U8409 (N_8409,N_7984,N_7823);
or U8410 (N_8410,N_7946,N_7877);
and U8411 (N_8411,N_7654,N_7621);
xnor U8412 (N_8412,N_7736,N_7601);
nand U8413 (N_8413,N_7648,N_7942);
and U8414 (N_8414,N_7859,N_7970);
and U8415 (N_8415,N_7906,N_7778);
and U8416 (N_8416,N_7985,N_7737);
nand U8417 (N_8417,N_7899,N_7749);
nand U8418 (N_8418,N_7565,N_7625);
nor U8419 (N_8419,N_7941,N_7999);
nor U8420 (N_8420,N_7688,N_7743);
and U8421 (N_8421,N_7702,N_7882);
nor U8422 (N_8422,N_7693,N_7746);
nand U8423 (N_8423,N_7538,N_7976);
or U8424 (N_8424,N_7853,N_7891);
and U8425 (N_8425,N_7625,N_7893);
nor U8426 (N_8426,N_7689,N_7967);
nor U8427 (N_8427,N_7788,N_7637);
or U8428 (N_8428,N_7785,N_7542);
nor U8429 (N_8429,N_7949,N_7830);
or U8430 (N_8430,N_7777,N_7662);
nand U8431 (N_8431,N_7972,N_7754);
and U8432 (N_8432,N_7949,N_7876);
nor U8433 (N_8433,N_7895,N_7872);
or U8434 (N_8434,N_7825,N_7919);
xor U8435 (N_8435,N_7735,N_7553);
or U8436 (N_8436,N_7813,N_7897);
and U8437 (N_8437,N_7901,N_7718);
or U8438 (N_8438,N_7861,N_7840);
or U8439 (N_8439,N_7955,N_7907);
and U8440 (N_8440,N_7917,N_7824);
xnor U8441 (N_8441,N_7541,N_7857);
nand U8442 (N_8442,N_7886,N_7770);
nor U8443 (N_8443,N_7530,N_7894);
and U8444 (N_8444,N_7637,N_7900);
nand U8445 (N_8445,N_7687,N_7936);
nand U8446 (N_8446,N_7623,N_7508);
and U8447 (N_8447,N_7676,N_7896);
nor U8448 (N_8448,N_7947,N_7603);
nor U8449 (N_8449,N_7865,N_7579);
nor U8450 (N_8450,N_7774,N_7543);
nand U8451 (N_8451,N_7807,N_7699);
or U8452 (N_8452,N_7862,N_7774);
nor U8453 (N_8453,N_7994,N_7743);
nor U8454 (N_8454,N_7657,N_7863);
and U8455 (N_8455,N_7975,N_7854);
nand U8456 (N_8456,N_7761,N_7702);
nor U8457 (N_8457,N_7782,N_7531);
nand U8458 (N_8458,N_7611,N_7691);
nor U8459 (N_8459,N_7539,N_7575);
xnor U8460 (N_8460,N_7670,N_7868);
nand U8461 (N_8461,N_7533,N_7638);
nor U8462 (N_8462,N_7695,N_7704);
nand U8463 (N_8463,N_7987,N_7839);
and U8464 (N_8464,N_7587,N_7693);
nand U8465 (N_8465,N_7699,N_7531);
nor U8466 (N_8466,N_7607,N_7975);
and U8467 (N_8467,N_7982,N_7708);
and U8468 (N_8468,N_7801,N_7807);
nand U8469 (N_8469,N_7732,N_7850);
or U8470 (N_8470,N_7959,N_7797);
or U8471 (N_8471,N_7863,N_7678);
nand U8472 (N_8472,N_7769,N_7830);
and U8473 (N_8473,N_7903,N_7792);
nand U8474 (N_8474,N_7552,N_7755);
nand U8475 (N_8475,N_7532,N_7891);
and U8476 (N_8476,N_7715,N_7555);
nor U8477 (N_8477,N_7900,N_7563);
nor U8478 (N_8478,N_7646,N_7506);
and U8479 (N_8479,N_7676,N_7775);
or U8480 (N_8480,N_7544,N_7863);
or U8481 (N_8481,N_7553,N_7740);
nand U8482 (N_8482,N_7644,N_7575);
and U8483 (N_8483,N_7545,N_7860);
nand U8484 (N_8484,N_7617,N_7735);
nor U8485 (N_8485,N_7575,N_7823);
nand U8486 (N_8486,N_7676,N_7693);
or U8487 (N_8487,N_7864,N_7639);
xor U8488 (N_8488,N_7624,N_7584);
or U8489 (N_8489,N_7549,N_7985);
or U8490 (N_8490,N_7899,N_7724);
or U8491 (N_8491,N_7550,N_7561);
nand U8492 (N_8492,N_7999,N_7698);
nor U8493 (N_8493,N_7691,N_7930);
nor U8494 (N_8494,N_7824,N_7885);
and U8495 (N_8495,N_7610,N_7706);
nor U8496 (N_8496,N_7523,N_7740);
nor U8497 (N_8497,N_7923,N_7551);
and U8498 (N_8498,N_7704,N_7643);
xor U8499 (N_8499,N_7772,N_7961);
or U8500 (N_8500,N_8284,N_8214);
or U8501 (N_8501,N_8304,N_8470);
xor U8502 (N_8502,N_8326,N_8142);
and U8503 (N_8503,N_8167,N_8150);
xnor U8504 (N_8504,N_8231,N_8385);
nand U8505 (N_8505,N_8416,N_8067);
xnor U8506 (N_8506,N_8481,N_8082);
and U8507 (N_8507,N_8371,N_8260);
nand U8508 (N_8508,N_8316,N_8406);
and U8509 (N_8509,N_8490,N_8203);
or U8510 (N_8510,N_8084,N_8045);
nand U8511 (N_8511,N_8215,N_8375);
or U8512 (N_8512,N_8110,N_8471);
and U8513 (N_8513,N_8341,N_8468);
nor U8514 (N_8514,N_8227,N_8296);
or U8515 (N_8515,N_8455,N_8223);
nand U8516 (N_8516,N_8016,N_8238);
nand U8517 (N_8517,N_8083,N_8319);
xor U8518 (N_8518,N_8065,N_8099);
nor U8519 (N_8519,N_8415,N_8282);
and U8520 (N_8520,N_8201,N_8002);
or U8521 (N_8521,N_8191,N_8365);
and U8522 (N_8522,N_8262,N_8056);
or U8523 (N_8523,N_8437,N_8448);
nor U8524 (N_8524,N_8176,N_8347);
nand U8525 (N_8525,N_8394,N_8337);
nor U8526 (N_8526,N_8152,N_8332);
nand U8527 (N_8527,N_8410,N_8439);
or U8528 (N_8528,N_8348,N_8087);
nor U8529 (N_8529,N_8333,N_8369);
or U8530 (N_8530,N_8381,N_8431);
or U8531 (N_8531,N_8279,N_8386);
or U8532 (N_8532,N_8270,N_8310);
nor U8533 (N_8533,N_8435,N_8198);
or U8534 (N_8534,N_8117,N_8138);
nor U8535 (N_8535,N_8209,N_8374);
nand U8536 (N_8536,N_8382,N_8104);
nand U8537 (N_8537,N_8389,N_8071);
or U8538 (N_8538,N_8093,N_8392);
or U8539 (N_8539,N_8486,N_8403);
and U8540 (N_8540,N_8004,N_8135);
nand U8541 (N_8541,N_8463,N_8059);
and U8542 (N_8542,N_8302,N_8325);
nor U8543 (N_8543,N_8134,N_8050);
or U8544 (N_8544,N_8060,N_8047);
or U8545 (N_8545,N_8208,N_8048);
nand U8546 (N_8546,N_8131,N_8109);
or U8547 (N_8547,N_8197,N_8465);
nand U8548 (N_8548,N_8009,N_8189);
nor U8549 (N_8549,N_8261,N_8187);
and U8550 (N_8550,N_8088,N_8275);
nor U8551 (N_8551,N_8393,N_8119);
or U8552 (N_8552,N_8021,N_8474);
nand U8553 (N_8553,N_8295,N_8454);
and U8554 (N_8554,N_8165,N_8411);
nand U8555 (N_8555,N_8402,N_8140);
nand U8556 (N_8556,N_8210,N_8200);
or U8557 (N_8557,N_8344,N_8343);
nand U8558 (N_8558,N_8354,N_8268);
or U8559 (N_8559,N_8349,N_8323);
nand U8560 (N_8560,N_8064,N_8230);
nand U8561 (N_8561,N_8440,N_8441);
nand U8562 (N_8562,N_8058,N_8040);
or U8563 (N_8563,N_8383,N_8281);
nor U8564 (N_8564,N_8364,N_8073);
nor U8565 (N_8565,N_8265,N_8405);
nand U8566 (N_8566,N_8467,N_8396);
nand U8567 (N_8567,N_8240,N_8458);
nor U8568 (N_8568,N_8242,N_8428);
and U8569 (N_8569,N_8206,N_8163);
or U8570 (N_8570,N_8130,N_8445);
and U8571 (N_8571,N_8026,N_8070);
nor U8572 (N_8572,N_8054,N_8161);
xnor U8573 (N_8573,N_8185,N_8037);
or U8574 (N_8574,N_8211,N_8317);
nor U8575 (N_8575,N_8379,N_8308);
or U8576 (N_8576,N_8010,N_8311);
and U8577 (N_8577,N_8205,N_8327);
or U8578 (N_8578,N_8178,N_8264);
or U8579 (N_8579,N_8126,N_8247);
nand U8580 (N_8580,N_8464,N_8252);
or U8581 (N_8581,N_8014,N_8100);
nor U8582 (N_8582,N_8487,N_8266);
nand U8583 (N_8583,N_8043,N_8034);
nor U8584 (N_8584,N_8390,N_8409);
and U8585 (N_8585,N_8460,N_8484);
and U8586 (N_8586,N_8235,N_8169);
and U8587 (N_8587,N_8305,N_8062);
nand U8588 (N_8588,N_8340,N_8219);
nor U8589 (N_8589,N_8145,N_8280);
nor U8590 (N_8590,N_8132,N_8444);
and U8591 (N_8591,N_8212,N_8251);
or U8592 (N_8592,N_8388,N_8408);
xor U8593 (N_8593,N_8077,N_8139);
and U8594 (N_8594,N_8233,N_8075);
or U8595 (N_8595,N_8180,N_8494);
nor U8596 (N_8596,N_8186,N_8461);
nor U8597 (N_8597,N_8029,N_8288);
nor U8598 (N_8598,N_8147,N_8477);
nand U8599 (N_8599,N_8286,N_8309);
nand U8600 (N_8600,N_8015,N_8172);
nor U8601 (N_8601,N_8112,N_8220);
or U8602 (N_8602,N_8378,N_8174);
and U8603 (N_8603,N_8051,N_8153);
xor U8604 (N_8604,N_8345,N_8120);
nor U8605 (N_8605,N_8278,N_8063);
and U8606 (N_8606,N_8188,N_8492);
nand U8607 (N_8607,N_8489,N_8194);
and U8608 (N_8608,N_8373,N_8190);
and U8609 (N_8609,N_8417,N_8450);
and U8610 (N_8610,N_8250,N_8496);
nor U8611 (N_8611,N_8272,N_8277);
or U8612 (N_8612,N_8199,N_8245);
and U8613 (N_8613,N_8068,N_8107);
nor U8614 (N_8614,N_8446,N_8336);
or U8615 (N_8615,N_8377,N_8129);
nor U8616 (N_8616,N_8306,N_8006);
or U8617 (N_8617,N_8495,N_8404);
or U8618 (N_8618,N_8241,N_8177);
and U8619 (N_8619,N_8181,N_8222);
or U8620 (N_8620,N_8133,N_8159);
nand U8621 (N_8621,N_8456,N_8207);
nand U8622 (N_8622,N_8384,N_8137);
and U8623 (N_8623,N_8469,N_8475);
and U8624 (N_8624,N_8413,N_8017);
or U8625 (N_8625,N_8228,N_8269);
nor U8626 (N_8626,N_8027,N_8192);
nand U8627 (N_8627,N_8482,N_8274);
nor U8628 (N_8628,N_8234,N_8011);
or U8629 (N_8629,N_8038,N_8196);
and U8630 (N_8630,N_8221,N_8338);
and U8631 (N_8631,N_8401,N_8108);
nand U8632 (N_8632,N_8363,N_8313);
xnor U8633 (N_8633,N_8053,N_8156);
or U8634 (N_8634,N_8438,N_8303);
or U8635 (N_8635,N_8499,N_8483);
or U8636 (N_8636,N_8023,N_8432);
and U8637 (N_8637,N_8273,N_8036);
nand U8638 (N_8638,N_8330,N_8155);
nand U8639 (N_8639,N_8491,N_8294);
nand U8640 (N_8640,N_8125,N_8255);
nor U8641 (N_8641,N_8000,N_8328);
or U8642 (N_8642,N_8044,N_8462);
nand U8643 (N_8643,N_8407,N_8086);
nand U8644 (N_8644,N_8061,N_8287);
xor U8645 (N_8645,N_8442,N_8046);
xnor U8646 (N_8646,N_8158,N_8397);
and U8647 (N_8647,N_8076,N_8168);
xor U8648 (N_8648,N_8368,N_8204);
or U8649 (N_8649,N_8127,N_8113);
nor U8650 (N_8650,N_8019,N_8020);
nand U8651 (N_8651,N_8097,N_8146);
nor U8652 (N_8652,N_8123,N_8078);
and U8653 (N_8653,N_8488,N_8098);
nor U8654 (N_8654,N_8253,N_8193);
nand U8655 (N_8655,N_8380,N_8012);
nand U8656 (N_8656,N_8074,N_8298);
and U8657 (N_8657,N_8069,N_8143);
nand U8658 (N_8658,N_8419,N_8106);
and U8659 (N_8659,N_8018,N_8315);
or U8660 (N_8660,N_8248,N_8128);
or U8661 (N_8661,N_8182,N_8451);
nand U8662 (N_8662,N_8285,N_8149);
nand U8663 (N_8663,N_8370,N_8160);
nand U8664 (N_8664,N_8425,N_8144);
nor U8665 (N_8665,N_8094,N_8299);
and U8666 (N_8666,N_8391,N_8434);
nand U8667 (N_8667,N_8111,N_8359);
nor U8668 (N_8668,N_8291,N_8430);
nor U8669 (N_8669,N_8433,N_8052);
nand U8670 (N_8670,N_8141,N_8424);
nor U8671 (N_8671,N_8162,N_8289);
nor U8672 (N_8672,N_8367,N_8257);
and U8673 (N_8673,N_8072,N_8473);
xor U8674 (N_8674,N_8357,N_8423);
and U8675 (N_8675,N_8307,N_8351);
nor U8676 (N_8676,N_8246,N_8334);
and U8677 (N_8677,N_8173,N_8249);
or U8678 (N_8678,N_8089,N_8376);
nand U8679 (N_8679,N_8041,N_8259);
or U8680 (N_8680,N_8362,N_8447);
nor U8681 (N_8681,N_8118,N_8151);
nand U8682 (N_8682,N_8422,N_8085);
nand U8683 (N_8683,N_8360,N_8297);
xor U8684 (N_8684,N_8008,N_8300);
nand U8685 (N_8685,N_8005,N_8080);
nand U8686 (N_8686,N_8271,N_8331);
nand U8687 (N_8687,N_8472,N_8480);
and U8688 (N_8688,N_8318,N_8179);
nand U8689 (N_8689,N_8102,N_8124);
xnor U8690 (N_8690,N_8032,N_8157);
nor U8691 (N_8691,N_8342,N_8358);
and U8692 (N_8692,N_8025,N_8195);
and U8693 (N_8693,N_8312,N_8183);
nor U8694 (N_8694,N_8293,N_8372);
nor U8695 (N_8695,N_8091,N_8283);
nor U8696 (N_8696,N_8013,N_8081);
or U8697 (N_8697,N_8414,N_8267);
nand U8698 (N_8698,N_8175,N_8170);
and U8699 (N_8699,N_8314,N_8361);
nor U8700 (N_8700,N_8387,N_8095);
and U8701 (N_8701,N_8399,N_8350);
or U8702 (N_8702,N_8236,N_8346);
and U8703 (N_8703,N_8244,N_8042);
or U8704 (N_8704,N_8476,N_8035);
or U8705 (N_8705,N_8122,N_8452);
and U8706 (N_8706,N_8001,N_8030);
nor U8707 (N_8707,N_8479,N_8031);
and U8708 (N_8708,N_8493,N_8320);
and U8709 (N_8709,N_8092,N_8202);
nor U8710 (N_8710,N_8079,N_8418);
nand U8711 (N_8711,N_8321,N_8400);
nand U8712 (N_8712,N_8096,N_8366);
nand U8713 (N_8713,N_8420,N_8003);
nand U8714 (N_8714,N_8213,N_8090);
nor U8715 (N_8715,N_8478,N_8352);
nand U8716 (N_8716,N_8224,N_8443);
or U8717 (N_8717,N_8449,N_8436);
and U8718 (N_8718,N_8459,N_8115);
xor U8719 (N_8719,N_8049,N_8226);
nor U8720 (N_8720,N_8498,N_8395);
nor U8721 (N_8721,N_8148,N_8007);
xnor U8722 (N_8722,N_8039,N_8356);
nor U8723 (N_8723,N_8335,N_8164);
nor U8724 (N_8724,N_8263,N_8232);
nand U8725 (N_8725,N_8121,N_8329);
nand U8726 (N_8726,N_8237,N_8258);
nand U8727 (N_8727,N_8429,N_8497);
or U8728 (N_8728,N_8301,N_8426);
nand U8729 (N_8729,N_8057,N_8022);
xnor U8730 (N_8730,N_8290,N_8033);
nand U8731 (N_8731,N_8225,N_8171);
or U8732 (N_8732,N_8028,N_8114);
nand U8733 (N_8733,N_8136,N_8239);
or U8734 (N_8734,N_8485,N_8339);
and U8735 (N_8735,N_8116,N_8101);
or U8736 (N_8736,N_8427,N_8353);
nor U8737 (N_8737,N_8243,N_8216);
and U8738 (N_8738,N_8154,N_8254);
nor U8739 (N_8739,N_8066,N_8421);
nor U8740 (N_8740,N_8322,N_8256);
xor U8741 (N_8741,N_8166,N_8217);
nor U8742 (N_8742,N_8292,N_8453);
or U8743 (N_8743,N_8024,N_8218);
and U8744 (N_8744,N_8055,N_8103);
nand U8745 (N_8745,N_8398,N_8466);
nor U8746 (N_8746,N_8457,N_8412);
nand U8747 (N_8747,N_8229,N_8355);
xnor U8748 (N_8748,N_8276,N_8184);
xor U8749 (N_8749,N_8105,N_8324);
or U8750 (N_8750,N_8083,N_8282);
xnor U8751 (N_8751,N_8160,N_8425);
or U8752 (N_8752,N_8010,N_8294);
and U8753 (N_8753,N_8311,N_8054);
or U8754 (N_8754,N_8031,N_8275);
and U8755 (N_8755,N_8072,N_8314);
and U8756 (N_8756,N_8030,N_8092);
or U8757 (N_8757,N_8479,N_8123);
nand U8758 (N_8758,N_8384,N_8152);
nand U8759 (N_8759,N_8252,N_8425);
or U8760 (N_8760,N_8367,N_8015);
nor U8761 (N_8761,N_8403,N_8184);
nand U8762 (N_8762,N_8232,N_8277);
nand U8763 (N_8763,N_8001,N_8129);
and U8764 (N_8764,N_8026,N_8439);
nor U8765 (N_8765,N_8254,N_8102);
xnor U8766 (N_8766,N_8219,N_8353);
and U8767 (N_8767,N_8334,N_8300);
or U8768 (N_8768,N_8171,N_8243);
nor U8769 (N_8769,N_8411,N_8456);
nand U8770 (N_8770,N_8218,N_8489);
nor U8771 (N_8771,N_8002,N_8304);
nand U8772 (N_8772,N_8317,N_8307);
nor U8773 (N_8773,N_8493,N_8072);
nor U8774 (N_8774,N_8002,N_8097);
and U8775 (N_8775,N_8229,N_8274);
and U8776 (N_8776,N_8120,N_8279);
nand U8777 (N_8777,N_8154,N_8102);
nor U8778 (N_8778,N_8370,N_8029);
and U8779 (N_8779,N_8456,N_8111);
and U8780 (N_8780,N_8066,N_8300);
xnor U8781 (N_8781,N_8465,N_8046);
nand U8782 (N_8782,N_8003,N_8318);
nor U8783 (N_8783,N_8030,N_8074);
or U8784 (N_8784,N_8286,N_8141);
xnor U8785 (N_8785,N_8297,N_8337);
or U8786 (N_8786,N_8129,N_8220);
nor U8787 (N_8787,N_8010,N_8296);
or U8788 (N_8788,N_8148,N_8260);
nor U8789 (N_8789,N_8226,N_8105);
or U8790 (N_8790,N_8117,N_8202);
nor U8791 (N_8791,N_8373,N_8400);
xor U8792 (N_8792,N_8179,N_8010);
or U8793 (N_8793,N_8086,N_8471);
xnor U8794 (N_8794,N_8172,N_8192);
and U8795 (N_8795,N_8167,N_8444);
nor U8796 (N_8796,N_8386,N_8093);
nand U8797 (N_8797,N_8049,N_8092);
nand U8798 (N_8798,N_8455,N_8255);
and U8799 (N_8799,N_8381,N_8234);
nor U8800 (N_8800,N_8080,N_8011);
or U8801 (N_8801,N_8125,N_8123);
or U8802 (N_8802,N_8149,N_8152);
nor U8803 (N_8803,N_8266,N_8147);
nor U8804 (N_8804,N_8248,N_8018);
nor U8805 (N_8805,N_8172,N_8135);
nor U8806 (N_8806,N_8285,N_8090);
or U8807 (N_8807,N_8056,N_8135);
nand U8808 (N_8808,N_8352,N_8476);
and U8809 (N_8809,N_8385,N_8074);
and U8810 (N_8810,N_8420,N_8465);
nand U8811 (N_8811,N_8226,N_8460);
or U8812 (N_8812,N_8313,N_8015);
nor U8813 (N_8813,N_8395,N_8468);
nor U8814 (N_8814,N_8060,N_8099);
nor U8815 (N_8815,N_8290,N_8006);
or U8816 (N_8816,N_8476,N_8065);
nand U8817 (N_8817,N_8262,N_8376);
or U8818 (N_8818,N_8018,N_8403);
nor U8819 (N_8819,N_8442,N_8279);
and U8820 (N_8820,N_8257,N_8089);
nand U8821 (N_8821,N_8427,N_8081);
xor U8822 (N_8822,N_8138,N_8304);
nand U8823 (N_8823,N_8007,N_8149);
nor U8824 (N_8824,N_8252,N_8080);
nand U8825 (N_8825,N_8360,N_8026);
and U8826 (N_8826,N_8099,N_8338);
xnor U8827 (N_8827,N_8089,N_8155);
xnor U8828 (N_8828,N_8087,N_8217);
or U8829 (N_8829,N_8302,N_8189);
nor U8830 (N_8830,N_8324,N_8497);
nand U8831 (N_8831,N_8107,N_8149);
nor U8832 (N_8832,N_8443,N_8347);
nor U8833 (N_8833,N_8217,N_8422);
xor U8834 (N_8834,N_8176,N_8342);
nor U8835 (N_8835,N_8411,N_8310);
nor U8836 (N_8836,N_8189,N_8239);
and U8837 (N_8837,N_8019,N_8476);
and U8838 (N_8838,N_8006,N_8250);
or U8839 (N_8839,N_8308,N_8467);
and U8840 (N_8840,N_8178,N_8312);
nand U8841 (N_8841,N_8334,N_8101);
nor U8842 (N_8842,N_8322,N_8048);
and U8843 (N_8843,N_8107,N_8476);
or U8844 (N_8844,N_8365,N_8298);
or U8845 (N_8845,N_8345,N_8295);
nor U8846 (N_8846,N_8380,N_8169);
nand U8847 (N_8847,N_8050,N_8274);
or U8848 (N_8848,N_8257,N_8328);
and U8849 (N_8849,N_8288,N_8219);
and U8850 (N_8850,N_8112,N_8177);
and U8851 (N_8851,N_8451,N_8176);
nand U8852 (N_8852,N_8212,N_8411);
nor U8853 (N_8853,N_8234,N_8157);
and U8854 (N_8854,N_8042,N_8216);
or U8855 (N_8855,N_8179,N_8487);
nand U8856 (N_8856,N_8186,N_8331);
nor U8857 (N_8857,N_8250,N_8284);
or U8858 (N_8858,N_8339,N_8383);
xor U8859 (N_8859,N_8352,N_8190);
nor U8860 (N_8860,N_8069,N_8271);
nand U8861 (N_8861,N_8206,N_8335);
nand U8862 (N_8862,N_8084,N_8319);
or U8863 (N_8863,N_8136,N_8468);
nand U8864 (N_8864,N_8214,N_8478);
nor U8865 (N_8865,N_8145,N_8183);
and U8866 (N_8866,N_8160,N_8449);
or U8867 (N_8867,N_8408,N_8175);
or U8868 (N_8868,N_8418,N_8177);
nand U8869 (N_8869,N_8114,N_8182);
nand U8870 (N_8870,N_8061,N_8028);
or U8871 (N_8871,N_8108,N_8118);
nor U8872 (N_8872,N_8291,N_8118);
nand U8873 (N_8873,N_8226,N_8016);
and U8874 (N_8874,N_8490,N_8056);
xnor U8875 (N_8875,N_8036,N_8078);
xor U8876 (N_8876,N_8311,N_8322);
nor U8877 (N_8877,N_8073,N_8494);
or U8878 (N_8878,N_8301,N_8384);
or U8879 (N_8879,N_8305,N_8123);
or U8880 (N_8880,N_8294,N_8496);
xnor U8881 (N_8881,N_8468,N_8356);
and U8882 (N_8882,N_8046,N_8374);
nor U8883 (N_8883,N_8328,N_8096);
or U8884 (N_8884,N_8237,N_8172);
or U8885 (N_8885,N_8202,N_8348);
or U8886 (N_8886,N_8206,N_8285);
or U8887 (N_8887,N_8348,N_8165);
and U8888 (N_8888,N_8143,N_8339);
or U8889 (N_8889,N_8192,N_8483);
or U8890 (N_8890,N_8140,N_8184);
nor U8891 (N_8891,N_8365,N_8007);
nand U8892 (N_8892,N_8243,N_8403);
nand U8893 (N_8893,N_8235,N_8180);
xor U8894 (N_8894,N_8379,N_8075);
nand U8895 (N_8895,N_8310,N_8272);
nor U8896 (N_8896,N_8152,N_8354);
nor U8897 (N_8897,N_8026,N_8259);
and U8898 (N_8898,N_8452,N_8128);
nor U8899 (N_8899,N_8454,N_8278);
nand U8900 (N_8900,N_8275,N_8458);
or U8901 (N_8901,N_8484,N_8228);
and U8902 (N_8902,N_8208,N_8221);
nor U8903 (N_8903,N_8428,N_8138);
and U8904 (N_8904,N_8082,N_8432);
xor U8905 (N_8905,N_8172,N_8077);
xnor U8906 (N_8906,N_8140,N_8089);
and U8907 (N_8907,N_8144,N_8183);
nand U8908 (N_8908,N_8397,N_8323);
xnor U8909 (N_8909,N_8152,N_8130);
or U8910 (N_8910,N_8483,N_8298);
xor U8911 (N_8911,N_8299,N_8466);
nand U8912 (N_8912,N_8257,N_8434);
and U8913 (N_8913,N_8293,N_8056);
nand U8914 (N_8914,N_8424,N_8211);
nand U8915 (N_8915,N_8381,N_8110);
or U8916 (N_8916,N_8279,N_8119);
nand U8917 (N_8917,N_8058,N_8205);
or U8918 (N_8918,N_8265,N_8187);
nand U8919 (N_8919,N_8300,N_8275);
and U8920 (N_8920,N_8070,N_8371);
or U8921 (N_8921,N_8213,N_8164);
and U8922 (N_8922,N_8033,N_8114);
nand U8923 (N_8923,N_8269,N_8139);
nor U8924 (N_8924,N_8081,N_8443);
nand U8925 (N_8925,N_8320,N_8002);
nand U8926 (N_8926,N_8489,N_8364);
xnor U8927 (N_8927,N_8454,N_8489);
or U8928 (N_8928,N_8320,N_8267);
nand U8929 (N_8929,N_8056,N_8318);
or U8930 (N_8930,N_8483,N_8020);
nor U8931 (N_8931,N_8216,N_8334);
and U8932 (N_8932,N_8203,N_8476);
nand U8933 (N_8933,N_8437,N_8334);
nand U8934 (N_8934,N_8401,N_8490);
and U8935 (N_8935,N_8050,N_8345);
nand U8936 (N_8936,N_8375,N_8125);
or U8937 (N_8937,N_8008,N_8225);
or U8938 (N_8938,N_8275,N_8215);
nor U8939 (N_8939,N_8079,N_8018);
and U8940 (N_8940,N_8226,N_8024);
nand U8941 (N_8941,N_8130,N_8104);
or U8942 (N_8942,N_8341,N_8498);
and U8943 (N_8943,N_8045,N_8362);
or U8944 (N_8944,N_8035,N_8301);
nor U8945 (N_8945,N_8087,N_8027);
and U8946 (N_8946,N_8055,N_8020);
and U8947 (N_8947,N_8112,N_8185);
nand U8948 (N_8948,N_8326,N_8156);
nand U8949 (N_8949,N_8110,N_8211);
xnor U8950 (N_8950,N_8062,N_8299);
and U8951 (N_8951,N_8061,N_8109);
nand U8952 (N_8952,N_8391,N_8157);
nand U8953 (N_8953,N_8006,N_8048);
xor U8954 (N_8954,N_8296,N_8375);
xnor U8955 (N_8955,N_8035,N_8485);
nor U8956 (N_8956,N_8305,N_8054);
and U8957 (N_8957,N_8454,N_8398);
nor U8958 (N_8958,N_8336,N_8484);
xor U8959 (N_8959,N_8004,N_8222);
nor U8960 (N_8960,N_8085,N_8036);
or U8961 (N_8961,N_8060,N_8286);
or U8962 (N_8962,N_8192,N_8042);
nand U8963 (N_8963,N_8069,N_8128);
or U8964 (N_8964,N_8491,N_8176);
nor U8965 (N_8965,N_8299,N_8396);
nand U8966 (N_8966,N_8166,N_8203);
or U8967 (N_8967,N_8042,N_8412);
or U8968 (N_8968,N_8211,N_8170);
nand U8969 (N_8969,N_8155,N_8208);
nor U8970 (N_8970,N_8142,N_8416);
or U8971 (N_8971,N_8385,N_8442);
or U8972 (N_8972,N_8165,N_8449);
nor U8973 (N_8973,N_8024,N_8488);
nand U8974 (N_8974,N_8235,N_8116);
and U8975 (N_8975,N_8356,N_8011);
nor U8976 (N_8976,N_8154,N_8240);
nor U8977 (N_8977,N_8249,N_8457);
nor U8978 (N_8978,N_8478,N_8294);
nor U8979 (N_8979,N_8346,N_8269);
nand U8980 (N_8980,N_8182,N_8424);
and U8981 (N_8981,N_8141,N_8323);
or U8982 (N_8982,N_8214,N_8144);
or U8983 (N_8983,N_8113,N_8214);
nor U8984 (N_8984,N_8245,N_8250);
xnor U8985 (N_8985,N_8180,N_8092);
and U8986 (N_8986,N_8433,N_8119);
and U8987 (N_8987,N_8001,N_8076);
and U8988 (N_8988,N_8386,N_8329);
or U8989 (N_8989,N_8102,N_8056);
or U8990 (N_8990,N_8488,N_8012);
nor U8991 (N_8991,N_8081,N_8279);
and U8992 (N_8992,N_8340,N_8019);
or U8993 (N_8993,N_8059,N_8305);
nor U8994 (N_8994,N_8332,N_8333);
or U8995 (N_8995,N_8188,N_8331);
and U8996 (N_8996,N_8298,N_8162);
nand U8997 (N_8997,N_8150,N_8349);
and U8998 (N_8998,N_8173,N_8343);
and U8999 (N_8999,N_8014,N_8072);
and U9000 (N_9000,N_8645,N_8656);
nor U9001 (N_9001,N_8722,N_8578);
or U9002 (N_9002,N_8883,N_8876);
or U9003 (N_9003,N_8516,N_8840);
or U9004 (N_9004,N_8556,N_8568);
nand U9005 (N_9005,N_8592,N_8905);
and U9006 (N_9006,N_8533,N_8659);
nor U9007 (N_9007,N_8671,N_8717);
nor U9008 (N_9008,N_8588,N_8963);
and U9009 (N_9009,N_8683,N_8901);
or U9010 (N_9010,N_8941,N_8824);
nor U9011 (N_9011,N_8687,N_8816);
and U9012 (N_9012,N_8637,N_8991);
or U9013 (N_9013,N_8718,N_8648);
nand U9014 (N_9014,N_8909,N_8910);
or U9015 (N_9015,N_8721,N_8693);
nand U9016 (N_9016,N_8647,N_8965);
and U9017 (N_9017,N_8778,N_8799);
xnor U9018 (N_9018,N_8789,N_8943);
xor U9019 (N_9019,N_8567,N_8747);
and U9020 (N_9020,N_8775,N_8733);
or U9021 (N_9021,N_8615,N_8700);
nand U9022 (N_9022,N_8967,N_8825);
or U9023 (N_9023,N_8852,N_8916);
nand U9024 (N_9024,N_8537,N_8593);
nor U9025 (N_9025,N_8996,N_8969);
xnor U9026 (N_9026,N_8971,N_8552);
xor U9027 (N_9027,N_8680,N_8940);
nand U9028 (N_9028,N_8815,N_8538);
nand U9029 (N_9029,N_8528,N_8893);
or U9030 (N_9030,N_8932,N_8841);
or U9031 (N_9031,N_8754,N_8844);
or U9032 (N_9032,N_8569,N_8622);
and U9033 (N_9033,N_8701,N_8741);
and U9034 (N_9034,N_8633,N_8895);
nor U9035 (N_9035,N_8939,N_8655);
nor U9036 (N_9036,N_8676,N_8699);
nor U9037 (N_9037,N_8880,N_8510);
nor U9038 (N_9038,N_8731,N_8817);
and U9039 (N_9039,N_8867,N_8842);
nor U9040 (N_9040,N_8650,N_8564);
or U9041 (N_9041,N_8604,N_8511);
and U9042 (N_9042,N_8755,N_8752);
nor U9043 (N_9043,N_8508,N_8649);
nor U9044 (N_9044,N_8989,N_8773);
and U9045 (N_9045,N_8850,N_8677);
nor U9046 (N_9046,N_8805,N_8808);
nand U9047 (N_9047,N_8559,N_8502);
and U9048 (N_9048,N_8781,N_8782);
nor U9049 (N_9049,N_8685,N_8864);
nor U9050 (N_9050,N_8549,N_8684);
nor U9051 (N_9051,N_8667,N_8625);
and U9052 (N_9052,N_8575,N_8545);
nor U9053 (N_9053,N_8660,N_8813);
nor U9054 (N_9054,N_8597,N_8602);
or U9055 (N_9055,N_8924,N_8703);
nand U9056 (N_9056,N_8705,N_8964);
xnor U9057 (N_9057,N_8746,N_8935);
and U9058 (N_9058,N_8740,N_8823);
or U9059 (N_9059,N_8620,N_8665);
or U9060 (N_9060,N_8957,N_8580);
nor U9061 (N_9061,N_8523,N_8838);
or U9062 (N_9062,N_8889,N_8504);
and U9063 (N_9063,N_8662,N_8669);
xnor U9064 (N_9064,N_8535,N_8945);
and U9065 (N_9065,N_8692,N_8832);
nor U9066 (N_9066,N_8636,N_8628);
nor U9067 (N_9067,N_8809,N_8713);
nand U9068 (N_9068,N_8818,N_8942);
nor U9069 (N_9069,N_8554,N_8888);
nor U9070 (N_9070,N_8952,N_8987);
nand U9071 (N_9071,N_8710,N_8860);
and U9072 (N_9072,N_8953,N_8617);
nor U9073 (N_9073,N_8834,N_8576);
and U9074 (N_9074,N_8854,N_8981);
xor U9075 (N_9075,N_8959,N_8506);
or U9076 (N_9076,N_8931,N_8724);
nand U9077 (N_9077,N_8513,N_8806);
or U9078 (N_9078,N_8811,N_8727);
nor U9079 (N_9079,N_8837,N_8798);
nand U9080 (N_9080,N_8946,N_8877);
and U9081 (N_9081,N_8890,N_8595);
or U9082 (N_9082,N_8779,N_8652);
nor U9083 (N_9083,N_8723,N_8956);
nor U9084 (N_9084,N_8530,N_8846);
nand U9085 (N_9085,N_8546,N_8878);
and U9086 (N_9086,N_8682,N_8827);
or U9087 (N_9087,N_8581,N_8830);
nand U9088 (N_9088,N_8715,N_8766);
and U9089 (N_9089,N_8978,N_8947);
or U9090 (N_9090,N_8785,N_8608);
or U9091 (N_9091,N_8630,N_8758);
or U9092 (N_9092,N_8536,N_8734);
and U9093 (N_9093,N_8992,N_8771);
nor U9094 (N_9094,N_8547,N_8560);
nor U9095 (N_9095,N_8904,N_8810);
nor U9096 (N_9096,N_8875,N_8606);
or U9097 (N_9097,N_8930,N_8761);
nand U9098 (N_9098,N_8619,N_8562);
nand U9099 (N_9099,N_8640,N_8541);
and U9100 (N_9100,N_8632,N_8828);
and U9101 (N_9101,N_8661,N_8979);
nand U9102 (N_9102,N_8975,N_8928);
and U9103 (N_9103,N_8995,N_8960);
nand U9104 (N_9104,N_8836,N_8600);
nand U9105 (N_9105,N_8749,N_8599);
and U9106 (N_9106,N_8814,N_8988);
or U9107 (N_9107,N_8977,N_8641);
or U9108 (N_9108,N_8925,N_8524);
xnor U9109 (N_9109,N_8797,N_8833);
nand U9110 (N_9110,N_8743,N_8871);
and U9111 (N_9111,N_8673,N_8745);
nor U9112 (N_9112,N_8984,N_8514);
or U9113 (N_9113,N_8885,N_8865);
and U9114 (N_9114,N_8638,N_8635);
nor U9115 (N_9115,N_8561,N_8732);
nor U9116 (N_9116,N_8920,N_8627);
and U9117 (N_9117,N_8738,N_8621);
nor U9118 (N_9118,N_8804,N_8565);
nor U9119 (N_9119,N_8949,N_8594);
and U9120 (N_9120,N_8589,N_8708);
nor U9121 (N_9121,N_8879,N_8726);
and U9122 (N_9122,N_8634,N_8794);
nor U9123 (N_9123,N_8861,N_8847);
and U9124 (N_9124,N_8590,N_8826);
xnor U9125 (N_9125,N_8739,N_8614);
or U9126 (N_9126,N_8881,N_8674);
or U9127 (N_9127,N_8767,N_8571);
or U9128 (N_9128,N_8643,N_8917);
nand U9129 (N_9129,N_8657,N_8985);
nand U9130 (N_9130,N_8672,N_8906);
or U9131 (N_9131,N_8972,N_8911);
xnor U9132 (N_9132,N_8938,N_8736);
or U9133 (N_9133,N_8500,N_8531);
and U9134 (N_9134,N_8585,N_8927);
and U9135 (N_9135,N_8800,N_8651);
and U9136 (N_9136,N_8777,N_8756);
or U9137 (N_9137,N_8955,N_8821);
nand U9138 (N_9138,N_8873,N_8714);
or U9139 (N_9139,N_8866,N_8712);
or U9140 (N_9140,N_8919,N_8768);
nand U9141 (N_9141,N_8729,N_8848);
nor U9142 (N_9142,N_8521,N_8646);
and U9143 (N_9143,N_8558,N_8937);
or U9144 (N_9144,N_8970,N_8596);
or U9145 (N_9145,N_8764,N_8954);
xor U9146 (N_9146,N_8760,N_8509);
nor U9147 (N_9147,N_8696,N_8923);
nand U9148 (N_9148,N_8572,N_8934);
nor U9149 (N_9149,N_8644,N_8796);
nand U9150 (N_9150,N_8570,N_8757);
or U9151 (N_9151,N_8610,N_8983);
or U9152 (N_9152,N_8618,N_8835);
or U9153 (N_9153,N_8612,N_8605);
nand U9154 (N_9154,N_8582,N_8759);
nor U9155 (N_9155,N_8962,N_8642);
xnor U9156 (N_9156,N_8573,N_8550);
nand U9157 (N_9157,N_8668,N_8613);
nor U9158 (N_9158,N_8742,N_8994);
nand U9159 (N_9159,N_8503,N_8772);
or U9160 (N_9160,N_8831,N_8664);
or U9161 (N_9161,N_8525,N_8858);
nand U9162 (N_9162,N_8540,N_8851);
nor U9163 (N_9163,N_8587,N_8654);
nor U9164 (N_9164,N_8702,N_8999);
nand U9165 (N_9165,N_8584,N_8863);
nand U9166 (N_9166,N_8929,N_8522);
nor U9167 (N_9167,N_8856,N_8998);
nor U9168 (N_9168,N_8539,N_8859);
nor U9169 (N_9169,N_8770,N_8719);
or U9170 (N_9170,N_8790,N_8902);
nor U9171 (N_9171,N_8529,N_8926);
nor U9172 (N_9172,N_8542,N_8780);
nand U9173 (N_9173,N_8598,N_8744);
nor U9174 (N_9174,N_8944,N_8855);
or U9175 (N_9175,N_8519,N_8591);
or U9176 (N_9176,N_8872,N_8505);
nor U9177 (N_9177,N_8544,N_8534);
nand U9178 (N_9178,N_8795,N_8517);
or U9179 (N_9179,N_8765,N_8912);
nor U9180 (N_9180,N_8896,N_8958);
nor U9181 (N_9181,N_8857,N_8900);
nor U9182 (N_9182,N_8557,N_8913);
xnor U9183 (N_9183,N_8518,N_8526);
nor U9184 (N_9184,N_8907,N_8936);
and U9185 (N_9185,N_8976,N_8974);
or U9186 (N_9186,N_8611,N_8698);
or U9187 (N_9187,N_8653,N_8512);
nand U9188 (N_9188,N_8769,N_8691);
nand U9189 (N_9189,N_8884,N_8898);
nand U9190 (N_9190,N_8762,N_8753);
and U9191 (N_9191,N_8786,N_8709);
and U9192 (N_9192,N_8829,N_8787);
xnor U9193 (N_9193,N_8675,N_8555);
or U9194 (N_9194,N_8922,N_8689);
or U9195 (N_9195,N_8601,N_8603);
nor U9196 (N_9196,N_8706,N_8574);
nand U9197 (N_9197,N_8725,N_8807);
nor U9198 (N_9198,N_8870,N_8982);
or U9199 (N_9199,N_8891,N_8933);
nor U9200 (N_9200,N_8914,N_8792);
nand U9201 (N_9201,N_8822,N_8763);
and U9202 (N_9202,N_8686,N_8894);
xor U9203 (N_9203,N_8980,N_8666);
nor U9204 (N_9204,N_8532,N_8820);
or U9205 (N_9205,N_8882,N_8629);
and U9206 (N_9206,N_8681,N_8948);
xor U9207 (N_9207,N_8750,N_8819);
and U9208 (N_9208,N_8951,N_8791);
nand U9209 (N_9209,N_8678,N_8961);
and U9210 (N_9210,N_8774,N_8973);
nand U9211 (N_9211,N_8950,N_8801);
xnor U9212 (N_9212,N_8688,N_8968);
nor U9213 (N_9213,N_8577,N_8694);
nand U9214 (N_9214,N_8515,N_8553);
and U9215 (N_9215,N_8784,N_8583);
and U9216 (N_9216,N_8869,N_8623);
or U9217 (N_9217,N_8507,N_8783);
xnor U9218 (N_9218,N_8501,N_8616);
and U9219 (N_9219,N_8711,N_8839);
and U9220 (N_9220,N_8639,N_8735);
nand U9221 (N_9221,N_8566,N_8663);
nor U9222 (N_9222,N_8849,N_8737);
and U9223 (N_9223,N_8899,N_8966);
nand U9224 (N_9224,N_8658,N_8579);
nor U9225 (N_9225,N_8776,N_8728);
nor U9226 (N_9226,N_8986,N_8631);
or U9227 (N_9227,N_8887,N_8697);
and U9228 (N_9228,N_8543,N_8563);
nor U9229 (N_9229,N_8803,N_8812);
or U9230 (N_9230,N_8751,N_8997);
nor U9231 (N_9231,N_8626,N_8716);
or U9232 (N_9232,N_8845,N_8874);
and U9233 (N_9233,N_8788,N_8853);
or U9234 (N_9234,N_8921,N_8862);
and U9235 (N_9235,N_8609,N_8868);
nor U9236 (N_9236,N_8704,N_8793);
or U9237 (N_9237,N_8679,N_8720);
xnor U9238 (N_9238,N_8670,N_8520);
nand U9239 (N_9239,N_8748,N_8695);
nor U9240 (N_9240,N_8908,N_8586);
or U9241 (N_9241,N_8624,N_8843);
nor U9242 (N_9242,N_8548,N_8690);
nand U9243 (N_9243,N_8607,N_8915);
nand U9244 (N_9244,N_8990,N_8527);
nor U9245 (N_9245,N_8892,N_8897);
or U9246 (N_9246,N_8707,N_8730);
nand U9247 (N_9247,N_8802,N_8993);
and U9248 (N_9248,N_8918,N_8903);
and U9249 (N_9249,N_8886,N_8551);
or U9250 (N_9250,N_8694,N_8820);
or U9251 (N_9251,N_8879,N_8605);
xor U9252 (N_9252,N_8740,N_8893);
and U9253 (N_9253,N_8586,N_8556);
xor U9254 (N_9254,N_8609,N_8576);
and U9255 (N_9255,N_8684,N_8776);
nand U9256 (N_9256,N_8683,N_8966);
nand U9257 (N_9257,N_8619,N_8845);
nor U9258 (N_9258,N_8762,N_8607);
nand U9259 (N_9259,N_8929,N_8895);
nand U9260 (N_9260,N_8972,N_8864);
or U9261 (N_9261,N_8774,N_8737);
or U9262 (N_9262,N_8948,N_8779);
nor U9263 (N_9263,N_8811,N_8863);
and U9264 (N_9264,N_8627,N_8944);
xor U9265 (N_9265,N_8525,N_8504);
nand U9266 (N_9266,N_8537,N_8867);
and U9267 (N_9267,N_8853,N_8984);
or U9268 (N_9268,N_8933,N_8596);
or U9269 (N_9269,N_8600,N_8941);
nor U9270 (N_9270,N_8702,N_8863);
nor U9271 (N_9271,N_8966,N_8878);
and U9272 (N_9272,N_8811,N_8874);
and U9273 (N_9273,N_8878,N_8879);
or U9274 (N_9274,N_8529,N_8604);
nand U9275 (N_9275,N_8619,N_8778);
nor U9276 (N_9276,N_8643,N_8972);
and U9277 (N_9277,N_8512,N_8633);
or U9278 (N_9278,N_8640,N_8866);
nor U9279 (N_9279,N_8754,N_8528);
nor U9280 (N_9280,N_8813,N_8925);
nand U9281 (N_9281,N_8542,N_8995);
nor U9282 (N_9282,N_8925,N_8516);
or U9283 (N_9283,N_8867,N_8791);
and U9284 (N_9284,N_8615,N_8787);
and U9285 (N_9285,N_8525,N_8657);
and U9286 (N_9286,N_8549,N_8870);
and U9287 (N_9287,N_8898,N_8542);
or U9288 (N_9288,N_8814,N_8845);
or U9289 (N_9289,N_8808,N_8698);
nor U9290 (N_9290,N_8519,N_8939);
and U9291 (N_9291,N_8818,N_8871);
nor U9292 (N_9292,N_8921,N_8550);
nor U9293 (N_9293,N_8802,N_8989);
xnor U9294 (N_9294,N_8932,N_8877);
or U9295 (N_9295,N_8762,N_8728);
nor U9296 (N_9296,N_8804,N_8877);
nor U9297 (N_9297,N_8993,N_8950);
nand U9298 (N_9298,N_8769,N_8940);
nor U9299 (N_9299,N_8649,N_8951);
nor U9300 (N_9300,N_8952,N_8647);
nand U9301 (N_9301,N_8737,N_8910);
nand U9302 (N_9302,N_8687,N_8987);
and U9303 (N_9303,N_8807,N_8648);
nand U9304 (N_9304,N_8945,N_8909);
nand U9305 (N_9305,N_8750,N_8832);
and U9306 (N_9306,N_8652,N_8616);
and U9307 (N_9307,N_8742,N_8519);
nand U9308 (N_9308,N_8948,N_8533);
or U9309 (N_9309,N_8679,N_8508);
and U9310 (N_9310,N_8908,N_8513);
nor U9311 (N_9311,N_8557,N_8539);
and U9312 (N_9312,N_8942,N_8690);
nor U9313 (N_9313,N_8533,N_8520);
or U9314 (N_9314,N_8686,N_8727);
and U9315 (N_9315,N_8729,N_8789);
xor U9316 (N_9316,N_8530,N_8835);
xnor U9317 (N_9317,N_8860,N_8728);
or U9318 (N_9318,N_8549,N_8625);
and U9319 (N_9319,N_8923,N_8906);
nand U9320 (N_9320,N_8683,N_8707);
nor U9321 (N_9321,N_8520,N_8511);
or U9322 (N_9322,N_8745,N_8620);
and U9323 (N_9323,N_8820,N_8840);
nand U9324 (N_9324,N_8545,N_8778);
nand U9325 (N_9325,N_8676,N_8817);
and U9326 (N_9326,N_8919,N_8597);
nand U9327 (N_9327,N_8830,N_8896);
nand U9328 (N_9328,N_8829,N_8982);
nand U9329 (N_9329,N_8664,N_8632);
and U9330 (N_9330,N_8960,N_8893);
nand U9331 (N_9331,N_8838,N_8652);
and U9332 (N_9332,N_8709,N_8968);
nand U9333 (N_9333,N_8814,N_8576);
nor U9334 (N_9334,N_8931,N_8819);
or U9335 (N_9335,N_8972,N_8724);
xnor U9336 (N_9336,N_8561,N_8819);
or U9337 (N_9337,N_8537,N_8948);
and U9338 (N_9338,N_8771,N_8793);
or U9339 (N_9339,N_8787,N_8531);
and U9340 (N_9340,N_8745,N_8549);
nand U9341 (N_9341,N_8727,N_8678);
nor U9342 (N_9342,N_8863,N_8983);
or U9343 (N_9343,N_8862,N_8660);
or U9344 (N_9344,N_8564,N_8631);
nor U9345 (N_9345,N_8714,N_8573);
nand U9346 (N_9346,N_8646,N_8849);
and U9347 (N_9347,N_8753,N_8749);
nor U9348 (N_9348,N_8802,N_8767);
nand U9349 (N_9349,N_8569,N_8992);
nor U9350 (N_9350,N_8503,N_8987);
nand U9351 (N_9351,N_8611,N_8749);
xor U9352 (N_9352,N_8841,N_8868);
nor U9353 (N_9353,N_8770,N_8956);
and U9354 (N_9354,N_8576,N_8581);
nor U9355 (N_9355,N_8971,N_8748);
nor U9356 (N_9356,N_8814,N_8530);
nor U9357 (N_9357,N_8682,N_8998);
xnor U9358 (N_9358,N_8520,N_8566);
nand U9359 (N_9359,N_8917,N_8875);
or U9360 (N_9360,N_8824,N_8634);
or U9361 (N_9361,N_8530,N_8668);
nor U9362 (N_9362,N_8684,N_8720);
nand U9363 (N_9363,N_8750,N_8554);
nor U9364 (N_9364,N_8685,N_8701);
or U9365 (N_9365,N_8600,N_8625);
and U9366 (N_9366,N_8701,N_8681);
nand U9367 (N_9367,N_8851,N_8706);
nor U9368 (N_9368,N_8533,N_8710);
nand U9369 (N_9369,N_8822,N_8814);
and U9370 (N_9370,N_8599,N_8709);
nor U9371 (N_9371,N_8905,N_8873);
nor U9372 (N_9372,N_8630,N_8896);
and U9373 (N_9373,N_8782,N_8844);
xor U9374 (N_9374,N_8993,N_8862);
or U9375 (N_9375,N_8683,N_8660);
nand U9376 (N_9376,N_8530,N_8893);
nand U9377 (N_9377,N_8831,N_8653);
and U9378 (N_9378,N_8833,N_8675);
or U9379 (N_9379,N_8501,N_8839);
and U9380 (N_9380,N_8594,N_8922);
and U9381 (N_9381,N_8745,N_8606);
nand U9382 (N_9382,N_8882,N_8704);
nor U9383 (N_9383,N_8532,N_8613);
nand U9384 (N_9384,N_8744,N_8590);
nor U9385 (N_9385,N_8769,N_8704);
and U9386 (N_9386,N_8562,N_8862);
and U9387 (N_9387,N_8545,N_8714);
nand U9388 (N_9388,N_8724,N_8844);
or U9389 (N_9389,N_8949,N_8976);
and U9390 (N_9390,N_8777,N_8819);
or U9391 (N_9391,N_8961,N_8666);
and U9392 (N_9392,N_8613,N_8941);
nor U9393 (N_9393,N_8741,N_8682);
nand U9394 (N_9394,N_8512,N_8637);
and U9395 (N_9395,N_8576,N_8802);
nand U9396 (N_9396,N_8575,N_8714);
or U9397 (N_9397,N_8768,N_8884);
xnor U9398 (N_9398,N_8500,N_8850);
or U9399 (N_9399,N_8531,N_8713);
or U9400 (N_9400,N_8922,N_8905);
nand U9401 (N_9401,N_8511,N_8579);
nand U9402 (N_9402,N_8695,N_8581);
or U9403 (N_9403,N_8920,N_8561);
or U9404 (N_9404,N_8876,N_8722);
nor U9405 (N_9405,N_8681,N_8597);
and U9406 (N_9406,N_8599,N_8884);
nand U9407 (N_9407,N_8682,N_8877);
nor U9408 (N_9408,N_8710,N_8524);
and U9409 (N_9409,N_8676,N_8831);
nand U9410 (N_9410,N_8944,N_8701);
or U9411 (N_9411,N_8748,N_8537);
nand U9412 (N_9412,N_8893,N_8544);
or U9413 (N_9413,N_8599,N_8579);
nand U9414 (N_9414,N_8548,N_8705);
or U9415 (N_9415,N_8582,N_8855);
and U9416 (N_9416,N_8866,N_8657);
nor U9417 (N_9417,N_8764,N_8726);
or U9418 (N_9418,N_8991,N_8812);
nor U9419 (N_9419,N_8946,N_8882);
or U9420 (N_9420,N_8930,N_8513);
xor U9421 (N_9421,N_8604,N_8976);
nand U9422 (N_9422,N_8914,N_8542);
nor U9423 (N_9423,N_8854,N_8939);
nand U9424 (N_9424,N_8595,N_8735);
and U9425 (N_9425,N_8523,N_8731);
nor U9426 (N_9426,N_8649,N_8612);
and U9427 (N_9427,N_8856,N_8821);
nand U9428 (N_9428,N_8718,N_8891);
nand U9429 (N_9429,N_8881,N_8820);
or U9430 (N_9430,N_8938,N_8535);
and U9431 (N_9431,N_8968,N_8983);
or U9432 (N_9432,N_8920,N_8771);
or U9433 (N_9433,N_8851,N_8944);
and U9434 (N_9434,N_8864,N_8836);
xnor U9435 (N_9435,N_8586,N_8642);
nor U9436 (N_9436,N_8853,N_8527);
xnor U9437 (N_9437,N_8992,N_8792);
nand U9438 (N_9438,N_8730,N_8917);
nor U9439 (N_9439,N_8608,N_8936);
or U9440 (N_9440,N_8522,N_8830);
nand U9441 (N_9441,N_8681,N_8572);
or U9442 (N_9442,N_8726,N_8520);
nor U9443 (N_9443,N_8723,N_8862);
and U9444 (N_9444,N_8742,N_8866);
and U9445 (N_9445,N_8768,N_8944);
xor U9446 (N_9446,N_8991,N_8646);
or U9447 (N_9447,N_8547,N_8704);
or U9448 (N_9448,N_8685,N_8524);
and U9449 (N_9449,N_8536,N_8859);
and U9450 (N_9450,N_8978,N_8850);
xnor U9451 (N_9451,N_8513,N_8911);
nor U9452 (N_9452,N_8501,N_8610);
or U9453 (N_9453,N_8893,N_8963);
or U9454 (N_9454,N_8609,N_8951);
or U9455 (N_9455,N_8904,N_8851);
or U9456 (N_9456,N_8988,N_8520);
nor U9457 (N_9457,N_8706,N_8923);
nand U9458 (N_9458,N_8911,N_8597);
xor U9459 (N_9459,N_8717,N_8850);
nand U9460 (N_9460,N_8601,N_8919);
or U9461 (N_9461,N_8999,N_8640);
nand U9462 (N_9462,N_8834,N_8747);
nand U9463 (N_9463,N_8595,N_8871);
and U9464 (N_9464,N_8570,N_8751);
nor U9465 (N_9465,N_8826,N_8711);
or U9466 (N_9466,N_8512,N_8715);
or U9467 (N_9467,N_8679,N_8772);
or U9468 (N_9468,N_8607,N_8991);
or U9469 (N_9469,N_8846,N_8784);
xor U9470 (N_9470,N_8850,N_8872);
xnor U9471 (N_9471,N_8882,N_8568);
and U9472 (N_9472,N_8620,N_8940);
and U9473 (N_9473,N_8664,N_8593);
xor U9474 (N_9474,N_8583,N_8616);
nand U9475 (N_9475,N_8503,N_8971);
and U9476 (N_9476,N_8992,N_8930);
nand U9477 (N_9477,N_8792,N_8955);
or U9478 (N_9478,N_8606,N_8587);
nor U9479 (N_9479,N_8711,N_8525);
and U9480 (N_9480,N_8948,N_8845);
nor U9481 (N_9481,N_8765,N_8850);
and U9482 (N_9482,N_8557,N_8940);
or U9483 (N_9483,N_8509,N_8533);
nor U9484 (N_9484,N_8782,N_8599);
nand U9485 (N_9485,N_8767,N_8887);
nor U9486 (N_9486,N_8927,N_8638);
nor U9487 (N_9487,N_8763,N_8783);
nand U9488 (N_9488,N_8620,N_8758);
nand U9489 (N_9489,N_8694,N_8927);
nor U9490 (N_9490,N_8918,N_8735);
nand U9491 (N_9491,N_8526,N_8917);
or U9492 (N_9492,N_8520,N_8936);
nor U9493 (N_9493,N_8888,N_8921);
or U9494 (N_9494,N_8746,N_8660);
or U9495 (N_9495,N_8727,N_8897);
xor U9496 (N_9496,N_8759,N_8878);
nor U9497 (N_9497,N_8809,N_8893);
nor U9498 (N_9498,N_8953,N_8534);
nor U9499 (N_9499,N_8562,N_8750);
and U9500 (N_9500,N_9093,N_9228);
nand U9501 (N_9501,N_9253,N_9432);
or U9502 (N_9502,N_9124,N_9383);
nor U9503 (N_9503,N_9359,N_9152);
or U9504 (N_9504,N_9068,N_9151);
nor U9505 (N_9505,N_9435,N_9381);
or U9506 (N_9506,N_9287,N_9025);
and U9507 (N_9507,N_9133,N_9330);
or U9508 (N_9508,N_9310,N_9398);
nand U9509 (N_9509,N_9465,N_9146);
nor U9510 (N_9510,N_9247,N_9453);
nand U9511 (N_9511,N_9106,N_9041);
nand U9512 (N_9512,N_9008,N_9427);
nand U9513 (N_9513,N_9457,N_9299);
nand U9514 (N_9514,N_9372,N_9006);
or U9515 (N_9515,N_9073,N_9061);
nand U9516 (N_9516,N_9480,N_9063);
nand U9517 (N_9517,N_9026,N_9069);
nor U9518 (N_9518,N_9312,N_9187);
nor U9519 (N_9519,N_9293,N_9373);
nor U9520 (N_9520,N_9308,N_9346);
nor U9521 (N_9521,N_9119,N_9362);
nand U9522 (N_9522,N_9281,N_9391);
and U9523 (N_9523,N_9379,N_9186);
nand U9524 (N_9524,N_9343,N_9114);
or U9525 (N_9525,N_9035,N_9046);
and U9526 (N_9526,N_9331,N_9324);
nand U9527 (N_9527,N_9080,N_9156);
nand U9528 (N_9528,N_9323,N_9497);
nand U9529 (N_9529,N_9263,N_9364);
xnor U9530 (N_9530,N_9153,N_9447);
and U9531 (N_9531,N_9023,N_9126);
and U9532 (N_9532,N_9201,N_9221);
nor U9533 (N_9533,N_9135,N_9335);
nor U9534 (N_9534,N_9204,N_9474);
and U9535 (N_9535,N_9207,N_9486);
or U9536 (N_9536,N_9386,N_9129);
or U9537 (N_9537,N_9016,N_9467);
or U9538 (N_9538,N_9066,N_9236);
nand U9539 (N_9539,N_9258,N_9367);
nor U9540 (N_9540,N_9326,N_9077);
and U9541 (N_9541,N_9471,N_9036);
or U9542 (N_9542,N_9134,N_9431);
or U9543 (N_9543,N_9316,N_9222);
xor U9544 (N_9544,N_9402,N_9214);
or U9545 (N_9545,N_9065,N_9138);
nor U9546 (N_9546,N_9302,N_9169);
nor U9547 (N_9547,N_9078,N_9081);
xor U9548 (N_9548,N_9105,N_9412);
nor U9549 (N_9549,N_9039,N_9271);
xor U9550 (N_9550,N_9469,N_9085);
xnor U9551 (N_9551,N_9015,N_9244);
nand U9552 (N_9552,N_9366,N_9354);
or U9553 (N_9553,N_9190,N_9418);
and U9554 (N_9554,N_9032,N_9425);
nand U9555 (N_9555,N_9056,N_9405);
nor U9556 (N_9556,N_9002,N_9357);
or U9557 (N_9557,N_9220,N_9136);
or U9558 (N_9558,N_9231,N_9421);
nand U9559 (N_9559,N_9140,N_9194);
xor U9560 (N_9560,N_9481,N_9347);
nor U9561 (N_9561,N_9090,N_9234);
nor U9562 (N_9562,N_9493,N_9157);
xnor U9563 (N_9563,N_9147,N_9202);
and U9564 (N_9564,N_9091,N_9177);
nor U9565 (N_9565,N_9086,N_9175);
and U9566 (N_9566,N_9337,N_9400);
nor U9567 (N_9567,N_9416,N_9322);
xor U9568 (N_9568,N_9473,N_9475);
and U9569 (N_9569,N_9230,N_9328);
xnor U9570 (N_9570,N_9482,N_9254);
nand U9571 (N_9571,N_9104,N_9332);
or U9572 (N_9572,N_9243,N_9092);
nor U9573 (N_9573,N_9076,N_9161);
nor U9574 (N_9574,N_9446,N_9336);
nand U9575 (N_9575,N_9205,N_9297);
and U9576 (N_9576,N_9249,N_9371);
nand U9577 (N_9577,N_9100,N_9437);
and U9578 (N_9578,N_9246,N_9352);
and U9579 (N_9579,N_9392,N_9494);
nor U9580 (N_9580,N_9298,N_9223);
xor U9581 (N_9581,N_9479,N_9178);
and U9582 (N_9582,N_9001,N_9239);
and U9583 (N_9583,N_9195,N_9004);
or U9584 (N_9584,N_9052,N_9111);
or U9585 (N_9585,N_9484,N_9213);
and U9586 (N_9586,N_9266,N_9314);
nand U9587 (N_9587,N_9459,N_9179);
or U9588 (N_9588,N_9462,N_9252);
and U9589 (N_9589,N_9487,N_9245);
xnor U9590 (N_9590,N_9050,N_9313);
xor U9591 (N_9591,N_9227,N_9142);
nor U9592 (N_9592,N_9014,N_9044);
xor U9593 (N_9593,N_9103,N_9436);
or U9594 (N_9594,N_9338,N_9042);
nor U9595 (N_9595,N_9062,N_9451);
and U9596 (N_9596,N_9200,N_9477);
and U9597 (N_9597,N_9466,N_9098);
xnor U9598 (N_9598,N_9376,N_9034);
nor U9599 (N_9599,N_9321,N_9225);
and U9600 (N_9600,N_9208,N_9305);
or U9601 (N_9601,N_9498,N_9210);
or U9602 (N_9602,N_9340,N_9408);
or U9603 (N_9603,N_9422,N_9311);
or U9604 (N_9604,N_9374,N_9072);
or U9605 (N_9605,N_9361,N_9264);
nand U9606 (N_9606,N_9040,N_9250);
or U9607 (N_9607,N_9184,N_9449);
and U9608 (N_9608,N_9087,N_9168);
nand U9609 (N_9609,N_9309,N_9096);
and U9610 (N_9610,N_9251,N_9382);
or U9611 (N_9611,N_9430,N_9443);
nor U9612 (N_9612,N_9012,N_9053);
and U9613 (N_9613,N_9388,N_9351);
or U9614 (N_9614,N_9496,N_9203);
nand U9615 (N_9615,N_9292,N_9334);
and U9616 (N_9616,N_9164,N_9370);
and U9617 (N_9617,N_9289,N_9199);
and U9618 (N_9618,N_9452,N_9420);
nand U9619 (N_9619,N_9294,N_9438);
or U9620 (N_9620,N_9235,N_9472);
nand U9621 (N_9621,N_9083,N_9433);
and U9622 (N_9622,N_9403,N_9127);
nor U9623 (N_9623,N_9256,N_9478);
xor U9624 (N_9624,N_9257,N_9218);
nand U9625 (N_9625,N_9407,N_9132);
and U9626 (N_9626,N_9058,N_9282);
xor U9627 (N_9627,N_9180,N_9277);
nand U9628 (N_9628,N_9048,N_9043);
nor U9629 (N_9629,N_9176,N_9279);
or U9630 (N_9630,N_9095,N_9434);
nor U9631 (N_9631,N_9000,N_9079);
or U9632 (N_9632,N_9306,N_9455);
nor U9633 (N_9633,N_9120,N_9055);
and U9634 (N_9634,N_9182,N_9355);
nor U9635 (N_9635,N_9415,N_9464);
or U9636 (N_9636,N_9375,N_9206);
xnor U9637 (N_9637,N_9089,N_9303);
or U9638 (N_9638,N_9394,N_9229);
or U9639 (N_9639,N_9270,N_9356);
and U9640 (N_9640,N_9448,N_9107);
nand U9641 (N_9641,N_9024,N_9145);
or U9642 (N_9642,N_9007,N_9108);
nor U9643 (N_9643,N_9275,N_9224);
and U9644 (N_9644,N_9369,N_9099);
nor U9645 (N_9645,N_9342,N_9020);
nor U9646 (N_9646,N_9278,N_9211);
nor U9647 (N_9647,N_9242,N_9174);
or U9648 (N_9648,N_9049,N_9353);
or U9649 (N_9649,N_9037,N_9189);
or U9650 (N_9650,N_9395,N_9488);
or U9651 (N_9651,N_9296,N_9377);
or U9652 (N_9652,N_9128,N_9315);
xnor U9653 (N_9653,N_9350,N_9188);
and U9654 (N_9654,N_9196,N_9470);
xnor U9655 (N_9655,N_9365,N_9067);
xor U9656 (N_9656,N_9209,N_9123);
or U9657 (N_9657,N_9409,N_9348);
nor U9658 (N_9658,N_9232,N_9215);
xnor U9659 (N_9659,N_9265,N_9273);
or U9660 (N_9660,N_9021,N_9378);
nand U9661 (N_9661,N_9274,N_9018);
and U9662 (N_9662,N_9461,N_9406);
and U9663 (N_9663,N_9262,N_9149);
or U9664 (N_9664,N_9110,N_9118);
nand U9665 (N_9665,N_9307,N_9304);
nand U9666 (N_9666,N_9181,N_9360);
and U9667 (N_9667,N_9150,N_9476);
or U9668 (N_9668,N_9460,N_9413);
or U9669 (N_9669,N_9094,N_9414);
and U9670 (N_9670,N_9269,N_9341);
or U9671 (N_9671,N_9499,N_9070);
nor U9672 (N_9672,N_9117,N_9295);
nand U9673 (N_9673,N_9489,N_9385);
and U9674 (N_9674,N_9197,N_9329);
nand U9675 (N_9675,N_9440,N_9162);
and U9676 (N_9676,N_9139,N_9283);
or U9677 (N_9677,N_9259,N_9238);
and U9678 (N_9678,N_9419,N_9029);
nand U9679 (N_9679,N_9130,N_9368);
or U9680 (N_9680,N_9059,N_9495);
nand U9681 (N_9681,N_9165,N_9011);
or U9682 (N_9682,N_9280,N_9288);
nor U9683 (N_9683,N_9017,N_9102);
or U9684 (N_9684,N_9284,N_9064);
and U9685 (N_9685,N_9047,N_9028);
or U9686 (N_9686,N_9339,N_9393);
and U9687 (N_9687,N_9003,N_9390);
nor U9688 (N_9688,N_9113,N_9155);
and U9689 (N_9689,N_9082,N_9141);
nand U9690 (N_9690,N_9071,N_9411);
nand U9691 (N_9691,N_9137,N_9019);
and U9692 (N_9692,N_9075,N_9424);
or U9693 (N_9693,N_9492,N_9333);
or U9694 (N_9694,N_9226,N_9417);
nor U9695 (N_9695,N_9276,N_9033);
nand U9696 (N_9696,N_9384,N_9444);
or U9697 (N_9697,N_9185,N_9468);
and U9698 (N_9698,N_9237,N_9445);
or U9699 (N_9699,N_9084,N_9154);
or U9700 (N_9700,N_9159,N_9115);
nand U9701 (N_9701,N_9125,N_9439);
or U9702 (N_9702,N_9112,N_9320);
xnor U9703 (N_9703,N_9248,N_9301);
xnor U9704 (N_9704,N_9255,N_9490);
or U9705 (N_9705,N_9088,N_9217);
xor U9706 (N_9706,N_9442,N_9463);
xor U9707 (N_9707,N_9170,N_9013);
and U9708 (N_9708,N_9010,N_9387);
nand U9709 (N_9709,N_9358,N_9172);
or U9710 (N_9710,N_9038,N_9300);
and U9711 (N_9711,N_9219,N_9173);
and U9712 (N_9712,N_9423,N_9109);
nor U9713 (N_9713,N_9122,N_9344);
nor U9714 (N_9714,N_9260,N_9097);
nor U9715 (N_9715,N_9290,N_9198);
nor U9716 (N_9716,N_9426,N_9456);
xor U9717 (N_9717,N_9131,N_9429);
and U9718 (N_9718,N_9428,N_9009);
nand U9719 (N_9719,N_9345,N_9054);
and U9720 (N_9720,N_9410,N_9193);
or U9721 (N_9721,N_9171,N_9485);
nand U9722 (N_9722,N_9318,N_9491);
and U9723 (N_9723,N_9327,N_9027);
and U9724 (N_9724,N_9286,N_9317);
nor U9725 (N_9725,N_9045,N_9349);
nand U9726 (N_9726,N_9399,N_9116);
nand U9727 (N_9727,N_9158,N_9192);
and U9728 (N_9728,N_9143,N_9057);
nand U9729 (N_9729,N_9144,N_9397);
nand U9730 (N_9730,N_9212,N_9325);
nor U9731 (N_9731,N_9363,N_9454);
nand U9732 (N_9732,N_9051,N_9261);
xnor U9733 (N_9733,N_9380,N_9074);
and U9734 (N_9734,N_9291,N_9022);
nor U9735 (N_9735,N_9450,N_9101);
nor U9736 (N_9736,N_9404,N_9268);
nor U9737 (N_9737,N_9285,N_9191);
and U9738 (N_9738,N_9160,N_9233);
or U9739 (N_9739,N_9458,N_9166);
or U9740 (N_9740,N_9319,N_9005);
and U9741 (N_9741,N_9401,N_9148);
or U9742 (N_9742,N_9272,N_9216);
and U9743 (N_9743,N_9031,N_9241);
and U9744 (N_9744,N_9267,N_9240);
or U9745 (N_9745,N_9396,N_9389);
or U9746 (N_9746,N_9441,N_9167);
nor U9747 (N_9747,N_9121,N_9060);
nor U9748 (N_9748,N_9483,N_9030);
xnor U9749 (N_9749,N_9163,N_9183);
and U9750 (N_9750,N_9429,N_9093);
and U9751 (N_9751,N_9296,N_9479);
or U9752 (N_9752,N_9206,N_9065);
or U9753 (N_9753,N_9205,N_9180);
nand U9754 (N_9754,N_9315,N_9182);
nand U9755 (N_9755,N_9272,N_9453);
and U9756 (N_9756,N_9266,N_9139);
nor U9757 (N_9757,N_9262,N_9032);
nand U9758 (N_9758,N_9344,N_9001);
or U9759 (N_9759,N_9379,N_9251);
nor U9760 (N_9760,N_9284,N_9322);
or U9761 (N_9761,N_9364,N_9360);
or U9762 (N_9762,N_9197,N_9171);
nand U9763 (N_9763,N_9411,N_9086);
nand U9764 (N_9764,N_9442,N_9257);
and U9765 (N_9765,N_9273,N_9142);
nor U9766 (N_9766,N_9385,N_9257);
or U9767 (N_9767,N_9357,N_9284);
nor U9768 (N_9768,N_9237,N_9368);
or U9769 (N_9769,N_9324,N_9273);
nor U9770 (N_9770,N_9007,N_9406);
or U9771 (N_9771,N_9131,N_9044);
and U9772 (N_9772,N_9014,N_9252);
and U9773 (N_9773,N_9421,N_9240);
xnor U9774 (N_9774,N_9405,N_9188);
nor U9775 (N_9775,N_9359,N_9381);
nor U9776 (N_9776,N_9489,N_9203);
or U9777 (N_9777,N_9033,N_9257);
xor U9778 (N_9778,N_9450,N_9206);
xor U9779 (N_9779,N_9077,N_9198);
or U9780 (N_9780,N_9113,N_9287);
nor U9781 (N_9781,N_9011,N_9413);
or U9782 (N_9782,N_9277,N_9236);
and U9783 (N_9783,N_9372,N_9118);
and U9784 (N_9784,N_9329,N_9380);
xor U9785 (N_9785,N_9497,N_9185);
and U9786 (N_9786,N_9331,N_9421);
or U9787 (N_9787,N_9208,N_9241);
or U9788 (N_9788,N_9498,N_9221);
nand U9789 (N_9789,N_9358,N_9492);
and U9790 (N_9790,N_9279,N_9156);
and U9791 (N_9791,N_9474,N_9236);
nand U9792 (N_9792,N_9119,N_9037);
nor U9793 (N_9793,N_9048,N_9295);
and U9794 (N_9794,N_9325,N_9273);
nor U9795 (N_9795,N_9481,N_9082);
and U9796 (N_9796,N_9143,N_9222);
or U9797 (N_9797,N_9215,N_9078);
or U9798 (N_9798,N_9134,N_9443);
or U9799 (N_9799,N_9130,N_9306);
or U9800 (N_9800,N_9332,N_9364);
or U9801 (N_9801,N_9059,N_9200);
xor U9802 (N_9802,N_9310,N_9126);
and U9803 (N_9803,N_9089,N_9270);
or U9804 (N_9804,N_9127,N_9484);
nor U9805 (N_9805,N_9022,N_9351);
or U9806 (N_9806,N_9482,N_9075);
and U9807 (N_9807,N_9082,N_9145);
nor U9808 (N_9808,N_9476,N_9076);
xor U9809 (N_9809,N_9155,N_9123);
or U9810 (N_9810,N_9444,N_9124);
nand U9811 (N_9811,N_9335,N_9063);
and U9812 (N_9812,N_9282,N_9391);
nand U9813 (N_9813,N_9487,N_9337);
and U9814 (N_9814,N_9316,N_9031);
and U9815 (N_9815,N_9290,N_9228);
xor U9816 (N_9816,N_9150,N_9184);
nor U9817 (N_9817,N_9012,N_9448);
and U9818 (N_9818,N_9254,N_9190);
nand U9819 (N_9819,N_9482,N_9476);
nor U9820 (N_9820,N_9125,N_9150);
nor U9821 (N_9821,N_9497,N_9382);
and U9822 (N_9822,N_9401,N_9285);
and U9823 (N_9823,N_9008,N_9214);
xor U9824 (N_9824,N_9385,N_9074);
and U9825 (N_9825,N_9424,N_9361);
xnor U9826 (N_9826,N_9423,N_9455);
nand U9827 (N_9827,N_9056,N_9072);
or U9828 (N_9828,N_9123,N_9210);
nor U9829 (N_9829,N_9004,N_9234);
nand U9830 (N_9830,N_9269,N_9373);
and U9831 (N_9831,N_9456,N_9276);
or U9832 (N_9832,N_9067,N_9363);
nor U9833 (N_9833,N_9350,N_9268);
nand U9834 (N_9834,N_9233,N_9208);
or U9835 (N_9835,N_9370,N_9177);
xnor U9836 (N_9836,N_9019,N_9008);
nand U9837 (N_9837,N_9118,N_9445);
and U9838 (N_9838,N_9019,N_9334);
nor U9839 (N_9839,N_9272,N_9004);
nand U9840 (N_9840,N_9109,N_9011);
nand U9841 (N_9841,N_9060,N_9430);
nand U9842 (N_9842,N_9149,N_9362);
xor U9843 (N_9843,N_9398,N_9092);
nor U9844 (N_9844,N_9392,N_9260);
nand U9845 (N_9845,N_9379,N_9384);
and U9846 (N_9846,N_9312,N_9177);
and U9847 (N_9847,N_9240,N_9008);
nor U9848 (N_9848,N_9152,N_9239);
nor U9849 (N_9849,N_9030,N_9050);
and U9850 (N_9850,N_9438,N_9382);
xnor U9851 (N_9851,N_9415,N_9109);
nand U9852 (N_9852,N_9136,N_9315);
nor U9853 (N_9853,N_9300,N_9306);
or U9854 (N_9854,N_9402,N_9291);
and U9855 (N_9855,N_9394,N_9159);
and U9856 (N_9856,N_9490,N_9140);
nand U9857 (N_9857,N_9227,N_9392);
and U9858 (N_9858,N_9314,N_9180);
nand U9859 (N_9859,N_9240,N_9138);
nor U9860 (N_9860,N_9077,N_9213);
nor U9861 (N_9861,N_9321,N_9166);
or U9862 (N_9862,N_9292,N_9179);
nand U9863 (N_9863,N_9158,N_9085);
and U9864 (N_9864,N_9490,N_9215);
nor U9865 (N_9865,N_9007,N_9172);
xnor U9866 (N_9866,N_9152,N_9124);
xnor U9867 (N_9867,N_9130,N_9186);
and U9868 (N_9868,N_9430,N_9024);
or U9869 (N_9869,N_9310,N_9092);
and U9870 (N_9870,N_9293,N_9312);
nor U9871 (N_9871,N_9002,N_9313);
or U9872 (N_9872,N_9075,N_9409);
nor U9873 (N_9873,N_9022,N_9315);
or U9874 (N_9874,N_9432,N_9258);
and U9875 (N_9875,N_9223,N_9246);
or U9876 (N_9876,N_9131,N_9215);
xnor U9877 (N_9877,N_9481,N_9097);
and U9878 (N_9878,N_9031,N_9384);
or U9879 (N_9879,N_9092,N_9155);
nand U9880 (N_9880,N_9060,N_9275);
and U9881 (N_9881,N_9036,N_9344);
or U9882 (N_9882,N_9246,N_9457);
nor U9883 (N_9883,N_9099,N_9100);
or U9884 (N_9884,N_9144,N_9338);
and U9885 (N_9885,N_9014,N_9353);
and U9886 (N_9886,N_9004,N_9030);
nand U9887 (N_9887,N_9154,N_9166);
and U9888 (N_9888,N_9016,N_9439);
and U9889 (N_9889,N_9272,N_9423);
nor U9890 (N_9890,N_9292,N_9313);
and U9891 (N_9891,N_9436,N_9474);
and U9892 (N_9892,N_9262,N_9317);
and U9893 (N_9893,N_9019,N_9268);
nand U9894 (N_9894,N_9069,N_9294);
nand U9895 (N_9895,N_9465,N_9097);
or U9896 (N_9896,N_9376,N_9093);
or U9897 (N_9897,N_9040,N_9055);
nand U9898 (N_9898,N_9439,N_9107);
xnor U9899 (N_9899,N_9352,N_9408);
nor U9900 (N_9900,N_9311,N_9273);
nand U9901 (N_9901,N_9278,N_9219);
or U9902 (N_9902,N_9045,N_9459);
nor U9903 (N_9903,N_9481,N_9049);
xnor U9904 (N_9904,N_9084,N_9258);
or U9905 (N_9905,N_9403,N_9390);
nor U9906 (N_9906,N_9089,N_9144);
or U9907 (N_9907,N_9183,N_9101);
and U9908 (N_9908,N_9042,N_9117);
and U9909 (N_9909,N_9084,N_9368);
nand U9910 (N_9910,N_9231,N_9324);
or U9911 (N_9911,N_9278,N_9361);
and U9912 (N_9912,N_9174,N_9113);
xnor U9913 (N_9913,N_9261,N_9156);
or U9914 (N_9914,N_9252,N_9174);
nand U9915 (N_9915,N_9453,N_9254);
and U9916 (N_9916,N_9460,N_9355);
or U9917 (N_9917,N_9157,N_9485);
or U9918 (N_9918,N_9160,N_9412);
nor U9919 (N_9919,N_9397,N_9425);
or U9920 (N_9920,N_9223,N_9485);
or U9921 (N_9921,N_9484,N_9243);
nor U9922 (N_9922,N_9405,N_9450);
nor U9923 (N_9923,N_9497,N_9252);
nor U9924 (N_9924,N_9497,N_9030);
nand U9925 (N_9925,N_9319,N_9247);
and U9926 (N_9926,N_9327,N_9489);
and U9927 (N_9927,N_9391,N_9269);
nor U9928 (N_9928,N_9188,N_9221);
and U9929 (N_9929,N_9027,N_9392);
nor U9930 (N_9930,N_9497,N_9266);
or U9931 (N_9931,N_9031,N_9030);
nand U9932 (N_9932,N_9484,N_9170);
or U9933 (N_9933,N_9497,N_9118);
and U9934 (N_9934,N_9188,N_9239);
nand U9935 (N_9935,N_9075,N_9388);
nand U9936 (N_9936,N_9138,N_9054);
and U9937 (N_9937,N_9029,N_9271);
nor U9938 (N_9938,N_9193,N_9323);
xnor U9939 (N_9939,N_9358,N_9148);
and U9940 (N_9940,N_9225,N_9317);
nand U9941 (N_9941,N_9306,N_9434);
and U9942 (N_9942,N_9335,N_9103);
and U9943 (N_9943,N_9429,N_9028);
or U9944 (N_9944,N_9150,N_9096);
nand U9945 (N_9945,N_9185,N_9161);
or U9946 (N_9946,N_9389,N_9324);
nor U9947 (N_9947,N_9485,N_9358);
nand U9948 (N_9948,N_9010,N_9285);
and U9949 (N_9949,N_9169,N_9364);
nand U9950 (N_9950,N_9493,N_9016);
or U9951 (N_9951,N_9192,N_9401);
nor U9952 (N_9952,N_9188,N_9352);
or U9953 (N_9953,N_9168,N_9496);
nand U9954 (N_9954,N_9402,N_9042);
and U9955 (N_9955,N_9314,N_9327);
nand U9956 (N_9956,N_9437,N_9126);
and U9957 (N_9957,N_9258,N_9015);
or U9958 (N_9958,N_9214,N_9088);
nand U9959 (N_9959,N_9455,N_9408);
or U9960 (N_9960,N_9391,N_9202);
or U9961 (N_9961,N_9270,N_9488);
or U9962 (N_9962,N_9036,N_9483);
nor U9963 (N_9963,N_9495,N_9232);
or U9964 (N_9964,N_9225,N_9340);
nor U9965 (N_9965,N_9140,N_9321);
and U9966 (N_9966,N_9066,N_9078);
nor U9967 (N_9967,N_9388,N_9085);
or U9968 (N_9968,N_9338,N_9015);
xor U9969 (N_9969,N_9295,N_9073);
xnor U9970 (N_9970,N_9153,N_9174);
or U9971 (N_9971,N_9319,N_9000);
xnor U9972 (N_9972,N_9256,N_9008);
or U9973 (N_9973,N_9101,N_9027);
nor U9974 (N_9974,N_9244,N_9404);
or U9975 (N_9975,N_9389,N_9067);
nor U9976 (N_9976,N_9059,N_9313);
nand U9977 (N_9977,N_9088,N_9381);
nand U9978 (N_9978,N_9445,N_9366);
nand U9979 (N_9979,N_9023,N_9199);
nor U9980 (N_9980,N_9106,N_9085);
nor U9981 (N_9981,N_9068,N_9010);
xor U9982 (N_9982,N_9492,N_9158);
and U9983 (N_9983,N_9153,N_9305);
or U9984 (N_9984,N_9175,N_9393);
nor U9985 (N_9985,N_9043,N_9202);
nor U9986 (N_9986,N_9248,N_9360);
and U9987 (N_9987,N_9142,N_9196);
or U9988 (N_9988,N_9286,N_9093);
and U9989 (N_9989,N_9264,N_9313);
and U9990 (N_9990,N_9229,N_9206);
nor U9991 (N_9991,N_9123,N_9419);
or U9992 (N_9992,N_9068,N_9368);
or U9993 (N_9993,N_9298,N_9305);
nor U9994 (N_9994,N_9053,N_9235);
xor U9995 (N_9995,N_9380,N_9251);
nand U9996 (N_9996,N_9135,N_9291);
nand U9997 (N_9997,N_9123,N_9207);
nand U9998 (N_9998,N_9340,N_9234);
xnor U9999 (N_9999,N_9002,N_9374);
and UO_0 (O_0,N_9619,N_9655);
nand UO_1 (O_1,N_9736,N_9600);
nor UO_2 (O_2,N_9886,N_9917);
nand UO_3 (O_3,N_9972,N_9591);
nor UO_4 (O_4,N_9661,N_9968);
or UO_5 (O_5,N_9855,N_9926);
or UO_6 (O_6,N_9740,N_9808);
nor UO_7 (O_7,N_9509,N_9675);
or UO_8 (O_8,N_9853,N_9759);
and UO_9 (O_9,N_9648,N_9801);
and UO_10 (O_10,N_9758,N_9515);
and UO_11 (O_11,N_9962,N_9838);
and UO_12 (O_12,N_9575,N_9942);
nor UO_13 (O_13,N_9796,N_9843);
nor UO_14 (O_14,N_9522,N_9870);
nor UO_15 (O_15,N_9680,N_9896);
nor UO_16 (O_16,N_9948,N_9679);
nand UO_17 (O_17,N_9792,N_9845);
nor UO_18 (O_18,N_9703,N_9863);
nor UO_19 (O_19,N_9724,N_9623);
and UO_20 (O_20,N_9780,N_9745);
xnor UO_21 (O_21,N_9852,N_9577);
or UO_22 (O_22,N_9606,N_9588);
and UO_23 (O_23,N_9663,N_9586);
or UO_24 (O_24,N_9932,N_9873);
nor UO_25 (O_25,N_9563,N_9860);
or UO_26 (O_26,N_9894,N_9971);
nand UO_27 (O_27,N_9823,N_9597);
and UO_28 (O_28,N_9874,N_9766);
xnor UO_29 (O_29,N_9908,N_9840);
or UO_30 (O_30,N_9535,N_9533);
xor UO_31 (O_31,N_9628,N_9634);
and UO_32 (O_32,N_9502,N_9632);
xnor UO_33 (O_33,N_9775,N_9543);
and UO_34 (O_34,N_9892,N_9990);
nand UO_35 (O_35,N_9985,N_9698);
and UO_36 (O_36,N_9903,N_9564);
nor UO_37 (O_37,N_9737,N_9817);
nand UO_38 (O_38,N_9620,N_9829);
or UO_39 (O_39,N_9975,N_9602);
xor UO_40 (O_40,N_9692,N_9658);
and UO_41 (O_41,N_9681,N_9691);
nand UO_42 (O_42,N_9982,N_9694);
xnor UO_43 (O_43,N_9621,N_9559);
or UO_44 (O_44,N_9517,N_9955);
xnor UO_45 (O_45,N_9704,N_9640);
nand UO_46 (O_46,N_9572,N_9866);
nor UO_47 (O_47,N_9888,N_9919);
or UO_48 (O_48,N_9986,N_9773);
nor UO_49 (O_49,N_9929,N_9659);
or UO_50 (O_50,N_9776,N_9783);
and UO_51 (O_51,N_9754,N_9806);
nor UO_52 (O_52,N_9665,N_9699);
and UO_53 (O_53,N_9581,N_9654);
nand UO_54 (O_54,N_9700,N_9741);
nand UO_55 (O_55,N_9749,N_9842);
nand UO_56 (O_56,N_9925,N_9916);
nor UO_57 (O_57,N_9992,N_9904);
nor UO_58 (O_58,N_9707,N_9831);
and UO_59 (O_59,N_9733,N_9875);
nand UO_60 (O_60,N_9771,N_9539);
nand UO_61 (O_61,N_9798,N_9906);
nor UO_62 (O_62,N_9824,N_9983);
and UO_63 (O_63,N_9958,N_9551);
nor UO_64 (O_64,N_9996,N_9630);
and UO_65 (O_65,N_9593,N_9960);
nand UO_66 (O_66,N_9729,N_9697);
or UO_67 (O_67,N_9909,N_9585);
and UO_68 (O_68,N_9869,N_9604);
and UO_69 (O_69,N_9558,N_9701);
and UO_70 (O_70,N_9708,N_9565);
xor UO_71 (O_71,N_9599,N_9859);
nand UO_72 (O_72,N_9921,N_9877);
or UO_73 (O_73,N_9715,N_9684);
nand UO_74 (O_74,N_9998,N_9835);
nand UO_75 (O_75,N_9718,N_9850);
nor UO_76 (O_76,N_9614,N_9747);
or UO_77 (O_77,N_9503,N_9629);
and UO_78 (O_78,N_9910,N_9989);
xnor UO_79 (O_79,N_9978,N_9721);
nand UO_80 (O_80,N_9646,N_9893);
or UO_81 (O_81,N_9598,N_9887);
nor UO_82 (O_82,N_9664,N_9966);
and UO_83 (O_83,N_9936,N_9711);
and UO_84 (O_84,N_9651,N_9549);
and UO_85 (O_85,N_9956,N_9912);
nor UO_86 (O_86,N_9822,N_9653);
nand UO_87 (O_87,N_9935,N_9723);
or UO_88 (O_88,N_9770,N_9867);
nand UO_89 (O_89,N_9545,N_9809);
nor UO_90 (O_90,N_9889,N_9821);
or UO_91 (O_91,N_9899,N_9902);
or UO_92 (O_92,N_9952,N_9612);
nand UO_93 (O_93,N_9778,N_9927);
or UO_94 (O_94,N_9970,N_9947);
nand UO_95 (O_95,N_9964,N_9981);
nor UO_96 (O_96,N_9584,N_9616);
or UO_97 (O_97,N_9871,N_9514);
or UO_98 (O_98,N_9895,N_9524);
or UO_99 (O_99,N_9735,N_9748);
and UO_100 (O_100,N_9761,N_9650);
and UO_101 (O_101,N_9924,N_9594);
and UO_102 (O_102,N_9731,N_9969);
or UO_103 (O_103,N_9687,N_9764);
or UO_104 (O_104,N_9676,N_9945);
xor UO_105 (O_105,N_9529,N_9865);
nand UO_106 (O_106,N_9568,N_9580);
and UO_107 (O_107,N_9518,N_9790);
xnor UO_108 (O_108,N_9784,N_9841);
and UO_109 (O_109,N_9751,N_9541);
or UO_110 (O_110,N_9782,N_9878);
and UO_111 (O_111,N_9768,N_9803);
nand UO_112 (O_112,N_9526,N_9636);
nor UO_113 (O_113,N_9763,N_9941);
nand UO_114 (O_114,N_9819,N_9995);
nor UO_115 (O_115,N_9720,N_9795);
nand UO_116 (O_116,N_9846,N_9605);
and UO_117 (O_117,N_9712,N_9674);
and UO_118 (O_118,N_9561,N_9693);
or UO_119 (O_119,N_9501,N_9554);
or UO_120 (O_120,N_9574,N_9967);
and UO_121 (O_121,N_9552,N_9901);
and UO_122 (O_122,N_9557,N_9744);
nor UO_123 (O_123,N_9811,N_9802);
xnor UO_124 (O_124,N_9500,N_9911);
or UO_125 (O_125,N_9544,N_9789);
nand UO_126 (O_126,N_9622,N_9555);
nor UO_127 (O_127,N_9818,N_9923);
nor UO_128 (O_128,N_9856,N_9506);
and UO_129 (O_129,N_9530,N_9669);
nand UO_130 (O_130,N_9717,N_9825);
and UO_131 (O_131,N_9965,N_9772);
nor UO_132 (O_132,N_9938,N_9637);
or UO_133 (O_133,N_9510,N_9750);
nor UO_134 (O_134,N_9800,N_9611);
xnor UO_135 (O_135,N_9940,N_9984);
and UO_136 (O_136,N_9987,N_9848);
and UO_137 (O_137,N_9668,N_9576);
nand UO_138 (O_138,N_9710,N_9815);
nand UO_139 (O_139,N_9814,N_9579);
nand UO_140 (O_140,N_9713,N_9726);
nand UO_141 (O_141,N_9779,N_9949);
nor UO_142 (O_142,N_9900,N_9682);
nor UO_143 (O_143,N_9973,N_9787);
nand UO_144 (O_144,N_9596,N_9608);
or UO_145 (O_145,N_9706,N_9826);
or UO_146 (O_146,N_9880,N_9610);
or UO_147 (O_147,N_9666,N_9939);
and UO_148 (O_148,N_9647,N_9857);
nand UO_149 (O_149,N_9786,N_9953);
nor UO_150 (O_150,N_9553,N_9793);
or UO_151 (O_151,N_9864,N_9743);
nor UO_152 (O_152,N_9644,N_9891);
and UO_153 (O_153,N_9788,N_9702);
nor UO_154 (O_154,N_9851,N_9537);
nand UO_155 (O_155,N_9974,N_9872);
and UO_156 (O_156,N_9570,N_9876);
nand UO_157 (O_157,N_9999,N_9532);
nand UO_158 (O_158,N_9762,N_9667);
nand UO_159 (O_159,N_9977,N_9933);
or UO_160 (O_160,N_9635,N_9997);
and UO_161 (O_161,N_9858,N_9810);
nor UO_162 (O_162,N_9504,N_9673);
nor UO_163 (O_163,N_9813,N_9672);
nor UO_164 (O_164,N_9538,N_9677);
or UO_165 (O_165,N_9683,N_9799);
or UO_166 (O_166,N_9993,N_9862);
or UO_167 (O_167,N_9573,N_9915);
nand UO_168 (O_168,N_9950,N_9807);
and UO_169 (O_169,N_9678,N_9625);
or UO_170 (O_170,N_9930,N_9854);
and UO_171 (O_171,N_9617,N_9979);
and UO_172 (O_172,N_9928,N_9907);
or UO_173 (O_173,N_9719,N_9695);
or UO_174 (O_174,N_9905,N_9516);
or UO_175 (O_175,N_9734,N_9791);
nand UO_176 (O_176,N_9756,N_9785);
nand UO_177 (O_177,N_9918,N_9994);
nand UO_178 (O_178,N_9686,N_9660);
nor UO_179 (O_179,N_9550,N_9523);
nor UO_180 (O_180,N_9781,N_9671);
or UO_181 (O_181,N_9519,N_9587);
and UO_182 (O_182,N_9883,N_9601);
or UO_183 (O_183,N_9959,N_9649);
or UO_184 (O_184,N_9954,N_9582);
nand UO_185 (O_185,N_9957,N_9839);
nor UO_186 (O_186,N_9566,N_9547);
nor UO_187 (O_187,N_9583,N_9613);
nor UO_188 (O_188,N_9560,N_9988);
nand UO_189 (O_189,N_9777,N_9595);
nand UO_190 (O_190,N_9609,N_9847);
nand UO_191 (O_191,N_9820,N_9881);
xor UO_192 (O_192,N_9639,N_9615);
nand UO_193 (O_193,N_9805,N_9742);
or UO_194 (O_194,N_9511,N_9638);
or UO_195 (O_195,N_9879,N_9937);
nand UO_196 (O_196,N_9728,N_9657);
and UO_197 (O_197,N_9898,N_9688);
and UO_198 (O_198,N_9961,N_9944);
nor UO_199 (O_199,N_9951,N_9508);
and UO_200 (O_200,N_9589,N_9548);
nand UO_201 (O_201,N_9738,N_9830);
and UO_202 (O_202,N_9920,N_9836);
nor UO_203 (O_203,N_9963,N_9914);
nor UO_204 (O_204,N_9520,N_9753);
or UO_205 (O_205,N_9652,N_9714);
nand UO_206 (O_206,N_9643,N_9569);
nor UO_207 (O_207,N_9603,N_9844);
and UO_208 (O_208,N_9828,N_9837);
xnor UO_209 (O_209,N_9705,N_9882);
nand UO_210 (O_210,N_9774,N_9571);
nor UO_211 (O_211,N_9709,N_9833);
nor UO_212 (O_212,N_9722,N_9760);
xor UO_213 (O_213,N_9513,N_9897);
or UO_214 (O_214,N_9767,N_9505);
nor UO_215 (O_215,N_9567,N_9885);
nand UO_216 (O_216,N_9512,N_9527);
or UO_217 (O_217,N_9542,N_9562);
and UO_218 (O_218,N_9645,N_9834);
and UO_219 (O_219,N_9531,N_9757);
or UO_220 (O_220,N_9556,N_9943);
nand UO_221 (O_221,N_9578,N_9934);
nand UO_222 (O_222,N_9618,N_9642);
nand UO_223 (O_223,N_9525,N_9590);
and UO_224 (O_224,N_9922,N_9752);
and UO_225 (O_225,N_9507,N_9534);
or UO_226 (O_226,N_9546,N_9690);
nor UO_227 (O_227,N_9592,N_9528);
or UO_228 (O_228,N_9980,N_9746);
xnor UO_229 (O_229,N_9670,N_9849);
or UO_230 (O_230,N_9739,N_9991);
xor UO_231 (O_231,N_9816,N_9765);
or UO_232 (O_232,N_9656,N_9890);
nand UO_233 (O_233,N_9521,N_9861);
xnor UO_234 (O_234,N_9931,N_9755);
and UO_235 (O_235,N_9797,N_9976);
and UO_236 (O_236,N_9769,N_9804);
nor UO_237 (O_237,N_9730,N_9725);
nor UO_238 (O_238,N_9626,N_9540);
nand UO_239 (O_239,N_9827,N_9641);
and UO_240 (O_240,N_9832,N_9716);
xnor UO_241 (O_241,N_9689,N_9946);
and UO_242 (O_242,N_9884,N_9794);
nor UO_243 (O_243,N_9631,N_9627);
nand UO_244 (O_244,N_9696,N_9732);
nand UO_245 (O_245,N_9913,N_9536);
or UO_246 (O_246,N_9624,N_9607);
and UO_247 (O_247,N_9727,N_9633);
nor UO_248 (O_248,N_9662,N_9685);
or UO_249 (O_249,N_9868,N_9812);
nand UO_250 (O_250,N_9512,N_9714);
or UO_251 (O_251,N_9849,N_9763);
and UO_252 (O_252,N_9774,N_9522);
nor UO_253 (O_253,N_9854,N_9969);
or UO_254 (O_254,N_9700,N_9573);
nand UO_255 (O_255,N_9540,N_9761);
nor UO_256 (O_256,N_9751,N_9947);
nand UO_257 (O_257,N_9872,N_9700);
or UO_258 (O_258,N_9893,N_9568);
or UO_259 (O_259,N_9708,N_9837);
nor UO_260 (O_260,N_9801,N_9513);
nand UO_261 (O_261,N_9733,N_9660);
or UO_262 (O_262,N_9932,N_9564);
or UO_263 (O_263,N_9900,N_9585);
xnor UO_264 (O_264,N_9590,N_9870);
xor UO_265 (O_265,N_9662,N_9745);
or UO_266 (O_266,N_9988,N_9798);
and UO_267 (O_267,N_9532,N_9901);
nor UO_268 (O_268,N_9522,N_9734);
or UO_269 (O_269,N_9659,N_9717);
nand UO_270 (O_270,N_9671,N_9979);
or UO_271 (O_271,N_9814,N_9825);
or UO_272 (O_272,N_9997,N_9846);
or UO_273 (O_273,N_9856,N_9760);
nand UO_274 (O_274,N_9620,N_9897);
and UO_275 (O_275,N_9919,N_9763);
or UO_276 (O_276,N_9545,N_9833);
nand UO_277 (O_277,N_9638,N_9814);
nor UO_278 (O_278,N_9563,N_9688);
or UO_279 (O_279,N_9684,N_9700);
xnor UO_280 (O_280,N_9739,N_9596);
or UO_281 (O_281,N_9592,N_9638);
nand UO_282 (O_282,N_9552,N_9666);
nor UO_283 (O_283,N_9609,N_9763);
nor UO_284 (O_284,N_9785,N_9603);
nor UO_285 (O_285,N_9770,N_9981);
or UO_286 (O_286,N_9546,N_9731);
nand UO_287 (O_287,N_9938,N_9767);
nor UO_288 (O_288,N_9766,N_9909);
and UO_289 (O_289,N_9686,N_9573);
nand UO_290 (O_290,N_9731,N_9839);
nand UO_291 (O_291,N_9532,N_9971);
and UO_292 (O_292,N_9866,N_9534);
nand UO_293 (O_293,N_9723,N_9648);
or UO_294 (O_294,N_9512,N_9978);
nor UO_295 (O_295,N_9717,N_9744);
or UO_296 (O_296,N_9573,N_9688);
nand UO_297 (O_297,N_9804,N_9851);
nand UO_298 (O_298,N_9614,N_9834);
and UO_299 (O_299,N_9776,N_9775);
or UO_300 (O_300,N_9989,N_9827);
nand UO_301 (O_301,N_9613,N_9909);
or UO_302 (O_302,N_9725,N_9655);
nor UO_303 (O_303,N_9874,N_9774);
and UO_304 (O_304,N_9764,N_9688);
and UO_305 (O_305,N_9720,N_9638);
xnor UO_306 (O_306,N_9870,N_9706);
or UO_307 (O_307,N_9518,N_9868);
or UO_308 (O_308,N_9524,N_9902);
nor UO_309 (O_309,N_9610,N_9721);
or UO_310 (O_310,N_9520,N_9613);
and UO_311 (O_311,N_9748,N_9948);
and UO_312 (O_312,N_9536,N_9655);
nand UO_313 (O_313,N_9961,N_9752);
and UO_314 (O_314,N_9539,N_9672);
or UO_315 (O_315,N_9800,N_9805);
nand UO_316 (O_316,N_9974,N_9558);
nor UO_317 (O_317,N_9716,N_9917);
and UO_318 (O_318,N_9661,N_9914);
nand UO_319 (O_319,N_9735,N_9623);
and UO_320 (O_320,N_9525,N_9642);
xor UO_321 (O_321,N_9562,N_9624);
nand UO_322 (O_322,N_9530,N_9563);
or UO_323 (O_323,N_9511,N_9971);
and UO_324 (O_324,N_9537,N_9575);
nand UO_325 (O_325,N_9615,N_9562);
xnor UO_326 (O_326,N_9737,N_9863);
and UO_327 (O_327,N_9901,N_9694);
nand UO_328 (O_328,N_9917,N_9752);
nor UO_329 (O_329,N_9564,N_9955);
or UO_330 (O_330,N_9671,N_9597);
nor UO_331 (O_331,N_9570,N_9852);
and UO_332 (O_332,N_9956,N_9915);
xnor UO_333 (O_333,N_9559,N_9759);
nor UO_334 (O_334,N_9763,N_9746);
xor UO_335 (O_335,N_9998,N_9912);
or UO_336 (O_336,N_9766,N_9685);
nor UO_337 (O_337,N_9658,N_9591);
and UO_338 (O_338,N_9733,N_9768);
nand UO_339 (O_339,N_9822,N_9756);
and UO_340 (O_340,N_9507,N_9555);
or UO_341 (O_341,N_9605,N_9935);
nor UO_342 (O_342,N_9581,N_9750);
nor UO_343 (O_343,N_9773,N_9535);
nor UO_344 (O_344,N_9973,N_9610);
and UO_345 (O_345,N_9611,N_9778);
nand UO_346 (O_346,N_9977,N_9859);
nor UO_347 (O_347,N_9957,N_9549);
and UO_348 (O_348,N_9986,N_9538);
nand UO_349 (O_349,N_9793,N_9630);
or UO_350 (O_350,N_9851,N_9895);
and UO_351 (O_351,N_9982,N_9854);
xor UO_352 (O_352,N_9862,N_9822);
nand UO_353 (O_353,N_9674,N_9822);
nor UO_354 (O_354,N_9841,N_9647);
and UO_355 (O_355,N_9970,N_9784);
and UO_356 (O_356,N_9750,N_9615);
nand UO_357 (O_357,N_9921,N_9988);
or UO_358 (O_358,N_9958,N_9799);
and UO_359 (O_359,N_9797,N_9756);
nor UO_360 (O_360,N_9657,N_9719);
or UO_361 (O_361,N_9658,N_9592);
nand UO_362 (O_362,N_9823,N_9503);
and UO_363 (O_363,N_9695,N_9761);
or UO_364 (O_364,N_9912,N_9597);
nand UO_365 (O_365,N_9994,N_9621);
or UO_366 (O_366,N_9869,N_9929);
or UO_367 (O_367,N_9985,N_9614);
nand UO_368 (O_368,N_9776,N_9949);
xor UO_369 (O_369,N_9877,N_9620);
nor UO_370 (O_370,N_9837,N_9798);
nor UO_371 (O_371,N_9786,N_9694);
nor UO_372 (O_372,N_9917,N_9642);
or UO_373 (O_373,N_9745,N_9750);
and UO_374 (O_374,N_9702,N_9879);
nor UO_375 (O_375,N_9891,N_9517);
xor UO_376 (O_376,N_9587,N_9616);
nor UO_377 (O_377,N_9834,N_9737);
and UO_378 (O_378,N_9583,N_9715);
xor UO_379 (O_379,N_9815,N_9706);
nand UO_380 (O_380,N_9628,N_9820);
and UO_381 (O_381,N_9657,N_9945);
and UO_382 (O_382,N_9917,N_9625);
nand UO_383 (O_383,N_9633,N_9710);
nor UO_384 (O_384,N_9909,N_9684);
nor UO_385 (O_385,N_9707,N_9711);
nand UO_386 (O_386,N_9713,N_9656);
or UO_387 (O_387,N_9730,N_9700);
nand UO_388 (O_388,N_9822,N_9694);
xor UO_389 (O_389,N_9613,N_9862);
nor UO_390 (O_390,N_9975,N_9728);
nand UO_391 (O_391,N_9892,N_9559);
nor UO_392 (O_392,N_9713,N_9943);
nand UO_393 (O_393,N_9826,N_9732);
nor UO_394 (O_394,N_9526,N_9940);
or UO_395 (O_395,N_9551,N_9894);
nand UO_396 (O_396,N_9821,N_9716);
nand UO_397 (O_397,N_9881,N_9682);
and UO_398 (O_398,N_9580,N_9975);
nand UO_399 (O_399,N_9847,N_9768);
nor UO_400 (O_400,N_9605,N_9754);
or UO_401 (O_401,N_9927,N_9712);
xnor UO_402 (O_402,N_9890,N_9927);
xnor UO_403 (O_403,N_9575,N_9693);
or UO_404 (O_404,N_9571,N_9825);
and UO_405 (O_405,N_9763,N_9873);
xnor UO_406 (O_406,N_9792,N_9812);
and UO_407 (O_407,N_9578,N_9766);
or UO_408 (O_408,N_9824,N_9583);
xor UO_409 (O_409,N_9708,N_9652);
and UO_410 (O_410,N_9670,N_9723);
or UO_411 (O_411,N_9637,N_9623);
nand UO_412 (O_412,N_9872,N_9583);
or UO_413 (O_413,N_9986,N_9988);
xor UO_414 (O_414,N_9870,N_9980);
or UO_415 (O_415,N_9951,N_9853);
xor UO_416 (O_416,N_9632,N_9647);
and UO_417 (O_417,N_9881,N_9751);
or UO_418 (O_418,N_9858,N_9763);
nor UO_419 (O_419,N_9638,N_9913);
nor UO_420 (O_420,N_9635,N_9534);
nor UO_421 (O_421,N_9923,N_9934);
or UO_422 (O_422,N_9998,N_9944);
nor UO_423 (O_423,N_9727,N_9568);
and UO_424 (O_424,N_9810,N_9550);
or UO_425 (O_425,N_9921,N_9607);
and UO_426 (O_426,N_9565,N_9780);
and UO_427 (O_427,N_9569,N_9525);
or UO_428 (O_428,N_9732,N_9561);
nand UO_429 (O_429,N_9726,N_9611);
or UO_430 (O_430,N_9555,N_9830);
and UO_431 (O_431,N_9667,N_9821);
nand UO_432 (O_432,N_9763,N_9713);
and UO_433 (O_433,N_9774,N_9989);
and UO_434 (O_434,N_9544,N_9951);
nand UO_435 (O_435,N_9773,N_9835);
nor UO_436 (O_436,N_9814,N_9794);
nor UO_437 (O_437,N_9764,N_9674);
xor UO_438 (O_438,N_9884,N_9648);
nand UO_439 (O_439,N_9937,N_9576);
and UO_440 (O_440,N_9876,N_9646);
nand UO_441 (O_441,N_9643,N_9916);
nor UO_442 (O_442,N_9797,N_9678);
nor UO_443 (O_443,N_9562,N_9800);
and UO_444 (O_444,N_9841,N_9937);
nor UO_445 (O_445,N_9637,N_9773);
and UO_446 (O_446,N_9993,N_9555);
or UO_447 (O_447,N_9778,N_9801);
xnor UO_448 (O_448,N_9623,N_9924);
nand UO_449 (O_449,N_9518,N_9737);
or UO_450 (O_450,N_9658,N_9512);
nor UO_451 (O_451,N_9817,N_9883);
and UO_452 (O_452,N_9775,N_9916);
nor UO_453 (O_453,N_9796,N_9719);
nand UO_454 (O_454,N_9664,N_9989);
nand UO_455 (O_455,N_9868,N_9887);
nor UO_456 (O_456,N_9525,N_9611);
xor UO_457 (O_457,N_9550,N_9571);
or UO_458 (O_458,N_9541,N_9505);
and UO_459 (O_459,N_9513,N_9674);
nor UO_460 (O_460,N_9857,N_9992);
or UO_461 (O_461,N_9551,N_9562);
nor UO_462 (O_462,N_9724,N_9505);
and UO_463 (O_463,N_9559,N_9758);
or UO_464 (O_464,N_9741,N_9692);
and UO_465 (O_465,N_9811,N_9892);
nand UO_466 (O_466,N_9713,N_9894);
nand UO_467 (O_467,N_9821,N_9560);
nand UO_468 (O_468,N_9819,N_9973);
nor UO_469 (O_469,N_9879,N_9573);
nor UO_470 (O_470,N_9803,N_9550);
or UO_471 (O_471,N_9513,N_9887);
nor UO_472 (O_472,N_9754,N_9562);
xnor UO_473 (O_473,N_9648,N_9677);
nor UO_474 (O_474,N_9968,N_9617);
or UO_475 (O_475,N_9703,N_9902);
nand UO_476 (O_476,N_9634,N_9524);
or UO_477 (O_477,N_9653,N_9964);
and UO_478 (O_478,N_9941,N_9652);
or UO_479 (O_479,N_9736,N_9571);
and UO_480 (O_480,N_9984,N_9680);
nor UO_481 (O_481,N_9625,N_9851);
nand UO_482 (O_482,N_9787,N_9579);
or UO_483 (O_483,N_9631,N_9669);
nor UO_484 (O_484,N_9847,N_9913);
nor UO_485 (O_485,N_9680,N_9794);
and UO_486 (O_486,N_9936,N_9928);
nor UO_487 (O_487,N_9666,N_9811);
or UO_488 (O_488,N_9677,N_9504);
or UO_489 (O_489,N_9679,N_9984);
and UO_490 (O_490,N_9533,N_9659);
xor UO_491 (O_491,N_9633,N_9995);
and UO_492 (O_492,N_9668,N_9748);
or UO_493 (O_493,N_9866,N_9815);
nand UO_494 (O_494,N_9781,N_9641);
and UO_495 (O_495,N_9941,N_9542);
or UO_496 (O_496,N_9552,N_9681);
nand UO_497 (O_497,N_9851,N_9907);
nand UO_498 (O_498,N_9665,N_9837);
or UO_499 (O_499,N_9796,N_9679);
nand UO_500 (O_500,N_9572,N_9638);
nand UO_501 (O_501,N_9634,N_9869);
or UO_502 (O_502,N_9645,N_9788);
and UO_503 (O_503,N_9996,N_9892);
nand UO_504 (O_504,N_9750,N_9742);
and UO_505 (O_505,N_9714,N_9854);
nand UO_506 (O_506,N_9852,N_9943);
nand UO_507 (O_507,N_9848,N_9596);
or UO_508 (O_508,N_9680,N_9663);
xor UO_509 (O_509,N_9873,N_9675);
nor UO_510 (O_510,N_9717,N_9836);
and UO_511 (O_511,N_9900,N_9614);
nor UO_512 (O_512,N_9605,N_9529);
xor UO_513 (O_513,N_9932,N_9730);
xor UO_514 (O_514,N_9820,N_9559);
and UO_515 (O_515,N_9883,N_9912);
nand UO_516 (O_516,N_9665,N_9807);
nor UO_517 (O_517,N_9960,N_9955);
or UO_518 (O_518,N_9548,N_9979);
or UO_519 (O_519,N_9652,N_9741);
nand UO_520 (O_520,N_9737,N_9701);
and UO_521 (O_521,N_9559,N_9749);
and UO_522 (O_522,N_9820,N_9773);
or UO_523 (O_523,N_9990,N_9632);
xor UO_524 (O_524,N_9678,N_9624);
xor UO_525 (O_525,N_9550,N_9616);
or UO_526 (O_526,N_9519,N_9725);
nand UO_527 (O_527,N_9850,N_9838);
or UO_528 (O_528,N_9717,N_9745);
and UO_529 (O_529,N_9700,N_9883);
nand UO_530 (O_530,N_9596,N_9904);
nor UO_531 (O_531,N_9803,N_9869);
and UO_532 (O_532,N_9720,N_9784);
nor UO_533 (O_533,N_9995,N_9873);
or UO_534 (O_534,N_9768,N_9781);
nor UO_535 (O_535,N_9911,N_9902);
xor UO_536 (O_536,N_9934,N_9993);
nand UO_537 (O_537,N_9909,N_9857);
xnor UO_538 (O_538,N_9878,N_9552);
nand UO_539 (O_539,N_9839,N_9944);
xor UO_540 (O_540,N_9861,N_9778);
nor UO_541 (O_541,N_9824,N_9753);
or UO_542 (O_542,N_9765,N_9667);
and UO_543 (O_543,N_9641,N_9822);
xor UO_544 (O_544,N_9510,N_9549);
and UO_545 (O_545,N_9778,N_9649);
nor UO_546 (O_546,N_9761,N_9944);
and UO_547 (O_547,N_9607,N_9832);
xor UO_548 (O_548,N_9782,N_9588);
and UO_549 (O_549,N_9759,N_9788);
nor UO_550 (O_550,N_9997,N_9834);
or UO_551 (O_551,N_9717,N_9695);
and UO_552 (O_552,N_9911,N_9979);
or UO_553 (O_553,N_9760,N_9598);
or UO_554 (O_554,N_9961,N_9758);
or UO_555 (O_555,N_9695,N_9548);
nor UO_556 (O_556,N_9551,N_9737);
nand UO_557 (O_557,N_9638,N_9916);
nand UO_558 (O_558,N_9687,N_9906);
nor UO_559 (O_559,N_9640,N_9637);
nor UO_560 (O_560,N_9942,N_9523);
nand UO_561 (O_561,N_9801,N_9828);
nand UO_562 (O_562,N_9838,N_9595);
and UO_563 (O_563,N_9853,N_9720);
and UO_564 (O_564,N_9587,N_9540);
or UO_565 (O_565,N_9694,N_9819);
or UO_566 (O_566,N_9536,N_9901);
and UO_567 (O_567,N_9901,N_9574);
xnor UO_568 (O_568,N_9843,N_9791);
xor UO_569 (O_569,N_9567,N_9802);
or UO_570 (O_570,N_9512,N_9756);
and UO_571 (O_571,N_9781,N_9815);
or UO_572 (O_572,N_9908,N_9767);
nor UO_573 (O_573,N_9990,N_9579);
nor UO_574 (O_574,N_9631,N_9840);
or UO_575 (O_575,N_9624,N_9548);
or UO_576 (O_576,N_9963,N_9955);
and UO_577 (O_577,N_9821,N_9987);
nor UO_578 (O_578,N_9776,N_9971);
nand UO_579 (O_579,N_9988,N_9929);
xor UO_580 (O_580,N_9725,N_9794);
nor UO_581 (O_581,N_9998,N_9965);
and UO_582 (O_582,N_9794,N_9625);
or UO_583 (O_583,N_9965,N_9804);
xnor UO_584 (O_584,N_9632,N_9832);
and UO_585 (O_585,N_9562,N_9683);
nand UO_586 (O_586,N_9675,N_9555);
or UO_587 (O_587,N_9801,N_9623);
nor UO_588 (O_588,N_9998,N_9679);
nor UO_589 (O_589,N_9533,N_9598);
nand UO_590 (O_590,N_9582,N_9897);
nor UO_591 (O_591,N_9574,N_9713);
and UO_592 (O_592,N_9651,N_9544);
nor UO_593 (O_593,N_9808,N_9861);
nand UO_594 (O_594,N_9765,N_9810);
nand UO_595 (O_595,N_9797,N_9545);
and UO_596 (O_596,N_9894,N_9957);
or UO_597 (O_597,N_9697,N_9665);
or UO_598 (O_598,N_9819,N_9564);
or UO_599 (O_599,N_9735,N_9812);
or UO_600 (O_600,N_9775,N_9989);
nor UO_601 (O_601,N_9997,N_9641);
nor UO_602 (O_602,N_9667,N_9674);
and UO_603 (O_603,N_9589,N_9744);
or UO_604 (O_604,N_9947,N_9890);
xnor UO_605 (O_605,N_9764,N_9946);
and UO_606 (O_606,N_9722,N_9619);
nand UO_607 (O_607,N_9809,N_9771);
nand UO_608 (O_608,N_9889,N_9905);
xor UO_609 (O_609,N_9947,N_9909);
xor UO_610 (O_610,N_9913,N_9686);
and UO_611 (O_611,N_9649,N_9945);
or UO_612 (O_612,N_9725,N_9904);
and UO_613 (O_613,N_9756,N_9709);
or UO_614 (O_614,N_9504,N_9655);
nand UO_615 (O_615,N_9675,N_9668);
nor UO_616 (O_616,N_9684,N_9667);
xnor UO_617 (O_617,N_9538,N_9643);
nor UO_618 (O_618,N_9597,N_9585);
or UO_619 (O_619,N_9809,N_9932);
nand UO_620 (O_620,N_9875,N_9865);
nand UO_621 (O_621,N_9655,N_9537);
nor UO_622 (O_622,N_9626,N_9687);
nand UO_623 (O_623,N_9524,N_9938);
nand UO_624 (O_624,N_9671,N_9674);
and UO_625 (O_625,N_9593,N_9767);
or UO_626 (O_626,N_9682,N_9773);
nand UO_627 (O_627,N_9506,N_9593);
and UO_628 (O_628,N_9541,N_9923);
nand UO_629 (O_629,N_9643,N_9652);
nand UO_630 (O_630,N_9884,N_9672);
and UO_631 (O_631,N_9895,N_9626);
nand UO_632 (O_632,N_9912,N_9592);
nand UO_633 (O_633,N_9756,N_9887);
nand UO_634 (O_634,N_9717,N_9740);
nor UO_635 (O_635,N_9653,N_9899);
nand UO_636 (O_636,N_9910,N_9873);
nor UO_637 (O_637,N_9828,N_9604);
and UO_638 (O_638,N_9958,N_9949);
or UO_639 (O_639,N_9837,N_9620);
and UO_640 (O_640,N_9629,N_9776);
and UO_641 (O_641,N_9886,N_9777);
nand UO_642 (O_642,N_9828,N_9668);
nand UO_643 (O_643,N_9771,N_9932);
or UO_644 (O_644,N_9591,N_9815);
and UO_645 (O_645,N_9596,N_9826);
nor UO_646 (O_646,N_9979,N_9692);
and UO_647 (O_647,N_9969,N_9956);
or UO_648 (O_648,N_9558,N_9745);
or UO_649 (O_649,N_9754,N_9672);
or UO_650 (O_650,N_9904,N_9856);
or UO_651 (O_651,N_9998,N_9852);
nor UO_652 (O_652,N_9823,N_9884);
nor UO_653 (O_653,N_9975,N_9859);
nand UO_654 (O_654,N_9946,N_9846);
nor UO_655 (O_655,N_9792,N_9861);
nand UO_656 (O_656,N_9679,N_9599);
or UO_657 (O_657,N_9798,N_9885);
nor UO_658 (O_658,N_9673,N_9903);
nand UO_659 (O_659,N_9646,N_9791);
and UO_660 (O_660,N_9711,N_9943);
or UO_661 (O_661,N_9747,N_9765);
and UO_662 (O_662,N_9897,N_9667);
nand UO_663 (O_663,N_9974,N_9506);
nor UO_664 (O_664,N_9938,N_9758);
nand UO_665 (O_665,N_9801,N_9686);
nand UO_666 (O_666,N_9861,N_9628);
xor UO_667 (O_667,N_9895,N_9929);
nor UO_668 (O_668,N_9614,N_9786);
nand UO_669 (O_669,N_9832,N_9946);
nand UO_670 (O_670,N_9984,N_9924);
nand UO_671 (O_671,N_9857,N_9788);
nor UO_672 (O_672,N_9663,N_9532);
nand UO_673 (O_673,N_9583,N_9759);
nand UO_674 (O_674,N_9862,N_9556);
nand UO_675 (O_675,N_9527,N_9833);
or UO_676 (O_676,N_9638,N_9805);
or UO_677 (O_677,N_9806,N_9529);
or UO_678 (O_678,N_9920,N_9947);
or UO_679 (O_679,N_9531,N_9834);
nand UO_680 (O_680,N_9713,N_9559);
nor UO_681 (O_681,N_9832,N_9595);
or UO_682 (O_682,N_9648,N_9854);
nand UO_683 (O_683,N_9581,N_9852);
and UO_684 (O_684,N_9960,N_9626);
and UO_685 (O_685,N_9565,N_9963);
nor UO_686 (O_686,N_9556,N_9638);
nor UO_687 (O_687,N_9973,N_9577);
nor UO_688 (O_688,N_9678,N_9947);
nor UO_689 (O_689,N_9815,N_9844);
nor UO_690 (O_690,N_9967,N_9753);
nor UO_691 (O_691,N_9721,N_9983);
and UO_692 (O_692,N_9917,N_9946);
and UO_693 (O_693,N_9831,N_9895);
and UO_694 (O_694,N_9705,N_9760);
nor UO_695 (O_695,N_9881,N_9731);
or UO_696 (O_696,N_9938,N_9700);
or UO_697 (O_697,N_9808,N_9961);
nand UO_698 (O_698,N_9774,N_9867);
or UO_699 (O_699,N_9657,N_9861);
or UO_700 (O_700,N_9500,N_9890);
nand UO_701 (O_701,N_9869,N_9536);
or UO_702 (O_702,N_9887,N_9861);
nor UO_703 (O_703,N_9851,N_9991);
or UO_704 (O_704,N_9777,N_9761);
nand UO_705 (O_705,N_9603,N_9787);
nand UO_706 (O_706,N_9727,N_9786);
or UO_707 (O_707,N_9582,N_9913);
and UO_708 (O_708,N_9719,N_9784);
or UO_709 (O_709,N_9817,N_9984);
nand UO_710 (O_710,N_9761,N_9910);
or UO_711 (O_711,N_9658,N_9854);
xnor UO_712 (O_712,N_9785,N_9618);
nor UO_713 (O_713,N_9951,N_9960);
nand UO_714 (O_714,N_9617,N_9590);
and UO_715 (O_715,N_9782,N_9730);
and UO_716 (O_716,N_9573,N_9523);
xor UO_717 (O_717,N_9770,N_9598);
nor UO_718 (O_718,N_9706,N_9844);
nand UO_719 (O_719,N_9905,N_9933);
and UO_720 (O_720,N_9976,N_9873);
or UO_721 (O_721,N_9818,N_9577);
nand UO_722 (O_722,N_9722,N_9719);
or UO_723 (O_723,N_9504,N_9820);
xor UO_724 (O_724,N_9635,N_9881);
nor UO_725 (O_725,N_9891,N_9611);
or UO_726 (O_726,N_9744,N_9900);
nand UO_727 (O_727,N_9715,N_9555);
nor UO_728 (O_728,N_9887,N_9718);
nor UO_729 (O_729,N_9829,N_9541);
or UO_730 (O_730,N_9659,N_9828);
or UO_731 (O_731,N_9854,N_9729);
nand UO_732 (O_732,N_9777,N_9935);
or UO_733 (O_733,N_9597,N_9827);
and UO_734 (O_734,N_9658,N_9555);
xor UO_735 (O_735,N_9769,N_9665);
nor UO_736 (O_736,N_9564,N_9795);
and UO_737 (O_737,N_9815,N_9853);
or UO_738 (O_738,N_9515,N_9620);
or UO_739 (O_739,N_9901,N_9640);
or UO_740 (O_740,N_9729,N_9583);
nand UO_741 (O_741,N_9744,N_9929);
nor UO_742 (O_742,N_9578,N_9763);
and UO_743 (O_743,N_9624,N_9843);
or UO_744 (O_744,N_9683,N_9611);
and UO_745 (O_745,N_9705,N_9999);
nor UO_746 (O_746,N_9935,N_9776);
and UO_747 (O_747,N_9767,N_9564);
xor UO_748 (O_748,N_9725,N_9580);
and UO_749 (O_749,N_9993,N_9625);
nand UO_750 (O_750,N_9881,N_9533);
xor UO_751 (O_751,N_9842,N_9573);
or UO_752 (O_752,N_9642,N_9666);
nor UO_753 (O_753,N_9730,N_9791);
or UO_754 (O_754,N_9839,N_9656);
and UO_755 (O_755,N_9543,N_9650);
nor UO_756 (O_756,N_9950,N_9514);
and UO_757 (O_757,N_9623,N_9896);
nand UO_758 (O_758,N_9724,N_9918);
and UO_759 (O_759,N_9686,N_9525);
or UO_760 (O_760,N_9943,N_9933);
and UO_761 (O_761,N_9922,N_9703);
and UO_762 (O_762,N_9902,N_9713);
nand UO_763 (O_763,N_9701,N_9835);
or UO_764 (O_764,N_9821,N_9864);
and UO_765 (O_765,N_9560,N_9881);
nor UO_766 (O_766,N_9760,N_9549);
nand UO_767 (O_767,N_9834,N_9556);
xor UO_768 (O_768,N_9609,N_9911);
nor UO_769 (O_769,N_9956,N_9747);
and UO_770 (O_770,N_9561,N_9913);
and UO_771 (O_771,N_9891,N_9626);
nor UO_772 (O_772,N_9708,N_9534);
or UO_773 (O_773,N_9682,N_9850);
or UO_774 (O_774,N_9834,N_9813);
and UO_775 (O_775,N_9586,N_9781);
nand UO_776 (O_776,N_9576,N_9911);
or UO_777 (O_777,N_9570,N_9828);
or UO_778 (O_778,N_9548,N_9724);
nand UO_779 (O_779,N_9919,N_9760);
nand UO_780 (O_780,N_9522,N_9504);
xnor UO_781 (O_781,N_9932,N_9795);
and UO_782 (O_782,N_9848,N_9923);
and UO_783 (O_783,N_9883,N_9729);
and UO_784 (O_784,N_9794,N_9984);
and UO_785 (O_785,N_9947,N_9860);
or UO_786 (O_786,N_9524,N_9898);
nor UO_787 (O_787,N_9755,N_9764);
nand UO_788 (O_788,N_9792,N_9548);
nor UO_789 (O_789,N_9921,N_9763);
nand UO_790 (O_790,N_9940,N_9928);
and UO_791 (O_791,N_9525,N_9724);
or UO_792 (O_792,N_9704,N_9775);
and UO_793 (O_793,N_9547,N_9540);
nor UO_794 (O_794,N_9766,N_9616);
or UO_795 (O_795,N_9945,N_9813);
nor UO_796 (O_796,N_9974,N_9646);
nand UO_797 (O_797,N_9761,N_9845);
and UO_798 (O_798,N_9717,N_9634);
nor UO_799 (O_799,N_9622,N_9970);
nor UO_800 (O_800,N_9528,N_9764);
or UO_801 (O_801,N_9640,N_9563);
and UO_802 (O_802,N_9525,N_9500);
xnor UO_803 (O_803,N_9823,N_9943);
or UO_804 (O_804,N_9654,N_9889);
and UO_805 (O_805,N_9842,N_9832);
nand UO_806 (O_806,N_9946,N_9631);
and UO_807 (O_807,N_9911,N_9932);
or UO_808 (O_808,N_9646,N_9877);
and UO_809 (O_809,N_9783,N_9738);
and UO_810 (O_810,N_9667,N_9587);
or UO_811 (O_811,N_9944,N_9943);
or UO_812 (O_812,N_9985,N_9547);
or UO_813 (O_813,N_9950,N_9620);
and UO_814 (O_814,N_9615,N_9957);
and UO_815 (O_815,N_9716,N_9621);
and UO_816 (O_816,N_9857,N_9937);
nand UO_817 (O_817,N_9780,N_9812);
nand UO_818 (O_818,N_9710,N_9938);
nor UO_819 (O_819,N_9640,N_9753);
xor UO_820 (O_820,N_9778,N_9915);
nor UO_821 (O_821,N_9953,N_9519);
nand UO_822 (O_822,N_9964,N_9525);
nand UO_823 (O_823,N_9569,N_9505);
or UO_824 (O_824,N_9846,N_9732);
nor UO_825 (O_825,N_9593,N_9936);
or UO_826 (O_826,N_9949,N_9816);
or UO_827 (O_827,N_9805,N_9813);
or UO_828 (O_828,N_9797,N_9503);
nor UO_829 (O_829,N_9646,N_9778);
and UO_830 (O_830,N_9617,N_9953);
xor UO_831 (O_831,N_9575,N_9675);
and UO_832 (O_832,N_9945,N_9584);
or UO_833 (O_833,N_9801,N_9632);
nand UO_834 (O_834,N_9625,N_9850);
nand UO_835 (O_835,N_9855,N_9700);
or UO_836 (O_836,N_9738,N_9912);
nand UO_837 (O_837,N_9722,N_9716);
and UO_838 (O_838,N_9866,N_9975);
nor UO_839 (O_839,N_9805,N_9838);
and UO_840 (O_840,N_9899,N_9618);
and UO_841 (O_841,N_9660,N_9637);
xnor UO_842 (O_842,N_9532,N_9769);
xor UO_843 (O_843,N_9595,N_9961);
nand UO_844 (O_844,N_9673,N_9923);
nor UO_845 (O_845,N_9911,N_9735);
nand UO_846 (O_846,N_9996,N_9915);
nand UO_847 (O_847,N_9738,N_9743);
nor UO_848 (O_848,N_9872,N_9620);
nand UO_849 (O_849,N_9921,N_9842);
and UO_850 (O_850,N_9998,N_9895);
or UO_851 (O_851,N_9528,N_9987);
and UO_852 (O_852,N_9816,N_9679);
or UO_853 (O_853,N_9846,N_9693);
nor UO_854 (O_854,N_9627,N_9634);
and UO_855 (O_855,N_9760,N_9955);
and UO_856 (O_856,N_9547,N_9986);
nand UO_857 (O_857,N_9539,N_9572);
and UO_858 (O_858,N_9864,N_9784);
or UO_859 (O_859,N_9984,N_9603);
or UO_860 (O_860,N_9529,N_9992);
and UO_861 (O_861,N_9660,N_9525);
nor UO_862 (O_862,N_9741,N_9672);
nor UO_863 (O_863,N_9580,N_9935);
nor UO_864 (O_864,N_9504,N_9944);
or UO_865 (O_865,N_9744,N_9974);
nor UO_866 (O_866,N_9909,N_9657);
or UO_867 (O_867,N_9876,N_9885);
nand UO_868 (O_868,N_9680,N_9562);
and UO_869 (O_869,N_9743,N_9795);
nand UO_870 (O_870,N_9637,N_9675);
or UO_871 (O_871,N_9802,N_9699);
or UO_872 (O_872,N_9796,N_9658);
nor UO_873 (O_873,N_9795,N_9882);
xnor UO_874 (O_874,N_9945,N_9593);
or UO_875 (O_875,N_9680,N_9824);
nand UO_876 (O_876,N_9577,N_9640);
and UO_877 (O_877,N_9613,N_9917);
nor UO_878 (O_878,N_9697,N_9850);
nand UO_879 (O_879,N_9734,N_9868);
xnor UO_880 (O_880,N_9564,N_9849);
nand UO_881 (O_881,N_9697,N_9505);
or UO_882 (O_882,N_9837,N_9683);
nand UO_883 (O_883,N_9757,N_9682);
nor UO_884 (O_884,N_9561,N_9924);
nand UO_885 (O_885,N_9794,N_9632);
nand UO_886 (O_886,N_9561,N_9961);
or UO_887 (O_887,N_9570,N_9541);
or UO_888 (O_888,N_9952,N_9583);
and UO_889 (O_889,N_9673,N_9848);
or UO_890 (O_890,N_9600,N_9501);
nor UO_891 (O_891,N_9565,N_9806);
nor UO_892 (O_892,N_9816,N_9914);
xor UO_893 (O_893,N_9926,N_9546);
nand UO_894 (O_894,N_9740,N_9655);
xor UO_895 (O_895,N_9668,N_9637);
nor UO_896 (O_896,N_9622,N_9903);
nand UO_897 (O_897,N_9972,N_9801);
nand UO_898 (O_898,N_9788,N_9703);
nand UO_899 (O_899,N_9532,N_9750);
or UO_900 (O_900,N_9975,N_9680);
nor UO_901 (O_901,N_9546,N_9884);
nand UO_902 (O_902,N_9592,N_9692);
and UO_903 (O_903,N_9606,N_9524);
nand UO_904 (O_904,N_9969,N_9939);
or UO_905 (O_905,N_9642,N_9698);
or UO_906 (O_906,N_9657,N_9749);
nor UO_907 (O_907,N_9594,N_9940);
nor UO_908 (O_908,N_9880,N_9872);
nor UO_909 (O_909,N_9912,N_9825);
and UO_910 (O_910,N_9995,N_9855);
or UO_911 (O_911,N_9896,N_9688);
or UO_912 (O_912,N_9581,N_9841);
nand UO_913 (O_913,N_9921,N_9628);
xor UO_914 (O_914,N_9811,N_9810);
nor UO_915 (O_915,N_9522,N_9578);
nor UO_916 (O_916,N_9537,N_9816);
nand UO_917 (O_917,N_9628,N_9840);
or UO_918 (O_918,N_9753,N_9724);
and UO_919 (O_919,N_9882,N_9546);
and UO_920 (O_920,N_9987,N_9502);
and UO_921 (O_921,N_9678,N_9802);
nor UO_922 (O_922,N_9889,N_9822);
and UO_923 (O_923,N_9814,N_9521);
and UO_924 (O_924,N_9566,N_9750);
and UO_925 (O_925,N_9849,N_9673);
nor UO_926 (O_926,N_9719,N_9983);
nor UO_927 (O_927,N_9978,N_9932);
nand UO_928 (O_928,N_9954,N_9792);
nor UO_929 (O_929,N_9803,N_9780);
and UO_930 (O_930,N_9924,N_9520);
nor UO_931 (O_931,N_9522,N_9843);
nor UO_932 (O_932,N_9729,N_9681);
or UO_933 (O_933,N_9706,N_9828);
or UO_934 (O_934,N_9637,N_9647);
nor UO_935 (O_935,N_9694,N_9595);
or UO_936 (O_936,N_9774,N_9942);
and UO_937 (O_937,N_9763,N_9830);
nor UO_938 (O_938,N_9616,N_9657);
nand UO_939 (O_939,N_9969,N_9702);
or UO_940 (O_940,N_9896,N_9876);
and UO_941 (O_941,N_9950,N_9894);
and UO_942 (O_942,N_9969,N_9944);
nor UO_943 (O_943,N_9781,N_9881);
nor UO_944 (O_944,N_9752,N_9880);
nor UO_945 (O_945,N_9919,N_9513);
or UO_946 (O_946,N_9641,N_9983);
or UO_947 (O_947,N_9884,N_9644);
nor UO_948 (O_948,N_9732,N_9880);
nand UO_949 (O_949,N_9829,N_9825);
nor UO_950 (O_950,N_9807,N_9664);
nor UO_951 (O_951,N_9888,N_9972);
xnor UO_952 (O_952,N_9593,N_9610);
or UO_953 (O_953,N_9510,N_9875);
nor UO_954 (O_954,N_9961,N_9993);
nand UO_955 (O_955,N_9566,N_9533);
nor UO_956 (O_956,N_9575,N_9790);
or UO_957 (O_957,N_9979,N_9869);
and UO_958 (O_958,N_9756,N_9903);
nand UO_959 (O_959,N_9532,N_9851);
nand UO_960 (O_960,N_9943,N_9843);
nand UO_961 (O_961,N_9605,N_9988);
or UO_962 (O_962,N_9563,N_9924);
nor UO_963 (O_963,N_9585,N_9513);
xnor UO_964 (O_964,N_9968,N_9782);
or UO_965 (O_965,N_9703,N_9947);
or UO_966 (O_966,N_9597,N_9543);
and UO_967 (O_967,N_9971,N_9672);
and UO_968 (O_968,N_9672,N_9856);
and UO_969 (O_969,N_9937,N_9631);
or UO_970 (O_970,N_9678,N_9569);
nor UO_971 (O_971,N_9850,N_9642);
nand UO_972 (O_972,N_9578,N_9923);
or UO_973 (O_973,N_9857,N_9878);
or UO_974 (O_974,N_9616,N_9737);
or UO_975 (O_975,N_9833,N_9955);
or UO_976 (O_976,N_9895,N_9959);
and UO_977 (O_977,N_9831,N_9642);
nand UO_978 (O_978,N_9864,N_9871);
or UO_979 (O_979,N_9648,N_9903);
and UO_980 (O_980,N_9645,N_9725);
nor UO_981 (O_981,N_9716,N_9565);
and UO_982 (O_982,N_9889,N_9974);
and UO_983 (O_983,N_9910,N_9809);
xor UO_984 (O_984,N_9990,N_9707);
nor UO_985 (O_985,N_9705,N_9550);
or UO_986 (O_986,N_9963,N_9979);
or UO_987 (O_987,N_9683,N_9952);
nor UO_988 (O_988,N_9810,N_9968);
nand UO_989 (O_989,N_9858,N_9666);
or UO_990 (O_990,N_9550,N_9765);
and UO_991 (O_991,N_9682,N_9610);
or UO_992 (O_992,N_9711,N_9714);
nand UO_993 (O_993,N_9901,N_9835);
and UO_994 (O_994,N_9923,N_9762);
nand UO_995 (O_995,N_9869,N_9851);
nand UO_996 (O_996,N_9911,N_9887);
nor UO_997 (O_997,N_9602,N_9848);
nand UO_998 (O_998,N_9949,N_9672);
or UO_999 (O_999,N_9589,N_9773);
or UO_1000 (O_1000,N_9576,N_9888);
or UO_1001 (O_1001,N_9604,N_9993);
nor UO_1002 (O_1002,N_9954,N_9538);
and UO_1003 (O_1003,N_9558,N_9960);
or UO_1004 (O_1004,N_9658,N_9519);
nand UO_1005 (O_1005,N_9706,N_9930);
nand UO_1006 (O_1006,N_9561,N_9642);
nor UO_1007 (O_1007,N_9776,N_9651);
or UO_1008 (O_1008,N_9782,N_9650);
or UO_1009 (O_1009,N_9702,N_9916);
and UO_1010 (O_1010,N_9534,N_9910);
or UO_1011 (O_1011,N_9577,N_9723);
or UO_1012 (O_1012,N_9956,N_9576);
nand UO_1013 (O_1013,N_9972,N_9692);
nand UO_1014 (O_1014,N_9621,N_9670);
nand UO_1015 (O_1015,N_9530,N_9564);
nand UO_1016 (O_1016,N_9677,N_9739);
nand UO_1017 (O_1017,N_9769,N_9943);
and UO_1018 (O_1018,N_9983,N_9717);
nor UO_1019 (O_1019,N_9863,N_9528);
nand UO_1020 (O_1020,N_9533,N_9555);
nand UO_1021 (O_1021,N_9615,N_9855);
and UO_1022 (O_1022,N_9745,N_9960);
nand UO_1023 (O_1023,N_9897,N_9718);
xnor UO_1024 (O_1024,N_9797,N_9980);
and UO_1025 (O_1025,N_9975,N_9615);
and UO_1026 (O_1026,N_9686,N_9547);
nand UO_1027 (O_1027,N_9528,N_9946);
nor UO_1028 (O_1028,N_9567,N_9828);
nor UO_1029 (O_1029,N_9755,N_9989);
xnor UO_1030 (O_1030,N_9869,N_9594);
and UO_1031 (O_1031,N_9767,N_9588);
or UO_1032 (O_1032,N_9685,N_9965);
xnor UO_1033 (O_1033,N_9741,N_9974);
nor UO_1034 (O_1034,N_9622,N_9706);
and UO_1035 (O_1035,N_9879,N_9819);
or UO_1036 (O_1036,N_9964,N_9640);
nand UO_1037 (O_1037,N_9912,N_9719);
nor UO_1038 (O_1038,N_9707,N_9649);
xnor UO_1039 (O_1039,N_9839,N_9605);
or UO_1040 (O_1040,N_9645,N_9904);
or UO_1041 (O_1041,N_9554,N_9790);
and UO_1042 (O_1042,N_9872,N_9604);
and UO_1043 (O_1043,N_9812,N_9927);
and UO_1044 (O_1044,N_9585,N_9680);
xnor UO_1045 (O_1045,N_9534,N_9982);
and UO_1046 (O_1046,N_9578,N_9736);
or UO_1047 (O_1047,N_9590,N_9744);
or UO_1048 (O_1048,N_9985,N_9952);
nor UO_1049 (O_1049,N_9663,N_9708);
or UO_1050 (O_1050,N_9570,N_9729);
and UO_1051 (O_1051,N_9508,N_9563);
and UO_1052 (O_1052,N_9584,N_9639);
nor UO_1053 (O_1053,N_9764,N_9914);
or UO_1054 (O_1054,N_9739,N_9654);
nand UO_1055 (O_1055,N_9941,N_9564);
and UO_1056 (O_1056,N_9667,N_9656);
xor UO_1057 (O_1057,N_9717,N_9612);
nor UO_1058 (O_1058,N_9538,N_9834);
and UO_1059 (O_1059,N_9867,N_9933);
nand UO_1060 (O_1060,N_9701,N_9593);
nand UO_1061 (O_1061,N_9901,N_9557);
or UO_1062 (O_1062,N_9581,N_9784);
nor UO_1063 (O_1063,N_9662,N_9816);
and UO_1064 (O_1064,N_9923,N_9985);
xnor UO_1065 (O_1065,N_9997,N_9714);
xor UO_1066 (O_1066,N_9656,N_9640);
nand UO_1067 (O_1067,N_9859,N_9519);
xnor UO_1068 (O_1068,N_9827,N_9900);
nand UO_1069 (O_1069,N_9584,N_9630);
xor UO_1070 (O_1070,N_9924,N_9975);
or UO_1071 (O_1071,N_9562,N_9690);
and UO_1072 (O_1072,N_9854,N_9772);
nand UO_1073 (O_1073,N_9977,N_9698);
nand UO_1074 (O_1074,N_9535,N_9615);
nand UO_1075 (O_1075,N_9824,N_9778);
or UO_1076 (O_1076,N_9982,N_9821);
xnor UO_1077 (O_1077,N_9634,N_9671);
nor UO_1078 (O_1078,N_9985,N_9669);
or UO_1079 (O_1079,N_9763,N_9586);
nand UO_1080 (O_1080,N_9559,N_9960);
and UO_1081 (O_1081,N_9718,N_9601);
nand UO_1082 (O_1082,N_9939,N_9928);
or UO_1083 (O_1083,N_9757,N_9629);
nor UO_1084 (O_1084,N_9529,N_9956);
or UO_1085 (O_1085,N_9961,N_9791);
nor UO_1086 (O_1086,N_9606,N_9555);
and UO_1087 (O_1087,N_9500,N_9958);
nor UO_1088 (O_1088,N_9991,N_9790);
xor UO_1089 (O_1089,N_9842,N_9821);
nor UO_1090 (O_1090,N_9799,N_9953);
or UO_1091 (O_1091,N_9891,N_9822);
and UO_1092 (O_1092,N_9764,N_9646);
and UO_1093 (O_1093,N_9686,N_9772);
xnor UO_1094 (O_1094,N_9654,N_9613);
and UO_1095 (O_1095,N_9558,N_9607);
xor UO_1096 (O_1096,N_9860,N_9503);
nand UO_1097 (O_1097,N_9919,N_9817);
or UO_1098 (O_1098,N_9843,N_9514);
and UO_1099 (O_1099,N_9904,N_9953);
nor UO_1100 (O_1100,N_9544,N_9839);
and UO_1101 (O_1101,N_9668,N_9551);
nand UO_1102 (O_1102,N_9860,N_9534);
xor UO_1103 (O_1103,N_9793,N_9974);
and UO_1104 (O_1104,N_9592,N_9834);
xnor UO_1105 (O_1105,N_9738,N_9999);
nor UO_1106 (O_1106,N_9693,N_9680);
nor UO_1107 (O_1107,N_9777,N_9797);
or UO_1108 (O_1108,N_9793,N_9809);
nand UO_1109 (O_1109,N_9726,N_9687);
nand UO_1110 (O_1110,N_9638,N_9996);
nand UO_1111 (O_1111,N_9705,N_9519);
nand UO_1112 (O_1112,N_9580,N_9625);
nand UO_1113 (O_1113,N_9582,N_9858);
xor UO_1114 (O_1114,N_9682,N_9604);
or UO_1115 (O_1115,N_9714,N_9783);
or UO_1116 (O_1116,N_9936,N_9538);
xnor UO_1117 (O_1117,N_9779,N_9761);
nand UO_1118 (O_1118,N_9846,N_9819);
xor UO_1119 (O_1119,N_9673,N_9659);
or UO_1120 (O_1120,N_9726,N_9664);
nor UO_1121 (O_1121,N_9840,N_9799);
nor UO_1122 (O_1122,N_9862,N_9749);
and UO_1123 (O_1123,N_9942,N_9703);
or UO_1124 (O_1124,N_9834,N_9815);
xor UO_1125 (O_1125,N_9598,N_9543);
nand UO_1126 (O_1126,N_9685,N_9574);
or UO_1127 (O_1127,N_9501,N_9712);
nor UO_1128 (O_1128,N_9814,N_9963);
xnor UO_1129 (O_1129,N_9767,N_9625);
nor UO_1130 (O_1130,N_9800,N_9559);
nand UO_1131 (O_1131,N_9893,N_9823);
or UO_1132 (O_1132,N_9975,N_9757);
nand UO_1133 (O_1133,N_9507,N_9895);
nand UO_1134 (O_1134,N_9535,N_9912);
or UO_1135 (O_1135,N_9516,N_9712);
and UO_1136 (O_1136,N_9844,N_9646);
nand UO_1137 (O_1137,N_9606,N_9717);
nor UO_1138 (O_1138,N_9873,N_9706);
nor UO_1139 (O_1139,N_9634,N_9984);
nor UO_1140 (O_1140,N_9810,N_9913);
and UO_1141 (O_1141,N_9812,N_9580);
nand UO_1142 (O_1142,N_9733,N_9584);
and UO_1143 (O_1143,N_9956,N_9887);
and UO_1144 (O_1144,N_9835,N_9866);
nor UO_1145 (O_1145,N_9593,N_9771);
and UO_1146 (O_1146,N_9860,N_9675);
or UO_1147 (O_1147,N_9553,N_9534);
nand UO_1148 (O_1148,N_9669,N_9749);
nor UO_1149 (O_1149,N_9659,N_9642);
nand UO_1150 (O_1150,N_9861,N_9750);
nor UO_1151 (O_1151,N_9744,N_9568);
xor UO_1152 (O_1152,N_9611,N_9764);
or UO_1153 (O_1153,N_9836,N_9816);
and UO_1154 (O_1154,N_9714,N_9672);
nor UO_1155 (O_1155,N_9579,N_9783);
and UO_1156 (O_1156,N_9777,N_9712);
nand UO_1157 (O_1157,N_9983,N_9738);
or UO_1158 (O_1158,N_9814,N_9759);
nand UO_1159 (O_1159,N_9694,N_9686);
nand UO_1160 (O_1160,N_9853,N_9677);
or UO_1161 (O_1161,N_9516,N_9806);
and UO_1162 (O_1162,N_9987,N_9920);
xor UO_1163 (O_1163,N_9649,N_9708);
nor UO_1164 (O_1164,N_9756,N_9875);
or UO_1165 (O_1165,N_9821,N_9828);
or UO_1166 (O_1166,N_9755,N_9749);
nand UO_1167 (O_1167,N_9692,N_9913);
and UO_1168 (O_1168,N_9975,N_9750);
nor UO_1169 (O_1169,N_9823,N_9783);
nand UO_1170 (O_1170,N_9839,N_9958);
xor UO_1171 (O_1171,N_9954,N_9734);
nor UO_1172 (O_1172,N_9914,N_9739);
and UO_1173 (O_1173,N_9614,N_9809);
xnor UO_1174 (O_1174,N_9683,N_9766);
nand UO_1175 (O_1175,N_9985,N_9787);
or UO_1176 (O_1176,N_9632,N_9921);
nand UO_1177 (O_1177,N_9570,N_9835);
and UO_1178 (O_1178,N_9734,N_9995);
nand UO_1179 (O_1179,N_9986,N_9641);
nand UO_1180 (O_1180,N_9924,N_9988);
xor UO_1181 (O_1181,N_9807,N_9684);
xor UO_1182 (O_1182,N_9749,N_9981);
or UO_1183 (O_1183,N_9634,N_9708);
or UO_1184 (O_1184,N_9579,N_9700);
or UO_1185 (O_1185,N_9625,N_9954);
or UO_1186 (O_1186,N_9819,N_9864);
nand UO_1187 (O_1187,N_9685,N_9788);
and UO_1188 (O_1188,N_9769,N_9724);
nor UO_1189 (O_1189,N_9821,N_9919);
or UO_1190 (O_1190,N_9570,N_9647);
nand UO_1191 (O_1191,N_9776,N_9885);
nor UO_1192 (O_1192,N_9646,N_9969);
nand UO_1193 (O_1193,N_9925,N_9970);
xor UO_1194 (O_1194,N_9730,N_9560);
nor UO_1195 (O_1195,N_9851,N_9878);
nor UO_1196 (O_1196,N_9911,N_9741);
and UO_1197 (O_1197,N_9708,N_9614);
or UO_1198 (O_1198,N_9968,N_9852);
nand UO_1199 (O_1199,N_9936,N_9808);
nand UO_1200 (O_1200,N_9731,N_9748);
nand UO_1201 (O_1201,N_9868,N_9939);
nand UO_1202 (O_1202,N_9602,N_9805);
nor UO_1203 (O_1203,N_9700,N_9633);
or UO_1204 (O_1204,N_9538,N_9557);
or UO_1205 (O_1205,N_9643,N_9709);
nand UO_1206 (O_1206,N_9837,N_9841);
nand UO_1207 (O_1207,N_9841,N_9709);
and UO_1208 (O_1208,N_9554,N_9707);
nor UO_1209 (O_1209,N_9874,N_9964);
or UO_1210 (O_1210,N_9694,N_9550);
xor UO_1211 (O_1211,N_9956,N_9737);
nor UO_1212 (O_1212,N_9810,N_9544);
nor UO_1213 (O_1213,N_9593,N_9627);
or UO_1214 (O_1214,N_9890,N_9705);
nand UO_1215 (O_1215,N_9610,N_9542);
nand UO_1216 (O_1216,N_9923,N_9558);
or UO_1217 (O_1217,N_9979,N_9748);
nand UO_1218 (O_1218,N_9844,N_9976);
nor UO_1219 (O_1219,N_9907,N_9944);
and UO_1220 (O_1220,N_9802,N_9771);
nand UO_1221 (O_1221,N_9554,N_9969);
or UO_1222 (O_1222,N_9622,N_9798);
nor UO_1223 (O_1223,N_9839,N_9756);
nor UO_1224 (O_1224,N_9853,N_9628);
and UO_1225 (O_1225,N_9679,N_9758);
or UO_1226 (O_1226,N_9958,N_9830);
or UO_1227 (O_1227,N_9590,N_9881);
or UO_1228 (O_1228,N_9771,N_9753);
nor UO_1229 (O_1229,N_9843,N_9811);
nor UO_1230 (O_1230,N_9747,N_9906);
and UO_1231 (O_1231,N_9863,N_9950);
or UO_1232 (O_1232,N_9984,N_9587);
or UO_1233 (O_1233,N_9967,N_9715);
nor UO_1234 (O_1234,N_9763,N_9768);
or UO_1235 (O_1235,N_9778,N_9535);
or UO_1236 (O_1236,N_9776,N_9751);
or UO_1237 (O_1237,N_9643,N_9815);
nand UO_1238 (O_1238,N_9735,N_9701);
nand UO_1239 (O_1239,N_9966,N_9826);
nor UO_1240 (O_1240,N_9685,N_9817);
nor UO_1241 (O_1241,N_9643,N_9642);
nor UO_1242 (O_1242,N_9897,N_9595);
and UO_1243 (O_1243,N_9965,N_9516);
xnor UO_1244 (O_1244,N_9834,N_9947);
or UO_1245 (O_1245,N_9623,N_9844);
or UO_1246 (O_1246,N_9936,N_9535);
or UO_1247 (O_1247,N_9584,N_9649);
and UO_1248 (O_1248,N_9842,N_9557);
and UO_1249 (O_1249,N_9694,N_9806);
or UO_1250 (O_1250,N_9857,N_9673);
or UO_1251 (O_1251,N_9924,N_9615);
nor UO_1252 (O_1252,N_9607,N_9620);
nand UO_1253 (O_1253,N_9696,N_9835);
nand UO_1254 (O_1254,N_9807,N_9935);
nand UO_1255 (O_1255,N_9689,N_9851);
nor UO_1256 (O_1256,N_9963,N_9803);
and UO_1257 (O_1257,N_9730,N_9581);
nand UO_1258 (O_1258,N_9740,N_9949);
nor UO_1259 (O_1259,N_9903,N_9687);
and UO_1260 (O_1260,N_9574,N_9875);
nor UO_1261 (O_1261,N_9502,N_9659);
nand UO_1262 (O_1262,N_9632,N_9590);
and UO_1263 (O_1263,N_9502,N_9990);
nand UO_1264 (O_1264,N_9682,N_9509);
nor UO_1265 (O_1265,N_9710,N_9838);
xor UO_1266 (O_1266,N_9656,N_9843);
and UO_1267 (O_1267,N_9872,N_9988);
nand UO_1268 (O_1268,N_9806,N_9505);
or UO_1269 (O_1269,N_9969,N_9590);
and UO_1270 (O_1270,N_9559,N_9576);
nor UO_1271 (O_1271,N_9728,N_9750);
and UO_1272 (O_1272,N_9519,N_9882);
nor UO_1273 (O_1273,N_9683,N_9664);
xor UO_1274 (O_1274,N_9679,N_9884);
nor UO_1275 (O_1275,N_9502,N_9542);
or UO_1276 (O_1276,N_9846,N_9663);
nand UO_1277 (O_1277,N_9730,N_9787);
nand UO_1278 (O_1278,N_9880,N_9708);
and UO_1279 (O_1279,N_9927,N_9552);
nand UO_1280 (O_1280,N_9686,N_9735);
nand UO_1281 (O_1281,N_9601,N_9669);
xnor UO_1282 (O_1282,N_9986,N_9827);
and UO_1283 (O_1283,N_9685,N_9687);
nor UO_1284 (O_1284,N_9523,N_9580);
xnor UO_1285 (O_1285,N_9919,N_9673);
nand UO_1286 (O_1286,N_9862,N_9946);
and UO_1287 (O_1287,N_9609,N_9543);
or UO_1288 (O_1288,N_9772,N_9810);
nand UO_1289 (O_1289,N_9926,N_9837);
nor UO_1290 (O_1290,N_9621,N_9770);
nand UO_1291 (O_1291,N_9882,N_9834);
nand UO_1292 (O_1292,N_9773,N_9767);
or UO_1293 (O_1293,N_9991,N_9553);
xnor UO_1294 (O_1294,N_9810,N_9997);
and UO_1295 (O_1295,N_9769,N_9582);
xor UO_1296 (O_1296,N_9962,N_9716);
and UO_1297 (O_1297,N_9679,N_9875);
or UO_1298 (O_1298,N_9808,N_9911);
or UO_1299 (O_1299,N_9693,N_9625);
nor UO_1300 (O_1300,N_9873,N_9724);
xnor UO_1301 (O_1301,N_9702,N_9587);
and UO_1302 (O_1302,N_9514,N_9613);
or UO_1303 (O_1303,N_9855,N_9769);
nor UO_1304 (O_1304,N_9878,N_9884);
and UO_1305 (O_1305,N_9858,N_9640);
nor UO_1306 (O_1306,N_9753,N_9988);
or UO_1307 (O_1307,N_9809,N_9996);
nor UO_1308 (O_1308,N_9616,N_9644);
and UO_1309 (O_1309,N_9675,N_9764);
xnor UO_1310 (O_1310,N_9590,N_9634);
and UO_1311 (O_1311,N_9802,N_9901);
nand UO_1312 (O_1312,N_9615,N_9885);
nor UO_1313 (O_1313,N_9998,N_9979);
nor UO_1314 (O_1314,N_9714,N_9973);
and UO_1315 (O_1315,N_9590,N_9666);
and UO_1316 (O_1316,N_9584,N_9882);
nor UO_1317 (O_1317,N_9694,N_9580);
or UO_1318 (O_1318,N_9906,N_9719);
and UO_1319 (O_1319,N_9553,N_9786);
xnor UO_1320 (O_1320,N_9757,N_9899);
or UO_1321 (O_1321,N_9848,N_9813);
nor UO_1322 (O_1322,N_9976,N_9754);
and UO_1323 (O_1323,N_9632,N_9638);
xor UO_1324 (O_1324,N_9522,N_9884);
or UO_1325 (O_1325,N_9848,N_9925);
nor UO_1326 (O_1326,N_9550,N_9876);
or UO_1327 (O_1327,N_9762,N_9630);
nor UO_1328 (O_1328,N_9830,N_9829);
xnor UO_1329 (O_1329,N_9874,N_9894);
nand UO_1330 (O_1330,N_9563,N_9949);
or UO_1331 (O_1331,N_9836,N_9931);
and UO_1332 (O_1332,N_9727,N_9740);
nand UO_1333 (O_1333,N_9896,N_9760);
or UO_1334 (O_1334,N_9921,N_9703);
nand UO_1335 (O_1335,N_9826,N_9718);
or UO_1336 (O_1336,N_9810,N_9597);
nand UO_1337 (O_1337,N_9572,N_9702);
and UO_1338 (O_1338,N_9548,N_9697);
nor UO_1339 (O_1339,N_9872,N_9946);
nand UO_1340 (O_1340,N_9948,N_9931);
nand UO_1341 (O_1341,N_9947,N_9992);
nand UO_1342 (O_1342,N_9609,N_9942);
nor UO_1343 (O_1343,N_9999,N_9924);
and UO_1344 (O_1344,N_9899,N_9790);
or UO_1345 (O_1345,N_9522,N_9689);
and UO_1346 (O_1346,N_9774,N_9826);
nand UO_1347 (O_1347,N_9613,N_9794);
or UO_1348 (O_1348,N_9934,N_9567);
or UO_1349 (O_1349,N_9964,N_9588);
or UO_1350 (O_1350,N_9692,N_9624);
xnor UO_1351 (O_1351,N_9888,N_9785);
and UO_1352 (O_1352,N_9733,N_9596);
and UO_1353 (O_1353,N_9871,N_9715);
nor UO_1354 (O_1354,N_9740,N_9530);
and UO_1355 (O_1355,N_9742,N_9927);
nor UO_1356 (O_1356,N_9865,N_9901);
or UO_1357 (O_1357,N_9557,N_9762);
or UO_1358 (O_1358,N_9928,N_9983);
and UO_1359 (O_1359,N_9992,N_9932);
or UO_1360 (O_1360,N_9708,N_9670);
or UO_1361 (O_1361,N_9915,N_9589);
nand UO_1362 (O_1362,N_9638,N_9623);
nor UO_1363 (O_1363,N_9565,N_9581);
or UO_1364 (O_1364,N_9786,N_9842);
and UO_1365 (O_1365,N_9643,N_9653);
and UO_1366 (O_1366,N_9740,N_9928);
and UO_1367 (O_1367,N_9577,N_9769);
nor UO_1368 (O_1368,N_9625,N_9543);
or UO_1369 (O_1369,N_9546,N_9869);
or UO_1370 (O_1370,N_9550,N_9670);
xor UO_1371 (O_1371,N_9880,N_9777);
nand UO_1372 (O_1372,N_9755,N_9832);
or UO_1373 (O_1373,N_9709,N_9897);
or UO_1374 (O_1374,N_9987,N_9552);
nand UO_1375 (O_1375,N_9786,N_9709);
and UO_1376 (O_1376,N_9664,N_9994);
xnor UO_1377 (O_1377,N_9976,N_9962);
nand UO_1378 (O_1378,N_9607,N_9548);
and UO_1379 (O_1379,N_9506,N_9961);
nor UO_1380 (O_1380,N_9722,N_9846);
nand UO_1381 (O_1381,N_9769,N_9560);
nand UO_1382 (O_1382,N_9512,N_9992);
nand UO_1383 (O_1383,N_9622,N_9975);
nor UO_1384 (O_1384,N_9533,N_9574);
xnor UO_1385 (O_1385,N_9512,N_9987);
or UO_1386 (O_1386,N_9957,N_9518);
or UO_1387 (O_1387,N_9664,N_9631);
nand UO_1388 (O_1388,N_9761,N_9726);
and UO_1389 (O_1389,N_9526,N_9733);
and UO_1390 (O_1390,N_9555,N_9681);
nor UO_1391 (O_1391,N_9802,N_9885);
nand UO_1392 (O_1392,N_9767,N_9967);
or UO_1393 (O_1393,N_9694,N_9501);
and UO_1394 (O_1394,N_9837,N_9701);
nor UO_1395 (O_1395,N_9847,N_9659);
nand UO_1396 (O_1396,N_9754,N_9579);
or UO_1397 (O_1397,N_9580,N_9624);
and UO_1398 (O_1398,N_9823,N_9551);
and UO_1399 (O_1399,N_9721,N_9884);
and UO_1400 (O_1400,N_9839,N_9814);
and UO_1401 (O_1401,N_9790,N_9551);
xnor UO_1402 (O_1402,N_9626,N_9612);
and UO_1403 (O_1403,N_9925,N_9734);
and UO_1404 (O_1404,N_9916,N_9979);
nand UO_1405 (O_1405,N_9778,N_9790);
or UO_1406 (O_1406,N_9776,N_9833);
or UO_1407 (O_1407,N_9990,N_9549);
or UO_1408 (O_1408,N_9553,N_9804);
nand UO_1409 (O_1409,N_9629,N_9749);
nand UO_1410 (O_1410,N_9900,N_9730);
nand UO_1411 (O_1411,N_9992,N_9680);
or UO_1412 (O_1412,N_9987,N_9798);
nor UO_1413 (O_1413,N_9592,N_9596);
nor UO_1414 (O_1414,N_9894,N_9682);
or UO_1415 (O_1415,N_9935,N_9669);
or UO_1416 (O_1416,N_9586,N_9947);
or UO_1417 (O_1417,N_9638,N_9886);
or UO_1418 (O_1418,N_9959,N_9969);
nand UO_1419 (O_1419,N_9923,N_9707);
nor UO_1420 (O_1420,N_9630,N_9779);
and UO_1421 (O_1421,N_9686,N_9577);
nand UO_1422 (O_1422,N_9726,N_9767);
nand UO_1423 (O_1423,N_9743,N_9708);
or UO_1424 (O_1424,N_9858,N_9625);
nand UO_1425 (O_1425,N_9908,N_9816);
and UO_1426 (O_1426,N_9697,N_9809);
and UO_1427 (O_1427,N_9883,N_9661);
nor UO_1428 (O_1428,N_9806,N_9987);
or UO_1429 (O_1429,N_9917,N_9827);
and UO_1430 (O_1430,N_9652,N_9640);
and UO_1431 (O_1431,N_9981,N_9804);
and UO_1432 (O_1432,N_9798,N_9663);
and UO_1433 (O_1433,N_9582,N_9621);
and UO_1434 (O_1434,N_9618,N_9789);
nand UO_1435 (O_1435,N_9629,N_9676);
xor UO_1436 (O_1436,N_9931,N_9909);
nor UO_1437 (O_1437,N_9627,N_9723);
xor UO_1438 (O_1438,N_9801,N_9716);
and UO_1439 (O_1439,N_9523,N_9968);
and UO_1440 (O_1440,N_9999,N_9670);
nand UO_1441 (O_1441,N_9877,N_9783);
nand UO_1442 (O_1442,N_9586,N_9937);
xnor UO_1443 (O_1443,N_9607,N_9922);
nand UO_1444 (O_1444,N_9606,N_9735);
nand UO_1445 (O_1445,N_9920,N_9958);
nor UO_1446 (O_1446,N_9568,N_9977);
nor UO_1447 (O_1447,N_9964,N_9842);
and UO_1448 (O_1448,N_9996,N_9768);
or UO_1449 (O_1449,N_9595,N_9720);
nor UO_1450 (O_1450,N_9528,N_9790);
and UO_1451 (O_1451,N_9668,N_9647);
or UO_1452 (O_1452,N_9548,N_9500);
xor UO_1453 (O_1453,N_9855,N_9759);
or UO_1454 (O_1454,N_9644,N_9786);
nand UO_1455 (O_1455,N_9743,N_9837);
nand UO_1456 (O_1456,N_9811,N_9501);
and UO_1457 (O_1457,N_9872,N_9565);
and UO_1458 (O_1458,N_9854,N_9962);
or UO_1459 (O_1459,N_9676,N_9722);
nand UO_1460 (O_1460,N_9515,N_9505);
or UO_1461 (O_1461,N_9689,N_9544);
nor UO_1462 (O_1462,N_9541,N_9919);
and UO_1463 (O_1463,N_9958,N_9775);
nand UO_1464 (O_1464,N_9510,N_9832);
or UO_1465 (O_1465,N_9888,N_9857);
or UO_1466 (O_1466,N_9521,N_9737);
xor UO_1467 (O_1467,N_9811,N_9913);
nand UO_1468 (O_1468,N_9731,N_9834);
nor UO_1469 (O_1469,N_9607,N_9920);
nand UO_1470 (O_1470,N_9802,N_9965);
nor UO_1471 (O_1471,N_9750,N_9804);
and UO_1472 (O_1472,N_9932,N_9531);
nand UO_1473 (O_1473,N_9925,N_9777);
nand UO_1474 (O_1474,N_9937,N_9900);
and UO_1475 (O_1475,N_9775,N_9974);
nor UO_1476 (O_1476,N_9911,N_9738);
or UO_1477 (O_1477,N_9928,N_9714);
and UO_1478 (O_1478,N_9663,N_9852);
or UO_1479 (O_1479,N_9837,N_9519);
and UO_1480 (O_1480,N_9566,N_9692);
or UO_1481 (O_1481,N_9583,N_9931);
or UO_1482 (O_1482,N_9986,N_9616);
nor UO_1483 (O_1483,N_9738,N_9798);
nand UO_1484 (O_1484,N_9955,N_9891);
nand UO_1485 (O_1485,N_9993,N_9745);
nand UO_1486 (O_1486,N_9796,N_9551);
nor UO_1487 (O_1487,N_9725,N_9567);
nor UO_1488 (O_1488,N_9663,N_9960);
or UO_1489 (O_1489,N_9794,N_9667);
nor UO_1490 (O_1490,N_9596,N_9726);
and UO_1491 (O_1491,N_9804,N_9510);
nor UO_1492 (O_1492,N_9507,N_9715);
or UO_1493 (O_1493,N_9829,N_9682);
nand UO_1494 (O_1494,N_9865,N_9893);
xnor UO_1495 (O_1495,N_9855,N_9763);
and UO_1496 (O_1496,N_9799,N_9786);
and UO_1497 (O_1497,N_9513,N_9960);
nor UO_1498 (O_1498,N_9825,N_9994);
or UO_1499 (O_1499,N_9884,N_9879);
endmodule