module basic_500_3000_500_30_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_215,In_156);
nor U1 (N_1,In_285,In_35);
or U2 (N_2,In_149,In_408);
nand U3 (N_3,In_154,In_299);
nand U4 (N_4,In_270,In_324);
nor U5 (N_5,In_456,In_337);
and U6 (N_6,In_437,In_216);
nor U7 (N_7,In_90,In_231);
nand U8 (N_8,In_471,In_10);
and U9 (N_9,In_110,In_22);
or U10 (N_10,In_114,In_463);
nand U11 (N_11,In_201,In_21);
xnor U12 (N_12,In_58,In_125);
xnor U13 (N_13,In_448,In_61);
or U14 (N_14,In_287,In_459);
nor U15 (N_15,In_491,In_445);
xnor U16 (N_16,In_19,In_382);
and U17 (N_17,In_343,In_160);
and U18 (N_18,In_133,In_138);
and U19 (N_19,In_288,In_259);
nor U20 (N_20,In_248,In_2);
nor U21 (N_21,In_15,In_427);
or U22 (N_22,In_59,In_66);
nor U23 (N_23,In_196,In_129);
nand U24 (N_24,In_174,In_268);
nand U25 (N_25,In_481,In_69);
nand U26 (N_26,In_442,In_294);
and U27 (N_27,In_454,In_296);
nor U28 (N_28,In_419,In_6);
nor U29 (N_29,In_474,In_49);
nor U30 (N_30,In_464,In_495);
nor U31 (N_31,In_412,In_168);
and U32 (N_32,In_346,In_476);
xor U33 (N_33,In_109,In_339);
nand U34 (N_34,In_79,In_193);
xor U35 (N_35,In_54,In_390);
nor U36 (N_36,In_43,In_281);
or U37 (N_37,In_5,In_153);
xnor U38 (N_38,In_98,In_267);
and U39 (N_39,In_399,In_290);
nand U40 (N_40,In_189,In_473);
or U41 (N_41,In_104,In_391);
nand U42 (N_42,In_101,In_308);
nor U43 (N_43,In_327,In_465);
or U44 (N_44,In_468,In_276);
and U45 (N_45,In_317,In_127);
xor U46 (N_46,In_302,In_88);
nor U47 (N_47,In_275,In_432);
and U48 (N_48,In_254,In_374);
xor U49 (N_49,In_286,In_410);
nor U50 (N_50,In_210,In_207);
or U51 (N_51,In_148,In_284);
nand U52 (N_52,In_159,In_400);
xor U53 (N_53,In_365,In_393);
nor U54 (N_54,In_181,In_62);
nor U55 (N_55,In_3,In_177);
nand U56 (N_56,In_232,In_492);
nand U57 (N_57,In_426,In_440);
and U58 (N_58,In_124,In_175);
or U59 (N_59,In_84,In_455);
or U60 (N_60,In_352,In_439);
nand U61 (N_61,In_441,In_310);
or U62 (N_62,In_496,In_187);
or U63 (N_63,In_63,In_401);
or U64 (N_64,In_490,In_239);
nand U65 (N_65,In_306,In_165);
and U66 (N_66,In_394,In_244);
nand U67 (N_67,In_57,In_217);
or U68 (N_68,In_213,In_349);
nor U69 (N_69,In_146,In_141);
xnor U70 (N_70,In_199,In_81);
nand U71 (N_71,In_458,In_155);
nor U72 (N_72,In_258,In_85);
nand U73 (N_73,In_245,In_421);
xor U74 (N_74,In_184,In_424);
or U75 (N_75,In_326,In_227);
and U76 (N_76,In_253,In_23);
and U77 (N_77,In_416,In_345);
and U78 (N_78,In_182,In_344);
nor U79 (N_79,In_291,In_307);
nand U80 (N_80,In_485,In_369);
and U81 (N_81,In_18,In_354);
nor U82 (N_82,In_30,In_357);
nor U83 (N_83,In_122,In_484);
nor U84 (N_84,In_332,In_272);
nand U85 (N_85,In_33,In_257);
or U86 (N_86,In_222,In_397);
nor U87 (N_87,In_434,In_76);
nand U88 (N_88,In_100,In_13);
xnor U89 (N_89,In_261,In_48);
nand U90 (N_90,In_224,In_470);
xnor U91 (N_91,In_37,In_102);
xor U92 (N_92,In_255,In_355);
and U93 (N_93,In_1,In_309);
xor U94 (N_94,In_94,In_269);
and U95 (N_95,In_404,In_65);
and U96 (N_96,In_14,In_180);
or U97 (N_97,In_428,In_237);
nor U98 (N_98,In_411,In_420);
and U99 (N_99,In_73,In_55);
nand U100 (N_100,In_137,N_98);
nor U101 (N_101,In_359,In_42);
xor U102 (N_102,In_96,In_46);
and U103 (N_103,In_116,In_50);
and U104 (N_104,N_89,N_25);
or U105 (N_105,In_236,In_303);
nand U106 (N_106,In_120,In_277);
or U107 (N_107,N_93,In_147);
and U108 (N_108,In_134,In_403);
nand U109 (N_109,N_95,In_91);
nand U110 (N_110,In_220,In_142);
nor U111 (N_111,In_320,In_51);
nor U112 (N_112,In_319,In_368);
and U113 (N_113,In_435,N_96);
xnor U114 (N_114,In_370,In_353);
or U115 (N_115,N_27,N_79);
xor U116 (N_116,In_321,In_99);
nor U117 (N_117,In_25,In_67);
xnor U118 (N_118,In_242,In_95);
and U119 (N_119,N_77,In_162);
and U120 (N_120,In_386,N_78);
nor U121 (N_121,N_36,In_27);
xnor U122 (N_122,N_61,N_88);
xnor U123 (N_123,In_223,In_301);
and U124 (N_124,In_243,N_75);
nand U125 (N_125,In_383,In_388);
nor U126 (N_126,In_375,In_389);
xnor U127 (N_127,In_64,In_188);
nor U128 (N_128,In_499,In_493);
or U129 (N_129,In_163,N_38);
xnor U130 (N_130,N_8,N_40);
nand U131 (N_131,In_45,In_115);
xnor U132 (N_132,In_333,In_479);
xor U133 (N_133,N_1,N_73);
and U134 (N_134,N_21,In_415);
and U135 (N_135,N_67,In_170);
xor U136 (N_136,N_37,In_238);
or U137 (N_137,In_111,In_131);
and U138 (N_138,In_44,In_487);
and U139 (N_139,N_81,N_54);
xnor U140 (N_140,In_219,In_24);
nor U141 (N_141,In_38,In_422);
nor U142 (N_142,In_356,In_234);
or U143 (N_143,In_398,In_186);
or U144 (N_144,N_14,In_77);
and U145 (N_145,N_0,In_26);
nor U146 (N_146,In_430,In_225);
xor U147 (N_147,In_12,In_449);
nand U148 (N_148,In_380,In_497);
xor U149 (N_149,In_376,In_328);
and U150 (N_150,N_11,N_5);
nand U151 (N_151,N_92,In_392);
and U152 (N_152,In_52,In_452);
or U153 (N_153,N_83,N_45);
and U154 (N_154,N_55,In_71);
nand U155 (N_155,In_151,In_364);
nand U156 (N_156,In_233,In_203);
or U157 (N_157,N_47,In_477);
xnor U158 (N_158,In_264,N_71);
nor U159 (N_159,In_218,In_314);
nand U160 (N_160,In_443,In_208);
and U161 (N_161,In_7,In_9);
and U162 (N_162,In_300,N_59);
xor U163 (N_163,In_143,In_118);
or U164 (N_164,In_316,N_74);
nor U165 (N_165,In_209,N_51);
xnor U166 (N_166,In_250,N_42);
xnor U167 (N_167,In_282,N_70);
nor U168 (N_168,In_93,In_280);
or U169 (N_169,In_70,In_265);
and U170 (N_170,In_128,In_123);
nor U171 (N_171,In_32,In_358);
nor U172 (N_172,In_106,In_164);
or U173 (N_173,In_256,N_69);
xor U174 (N_174,N_57,In_498);
nand U175 (N_175,In_113,In_478);
nand U176 (N_176,N_34,N_43);
xor U177 (N_177,In_330,In_145);
or U178 (N_178,In_252,In_461);
nor U179 (N_179,In_289,N_28);
xnor U180 (N_180,In_246,In_409);
xor U181 (N_181,In_460,In_395);
nor U182 (N_182,N_49,N_62);
xnor U183 (N_183,In_466,In_431);
and U184 (N_184,In_16,In_34);
and U185 (N_185,In_447,N_3);
or U186 (N_186,N_56,In_108);
xnor U187 (N_187,N_97,In_486);
nand U188 (N_188,N_60,In_39);
xnor U189 (N_189,In_103,In_204);
and U190 (N_190,N_19,In_425);
or U191 (N_191,In_387,In_28);
and U192 (N_192,In_190,In_87);
or U193 (N_193,In_229,In_366);
and U194 (N_194,In_423,In_361);
nor U195 (N_195,In_407,In_329);
or U196 (N_196,In_367,In_402);
xnor U197 (N_197,In_489,N_6);
nor U198 (N_198,N_48,In_72);
nor U199 (N_199,In_323,In_417);
nand U200 (N_200,N_123,N_168);
nor U201 (N_201,In_274,N_126);
nand U202 (N_202,In_260,In_192);
nand U203 (N_203,In_271,In_214);
xor U204 (N_204,In_262,N_183);
or U205 (N_205,N_136,N_167);
xor U206 (N_206,In_97,In_273);
and U207 (N_207,In_17,In_313);
or U208 (N_208,N_90,N_151);
or U209 (N_209,N_143,In_292);
nor U210 (N_210,N_80,In_446);
nand U211 (N_211,In_132,N_178);
xor U212 (N_212,In_331,N_161);
or U213 (N_213,N_124,In_179);
nand U214 (N_214,N_130,In_247);
and U215 (N_215,In_305,N_29);
nor U216 (N_216,In_121,N_147);
xnor U217 (N_217,In_413,In_202);
and U218 (N_218,N_86,N_165);
or U219 (N_219,In_20,N_191);
nor U220 (N_220,N_105,In_212);
and U221 (N_221,In_467,N_32);
and U222 (N_222,N_194,In_166);
xnor U223 (N_223,In_167,N_177);
nand U224 (N_224,N_157,N_196);
and U225 (N_225,In_53,In_41);
nor U226 (N_226,N_142,N_64);
nor U227 (N_227,In_293,N_169);
or U228 (N_228,N_175,In_47);
and U229 (N_229,In_144,N_17);
xor U230 (N_230,N_186,In_475);
and U231 (N_231,In_342,In_4);
xnor U232 (N_232,In_117,N_188);
nand U233 (N_233,In_450,In_60);
xor U234 (N_234,N_199,N_18);
nor U235 (N_235,In_150,N_76);
nor U236 (N_236,N_102,N_192);
or U237 (N_237,In_347,In_436);
and U238 (N_238,N_132,N_138);
or U239 (N_239,In_195,In_206);
and U240 (N_240,N_35,In_295);
xnor U241 (N_241,N_190,In_172);
and U242 (N_242,In_371,In_322);
or U243 (N_243,In_176,In_11);
nand U244 (N_244,N_107,N_101);
or U245 (N_245,N_134,N_181);
nand U246 (N_246,In_157,In_480);
or U247 (N_247,N_31,N_148);
or U248 (N_248,In_75,N_68);
or U249 (N_249,N_153,N_137);
and U250 (N_250,N_30,In_341);
xnor U251 (N_251,In_183,N_65);
or U252 (N_252,N_146,N_185);
nor U253 (N_253,N_141,In_494);
nand U254 (N_254,N_133,N_135);
or U255 (N_255,In_266,In_278);
and U256 (N_256,N_116,N_63);
or U257 (N_257,In_315,N_52);
or U258 (N_258,N_125,In_198);
nand U259 (N_259,N_182,N_112);
and U260 (N_260,N_53,In_405);
and U261 (N_261,N_94,N_119);
nand U262 (N_262,In_200,In_78);
or U263 (N_263,In_251,N_2);
nor U264 (N_264,In_126,In_414);
or U265 (N_265,N_46,In_152);
xor U266 (N_266,In_482,In_338);
xor U267 (N_267,In_68,In_226);
nand U268 (N_268,In_453,In_241);
xor U269 (N_269,N_22,N_72);
and U270 (N_270,In_334,N_166);
or U271 (N_271,In_205,N_197);
nor U272 (N_272,In_488,N_131);
nand U273 (N_273,N_156,In_158);
nand U274 (N_274,N_103,N_170);
nand U275 (N_275,N_174,In_350);
xor U276 (N_276,In_36,In_107);
and U277 (N_277,N_33,N_149);
nand U278 (N_278,In_197,N_84);
nand U279 (N_279,N_23,N_198);
nand U280 (N_280,N_13,N_122);
nand U281 (N_281,N_4,In_283);
and U282 (N_282,N_104,In_82);
xnor U283 (N_283,In_185,N_12);
nand U284 (N_284,In_119,N_24);
nor U285 (N_285,N_85,In_384);
nand U286 (N_286,N_99,In_105);
or U287 (N_287,N_164,N_106);
and U288 (N_288,In_221,In_173);
nor U289 (N_289,N_127,In_396);
or U290 (N_290,In_31,N_50);
or U291 (N_291,In_444,In_240);
or U292 (N_292,N_139,N_82);
nor U293 (N_293,In_373,N_187);
and U294 (N_294,In_136,In_161);
and U295 (N_295,In_381,N_109);
or U296 (N_296,N_154,In_194);
nor U297 (N_297,In_318,In_348);
nand U298 (N_298,In_263,In_191);
nand U299 (N_299,N_7,In_363);
nor U300 (N_300,N_229,N_244);
xnor U301 (N_301,N_160,N_193);
xnor U302 (N_302,N_256,N_286);
or U303 (N_303,In_377,N_41);
xor U304 (N_304,N_252,N_214);
xnor U305 (N_305,In_335,In_418);
xnor U306 (N_306,N_163,N_129);
nor U307 (N_307,N_218,N_117);
and U308 (N_308,N_211,In_171);
or U309 (N_309,N_203,N_212);
nor U310 (N_310,N_276,N_222);
or U311 (N_311,N_152,In_135);
and U312 (N_312,N_227,N_208);
or U313 (N_313,N_294,In_112);
nand U314 (N_314,In_249,In_169);
and U315 (N_315,N_257,N_180);
or U316 (N_316,N_219,N_121);
and U317 (N_317,N_236,N_115);
xnor U318 (N_318,N_278,N_162);
or U319 (N_319,In_279,N_173);
xnor U320 (N_320,N_128,N_242);
xnor U321 (N_321,N_206,N_140);
nand U322 (N_322,In_379,N_66);
and U323 (N_323,N_113,In_228);
and U324 (N_324,N_282,N_44);
nand U325 (N_325,N_296,N_224);
xnor U326 (N_326,N_290,N_250);
nor U327 (N_327,N_20,N_246);
or U328 (N_328,In_378,N_189);
xor U329 (N_329,N_260,N_213);
nor U330 (N_330,In_140,In_372);
nor U331 (N_331,N_207,In_438);
and U332 (N_332,In_457,N_220);
or U333 (N_333,N_10,N_201);
nor U334 (N_334,In_89,N_120);
nand U335 (N_335,N_171,In_230);
nor U336 (N_336,N_289,N_248);
or U337 (N_337,In_178,N_172);
xor U338 (N_338,In_298,N_259);
xor U339 (N_339,N_91,N_299);
nand U340 (N_340,N_144,N_195);
xor U341 (N_341,N_235,In_462);
xor U342 (N_342,N_110,In_351);
nor U343 (N_343,In_139,In_469);
xor U344 (N_344,In_83,N_287);
nor U345 (N_345,In_29,N_145);
nand U346 (N_346,N_111,N_298);
nand U347 (N_347,N_251,N_273);
nor U348 (N_348,N_231,N_274);
or U349 (N_349,N_253,N_284);
xnor U350 (N_350,N_272,N_263);
nand U351 (N_351,N_247,N_184);
nor U352 (N_352,N_225,N_292);
xor U353 (N_353,N_205,In_311);
xor U354 (N_354,In_483,N_108);
xnor U355 (N_355,N_258,In_451);
and U356 (N_356,N_228,N_237);
nand U357 (N_357,N_39,N_150);
nand U358 (N_358,N_270,N_243);
nand U359 (N_359,N_155,N_262);
and U360 (N_360,In_86,N_9);
and U361 (N_361,N_176,N_269);
xnor U362 (N_362,N_261,N_275);
nand U363 (N_363,N_179,N_281);
nand U364 (N_364,N_114,In_429);
nand U365 (N_365,N_265,N_230);
and U366 (N_366,N_283,N_221);
and U367 (N_367,N_291,N_245);
and U368 (N_368,N_285,N_234);
nor U369 (N_369,In_360,N_271);
nor U370 (N_370,N_87,N_226);
xnor U371 (N_371,In_406,In_211);
nand U372 (N_372,N_240,In_325);
and U373 (N_373,In_362,In_92);
and U374 (N_374,N_158,In_312);
and U375 (N_375,N_15,In_8);
and U376 (N_376,N_266,N_209);
and U377 (N_377,N_254,N_238);
xnor U378 (N_378,N_26,N_295);
or U379 (N_379,In_40,In_80);
or U380 (N_380,N_280,N_215);
or U381 (N_381,In_304,N_202);
and U382 (N_382,N_58,In_340);
xor U383 (N_383,N_288,In_130);
and U384 (N_384,N_264,N_277);
or U385 (N_385,N_100,N_118);
and U386 (N_386,N_268,N_239);
or U387 (N_387,N_200,N_223);
or U388 (N_388,In_297,N_216);
or U389 (N_389,In_433,N_249);
or U390 (N_390,N_241,In_56);
nand U391 (N_391,N_232,N_255);
nor U392 (N_392,N_159,N_217);
nor U393 (N_393,In_385,N_16);
nor U394 (N_394,N_210,In_0);
nand U395 (N_395,In_235,In_74);
xor U396 (N_396,N_204,N_293);
and U397 (N_397,N_279,In_472);
nand U398 (N_398,N_297,N_267);
and U399 (N_399,In_336,N_233);
and U400 (N_400,N_397,N_359);
or U401 (N_401,N_339,N_357);
nand U402 (N_402,N_349,N_338);
nand U403 (N_403,N_307,N_389);
nor U404 (N_404,N_370,N_303);
xor U405 (N_405,N_316,N_396);
nor U406 (N_406,N_308,N_361);
nor U407 (N_407,N_333,N_358);
or U408 (N_408,N_385,N_393);
and U409 (N_409,N_345,N_356);
xnor U410 (N_410,N_350,N_337);
nor U411 (N_411,N_363,N_372);
and U412 (N_412,N_341,N_330);
nor U413 (N_413,N_381,N_335);
nand U414 (N_414,N_318,N_384);
or U415 (N_415,N_378,N_347);
nor U416 (N_416,N_394,N_355);
or U417 (N_417,N_353,N_329);
nor U418 (N_418,N_391,N_314);
xor U419 (N_419,N_386,N_312);
xor U420 (N_420,N_301,N_376);
nand U421 (N_421,N_354,N_327);
or U422 (N_422,N_374,N_371);
or U423 (N_423,N_323,N_383);
or U424 (N_424,N_342,N_368);
or U425 (N_425,N_328,N_336);
or U426 (N_426,N_380,N_352);
and U427 (N_427,N_364,N_321);
or U428 (N_428,N_319,N_399);
and U429 (N_429,N_346,N_324);
nor U430 (N_430,N_382,N_317);
or U431 (N_431,N_302,N_343);
or U432 (N_432,N_332,N_367);
nor U433 (N_433,N_390,N_348);
xor U434 (N_434,N_300,N_392);
or U435 (N_435,N_351,N_331);
xnor U436 (N_436,N_387,N_375);
nand U437 (N_437,N_369,N_310);
nor U438 (N_438,N_315,N_306);
nor U439 (N_439,N_395,N_377);
nand U440 (N_440,N_373,N_398);
nand U441 (N_441,N_344,N_304);
nand U442 (N_442,N_360,N_325);
nand U443 (N_443,N_362,N_326);
xor U444 (N_444,N_388,N_379);
or U445 (N_445,N_313,N_334);
nand U446 (N_446,N_322,N_365);
xnor U447 (N_447,N_309,N_305);
nand U448 (N_448,N_311,N_340);
nor U449 (N_449,N_320,N_366);
and U450 (N_450,N_354,N_312);
nand U451 (N_451,N_337,N_319);
xor U452 (N_452,N_374,N_359);
or U453 (N_453,N_322,N_376);
and U454 (N_454,N_394,N_379);
xnor U455 (N_455,N_314,N_310);
xor U456 (N_456,N_326,N_314);
nand U457 (N_457,N_386,N_323);
and U458 (N_458,N_383,N_361);
nand U459 (N_459,N_321,N_397);
nor U460 (N_460,N_357,N_380);
nor U461 (N_461,N_345,N_398);
nor U462 (N_462,N_371,N_318);
nor U463 (N_463,N_384,N_324);
xnor U464 (N_464,N_352,N_346);
and U465 (N_465,N_395,N_392);
nor U466 (N_466,N_317,N_357);
nand U467 (N_467,N_346,N_331);
nor U468 (N_468,N_386,N_315);
and U469 (N_469,N_304,N_360);
or U470 (N_470,N_384,N_397);
nand U471 (N_471,N_383,N_396);
xnor U472 (N_472,N_314,N_357);
or U473 (N_473,N_300,N_349);
or U474 (N_474,N_346,N_356);
or U475 (N_475,N_323,N_306);
nor U476 (N_476,N_346,N_340);
and U477 (N_477,N_327,N_373);
or U478 (N_478,N_351,N_359);
nor U479 (N_479,N_398,N_321);
or U480 (N_480,N_343,N_347);
xnor U481 (N_481,N_382,N_386);
nor U482 (N_482,N_337,N_363);
or U483 (N_483,N_397,N_346);
and U484 (N_484,N_365,N_391);
or U485 (N_485,N_362,N_345);
or U486 (N_486,N_311,N_369);
and U487 (N_487,N_390,N_384);
or U488 (N_488,N_337,N_320);
and U489 (N_489,N_395,N_312);
nor U490 (N_490,N_358,N_328);
xnor U491 (N_491,N_391,N_376);
xnor U492 (N_492,N_329,N_372);
nand U493 (N_493,N_349,N_372);
nand U494 (N_494,N_339,N_364);
nand U495 (N_495,N_397,N_322);
nor U496 (N_496,N_398,N_365);
nor U497 (N_497,N_389,N_328);
or U498 (N_498,N_334,N_365);
or U499 (N_499,N_364,N_322);
nand U500 (N_500,N_415,N_452);
xor U501 (N_501,N_445,N_407);
xor U502 (N_502,N_493,N_484);
xor U503 (N_503,N_435,N_444);
or U504 (N_504,N_454,N_431);
nor U505 (N_505,N_460,N_439);
nor U506 (N_506,N_489,N_464);
or U507 (N_507,N_455,N_462);
xor U508 (N_508,N_410,N_457);
and U509 (N_509,N_495,N_430);
and U510 (N_510,N_440,N_448);
and U511 (N_511,N_465,N_404);
xor U512 (N_512,N_429,N_483);
and U513 (N_513,N_478,N_411);
and U514 (N_514,N_432,N_419);
or U515 (N_515,N_461,N_469);
nor U516 (N_516,N_485,N_477);
and U517 (N_517,N_424,N_403);
nand U518 (N_518,N_491,N_417);
and U519 (N_519,N_458,N_436);
nand U520 (N_520,N_438,N_459);
nor U521 (N_521,N_408,N_447);
nor U522 (N_522,N_467,N_453);
or U523 (N_523,N_481,N_421);
xor U524 (N_524,N_437,N_473);
or U525 (N_525,N_413,N_456);
or U526 (N_526,N_423,N_488);
and U527 (N_527,N_426,N_442);
or U528 (N_528,N_482,N_497);
nor U529 (N_529,N_425,N_496);
or U530 (N_530,N_499,N_476);
or U531 (N_531,N_479,N_492);
xnor U532 (N_532,N_451,N_486);
nor U533 (N_533,N_498,N_428);
xnor U534 (N_534,N_468,N_409);
or U535 (N_535,N_480,N_414);
nand U536 (N_536,N_472,N_490);
nor U537 (N_537,N_418,N_475);
nor U538 (N_538,N_405,N_401);
and U539 (N_539,N_412,N_427);
xor U540 (N_540,N_422,N_487);
nor U541 (N_541,N_443,N_400);
nor U542 (N_542,N_449,N_474);
or U543 (N_543,N_402,N_433);
nor U544 (N_544,N_441,N_416);
nor U545 (N_545,N_450,N_466);
or U546 (N_546,N_494,N_406);
xnor U547 (N_547,N_470,N_446);
or U548 (N_548,N_434,N_463);
nor U549 (N_549,N_471,N_420);
xnor U550 (N_550,N_420,N_439);
xor U551 (N_551,N_483,N_433);
nand U552 (N_552,N_446,N_440);
and U553 (N_553,N_475,N_420);
nor U554 (N_554,N_487,N_404);
xor U555 (N_555,N_406,N_451);
xor U556 (N_556,N_492,N_481);
nor U557 (N_557,N_432,N_441);
nor U558 (N_558,N_481,N_485);
xnor U559 (N_559,N_440,N_416);
nand U560 (N_560,N_465,N_408);
xor U561 (N_561,N_483,N_428);
and U562 (N_562,N_484,N_468);
and U563 (N_563,N_409,N_403);
or U564 (N_564,N_475,N_446);
and U565 (N_565,N_455,N_490);
xor U566 (N_566,N_426,N_462);
nor U567 (N_567,N_432,N_467);
or U568 (N_568,N_425,N_429);
and U569 (N_569,N_432,N_445);
or U570 (N_570,N_484,N_471);
or U571 (N_571,N_411,N_462);
or U572 (N_572,N_468,N_458);
nor U573 (N_573,N_475,N_402);
or U574 (N_574,N_468,N_411);
nand U575 (N_575,N_431,N_483);
or U576 (N_576,N_483,N_408);
xnor U577 (N_577,N_494,N_416);
xnor U578 (N_578,N_426,N_494);
xor U579 (N_579,N_488,N_449);
xnor U580 (N_580,N_457,N_451);
nor U581 (N_581,N_434,N_417);
nor U582 (N_582,N_440,N_438);
and U583 (N_583,N_467,N_415);
nor U584 (N_584,N_405,N_460);
and U585 (N_585,N_473,N_407);
nand U586 (N_586,N_465,N_467);
or U587 (N_587,N_478,N_425);
or U588 (N_588,N_456,N_449);
xor U589 (N_589,N_447,N_473);
and U590 (N_590,N_413,N_484);
and U591 (N_591,N_459,N_474);
nor U592 (N_592,N_497,N_419);
xor U593 (N_593,N_416,N_474);
nand U594 (N_594,N_422,N_464);
xnor U595 (N_595,N_436,N_445);
or U596 (N_596,N_409,N_480);
nor U597 (N_597,N_424,N_470);
or U598 (N_598,N_460,N_480);
nor U599 (N_599,N_494,N_491);
or U600 (N_600,N_577,N_579);
nor U601 (N_601,N_552,N_580);
nand U602 (N_602,N_574,N_553);
or U603 (N_603,N_535,N_558);
or U604 (N_604,N_589,N_526);
or U605 (N_605,N_538,N_583);
or U606 (N_606,N_575,N_590);
and U607 (N_607,N_510,N_550);
nor U608 (N_608,N_508,N_528);
or U609 (N_609,N_554,N_505);
or U610 (N_610,N_547,N_507);
nand U611 (N_611,N_562,N_521);
or U612 (N_612,N_572,N_546);
and U613 (N_613,N_519,N_566);
and U614 (N_614,N_585,N_576);
xnor U615 (N_615,N_511,N_544);
and U616 (N_616,N_581,N_537);
nand U617 (N_617,N_500,N_536);
and U618 (N_618,N_549,N_570);
or U619 (N_619,N_565,N_520);
nand U620 (N_620,N_595,N_504);
xnor U621 (N_621,N_530,N_545);
or U622 (N_622,N_513,N_557);
or U623 (N_623,N_582,N_563);
nor U624 (N_624,N_541,N_517);
xor U625 (N_625,N_596,N_533);
nand U626 (N_626,N_534,N_543);
nor U627 (N_627,N_509,N_567);
nand U628 (N_628,N_542,N_512);
xor U629 (N_629,N_560,N_591);
nand U630 (N_630,N_523,N_559);
xor U631 (N_631,N_597,N_568);
nand U632 (N_632,N_503,N_569);
nand U633 (N_633,N_548,N_527);
nor U634 (N_634,N_564,N_522);
nor U635 (N_635,N_594,N_593);
nand U636 (N_636,N_514,N_571);
xnor U637 (N_637,N_586,N_525);
nand U638 (N_638,N_506,N_584);
nor U639 (N_639,N_531,N_529);
xnor U640 (N_640,N_578,N_598);
xor U641 (N_641,N_556,N_539);
xor U642 (N_642,N_573,N_592);
nor U643 (N_643,N_551,N_555);
or U644 (N_644,N_518,N_532);
nand U645 (N_645,N_524,N_599);
and U646 (N_646,N_587,N_540);
xnor U647 (N_647,N_516,N_588);
nand U648 (N_648,N_501,N_515);
and U649 (N_649,N_502,N_561);
or U650 (N_650,N_524,N_503);
and U651 (N_651,N_516,N_544);
or U652 (N_652,N_576,N_532);
and U653 (N_653,N_546,N_530);
xor U654 (N_654,N_564,N_582);
xor U655 (N_655,N_571,N_569);
xor U656 (N_656,N_584,N_521);
xor U657 (N_657,N_546,N_598);
or U658 (N_658,N_503,N_518);
xnor U659 (N_659,N_560,N_531);
nor U660 (N_660,N_597,N_596);
and U661 (N_661,N_549,N_584);
or U662 (N_662,N_503,N_510);
nor U663 (N_663,N_522,N_533);
nor U664 (N_664,N_510,N_584);
and U665 (N_665,N_578,N_517);
nand U666 (N_666,N_533,N_508);
nor U667 (N_667,N_542,N_570);
xnor U668 (N_668,N_503,N_583);
xnor U669 (N_669,N_506,N_536);
nand U670 (N_670,N_564,N_518);
nand U671 (N_671,N_539,N_546);
nor U672 (N_672,N_581,N_561);
or U673 (N_673,N_591,N_556);
and U674 (N_674,N_579,N_524);
nand U675 (N_675,N_593,N_515);
and U676 (N_676,N_529,N_574);
or U677 (N_677,N_537,N_508);
or U678 (N_678,N_532,N_529);
or U679 (N_679,N_582,N_510);
or U680 (N_680,N_560,N_557);
or U681 (N_681,N_533,N_547);
xnor U682 (N_682,N_569,N_508);
xnor U683 (N_683,N_566,N_561);
and U684 (N_684,N_573,N_538);
nor U685 (N_685,N_524,N_537);
and U686 (N_686,N_561,N_546);
xor U687 (N_687,N_562,N_533);
nor U688 (N_688,N_560,N_554);
and U689 (N_689,N_538,N_564);
nor U690 (N_690,N_571,N_538);
xnor U691 (N_691,N_524,N_501);
nand U692 (N_692,N_539,N_584);
and U693 (N_693,N_530,N_598);
nand U694 (N_694,N_556,N_520);
and U695 (N_695,N_525,N_581);
nand U696 (N_696,N_535,N_560);
nor U697 (N_697,N_546,N_592);
xor U698 (N_698,N_514,N_510);
xnor U699 (N_699,N_533,N_574);
xor U700 (N_700,N_649,N_621);
xor U701 (N_701,N_617,N_610);
and U702 (N_702,N_605,N_673);
nor U703 (N_703,N_644,N_660);
or U704 (N_704,N_634,N_630);
nor U705 (N_705,N_640,N_616);
and U706 (N_706,N_684,N_631);
and U707 (N_707,N_613,N_670);
and U708 (N_708,N_662,N_638);
xnor U709 (N_709,N_661,N_694);
xor U710 (N_710,N_622,N_609);
nor U711 (N_711,N_645,N_623);
xor U712 (N_712,N_606,N_632);
nor U713 (N_713,N_641,N_646);
and U714 (N_714,N_683,N_658);
or U715 (N_715,N_626,N_675);
nor U716 (N_716,N_691,N_671);
or U717 (N_717,N_627,N_656);
nand U718 (N_718,N_657,N_654);
and U719 (N_719,N_697,N_692);
or U720 (N_720,N_636,N_696);
or U721 (N_721,N_672,N_642);
and U722 (N_722,N_682,N_619);
or U723 (N_723,N_633,N_680);
nand U724 (N_724,N_659,N_625);
xnor U725 (N_725,N_615,N_674);
nor U726 (N_726,N_689,N_611);
nand U727 (N_727,N_686,N_655);
and U728 (N_728,N_665,N_679);
nor U729 (N_729,N_637,N_614);
and U730 (N_730,N_681,N_699);
nor U731 (N_731,N_647,N_629);
and U732 (N_732,N_678,N_667);
nand U733 (N_733,N_676,N_650);
or U734 (N_734,N_669,N_612);
nor U735 (N_735,N_695,N_601);
nand U736 (N_736,N_603,N_608);
nand U737 (N_737,N_607,N_653);
or U738 (N_738,N_648,N_624);
or U739 (N_739,N_666,N_668);
and U740 (N_740,N_602,N_690);
xor U741 (N_741,N_635,N_600);
and U742 (N_742,N_693,N_685);
or U743 (N_743,N_652,N_639);
and U744 (N_744,N_643,N_618);
or U745 (N_745,N_688,N_620);
nor U746 (N_746,N_604,N_663);
xor U747 (N_747,N_628,N_677);
xor U748 (N_748,N_664,N_687);
nor U749 (N_749,N_698,N_651);
nand U750 (N_750,N_655,N_636);
nor U751 (N_751,N_692,N_661);
and U752 (N_752,N_657,N_606);
or U753 (N_753,N_668,N_659);
nand U754 (N_754,N_624,N_629);
nand U755 (N_755,N_687,N_685);
xnor U756 (N_756,N_663,N_622);
and U757 (N_757,N_656,N_675);
xor U758 (N_758,N_614,N_629);
or U759 (N_759,N_642,N_619);
nor U760 (N_760,N_618,N_608);
or U761 (N_761,N_674,N_617);
xnor U762 (N_762,N_621,N_601);
xor U763 (N_763,N_604,N_674);
nor U764 (N_764,N_626,N_621);
nor U765 (N_765,N_656,N_618);
and U766 (N_766,N_679,N_626);
nand U767 (N_767,N_625,N_628);
xor U768 (N_768,N_677,N_662);
xor U769 (N_769,N_619,N_602);
nand U770 (N_770,N_639,N_664);
and U771 (N_771,N_631,N_677);
nor U772 (N_772,N_675,N_691);
xnor U773 (N_773,N_670,N_637);
and U774 (N_774,N_685,N_605);
or U775 (N_775,N_616,N_635);
nor U776 (N_776,N_604,N_672);
nor U777 (N_777,N_605,N_632);
nor U778 (N_778,N_633,N_609);
nand U779 (N_779,N_650,N_651);
or U780 (N_780,N_609,N_628);
or U781 (N_781,N_600,N_695);
and U782 (N_782,N_602,N_612);
xor U783 (N_783,N_617,N_623);
and U784 (N_784,N_627,N_638);
and U785 (N_785,N_661,N_677);
nor U786 (N_786,N_686,N_630);
nor U787 (N_787,N_672,N_654);
nor U788 (N_788,N_637,N_686);
and U789 (N_789,N_663,N_676);
xnor U790 (N_790,N_676,N_682);
or U791 (N_791,N_633,N_608);
or U792 (N_792,N_625,N_620);
nand U793 (N_793,N_686,N_610);
nor U794 (N_794,N_633,N_621);
or U795 (N_795,N_633,N_643);
and U796 (N_796,N_657,N_655);
xnor U797 (N_797,N_601,N_665);
nor U798 (N_798,N_656,N_685);
nor U799 (N_799,N_640,N_696);
nor U800 (N_800,N_772,N_782);
and U801 (N_801,N_785,N_784);
nor U802 (N_802,N_791,N_757);
or U803 (N_803,N_769,N_786);
nor U804 (N_804,N_755,N_723);
xnor U805 (N_805,N_798,N_708);
nor U806 (N_806,N_732,N_710);
and U807 (N_807,N_794,N_730);
xnor U808 (N_808,N_722,N_727);
or U809 (N_809,N_789,N_756);
and U810 (N_810,N_781,N_718);
or U811 (N_811,N_712,N_709);
nand U812 (N_812,N_795,N_790);
nand U813 (N_813,N_734,N_736);
xnor U814 (N_814,N_776,N_719);
xor U815 (N_815,N_753,N_768);
nand U816 (N_816,N_737,N_778);
nor U817 (N_817,N_751,N_773);
and U818 (N_818,N_735,N_780);
and U819 (N_819,N_766,N_725);
xnor U820 (N_820,N_783,N_740);
and U821 (N_821,N_752,N_716);
nor U822 (N_822,N_797,N_770);
and U823 (N_823,N_774,N_724);
nand U824 (N_824,N_771,N_777);
or U825 (N_825,N_704,N_706);
nor U826 (N_826,N_796,N_739);
nor U827 (N_827,N_763,N_779);
and U828 (N_828,N_720,N_749);
and U829 (N_829,N_711,N_715);
or U830 (N_830,N_787,N_703);
xor U831 (N_831,N_788,N_792);
or U832 (N_832,N_764,N_761);
or U833 (N_833,N_731,N_745);
nor U834 (N_834,N_741,N_750);
xor U835 (N_835,N_742,N_738);
xor U836 (N_836,N_714,N_746);
and U837 (N_837,N_700,N_743);
nor U838 (N_838,N_733,N_759);
nand U839 (N_839,N_748,N_702);
or U840 (N_840,N_762,N_701);
nor U841 (N_841,N_721,N_729);
xor U842 (N_842,N_767,N_758);
xor U843 (N_843,N_728,N_717);
or U844 (N_844,N_707,N_744);
or U845 (N_845,N_747,N_793);
or U846 (N_846,N_799,N_726);
xor U847 (N_847,N_775,N_754);
nand U848 (N_848,N_713,N_705);
or U849 (N_849,N_765,N_760);
or U850 (N_850,N_704,N_767);
nor U851 (N_851,N_763,N_781);
and U852 (N_852,N_709,N_795);
and U853 (N_853,N_720,N_783);
nor U854 (N_854,N_761,N_768);
xnor U855 (N_855,N_781,N_713);
and U856 (N_856,N_734,N_796);
nand U857 (N_857,N_729,N_776);
nand U858 (N_858,N_768,N_738);
and U859 (N_859,N_736,N_799);
nand U860 (N_860,N_721,N_712);
nor U861 (N_861,N_724,N_751);
nand U862 (N_862,N_712,N_785);
or U863 (N_863,N_756,N_791);
nand U864 (N_864,N_700,N_746);
and U865 (N_865,N_786,N_716);
or U866 (N_866,N_746,N_705);
and U867 (N_867,N_723,N_776);
xor U868 (N_868,N_704,N_797);
xnor U869 (N_869,N_781,N_774);
or U870 (N_870,N_735,N_726);
or U871 (N_871,N_786,N_719);
nand U872 (N_872,N_781,N_730);
xor U873 (N_873,N_774,N_710);
nor U874 (N_874,N_732,N_726);
and U875 (N_875,N_708,N_738);
nand U876 (N_876,N_776,N_701);
xor U877 (N_877,N_764,N_703);
xnor U878 (N_878,N_730,N_742);
xor U879 (N_879,N_790,N_706);
and U880 (N_880,N_715,N_726);
nor U881 (N_881,N_714,N_758);
and U882 (N_882,N_775,N_739);
or U883 (N_883,N_755,N_748);
or U884 (N_884,N_771,N_767);
or U885 (N_885,N_759,N_710);
xor U886 (N_886,N_790,N_737);
or U887 (N_887,N_703,N_757);
xor U888 (N_888,N_702,N_785);
xor U889 (N_889,N_785,N_744);
and U890 (N_890,N_785,N_797);
nand U891 (N_891,N_740,N_779);
nor U892 (N_892,N_781,N_741);
xor U893 (N_893,N_789,N_757);
or U894 (N_894,N_739,N_762);
and U895 (N_895,N_738,N_772);
or U896 (N_896,N_785,N_700);
xnor U897 (N_897,N_772,N_742);
and U898 (N_898,N_760,N_748);
nand U899 (N_899,N_735,N_755);
and U900 (N_900,N_839,N_803);
nand U901 (N_901,N_832,N_825);
xnor U902 (N_902,N_816,N_876);
or U903 (N_903,N_844,N_870);
or U904 (N_904,N_850,N_887);
xor U905 (N_905,N_800,N_805);
or U906 (N_906,N_829,N_827);
xor U907 (N_907,N_801,N_863);
nand U908 (N_908,N_820,N_828);
xnor U909 (N_909,N_809,N_858);
or U910 (N_910,N_866,N_834);
xor U911 (N_911,N_835,N_867);
nand U912 (N_912,N_895,N_852);
and U913 (N_913,N_881,N_879);
or U914 (N_914,N_822,N_886);
xnor U915 (N_915,N_859,N_896);
and U916 (N_916,N_812,N_890);
nor U917 (N_917,N_899,N_877);
nand U918 (N_918,N_885,N_855);
xor U919 (N_919,N_836,N_868);
or U920 (N_920,N_889,N_857);
and U921 (N_921,N_838,N_845);
nand U922 (N_922,N_874,N_891);
nand U923 (N_923,N_875,N_819);
nor U924 (N_924,N_888,N_861);
nand U925 (N_925,N_860,N_854);
or U926 (N_926,N_833,N_893);
nand U927 (N_927,N_830,N_808);
xnor U928 (N_928,N_862,N_848);
nand U929 (N_929,N_818,N_806);
nor U930 (N_930,N_873,N_837);
nor U931 (N_931,N_892,N_841);
nor U932 (N_932,N_807,N_856);
nor U933 (N_933,N_880,N_871);
and U934 (N_934,N_826,N_884);
nor U935 (N_935,N_824,N_865);
nor U936 (N_936,N_883,N_853);
nand U937 (N_937,N_882,N_823);
nand U938 (N_938,N_898,N_849);
or U939 (N_939,N_810,N_811);
and U940 (N_940,N_864,N_802);
and U941 (N_941,N_817,N_843);
and U942 (N_942,N_814,N_815);
and U943 (N_943,N_851,N_821);
or U944 (N_944,N_842,N_813);
nor U945 (N_945,N_878,N_804);
nor U946 (N_946,N_847,N_894);
xor U947 (N_947,N_872,N_846);
and U948 (N_948,N_831,N_840);
and U949 (N_949,N_897,N_869);
or U950 (N_950,N_851,N_891);
and U951 (N_951,N_883,N_848);
and U952 (N_952,N_834,N_874);
or U953 (N_953,N_861,N_880);
and U954 (N_954,N_832,N_843);
or U955 (N_955,N_854,N_826);
nand U956 (N_956,N_850,N_854);
nand U957 (N_957,N_850,N_800);
or U958 (N_958,N_816,N_818);
and U959 (N_959,N_853,N_888);
and U960 (N_960,N_882,N_803);
nor U961 (N_961,N_836,N_808);
nor U962 (N_962,N_865,N_820);
nand U963 (N_963,N_852,N_867);
xnor U964 (N_964,N_842,N_884);
or U965 (N_965,N_864,N_898);
xnor U966 (N_966,N_815,N_862);
nor U967 (N_967,N_866,N_896);
nor U968 (N_968,N_809,N_896);
or U969 (N_969,N_801,N_848);
and U970 (N_970,N_816,N_897);
xnor U971 (N_971,N_820,N_883);
xor U972 (N_972,N_874,N_863);
and U973 (N_973,N_831,N_810);
xnor U974 (N_974,N_876,N_891);
and U975 (N_975,N_872,N_870);
xnor U976 (N_976,N_824,N_869);
xor U977 (N_977,N_825,N_807);
nor U978 (N_978,N_876,N_890);
and U979 (N_979,N_834,N_836);
or U980 (N_980,N_821,N_888);
and U981 (N_981,N_856,N_874);
xnor U982 (N_982,N_838,N_825);
nand U983 (N_983,N_807,N_833);
or U984 (N_984,N_832,N_814);
nand U985 (N_985,N_811,N_857);
and U986 (N_986,N_839,N_816);
nand U987 (N_987,N_892,N_875);
and U988 (N_988,N_830,N_823);
nor U989 (N_989,N_875,N_834);
xor U990 (N_990,N_822,N_847);
and U991 (N_991,N_881,N_808);
nor U992 (N_992,N_806,N_837);
xor U993 (N_993,N_848,N_875);
nand U994 (N_994,N_814,N_844);
nor U995 (N_995,N_829,N_854);
and U996 (N_996,N_846,N_845);
and U997 (N_997,N_816,N_866);
xnor U998 (N_998,N_884,N_873);
nand U999 (N_999,N_865,N_846);
nor U1000 (N_1000,N_977,N_981);
nor U1001 (N_1001,N_935,N_909);
nand U1002 (N_1002,N_984,N_970);
xor U1003 (N_1003,N_913,N_933);
and U1004 (N_1004,N_945,N_903);
nand U1005 (N_1005,N_922,N_963);
nor U1006 (N_1006,N_941,N_901);
nor U1007 (N_1007,N_985,N_976);
nor U1008 (N_1008,N_926,N_919);
nor U1009 (N_1009,N_978,N_910);
or U1010 (N_1010,N_902,N_923);
xor U1011 (N_1011,N_906,N_967);
or U1012 (N_1012,N_940,N_959);
or U1013 (N_1013,N_988,N_912);
nor U1014 (N_1014,N_917,N_949);
xor U1015 (N_1015,N_980,N_952);
and U1016 (N_1016,N_937,N_921);
xor U1017 (N_1017,N_960,N_992);
nor U1018 (N_1018,N_918,N_974);
xor U1019 (N_1019,N_966,N_964);
and U1020 (N_1020,N_931,N_953);
and U1021 (N_1021,N_954,N_915);
nand U1022 (N_1022,N_911,N_928);
nor U1023 (N_1023,N_956,N_948);
xnor U1024 (N_1024,N_950,N_997);
or U1025 (N_1025,N_968,N_936);
nor U1026 (N_1026,N_932,N_955);
or U1027 (N_1027,N_993,N_999);
nand U1028 (N_1028,N_905,N_939);
and U1029 (N_1029,N_975,N_969);
nand U1030 (N_1030,N_965,N_942);
nand U1031 (N_1031,N_983,N_904);
nor U1032 (N_1032,N_947,N_900);
and U1033 (N_1033,N_938,N_962);
and U1034 (N_1034,N_957,N_925);
nor U1035 (N_1035,N_971,N_982);
nor U1036 (N_1036,N_946,N_987);
and U1037 (N_1037,N_979,N_929);
nand U1038 (N_1038,N_951,N_907);
or U1039 (N_1039,N_930,N_961);
or U1040 (N_1040,N_991,N_920);
or U1041 (N_1041,N_990,N_927);
nand U1042 (N_1042,N_944,N_924);
xnor U1043 (N_1043,N_994,N_958);
nand U1044 (N_1044,N_943,N_972);
nor U1045 (N_1045,N_973,N_989);
and U1046 (N_1046,N_916,N_995);
or U1047 (N_1047,N_914,N_908);
nand U1048 (N_1048,N_986,N_934);
nand U1049 (N_1049,N_996,N_998);
nand U1050 (N_1050,N_958,N_906);
and U1051 (N_1051,N_902,N_911);
or U1052 (N_1052,N_990,N_925);
or U1053 (N_1053,N_928,N_909);
xor U1054 (N_1054,N_930,N_957);
or U1055 (N_1055,N_930,N_902);
and U1056 (N_1056,N_983,N_939);
nor U1057 (N_1057,N_970,N_939);
and U1058 (N_1058,N_944,N_948);
xnor U1059 (N_1059,N_956,N_983);
nor U1060 (N_1060,N_991,N_947);
or U1061 (N_1061,N_921,N_999);
or U1062 (N_1062,N_917,N_903);
nand U1063 (N_1063,N_903,N_926);
and U1064 (N_1064,N_931,N_973);
nand U1065 (N_1065,N_924,N_982);
and U1066 (N_1066,N_939,N_989);
or U1067 (N_1067,N_931,N_916);
xor U1068 (N_1068,N_956,N_917);
and U1069 (N_1069,N_959,N_970);
xor U1070 (N_1070,N_939,N_979);
and U1071 (N_1071,N_918,N_958);
or U1072 (N_1072,N_989,N_960);
nand U1073 (N_1073,N_956,N_930);
nand U1074 (N_1074,N_907,N_954);
and U1075 (N_1075,N_932,N_977);
or U1076 (N_1076,N_936,N_933);
or U1077 (N_1077,N_941,N_925);
xor U1078 (N_1078,N_967,N_918);
nand U1079 (N_1079,N_980,N_985);
or U1080 (N_1080,N_914,N_974);
or U1081 (N_1081,N_904,N_993);
or U1082 (N_1082,N_985,N_917);
xor U1083 (N_1083,N_979,N_975);
nand U1084 (N_1084,N_980,N_958);
nor U1085 (N_1085,N_975,N_932);
nand U1086 (N_1086,N_929,N_992);
and U1087 (N_1087,N_969,N_982);
nor U1088 (N_1088,N_984,N_936);
nand U1089 (N_1089,N_968,N_957);
or U1090 (N_1090,N_964,N_960);
or U1091 (N_1091,N_974,N_950);
nor U1092 (N_1092,N_930,N_937);
xor U1093 (N_1093,N_920,N_925);
and U1094 (N_1094,N_950,N_999);
nand U1095 (N_1095,N_948,N_919);
nand U1096 (N_1096,N_940,N_941);
nand U1097 (N_1097,N_925,N_933);
nand U1098 (N_1098,N_905,N_945);
or U1099 (N_1099,N_979,N_909);
xor U1100 (N_1100,N_1014,N_1003);
or U1101 (N_1101,N_1036,N_1095);
nor U1102 (N_1102,N_1051,N_1034);
xnor U1103 (N_1103,N_1057,N_1011);
and U1104 (N_1104,N_1056,N_1087);
nand U1105 (N_1105,N_1020,N_1035);
or U1106 (N_1106,N_1059,N_1029);
nand U1107 (N_1107,N_1002,N_1065);
nor U1108 (N_1108,N_1008,N_1047);
or U1109 (N_1109,N_1061,N_1060);
and U1110 (N_1110,N_1090,N_1018);
or U1111 (N_1111,N_1009,N_1081);
xor U1112 (N_1112,N_1015,N_1092);
xnor U1113 (N_1113,N_1079,N_1041);
and U1114 (N_1114,N_1054,N_1075);
or U1115 (N_1115,N_1019,N_1044);
or U1116 (N_1116,N_1074,N_1052);
nand U1117 (N_1117,N_1048,N_1030);
and U1118 (N_1118,N_1082,N_1099);
xnor U1119 (N_1119,N_1032,N_1031);
and U1120 (N_1120,N_1023,N_1037);
nor U1121 (N_1121,N_1088,N_1049);
xor U1122 (N_1122,N_1022,N_1038);
and U1123 (N_1123,N_1089,N_1026);
xnor U1124 (N_1124,N_1062,N_1013);
nor U1125 (N_1125,N_1085,N_1042);
and U1126 (N_1126,N_1001,N_1093);
or U1127 (N_1127,N_1055,N_1078);
and U1128 (N_1128,N_1040,N_1004);
or U1129 (N_1129,N_1096,N_1094);
xnor U1130 (N_1130,N_1086,N_1000);
xor U1131 (N_1131,N_1025,N_1039);
xnor U1132 (N_1132,N_1097,N_1033);
nor U1133 (N_1133,N_1080,N_1064);
nor U1134 (N_1134,N_1006,N_1024);
nand U1135 (N_1135,N_1084,N_1058);
xnor U1136 (N_1136,N_1067,N_1070);
nor U1137 (N_1137,N_1010,N_1050);
and U1138 (N_1138,N_1083,N_1071);
nand U1139 (N_1139,N_1005,N_1027);
nand U1140 (N_1140,N_1098,N_1068);
nand U1141 (N_1141,N_1073,N_1053);
nor U1142 (N_1142,N_1046,N_1063);
xnor U1143 (N_1143,N_1043,N_1017);
nor U1144 (N_1144,N_1021,N_1028);
or U1145 (N_1145,N_1016,N_1091);
or U1146 (N_1146,N_1007,N_1069);
or U1147 (N_1147,N_1045,N_1077);
xnor U1148 (N_1148,N_1012,N_1076);
nand U1149 (N_1149,N_1072,N_1066);
nor U1150 (N_1150,N_1006,N_1098);
xor U1151 (N_1151,N_1048,N_1062);
xor U1152 (N_1152,N_1004,N_1095);
and U1153 (N_1153,N_1042,N_1077);
xnor U1154 (N_1154,N_1095,N_1023);
and U1155 (N_1155,N_1080,N_1089);
and U1156 (N_1156,N_1005,N_1067);
or U1157 (N_1157,N_1087,N_1005);
xor U1158 (N_1158,N_1068,N_1047);
xor U1159 (N_1159,N_1064,N_1095);
and U1160 (N_1160,N_1012,N_1061);
and U1161 (N_1161,N_1097,N_1070);
xnor U1162 (N_1162,N_1012,N_1072);
nand U1163 (N_1163,N_1094,N_1089);
or U1164 (N_1164,N_1069,N_1004);
xor U1165 (N_1165,N_1013,N_1086);
and U1166 (N_1166,N_1066,N_1011);
and U1167 (N_1167,N_1035,N_1093);
or U1168 (N_1168,N_1008,N_1062);
nand U1169 (N_1169,N_1052,N_1065);
and U1170 (N_1170,N_1093,N_1018);
xnor U1171 (N_1171,N_1068,N_1032);
or U1172 (N_1172,N_1030,N_1036);
or U1173 (N_1173,N_1020,N_1063);
xnor U1174 (N_1174,N_1055,N_1014);
xor U1175 (N_1175,N_1058,N_1015);
nor U1176 (N_1176,N_1065,N_1081);
and U1177 (N_1177,N_1035,N_1069);
and U1178 (N_1178,N_1025,N_1040);
xnor U1179 (N_1179,N_1037,N_1011);
and U1180 (N_1180,N_1081,N_1068);
and U1181 (N_1181,N_1074,N_1030);
and U1182 (N_1182,N_1065,N_1048);
nand U1183 (N_1183,N_1032,N_1057);
nor U1184 (N_1184,N_1058,N_1097);
nor U1185 (N_1185,N_1055,N_1031);
and U1186 (N_1186,N_1057,N_1065);
nor U1187 (N_1187,N_1013,N_1035);
and U1188 (N_1188,N_1043,N_1065);
and U1189 (N_1189,N_1090,N_1022);
or U1190 (N_1190,N_1082,N_1024);
nor U1191 (N_1191,N_1082,N_1076);
and U1192 (N_1192,N_1002,N_1070);
nand U1193 (N_1193,N_1090,N_1082);
xnor U1194 (N_1194,N_1055,N_1060);
nand U1195 (N_1195,N_1064,N_1024);
or U1196 (N_1196,N_1084,N_1037);
xnor U1197 (N_1197,N_1091,N_1074);
or U1198 (N_1198,N_1017,N_1021);
nor U1199 (N_1199,N_1000,N_1062);
or U1200 (N_1200,N_1153,N_1103);
xor U1201 (N_1201,N_1112,N_1132);
nor U1202 (N_1202,N_1136,N_1137);
xor U1203 (N_1203,N_1100,N_1186);
or U1204 (N_1204,N_1115,N_1162);
nand U1205 (N_1205,N_1128,N_1148);
and U1206 (N_1206,N_1196,N_1160);
and U1207 (N_1207,N_1130,N_1142);
nor U1208 (N_1208,N_1183,N_1182);
nand U1209 (N_1209,N_1113,N_1114);
and U1210 (N_1210,N_1116,N_1140);
nand U1211 (N_1211,N_1181,N_1191);
or U1212 (N_1212,N_1170,N_1133);
and U1213 (N_1213,N_1171,N_1194);
and U1214 (N_1214,N_1134,N_1144);
and U1215 (N_1215,N_1157,N_1105);
or U1216 (N_1216,N_1120,N_1131);
xor U1217 (N_1217,N_1168,N_1117);
and U1218 (N_1218,N_1159,N_1122);
xnor U1219 (N_1219,N_1192,N_1158);
and U1220 (N_1220,N_1107,N_1173);
nand U1221 (N_1221,N_1184,N_1138);
or U1222 (N_1222,N_1155,N_1172);
xnor U1223 (N_1223,N_1195,N_1106);
nand U1224 (N_1224,N_1164,N_1193);
nor U1225 (N_1225,N_1166,N_1176);
nor U1226 (N_1226,N_1188,N_1152);
nand U1227 (N_1227,N_1187,N_1161);
xnor U1228 (N_1228,N_1150,N_1108);
xor U1229 (N_1229,N_1141,N_1175);
nor U1230 (N_1230,N_1111,N_1154);
nor U1231 (N_1231,N_1199,N_1109);
nand U1232 (N_1232,N_1174,N_1198);
nand U1233 (N_1233,N_1151,N_1104);
nor U1234 (N_1234,N_1147,N_1126);
and U1235 (N_1235,N_1118,N_1125);
and U1236 (N_1236,N_1189,N_1139);
nor U1237 (N_1237,N_1167,N_1123);
nor U1238 (N_1238,N_1129,N_1190);
and U1239 (N_1239,N_1124,N_1180);
and U1240 (N_1240,N_1127,N_1102);
nand U1241 (N_1241,N_1121,N_1146);
or U1242 (N_1242,N_1179,N_1178);
nor U1243 (N_1243,N_1101,N_1169);
nor U1244 (N_1244,N_1156,N_1163);
xnor U1245 (N_1245,N_1145,N_1197);
and U1246 (N_1246,N_1185,N_1149);
and U1247 (N_1247,N_1110,N_1135);
nand U1248 (N_1248,N_1177,N_1165);
or U1249 (N_1249,N_1143,N_1119);
and U1250 (N_1250,N_1178,N_1166);
xnor U1251 (N_1251,N_1152,N_1172);
and U1252 (N_1252,N_1145,N_1130);
nor U1253 (N_1253,N_1119,N_1124);
and U1254 (N_1254,N_1179,N_1180);
and U1255 (N_1255,N_1192,N_1102);
or U1256 (N_1256,N_1116,N_1194);
nand U1257 (N_1257,N_1183,N_1159);
xnor U1258 (N_1258,N_1144,N_1141);
nor U1259 (N_1259,N_1179,N_1124);
nand U1260 (N_1260,N_1106,N_1193);
nor U1261 (N_1261,N_1106,N_1105);
or U1262 (N_1262,N_1170,N_1160);
xor U1263 (N_1263,N_1192,N_1199);
or U1264 (N_1264,N_1171,N_1187);
or U1265 (N_1265,N_1108,N_1158);
xnor U1266 (N_1266,N_1108,N_1114);
xnor U1267 (N_1267,N_1120,N_1103);
nand U1268 (N_1268,N_1106,N_1178);
nor U1269 (N_1269,N_1185,N_1157);
or U1270 (N_1270,N_1103,N_1167);
nand U1271 (N_1271,N_1123,N_1184);
nand U1272 (N_1272,N_1113,N_1120);
nor U1273 (N_1273,N_1146,N_1100);
and U1274 (N_1274,N_1132,N_1198);
nor U1275 (N_1275,N_1148,N_1157);
xor U1276 (N_1276,N_1161,N_1167);
nor U1277 (N_1277,N_1157,N_1159);
and U1278 (N_1278,N_1123,N_1197);
and U1279 (N_1279,N_1157,N_1173);
or U1280 (N_1280,N_1178,N_1165);
and U1281 (N_1281,N_1119,N_1184);
xnor U1282 (N_1282,N_1100,N_1106);
nand U1283 (N_1283,N_1124,N_1131);
or U1284 (N_1284,N_1108,N_1117);
and U1285 (N_1285,N_1125,N_1149);
or U1286 (N_1286,N_1168,N_1105);
xor U1287 (N_1287,N_1195,N_1124);
and U1288 (N_1288,N_1112,N_1104);
xor U1289 (N_1289,N_1171,N_1129);
or U1290 (N_1290,N_1170,N_1176);
nand U1291 (N_1291,N_1113,N_1140);
nand U1292 (N_1292,N_1152,N_1135);
or U1293 (N_1293,N_1164,N_1131);
and U1294 (N_1294,N_1161,N_1178);
or U1295 (N_1295,N_1103,N_1184);
nand U1296 (N_1296,N_1127,N_1123);
or U1297 (N_1297,N_1186,N_1129);
and U1298 (N_1298,N_1121,N_1161);
and U1299 (N_1299,N_1150,N_1193);
and U1300 (N_1300,N_1200,N_1287);
nor U1301 (N_1301,N_1201,N_1214);
or U1302 (N_1302,N_1245,N_1247);
or U1303 (N_1303,N_1221,N_1234);
and U1304 (N_1304,N_1225,N_1290);
or U1305 (N_1305,N_1226,N_1281);
nand U1306 (N_1306,N_1278,N_1264);
or U1307 (N_1307,N_1266,N_1277);
and U1308 (N_1308,N_1293,N_1212);
xnor U1309 (N_1309,N_1217,N_1242);
or U1310 (N_1310,N_1253,N_1294);
nor U1311 (N_1311,N_1205,N_1233);
xor U1312 (N_1312,N_1215,N_1283);
and U1313 (N_1313,N_1257,N_1260);
or U1314 (N_1314,N_1238,N_1298);
nand U1315 (N_1315,N_1286,N_1258);
nand U1316 (N_1316,N_1222,N_1259);
nand U1317 (N_1317,N_1244,N_1231);
nor U1318 (N_1318,N_1268,N_1219);
nand U1319 (N_1319,N_1273,N_1209);
xor U1320 (N_1320,N_1211,N_1241);
or U1321 (N_1321,N_1246,N_1292);
nor U1322 (N_1322,N_1295,N_1208);
and U1323 (N_1323,N_1288,N_1213);
xnor U1324 (N_1324,N_1236,N_1269);
xor U1325 (N_1325,N_1285,N_1249);
or U1326 (N_1326,N_1227,N_1250);
nand U1327 (N_1327,N_1252,N_1239);
nor U1328 (N_1328,N_1223,N_1203);
xnor U1329 (N_1329,N_1228,N_1240);
nand U1330 (N_1330,N_1271,N_1279);
xnor U1331 (N_1331,N_1262,N_1291);
and U1332 (N_1332,N_1220,N_1216);
xnor U1333 (N_1333,N_1263,N_1267);
and U1334 (N_1334,N_1272,N_1280);
or U1335 (N_1335,N_1251,N_1289);
xor U1336 (N_1336,N_1297,N_1235);
and U1337 (N_1337,N_1275,N_1230);
xor U1338 (N_1338,N_1254,N_1206);
nor U1339 (N_1339,N_1270,N_1237);
and U1340 (N_1340,N_1229,N_1232);
and U1341 (N_1341,N_1248,N_1282);
nor U1342 (N_1342,N_1261,N_1207);
and U1343 (N_1343,N_1284,N_1274);
and U1344 (N_1344,N_1276,N_1218);
or U1345 (N_1345,N_1256,N_1299);
or U1346 (N_1346,N_1224,N_1265);
nand U1347 (N_1347,N_1243,N_1202);
nor U1348 (N_1348,N_1255,N_1204);
and U1349 (N_1349,N_1210,N_1296);
nor U1350 (N_1350,N_1277,N_1285);
nand U1351 (N_1351,N_1217,N_1246);
and U1352 (N_1352,N_1269,N_1216);
xor U1353 (N_1353,N_1284,N_1261);
xnor U1354 (N_1354,N_1274,N_1228);
and U1355 (N_1355,N_1233,N_1209);
xor U1356 (N_1356,N_1266,N_1259);
xnor U1357 (N_1357,N_1217,N_1247);
and U1358 (N_1358,N_1227,N_1293);
and U1359 (N_1359,N_1275,N_1216);
and U1360 (N_1360,N_1244,N_1292);
nor U1361 (N_1361,N_1238,N_1232);
nand U1362 (N_1362,N_1209,N_1243);
xnor U1363 (N_1363,N_1275,N_1225);
xnor U1364 (N_1364,N_1270,N_1216);
nor U1365 (N_1365,N_1290,N_1287);
nand U1366 (N_1366,N_1231,N_1239);
nor U1367 (N_1367,N_1254,N_1293);
and U1368 (N_1368,N_1286,N_1261);
nor U1369 (N_1369,N_1201,N_1221);
nand U1370 (N_1370,N_1211,N_1242);
and U1371 (N_1371,N_1288,N_1266);
nand U1372 (N_1372,N_1246,N_1223);
or U1373 (N_1373,N_1211,N_1255);
and U1374 (N_1374,N_1230,N_1299);
or U1375 (N_1375,N_1256,N_1297);
or U1376 (N_1376,N_1231,N_1200);
xnor U1377 (N_1377,N_1203,N_1252);
and U1378 (N_1378,N_1228,N_1202);
or U1379 (N_1379,N_1234,N_1233);
nor U1380 (N_1380,N_1221,N_1292);
or U1381 (N_1381,N_1216,N_1279);
nor U1382 (N_1382,N_1274,N_1243);
and U1383 (N_1383,N_1244,N_1260);
nand U1384 (N_1384,N_1234,N_1215);
nor U1385 (N_1385,N_1269,N_1215);
nand U1386 (N_1386,N_1218,N_1290);
or U1387 (N_1387,N_1225,N_1293);
nand U1388 (N_1388,N_1237,N_1298);
or U1389 (N_1389,N_1247,N_1299);
nand U1390 (N_1390,N_1259,N_1297);
nor U1391 (N_1391,N_1289,N_1240);
and U1392 (N_1392,N_1212,N_1249);
and U1393 (N_1393,N_1242,N_1226);
xor U1394 (N_1394,N_1209,N_1295);
xor U1395 (N_1395,N_1268,N_1227);
xor U1396 (N_1396,N_1272,N_1210);
and U1397 (N_1397,N_1261,N_1263);
or U1398 (N_1398,N_1270,N_1279);
and U1399 (N_1399,N_1275,N_1243);
or U1400 (N_1400,N_1328,N_1362);
xor U1401 (N_1401,N_1386,N_1309);
and U1402 (N_1402,N_1383,N_1338);
or U1403 (N_1403,N_1391,N_1342);
and U1404 (N_1404,N_1381,N_1398);
nand U1405 (N_1405,N_1315,N_1316);
nor U1406 (N_1406,N_1301,N_1324);
and U1407 (N_1407,N_1339,N_1341);
nor U1408 (N_1408,N_1300,N_1311);
nand U1409 (N_1409,N_1390,N_1333);
and U1410 (N_1410,N_1363,N_1367);
or U1411 (N_1411,N_1394,N_1376);
xnor U1412 (N_1412,N_1352,N_1382);
or U1413 (N_1413,N_1335,N_1392);
or U1414 (N_1414,N_1380,N_1350);
xnor U1415 (N_1415,N_1320,N_1322);
or U1416 (N_1416,N_1357,N_1347);
and U1417 (N_1417,N_1374,N_1359);
or U1418 (N_1418,N_1340,N_1336);
and U1419 (N_1419,N_1317,N_1348);
or U1420 (N_1420,N_1389,N_1349);
and U1421 (N_1421,N_1393,N_1368);
nand U1422 (N_1422,N_1313,N_1303);
nand U1423 (N_1423,N_1318,N_1356);
or U1424 (N_1424,N_1369,N_1325);
nand U1425 (N_1425,N_1304,N_1344);
and U1426 (N_1426,N_1345,N_1378);
nand U1427 (N_1427,N_1365,N_1358);
and U1428 (N_1428,N_1307,N_1310);
nor U1429 (N_1429,N_1334,N_1314);
xnor U1430 (N_1430,N_1330,N_1351);
nor U1431 (N_1431,N_1355,N_1361);
or U1432 (N_1432,N_1327,N_1379);
xor U1433 (N_1433,N_1370,N_1331);
nor U1434 (N_1434,N_1396,N_1308);
nand U1435 (N_1435,N_1373,N_1353);
nor U1436 (N_1436,N_1360,N_1371);
nor U1437 (N_1437,N_1319,N_1377);
nor U1438 (N_1438,N_1364,N_1354);
and U1439 (N_1439,N_1302,N_1329);
or U1440 (N_1440,N_1343,N_1395);
or U1441 (N_1441,N_1337,N_1366);
or U1442 (N_1442,N_1384,N_1306);
nor U1443 (N_1443,N_1388,N_1375);
xnor U1444 (N_1444,N_1312,N_1326);
and U1445 (N_1445,N_1346,N_1397);
or U1446 (N_1446,N_1305,N_1387);
nor U1447 (N_1447,N_1372,N_1323);
nand U1448 (N_1448,N_1399,N_1385);
xor U1449 (N_1449,N_1332,N_1321);
nand U1450 (N_1450,N_1347,N_1348);
nor U1451 (N_1451,N_1386,N_1366);
or U1452 (N_1452,N_1301,N_1351);
and U1453 (N_1453,N_1356,N_1323);
xnor U1454 (N_1454,N_1344,N_1394);
nor U1455 (N_1455,N_1374,N_1332);
or U1456 (N_1456,N_1311,N_1347);
nand U1457 (N_1457,N_1360,N_1359);
nand U1458 (N_1458,N_1398,N_1393);
or U1459 (N_1459,N_1317,N_1360);
xnor U1460 (N_1460,N_1370,N_1313);
and U1461 (N_1461,N_1386,N_1385);
xnor U1462 (N_1462,N_1319,N_1383);
or U1463 (N_1463,N_1352,N_1348);
nor U1464 (N_1464,N_1373,N_1379);
nand U1465 (N_1465,N_1341,N_1399);
or U1466 (N_1466,N_1383,N_1362);
or U1467 (N_1467,N_1395,N_1389);
nor U1468 (N_1468,N_1380,N_1322);
and U1469 (N_1469,N_1309,N_1312);
nor U1470 (N_1470,N_1306,N_1328);
nor U1471 (N_1471,N_1374,N_1308);
nor U1472 (N_1472,N_1384,N_1386);
nand U1473 (N_1473,N_1313,N_1379);
nand U1474 (N_1474,N_1328,N_1347);
nand U1475 (N_1475,N_1310,N_1360);
and U1476 (N_1476,N_1384,N_1393);
nand U1477 (N_1477,N_1361,N_1390);
nor U1478 (N_1478,N_1367,N_1322);
or U1479 (N_1479,N_1317,N_1395);
xor U1480 (N_1480,N_1333,N_1325);
nor U1481 (N_1481,N_1302,N_1380);
nand U1482 (N_1482,N_1391,N_1338);
or U1483 (N_1483,N_1301,N_1308);
and U1484 (N_1484,N_1342,N_1308);
nand U1485 (N_1485,N_1398,N_1336);
and U1486 (N_1486,N_1337,N_1306);
nor U1487 (N_1487,N_1365,N_1317);
or U1488 (N_1488,N_1356,N_1378);
and U1489 (N_1489,N_1354,N_1318);
nand U1490 (N_1490,N_1338,N_1371);
and U1491 (N_1491,N_1379,N_1333);
nand U1492 (N_1492,N_1358,N_1324);
or U1493 (N_1493,N_1323,N_1367);
nor U1494 (N_1494,N_1353,N_1377);
or U1495 (N_1495,N_1325,N_1323);
and U1496 (N_1496,N_1389,N_1336);
or U1497 (N_1497,N_1349,N_1327);
nand U1498 (N_1498,N_1364,N_1308);
nand U1499 (N_1499,N_1354,N_1352);
xor U1500 (N_1500,N_1435,N_1452);
and U1501 (N_1501,N_1444,N_1430);
or U1502 (N_1502,N_1409,N_1406);
xor U1503 (N_1503,N_1499,N_1479);
or U1504 (N_1504,N_1410,N_1433);
nor U1505 (N_1505,N_1493,N_1462);
and U1506 (N_1506,N_1428,N_1456);
xnor U1507 (N_1507,N_1424,N_1466);
or U1508 (N_1508,N_1472,N_1415);
and U1509 (N_1509,N_1441,N_1443);
nand U1510 (N_1510,N_1455,N_1494);
or U1511 (N_1511,N_1483,N_1402);
nand U1512 (N_1512,N_1491,N_1457);
or U1513 (N_1513,N_1434,N_1445);
xor U1514 (N_1514,N_1438,N_1440);
xor U1515 (N_1515,N_1454,N_1416);
and U1516 (N_1516,N_1431,N_1403);
or U1517 (N_1517,N_1404,N_1484);
and U1518 (N_1518,N_1461,N_1463);
or U1519 (N_1519,N_1451,N_1471);
or U1520 (N_1520,N_1458,N_1478);
or U1521 (N_1521,N_1460,N_1486);
nand U1522 (N_1522,N_1498,N_1487);
or U1523 (N_1523,N_1436,N_1418);
and U1524 (N_1524,N_1467,N_1423);
or U1525 (N_1525,N_1449,N_1468);
nor U1526 (N_1526,N_1490,N_1422);
and U1527 (N_1527,N_1401,N_1442);
nor U1528 (N_1528,N_1495,N_1474);
nor U1529 (N_1529,N_1453,N_1480);
nand U1530 (N_1530,N_1405,N_1482);
nand U1531 (N_1531,N_1425,N_1476);
and U1532 (N_1532,N_1473,N_1496);
and U1533 (N_1533,N_1470,N_1448);
nand U1534 (N_1534,N_1432,N_1427);
nand U1535 (N_1535,N_1419,N_1488);
xnor U1536 (N_1536,N_1414,N_1408);
nor U1537 (N_1537,N_1417,N_1411);
nand U1538 (N_1538,N_1412,N_1420);
xor U1539 (N_1539,N_1413,N_1489);
nor U1540 (N_1540,N_1439,N_1492);
and U1541 (N_1541,N_1407,N_1450);
xnor U1542 (N_1542,N_1447,N_1464);
nand U1543 (N_1543,N_1429,N_1485);
nand U1544 (N_1544,N_1459,N_1400);
and U1545 (N_1545,N_1437,N_1421);
nor U1546 (N_1546,N_1465,N_1475);
and U1547 (N_1547,N_1477,N_1469);
xor U1548 (N_1548,N_1497,N_1481);
xor U1549 (N_1549,N_1446,N_1426);
xnor U1550 (N_1550,N_1487,N_1431);
xor U1551 (N_1551,N_1440,N_1416);
or U1552 (N_1552,N_1462,N_1418);
xor U1553 (N_1553,N_1457,N_1434);
and U1554 (N_1554,N_1441,N_1438);
and U1555 (N_1555,N_1483,N_1422);
or U1556 (N_1556,N_1449,N_1420);
or U1557 (N_1557,N_1475,N_1490);
nor U1558 (N_1558,N_1444,N_1452);
nand U1559 (N_1559,N_1483,N_1424);
xor U1560 (N_1560,N_1435,N_1489);
xor U1561 (N_1561,N_1400,N_1432);
or U1562 (N_1562,N_1464,N_1495);
nand U1563 (N_1563,N_1499,N_1431);
and U1564 (N_1564,N_1455,N_1450);
xnor U1565 (N_1565,N_1422,N_1456);
nor U1566 (N_1566,N_1460,N_1451);
and U1567 (N_1567,N_1479,N_1462);
and U1568 (N_1568,N_1447,N_1458);
or U1569 (N_1569,N_1487,N_1491);
and U1570 (N_1570,N_1480,N_1496);
xor U1571 (N_1571,N_1487,N_1407);
xnor U1572 (N_1572,N_1406,N_1481);
xor U1573 (N_1573,N_1403,N_1415);
and U1574 (N_1574,N_1428,N_1451);
nand U1575 (N_1575,N_1460,N_1438);
or U1576 (N_1576,N_1400,N_1475);
nand U1577 (N_1577,N_1496,N_1474);
or U1578 (N_1578,N_1473,N_1454);
and U1579 (N_1579,N_1444,N_1425);
xnor U1580 (N_1580,N_1432,N_1477);
xnor U1581 (N_1581,N_1473,N_1478);
nand U1582 (N_1582,N_1482,N_1454);
nand U1583 (N_1583,N_1411,N_1463);
and U1584 (N_1584,N_1492,N_1471);
or U1585 (N_1585,N_1430,N_1443);
xnor U1586 (N_1586,N_1404,N_1443);
or U1587 (N_1587,N_1492,N_1466);
and U1588 (N_1588,N_1475,N_1447);
nand U1589 (N_1589,N_1456,N_1442);
xnor U1590 (N_1590,N_1438,N_1404);
and U1591 (N_1591,N_1496,N_1457);
nand U1592 (N_1592,N_1418,N_1476);
or U1593 (N_1593,N_1467,N_1436);
nand U1594 (N_1594,N_1492,N_1488);
or U1595 (N_1595,N_1495,N_1440);
nand U1596 (N_1596,N_1410,N_1493);
xor U1597 (N_1597,N_1419,N_1499);
nand U1598 (N_1598,N_1411,N_1434);
nor U1599 (N_1599,N_1469,N_1450);
or U1600 (N_1600,N_1567,N_1524);
or U1601 (N_1601,N_1553,N_1506);
and U1602 (N_1602,N_1580,N_1508);
or U1603 (N_1603,N_1575,N_1531);
and U1604 (N_1604,N_1502,N_1535);
nor U1605 (N_1605,N_1544,N_1523);
and U1606 (N_1606,N_1505,N_1551);
xnor U1607 (N_1607,N_1533,N_1543);
nor U1608 (N_1608,N_1564,N_1563);
and U1609 (N_1609,N_1569,N_1530);
nor U1610 (N_1610,N_1512,N_1529);
xnor U1611 (N_1611,N_1582,N_1577);
nor U1612 (N_1612,N_1588,N_1566);
xor U1613 (N_1613,N_1542,N_1534);
xor U1614 (N_1614,N_1537,N_1519);
xor U1615 (N_1615,N_1558,N_1547);
or U1616 (N_1616,N_1546,N_1538);
xnor U1617 (N_1617,N_1503,N_1521);
nand U1618 (N_1618,N_1541,N_1510);
and U1619 (N_1619,N_1592,N_1554);
or U1620 (N_1620,N_1578,N_1526);
xnor U1621 (N_1621,N_1527,N_1555);
nor U1622 (N_1622,N_1504,N_1576);
or U1623 (N_1623,N_1573,N_1568);
and U1624 (N_1624,N_1539,N_1518);
xnor U1625 (N_1625,N_1548,N_1590);
and U1626 (N_1626,N_1532,N_1549);
nand U1627 (N_1627,N_1587,N_1517);
nand U1628 (N_1628,N_1507,N_1584);
nor U1629 (N_1629,N_1585,N_1599);
and U1630 (N_1630,N_1515,N_1594);
xnor U1631 (N_1631,N_1556,N_1562);
and U1632 (N_1632,N_1597,N_1528);
and U1633 (N_1633,N_1565,N_1525);
and U1634 (N_1634,N_1581,N_1579);
nand U1635 (N_1635,N_1596,N_1571);
xor U1636 (N_1636,N_1550,N_1591);
or U1637 (N_1637,N_1598,N_1561);
nand U1638 (N_1638,N_1545,N_1559);
or U1639 (N_1639,N_1593,N_1560);
or U1640 (N_1640,N_1511,N_1514);
and U1641 (N_1641,N_1501,N_1583);
or U1642 (N_1642,N_1509,N_1572);
and U1643 (N_1643,N_1595,N_1574);
nor U1644 (N_1644,N_1557,N_1522);
xor U1645 (N_1645,N_1520,N_1516);
or U1646 (N_1646,N_1500,N_1536);
and U1647 (N_1647,N_1589,N_1586);
and U1648 (N_1648,N_1570,N_1552);
and U1649 (N_1649,N_1513,N_1540);
and U1650 (N_1650,N_1560,N_1584);
or U1651 (N_1651,N_1521,N_1571);
or U1652 (N_1652,N_1535,N_1558);
or U1653 (N_1653,N_1520,N_1545);
nand U1654 (N_1654,N_1529,N_1573);
or U1655 (N_1655,N_1508,N_1592);
or U1656 (N_1656,N_1589,N_1560);
xor U1657 (N_1657,N_1510,N_1575);
nand U1658 (N_1658,N_1540,N_1568);
and U1659 (N_1659,N_1573,N_1547);
nand U1660 (N_1660,N_1556,N_1501);
or U1661 (N_1661,N_1560,N_1549);
nor U1662 (N_1662,N_1555,N_1517);
or U1663 (N_1663,N_1588,N_1510);
xor U1664 (N_1664,N_1598,N_1565);
nand U1665 (N_1665,N_1522,N_1515);
nor U1666 (N_1666,N_1578,N_1584);
xnor U1667 (N_1667,N_1516,N_1574);
or U1668 (N_1668,N_1590,N_1599);
nor U1669 (N_1669,N_1588,N_1584);
and U1670 (N_1670,N_1594,N_1554);
xnor U1671 (N_1671,N_1587,N_1589);
or U1672 (N_1672,N_1595,N_1590);
and U1673 (N_1673,N_1582,N_1574);
nand U1674 (N_1674,N_1535,N_1567);
and U1675 (N_1675,N_1521,N_1548);
nor U1676 (N_1676,N_1575,N_1513);
xor U1677 (N_1677,N_1559,N_1586);
or U1678 (N_1678,N_1582,N_1569);
xor U1679 (N_1679,N_1586,N_1571);
xor U1680 (N_1680,N_1598,N_1532);
and U1681 (N_1681,N_1577,N_1506);
xor U1682 (N_1682,N_1599,N_1539);
nor U1683 (N_1683,N_1545,N_1558);
nor U1684 (N_1684,N_1582,N_1545);
and U1685 (N_1685,N_1548,N_1574);
nand U1686 (N_1686,N_1501,N_1539);
and U1687 (N_1687,N_1502,N_1582);
and U1688 (N_1688,N_1505,N_1507);
nor U1689 (N_1689,N_1553,N_1596);
nand U1690 (N_1690,N_1505,N_1552);
or U1691 (N_1691,N_1550,N_1515);
and U1692 (N_1692,N_1518,N_1570);
nor U1693 (N_1693,N_1542,N_1566);
nand U1694 (N_1694,N_1531,N_1580);
xnor U1695 (N_1695,N_1552,N_1554);
and U1696 (N_1696,N_1562,N_1517);
and U1697 (N_1697,N_1563,N_1588);
nand U1698 (N_1698,N_1577,N_1536);
nand U1699 (N_1699,N_1538,N_1535);
or U1700 (N_1700,N_1683,N_1665);
or U1701 (N_1701,N_1649,N_1667);
nand U1702 (N_1702,N_1618,N_1691);
nor U1703 (N_1703,N_1600,N_1635);
xor U1704 (N_1704,N_1640,N_1620);
and U1705 (N_1705,N_1647,N_1673);
or U1706 (N_1706,N_1676,N_1668);
and U1707 (N_1707,N_1613,N_1682);
nand U1708 (N_1708,N_1650,N_1612);
nor U1709 (N_1709,N_1690,N_1608);
xor U1710 (N_1710,N_1664,N_1684);
and U1711 (N_1711,N_1697,N_1675);
nor U1712 (N_1712,N_1662,N_1645);
or U1713 (N_1713,N_1679,N_1621);
and U1714 (N_1714,N_1637,N_1652);
xnor U1715 (N_1715,N_1615,N_1656);
xor U1716 (N_1716,N_1678,N_1651);
and U1717 (N_1717,N_1619,N_1625);
nand U1718 (N_1718,N_1693,N_1669);
and U1719 (N_1719,N_1688,N_1602);
nor U1720 (N_1720,N_1674,N_1606);
xor U1721 (N_1721,N_1629,N_1692);
nand U1722 (N_1722,N_1666,N_1643);
nor U1723 (N_1723,N_1689,N_1699);
xor U1724 (N_1724,N_1617,N_1642);
nor U1725 (N_1725,N_1695,N_1610);
nand U1726 (N_1726,N_1671,N_1648);
and U1727 (N_1727,N_1630,N_1654);
xor U1728 (N_1728,N_1680,N_1604);
or U1729 (N_1729,N_1601,N_1623);
nand U1730 (N_1730,N_1698,N_1655);
nand U1731 (N_1731,N_1605,N_1603);
or U1732 (N_1732,N_1636,N_1644);
or U1733 (N_1733,N_1634,N_1614);
xnor U1734 (N_1734,N_1607,N_1687);
and U1735 (N_1735,N_1696,N_1631);
nand U1736 (N_1736,N_1632,N_1627);
nor U1737 (N_1737,N_1660,N_1670);
xor U1738 (N_1738,N_1685,N_1672);
nand U1739 (N_1739,N_1663,N_1653);
or U1740 (N_1740,N_1686,N_1624);
nand U1741 (N_1741,N_1646,N_1658);
xor U1742 (N_1742,N_1681,N_1611);
or U1743 (N_1743,N_1622,N_1639);
xnor U1744 (N_1744,N_1641,N_1633);
xor U1745 (N_1745,N_1657,N_1628);
or U1746 (N_1746,N_1638,N_1661);
and U1747 (N_1747,N_1626,N_1616);
xnor U1748 (N_1748,N_1609,N_1659);
nand U1749 (N_1749,N_1694,N_1677);
nand U1750 (N_1750,N_1691,N_1636);
or U1751 (N_1751,N_1654,N_1625);
or U1752 (N_1752,N_1693,N_1689);
and U1753 (N_1753,N_1619,N_1647);
or U1754 (N_1754,N_1677,N_1673);
and U1755 (N_1755,N_1677,N_1620);
or U1756 (N_1756,N_1629,N_1603);
nand U1757 (N_1757,N_1697,N_1665);
xnor U1758 (N_1758,N_1608,N_1686);
nor U1759 (N_1759,N_1626,N_1685);
nand U1760 (N_1760,N_1691,N_1656);
xor U1761 (N_1761,N_1681,N_1610);
xnor U1762 (N_1762,N_1636,N_1645);
nand U1763 (N_1763,N_1686,N_1640);
xor U1764 (N_1764,N_1604,N_1653);
or U1765 (N_1765,N_1628,N_1655);
nor U1766 (N_1766,N_1605,N_1671);
or U1767 (N_1767,N_1666,N_1640);
xnor U1768 (N_1768,N_1635,N_1621);
or U1769 (N_1769,N_1653,N_1640);
nor U1770 (N_1770,N_1651,N_1615);
xnor U1771 (N_1771,N_1627,N_1621);
and U1772 (N_1772,N_1619,N_1600);
and U1773 (N_1773,N_1673,N_1636);
nor U1774 (N_1774,N_1674,N_1672);
or U1775 (N_1775,N_1631,N_1651);
nand U1776 (N_1776,N_1647,N_1601);
and U1777 (N_1777,N_1629,N_1695);
or U1778 (N_1778,N_1647,N_1697);
nand U1779 (N_1779,N_1669,N_1643);
nand U1780 (N_1780,N_1624,N_1680);
nand U1781 (N_1781,N_1639,N_1659);
nor U1782 (N_1782,N_1690,N_1650);
and U1783 (N_1783,N_1687,N_1655);
or U1784 (N_1784,N_1697,N_1682);
nand U1785 (N_1785,N_1693,N_1635);
xnor U1786 (N_1786,N_1643,N_1659);
or U1787 (N_1787,N_1681,N_1661);
or U1788 (N_1788,N_1631,N_1694);
and U1789 (N_1789,N_1660,N_1607);
nor U1790 (N_1790,N_1665,N_1681);
nor U1791 (N_1791,N_1678,N_1623);
xnor U1792 (N_1792,N_1620,N_1630);
or U1793 (N_1793,N_1609,N_1639);
xor U1794 (N_1794,N_1672,N_1647);
nor U1795 (N_1795,N_1669,N_1679);
or U1796 (N_1796,N_1605,N_1618);
xnor U1797 (N_1797,N_1652,N_1661);
nand U1798 (N_1798,N_1699,N_1673);
nor U1799 (N_1799,N_1677,N_1646);
nand U1800 (N_1800,N_1742,N_1782);
nor U1801 (N_1801,N_1761,N_1713);
and U1802 (N_1802,N_1703,N_1741);
and U1803 (N_1803,N_1781,N_1785);
nor U1804 (N_1804,N_1734,N_1736);
nor U1805 (N_1805,N_1752,N_1774);
nor U1806 (N_1806,N_1706,N_1711);
nand U1807 (N_1807,N_1702,N_1733);
nand U1808 (N_1808,N_1796,N_1795);
nand U1809 (N_1809,N_1759,N_1794);
or U1810 (N_1810,N_1749,N_1788);
xnor U1811 (N_1811,N_1767,N_1727);
nor U1812 (N_1812,N_1790,N_1719);
and U1813 (N_1813,N_1776,N_1709);
nand U1814 (N_1814,N_1704,N_1760);
nand U1815 (N_1815,N_1770,N_1747);
nand U1816 (N_1816,N_1754,N_1739);
xnor U1817 (N_1817,N_1715,N_1777);
and U1818 (N_1818,N_1764,N_1769);
or U1819 (N_1819,N_1740,N_1707);
and U1820 (N_1820,N_1705,N_1700);
xnor U1821 (N_1821,N_1756,N_1793);
nand U1822 (N_1822,N_1780,N_1787);
xor U1823 (N_1823,N_1710,N_1768);
or U1824 (N_1824,N_1745,N_1744);
or U1825 (N_1825,N_1798,N_1714);
nor U1826 (N_1826,N_1786,N_1779);
or U1827 (N_1827,N_1724,N_1721);
xor U1828 (N_1828,N_1789,N_1737);
nand U1829 (N_1829,N_1775,N_1746);
nor U1830 (N_1830,N_1731,N_1757);
and U1831 (N_1831,N_1743,N_1791);
xor U1832 (N_1832,N_1751,N_1723);
or U1833 (N_1833,N_1797,N_1778);
nand U1834 (N_1834,N_1728,N_1753);
nand U1835 (N_1835,N_1718,N_1750);
nand U1836 (N_1836,N_1799,N_1716);
or U1837 (N_1837,N_1726,N_1792);
xnor U1838 (N_1838,N_1725,N_1773);
xnor U1839 (N_1839,N_1729,N_1755);
nand U1840 (N_1840,N_1772,N_1732);
and U1841 (N_1841,N_1763,N_1771);
or U1842 (N_1842,N_1784,N_1783);
or U1843 (N_1843,N_1762,N_1722);
nor U1844 (N_1844,N_1766,N_1758);
or U1845 (N_1845,N_1717,N_1748);
nand U1846 (N_1846,N_1735,N_1765);
nand U1847 (N_1847,N_1720,N_1712);
nor U1848 (N_1848,N_1708,N_1738);
nor U1849 (N_1849,N_1730,N_1701);
nand U1850 (N_1850,N_1799,N_1743);
and U1851 (N_1851,N_1781,N_1723);
or U1852 (N_1852,N_1793,N_1755);
xor U1853 (N_1853,N_1792,N_1769);
and U1854 (N_1854,N_1793,N_1780);
nor U1855 (N_1855,N_1713,N_1725);
nand U1856 (N_1856,N_1753,N_1721);
nor U1857 (N_1857,N_1707,N_1705);
nand U1858 (N_1858,N_1742,N_1716);
nor U1859 (N_1859,N_1713,N_1733);
nand U1860 (N_1860,N_1712,N_1751);
nand U1861 (N_1861,N_1765,N_1777);
and U1862 (N_1862,N_1770,N_1793);
or U1863 (N_1863,N_1726,N_1791);
and U1864 (N_1864,N_1794,N_1779);
nand U1865 (N_1865,N_1729,N_1766);
nand U1866 (N_1866,N_1705,N_1789);
and U1867 (N_1867,N_1768,N_1726);
nand U1868 (N_1868,N_1797,N_1709);
xor U1869 (N_1869,N_1713,N_1742);
xor U1870 (N_1870,N_1744,N_1758);
nor U1871 (N_1871,N_1753,N_1794);
xor U1872 (N_1872,N_1793,N_1726);
xnor U1873 (N_1873,N_1755,N_1726);
nand U1874 (N_1874,N_1712,N_1757);
or U1875 (N_1875,N_1781,N_1772);
or U1876 (N_1876,N_1790,N_1745);
nor U1877 (N_1877,N_1745,N_1763);
nor U1878 (N_1878,N_1712,N_1726);
or U1879 (N_1879,N_1749,N_1772);
and U1880 (N_1880,N_1761,N_1746);
xor U1881 (N_1881,N_1774,N_1734);
or U1882 (N_1882,N_1783,N_1712);
or U1883 (N_1883,N_1773,N_1788);
xor U1884 (N_1884,N_1714,N_1753);
nor U1885 (N_1885,N_1700,N_1733);
or U1886 (N_1886,N_1730,N_1729);
or U1887 (N_1887,N_1775,N_1709);
nand U1888 (N_1888,N_1729,N_1772);
or U1889 (N_1889,N_1724,N_1776);
xor U1890 (N_1890,N_1784,N_1744);
xor U1891 (N_1891,N_1739,N_1795);
and U1892 (N_1892,N_1716,N_1787);
nor U1893 (N_1893,N_1798,N_1736);
xor U1894 (N_1894,N_1731,N_1779);
nand U1895 (N_1895,N_1756,N_1795);
and U1896 (N_1896,N_1723,N_1797);
and U1897 (N_1897,N_1701,N_1773);
and U1898 (N_1898,N_1715,N_1737);
or U1899 (N_1899,N_1752,N_1731);
and U1900 (N_1900,N_1884,N_1886);
nand U1901 (N_1901,N_1842,N_1831);
nor U1902 (N_1902,N_1850,N_1881);
and U1903 (N_1903,N_1823,N_1876);
nand U1904 (N_1904,N_1851,N_1804);
xor U1905 (N_1905,N_1805,N_1813);
nand U1906 (N_1906,N_1858,N_1830);
nand U1907 (N_1907,N_1869,N_1807);
and U1908 (N_1908,N_1873,N_1892);
or U1909 (N_1909,N_1897,N_1847);
or U1910 (N_1910,N_1810,N_1874);
nand U1911 (N_1911,N_1814,N_1828);
or U1912 (N_1912,N_1853,N_1848);
nor U1913 (N_1913,N_1829,N_1809);
nand U1914 (N_1914,N_1885,N_1838);
xnor U1915 (N_1915,N_1890,N_1821);
xnor U1916 (N_1916,N_1877,N_1864);
and U1917 (N_1917,N_1812,N_1840);
xnor U1918 (N_1918,N_1887,N_1861);
xor U1919 (N_1919,N_1891,N_1862);
or U1920 (N_1920,N_1815,N_1803);
xor U1921 (N_1921,N_1837,N_1801);
nand U1922 (N_1922,N_1880,N_1820);
nor U1923 (N_1923,N_1836,N_1899);
and U1924 (N_1924,N_1802,N_1825);
nand U1925 (N_1925,N_1894,N_1819);
xnor U1926 (N_1926,N_1882,N_1875);
nor U1927 (N_1927,N_1868,N_1872);
and U1928 (N_1928,N_1816,N_1879);
and U1929 (N_1929,N_1883,N_1839);
and U1930 (N_1930,N_1835,N_1846);
nor U1931 (N_1931,N_1817,N_1855);
nand U1932 (N_1932,N_1843,N_1824);
and U1933 (N_1933,N_1800,N_1870);
xnor U1934 (N_1934,N_1806,N_1867);
xnor U1935 (N_1935,N_1849,N_1888);
or U1936 (N_1936,N_1827,N_1826);
xor U1937 (N_1937,N_1852,N_1863);
or U1938 (N_1938,N_1857,N_1856);
nand U1939 (N_1939,N_1893,N_1878);
xor U1940 (N_1940,N_1859,N_1808);
and U1941 (N_1941,N_1860,N_1865);
nor U1942 (N_1942,N_1889,N_1895);
nor U1943 (N_1943,N_1866,N_1818);
and U1944 (N_1944,N_1871,N_1832);
nand U1945 (N_1945,N_1834,N_1845);
and U1946 (N_1946,N_1811,N_1854);
xnor U1947 (N_1947,N_1844,N_1896);
xnor U1948 (N_1948,N_1822,N_1841);
xor U1949 (N_1949,N_1898,N_1833);
xnor U1950 (N_1950,N_1895,N_1887);
and U1951 (N_1951,N_1865,N_1895);
nor U1952 (N_1952,N_1863,N_1830);
nor U1953 (N_1953,N_1828,N_1869);
xor U1954 (N_1954,N_1880,N_1858);
and U1955 (N_1955,N_1856,N_1861);
xnor U1956 (N_1956,N_1893,N_1807);
nor U1957 (N_1957,N_1845,N_1859);
xnor U1958 (N_1958,N_1836,N_1824);
nand U1959 (N_1959,N_1814,N_1806);
and U1960 (N_1960,N_1867,N_1892);
and U1961 (N_1961,N_1805,N_1841);
nand U1962 (N_1962,N_1800,N_1877);
nor U1963 (N_1963,N_1891,N_1852);
nor U1964 (N_1964,N_1857,N_1818);
xnor U1965 (N_1965,N_1863,N_1871);
xor U1966 (N_1966,N_1833,N_1810);
xnor U1967 (N_1967,N_1867,N_1826);
nand U1968 (N_1968,N_1896,N_1853);
xor U1969 (N_1969,N_1877,N_1838);
xnor U1970 (N_1970,N_1875,N_1854);
and U1971 (N_1971,N_1894,N_1804);
nand U1972 (N_1972,N_1863,N_1809);
nor U1973 (N_1973,N_1815,N_1893);
nor U1974 (N_1974,N_1864,N_1814);
or U1975 (N_1975,N_1894,N_1812);
and U1976 (N_1976,N_1802,N_1897);
or U1977 (N_1977,N_1839,N_1866);
or U1978 (N_1978,N_1865,N_1804);
nor U1979 (N_1979,N_1860,N_1895);
nand U1980 (N_1980,N_1875,N_1842);
or U1981 (N_1981,N_1886,N_1854);
nor U1982 (N_1982,N_1890,N_1838);
nand U1983 (N_1983,N_1819,N_1827);
and U1984 (N_1984,N_1808,N_1827);
or U1985 (N_1985,N_1857,N_1806);
or U1986 (N_1986,N_1872,N_1860);
or U1987 (N_1987,N_1828,N_1810);
xnor U1988 (N_1988,N_1811,N_1838);
nand U1989 (N_1989,N_1806,N_1822);
and U1990 (N_1990,N_1835,N_1804);
or U1991 (N_1991,N_1856,N_1896);
or U1992 (N_1992,N_1840,N_1871);
xnor U1993 (N_1993,N_1882,N_1857);
nor U1994 (N_1994,N_1894,N_1862);
xor U1995 (N_1995,N_1889,N_1838);
nor U1996 (N_1996,N_1814,N_1843);
nand U1997 (N_1997,N_1877,N_1835);
nor U1998 (N_1998,N_1858,N_1810);
xnor U1999 (N_1999,N_1876,N_1840);
nor U2000 (N_2000,N_1945,N_1906);
or U2001 (N_2001,N_1930,N_1913);
xnor U2002 (N_2002,N_1905,N_1931);
nand U2003 (N_2003,N_1982,N_1940);
nor U2004 (N_2004,N_1944,N_1977);
nand U2005 (N_2005,N_1914,N_1968);
and U2006 (N_2006,N_1973,N_1919);
nor U2007 (N_2007,N_1989,N_1917);
and U2008 (N_2008,N_1958,N_1939);
and U2009 (N_2009,N_1986,N_1932);
and U2010 (N_2010,N_1963,N_1970);
xnor U2011 (N_2011,N_1996,N_1953);
nand U2012 (N_2012,N_1916,N_1947);
nand U2013 (N_2013,N_1964,N_1990);
xnor U2014 (N_2014,N_1926,N_1918);
xnor U2015 (N_2015,N_1983,N_1988);
nor U2016 (N_2016,N_1938,N_1995);
nor U2017 (N_2017,N_1998,N_1911);
xor U2018 (N_2018,N_1942,N_1959);
nand U2019 (N_2019,N_1987,N_1962);
xor U2020 (N_2020,N_1933,N_1927);
nand U2021 (N_2021,N_1925,N_1912);
nand U2022 (N_2022,N_1975,N_1915);
and U2023 (N_2023,N_1965,N_1967);
nor U2024 (N_2024,N_1941,N_1923);
nand U2025 (N_2025,N_1929,N_1900);
nor U2026 (N_2026,N_1937,N_1908);
or U2027 (N_2027,N_1984,N_1991);
xnor U2028 (N_2028,N_1985,N_1921);
nand U2029 (N_2029,N_1979,N_1935);
and U2030 (N_2030,N_1928,N_1960);
nand U2031 (N_2031,N_1981,N_1969);
xnor U2032 (N_2032,N_1978,N_1949);
xnor U2033 (N_2033,N_1934,N_1920);
nand U2034 (N_2034,N_1909,N_1961);
nor U2035 (N_2035,N_1936,N_1992);
nand U2036 (N_2036,N_1948,N_1904);
and U2037 (N_2037,N_1974,N_1902);
or U2038 (N_2038,N_1993,N_1954);
nand U2039 (N_2039,N_1957,N_1997);
xnor U2040 (N_2040,N_1971,N_1956);
xnor U2041 (N_2041,N_1976,N_1903);
and U2042 (N_2042,N_1950,N_1952);
and U2043 (N_2043,N_1943,N_1966);
nor U2044 (N_2044,N_1972,N_1924);
nor U2045 (N_2045,N_1946,N_1901);
xor U2046 (N_2046,N_1907,N_1922);
nand U2047 (N_2047,N_1999,N_1980);
or U2048 (N_2048,N_1951,N_1910);
xnor U2049 (N_2049,N_1955,N_1994);
nand U2050 (N_2050,N_1968,N_1907);
nor U2051 (N_2051,N_1902,N_1978);
xnor U2052 (N_2052,N_1954,N_1975);
or U2053 (N_2053,N_1929,N_1931);
and U2054 (N_2054,N_1986,N_1909);
and U2055 (N_2055,N_1971,N_1997);
and U2056 (N_2056,N_1963,N_1967);
nand U2057 (N_2057,N_1969,N_1907);
and U2058 (N_2058,N_1936,N_1954);
or U2059 (N_2059,N_1925,N_1961);
xor U2060 (N_2060,N_1928,N_1970);
xnor U2061 (N_2061,N_1998,N_1988);
nor U2062 (N_2062,N_1915,N_1929);
nor U2063 (N_2063,N_1951,N_1944);
or U2064 (N_2064,N_1986,N_1956);
or U2065 (N_2065,N_1905,N_1951);
and U2066 (N_2066,N_1930,N_1983);
and U2067 (N_2067,N_1915,N_1964);
xnor U2068 (N_2068,N_1928,N_1992);
nand U2069 (N_2069,N_1910,N_1967);
or U2070 (N_2070,N_1968,N_1954);
or U2071 (N_2071,N_1946,N_1980);
nor U2072 (N_2072,N_1994,N_1966);
or U2073 (N_2073,N_1924,N_1950);
nor U2074 (N_2074,N_1929,N_1902);
xnor U2075 (N_2075,N_1903,N_1925);
or U2076 (N_2076,N_1962,N_1917);
nor U2077 (N_2077,N_1971,N_1932);
or U2078 (N_2078,N_1929,N_1914);
nand U2079 (N_2079,N_1986,N_1980);
or U2080 (N_2080,N_1976,N_1935);
nor U2081 (N_2081,N_1987,N_1939);
or U2082 (N_2082,N_1963,N_1945);
and U2083 (N_2083,N_1938,N_1998);
nor U2084 (N_2084,N_1976,N_1978);
or U2085 (N_2085,N_1906,N_1999);
xor U2086 (N_2086,N_1943,N_1990);
xnor U2087 (N_2087,N_1961,N_1994);
or U2088 (N_2088,N_1912,N_1944);
and U2089 (N_2089,N_1967,N_1912);
nand U2090 (N_2090,N_1927,N_1907);
or U2091 (N_2091,N_1991,N_1969);
nand U2092 (N_2092,N_1933,N_1956);
nand U2093 (N_2093,N_1905,N_1935);
and U2094 (N_2094,N_1909,N_1956);
or U2095 (N_2095,N_1901,N_1909);
and U2096 (N_2096,N_1926,N_1959);
nor U2097 (N_2097,N_1913,N_1963);
xnor U2098 (N_2098,N_1969,N_1977);
nor U2099 (N_2099,N_1978,N_1991);
nand U2100 (N_2100,N_2028,N_2025);
or U2101 (N_2101,N_2056,N_2072);
and U2102 (N_2102,N_2086,N_2016);
and U2103 (N_2103,N_2023,N_2038);
and U2104 (N_2104,N_2009,N_2010);
xor U2105 (N_2105,N_2044,N_2014);
and U2106 (N_2106,N_2052,N_2068);
nor U2107 (N_2107,N_2047,N_2020);
nand U2108 (N_2108,N_2081,N_2031);
xnor U2109 (N_2109,N_2059,N_2034);
and U2110 (N_2110,N_2032,N_2045);
xnor U2111 (N_2111,N_2069,N_2035);
and U2112 (N_2112,N_2083,N_2004);
xnor U2113 (N_2113,N_2011,N_2079);
xor U2114 (N_2114,N_2097,N_2095);
and U2115 (N_2115,N_2062,N_2041);
nand U2116 (N_2116,N_2057,N_2061);
and U2117 (N_2117,N_2074,N_2087);
and U2118 (N_2118,N_2090,N_2021);
and U2119 (N_2119,N_2051,N_2029);
nor U2120 (N_2120,N_2024,N_2007);
or U2121 (N_2121,N_2048,N_2006);
and U2122 (N_2122,N_2065,N_2055);
and U2123 (N_2123,N_2037,N_2063);
or U2124 (N_2124,N_2026,N_2064);
nor U2125 (N_2125,N_2082,N_2098);
xor U2126 (N_2126,N_2066,N_2040);
xor U2127 (N_2127,N_2093,N_2085);
xnor U2128 (N_2128,N_2080,N_2049);
or U2129 (N_2129,N_2070,N_2027);
nand U2130 (N_2130,N_2099,N_2013);
nor U2131 (N_2131,N_2094,N_2077);
nand U2132 (N_2132,N_2067,N_2018);
nand U2133 (N_2133,N_2002,N_2092);
nor U2134 (N_2134,N_2053,N_2017);
or U2135 (N_2135,N_2050,N_2091);
nor U2136 (N_2136,N_2022,N_2012);
nor U2137 (N_2137,N_2042,N_2019);
or U2138 (N_2138,N_2039,N_2015);
nor U2139 (N_2139,N_2078,N_2043);
nor U2140 (N_2140,N_2036,N_2060);
nor U2141 (N_2141,N_2076,N_2075);
xnor U2142 (N_2142,N_2058,N_2046);
nand U2143 (N_2143,N_2084,N_2073);
or U2144 (N_2144,N_2008,N_2003);
and U2145 (N_2145,N_2088,N_2089);
nand U2146 (N_2146,N_2033,N_2005);
or U2147 (N_2147,N_2054,N_2030);
nor U2148 (N_2148,N_2001,N_2096);
xnor U2149 (N_2149,N_2000,N_2071);
nor U2150 (N_2150,N_2025,N_2059);
and U2151 (N_2151,N_2083,N_2092);
or U2152 (N_2152,N_2086,N_2068);
nor U2153 (N_2153,N_2020,N_2069);
or U2154 (N_2154,N_2027,N_2061);
nor U2155 (N_2155,N_2099,N_2057);
nand U2156 (N_2156,N_2016,N_2052);
nand U2157 (N_2157,N_2022,N_2003);
nand U2158 (N_2158,N_2025,N_2078);
xnor U2159 (N_2159,N_2085,N_2016);
nor U2160 (N_2160,N_2063,N_2020);
nor U2161 (N_2161,N_2013,N_2057);
nand U2162 (N_2162,N_2021,N_2024);
nor U2163 (N_2163,N_2095,N_2014);
or U2164 (N_2164,N_2081,N_2023);
nor U2165 (N_2165,N_2079,N_2056);
xnor U2166 (N_2166,N_2064,N_2030);
nand U2167 (N_2167,N_2035,N_2007);
and U2168 (N_2168,N_2092,N_2076);
or U2169 (N_2169,N_2012,N_2062);
xor U2170 (N_2170,N_2010,N_2064);
xnor U2171 (N_2171,N_2018,N_2019);
and U2172 (N_2172,N_2085,N_2010);
and U2173 (N_2173,N_2093,N_2089);
nand U2174 (N_2174,N_2062,N_2087);
or U2175 (N_2175,N_2067,N_2083);
or U2176 (N_2176,N_2039,N_2017);
nor U2177 (N_2177,N_2066,N_2075);
nand U2178 (N_2178,N_2079,N_2038);
nand U2179 (N_2179,N_2064,N_2051);
or U2180 (N_2180,N_2083,N_2056);
nor U2181 (N_2181,N_2081,N_2048);
or U2182 (N_2182,N_2095,N_2036);
xor U2183 (N_2183,N_2041,N_2051);
nor U2184 (N_2184,N_2050,N_2096);
xnor U2185 (N_2185,N_2077,N_2040);
nor U2186 (N_2186,N_2027,N_2022);
or U2187 (N_2187,N_2003,N_2028);
and U2188 (N_2188,N_2025,N_2058);
and U2189 (N_2189,N_2082,N_2016);
nand U2190 (N_2190,N_2065,N_2082);
nand U2191 (N_2191,N_2021,N_2081);
or U2192 (N_2192,N_2003,N_2097);
or U2193 (N_2193,N_2022,N_2089);
xor U2194 (N_2194,N_2069,N_2055);
nor U2195 (N_2195,N_2081,N_2094);
and U2196 (N_2196,N_2082,N_2002);
and U2197 (N_2197,N_2023,N_2063);
xor U2198 (N_2198,N_2006,N_2011);
or U2199 (N_2199,N_2042,N_2003);
nand U2200 (N_2200,N_2130,N_2194);
xor U2201 (N_2201,N_2122,N_2172);
or U2202 (N_2202,N_2109,N_2140);
xor U2203 (N_2203,N_2138,N_2123);
xnor U2204 (N_2204,N_2110,N_2115);
xor U2205 (N_2205,N_2136,N_2189);
nor U2206 (N_2206,N_2195,N_2184);
nand U2207 (N_2207,N_2191,N_2182);
and U2208 (N_2208,N_2160,N_2173);
nand U2209 (N_2209,N_2164,N_2170);
nand U2210 (N_2210,N_2114,N_2102);
and U2211 (N_2211,N_2101,N_2174);
nand U2212 (N_2212,N_2193,N_2100);
nand U2213 (N_2213,N_2186,N_2199);
and U2214 (N_2214,N_2176,N_2121);
nand U2215 (N_2215,N_2139,N_2132);
nor U2216 (N_2216,N_2108,N_2188);
xor U2217 (N_2217,N_2190,N_2157);
nand U2218 (N_2218,N_2158,N_2152);
and U2219 (N_2219,N_2116,N_2180);
nor U2220 (N_2220,N_2196,N_2149);
nand U2221 (N_2221,N_2126,N_2104);
xor U2222 (N_2222,N_2141,N_2133);
and U2223 (N_2223,N_2197,N_2181);
and U2224 (N_2224,N_2150,N_2178);
or U2225 (N_2225,N_2143,N_2168);
nand U2226 (N_2226,N_2120,N_2144);
or U2227 (N_2227,N_2145,N_2107);
or U2228 (N_2228,N_2118,N_2142);
xor U2229 (N_2229,N_2198,N_2135);
nand U2230 (N_2230,N_2111,N_2147);
xnor U2231 (N_2231,N_2159,N_2131);
nand U2232 (N_2232,N_2187,N_2156);
nor U2233 (N_2233,N_2154,N_2185);
xnor U2234 (N_2234,N_2192,N_2148);
or U2235 (N_2235,N_2166,N_2125);
nor U2236 (N_2236,N_2153,N_2124);
nand U2237 (N_2237,N_2119,N_2103);
or U2238 (N_2238,N_2177,N_2162);
nand U2239 (N_2239,N_2167,N_2183);
xor U2240 (N_2240,N_2127,N_2171);
nor U2241 (N_2241,N_2117,N_2128);
or U2242 (N_2242,N_2113,N_2163);
nor U2243 (N_2243,N_2155,N_2161);
nand U2244 (N_2244,N_2112,N_2137);
or U2245 (N_2245,N_2105,N_2129);
and U2246 (N_2246,N_2165,N_2175);
or U2247 (N_2247,N_2169,N_2179);
nand U2248 (N_2248,N_2106,N_2151);
nor U2249 (N_2249,N_2134,N_2146);
xnor U2250 (N_2250,N_2176,N_2132);
nor U2251 (N_2251,N_2188,N_2152);
or U2252 (N_2252,N_2196,N_2185);
nor U2253 (N_2253,N_2176,N_2182);
nor U2254 (N_2254,N_2154,N_2147);
and U2255 (N_2255,N_2124,N_2155);
nand U2256 (N_2256,N_2135,N_2192);
nand U2257 (N_2257,N_2118,N_2112);
or U2258 (N_2258,N_2101,N_2106);
and U2259 (N_2259,N_2138,N_2132);
and U2260 (N_2260,N_2116,N_2133);
or U2261 (N_2261,N_2138,N_2164);
or U2262 (N_2262,N_2152,N_2124);
nand U2263 (N_2263,N_2123,N_2195);
and U2264 (N_2264,N_2143,N_2122);
or U2265 (N_2265,N_2198,N_2151);
xor U2266 (N_2266,N_2192,N_2165);
nor U2267 (N_2267,N_2191,N_2138);
or U2268 (N_2268,N_2153,N_2196);
and U2269 (N_2269,N_2104,N_2109);
xnor U2270 (N_2270,N_2159,N_2161);
nand U2271 (N_2271,N_2186,N_2106);
nor U2272 (N_2272,N_2106,N_2138);
nand U2273 (N_2273,N_2139,N_2161);
xor U2274 (N_2274,N_2145,N_2148);
xor U2275 (N_2275,N_2142,N_2185);
and U2276 (N_2276,N_2185,N_2180);
or U2277 (N_2277,N_2142,N_2198);
nor U2278 (N_2278,N_2116,N_2153);
xor U2279 (N_2279,N_2142,N_2191);
nand U2280 (N_2280,N_2179,N_2190);
or U2281 (N_2281,N_2158,N_2154);
or U2282 (N_2282,N_2197,N_2133);
or U2283 (N_2283,N_2173,N_2164);
xnor U2284 (N_2284,N_2160,N_2132);
nor U2285 (N_2285,N_2164,N_2141);
nor U2286 (N_2286,N_2164,N_2199);
xor U2287 (N_2287,N_2130,N_2142);
nand U2288 (N_2288,N_2139,N_2146);
xor U2289 (N_2289,N_2154,N_2181);
nand U2290 (N_2290,N_2149,N_2162);
or U2291 (N_2291,N_2111,N_2117);
or U2292 (N_2292,N_2109,N_2120);
nand U2293 (N_2293,N_2127,N_2164);
nand U2294 (N_2294,N_2115,N_2111);
nor U2295 (N_2295,N_2177,N_2107);
xnor U2296 (N_2296,N_2191,N_2161);
xnor U2297 (N_2297,N_2185,N_2144);
nand U2298 (N_2298,N_2135,N_2109);
or U2299 (N_2299,N_2168,N_2131);
and U2300 (N_2300,N_2213,N_2278);
nand U2301 (N_2301,N_2259,N_2264);
or U2302 (N_2302,N_2260,N_2261);
nand U2303 (N_2303,N_2232,N_2291);
xor U2304 (N_2304,N_2252,N_2263);
nor U2305 (N_2305,N_2254,N_2237);
nand U2306 (N_2306,N_2242,N_2257);
and U2307 (N_2307,N_2274,N_2285);
nor U2308 (N_2308,N_2282,N_2297);
nor U2309 (N_2309,N_2265,N_2211);
nor U2310 (N_2310,N_2299,N_2202);
or U2311 (N_2311,N_2223,N_2272);
nand U2312 (N_2312,N_2294,N_2248);
or U2313 (N_2313,N_2286,N_2296);
nand U2314 (N_2314,N_2218,N_2224);
and U2315 (N_2315,N_2210,N_2239);
nor U2316 (N_2316,N_2243,N_2229);
nand U2317 (N_2317,N_2258,N_2233);
nor U2318 (N_2318,N_2219,N_2228);
and U2319 (N_2319,N_2268,N_2236);
and U2320 (N_2320,N_2217,N_2251);
nand U2321 (N_2321,N_2276,N_2283);
or U2322 (N_2322,N_2203,N_2214);
nand U2323 (N_2323,N_2284,N_2256);
nand U2324 (N_2324,N_2275,N_2281);
and U2325 (N_2325,N_2206,N_2288);
nand U2326 (N_2326,N_2200,N_2244);
nand U2327 (N_2327,N_2280,N_2250);
nor U2328 (N_2328,N_2212,N_2235);
nor U2329 (N_2329,N_2295,N_2289);
nand U2330 (N_2330,N_2225,N_2222);
or U2331 (N_2331,N_2207,N_2273);
nor U2332 (N_2332,N_2241,N_2287);
and U2333 (N_2333,N_2208,N_2201);
xnor U2334 (N_2334,N_2215,N_2220);
or U2335 (N_2335,N_2279,N_2292);
nor U2336 (N_2336,N_2209,N_2277);
xor U2337 (N_2337,N_2221,N_2262);
or U2338 (N_2338,N_2234,N_2216);
or U2339 (N_2339,N_2290,N_2293);
xnor U2340 (N_2340,N_2298,N_2231);
nor U2341 (N_2341,N_2247,N_2266);
xnor U2342 (N_2342,N_2230,N_2226);
xor U2343 (N_2343,N_2246,N_2240);
nor U2344 (N_2344,N_2245,N_2227);
nand U2345 (N_2345,N_2253,N_2270);
or U2346 (N_2346,N_2255,N_2205);
or U2347 (N_2347,N_2271,N_2269);
nand U2348 (N_2348,N_2204,N_2249);
nand U2349 (N_2349,N_2238,N_2267);
nand U2350 (N_2350,N_2201,N_2287);
nand U2351 (N_2351,N_2286,N_2294);
xor U2352 (N_2352,N_2233,N_2224);
xor U2353 (N_2353,N_2285,N_2240);
and U2354 (N_2354,N_2244,N_2214);
and U2355 (N_2355,N_2271,N_2200);
or U2356 (N_2356,N_2250,N_2273);
or U2357 (N_2357,N_2204,N_2275);
xor U2358 (N_2358,N_2232,N_2226);
or U2359 (N_2359,N_2230,N_2202);
nand U2360 (N_2360,N_2227,N_2286);
and U2361 (N_2361,N_2227,N_2222);
or U2362 (N_2362,N_2223,N_2262);
nor U2363 (N_2363,N_2267,N_2243);
nor U2364 (N_2364,N_2230,N_2275);
nor U2365 (N_2365,N_2243,N_2265);
nor U2366 (N_2366,N_2205,N_2297);
nor U2367 (N_2367,N_2241,N_2248);
or U2368 (N_2368,N_2202,N_2204);
xor U2369 (N_2369,N_2219,N_2200);
and U2370 (N_2370,N_2218,N_2209);
nand U2371 (N_2371,N_2241,N_2221);
nand U2372 (N_2372,N_2213,N_2253);
xnor U2373 (N_2373,N_2256,N_2228);
nand U2374 (N_2374,N_2226,N_2209);
nand U2375 (N_2375,N_2284,N_2223);
nor U2376 (N_2376,N_2214,N_2236);
nor U2377 (N_2377,N_2278,N_2237);
and U2378 (N_2378,N_2265,N_2287);
xnor U2379 (N_2379,N_2257,N_2240);
or U2380 (N_2380,N_2287,N_2259);
or U2381 (N_2381,N_2271,N_2265);
xor U2382 (N_2382,N_2267,N_2232);
and U2383 (N_2383,N_2265,N_2299);
nor U2384 (N_2384,N_2287,N_2273);
and U2385 (N_2385,N_2215,N_2279);
and U2386 (N_2386,N_2220,N_2240);
xor U2387 (N_2387,N_2214,N_2294);
nand U2388 (N_2388,N_2204,N_2258);
and U2389 (N_2389,N_2296,N_2218);
and U2390 (N_2390,N_2263,N_2243);
xnor U2391 (N_2391,N_2294,N_2260);
or U2392 (N_2392,N_2288,N_2243);
and U2393 (N_2393,N_2273,N_2202);
nor U2394 (N_2394,N_2280,N_2235);
nand U2395 (N_2395,N_2264,N_2205);
nand U2396 (N_2396,N_2268,N_2212);
nand U2397 (N_2397,N_2217,N_2286);
xnor U2398 (N_2398,N_2250,N_2240);
xor U2399 (N_2399,N_2205,N_2224);
xor U2400 (N_2400,N_2341,N_2316);
and U2401 (N_2401,N_2315,N_2338);
and U2402 (N_2402,N_2302,N_2384);
nor U2403 (N_2403,N_2343,N_2358);
nor U2404 (N_2404,N_2367,N_2339);
nand U2405 (N_2405,N_2371,N_2331);
nor U2406 (N_2406,N_2327,N_2373);
xor U2407 (N_2407,N_2354,N_2310);
xor U2408 (N_2408,N_2381,N_2333);
nand U2409 (N_2409,N_2318,N_2389);
nor U2410 (N_2410,N_2393,N_2363);
and U2411 (N_2411,N_2306,N_2323);
nor U2412 (N_2412,N_2382,N_2347);
nor U2413 (N_2413,N_2396,N_2311);
xnor U2414 (N_2414,N_2394,N_2355);
nor U2415 (N_2415,N_2377,N_2391);
nand U2416 (N_2416,N_2380,N_2345);
nand U2417 (N_2417,N_2376,N_2397);
or U2418 (N_2418,N_2390,N_2360);
nor U2419 (N_2419,N_2340,N_2342);
or U2420 (N_2420,N_2330,N_2308);
and U2421 (N_2421,N_2320,N_2353);
nand U2422 (N_2422,N_2326,N_2319);
nand U2423 (N_2423,N_2399,N_2303);
nor U2424 (N_2424,N_2361,N_2300);
xnor U2425 (N_2425,N_2301,N_2350);
nor U2426 (N_2426,N_2309,N_2313);
nand U2427 (N_2427,N_2392,N_2304);
nor U2428 (N_2428,N_2362,N_2337);
xor U2429 (N_2429,N_2357,N_2366);
nand U2430 (N_2430,N_2379,N_2372);
or U2431 (N_2431,N_2374,N_2349);
nand U2432 (N_2432,N_2324,N_2352);
or U2433 (N_2433,N_2348,N_2321);
xnor U2434 (N_2434,N_2346,N_2344);
and U2435 (N_2435,N_2378,N_2314);
or U2436 (N_2436,N_2369,N_2351);
nand U2437 (N_2437,N_2387,N_2312);
and U2438 (N_2438,N_2305,N_2335);
and U2439 (N_2439,N_2329,N_2336);
xnor U2440 (N_2440,N_2359,N_2317);
or U2441 (N_2441,N_2398,N_2375);
nand U2442 (N_2442,N_2386,N_2325);
nor U2443 (N_2443,N_2364,N_2328);
and U2444 (N_2444,N_2368,N_2356);
xor U2445 (N_2445,N_2307,N_2388);
or U2446 (N_2446,N_2383,N_2385);
nor U2447 (N_2447,N_2370,N_2395);
nand U2448 (N_2448,N_2322,N_2334);
nand U2449 (N_2449,N_2365,N_2332);
nand U2450 (N_2450,N_2325,N_2364);
or U2451 (N_2451,N_2325,N_2352);
or U2452 (N_2452,N_2322,N_2301);
xor U2453 (N_2453,N_2397,N_2320);
xor U2454 (N_2454,N_2322,N_2394);
nand U2455 (N_2455,N_2386,N_2306);
nand U2456 (N_2456,N_2339,N_2341);
and U2457 (N_2457,N_2368,N_2390);
and U2458 (N_2458,N_2360,N_2330);
or U2459 (N_2459,N_2350,N_2326);
or U2460 (N_2460,N_2373,N_2372);
nand U2461 (N_2461,N_2345,N_2325);
nor U2462 (N_2462,N_2353,N_2340);
and U2463 (N_2463,N_2313,N_2303);
xnor U2464 (N_2464,N_2372,N_2389);
or U2465 (N_2465,N_2383,N_2307);
and U2466 (N_2466,N_2347,N_2368);
xor U2467 (N_2467,N_2347,N_2397);
nor U2468 (N_2468,N_2305,N_2351);
or U2469 (N_2469,N_2367,N_2379);
xor U2470 (N_2470,N_2301,N_2329);
and U2471 (N_2471,N_2313,N_2323);
nand U2472 (N_2472,N_2328,N_2335);
nand U2473 (N_2473,N_2339,N_2385);
and U2474 (N_2474,N_2347,N_2307);
nor U2475 (N_2475,N_2316,N_2349);
nor U2476 (N_2476,N_2316,N_2356);
and U2477 (N_2477,N_2357,N_2316);
and U2478 (N_2478,N_2355,N_2388);
and U2479 (N_2479,N_2308,N_2313);
and U2480 (N_2480,N_2395,N_2399);
nor U2481 (N_2481,N_2396,N_2303);
xnor U2482 (N_2482,N_2395,N_2320);
or U2483 (N_2483,N_2376,N_2304);
nand U2484 (N_2484,N_2319,N_2322);
and U2485 (N_2485,N_2375,N_2326);
nor U2486 (N_2486,N_2357,N_2395);
nor U2487 (N_2487,N_2385,N_2310);
and U2488 (N_2488,N_2375,N_2376);
and U2489 (N_2489,N_2358,N_2378);
xor U2490 (N_2490,N_2303,N_2354);
and U2491 (N_2491,N_2316,N_2365);
nand U2492 (N_2492,N_2318,N_2381);
xnor U2493 (N_2493,N_2346,N_2375);
nor U2494 (N_2494,N_2312,N_2386);
or U2495 (N_2495,N_2373,N_2336);
nand U2496 (N_2496,N_2368,N_2363);
or U2497 (N_2497,N_2331,N_2309);
xnor U2498 (N_2498,N_2340,N_2341);
xor U2499 (N_2499,N_2382,N_2330);
xor U2500 (N_2500,N_2458,N_2441);
nor U2501 (N_2501,N_2421,N_2461);
and U2502 (N_2502,N_2487,N_2425);
nor U2503 (N_2503,N_2406,N_2435);
nand U2504 (N_2504,N_2477,N_2478);
xor U2505 (N_2505,N_2426,N_2463);
xnor U2506 (N_2506,N_2405,N_2430);
xor U2507 (N_2507,N_2448,N_2459);
nor U2508 (N_2508,N_2403,N_2431);
nand U2509 (N_2509,N_2470,N_2480);
or U2510 (N_2510,N_2409,N_2447);
or U2511 (N_2511,N_2494,N_2422);
nor U2512 (N_2512,N_2466,N_2473);
and U2513 (N_2513,N_2420,N_2481);
and U2514 (N_2514,N_2439,N_2412);
nand U2515 (N_2515,N_2476,N_2407);
and U2516 (N_2516,N_2451,N_2492);
nand U2517 (N_2517,N_2450,N_2429);
or U2518 (N_2518,N_2482,N_2468);
nor U2519 (N_2519,N_2428,N_2497);
and U2520 (N_2520,N_2456,N_2498);
nor U2521 (N_2521,N_2442,N_2491);
xor U2522 (N_2522,N_2415,N_2427);
and U2523 (N_2523,N_2460,N_2438);
or U2524 (N_2524,N_2417,N_2453);
or U2525 (N_2525,N_2404,N_2436);
nor U2526 (N_2526,N_2410,N_2474);
nand U2527 (N_2527,N_2433,N_2479);
nor U2528 (N_2528,N_2484,N_2490);
or U2529 (N_2529,N_2464,N_2444);
nand U2530 (N_2530,N_2452,N_2414);
xor U2531 (N_2531,N_2402,N_2423);
nor U2532 (N_2532,N_2418,N_2471);
nor U2533 (N_2533,N_2488,N_2437);
nor U2534 (N_2534,N_2499,N_2496);
or U2535 (N_2535,N_2411,N_2400);
xor U2536 (N_2536,N_2440,N_2401);
nand U2537 (N_2537,N_2457,N_2446);
xor U2538 (N_2538,N_2443,N_2475);
nand U2539 (N_2539,N_2454,N_2495);
and U2540 (N_2540,N_2413,N_2455);
and U2541 (N_2541,N_2486,N_2419);
xor U2542 (N_2542,N_2449,N_2465);
xnor U2543 (N_2543,N_2472,N_2432);
nor U2544 (N_2544,N_2434,N_2485);
nor U2545 (N_2545,N_2462,N_2483);
and U2546 (N_2546,N_2493,N_2489);
nand U2547 (N_2547,N_2445,N_2424);
nand U2548 (N_2548,N_2408,N_2416);
nand U2549 (N_2549,N_2469,N_2467);
or U2550 (N_2550,N_2492,N_2400);
and U2551 (N_2551,N_2490,N_2428);
and U2552 (N_2552,N_2483,N_2499);
nand U2553 (N_2553,N_2439,N_2423);
and U2554 (N_2554,N_2418,N_2406);
nor U2555 (N_2555,N_2415,N_2423);
nand U2556 (N_2556,N_2425,N_2445);
or U2557 (N_2557,N_2468,N_2486);
xor U2558 (N_2558,N_2474,N_2404);
xor U2559 (N_2559,N_2486,N_2437);
xor U2560 (N_2560,N_2466,N_2415);
nor U2561 (N_2561,N_2497,N_2449);
xnor U2562 (N_2562,N_2480,N_2401);
xnor U2563 (N_2563,N_2401,N_2454);
and U2564 (N_2564,N_2476,N_2405);
and U2565 (N_2565,N_2421,N_2476);
or U2566 (N_2566,N_2480,N_2472);
nor U2567 (N_2567,N_2497,N_2466);
nor U2568 (N_2568,N_2418,N_2466);
or U2569 (N_2569,N_2444,N_2478);
and U2570 (N_2570,N_2494,N_2452);
nand U2571 (N_2571,N_2482,N_2427);
nand U2572 (N_2572,N_2485,N_2462);
xor U2573 (N_2573,N_2472,N_2477);
or U2574 (N_2574,N_2427,N_2422);
or U2575 (N_2575,N_2447,N_2499);
or U2576 (N_2576,N_2430,N_2437);
nand U2577 (N_2577,N_2432,N_2416);
or U2578 (N_2578,N_2480,N_2400);
nand U2579 (N_2579,N_2409,N_2482);
and U2580 (N_2580,N_2447,N_2488);
and U2581 (N_2581,N_2466,N_2499);
or U2582 (N_2582,N_2430,N_2497);
nor U2583 (N_2583,N_2449,N_2469);
nand U2584 (N_2584,N_2490,N_2478);
xnor U2585 (N_2585,N_2468,N_2459);
and U2586 (N_2586,N_2474,N_2422);
nor U2587 (N_2587,N_2459,N_2439);
nand U2588 (N_2588,N_2465,N_2481);
nand U2589 (N_2589,N_2438,N_2484);
xnor U2590 (N_2590,N_2491,N_2463);
nor U2591 (N_2591,N_2435,N_2443);
nand U2592 (N_2592,N_2469,N_2409);
xnor U2593 (N_2593,N_2462,N_2488);
xor U2594 (N_2594,N_2446,N_2433);
nand U2595 (N_2595,N_2404,N_2469);
and U2596 (N_2596,N_2452,N_2461);
nor U2597 (N_2597,N_2485,N_2439);
or U2598 (N_2598,N_2428,N_2411);
nand U2599 (N_2599,N_2475,N_2454);
nand U2600 (N_2600,N_2555,N_2564);
nand U2601 (N_2601,N_2508,N_2557);
and U2602 (N_2602,N_2585,N_2528);
nor U2603 (N_2603,N_2535,N_2558);
nand U2604 (N_2604,N_2517,N_2570);
nor U2605 (N_2605,N_2547,N_2537);
nor U2606 (N_2606,N_2589,N_2516);
nand U2607 (N_2607,N_2510,N_2567);
or U2608 (N_2608,N_2526,N_2519);
nand U2609 (N_2609,N_2544,N_2522);
nand U2610 (N_2610,N_2520,N_2506);
or U2611 (N_2611,N_2529,N_2581);
and U2612 (N_2612,N_2550,N_2571);
nand U2613 (N_2613,N_2568,N_2539);
nor U2614 (N_2614,N_2572,N_2566);
nor U2615 (N_2615,N_2504,N_2543);
or U2616 (N_2616,N_2534,N_2562);
nand U2617 (N_2617,N_2592,N_2580);
xnor U2618 (N_2618,N_2561,N_2542);
xnor U2619 (N_2619,N_2521,N_2500);
or U2620 (N_2620,N_2503,N_2559);
xnor U2621 (N_2621,N_2586,N_2587);
nand U2622 (N_2622,N_2591,N_2512);
or U2623 (N_2623,N_2538,N_2584);
nor U2624 (N_2624,N_2598,N_2565);
nand U2625 (N_2625,N_2505,N_2560);
xnor U2626 (N_2626,N_2548,N_2525);
or U2627 (N_2627,N_2590,N_2536);
and U2628 (N_2628,N_2518,N_2514);
nor U2629 (N_2629,N_2574,N_2597);
and U2630 (N_2630,N_2594,N_2593);
xor U2631 (N_2631,N_2577,N_2549);
nor U2632 (N_2632,N_2532,N_2595);
nor U2633 (N_2633,N_2552,N_2513);
and U2634 (N_2634,N_2556,N_2527);
or U2635 (N_2635,N_2540,N_2588);
and U2636 (N_2636,N_2524,N_2563);
and U2637 (N_2637,N_2578,N_2576);
nor U2638 (N_2638,N_2579,N_2583);
xnor U2639 (N_2639,N_2553,N_2530);
or U2640 (N_2640,N_2575,N_2531);
nor U2641 (N_2641,N_2509,N_2551);
and U2642 (N_2642,N_2511,N_2546);
or U2643 (N_2643,N_2596,N_2501);
xnor U2644 (N_2644,N_2502,N_2523);
nand U2645 (N_2645,N_2515,N_2582);
and U2646 (N_2646,N_2507,N_2541);
and U2647 (N_2647,N_2569,N_2554);
xnor U2648 (N_2648,N_2599,N_2545);
and U2649 (N_2649,N_2533,N_2573);
or U2650 (N_2650,N_2539,N_2527);
nor U2651 (N_2651,N_2501,N_2597);
or U2652 (N_2652,N_2539,N_2510);
nor U2653 (N_2653,N_2571,N_2515);
and U2654 (N_2654,N_2590,N_2500);
nand U2655 (N_2655,N_2504,N_2598);
nor U2656 (N_2656,N_2550,N_2582);
nand U2657 (N_2657,N_2570,N_2503);
or U2658 (N_2658,N_2588,N_2593);
nor U2659 (N_2659,N_2504,N_2581);
nor U2660 (N_2660,N_2551,N_2532);
nand U2661 (N_2661,N_2537,N_2555);
and U2662 (N_2662,N_2575,N_2559);
xor U2663 (N_2663,N_2505,N_2574);
xnor U2664 (N_2664,N_2591,N_2577);
nor U2665 (N_2665,N_2561,N_2531);
nor U2666 (N_2666,N_2541,N_2526);
nand U2667 (N_2667,N_2543,N_2557);
xnor U2668 (N_2668,N_2518,N_2583);
and U2669 (N_2669,N_2591,N_2502);
nand U2670 (N_2670,N_2501,N_2570);
nor U2671 (N_2671,N_2584,N_2530);
and U2672 (N_2672,N_2580,N_2589);
or U2673 (N_2673,N_2555,N_2538);
xnor U2674 (N_2674,N_2539,N_2570);
or U2675 (N_2675,N_2522,N_2528);
xor U2676 (N_2676,N_2524,N_2542);
or U2677 (N_2677,N_2594,N_2566);
nand U2678 (N_2678,N_2570,N_2587);
nor U2679 (N_2679,N_2516,N_2578);
xnor U2680 (N_2680,N_2575,N_2549);
nor U2681 (N_2681,N_2564,N_2529);
and U2682 (N_2682,N_2507,N_2501);
nor U2683 (N_2683,N_2522,N_2526);
and U2684 (N_2684,N_2517,N_2535);
and U2685 (N_2685,N_2584,N_2512);
nor U2686 (N_2686,N_2580,N_2579);
nand U2687 (N_2687,N_2556,N_2567);
xor U2688 (N_2688,N_2550,N_2561);
and U2689 (N_2689,N_2542,N_2519);
nor U2690 (N_2690,N_2509,N_2573);
nor U2691 (N_2691,N_2568,N_2542);
nand U2692 (N_2692,N_2561,N_2526);
nor U2693 (N_2693,N_2588,N_2556);
nor U2694 (N_2694,N_2553,N_2584);
or U2695 (N_2695,N_2514,N_2545);
nor U2696 (N_2696,N_2551,N_2556);
xnor U2697 (N_2697,N_2514,N_2589);
and U2698 (N_2698,N_2549,N_2553);
and U2699 (N_2699,N_2508,N_2559);
nor U2700 (N_2700,N_2643,N_2658);
xor U2701 (N_2701,N_2654,N_2674);
nor U2702 (N_2702,N_2675,N_2616);
and U2703 (N_2703,N_2669,N_2696);
nand U2704 (N_2704,N_2629,N_2699);
or U2705 (N_2705,N_2660,N_2615);
and U2706 (N_2706,N_2614,N_2662);
and U2707 (N_2707,N_2644,N_2681);
nor U2708 (N_2708,N_2690,N_2620);
nor U2709 (N_2709,N_2628,N_2683);
nand U2710 (N_2710,N_2655,N_2619);
or U2711 (N_2711,N_2686,N_2639);
and U2712 (N_2712,N_2607,N_2693);
nor U2713 (N_2713,N_2664,N_2665);
and U2714 (N_2714,N_2651,N_2626);
and U2715 (N_2715,N_2601,N_2627);
and U2716 (N_2716,N_2612,N_2691);
xnor U2717 (N_2717,N_2631,N_2680);
and U2718 (N_2718,N_2625,N_2650);
or U2719 (N_2719,N_2688,N_2682);
or U2720 (N_2720,N_2671,N_2640);
and U2721 (N_2721,N_2666,N_2624);
nor U2722 (N_2722,N_2649,N_2668);
nor U2723 (N_2723,N_2630,N_2667);
and U2724 (N_2724,N_2657,N_2633);
nor U2725 (N_2725,N_2670,N_2645);
or U2726 (N_2726,N_2679,N_2689);
nor U2727 (N_2727,N_2678,N_2647);
or U2728 (N_2728,N_2606,N_2684);
or U2729 (N_2729,N_2610,N_2673);
or U2730 (N_2730,N_2636,N_2618);
or U2731 (N_2731,N_2697,N_2642);
nor U2732 (N_2732,N_2661,N_2602);
and U2733 (N_2733,N_2685,N_2687);
nand U2734 (N_2734,N_2617,N_2698);
and U2735 (N_2735,N_2648,N_2672);
xor U2736 (N_2736,N_2663,N_2677);
xor U2737 (N_2737,N_2609,N_2605);
nand U2738 (N_2738,N_2604,N_2653);
xnor U2739 (N_2739,N_2692,N_2632);
nor U2740 (N_2740,N_2676,N_2613);
nor U2741 (N_2741,N_2637,N_2641);
nor U2742 (N_2742,N_2635,N_2695);
nand U2743 (N_2743,N_2638,N_2646);
xnor U2744 (N_2744,N_2634,N_2621);
nand U2745 (N_2745,N_2659,N_2656);
and U2746 (N_2746,N_2652,N_2694);
xor U2747 (N_2747,N_2603,N_2600);
nand U2748 (N_2748,N_2608,N_2622);
nand U2749 (N_2749,N_2611,N_2623);
and U2750 (N_2750,N_2632,N_2663);
or U2751 (N_2751,N_2652,N_2658);
and U2752 (N_2752,N_2696,N_2611);
xor U2753 (N_2753,N_2613,N_2664);
and U2754 (N_2754,N_2668,N_2623);
nand U2755 (N_2755,N_2641,N_2642);
nand U2756 (N_2756,N_2698,N_2618);
nor U2757 (N_2757,N_2652,N_2696);
nor U2758 (N_2758,N_2699,N_2642);
or U2759 (N_2759,N_2630,N_2655);
or U2760 (N_2760,N_2685,N_2686);
xor U2761 (N_2761,N_2698,N_2623);
xnor U2762 (N_2762,N_2641,N_2666);
nand U2763 (N_2763,N_2657,N_2609);
nor U2764 (N_2764,N_2649,N_2680);
and U2765 (N_2765,N_2612,N_2696);
or U2766 (N_2766,N_2694,N_2671);
nor U2767 (N_2767,N_2677,N_2606);
or U2768 (N_2768,N_2699,N_2679);
or U2769 (N_2769,N_2691,N_2619);
nor U2770 (N_2770,N_2610,N_2604);
and U2771 (N_2771,N_2620,N_2614);
xor U2772 (N_2772,N_2642,N_2622);
xnor U2773 (N_2773,N_2644,N_2668);
and U2774 (N_2774,N_2627,N_2686);
or U2775 (N_2775,N_2665,N_2637);
xnor U2776 (N_2776,N_2684,N_2639);
xnor U2777 (N_2777,N_2611,N_2603);
xor U2778 (N_2778,N_2633,N_2662);
or U2779 (N_2779,N_2626,N_2615);
or U2780 (N_2780,N_2693,N_2631);
or U2781 (N_2781,N_2667,N_2601);
xor U2782 (N_2782,N_2672,N_2688);
or U2783 (N_2783,N_2667,N_2636);
nor U2784 (N_2784,N_2612,N_2613);
nor U2785 (N_2785,N_2628,N_2634);
xnor U2786 (N_2786,N_2681,N_2665);
or U2787 (N_2787,N_2651,N_2636);
nor U2788 (N_2788,N_2688,N_2690);
and U2789 (N_2789,N_2608,N_2606);
or U2790 (N_2790,N_2615,N_2623);
nor U2791 (N_2791,N_2661,N_2631);
nand U2792 (N_2792,N_2625,N_2621);
xnor U2793 (N_2793,N_2640,N_2610);
nand U2794 (N_2794,N_2682,N_2639);
nor U2795 (N_2795,N_2616,N_2659);
xor U2796 (N_2796,N_2618,N_2633);
xor U2797 (N_2797,N_2638,N_2684);
nand U2798 (N_2798,N_2629,N_2656);
and U2799 (N_2799,N_2653,N_2677);
xnor U2800 (N_2800,N_2777,N_2746);
nand U2801 (N_2801,N_2783,N_2747);
nor U2802 (N_2802,N_2788,N_2749);
and U2803 (N_2803,N_2753,N_2781);
nor U2804 (N_2804,N_2709,N_2795);
and U2805 (N_2805,N_2755,N_2763);
xor U2806 (N_2806,N_2798,N_2792);
nand U2807 (N_2807,N_2704,N_2791);
nor U2808 (N_2808,N_2725,N_2738);
nand U2809 (N_2809,N_2768,N_2700);
or U2810 (N_2810,N_2732,N_2707);
nand U2811 (N_2811,N_2720,N_2797);
nor U2812 (N_2812,N_2771,N_2784);
or U2813 (N_2813,N_2773,N_2754);
nor U2814 (N_2814,N_2750,N_2734);
and U2815 (N_2815,N_2724,N_2793);
nand U2816 (N_2816,N_2772,N_2718);
nand U2817 (N_2817,N_2702,N_2756);
nand U2818 (N_2818,N_2779,N_2790);
nor U2819 (N_2819,N_2731,N_2726);
or U2820 (N_2820,N_2710,N_2794);
nor U2821 (N_2821,N_2760,N_2785);
nor U2822 (N_2822,N_2742,N_2759);
or U2823 (N_2823,N_2729,N_2719);
nand U2824 (N_2824,N_2789,N_2736);
and U2825 (N_2825,N_2769,N_2730);
nand U2826 (N_2826,N_2723,N_2787);
and U2827 (N_2827,N_2767,N_2766);
and U2828 (N_2828,N_2737,N_2775);
nor U2829 (N_2829,N_2799,N_2735);
or U2830 (N_2830,N_2716,N_2703);
nor U2831 (N_2831,N_2758,N_2774);
xnor U2832 (N_2832,N_2776,N_2714);
nand U2833 (N_2833,N_2701,N_2752);
nand U2834 (N_2834,N_2757,N_2728);
or U2835 (N_2835,N_2765,N_2708);
or U2836 (N_2836,N_2740,N_2717);
or U2837 (N_2837,N_2761,N_2748);
xor U2838 (N_2838,N_2713,N_2745);
nor U2839 (N_2839,N_2764,N_2744);
xor U2840 (N_2840,N_2782,N_2705);
and U2841 (N_2841,N_2711,N_2739);
xnor U2842 (N_2842,N_2786,N_2770);
xor U2843 (N_2843,N_2733,N_2741);
xnor U2844 (N_2844,N_2796,N_2706);
xnor U2845 (N_2845,N_2762,N_2743);
xnor U2846 (N_2846,N_2721,N_2722);
or U2847 (N_2847,N_2751,N_2727);
nand U2848 (N_2848,N_2778,N_2780);
nand U2849 (N_2849,N_2715,N_2712);
xor U2850 (N_2850,N_2737,N_2777);
xor U2851 (N_2851,N_2735,N_2759);
and U2852 (N_2852,N_2728,N_2787);
nand U2853 (N_2853,N_2780,N_2726);
and U2854 (N_2854,N_2747,N_2791);
or U2855 (N_2855,N_2722,N_2772);
or U2856 (N_2856,N_2700,N_2787);
nand U2857 (N_2857,N_2790,N_2756);
nor U2858 (N_2858,N_2795,N_2755);
nand U2859 (N_2859,N_2745,N_2708);
and U2860 (N_2860,N_2775,N_2731);
xnor U2861 (N_2861,N_2785,N_2777);
nor U2862 (N_2862,N_2785,N_2788);
nand U2863 (N_2863,N_2717,N_2714);
nand U2864 (N_2864,N_2741,N_2773);
xor U2865 (N_2865,N_2743,N_2771);
xor U2866 (N_2866,N_2789,N_2742);
nor U2867 (N_2867,N_2777,N_2744);
or U2868 (N_2868,N_2791,N_2777);
xor U2869 (N_2869,N_2753,N_2747);
nor U2870 (N_2870,N_2770,N_2761);
xor U2871 (N_2871,N_2754,N_2708);
or U2872 (N_2872,N_2754,N_2712);
or U2873 (N_2873,N_2744,N_2799);
and U2874 (N_2874,N_2701,N_2742);
xnor U2875 (N_2875,N_2772,N_2758);
xnor U2876 (N_2876,N_2790,N_2770);
or U2877 (N_2877,N_2709,N_2733);
nand U2878 (N_2878,N_2757,N_2781);
xor U2879 (N_2879,N_2715,N_2726);
xnor U2880 (N_2880,N_2749,N_2704);
xor U2881 (N_2881,N_2719,N_2740);
xor U2882 (N_2882,N_2775,N_2798);
nand U2883 (N_2883,N_2761,N_2706);
nand U2884 (N_2884,N_2723,N_2718);
xnor U2885 (N_2885,N_2789,N_2738);
or U2886 (N_2886,N_2727,N_2772);
nor U2887 (N_2887,N_2797,N_2739);
nor U2888 (N_2888,N_2799,N_2795);
and U2889 (N_2889,N_2734,N_2786);
or U2890 (N_2890,N_2780,N_2772);
nand U2891 (N_2891,N_2719,N_2745);
or U2892 (N_2892,N_2780,N_2797);
nand U2893 (N_2893,N_2741,N_2715);
nand U2894 (N_2894,N_2707,N_2712);
or U2895 (N_2895,N_2737,N_2715);
or U2896 (N_2896,N_2768,N_2760);
and U2897 (N_2897,N_2701,N_2708);
nor U2898 (N_2898,N_2780,N_2714);
and U2899 (N_2899,N_2743,N_2774);
xnor U2900 (N_2900,N_2884,N_2892);
or U2901 (N_2901,N_2810,N_2844);
nand U2902 (N_2902,N_2881,N_2813);
and U2903 (N_2903,N_2811,N_2894);
nor U2904 (N_2904,N_2824,N_2871);
nor U2905 (N_2905,N_2817,N_2895);
or U2906 (N_2906,N_2823,N_2841);
or U2907 (N_2907,N_2875,N_2806);
nor U2908 (N_2908,N_2888,N_2865);
nand U2909 (N_2909,N_2826,N_2819);
nor U2910 (N_2910,N_2838,N_2863);
and U2911 (N_2911,N_2887,N_2880);
and U2912 (N_2912,N_2818,N_2803);
or U2913 (N_2913,N_2812,N_2893);
nor U2914 (N_2914,N_2890,N_2854);
xor U2915 (N_2915,N_2801,N_2874);
and U2916 (N_2916,N_2853,N_2847);
nor U2917 (N_2917,N_2883,N_2800);
and U2918 (N_2918,N_2859,N_2885);
and U2919 (N_2919,N_2808,N_2830);
and U2920 (N_2920,N_2867,N_2891);
or U2921 (N_2921,N_2833,N_2843);
nor U2922 (N_2922,N_2816,N_2845);
nand U2923 (N_2923,N_2831,N_2862);
and U2924 (N_2924,N_2815,N_2846);
or U2925 (N_2925,N_2842,N_2825);
or U2926 (N_2926,N_2861,N_2802);
nand U2927 (N_2927,N_2807,N_2835);
or U2928 (N_2928,N_2857,N_2829);
xor U2929 (N_2929,N_2851,N_2856);
nand U2930 (N_2930,N_2828,N_2848);
xor U2931 (N_2931,N_2869,N_2814);
nand U2932 (N_2932,N_2899,N_2873);
or U2933 (N_2933,N_2827,N_2809);
nand U2934 (N_2934,N_2898,N_2877);
and U2935 (N_2935,N_2886,N_2834);
nand U2936 (N_2936,N_2837,N_2872);
and U2937 (N_2937,N_2866,N_2879);
nor U2938 (N_2938,N_2878,N_2860);
and U2939 (N_2939,N_2850,N_2821);
nor U2940 (N_2940,N_2896,N_2876);
nand U2941 (N_2941,N_2805,N_2839);
xnor U2942 (N_2942,N_2897,N_2858);
nand U2943 (N_2943,N_2836,N_2868);
and U2944 (N_2944,N_2889,N_2822);
xor U2945 (N_2945,N_2882,N_2832);
xnor U2946 (N_2946,N_2852,N_2870);
nand U2947 (N_2947,N_2820,N_2804);
and U2948 (N_2948,N_2864,N_2855);
and U2949 (N_2949,N_2840,N_2849);
xor U2950 (N_2950,N_2840,N_2801);
and U2951 (N_2951,N_2852,N_2858);
xnor U2952 (N_2952,N_2840,N_2888);
xor U2953 (N_2953,N_2833,N_2866);
nand U2954 (N_2954,N_2840,N_2879);
xnor U2955 (N_2955,N_2864,N_2881);
xnor U2956 (N_2956,N_2889,N_2842);
xnor U2957 (N_2957,N_2836,N_2842);
xor U2958 (N_2958,N_2848,N_2815);
nor U2959 (N_2959,N_2889,N_2882);
xnor U2960 (N_2960,N_2867,N_2854);
nor U2961 (N_2961,N_2895,N_2896);
nor U2962 (N_2962,N_2840,N_2878);
nand U2963 (N_2963,N_2879,N_2807);
nand U2964 (N_2964,N_2831,N_2878);
or U2965 (N_2965,N_2849,N_2863);
or U2966 (N_2966,N_2801,N_2896);
nor U2967 (N_2967,N_2840,N_2869);
or U2968 (N_2968,N_2855,N_2848);
or U2969 (N_2969,N_2876,N_2870);
and U2970 (N_2970,N_2849,N_2821);
nor U2971 (N_2971,N_2837,N_2860);
or U2972 (N_2972,N_2844,N_2820);
nand U2973 (N_2973,N_2876,N_2872);
nor U2974 (N_2974,N_2886,N_2829);
or U2975 (N_2975,N_2882,N_2894);
xnor U2976 (N_2976,N_2800,N_2826);
nor U2977 (N_2977,N_2845,N_2823);
nor U2978 (N_2978,N_2846,N_2830);
or U2979 (N_2979,N_2815,N_2804);
nand U2980 (N_2980,N_2862,N_2816);
and U2981 (N_2981,N_2827,N_2819);
nand U2982 (N_2982,N_2898,N_2807);
nand U2983 (N_2983,N_2881,N_2808);
nand U2984 (N_2984,N_2828,N_2862);
or U2985 (N_2985,N_2865,N_2835);
nor U2986 (N_2986,N_2849,N_2845);
or U2987 (N_2987,N_2823,N_2876);
xnor U2988 (N_2988,N_2898,N_2899);
nand U2989 (N_2989,N_2842,N_2887);
nor U2990 (N_2990,N_2884,N_2890);
xnor U2991 (N_2991,N_2839,N_2856);
and U2992 (N_2992,N_2884,N_2830);
nor U2993 (N_2993,N_2856,N_2889);
and U2994 (N_2994,N_2891,N_2862);
xnor U2995 (N_2995,N_2834,N_2859);
and U2996 (N_2996,N_2847,N_2834);
xor U2997 (N_2997,N_2823,N_2826);
nand U2998 (N_2998,N_2806,N_2812);
xor U2999 (N_2999,N_2849,N_2864);
xor UO_0 (O_0,N_2927,N_2929);
or UO_1 (O_1,N_2902,N_2910);
xnor UO_2 (O_2,N_2968,N_2945);
and UO_3 (O_3,N_2900,N_2960);
nor UO_4 (O_4,N_2922,N_2939);
nor UO_5 (O_5,N_2967,N_2974);
xnor UO_6 (O_6,N_2937,N_2921);
xnor UO_7 (O_7,N_2957,N_2985);
and UO_8 (O_8,N_2924,N_2958);
and UO_9 (O_9,N_2946,N_2905);
or UO_10 (O_10,N_2949,N_2970);
nor UO_11 (O_11,N_2906,N_2935);
xnor UO_12 (O_12,N_2973,N_2969);
xnor UO_13 (O_13,N_2944,N_2904);
nor UO_14 (O_14,N_2961,N_2978);
or UO_15 (O_15,N_2918,N_2988);
nand UO_16 (O_16,N_2938,N_2954);
xnor UO_17 (O_17,N_2916,N_2920);
or UO_18 (O_18,N_2989,N_2952);
nor UO_19 (O_19,N_2940,N_2925);
and UO_20 (O_20,N_2948,N_2930);
nor UO_21 (O_21,N_2999,N_2934);
or UO_22 (O_22,N_2912,N_2941);
or UO_23 (O_23,N_2908,N_2976);
and UO_24 (O_24,N_2990,N_2980);
xor UO_25 (O_25,N_2975,N_2971);
and UO_26 (O_26,N_2992,N_2907);
nor UO_27 (O_27,N_2919,N_2928);
or UO_28 (O_28,N_2911,N_2981);
nand UO_29 (O_29,N_2986,N_2993);
or UO_30 (O_30,N_2947,N_2901);
nor UO_31 (O_31,N_2951,N_2995);
xnor UO_32 (O_32,N_2966,N_2972);
or UO_33 (O_33,N_2933,N_2959);
nor UO_34 (O_34,N_2932,N_2943);
xor UO_35 (O_35,N_2984,N_2998);
nand UO_36 (O_36,N_2994,N_2926);
nand UO_37 (O_37,N_2977,N_2913);
nor UO_38 (O_38,N_2953,N_2956);
or UO_39 (O_39,N_2923,N_2915);
or UO_40 (O_40,N_2942,N_2931);
or UO_41 (O_41,N_2909,N_2987);
nand UO_42 (O_42,N_2997,N_2979);
and UO_43 (O_43,N_2950,N_2936);
nor UO_44 (O_44,N_2965,N_2996);
nand UO_45 (O_45,N_2917,N_2955);
and UO_46 (O_46,N_2983,N_2982);
nor UO_47 (O_47,N_2962,N_2903);
nor UO_48 (O_48,N_2964,N_2963);
and UO_49 (O_49,N_2991,N_2914);
nand UO_50 (O_50,N_2908,N_2988);
xnor UO_51 (O_51,N_2922,N_2924);
nand UO_52 (O_52,N_2928,N_2986);
or UO_53 (O_53,N_2959,N_2991);
or UO_54 (O_54,N_2915,N_2922);
xnor UO_55 (O_55,N_2919,N_2901);
xnor UO_56 (O_56,N_2908,N_2936);
and UO_57 (O_57,N_2909,N_2942);
and UO_58 (O_58,N_2931,N_2954);
nand UO_59 (O_59,N_2980,N_2960);
xor UO_60 (O_60,N_2988,N_2932);
or UO_61 (O_61,N_2955,N_2961);
xnor UO_62 (O_62,N_2944,N_2996);
nor UO_63 (O_63,N_2995,N_2982);
nor UO_64 (O_64,N_2987,N_2981);
nand UO_65 (O_65,N_2937,N_2927);
nand UO_66 (O_66,N_2900,N_2920);
nand UO_67 (O_67,N_2953,N_2936);
nor UO_68 (O_68,N_2931,N_2950);
nor UO_69 (O_69,N_2972,N_2960);
or UO_70 (O_70,N_2981,N_2909);
or UO_71 (O_71,N_2946,N_2961);
or UO_72 (O_72,N_2905,N_2997);
or UO_73 (O_73,N_2997,N_2925);
xor UO_74 (O_74,N_2988,N_2977);
or UO_75 (O_75,N_2912,N_2983);
nand UO_76 (O_76,N_2954,N_2952);
nor UO_77 (O_77,N_2975,N_2923);
nand UO_78 (O_78,N_2983,N_2991);
nand UO_79 (O_79,N_2900,N_2941);
xnor UO_80 (O_80,N_2957,N_2963);
and UO_81 (O_81,N_2946,N_2913);
and UO_82 (O_82,N_2948,N_2912);
nor UO_83 (O_83,N_2915,N_2989);
and UO_84 (O_84,N_2902,N_2906);
and UO_85 (O_85,N_2996,N_2907);
or UO_86 (O_86,N_2963,N_2944);
and UO_87 (O_87,N_2906,N_2908);
and UO_88 (O_88,N_2929,N_2932);
or UO_89 (O_89,N_2917,N_2944);
and UO_90 (O_90,N_2922,N_2992);
xor UO_91 (O_91,N_2956,N_2979);
xnor UO_92 (O_92,N_2999,N_2980);
xor UO_93 (O_93,N_2939,N_2937);
and UO_94 (O_94,N_2956,N_2991);
or UO_95 (O_95,N_2979,N_2936);
nor UO_96 (O_96,N_2938,N_2928);
nand UO_97 (O_97,N_2953,N_2969);
and UO_98 (O_98,N_2938,N_2918);
nor UO_99 (O_99,N_2943,N_2982);
xor UO_100 (O_100,N_2972,N_2928);
xnor UO_101 (O_101,N_2964,N_2930);
nor UO_102 (O_102,N_2905,N_2974);
xnor UO_103 (O_103,N_2931,N_2998);
xor UO_104 (O_104,N_2934,N_2984);
xnor UO_105 (O_105,N_2943,N_2980);
nand UO_106 (O_106,N_2985,N_2905);
or UO_107 (O_107,N_2911,N_2944);
or UO_108 (O_108,N_2998,N_2945);
xnor UO_109 (O_109,N_2927,N_2930);
xnor UO_110 (O_110,N_2936,N_2957);
xor UO_111 (O_111,N_2946,N_2933);
or UO_112 (O_112,N_2992,N_2963);
or UO_113 (O_113,N_2997,N_2957);
nand UO_114 (O_114,N_2978,N_2928);
or UO_115 (O_115,N_2983,N_2940);
nand UO_116 (O_116,N_2938,N_2919);
or UO_117 (O_117,N_2947,N_2952);
or UO_118 (O_118,N_2939,N_2908);
nand UO_119 (O_119,N_2968,N_2993);
and UO_120 (O_120,N_2921,N_2949);
or UO_121 (O_121,N_2974,N_2997);
nor UO_122 (O_122,N_2919,N_2926);
or UO_123 (O_123,N_2973,N_2953);
or UO_124 (O_124,N_2917,N_2921);
or UO_125 (O_125,N_2926,N_2958);
xnor UO_126 (O_126,N_2937,N_2902);
and UO_127 (O_127,N_2996,N_2955);
and UO_128 (O_128,N_2990,N_2991);
nand UO_129 (O_129,N_2969,N_2929);
xor UO_130 (O_130,N_2952,N_2974);
or UO_131 (O_131,N_2987,N_2995);
and UO_132 (O_132,N_2903,N_2954);
nor UO_133 (O_133,N_2945,N_2962);
nand UO_134 (O_134,N_2944,N_2935);
nor UO_135 (O_135,N_2932,N_2905);
xnor UO_136 (O_136,N_2974,N_2965);
nand UO_137 (O_137,N_2963,N_2932);
and UO_138 (O_138,N_2957,N_2924);
nor UO_139 (O_139,N_2955,N_2926);
xor UO_140 (O_140,N_2948,N_2933);
xnor UO_141 (O_141,N_2982,N_2994);
nor UO_142 (O_142,N_2961,N_2929);
xnor UO_143 (O_143,N_2974,N_2912);
xnor UO_144 (O_144,N_2971,N_2918);
nor UO_145 (O_145,N_2968,N_2935);
xor UO_146 (O_146,N_2949,N_2994);
and UO_147 (O_147,N_2995,N_2976);
nand UO_148 (O_148,N_2986,N_2923);
and UO_149 (O_149,N_2997,N_2968);
xor UO_150 (O_150,N_2927,N_2973);
xnor UO_151 (O_151,N_2969,N_2981);
nand UO_152 (O_152,N_2910,N_2963);
nand UO_153 (O_153,N_2911,N_2988);
nor UO_154 (O_154,N_2962,N_2936);
nand UO_155 (O_155,N_2987,N_2941);
nand UO_156 (O_156,N_2940,N_2990);
xor UO_157 (O_157,N_2974,N_2935);
nand UO_158 (O_158,N_2923,N_2933);
nand UO_159 (O_159,N_2922,N_2976);
nand UO_160 (O_160,N_2936,N_2960);
xor UO_161 (O_161,N_2986,N_2991);
xor UO_162 (O_162,N_2982,N_2965);
nor UO_163 (O_163,N_2945,N_2905);
and UO_164 (O_164,N_2950,N_2940);
xnor UO_165 (O_165,N_2904,N_2961);
or UO_166 (O_166,N_2920,N_2973);
nor UO_167 (O_167,N_2975,N_2999);
and UO_168 (O_168,N_2950,N_2946);
nor UO_169 (O_169,N_2949,N_2990);
nand UO_170 (O_170,N_2999,N_2910);
nor UO_171 (O_171,N_2976,N_2931);
or UO_172 (O_172,N_2944,N_2961);
nor UO_173 (O_173,N_2933,N_2912);
xnor UO_174 (O_174,N_2977,N_2970);
nor UO_175 (O_175,N_2973,N_2916);
or UO_176 (O_176,N_2960,N_2998);
nor UO_177 (O_177,N_2916,N_2906);
nor UO_178 (O_178,N_2970,N_2933);
xnor UO_179 (O_179,N_2956,N_2982);
or UO_180 (O_180,N_2959,N_2927);
xnor UO_181 (O_181,N_2981,N_2931);
and UO_182 (O_182,N_2990,N_2924);
xnor UO_183 (O_183,N_2906,N_2951);
nor UO_184 (O_184,N_2956,N_2919);
and UO_185 (O_185,N_2935,N_2909);
xnor UO_186 (O_186,N_2954,N_2974);
xor UO_187 (O_187,N_2964,N_2900);
nor UO_188 (O_188,N_2908,N_2905);
or UO_189 (O_189,N_2922,N_2920);
xor UO_190 (O_190,N_2943,N_2974);
or UO_191 (O_191,N_2965,N_2962);
nor UO_192 (O_192,N_2980,N_2912);
xnor UO_193 (O_193,N_2907,N_2958);
or UO_194 (O_194,N_2944,N_2955);
xor UO_195 (O_195,N_2980,N_2924);
or UO_196 (O_196,N_2929,N_2919);
nor UO_197 (O_197,N_2955,N_2914);
nand UO_198 (O_198,N_2996,N_2922);
nand UO_199 (O_199,N_2918,N_2946);
or UO_200 (O_200,N_2934,N_2976);
and UO_201 (O_201,N_2901,N_2962);
or UO_202 (O_202,N_2915,N_2931);
or UO_203 (O_203,N_2999,N_2983);
or UO_204 (O_204,N_2981,N_2995);
or UO_205 (O_205,N_2990,N_2926);
and UO_206 (O_206,N_2901,N_2966);
nand UO_207 (O_207,N_2967,N_2945);
xor UO_208 (O_208,N_2928,N_2971);
xnor UO_209 (O_209,N_2954,N_2907);
or UO_210 (O_210,N_2964,N_2947);
xor UO_211 (O_211,N_2914,N_2968);
xor UO_212 (O_212,N_2919,N_2948);
or UO_213 (O_213,N_2947,N_2981);
nand UO_214 (O_214,N_2953,N_2980);
nand UO_215 (O_215,N_2985,N_2986);
or UO_216 (O_216,N_2956,N_2947);
xnor UO_217 (O_217,N_2929,N_2948);
xor UO_218 (O_218,N_2934,N_2986);
or UO_219 (O_219,N_2904,N_2939);
and UO_220 (O_220,N_2977,N_2934);
xor UO_221 (O_221,N_2915,N_2943);
nand UO_222 (O_222,N_2966,N_2954);
xor UO_223 (O_223,N_2913,N_2917);
nand UO_224 (O_224,N_2937,N_2981);
or UO_225 (O_225,N_2976,N_2911);
or UO_226 (O_226,N_2986,N_2918);
nor UO_227 (O_227,N_2926,N_2920);
and UO_228 (O_228,N_2954,N_2912);
and UO_229 (O_229,N_2995,N_2913);
and UO_230 (O_230,N_2981,N_2940);
nand UO_231 (O_231,N_2971,N_2934);
nand UO_232 (O_232,N_2956,N_2958);
xnor UO_233 (O_233,N_2940,N_2938);
nand UO_234 (O_234,N_2947,N_2959);
nor UO_235 (O_235,N_2937,N_2904);
nand UO_236 (O_236,N_2959,N_2948);
xnor UO_237 (O_237,N_2992,N_2980);
or UO_238 (O_238,N_2982,N_2966);
nand UO_239 (O_239,N_2908,N_2978);
or UO_240 (O_240,N_2994,N_2961);
xor UO_241 (O_241,N_2906,N_2960);
nand UO_242 (O_242,N_2908,N_2913);
or UO_243 (O_243,N_2969,N_2918);
or UO_244 (O_244,N_2942,N_2978);
or UO_245 (O_245,N_2999,N_2998);
and UO_246 (O_246,N_2973,N_2921);
and UO_247 (O_247,N_2956,N_2966);
nand UO_248 (O_248,N_2964,N_2924);
nand UO_249 (O_249,N_2956,N_2926);
and UO_250 (O_250,N_2917,N_2957);
xor UO_251 (O_251,N_2975,N_2964);
nand UO_252 (O_252,N_2940,N_2936);
xor UO_253 (O_253,N_2985,N_2969);
or UO_254 (O_254,N_2996,N_2909);
xor UO_255 (O_255,N_2983,N_2956);
and UO_256 (O_256,N_2935,N_2901);
xor UO_257 (O_257,N_2962,N_2997);
and UO_258 (O_258,N_2961,N_2977);
nor UO_259 (O_259,N_2958,N_2911);
nor UO_260 (O_260,N_2939,N_2926);
nor UO_261 (O_261,N_2971,N_2980);
nor UO_262 (O_262,N_2905,N_2967);
xor UO_263 (O_263,N_2974,N_2959);
and UO_264 (O_264,N_2964,N_2937);
xor UO_265 (O_265,N_2973,N_2947);
nand UO_266 (O_266,N_2900,N_2902);
nand UO_267 (O_267,N_2924,N_2997);
nor UO_268 (O_268,N_2922,N_2949);
nor UO_269 (O_269,N_2994,N_2991);
and UO_270 (O_270,N_2902,N_2974);
or UO_271 (O_271,N_2957,N_2910);
nor UO_272 (O_272,N_2926,N_2989);
nor UO_273 (O_273,N_2941,N_2925);
or UO_274 (O_274,N_2934,N_2911);
nor UO_275 (O_275,N_2960,N_2921);
and UO_276 (O_276,N_2945,N_2953);
and UO_277 (O_277,N_2952,N_2925);
nand UO_278 (O_278,N_2972,N_2941);
or UO_279 (O_279,N_2999,N_2935);
xor UO_280 (O_280,N_2905,N_2929);
nand UO_281 (O_281,N_2905,N_2980);
xnor UO_282 (O_282,N_2976,N_2902);
nand UO_283 (O_283,N_2936,N_2986);
or UO_284 (O_284,N_2991,N_2922);
or UO_285 (O_285,N_2914,N_2951);
or UO_286 (O_286,N_2900,N_2983);
nand UO_287 (O_287,N_2943,N_2936);
and UO_288 (O_288,N_2947,N_2954);
nor UO_289 (O_289,N_2964,N_2925);
and UO_290 (O_290,N_2905,N_2996);
or UO_291 (O_291,N_2911,N_2959);
xor UO_292 (O_292,N_2971,N_2992);
nor UO_293 (O_293,N_2951,N_2943);
nand UO_294 (O_294,N_2953,N_2923);
and UO_295 (O_295,N_2940,N_2934);
nor UO_296 (O_296,N_2992,N_2925);
and UO_297 (O_297,N_2903,N_2974);
and UO_298 (O_298,N_2991,N_2967);
nor UO_299 (O_299,N_2957,N_2967);
and UO_300 (O_300,N_2940,N_2927);
and UO_301 (O_301,N_2956,N_2929);
xor UO_302 (O_302,N_2961,N_2950);
or UO_303 (O_303,N_2931,N_2984);
or UO_304 (O_304,N_2980,N_2938);
nor UO_305 (O_305,N_2998,N_2911);
and UO_306 (O_306,N_2945,N_2907);
nor UO_307 (O_307,N_2942,N_2922);
or UO_308 (O_308,N_2945,N_2975);
and UO_309 (O_309,N_2962,N_2966);
nor UO_310 (O_310,N_2957,N_2941);
or UO_311 (O_311,N_2962,N_2917);
and UO_312 (O_312,N_2988,N_2957);
nor UO_313 (O_313,N_2980,N_2954);
or UO_314 (O_314,N_2964,N_2903);
nand UO_315 (O_315,N_2986,N_2983);
nor UO_316 (O_316,N_2946,N_2972);
nand UO_317 (O_317,N_2980,N_2937);
xor UO_318 (O_318,N_2921,N_2926);
xnor UO_319 (O_319,N_2942,N_2936);
nand UO_320 (O_320,N_2914,N_2917);
nor UO_321 (O_321,N_2951,N_2926);
nor UO_322 (O_322,N_2942,N_2960);
nor UO_323 (O_323,N_2900,N_2966);
nor UO_324 (O_324,N_2994,N_2984);
and UO_325 (O_325,N_2950,N_2969);
and UO_326 (O_326,N_2971,N_2993);
and UO_327 (O_327,N_2993,N_2913);
or UO_328 (O_328,N_2926,N_2933);
nand UO_329 (O_329,N_2975,N_2984);
xnor UO_330 (O_330,N_2906,N_2958);
nor UO_331 (O_331,N_2950,N_2984);
or UO_332 (O_332,N_2940,N_2963);
nor UO_333 (O_333,N_2931,N_2999);
and UO_334 (O_334,N_2979,N_2953);
nand UO_335 (O_335,N_2929,N_2960);
xor UO_336 (O_336,N_2990,N_2984);
or UO_337 (O_337,N_2997,N_2983);
nand UO_338 (O_338,N_2902,N_2909);
xor UO_339 (O_339,N_2983,N_2919);
nor UO_340 (O_340,N_2939,N_2907);
or UO_341 (O_341,N_2957,N_2909);
or UO_342 (O_342,N_2939,N_2946);
nor UO_343 (O_343,N_2909,N_2908);
and UO_344 (O_344,N_2916,N_2980);
nand UO_345 (O_345,N_2984,N_2971);
or UO_346 (O_346,N_2958,N_2989);
xor UO_347 (O_347,N_2984,N_2919);
or UO_348 (O_348,N_2993,N_2932);
and UO_349 (O_349,N_2932,N_2973);
xnor UO_350 (O_350,N_2914,N_2969);
and UO_351 (O_351,N_2913,N_2964);
nand UO_352 (O_352,N_2946,N_2958);
or UO_353 (O_353,N_2966,N_2955);
and UO_354 (O_354,N_2994,N_2922);
or UO_355 (O_355,N_2945,N_2987);
nor UO_356 (O_356,N_2996,N_2935);
and UO_357 (O_357,N_2939,N_2925);
nor UO_358 (O_358,N_2976,N_2903);
nand UO_359 (O_359,N_2983,N_2962);
and UO_360 (O_360,N_2989,N_2982);
nor UO_361 (O_361,N_2900,N_2917);
nor UO_362 (O_362,N_2904,N_2973);
xor UO_363 (O_363,N_2942,N_2952);
and UO_364 (O_364,N_2967,N_2901);
xnor UO_365 (O_365,N_2954,N_2996);
xor UO_366 (O_366,N_2953,N_2929);
nor UO_367 (O_367,N_2911,N_2994);
nor UO_368 (O_368,N_2917,N_2908);
nor UO_369 (O_369,N_2928,N_2905);
and UO_370 (O_370,N_2975,N_2921);
xnor UO_371 (O_371,N_2936,N_2922);
nor UO_372 (O_372,N_2934,N_2921);
nand UO_373 (O_373,N_2957,N_2969);
xnor UO_374 (O_374,N_2924,N_2906);
xnor UO_375 (O_375,N_2936,N_2939);
nand UO_376 (O_376,N_2934,N_2956);
and UO_377 (O_377,N_2948,N_2984);
nand UO_378 (O_378,N_2914,N_2986);
or UO_379 (O_379,N_2982,N_2998);
and UO_380 (O_380,N_2934,N_2989);
xor UO_381 (O_381,N_2979,N_2960);
nor UO_382 (O_382,N_2998,N_2970);
and UO_383 (O_383,N_2946,N_2973);
or UO_384 (O_384,N_2966,N_2949);
or UO_385 (O_385,N_2960,N_2922);
nand UO_386 (O_386,N_2938,N_2922);
nor UO_387 (O_387,N_2984,N_2969);
and UO_388 (O_388,N_2924,N_2927);
or UO_389 (O_389,N_2915,N_2920);
or UO_390 (O_390,N_2992,N_2906);
nand UO_391 (O_391,N_2960,N_2995);
and UO_392 (O_392,N_2997,N_2964);
nand UO_393 (O_393,N_2900,N_2954);
and UO_394 (O_394,N_2911,N_2954);
or UO_395 (O_395,N_2941,N_2919);
and UO_396 (O_396,N_2976,N_2954);
nor UO_397 (O_397,N_2940,N_2987);
nor UO_398 (O_398,N_2987,N_2939);
or UO_399 (O_399,N_2997,N_2977);
nand UO_400 (O_400,N_2911,N_2949);
nor UO_401 (O_401,N_2944,N_2965);
and UO_402 (O_402,N_2987,N_2933);
and UO_403 (O_403,N_2921,N_2948);
nand UO_404 (O_404,N_2970,N_2984);
nor UO_405 (O_405,N_2994,N_2908);
xor UO_406 (O_406,N_2925,N_2990);
nand UO_407 (O_407,N_2928,N_2914);
and UO_408 (O_408,N_2914,N_2931);
nor UO_409 (O_409,N_2959,N_2957);
nand UO_410 (O_410,N_2969,N_2980);
nor UO_411 (O_411,N_2995,N_2945);
or UO_412 (O_412,N_2971,N_2909);
xor UO_413 (O_413,N_2962,N_2926);
nor UO_414 (O_414,N_2972,N_2981);
or UO_415 (O_415,N_2922,N_2923);
or UO_416 (O_416,N_2993,N_2952);
nor UO_417 (O_417,N_2933,N_2915);
xnor UO_418 (O_418,N_2904,N_2956);
nor UO_419 (O_419,N_2993,N_2927);
and UO_420 (O_420,N_2986,N_2905);
xor UO_421 (O_421,N_2931,N_2983);
nand UO_422 (O_422,N_2945,N_2929);
and UO_423 (O_423,N_2972,N_2969);
and UO_424 (O_424,N_2988,N_2968);
or UO_425 (O_425,N_2965,N_2964);
nand UO_426 (O_426,N_2983,N_2904);
and UO_427 (O_427,N_2907,N_2901);
nor UO_428 (O_428,N_2979,N_2931);
xor UO_429 (O_429,N_2933,N_2900);
nand UO_430 (O_430,N_2960,N_2904);
and UO_431 (O_431,N_2990,N_2946);
nand UO_432 (O_432,N_2924,N_2911);
and UO_433 (O_433,N_2971,N_2981);
nor UO_434 (O_434,N_2937,N_2908);
nor UO_435 (O_435,N_2916,N_2991);
nor UO_436 (O_436,N_2932,N_2979);
nand UO_437 (O_437,N_2913,N_2967);
nand UO_438 (O_438,N_2928,N_2935);
xor UO_439 (O_439,N_2957,N_2986);
or UO_440 (O_440,N_2961,N_2942);
and UO_441 (O_441,N_2953,N_2982);
nand UO_442 (O_442,N_2975,N_2915);
and UO_443 (O_443,N_2911,N_2970);
and UO_444 (O_444,N_2954,N_2997);
and UO_445 (O_445,N_2937,N_2956);
or UO_446 (O_446,N_2932,N_2924);
or UO_447 (O_447,N_2902,N_2952);
xnor UO_448 (O_448,N_2982,N_2922);
and UO_449 (O_449,N_2977,N_2923);
or UO_450 (O_450,N_2990,N_2992);
or UO_451 (O_451,N_2944,N_2985);
and UO_452 (O_452,N_2950,N_2914);
nor UO_453 (O_453,N_2972,N_2912);
nor UO_454 (O_454,N_2996,N_2977);
nand UO_455 (O_455,N_2906,N_2927);
or UO_456 (O_456,N_2986,N_2921);
nor UO_457 (O_457,N_2921,N_2965);
xor UO_458 (O_458,N_2964,N_2927);
and UO_459 (O_459,N_2963,N_2916);
xor UO_460 (O_460,N_2971,N_2948);
or UO_461 (O_461,N_2993,N_2953);
and UO_462 (O_462,N_2941,N_2907);
and UO_463 (O_463,N_2978,N_2968);
nand UO_464 (O_464,N_2910,N_2946);
or UO_465 (O_465,N_2994,N_2919);
or UO_466 (O_466,N_2998,N_2913);
and UO_467 (O_467,N_2909,N_2990);
nand UO_468 (O_468,N_2910,N_2973);
or UO_469 (O_469,N_2953,N_2965);
or UO_470 (O_470,N_2985,N_2907);
xnor UO_471 (O_471,N_2902,N_2964);
or UO_472 (O_472,N_2940,N_2992);
or UO_473 (O_473,N_2948,N_2972);
or UO_474 (O_474,N_2987,N_2906);
nand UO_475 (O_475,N_2987,N_2908);
or UO_476 (O_476,N_2990,N_2905);
nand UO_477 (O_477,N_2964,N_2992);
nand UO_478 (O_478,N_2993,N_2995);
nand UO_479 (O_479,N_2986,N_2924);
and UO_480 (O_480,N_2959,N_2918);
nand UO_481 (O_481,N_2968,N_2970);
nand UO_482 (O_482,N_2973,N_2985);
xor UO_483 (O_483,N_2943,N_2959);
nor UO_484 (O_484,N_2935,N_2918);
nor UO_485 (O_485,N_2957,N_2978);
or UO_486 (O_486,N_2933,N_2943);
nand UO_487 (O_487,N_2917,N_2971);
xnor UO_488 (O_488,N_2951,N_2997);
and UO_489 (O_489,N_2940,N_2908);
xnor UO_490 (O_490,N_2948,N_2962);
xnor UO_491 (O_491,N_2917,N_2976);
nor UO_492 (O_492,N_2996,N_2948);
nand UO_493 (O_493,N_2954,N_2932);
or UO_494 (O_494,N_2999,N_2987);
xor UO_495 (O_495,N_2986,N_2980);
nor UO_496 (O_496,N_2902,N_2984);
or UO_497 (O_497,N_2932,N_2903);
xnor UO_498 (O_498,N_2916,N_2942);
nand UO_499 (O_499,N_2920,N_2951);
endmodule