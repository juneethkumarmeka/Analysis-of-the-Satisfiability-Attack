module basic_1500_15000_2000_75_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_1018,In_449);
xor U1 (N_1,In_63,In_1176);
nor U2 (N_2,In_13,In_959);
and U3 (N_3,In_254,In_1145);
nand U4 (N_4,In_1137,In_239);
and U5 (N_5,In_1143,In_1240);
or U6 (N_6,In_1299,In_87);
or U7 (N_7,In_1188,In_709);
nand U8 (N_8,In_174,In_19);
or U9 (N_9,In_981,In_197);
or U10 (N_10,In_4,In_88);
xor U11 (N_11,In_1051,In_527);
or U12 (N_12,In_1210,In_646);
xnor U13 (N_13,In_1469,In_894);
and U14 (N_14,In_1396,In_887);
nand U15 (N_15,In_1477,In_987);
nand U16 (N_16,In_1057,In_587);
nand U17 (N_17,In_274,In_191);
and U18 (N_18,In_1433,In_794);
nand U19 (N_19,In_602,In_1474);
nor U20 (N_20,In_1339,In_958);
nor U21 (N_21,In_1411,In_100);
nor U22 (N_22,In_360,In_864);
nor U23 (N_23,In_660,In_621);
or U24 (N_24,In_461,In_681);
xnor U25 (N_25,In_719,In_940);
nor U26 (N_26,In_640,In_653);
xnor U27 (N_27,In_1096,In_447);
or U28 (N_28,In_462,In_1330);
xnor U29 (N_29,In_608,In_1295);
or U30 (N_30,In_193,In_977);
xor U31 (N_31,In_976,In_223);
or U32 (N_32,In_1298,In_624);
xor U33 (N_33,In_213,In_217);
and U34 (N_34,In_346,In_91);
or U35 (N_35,In_993,In_1480);
or U36 (N_36,In_384,In_1164);
nand U37 (N_37,In_968,In_1211);
nor U38 (N_38,In_1226,In_1366);
nor U39 (N_39,In_943,In_1276);
nor U40 (N_40,In_249,In_1431);
nor U41 (N_41,In_1213,In_1268);
or U42 (N_42,In_588,In_1093);
nand U43 (N_43,In_356,In_1252);
xor U44 (N_44,In_130,In_122);
nand U45 (N_45,In_324,In_766);
or U46 (N_46,In_898,In_720);
nand U47 (N_47,In_378,In_158);
nand U48 (N_48,In_489,In_281);
nand U49 (N_49,In_181,In_634);
and U50 (N_50,In_851,In_259);
xor U51 (N_51,In_994,In_1462);
nand U52 (N_52,In_305,In_760);
xnor U53 (N_53,In_882,In_875);
and U54 (N_54,In_1418,In_1003);
or U55 (N_55,In_220,In_1364);
xor U56 (N_56,In_534,In_497);
or U57 (N_57,In_1373,In_62);
or U58 (N_58,In_54,In_1490);
xnor U59 (N_59,In_573,In_836);
and U60 (N_60,In_702,In_674);
and U61 (N_61,In_937,In_874);
nand U62 (N_62,In_800,In_370);
nand U63 (N_63,In_403,In_770);
xor U64 (N_64,In_1390,In_1494);
or U65 (N_65,In_765,In_1478);
xor U66 (N_66,In_1125,In_355);
nand U67 (N_67,In_435,In_1231);
nand U68 (N_68,In_715,In_811);
nor U69 (N_69,In_1269,In_1254);
and U70 (N_70,In_605,In_893);
or U71 (N_71,In_885,In_869);
nand U72 (N_72,In_164,In_503);
xor U73 (N_73,In_858,In_1363);
and U74 (N_74,In_1009,In_1283);
nor U75 (N_75,In_102,In_73);
xnor U76 (N_76,In_601,In_11);
and U77 (N_77,In_1230,In_843);
and U78 (N_78,In_1484,In_988);
nand U79 (N_79,In_647,In_219);
or U80 (N_80,In_593,In_7);
nand U81 (N_81,In_764,In_433);
and U82 (N_82,In_597,In_1380);
nand U83 (N_83,In_1225,In_756);
or U84 (N_84,In_275,In_973);
or U85 (N_85,In_157,In_545);
xor U86 (N_86,In_257,In_468);
and U87 (N_87,In_1090,In_498);
nand U88 (N_88,In_1289,In_1062);
nand U89 (N_89,In_300,In_1136);
or U90 (N_90,In_532,In_486);
or U91 (N_91,In_149,In_1346);
nand U92 (N_92,In_1201,In_758);
xor U93 (N_93,In_31,In_1098);
xor U94 (N_94,In_10,In_114);
nand U95 (N_95,In_1227,In_1453);
nand U96 (N_96,In_997,In_1050);
nand U97 (N_97,In_513,In_901);
xor U98 (N_98,In_404,In_1218);
or U99 (N_99,In_1250,In_746);
and U100 (N_100,In_628,In_1116);
nand U101 (N_101,In_1005,In_549);
xnor U102 (N_102,In_975,In_412);
nor U103 (N_103,In_1069,In_1306);
nor U104 (N_104,In_1497,In_721);
nor U105 (N_105,In_1401,In_670);
or U106 (N_106,In_312,In_866);
nor U107 (N_107,In_1161,In_294);
or U108 (N_108,In_1452,In_71);
nor U109 (N_109,In_1479,In_547);
xor U110 (N_110,In_451,In_1040);
xnor U111 (N_111,In_0,In_290);
nor U112 (N_112,In_1159,In_36);
nor U113 (N_113,In_878,In_853);
nor U114 (N_114,In_1142,In_590);
nand U115 (N_115,In_1312,In_38);
or U116 (N_116,In_1154,In_358);
nand U117 (N_117,In_1444,In_210);
nor U118 (N_118,In_339,In_829);
nor U119 (N_119,In_798,In_1436);
or U120 (N_120,In_94,In_134);
xnor U121 (N_121,In_753,In_82);
nand U122 (N_122,In_331,In_342);
and U123 (N_123,In_110,In_891);
xor U124 (N_124,In_790,In_662);
nor U125 (N_125,In_1456,In_1360);
nand U126 (N_126,In_292,In_938);
or U127 (N_127,In_852,In_778);
nor U128 (N_128,In_1322,In_881);
and U129 (N_129,In_454,In_242);
nor U130 (N_130,In_373,In_782);
nor U131 (N_131,In_791,In_802);
nand U132 (N_132,In_614,In_804);
nand U133 (N_133,In_345,In_326);
and U134 (N_134,In_1429,In_47);
xnor U135 (N_135,In_1180,In_491);
xnor U136 (N_136,In_84,In_1435);
xor U137 (N_137,In_734,In_1476);
or U138 (N_138,In_518,In_168);
nand U139 (N_139,In_1020,In_1190);
xnor U140 (N_140,In_850,In_320);
or U141 (N_141,In_1031,In_788);
nor U142 (N_142,In_1006,In_1427);
nor U143 (N_143,In_970,In_27);
or U144 (N_144,In_99,In_432);
and U145 (N_145,In_707,In_932);
nor U146 (N_146,In_904,In_1056);
and U147 (N_147,In_382,In_604);
xnor U148 (N_148,In_946,In_278);
or U149 (N_149,In_1319,In_317);
or U150 (N_150,In_1167,In_125);
xor U151 (N_151,In_437,In_1114);
nor U152 (N_152,In_1199,In_58);
nor U153 (N_153,In_934,In_1129);
or U154 (N_154,In_495,In_199);
or U155 (N_155,In_920,In_446);
and U156 (N_156,In_761,In_828);
xor U157 (N_157,In_786,In_944);
nor U158 (N_158,In_1459,In_809);
or U159 (N_159,In_1486,In_1148);
or U160 (N_160,In_550,In_1078);
or U161 (N_161,In_961,In_632);
and U162 (N_162,In_135,In_948);
and U163 (N_163,In_727,In_467);
and U164 (N_164,In_659,In_586);
and U165 (N_165,In_35,In_1035);
and U166 (N_166,In_66,In_733);
or U167 (N_167,In_309,In_949);
and U168 (N_168,In_1389,In_677);
nor U169 (N_169,In_1328,In_1237);
and U170 (N_170,In_827,In_673);
xnor U171 (N_171,In_53,In_424);
or U172 (N_172,In_444,In_178);
nand U173 (N_173,In_1214,In_1282);
xor U174 (N_174,In_921,In_595);
and U175 (N_175,In_1023,In_815);
nand U176 (N_176,In_907,In_1262);
nand U177 (N_177,In_1158,In_540);
or U178 (N_178,In_234,In_411);
nor U179 (N_179,In_289,In_385);
and U180 (N_180,In_9,In_1464);
or U181 (N_181,In_1068,In_631);
xor U182 (N_182,In_1160,In_162);
and U183 (N_183,In_147,In_1156);
or U184 (N_184,In_405,In_1202);
nand U185 (N_185,In_1080,In_426);
xor U186 (N_186,In_338,In_349);
or U187 (N_187,In_501,In_688);
and U188 (N_188,In_472,In_931);
nand U189 (N_189,In_1095,In_777);
or U190 (N_190,In_722,In_926);
nor U191 (N_191,In_1046,In_214);
xnor U192 (N_192,In_22,In_554);
and U193 (N_193,In_415,In_150);
nor U194 (N_194,In_256,In_1323);
xor U195 (N_195,In_839,In_916);
nor U196 (N_196,In_189,In_969);
nand U197 (N_197,In_1343,In_589);
or U198 (N_198,In_78,In_1404);
or U199 (N_199,In_801,In_179);
xor U200 (N_200,In_485,In_1384);
nand U201 (N_201,In_1382,In_45);
nor U202 (N_202,In_572,In_268);
nand U203 (N_203,In_354,In_1197);
and U204 (N_204,In_960,N_57);
nand U205 (N_205,In_129,In_111);
and U206 (N_206,N_80,In_1445);
or U207 (N_207,In_516,In_70);
or U208 (N_208,In_1087,In_1398);
nor U209 (N_209,In_103,In_156);
nor U210 (N_210,In_1263,In_711);
xor U211 (N_211,N_93,In_871);
xor U212 (N_212,In_701,In_398);
or U213 (N_213,In_1241,In_1126);
nand U214 (N_214,In_1152,In_1030);
xnor U215 (N_215,In_951,In_972);
nand U216 (N_216,N_175,In_522);
nor U217 (N_217,In_287,In_1165);
nor U218 (N_218,In_172,In_445);
nor U219 (N_219,In_971,In_1186);
nand U220 (N_220,In_144,In_854);
or U221 (N_221,N_192,N_131);
nor U222 (N_222,In_127,N_146);
nand U223 (N_223,N_199,In_1185);
and U224 (N_224,In_98,In_1178);
and U225 (N_225,N_60,In_1181);
nand U226 (N_226,In_1356,In_1272);
nor U227 (N_227,In_1244,In_425);
nand U228 (N_228,In_842,In_367);
xor U229 (N_229,In_1054,In_264);
nand U230 (N_230,In_194,In_666);
and U231 (N_231,In_1229,In_42);
or U232 (N_232,In_1454,In_479);
or U233 (N_233,N_124,N_92);
nor U234 (N_234,In_307,In_329);
nor U235 (N_235,In_979,In_422);
nor U236 (N_236,In_877,In_311);
nor U237 (N_237,In_24,In_237);
or U238 (N_238,N_73,In_569);
nor U239 (N_239,In_72,In_736);
nand U240 (N_240,In_1011,In_115);
and U241 (N_241,In_299,In_121);
nor U242 (N_242,N_174,In_402);
and U243 (N_243,N_104,In_542);
or U244 (N_244,N_62,In_1463);
nor U245 (N_245,In_1168,In_188);
and U246 (N_246,In_43,In_880);
and U247 (N_247,In_208,In_899);
xnor U248 (N_248,In_276,In_1318);
nor U249 (N_249,In_911,In_184);
and U250 (N_250,In_417,N_143);
nor U251 (N_251,In_1239,In_1097);
nor U252 (N_252,In_757,In_1488);
nand U253 (N_253,In_781,In_857);
nor U254 (N_254,In_763,In_206);
nor U255 (N_255,In_1491,N_19);
and U256 (N_256,In_1088,In_6);
xnor U257 (N_257,In_14,In_460);
and U258 (N_258,In_884,In_1495);
or U259 (N_259,In_641,N_153);
nor U260 (N_260,In_1203,In_224);
xor U261 (N_261,In_1403,In_151);
nor U262 (N_262,In_190,In_3);
or U263 (N_263,In_1208,In_1278);
xor U264 (N_264,In_1338,In_544);
nand U265 (N_265,In_1439,In_929);
xor U266 (N_266,In_250,N_89);
xor U267 (N_267,In_142,In_1409);
nand U268 (N_268,In_925,In_1205);
nor U269 (N_269,N_12,N_110);
and U270 (N_270,In_676,In_107);
and U271 (N_271,In_983,N_168);
and U272 (N_272,In_273,In_286);
or U273 (N_273,N_108,In_138);
nor U274 (N_274,In_663,N_158);
nand U275 (N_275,In_12,In_563);
or U276 (N_276,In_1473,In_52);
nand U277 (N_277,In_368,In_730);
or U278 (N_278,In_137,In_678);
nand U279 (N_279,N_49,In_992);
and U280 (N_280,In_780,In_1441);
xor U281 (N_281,N_101,In_668);
xor U282 (N_282,N_95,In_1169);
xnor U283 (N_283,In_1248,In_832);
and U284 (N_284,In_116,In_962);
nor U285 (N_285,In_1109,In_697);
nand U286 (N_286,In_1147,In_1415);
nor U287 (N_287,In_775,N_32);
and U288 (N_288,In_1027,N_186);
nor U289 (N_289,In_886,In_967);
and U290 (N_290,N_145,In_517);
nor U291 (N_291,In_935,In_222);
or U292 (N_292,In_363,In_748);
nand U293 (N_293,N_44,In_1107);
nor U294 (N_294,In_1238,In_1417);
and U295 (N_295,In_1077,In_906);
nand U296 (N_296,In_1449,In_1440);
nor U297 (N_297,In_557,In_436);
xor U298 (N_298,In_1194,In_1141);
xor U299 (N_299,In_258,In_118);
nor U300 (N_300,In_205,In_664);
or U301 (N_301,In_1483,In_636);
or U302 (N_302,N_169,In_1151);
nand U303 (N_303,In_551,In_470);
and U304 (N_304,In_823,In_1261);
or U305 (N_305,N_121,In_692);
and U306 (N_306,N_105,N_34);
xor U307 (N_307,In_431,In_396);
nand U308 (N_308,In_622,In_742);
xnor U309 (N_309,In_487,In_978);
and U310 (N_310,In_1461,In_1350);
and U311 (N_311,In_198,In_332);
nand U312 (N_312,In_936,In_37);
and U313 (N_313,In_277,In_1422);
nor U314 (N_314,N_82,In_803);
or U315 (N_315,In_963,In_694);
nand U316 (N_316,In_1184,In_26);
nand U317 (N_317,N_116,In_915);
xor U318 (N_318,In_443,In_1124);
nor U319 (N_319,In_609,In_1198);
nor U320 (N_320,In_180,In_270);
or U321 (N_321,In_996,In_1362);
nand U322 (N_322,N_144,In_1104);
xnor U323 (N_323,In_738,In_623);
nor U324 (N_324,In_1007,In_933);
nand U325 (N_325,In_728,In_166);
nor U326 (N_326,In_475,In_68);
nand U327 (N_327,In_562,In_95);
nor U328 (N_328,N_136,In_648);
nand U329 (N_329,In_1258,N_0);
nor U330 (N_330,In_288,In_1496);
nor U331 (N_331,In_1348,In_243);
nor U332 (N_332,In_558,In_556);
nand U333 (N_333,In_889,In_856);
or U334 (N_334,In_1399,In_630);
xnor U335 (N_335,In_942,In_1311);
nand U336 (N_336,In_1084,N_28);
and U337 (N_337,In_146,In_245);
xor U338 (N_338,In_302,In_335);
or U339 (N_339,In_718,In_855);
or U340 (N_340,In_1347,In_512);
or U341 (N_341,In_838,In_448);
xnor U342 (N_342,In_231,In_1412);
and U343 (N_343,In_539,In_153);
or U344 (N_344,In_261,In_1060);
nor U345 (N_345,In_1270,In_696);
nand U346 (N_346,In_870,In_1451);
or U347 (N_347,In_914,In_530);
nand U348 (N_348,In_1140,N_152);
xnor U349 (N_349,In_1305,In_1288);
and U350 (N_350,In_33,In_703);
and U351 (N_351,In_1423,In_1016);
nor U352 (N_352,In_560,N_165);
nor U353 (N_353,In_579,In_41);
xnor U354 (N_354,N_179,In_209);
xnor U355 (N_355,In_1317,In_700);
or U356 (N_356,In_89,N_5);
nand U357 (N_357,N_69,In_1207);
xnor U358 (N_358,In_1132,In_1174);
and U359 (N_359,In_524,N_118);
nand U360 (N_360,In_40,In_109);
nand U361 (N_361,In_533,In_44);
or U362 (N_362,N_147,In_919);
xnor U363 (N_363,In_1342,In_743);
xor U364 (N_364,In_418,In_1455);
nand U365 (N_365,In_1286,In_650);
or U366 (N_366,In_5,In_428);
nor U367 (N_367,In_900,In_152);
and U368 (N_368,In_1253,In_410);
xor U369 (N_369,In_1091,N_24);
and U370 (N_370,In_616,In_1414);
xor U371 (N_371,N_6,In_950);
or U372 (N_372,In_1071,In_555);
nor U373 (N_373,In_1105,In_691);
nor U374 (N_374,In_369,N_188);
nand U375 (N_375,In_671,In_1432);
xor U376 (N_376,In_296,In_685);
nor U377 (N_377,In_581,In_375);
xor U378 (N_378,In_859,In_148);
and U379 (N_379,In_1413,In_714);
or U380 (N_380,In_343,In_429);
xnor U381 (N_381,In_974,In_806);
and U382 (N_382,In_966,In_1232);
nand U383 (N_383,In_1206,In_822);
nand U384 (N_384,In_1192,In_985);
nand U385 (N_385,In_546,N_162);
or U386 (N_386,In_106,N_177);
nand U387 (N_387,In_229,In_515);
and U388 (N_388,In_314,In_1085);
and U389 (N_389,In_380,In_617);
or U390 (N_390,In_644,In_480);
or U391 (N_391,In_310,In_831);
xor U392 (N_392,In_139,In_265);
nand U393 (N_393,N_81,In_341);
and U394 (N_394,In_789,In_371);
nand U395 (N_395,In_930,In_509);
and U396 (N_396,In_1274,In_982);
or U397 (N_397,In_1471,In_1405);
xor U398 (N_398,In_340,In_330);
and U399 (N_399,In_173,In_1388);
or U400 (N_400,In_642,N_9);
or U401 (N_401,In_112,In_708);
xor U402 (N_402,In_578,In_917);
and U403 (N_403,N_54,N_21);
and U404 (N_404,In_774,In_1223);
or U405 (N_405,In_705,N_18);
or U406 (N_406,In_879,In_1304);
nand U407 (N_407,N_324,N_337);
nor U408 (N_408,N_3,In_357);
xor U409 (N_409,In_656,In_1246);
and U410 (N_410,In_862,In_1352);
nor U411 (N_411,In_990,In_1457);
xor U412 (N_412,In_201,In_596);
nor U413 (N_413,In_1426,In_392);
xor U414 (N_414,In_246,In_215);
or U415 (N_415,In_51,N_27);
xnor U416 (N_416,N_290,In_1326);
xor U417 (N_417,In_511,In_455);
nor U418 (N_418,N_134,In_1324);
nor U419 (N_419,In_119,In_334);
xnor U420 (N_420,N_138,In_1083);
nand U421 (N_421,In_808,In_717);
xor U422 (N_422,N_237,N_182);
nand U423 (N_423,N_323,In_729);
xnor U424 (N_424,In_945,N_83);
and U425 (N_425,In_18,In_1195);
nand U426 (N_426,N_245,In_750);
and U427 (N_427,In_1182,In_841);
xor U428 (N_428,N_71,In_469);
nand U429 (N_429,In_525,N_266);
nor U430 (N_430,In_1012,In_85);
and U431 (N_431,N_240,In_1155);
and U432 (N_432,In_771,N_265);
nor U433 (N_433,N_270,In_1081);
nand U434 (N_434,In_816,In_233);
nand U435 (N_435,N_201,In_440);
nand U436 (N_436,In_136,In_1166);
xor U437 (N_437,N_50,In_1117);
and U438 (N_438,In_1265,N_282);
or U439 (N_439,In_813,In_1467);
or U440 (N_440,In_416,In_154);
nand U441 (N_441,In_1383,In_767);
or U442 (N_442,In_584,In_452);
nor U443 (N_443,In_955,In_1123);
nand U444 (N_444,In_941,N_271);
and U445 (N_445,N_261,In_362);
xnor U446 (N_446,N_149,In_366);
and U447 (N_447,N_200,In_810);
nor U448 (N_448,N_132,In_167);
and U449 (N_449,N_37,N_313);
or U450 (N_450,In_1277,In_20);
and U451 (N_451,In_171,In_580);
nand U452 (N_452,In_406,N_59);
nand U453 (N_453,N_58,In_704);
and U454 (N_454,N_164,In_133);
and U455 (N_455,In_909,N_161);
xnor U456 (N_456,In_407,In_140);
xor U457 (N_457,In_1173,In_1301);
nand U458 (N_458,N_243,In_706);
nand U459 (N_459,N_51,In_1118);
or U460 (N_460,In_1365,In_1120);
nor U461 (N_461,N_269,In_381);
xor U462 (N_462,In_689,In_1222);
and U463 (N_463,In_401,In_1251);
nor U464 (N_464,In_922,In_1064);
nand U465 (N_465,In_520,N_254);
and U466 (N_466,In_386,In_1281);
nor U467 (N_467,In_483,N_234);
nand U468 (N_468,In_759,In_272);
nor U469 (N_469,N_388,N_112);
nor U470 (N_470,In_496,N_343);
xor U471 (N_471,In_1072,N_310);
nand U472 (N_472,N_20,In_1416);
and U473 (N_473,In_913,In_1419);
or U474 (N_474,In_1033,In_328);
nor U475 (N_475,In_1082,In_1065);
xor U476 (N_476,N_311,In_494);
or U477 (N_477,N_255,In_160);
and U478 (N_478,In_484,N_85);
or U479 (N_479,In_69,In_315);
xor U480 (N_480,In_575,In_131);
xor U481 (N_481,In_744,N_396);
nand U482 (N_482,In_1247,In_820);
nor U483 (N_483,In_301,In_1468);
xnor U484 (N_484,In_1001,In_559);
and U485 (N_485,In_833,In_1443);
or U486 (N_486,In_667,In_902);
and U487 (N_487,In_16,In_1099);
xnor U488 (N_488,In_1219,N_372);
and U489 (N_489,In_566,In_176);
nor U490 (N_490,In_1313,N_26);
or U491 (N_491,In_1335,N_142);
xnor U492 (N_492,In_868,In_897);
nand U493 (N_493,In_227,N_52);
xor U494 (N_494,In_1349,N_231);
nor U495 (N_495,N_305,N_206);
or U496 (N_496,In_492,In_536);
or U497 (N_497,In_365,In_1329);
nor U498 (N_498,In_645,N_249);
nor U499 (N_499,N_68,In_465);
xor U500 (N_500,N_383,In_1255);
nand U501 (N_501,In_1386,In_1070);
nor U502 (N_502,N_111,In_389);
nor U503 (N_503,N_214,In_606);
or U504 (N_504,In_861,N_98);
xnor U505 (N_505,In_244,In_1370);
or U506 (N_506,In_248,N_267);
and U507 (N_507,In_1017,N_326);
nand U508 (N_508,In_903,In_1357);
or U509 (N_509,N_96,In_799);
or U510 (N_510,In_478,N_197);
or U511 (N_511,N_157,In_427);
or U512 (N_512,In_1400,N_43);
nor U513 (N_513,In_514,In_768);
and U514 (N_514,In_779,In_655);
nor U515 (N_515,N_233,In_1372);
or U516 (N_516,N_256,In_450);
nor U517 (N_517,N_262,In_267);
nand U518 (N_518,In_837,In_769);
and U519 (N_519,In_170,In_735);
nand U520 (N_520,In_393,N_222);
nor U521 (N_521,In_883,In_690);
nand U522 (N_522,In_266,N_203);
nor U523 (N_523,In_999,In_1193);
nand U524 (N_524,In_1381,In_1221);
nand U525 (N_525,In_521,In_1287);
xnor U526 (N_526,In_1498,In_888);
xnor U527 (N_527,N_353,In_104);
and U528 (N_528,In_523,In_1022);
nand U529 (N_529,In_1428,In_1481);
and U530 (N_530,In_576,In_1008);
nor U531 (N_531,N_338,In_1157);
and U532 (N_532,N_97,N_373);
or U533 (N_533,In_716,N_22);
and U534 (N_534,N_318,In_413);
xnor U535 (N_535,In_388,In_995);
nand U536 (N_536,In_65,In_683);
xor U537 (N_537,N_347,In_1122);
and U538 (N_538,N_72,In_956);
nand U539 (N_539,In_863,In_583);
xor U540 (N_540,N_286,In_669);
or U541 (N_541,In_1310,In_998);
xnor U542 (N_542,In_693,N_309);
and U543 (N_543,N_185,In_241);
nor U544 (N_544,In_1242,In_269);
or U545 (N_545,In_1284,In_196);
xnor U546 (N_546,In_1358,In_638);
nor U547 (N_547,In_1465,N_377);
and U548 (N_548,N_258,N_301);
or U549 (N_549,In_657,In_391);
xnor U550 (N_550,In_1115,N_380);
xnor U551 (N_551,N_1,In_238);
xor U552 (N_552,N_14,In_49);
nand U553 (N_553,In_226,N_321);
or U554 (N_554,N_292,N_368);
xor U555 (N_555,In_908,N_4);
xnor U556 (N_556,In_280,In_1361);
xnor U557 (N_557,In_1291,N_327);
nand U558 (N_558,N_181,N_35);
and U559 (N_559,In_1189,N_322);
xnor U560 (N_560,In_1300,N_355);
nand U561 (N_561,In_1408,N_88);
xor U562 (N_562,N_342,In_552);
and U563 (N_563,N_103,In_1249);
or U564 (N_564,In_232,N_187);
xor U565 (N_565,N_70,N_226);
nand U566 (N_566,In_463,In_1374);
or U567 (N_567,N_160,In_1103);
and U568 (N_568,In_845,In_74);
nor U569 (N_569,In_351,In_626);
or U570 (N_570,In_80,In_61);
nor U571 (N_571,In_1111,In_846);
xnor U572 (N_572,In_303,N_167);
nor U573 (N_573,N_125,In_203);
or U574 (N_574,In_1407,N_374);
xor U575 (N_575,In_490,In_1353);
nor U576 (N_576,N_213,N_2);
or U577 (N_577,In_1163,In_235);
nor U578 (N_578,In_1376,N_384);
nand U579 (N_579,N_340,In_1204);
nand U580 (N_580,In_195,In_890);
xnor U581 (N_581,In_390,In_1391);
nand U582 (N_582,In_1220,N_320);
or U583 (N_583,N_196,N_253);
and U584 (N_584,N_223,In_17);
nand U585 (N_585,In_627,In_108);
nand U586 (N_586,In_1447,In_762);
nand U587 (N_587,In_740,N_91);
nand U588 (N_588,In_847,In_1297);
or U589 (N_589,In_745,In_1183);
or U590 (N_590,N_225,In_980);
or U591 (N_591,N_329,In_76);
xor U592 (N_592,In_991,N_178);
xnor U593 (N_593,N_180,In_81);
nand U594 (N_594,In_1337,In_784);
and U595 (N_595,In_710,In_1369);
nor U596 (N_596,In_643,In_1004);
or U597 (N_597,N_242,N_260);
and U598 (N_598,N_140,In_1149);
or U599 (N_599,In_474,In_200);
nor U600 (N_600,In_749,In_83);
xnor U601 (N_601,In_844,N_529);
nor U602 (N_602,In_1024,In_1228);
and U603 (N_603,In_1243,In_8);
xor U604 (N_604,N_598,N_278);
xor U605 (N_605,In_477,In_488);
nand U606 (N_606,In_1257,In_185);
nand U607 (N_607,In_353,N_288);
or U608 (N_608,N_519,N_314);
nand U609 (N_609,In_654,N_40);
and U610 (N_610,In_565,In_395);
nor U611 (N_611,In_553,N_545);
nor U612 (N_612,N_436,In_592);
nand U613 (N_613,N_367,In_25);
nor U614 (N_614,In_1340,In_1285);
nand U615 (N_615,N_339,In_1131);
and U616 (N_616,N_421,N_360);
nand U617 (N_617,In_113,N_407);
or U618 (N_618,In_1336,N_137);
or U619 (N_619,In_529,N_486);
and U620 (N_620,N_586,In_1010);
and U621 (N_621,N_190,N_516);
or U622 (N_622,In_599,N_594);
nand U623 (N_623,In_611,In_75);
and U624 (N_624,N_280,N_16);
or U625 (N_625,In_421,N_235);
xnor U626 (N_626,N_572,N_219);
xnor U627 (N_627,N_47,N_361);
or U628 (N_628,In_795,In_964);
nor U629 (N_629,In_325,In_649);
xor U630 (N_630,N_564,In_1235);
nand U631 (N_631,In_32,N_293);
or U632 (N_632,In_1303,In_739);
nor U633 (N_633,N_472,N_533);
nand U634 (N_634,In_1028,In_1048);
nand U635 (N_635,In_1015,In_1025);
nand U636 (N_636,In_283,In_1217);
nor U637 (N_637,N_395,In_528);
nand U638 (N_638,N_335,In_849);
and U639 (N_639,N_438,N_284);
nor U640 (N_640,N_535,In_1367);
or U641 (N_641,In_15,In_1101);
nand U642 (N_642,In_571,In_1153);
nor U643 (N_643,In_57,N_205);
nor U644 (N_644,N_263,In_726);
nor U645 (N_645,N_193,In_732);
xor U646 (N_646,N_163,N_129);
nand U647 (N_647,In_1113,N_102);
and U648 (N_648,N_107,In_161);
xor U649 (N_649,In_741,In_225);
or U650 (N_650,In_1133,In_526);
nand U651 (N_651,N_238,In_1036);
xor U652 (N_652,In_1368,In_651);
nand U653 (N_653,N_366,In_1002);
and U654 (N_654,In_336,In_947);
and U655 (N_655,In_459,N_549);
and U656 (N_656,In_59,N_349);
or U657 (N_657,N_114,In_724);
or U658 (N_658,N_487,In_1493);
or U659 (N_659,In_840,N_430);
nand U660 (N_660,In_686,In_1092);
xor U661 (N_661,In_1066,In_519);
or U662 (N_662,In_1013,In_177);
nand U663 (N_663,In_253,In_481);
nor U664 (N_664,N_76,In_1321);
nor U665 (N_665,N_381,N_582);
xnor U666 (N_666,In_23,In_1146);
nor U667 (N_667,In_155,N_408);
or U668 (N_668,In_86,In_1325);
and U669 (N_669,N_419,In_1038);
xor U670 (N_670,N_527,N_556);
and U671 (N_671,In_439,In_1487);
nand U672 (N_672,In_506,N_36);
and U673 (N_673,In_1273,N_589);
or U674 (N_674,In_399,N_466);
and U675 (N_675,In_92,N_25);
nand U676 (N_676,In_652,N_402);
and U677 (N_677,In_165,N_8);
xor U678 (N_678,In_1233,In_1359);
or U679 (N_679,In_1271,N_446);
and U680 (N_680,In_192,N_139);
and U681 (N_681,N_7,In_240);
nor U682 (N_682,In_1334,In_865);
or U683 (N_683,In_1460,In_1424);
or U684 (N_684,N_457,N_227);
or U685 (N_685,In_819,N_211);
xnor U686 (N_686,In_687,N_176);
nand U687 (N_687,N_420,N_120);
nor U688 (N_688,N_413,N_538);
nor U689 (N_689,In_316,N_294);
nand U690 (N_690,In_493,In_1100);
nor U691 (N_691,N_357,N_584);
and U692 (N_692,In_826,In_1043);
nor U693 (N_693,In_635,N_554);
and U694 (N_694,N_449,N_364);
nand U695 (N_695,In_965,In_141);
nand U696 (N_696,In_376,N_371);
nand U697 (N_697,In_419,In_344);
nand U698 (N_698,N_128,N_515);
xnor U699 (N_699,N_78,N_378);
xor U700 (N_700,In_1200,In_1499);
or U701 (N_701,N_48,In_187);
and U702 (N_702,In_910,In_1127);
or U703 (N_703,N_306,N_405);
and U704 (N_704,In_228,N_481);
nor U705 (N_705,In_1446,In_1052);
nand U706 (N_706,N_518,In_55);
nand U707 (N_707,In_1466,N_454);
nor U708 (N_708,N_100,N_414);
nand U709 (N_709,In_1089,N_325);
or U710 (N_710,In_615,N_450);
nand U711 (N_711,N_218,In_776);
nand U712 (N_712,In_374,N_39);
or U713 (N_713,N_148,In_712);
xnor U714 (N_714,In_21,In_1034);
or U715 (N_715,In_1393,N_422);
xnor U716 (N_716,In_279,In_755);
nand U717 (N_717,In_230,In_821);
nor U718 (N_718,N_590,In_1402);
nor U719 (N_719,In_1450,In_568);
nand U720 (N_720,In_1259,In_825);
nand U721 (N_721,In_1492,In_723);
nor U722 (N_722,In_124,N_259);
and U723 (N_723,In_359,N_184);
or U724 (N_724,In_1053,In_202);
xor U725 (N_725,In_924,In_101);
and U726 (N_726,N_415,N_296);
nand U727 (N_727,N_501,In_1075);
xnor U728 (N_728,N_424,N_379);
nand U729 (N_729,In_430,N_389);
xnor U730 (N_730,N_455,In_594);
nor U731 (N_731,N_251,N_38);
xor U732 (N_732,In_698,In_1179);
and U733 (N_733,N_308,In_860);
or U734 (N_734,N_532,N_246);
and U735 (N_735,In_1260,In_1430);
nand U736 (N_736,N_574,In_661);
xor U737 (N_737,In_60,N_510);
nand U738 (N_738,In_835,N_488);
nand U739 (N_739,N_106,In_1331);
and U740 (N_740,N_585,In_923);
xor U741 (N_741,N_561,N_536);
xnor U742 (N_742,N_31,N_207);
and U743 (N_743,N_534,In_1135);
xor U744 (N_744,In_1351,In_1245);
xor U745 (N_745,In_1139,In_327);
xnor U746 (N_746,In_502,In_751);
or U747 (N_747,N_403,N_540);
nand U748 (N_748,In_50,In_785);
nand U749 (N_749,In_306,N_587);
nand U750 (N_750,N_478,In_954);
or U751 (N_751,In_295,N_588);
and U752 (N_752,In_574,N_273);
nor U753 (N_753,In_90,N_485);
xnor U754 (N_754,In_2,In_1292);
and U755 (N_755,N_416,In_639);
and U756 (N_756,N_241,N_495);
or U757 (N_757,N_567,In_473);
nor U758 (N_758,N_558,In_46);
xnor U759 (N_759,N_470,In_48);
and U760 (N_760,N_441,In_1177);
or U761 (N_761,In_792,In_1187);
and U762 (N_762,N_435,In_1112);
xor U763 (N_763,N_239,In_817);
or U764 (N_764,N_489,In_159);
and U765 (N_765,In_1442,In_64);
and U766 (N_766,N_400,In_1130);
nand U767 (N_767,In_1079,In_1437);
nand U768 (N_768,N_189,In_1175);
nor U769 (N_769,N_382,In_1475);
or U770 (N_770,In_39,N_370);
and U771 (N_771,N_580,N_392);
nor U772 (N_772,In_204,N_456);
xor U773 (N_773,In_1234,N_555);
nor U774 (N_774,In_379,In_1485);
xor U775 (N_775,In_895,In_772);
or U776 (N_776,N_352,N_596);
and U777 (N_777,In_773,In_298);
and U778 (N_778,N_597,In_1029);
nor U779 (N_779,N_477,N_546);
nand U780 (N_780,N_406,In_163);
xnor U781 (N_781,N_99,In_1055);
xnor U782 (N_782,N_559,In_543);
nand U783 (N_783,N_443,N_291);
xor U784 (N_784,N_442,N_217);
and U785 (N_785,In_1076,In_1290);
xor U786 (N_786,In_1264,N_247);
nor U787 (N_787,In_313,N_453);
xor U788 (N_788,N_198,In_548);
and U789 (N_789,In_796,In_434);
or U790 (N_790,In_218,N_537);
nand U791 (N_791,N_498,In_912);
or U792 (N_792,In_1236,In_319);
nor U793 (N_793,In_56,In_713);
and U794 (N_794,In_308,In_928);
xor U795 (N_795,In_1302,N_363);
or U796 (N_796,In_986,In_1021);
nand U797 (N_797,In_1094,N_551);
nor U798 (N_798,In_984,In_1378);
xnor U799 (N_799,In_1108,In_438);
nand U800 (N_800,In_1150,In_361);
nand U801 (N_801,N_687,N_499);
nor U802 (N_802,N_668,N_647);
nor U803 (N_803,N_746,N_53);
nand U804 (N_804,N_600,N_754);
nand U805 (N_805,N_665,N_728);
xor U806 (N_806,N_528,In_510);
or U807 (N_807,N_41,N_530);
and U808 (N_808,N_621,In_132);
nor U809 (N_809,N_571,In_927);
or U810 (N_810,In_333,N_785);
nor U811 (N_811,N_606,N_725);
nand U812 (N_812,N_733,N_252);
nor U813 (N_813,N_445,N_622);
and U814 (N_814,N_741,N_663);
nand U815 (N_815,In_321,In_400);
and U816 (N_816,In_291,In_337);
and U817 (N_817,N_394,In_282);
or U818 (N_818,N_113,N_671);
and U819 (N_819,N_658,N_299);
xor U820 (N_820,N_742,N_609);
and U821 (N_821,N_281,N_715);
nand U822 (N_822,In_364,In_212);
xor U823 (N_823,N_509,N_399);
xnor U824 (N_824,In_67,N_640);
nand U825 (N_825,N_710,N_473);
nand U826 (N_826,In_1341,N_729);
nor U827 (N_827,N_738,N_636);
or U828 (N_828,N_151,N_482);
and U829 (N_829,N_602,N_504);
xnor U830 (N_830,N_159,N_15);
or U831 (N_831,In_252,In_582);
xnor U832 (N_832,N_707,In_442);
nand U833 (N_833,In_1394,N_776);
xnor U834 (N_834,N_719,N_618);
and U835 (N_835,In_271,In_255);
and U836 (N_836,In_1279,In_453);
and U837 (N_837,In_1073,N_216);
and U838 (N_838,N_714,N_468);
nor U839 (N_839,In_1307,In_377);
and U840 (N_840,In_1448,In_680);
nand U841 (N_841,In_1224,N_641);
or U842 (N_842,N_358,N_632);
xor U843 (N_843,N_65,N_474);
nand U844 (N_844,N_577,In_1397);
or U845 (N_845,N_362,N_397);
or U846 (N_846,N_751,N_657);
nor U847 (N_847,In_507,In_1275);
xnor U848 (N_848,N_334,N_475);
nand U849 (N_849,N_737,N_300);
nand U850 (N_850,N_215,In_260);
and U851 (N_851,In_1191,N_463);
or U852 (N_852,N_744,N_557);
nand U853 (N_853,N_11,N_459);
nand U854 (N_854,In_637,N_297);
or U855 (N_855,N_434,N_345);
or U856 (N_856,N_55,N_722);
nor U857 (N_857,In_585,In_747);
nand U858 (N_858,In_695,N_760);
and U859 (N_859,In_848,In_1063);
or U860 (N_860,N_541,N_717);
nand U861 (N_861,N_194,N_635);
xor U862 (N_862,In_1333,In_394);
or U863 (N_863,N_461,N_749);
nand U864 (N_864,In_1014,N_79);
nand U865 (N_865,In_625,N_702);
or U866 (N_866,In_873,N_705);
xor U867 (N_867,In_397,In_1106);
nor U868 (N_868,N_669,N_786);
nor U869 (N_869,N_758,N_505);
xor U870 (N_870,N_766,In_1294);
nand U871 (N_871,In_143,N_526);
nand U872 (N_872,In_126,In_1128);
nor U873 (N_873,N_748,N_779);
and U874 (N_874,N_56,N_631);
nand U875 (N_875,N_683,N_109);
and U876 (N_876,N_730,In_1256);
or U877 (N_877,N_667,N_328);
xor U878 (N_878,N_244,N_204);
nor U879 (N_879,In_1037,N_645);
xor U880 (N_880,In_793,N_797);
xnor U881 (N_881,N_30,In_1196);
or U882 (N_882,In_1280,N_709);
and U883 (N_883,N_675,In_77);
and U884 (N_884,N_115,N_656);
nor U885 (N_885,N_173,N_117);
nand U886 (N_886,N_490,N_661);
and U887 (N_887,In_1041,N_517);
nand U888 (N_888,N_581,In_737);
nor U889 (N_889,In_1406,In_221);
xnor U890 (N_890,In_263,N_316);
nand U891 (N_891,N_319,N_458);
nor U892 (N_892,N_697,In_1458);
nand U893 (N_893,N_789,In_1344);
xnor U894 (N_894,N_773,In_867);
and U895 (N_895,N_792,In_1309);
or U896 (N_896,N_156,In_814);
nor U897 (N_897,N_700,N_727);
and U898 (N_898,N_639,In_1067);
nor U899 (N_899,N_756,In_207);
xor U900 (N_900,In_538,N_778);
and U901 (N_901,N_494,N_212);
or U902 (N_902,In_989,N_695);
and U903 (N_903,N_230,N_791);
nor U904 (N_904,N_611,N_757);
nor U905 (N_905,In_1059,In_322);
xnor U906 (N_906,N_502,In_787);
xor U907 (N_907,In_805,In_182);
or U908 (N_908,In_284,N_761);
and U909 (N_909,N_573,N_404);
nand U910 (N_910,N_330,N_716);
nand U911 (N_911,In_1377,In_466);
and U912 (N_912,In_247,N_795);
and U913 (N_913,In_1395,N_283);
xnor U914 (N_914,N_670,In_145);
nor U915 (N_915,N_607,N_649);
xnor U916 (N_916,In_591,In_1170);
and U917 (N_917,N_677,In_537);
and U918 (N_918,In_567,N_692);
or U919 (N_919,In_684,N_209);
and U920 (N_920,N_550,In_607);
or U921 (N_921,N_782,In_613);
nor U922 (N_922,N_794,In_1371);
nor U923 (N_923,N_511,N_664);
xnor U924 (N_924,N_604,N_257);
xnor U925 (N_925,N_33,N_620);
or U926 (N_926,N_491,N_775);
nor U927 (N_927,In_408,In_1058);
xor U928 (N_928,N_629,N_42);
nor U929 (N_929,N_274,In_1296);
or U930 (N_930,In_1379,In_619);
xnor U931 (N_931,In_499,N_601);
or U932 (N_932,N_603,N_799);
and U933 (N_933,N_617,In_30);
xor U934 (N_934,N_390,In_672);
or U935 (N_935,N_229,In_918);
nand U936 (N_936,N_183,N_150);
nor U937 (N_937,In_1042,N_745);
and U938 (N_938,N_220,In_96);
nand U939 (N_939,N_90,N_264);
nand U940 (N_940,N_248,N_712);
nor U941 (N_941,N_506,N_548);
and U942 (N_942,N_565,In_679);
nand U943 (N_943,N_614,N_731);
nand U944 (N_944,N_578,N_460);
nand U945 (N_945,In_1000,N_503);
xor U946 (N_946,N_627,N_576);
nor U947 (N_947,N_788,N_287);
and U948 (N_948,N_769,N_593);
nand U949 (N_949,In_610,In_725);
nand U950 (N_950,In_731,N_525);
and U951 (N_951,N_643,N_170);
and U952 (N_952,N_331,N_250);
nand U953 (N_953,N_615,In_1216);
nand U954 (N_954,In_508,N_750);
and U955 (N_955,N_171,N_202);
nor U956 (N_956,In_93,N_762);
nand U957 (N_957,N_625,N_542);
and U958 (N_958,N_720,N_539);
nor U959 (N_959,In_754,N_483);
or U960 (N_960,In_1061,N_398);
or U961 (N_961,N_678,In_633);
nand U962 (N_962,N_610,N_753);
or U963 (N_963,N_385,In_629);
or U964 (N_964,In_1315,N_94);
or U965 (N_965,N_341,N_172);
xnor U966 (N_966,N_210,N_130);
nand U967 (N_967,N_568,In_1489);
and U968 (N_968,N_61,N_547);
nand U969 (N_969,In_456,N_492);
xor U970 (N_970,N_662,N_409);
and U971 (N_971,N_566,N_583);
and U972 (N_972,N_723,N_608);
xor U973 (N_973,In_1425,In_603);
xor U974 (N_974,In_675,N_452);
nand U975 (N_975,N_426,N_484);
or U976 (N_976,N_767,N_275);
and U977 (N_977,N_480,N_798);
or U978 (N_978,N_23,N_524);
or U979 (N_979,N_694,N_191);
and U980 (N_980,N_646,N_401);
and U981 (N_981,In_953,N_685);
xnor U982 (N_982,In_824,N_628);
xor U983 (N_983,In_564,In_441);
nor U984 (N_984,In_1134,N_612);
and U985 (N_985,In_541,N_29);
xnor U986 (N_986,N_122,In_1438);
nor U987 (N_987,N_513,N_302);
and U988 (N_988,N_298,N_690);
nand U989 (N_989,In_482,N_351);
or U990 (N_990,N_780,N_493);
or U991 (N_991,N_303,In_1026);
xnor U992 (N_992,N_682,N_763);
nor U993 (N_993,N_13,N_87);
nor U994 (N_994,N_653,In_423);
nand U995 (N_995,N_496,In_1293);
nand U996 (N_996,In_957,N_676);
nor U997 (N_997,N_706,In_186);
nand U998 (N_998,N_45,In_1209);
and U999 (N_999,N_784,N_332);
xnor U1000 (N_1000,N_701,N_651);
or U1001 (N_1001,In_1355,N_998);
xnor U1002 (N_1002,N_842,In_1039);
xnor U1003 (N_1003,N_734,N_279);
xnor U1004 (N_1004,N_881,N_221);
and U1005 (N_1005,N_476,N_166);
xnor U1006 (N_1006,N_801,In_905);
and U1007 (N_1007,N_500,In_1045);
and U1008 (N_1008,N_956,In_414);
or U1009 (N_1009,N_522,N_736);
nor U1010 (N_1010,In_471,N_977);
nand U1011 (N_1011,N_937,N_126);
xor U1012 (N_1012,N_819,N_864);
nand U1013 (N_1013,N_926,In_1410);
nor U1014 (N_1014,N_983,N_847);
and U1015 (N_1015,In_531,N_411);
xor U1016 (N_1016,N_289,N_155);
nor U1017 (N_1017,N_768,N_869);
nor U1018 (N_1018,N_354,N_807);
xnor U1019 (N_1019,N_947,N_972);
xor U1020 (N_1020,N_268,In_1472);
or U1021 (N_1021,N_830,N_994);
and U1022 (N_1022,N_884,N_790);
or U1023 (N_1023,In_304,N_285);
nand U1024 (N_1024,N_999,N_523);
nand U1025 (N_1025,N_681,N_895);
xor U1026 (N_1026,In_1162,N_135);
and U1027 (N_1027,N_666,N_858);
xnor U1028 (N_1028,N_448,N_344);
nor U1029 (N_1029,N_897,N_391);
or U1030 (N_1030,N_912,N_704);
xnor U1031 (N_1031,N_703,N_927);
and U1032 (N_1032,In_297,N_369);
nor U1033 (N_1033,N_992,N_119);
or U1034 (N_1034,N_560,N_975);
nand U1035 (N_1035,N_968,N_988);
nor U1036 (N_1036,N_879,N_521);
nor U1037 (N_1037,N_648,N_919);
or U1038 (N_1038,In_420,N_985);
xnor U1039 (N_1039,N_940,N_569);
xor U1040 (N_1040,In_29,N_127);
and U1041 (N_1041,In_120,N_948);
nand U1042 (N_1042,N_914,N_898);
nand U1043 (N_1043,N_154,In_323);
xor U1044 (N_1044,N_633,N_813);
and U1045 (N_1045,In_570,N_348);
or U1046 (N_1046,In_1215,N_644);
or U1047 (N_1047,N_553,In_1267);
and U1048 (N_1048,N_208,N_699);
or U1049 (N_1049,In_1420,N_837);
xor U1050 (N_1050,In_183,N_272);
and U1051 (N_1051,N_804,N_570);
and U1052 (N_1052,N_959,N_66);
and U1053 (N_1053,N_944,N_654);
nor U1054 (N_1054,N_915,N_777);
nand U1055 (N_1055,N_993,N_721);
nand U1056 (N_1056,N_356,N_508);
nand U1057 (N_1057,In_752,N_839);
or U1058 (N_1058,In_500,N_943);
nand U1059 (N_1059,N_925,In_476);
xnor U1060 (N_1060,N_507,N_979);
nand U1061 (N_1061,N_520,N_783);
and U1062 (N_1062,In_169,N_909);
or U1063 (N_1063,N_817,N_592);
nor U1064 (N_1064,N_806,N_899);
nor U1065 (N_1065,N_893,N_827);
xor U1066 (N_1066,N_921,N_659);
and U1067 (N_1067,In_123,In_97);
and U1068 (N_1068,N_851,N_970);
nor U1069 (N_1069,In_79,In_251);
nand U1070 (N_1070,N_859,In_464);
xor U1071 (N_1071,N_429,In_939);
and U1072 (N_1072,N_812,N_743);
and U1073 (N_1073,N_759,N_346);
or U1074 (N_1074,N_843,N_674);
nand U1075 (N_1075,N_923,N_307);
nor U1076 (N_1076,N_497,N_924);
nor U1077 (N_1077,In_1375,In_1308);
or U1078 (N_1078,N_63,N_809);
nand U1079 (N_1079,N_958,N_386);
nor U1080 (N_1080,N_902,N_978);
xor U1081 (N_1081,In_876,N_852);
nand U1082 (N_1082,In_1332,In_1074);
xnor U1083 (N_1083,N_563,N_444);
xnor U1084 (N_1084,N_650,N_825);
nand U1085 (N_1085,N_718,In_1086);
or U1086 (N_1086,In_812,N_818);
nor U1087 (N_1087,N_680,N_891);
nor U1088 (N_1088,N_512,N_991);
nand U1089 (N_1089,N_844,N_599);
xnor U1090 (N_1090,N_688,N_805);
and U1091 (N_1091,N_793,N_764);
nand U1092 (N_1092,N_984,In_211);
xor U1093 (N_1093,N_885,N_376);
nand U1094 (N_1094,In_783,N_315);
nor U1095 (N_1095,N_803,N_850);
xor U1096 (N_1096,N_630,N_829);
nand U1097 (N_1097,N_711,N_439);
nor U1098 (N_1098,In_561,N_930);
nor U1099 (N_1099,N_872,N_823);
or U1100 (N_1100,N_693,In_457);
and U1101 (N_1101,N_934,N_691);
xor U1102 (N_1102,In_598,In_383);
nand U1103 (N_1103,N_865,N_123);
xor U1104 (N_1104,N_552,N_920);
and U1105 (N_1105,In_1316,N_846);
nor U1106 (N_1106,In_620,N_822);
nand U1107 (N_1107,N_942,N_981);
xor U1108 (N_1108,N_946,N_74);
or U1109 (N_1109,N_966,In_1320);
nand U1110 (N_1110,N_228,N_660);
xnor U1111 (N_1111,N_359,N_894);
and U1112 (N_1112,N_955,N_892);
and U1113 (N_1113,N_824,N_689);
nor U1114 (N_1114,N_686,N_544);
and U1115 (N_1115,In_1345,N_365);
or U1116 (N_1116,N_996,N_579);
nor U1117 (N_1117,N_623,N_957);
and U1118 (N_1118,N_652,N_973);
nor U1119 (N_1119,N_479,In_577);
xnor U1120 (N_1120,In_818,In_612);
or U1121 (N_1121,N_619,N_841);
nand U1122 (N_1122,In_1354,N_605);
and U1123 (N_1123,N_916,N_232);
xnor U1124 (N_1124,N_740,N_431);
or U1125 (N_1125,N_708,N_437);
xor U1126 (N_1126,N_997,In_1392);
xor U1127 (N_1127,N_295,N_941);
or U1128 (N_1128,N_882,N_874);
nor U1129 (N_1129,N_857,N_856);
xor U1130 (N_1130,N_911,N_862);
and U1131 (N_1131,N_317,N_906);
nor U1132 (N_1132,N_735,N_875);
or U1133 (N_1133,N_989,N_928);
and U1134 (N_1134,N_938,N_333);
or U1135 (N_1135,N_808,N_967);
xor U1136 (N_1136,N_866,N_834);
or U1137 (N_1137,N_913,N_900);
nand U1138 (N_1138,In_1421,In_896);
and U1139 (N_1139,N_336,In_830);
nor U1140 (N_1140,N_873,N_853);
xnor U1141 (N_1141,N_613,N_861);
nand U1142 (N_1142,N_945,N_931);
and U1143 (N_1143,N_904,In_1102);
and U1144 (N_1144,N_575,N_964);
nor U1145 (N_1145,N_387,In_1387);
nor U1146 (N_1146,In_1212,N_418);
or U1147 (N_1147,In_1172,N_471);
nand U1148 (N_1148,N_917,In_262);
and U1149 (N_1149,N_713,N_860);
or U1150 (N_1150,In_665,N_672);
or U1151 (N_1151,N_276,N_908);
xor U1152 (N_1152,N_910,N_833);
nor U1153 (N_1153,In_318,N_637);
xor U1154 (N_1154,N_752,N_787);
nand U1155 (N_1155,N_965,N_86);
or U1156 (N_1156,N_412,In_409);
xor U1157 (N_1157,N_887,N_953);
nand U1158 (N_1158,N_929,N_642);
or U1159 (N_1159,In_1047,N_467);
xor U1160 (N_1160,N_831,N_918);
nand U1161 (N_1161,N_811,N_440);
nor U1162 (N_1162,N_781,In_348);
or U1163 (N_1163,N_75,N_821);
and U1164 (N_1164,N_684,In_372);
xor U1165 (N_1165,N_304,N_962);
xor U1166 (N_1166,In_347,N_935);
and U1167 (N_1167,N_739,N_698);
xnor U1168 (N_1168,N_939,In_1138);
xor U1169 (N_1169,N_655,In_1144);
nor U1170 (N_1170,N_433,N_17);
nor U1171 (N_1171,N_626,N_854);
or U1172 (N_1172,N_800,N_987);
xnor U1173 (N_1173,In_285,N_969);
and U1174 (N_1174,In_34,N_871);
xor U1175 (N_1175,N_747,In_952);
nand U1176 (N_1176,N_771,N_889);
and U1177 (N_1177,In_600,N_828);
xnor U1178 (N_1178,In_117,In_797);
nand U1179 (N_1179,In_872,N_469);
and U1180 (N_1180,N_949,N_673);
nand U1181 (N_1181,In_458,N_423);
or U1182 (N_1182,N_451,N_954);
nand U1183 (N_1183,In_807,N_432);
and U1184 (N_1184,N_393,N_732);
or U1185 (N_1185,N_427,N_543);
nand U1186 (N_1186,N_976,N_84);
xor U1187 (N_1187,N_755,In_350);
xor U1188 (N_1188,In_1171,N_465);
and U1189 (N_1189,N_638,N_133);
xor U1190 (N_1190,In_236,N_890);
and U1191 (N_1191,N_816,N_980);
and U1192 (N_1192,N_974,In_1019);
and U1193 (N_1193,N_634,N_447);
and U1194 (N_1194,N_462,N_849);
nor U1195 (N_1195,In_1434,N_770);
xor U1196 (N_1196,N_765,In_682);
or U1197 (N_1197,N_810,N_425);
nand U1198 (N_1198,In_535,N_375);
and U1199 (N_1199,N_312,N_616);
xnor U1200 (N_1200,N_1172,N_1041);
and U1201 (N_1201,N_1055,N_1132);
or U1202 (N_1202,N_995,N_1183);
xnor U1203 (N_1203,N_1077,N_836);
or U1204 (N_1204,N_1009,In_504);
nor U1205 (N_1205,N_1017,N_1150);
xor U1206 (N_1206,N_845,N_1130);
nand U1207 (N_1207,N_1060,N_1071);
or U1208 (N_1208,N_1065,In_699);
nand U1209 (N_1209,N_1152,In_1470);
and U1210 (N_1210,In_1,N_1053);
and U1211 (N_1211,N_832,N_1010);
and U1212 (N_1212,N_1040,N_1145);
and U1213 (N_1213,N_1194,N_1089);
or U1214 (N_1214,N_1054,N_1107);
xnor U1215 (N_1215,In_1482,N_1086);
or U1216 (N_1216,N_195,N_1104);
and U1217 (N_1217,N_1144,N_1101);
or U1218 (N_1218,N_1195,N_1005);
or U1219 (N_1219,N_1139,N_1118);
or U1220 (N_1220,N_1002,N_1154);
xor U1221 (N_1221,N_986,N_1022);
xnor U1222 (N_1222,N_961,N_1003);
xnor U1223 (N_1223,N_1033,N_726);
and U1224 (N_1224,N_840,N_1025);
nand U1225 (N_1225,N_1013,N_1142);
nand U1226 (N_1226,N_1133,N_870);
nand U1227 (N_1227,N_826,N_901);
nor U1228 (N_1228,N_595,N_1004);
and U1229 (N_1229,N_883,N_1109);
or U1230 (N_1230,N_10,N_1099);
or U1231 (N_1231,N_896,N_886);
nand U1232 (N_1232,N_1095,N_1131);
and U1233 (N_1233,N_428,N_64);
xor U1234 (N_1234,N_1184,N_1138);
nor U1235 (N_1235,N_1178,N_1090);
nor U1236 (N_1236,N_224,N_1128);
xor U1237 (N_1237,N_1157,N_1192);
nor U1238 (N_1238,N_1111,N_820);
nor U1239 (N_1239,N_1162,N_1064);
xnor U1240 (N_1240,N_1164,N_982);
and U1241 (N_1241,N_815,In_387);
xnor U1242 (N_1242,In_618,N_1076);
nand U1243 (N_1243,N_1043,N_1174);
xor U1244 (N_1244,N_1081,N_1011);
nor U1245 (N_1245,N_1069,N_835);
xor U1246 (N_1246,N_1180,N_1012);
and U1247 (N_1247,N_1082,N_1115);
xnor U1248 (N_1248,N_863,N_1050);
nor U1249 (N_1249,N_1102,N_1066);
nor U1250 (N_1250,N_1019,N_562);
nand U1251 (N_1251,N_46,N_1103);
or U1252 (N_1252,N_1035,N_1137);
nand U1253 (N_1253,N_1061,N_1148);
xnor U1254 (N_1254,N_1106,N_1116);
xnor U1255 (N_1255,In_1032,N_903);
or U1256 (N_1256,N_1015,N_1038);
or U1257 (N_1257,N_1188,N_1167);
nor U1258 (N_1258,N_1189,N_1143);
and U1259 (N_1259,In_105,N_1026);
xor U1260 (N_1260,N_1129,N_1023);
nand U1261 (N_1261,N_1155,N_1168);
nor U1262 (N_1262,N_932,N_1113);
nor U1263 (N_1263,In_28,N_1166);
or U1264 (N_1264,N_1074,N_1097);
and U1265 (N_1265,N_1039,N_1123);
and U1266 (N_1266,N_1190,N_1196);
and U1267 (N_1267,N_1117,N_867);
xnor U1268 (N_1268,N_1127,N_1193);
and U1269 (N_1269,N_1085,N_1126);
nor U1270 (N_1270,N_1000,N_1191);
nand U1271 (N_1271,N_796,N_77);
or U1272 (N_1272,N_1073,N_1059);
nor U1273 (N_1273,In_1049,N_1173);
and U1274 (N_1274,N_236,N_1087);
nand U1275 (N_1275,N_350,N_591);
xnor U1276 (N_1276,N_1018,N_1092);
nor U1277 (N_1277,N_1112,N_1119);
and U1278 (N_1278,N_696,N_1001);
and U1279 (N_1279,N_1031,N_1187);
nand U1280 (N_1280,N_1070,N_1068);
or U1281 (N_1281,N_963,N_1179);
nand U1282 (N_1282,N_936,N_1198);
or U1283 (N_1283,N_1042,N_1080);
nand U1284 (N_1284,N_774,N_1029);
nor U1285 (N_1285,N_1091,In_175);
nand U1286 (N_1286,N_1058,N_1125);
nor U1287 (N_1287,N_1176,N_1096);
xnor U1288 (N_1288,N_877,N_1110);
and U1289 (N_1289,N_971,N_1160);
nand U1290 (N_1290,N_679,N_1163);
nor U1291 (N_1291,N_1151,N_1141);
and U1292 (N_1292,N_1169,In_293);
nor U1293 (N_1293,In_1121,N_1149);
xor U1294 (N_1294,N_1120,N_1051);
and U1295 (N_1295,N_1052,N_1057);
nor U1296 (N_1296,N_1049,N_950);
and U1297 (N_1297,In_834,N_1185);
nand U1298 (N_1298,In_1314,N_1171);
and U1299 (N_1299,N_1161,N_1175);
nor U1300 (N_1300,N_724,N_1006);
nor U1301 (N_1301,N_1047,N_67);
and U1302 (N_1302,In_1110,N_888);
and U1303 (N_1303,N_1177,N_1146);
xor U1304 (N_1304,N_410,N_1034);
nand U1305 (N_1305,N_1114,N_514);
xnor U1306 (N_1306,N_1027,N_1016);
nor U1307 (N_1307,N_1108,N_141);
xor U1308 (N_1308,N_814,N_880);
nand U1309 (N_1309,N_1028,N_1181);
or U1310 (N_1310,N_960,N_1182);
and U1311 (N_1311,N_951,N_922);
nor U1312 (N_1312,N_1159,N_1122);
xnor U1313 (N_1313,N_1044,N_1124);
xor U1314 (N_1314,N_1079,N_1020);
xor U1315 (N_1315,N_277,N_1094);
and U1316 (N_1316,N_1136,N_1056);
nor U1317 (N_1317,In_505,N_1037);
nor U1318 (N_1318,N_1048,In_1119);
xor U1319 (N_1319,N_1199,N_1088);
nand U1320 (N_1320,N_878,N_1098);
and U1321 (N_1321,N_1134,In_1327);
or U1322 (N_1322,N_1067,N_1075);
nand U1323 (N_1323,N_907,N_1072);
or U1324 (N_1324,N_1083,N_1093);
and U1325 (N_1325,N_1045,N_1100);
or U1326 (N_1326,N_1153,N_1036);
and U1327 (N_1327,N_1165,N_1024);
and U1328 (N_1328,N_1007,N_1140);
nand U1329 (N_1329,N_838,N_417);
xor U1330 (N_1330,N_1121,N_1170);
and U1331 (N_1331,N_1032,N_1063);
xor U1332 (N_1332,N_1078,N_1021);
nor U1333 (N_1333,N_855,In_1385);
xnor U1334 (N_1334,N_868,In_1266);
nor U1335 (N_1335,In_658,N_1197);
nand U1336 (N_1336,N_802,In_352);
xor U1337 (N_1337,N_1008,N_990);
and U1338 (N_1338,N_1135,N_1046);
nor U1339 (N_1339,N_1105,N_1158);
xor U1340 (N_1340,N_933,N_876);
and U1341 (N_1341,N_1084,N_905);
or U1342 (N_1342,N_1014,N_464);
and U1343 (N_1343,N_1030,N_1156);
and U1344 (N_1344,N_848,N_1186);
or U1345 (N_1345,In_128,In_216);
nor U1346 (N_1346,In_1044,N_624);
and U1347 (N_1347,In_892,N_1062);
nand U1348 (N_1348,N_531,N_772);
xnor U1349 (N_1349,N_952,N_1147);
xnor U1350 (N_1350,N_903,N_1133);
xnor U1351 (N_1351,N_1066,N_1079);
or U1352 (N_1352,N_67,N_410);
and U1353 (N_1353,N_1105,N_1084);
xor U1354 (N_1354,N_845,N_1095);
nor U1355 (N_1355,N_1070,N_1140);
xnor U1356 (N_1356,N_1000,N_1100);
and U1357 (N_1357,N_1103,N_1036);
xnor U1358 (N_1358,N_1144,In_1044);
and U1359 (N_1359,N_1101,In_1385);
nand U1360 (N_1360,N_1006,In_387);
or U1361 (N_1361,N_1053,N_1139);
nand U1362 (N_1362,N_990,N_820);
and U1363 (N_1363,In_1327,N_888);
nand U1364 (N_1364,N_1130,N_1185);
nor U1365 (N_1365,N_896,N_1186);
and U1366 (N_1366,In_352,In_1266);
and U1367 (N_1367,N_1126,N_1073);
or U1368 (N_1368,In_1385,N_595);
nand U1369 (N_1369,In_352,N_141);
or U1370 (N_1370,N_1177,N_1092);
xnor U1371 (N_1371,N_1023,N_1062);
nand U1372 (N_1372,N_724,In_505);
nand U1373 (N_1373,N_1075,N_1034);
or U1374 (N_1374,N_1164,In_1119);
and U1375 (N_1375,N_1163,N_1017);
and U1376 (N_1376,N_679,N_1122);
and U1377 (N_1377,N_410,N_1006);
nor U1378 (N_1378,N_1195,N_936);
xnor U1379 (N_1379,N_726,N_1173);
nor U1380 (N_1380,N_1065,In_387);
or U1381 (N_1381,N_845,N_1045);
or U1382 (N_1382,N_195,N_1127);
nand U1383 (N_1383,N_1155,In_128);
or U1384 (N_1384,N_1179,N_1043);
or U1385 (N_1385,N_1072,N_1036);
xnor U1386 (N_1386,N_1130,N_1025);
xnor U1387 (N_1387,In_1110,N_952);
or U1388 (N_1388,N_1189,N_1191);
and U1389 (N_1389,N_1099,N_1135);
nor U1390 (N_1390,In_1327,N_1033);
and U1391 (N_1391,N_1074,N_1018);
nand U1392 (N_1392,N_933,N_195);
xnor U1393 (N_1393,N_1006,N_1183);
nand U1394 (N_1394,N_961,N_774);
xor U1395 (N_1395,N_1014,N_905);
and U1396 (N_1396,N_1134,N_1001);
nor U1397 (N_1397,N_1136,N_880);
and U1398 (N_1398,N_1195,N_1057);
nand U1399 (N_1399,N_863,N_10);
xor U1400 (N_1400,N_1274,N_1238);
or U1401 (N_1401,N_1313,N_1328);
and U1402 (N_1402,N_1312,N_1320);
nand U1403 (N_1403,N_1381,N_1205);
and U1404 (N_1404,N_1235,N_1366);
or U1405 (N_1405,N_1353,N_1321);
or U1406 (N_1406,N_1318,N_1332);
nand U1407 (N_1407,N_1260,N_1243);
nor U1408 (N_1408,N_1392,N_1391);
xor U1409 (N_1409,N_1300,N_1278);
and U1410 (N_1410,N_1293,N_1246);
and U1411 (N_1411,N_1254,N_1239);
and U1412 (N_1412,N_1292,N_1357);
nor U1413 (N_1413,N_1372,N_1302);
nor U1414 (N_1414,N_1240,N_1331);
nand U1415 (N_1415,N_1206,N_1327);
nor U1416 (N_1416,N_1216,N_1379);
xnor U1417 (N_1417,N_1296,N_1276);
xnor U1418 (N_1418,N_1314,N_1317);
or U1419 (N_1419,N_1242,N_1290);
or U1420 (N_1420,N_1384,N_1396);
and U1421 (N_1421,N_1201,N_1207);
and U1422 (N_1422,N_1291,N_1319);
and U1423 (N_1423,N_1255,N_1250);
nor U1424 (N_1424,N_1237,N_1252);
nand U1425 (N_1425,N_1344,N_1215);
and U1426 (N_1426,N_1299,N_1374);
nor U1427 (N_1427,N_1202,N_1288);
nand U1428 (N_1428,N_1244,N_1295);
xnor U1429 (N_1429,N_1225,N_1270);
xnor U1430 (N_1430,N_1315,N_1306);
or U1431 (N_1431,N_1211,N_1326);
and U1432 (N_1432,N_1347,N_1364);
or U1433 (N_1433,N_1277,N_1325);
nand U1434 (N_1434,N_1218,N_1351);
xor U1435 (N_1435,N_1261,N_1279);
xnor U1436 (N_1436,N_1236,N_1334);
and U1437 (N_1437,N_1375,N_1307);
nand U1438 (N_1438,N_1273,N_1247);
xor U1439 (N_1439,N_1231,N_1224);
and U1440 (N_1440,N_1287,N_1241);
nand U1441 (N_1441,N_1329,N_1387);
and U1442 (N_1442,N_1245,N_1265);
or U1443 (N_1443,N_1308,N_1281);
and U1444 (N_1444,N_1316,N_1219);
xor U1445 (N_1445,N_1249,N_1294);
and U1446 (N_1446,N_1337,N_1282);
and U1447 (N_1447,N_1297,N_1248);
nor U1448 (N_1448,N_1335,N_1266);
nor U1449 (N_1449,N_1272,N_1399);
nor U1450 (N_1450,N_1214,N_1209);
and U1451 (N_1451,N_1359,N_1355);
nand U1452 (N_1452,N_1386,N_1361);
xnor U1453 (N_1453,N_1253,N_1203);
xnor U1454 (N_1454,N_1275,N_1228);
or U1455 (N_1455,N_1298,N_1398);
or U1456 (N_1456,N_1264,N_1305);
or U1457 (N_1457,N_1378,N_1258);
nor U1458 (N_1458,N_1388,N_1232);
nor U1459 (N_1459,N_1286,N_1376);
or U1460 (N_1460,N_1358,N_1268);
or U1461 (N_1461,N_1222,N_1280);
nand U1462 (N_1462,N_1336,N_1251);
nand U1463 (N_1463,N_1352,N_1213);
nor U1464 (N_1464,N_1394,N_1269);
and U1465 (N_1465,N_1200,N_1289);
nand U1466 (N_1466,N_1229,N_1304);
or U1467 (N_1467,N_1283,N_1220);
xor U1468 (N_1468,N_1389,N_1370);
nand U1469 (N_1469,N_1323,N_1371);
nand U1470 (N_1470,N_1223,N_1369);
nand U1471 (N_1471,N_1257,N_1256);
nand U1472 (N_1472,N_1310,N_1385);
nand U1473 (N_1473,N_1330,N_1271);
nand U1474 (N_1474,N_1360,N_1227);
nor U1475 (N_1475,N_1212,N_1363);
and U1476 (N_1476,N_1267,N_1345);
or U1477 (N_1477,N_1348,N_1343);
or U1478 (N_1478,N_1380,N_1210);
nor U1479 (N_1479,N_1393,N_1373);
xor U1480 (N_1480,N_1284,N_1311);
nand U1481 (N_1481,N_1383,N_1259);
nand U1482 (N_1482,N_1263,N_1342);
or U1483 (N_1483,N_1340,N_1322);
or U1484 (N_1484,N_1217,N_1333);
or U1485 (N_1485,N_1362,N_1368);
nand U1486 (N_1486,N_1367,N_1226);
and U1487 (N_1487,N_1350,N_1390);
xnor U1488 (N_1488,N_1341,N_1233);
nand U1489 (N_1489,N_1356,N_1303);
nand U1490 (N_1490,N_1382,N_1338);
and U1491 (N_1491,N_1349,N_1285);
and U1492 (N_1492,N_1221,N_1309);
or U1493 (N_1493,N_1301,N_1234);
and U1494 (N_1494,N_1354,N_1324);
nor U1495 (N_1495,N_1208,N_1262);
xor U1496 (N_1496,N_1365,N_1346);
nor U1497 (N_1497,N_1204,N_1377);
nand U1498 (N_1498,N_1395,N_1339);
or U1499 (N_1499,N_1397,N_1230);
nand U1500 (N_1500,N_1232,N_1272);
or U1501 (N_1501,N_1366,N_1205);
nor U1502 (N_1502,N_1325,N_1367);
or U1503 (N_1503,N_1240,N_1271);
xnor U1504 (N_1504,N_1240,N_1345);
nand U1505 (N_1505,N_1228,N_1253);
nand U1506 (N_1506,N_1228,N_1324);
or U1507 (N_1507,N_1356,N_1232);
or U1508 (N_1508,N_1291,N_1204);
nor U1509 (N_1509,N_1268,N_1337);
nand U1510 (N_1510,N_1280,N_1247);
and U1511 (N_1511,N_1228,N_1224);
or U1512 (N_1512,N_1270,N_1253);
xor U1513 (N_1513,N_1272,N_1261);
or U1514 (N_1514,N_1320,N_1315);
xnor U1515 (N_1515,N_1367,N_1328);
and U1516 (N_1516,N_1232,N_1371);
or U1517 (N_1517,N_1250,N_1303);
nand U1518 (N_1518,N_1396,N_1246);
nor U1519 (N_1519,N_1259,N_1328);
nand U1520 (N_1520,N_1372,N_1388);
and U1521 (N_1521,N_1257,N_1295);
and U1522 (N_1522,N_1265,N_1242);
and U1523 (N_1523,N_1203,N_1245);
nand U1524 (N_1524,N_1295,N_1373);
nand U1525 (N_1525,N_1203,N_1312);
xor U1526 (N_1526,N_1345,N_1327);
nand U1527 (N_1527,N_1234,N_1230);
or U1528 (N_1528,N_1399,N_1362);
or U1529 (N_1529,N_1377,N_1337);
and U1530 (N_1530,N_1316,N_1221);
or U1531 (N_1531,N_1262,N_1209);
xor U1532 (N_1532,N_1393,N_1359);
xnor U1533 (N_1533,N_1344,N_1330);
xor U1534 (N_1534,N_1270,N_1305);
nand U1535 (N_1535,N_1391,N_1352);
and U1536 (N_1536,N_1371,N_1252);
xnor U1537 (N_1537,N_1376,N_1290);
xor U1538 (N_1538,N_1246,N_1241);
or U1539 (N_1539,N_1225,N_1392);
and U1540 (N_1540,N_1221,N_1294);
and U1541 (N_1541,N_1339,N_1320);
and U1542 (N_1542,N_1336,N_1211);
nor U1543 (N_1543,N_1398,N_1307);
nor U1544 (N_1544,N_1367,N_1372);
nor U1545 (N_1545,N_1399,N_1350);
nor U1546 (N_1546,N_1261,N_1253);
and U1547 (N_1547,N_1237,N_1201);
nand U1548 (N_1548,N_1358,N_1260);
nor U1549 (N_1549,N_1241,N_1361);
xnor U1550 (N_1550,N_1386,N_1316);
and U1551 (N_1551,N_1255,N_1264);
or U1552 (N_1552,N_1371,N_1383);
xor U1553 (N_1553,N_1241,N_1354);
nand U1554 (N_1554,N_1363,N_1314);
or U1555 (N_1555,N_1341,N_1323);
or U1556 (N_1556,N_1296,N_1271);
nor U1557 (N_1557,N_1328,N_1344);
and U1558 (N_1558,N_1377,N_1248);
and U1559 (N_1559,N_1298,N_1248);
nand U1560 (N_1560,N_1244,N_1314);
nor U1561 (N_1561,N_1369,N_1370);
nand U1562 (N_1562,N_1320,N_1241);
or U1563 (N_1563,N_1353,N_1352);
and U1564 (N_1564,N_1315,N_1358);
nand U1565 (N_1565,N_1239,N_1394);
and U1566 (N_1566,N_1361,N_1331);
nor U1567 (N_1567,N_1336,N_1265);
nor U1568 (N_1568,N_1342,N_1325);
and U1569 (N_1569,N_1258,N_1274);
nor U1570 (N_1570,N_1374,N_1375);
nor U1571 (N_1571,N_1375,N_1243);
and U1572 (N_1572,N_1339,N_1354);
xor U1573 (N_1573,N_1354,N_1396);
or U1574 (N_1574,N_1227,N_1214);
and U1575 (N_1575,N_1254,N_1368);
nor U1576 (N_1576,N_1245,N_1389);
and U1577 (N_1577,N_1259,N_1343);
nor U1578 (N_1578,N_1327,N_1392);
and U1579 (N_1579,N_1249,N_1214);
nor U1580 (N_1580,N_1232,N_1253);
or U1581 (N_1581,N_1332,N_1233);
nand U1582 (N_1582,N_1363,N_1315);
nor U1583 (N_1583,N_1274,N_1211);
and U1584 (N_1584,N_1334,N_1245);
or U1585 (N_1585,N_1332,N_1301);
or U1586 (N_1586,N_1286,N_1242);
nand U1587 (N_1587,N_1242,N_1205);
nor U1588 (N_1588,N_1333,N_1291);
and U1589 (N_1589,N_1308,N_1370);
or U1590 (N_1590,N_1255,N_1262);
nand U1591 (N_1591,N_1239,N_1327);
nand U1592 (N_1592,N_1370,N_1246);
nand U1593 (N_1593,N_1308,N_1236);
and U1594 (N_1594,N_1284,N_1245);
nand U1595 (N_1595,N_1315,N_1251);
nor U1596 (N_1596,N_1354,N_1281);
nand U1597 (N_1597,N_1208,N_1318);
or U1598 (N_1598,N_1203,N_1398);
nor U1599 (N_1599,N_1331,N_1280);
or U1600 (N_1600,N_1520,N_1577);
xnor U1601 (N_1601,N_1594,N_1427);
xor U1602 (N_1602,N_1470,N_1516);
or U1603 (N_1603,N_1551,N_1450);
or U1604 (N_1604,N_1558,N_1596);
nand U1605 (N_1605,N_1499,N_1403);
xnor U1606 (N_1606,N_1591,N_1574);
xnor U1607 (N_1607,N_1465,N_1421);
nor U1608 (N_1608,N_1428,N_1512);
or U1609 (N_1609,N_1480,N_1413);
and U1610 (N_1610,N_1419,N_1458);
or U1611 (N_1611,N_1595,N_1584);
and U1612 (N_1612,N_1505,N_1547);
nand U1613 (N_1613,N_1410,N_1473);
or U1614 (N_1614,N_1502,N_1579);
and U1615 (N_1615,N_1518,N_1400);
or U1616 (N_1616,N_1495,N_1441);
nand U1617 (N_1617,N_1416,N_1503);
nor U1618 (N_1618,N_1571,N_1501);
xor U1619 (N_1619,N_1424,N_1426);
and U1620 (N_1620,N_1570,N_1530);
nand U1621 (N_1621,N_1554,N_1529);
and U1622 (N_1622,N_1531,N_1408);
nand U1623 (N_1623,N_1477,N_1437);
nor U1624 (N_1624,N_1412,N_1468);
nand U1625 (N_1625,N_1542,N_1401);
xor U1626 (N_1626,N_1525,N_1515);
and U1627 (N_1627,N_1583,N_1455);
and U1628 (N_1628,N_1585,N_1500);
nor U1629 (N_1629,N_1418,N_1472);
xnor U1630 (N_1630,N_1507,N_1454);
xor U1631 (N_1631,N_1589,N_1576);
xnor U1632 (N_1632,N_1466,N_1405);
nand U1633 (N_1633,N_1463,N_1537);
xnor U1634 (N_1634,N_1479,N_1580);
nand U1635 (N_1635,N_1434,N_1453);
or U1636 (N_1636,N_1549,N_1557);
and U1637 (N_1637,N_1414,N_1487);
nor U1638 (N_1638,N_1544,N_1447);
xnor U1639 (N_1639,N_1578,N_1481);
nor U1640 (N_1640,N_1526,N_1429);
nor U1641 (N_1641,N_1435,N_1425);
and U1642 (N_1642,N_1522,N_1491);
and U1643 (N_1643,N_1467,N_1444);
xor U1644 (N_1644,N_1431,N_1432);
nor U1645 (N_1645,N_1469,N_1494);
xor U1646 (N_1646,N_1567,N_1508);
or U1647 (N_1647,N_1423,N_1485);
and U1648 (N_1648,N_1460,N_1433);
nand U1649 (N_1649,N_1451,N_1521);
or U1650 (N_1650,N_1540,N_1457);
nor U1651 (N_1651,N_1588,N_1556);
xnor U1652 (N_1652,N_1566,N_1486);
or U1653 (N_1653,N_1514,N_1440);
and U1654 (N_1654,N_1406,N_1517);
xor U1655 (N_1655,N_1476,N_1528);
nor U1656 (N_1656,N_1575,N_1541);
and U1657 (N_1657,N_1523,N_1543);
and U1658 (N_1658,N_1488,N_1404);
or U1659 (N_1659,N_1459,N_1545);
nor U1660 (N_1660,N_1442,N_1409);
or U1661 (N_1661,N_1561,N_1527);
or U1662 (N_1662,N_1436,N_1464);
or U1663 (N_1663,N_1498,N_1592);
and U1664 (N_1664,N_1446,N_1496);
nand U1665 (N_1665,N_1497,N_1555);
nand U1666 (N_1666,N_1534,N_1538);
or U1667 (N_1667,N_1510,N_1563);
nand U1668 (N_1668,N_1559,N_1402);
or U1669 (N_1669,N_1581,N_1415);
xor U1670 (N_1670,N_1471,N_1519);
nand U1671 (N_1671,N_1513,N_1532);
nand U1672 (N_1672,N_1482,N_1443);
or U1673 (N_1673,N_1587,N_1449);
nand U1674 (N_1674,N_1484,N_1417);
and U1675 (N_1675,N_1461,N_1572);
nand U1676 (N_1676,N_1539,N_1439);
nand U1677 (N_1677,N_1565,N_1483);
and U1678 (N_1678,N_1490,N_1420);
xnor U1679 (N_1679,N_1456,N_1552);
nand U1680 (N_1680,N_1511,N_1564);
nand U1681 (N_1681,N_1535,N_1548);
or U1682 (N_1682,N_1422,N_1573);
xnor U1683 (N_1683,N_1562,N_1590);
or U1684 (N_1684,N_1478,N_1452);
nand U1685 (N_1685,N_1504,N_1493);
nand U1686 (N_1686,N_1509,N_1462);
and U1687 (N_1687,N_1430,N_1586);
xnor U1688 (N_1688,N_1568,N_1546);
xor U1689 (N_1689,N_1489,N_1536);
nand U1690 (N_1690,N_1593,N_1492);
xnor U1691 (N_1691,N_1407,N_1597);
xnor U1692 (N_1692,N_1411,N_1438);
and U1693 (N_1693,N_1560,N_1553);
nor U1694 (N_1694,N_1506,N_1550);
and U1695 (N_1695,N_1569,N_1533);
xnor U1696 (N_1696,N_1524,N_1475);
xnor U1697 (N_1697,N_1474,N_1582);
xnor U1698 (N_1698,N_1445,N_1448);
and U1699 (N_1699,N_1598,N_1599);
nand U1700 (N_1700,N_1459,N_1494);
nor U1701 (N_1701,N_1546,N_1433);
or U1702 (N_1702,N_1562,N_1586);
xnor U1703 (N_1703,N_1570,N_1528);
nor U1704 (N_1704,N_1409,N_1550);
and U1705 (N_1705,N_1476,N_1489);
nor U1706 (N_1706,N_1446,N_1533);
xor U1707 (N_1707,N_1523,N_1481);
or U1708 (N_1708,N_1407,N_1454);
or U1709 (N_1709,N_1578,N_1453);
xor U1710 (N_1710,N_1519,N_1423);
and U1711 (N_1711,N_1541,N_1593);
nand U1712 (N_1712,N_1574,N_1522);
and U1713 (N_1713,N_1573,N_1425);
nand U1714 (N_1714,N_1462,N_1424);
nor U1715 (N_1715,N_1564,N_1468);
and U1716 (N_1716,N_1417,N_1413);
or U1717 (N_1717,N_1549,N_1456);
nand U1718 (N_1718,N_1510,N_1508);
nor U1719 (N_1719,N_1584,N_1576);
xnor U1720 (N_1720,N_1591,N_1511);
nor U1721 (N_1721,N_1439,N_1418);
xnor U1722 (N_1722,N_1457,N_1451);
and U1723 (N_1723,N_1487,N_1592);
nor U1724 (N_1724,N_1575,N_1598);
or U1725 (N_1725,N_1406,N_1533);
nand U1726 (N_1726,N_1452,N_1487);
or U1727 (N_1727,N_1576,N_1529);
xor U1728 (N_1728,N_1410,N_1564);
or U1729 (N_1729,N_1527,N_1567);
or U1730 (N_1730,N_1583,N_1428);
or U1731 (N_1731,N_1572,N_1521);
and U1732 (N_1732,N_1475,N_1590);
and U1733 (N_1733,N_1409,N_1423);
nand U1734 (N_1734,N_1450,N_1466);
nor U1735 (N_1735,N_1596,N_1446);
nand U1736 (N_1736,N_1443,N_1500);
xnor U1737 (N_1737,N_1489,N_1550);
and U1738 (N_1738,N_1547,N_1508);
nor U1739 (N_1739,N_1500,N_1440);
nand U1740 (N_1740,N_1532,N_1540);
and U1741 (N_1741,N_1555,N_1514);
nor U1742 (N_1742,N_1426,N_1475);
or U1743 (N_1743,N_1470,N_1416);
and U1744 (N_1744,N_1410,N_1459);
or U1745 (N_1745,N_1561,N_1471);
nand U1746 (N_1746,N_1475,N_1403);
or U1747 (N_1747,N_1582,N_1579);
and U1748 (N_1748,N_1556,N_1506);
nand U1749 (N_1749,N_1569,N_1597);
and U1750 (N_1750,N_1460,N_1533);
xor U1751 (N_1751,N_1592,N_1524);
and U1752 (N_1752,N_1503,N_1483);
or U1753 (N_1753,N_1512,N_1471);
nand U1754 (N_1754,N_1598,N_1554);
nand U1755 (N_1755,N_1568,N_1476);
nand U1756 (N_1756,N_1503,N_1412);
xor U1757 (N_1757,N_1551,N_1577);
and U1758 (N_1758,N_1539,N_1546);
xnor U1759 (N_1759,N_1496,N_1420);
or U1760 (N_1760,N_1444,N_1549);
nand U1761 (N_1761,N_1508,N_1518);
nand U1762 (N_1762,N_1551,N_1449);
nor U1763 (N_1763,N_1595,N_1461);
and U1764 (N_1764,N_1493,N_1548);
or U1765 (N_1765,N_1584,N_1551);
nand U1766 (N_1766,N_1485,N_1461);
xor U1767 (N_1767,N_1462,N_1558);
nand U1768 (N_1768,N_1545,N_1426);
and U1769 (N_1769,N_1503,N_1518);
or U1770 (N_1770,N_1521,N_1509);
nand U1771 (N_1771,N_1434,N_1546);
and U1772 (N_1772,N_1429,N_1511);
nand U1773 (N_1773,N_1509,N_1531);
and U1774 (N_1774,N_1495,N_1491);
xnor U1775 (N_1775,N_1509,N_1550);
xor U1776 (N_1776,N_1542,N_1488);
and U1777 (N_1777,N_1463,N_1557);
nor U1778 (N_1778,N_1497,N_1500);
xnor U1779 (N_1779,N_1523,N_1427);
and U1780 (N_1780,N_1568,N_1523);
and U1781 (N_1781,N_1489,N_1563);
nand U1782 (N_1782,N_1500,N_1421);
nand U1783 (N_1783,N_1528,N_1472);
and U1784 (N_1784,N_1578,N_1495);
nand U1785 (N_1785,N_1512,N_1582);
or U1786 (N_1786,N_1521,N_1454);
xnor U1787 (N_1787,N_1550,N_1473);
or U1788 (N_1788,N_1475,N_1534);
nor U1789 (N_1789,N_1512,N_1422);
nand U1790 (N_1790,N_1534,N_1467);
xnor U1791 (N_1791,N_1595,N_1481);
nand U1792 (N_1792,N_1563,N_1513);
nor U1793 (N_1793,N_1552,N_1441);
xor U1794 (N_1794,N_1424,N_1529);
or U1795 (N_1795,N_1450,N_1422);
nand U1796 (N_1796,N_1523,N_1467);
and U1797 (N_1797,N_1472,N_1463);
nor U1798 (N_1798,N_1443,N_1588);
xnor U1799 (N_1799,N_1429,N_1563);
nor U1800 (N_1800,N_1742,N_1730);
nand U1801 (N_1801,N_1754,N_1637);
and U1802 (N_1802,N_1632,N_1728);
or U1803 (N_1803,N_1723,N_1688);
nor U1804 (N_1804,N_1641,N_1691);
nor U1805 (N_1805,N_1602,N_1617);
xor U1806 (N_1806,N_1779,N_1702);
nor U1807 (N_1807,N_1638,N_1727);
xnor U1808 (N_1808,N_1701,N_1785);
nand U1809 (N_1809,N_1628,N_1650);
nor U1810 (N_1810,N_1680,N_1747);
nor U1811 (N_1811,N_1651,N_1794);
or U1812 (N_1812,N_1777,N_1662);
xnor U1813 (N_1813,N_1690,N_1738);
or U1814 (N_1814,N_1658,N_1741);
and U1815 (N_1815,N_1737,N_1645);
xnor U1816 (N_1816,N_1799,N_1603);
or U1817 (N_1817,N_1619,N_1614);
nand U1818 (N_1818,N_1761,N_1732);
nand U1819 (N_1819,N_1698,N_1715);
nor U1820 (N_1820,N_1610,N_1601);
nand U1821 (N_1821,N_1615,N_1788);
or U1822 (N_1822,N_1720,N_1669);
or U1823 (N_1823,N_1791,N_1739);
xor U1824 (N_1824,N_1616,N_1607);
nand U1825 (N_1825,N_1784,N_1623);
or U1826 (N_1826,N_1774,N_1697);
and U1827 (N_1827,N_1653,N_1656);
or U1828 (N_1828,N_1647,N_1795);
and U1829 (N_1829,N_1740,N_1709);
nand U1830 (N_1830,N_1765,N_1703);
nor U1831 (N_1831,N_1682,N_1776);
or U1832 (N_1832,N_1612,N_1636);
xor U1833 (N_1833,N_1724,N_1762);
xor U1834 (N_1834,N_1790,N_1604);
xnor U1835 (N_1835,N_1686,N_1700);
nand U1836 (N_1836,N_1640,N_1778);
nand U1837 (N_1837,N_1758,N_1683);
nand U1838 (N_1838,N_1675,N_1644);
xor U1839 (N_1839,N_1753,N_1664);
nor U1840 (N_1840,N_1764,N_1618);
nor U1841 (N_1841,N_1659,N_1770);
or U1842 (N_1842,N_1714,N_1671);
nor U1843 (N_1843,N_1633,N_1689);
nor U1844 (N_1844,N_1749,N_1755);
xor U1845 (N_1845,N_1626,N_1735);
nand U1846 (N_1846,N_1783,N_1781);
nand U1847 (N_1847,N_1726,N_1678);
nand U1848 (N_1848,N_1734,N_1699);
and U1849 (N_1849,N_1661,N_1608);
or U1850 (N_1850,N_1793,N_1635);
nand U1851 (N_1851,N_1771,N_1677);
nor U1852 (N_1852,N_1773,N_1622);
nor U1853 (N_1853,N_1706,N_1634);
or U1854 (N_1854,N_1796,N_1772);
nand U1855 (N_1855,N_1789,N_1694);
nor U1856 (N_1856,N_1696,N_1759);
and U1857 (N_1857,N_1655,N_1639);
and U1858 (N_1858,N_1695,N_1707);
and U1859 (N_1859,N_1775,N_1752);
xor U1860 (N_1860,N_1692,N_1668);
or U1861 (N_1861,N_1704,N_1798);
and U1862 (N_1862,N_1693,N_1681);
or U1863 (N_1863,N_1767,N_1663);
nand U1864 (N_1864,N_1600,N_1782);
xor U1865 (N_1865,N_1670,N_1712);
and U1866 (N_1866,N_1713,N_1672);
or U1867 (N_1867,N_1751,N_1743);
nand U1868 (N_1868,N_1792,N_1605);
nor U1869 (N_1869,N_1621,N_1642);
xnor U1870 (N_1870,N_1613,N_1630);
and U1871 (N_1871,N_1673,N_1666);
or U1872 (N_1872,N_1648,N_1708);
or U1873 (N_1873,N_1768,N_1705);
nand U1874 (N_1874,N_1780,N_1620);
and U1875 (N_1875,N_1652,N_1763);
or U1876 (N_1876,N_1611,N_1731);
or U1877 (N_1877,N_1625,N_1760);
or U1878 (N_1878,N_1711,N_1756);
and U1879 (N_1879,N_1721,N_1736);
nor U1880 (N_1880,N_1766,N_1654);
and U1881 (N_1881,N_1665,N_1733);
and U1882 (N_1882,N_1629,N_1609);
xor U1883 (N_1883,N_1729,N_1744);
or U1884 (N_1884,N_1718,N_1719);
and U1885 (N_1885,N_1716,N_1748);
nand U1886 (N_1886,N_1649,N_1606);
nor U1887 (N_1887,N_1660,N_1631);
and U1888 (N_1888,N_1722,N_1710);
nand U1889 (N_1889,N_1750,N_1687);
nor U1890 (N_1890,N_1643,N_1646);
xnor U1891 (N_1891,N_1627,N_1757);
nor U1892 (N_1892,N_1667,N_1725);
or U1893 (N_1893,N_1797,N_1685);
or U1894 (N_1894,N_1786,N_1684);
and U1895 (N_1895,N_1676,N_1674);
xor U1896 (N_1896,N_1769,N_1745);
and U1897 (N_1897,N_1787,N_1624);
and U1898 (N_1898,N_1657,N_1717);
nor U1899 (N_1899,N_1746,N_1679);
or U1900 (N_1900,N_1760,N_1790);
or U1901 (N_1901,N_1746,N_1707);
and U1902 (N_1902,N_1610,N_1790);
nor U1903 (N_1903,N_1708,N_1653);
and U1904 (N_1904,N_1672,N_1769);
nor U1905 (N_1905,N_1748,N_1759);
nor U1906 (N_1906,N_1654,N_1660);
and U1907 (N_1907,N_1724,N_1674);
or U1908 (N_1908,N_1710,N_1738);
or U1909 (N_1909,N_1731,N_1629);
or U1910 (N_1910,N_1631,N_1731);
nand U1911 (N_1911,N_1634,N_1608);
nor U1912 (N_1912,N_1756,N_1737);
and U1913 (N_1913,N_1608,N_1781);
nand U1914 (N_1914,N_1610,N_1721);
nor U1915 (N_1915,N_1793,N_1720);
or U1916 (N_1916,N_1775,N_1655);
or U1917 (N_1917,N_1760,N_1730);
and U1918 (N_1918,N_1701,N_1686);
xnor U1919 (N_1919,N_1682,N_1636);
nor U1920 (N_1920,N_1684,N_1673);
nand U1921 (N_1921,N_1764,N_1734);
nor U1922 (N_1922,N_1634,N_1755);
or U1923 (N_1923,N_1798,N_1667);
nor U1924 (N_1924,N_1753,N_1648);
and U1925 (N_1925,N_1657,N_1638);
xnor U1926 (N_1926,N_1611,N_1649);
xnor U1927 (N_1927,N_1709,N_1763);
nand U1928 (N_1928,N_1792,N_1708);
nand U1929 (N_1929,N_1725,N_1769);
and U1930 (N_1930,N_1697,N_1610);
and U1931 (N_1931,N_1699,N_1613);
or U1932 (N_1932,N_1702,N_1682);
and U1933 (N_1933,N_1794,N_1613);
nand U1934 (N_1934,N_1756,N_1680);
and U1935 (N_1935,N_1789,N_1687);
or U1936 (N_1936,N_1759,N_1640);
nor U1937 (N_1937,N_1781,N_1750);
nor U1938 (N_1938,N_1732,N_1745);
xor U1939 (N_1939,N_1752,N_1725);
nor U1940 (N_1940,N_1683,N_1753);
and U1941 (N_1941,N_1765,N_1688);
and U1942 (N_1942,N_1670,N_1708);
xnor U1943 (N_1943,N_1661,N_1766);
and U1944 (N_1944,N_1685,N_1794);
or U1945 (N_1945,N_1707,N_1749);
nand U1946 (N_1946,N_1764,N_1793);
nor U1947 (N_1947,N_1707,N_1618);
xor U1948 (N_1948,N_1742,N_1691);
and U1949 (N_1949,N_1666,N_1708);
nor U1950 (N_1950,N_1795,N_1777);
and U1951 (N_1951,N_1605,N_1771);
or U1952 (N_1952,N_1635,N_1679);
and U1953 (N_1953,N_1755,N_1789);
and U1954 (N_1954,N_1696,N_1620);
nand U1955 (N_1955,N_1720,N_1609);
or U1956 (N_1956,N_1680,N_1650);
xor U1957 (N_1957,N_1762,N_1632);
nand U1958 (N_1958,N_1760,N_1744);
or U1959 (N_1959,N_1655,N_1770);
nand U1960 (N_1960,N_1630,N_1627);
and U1961 (N_1961,N_1797,N_1615);
or U1962 (N_1962,N_1776,N_1616);
nand U1963 (N_1963,N_1664,N_1767);
and U1964 (N_1964,N_1634,N_1749);
or U1965 (N_1965,N_1741,N_1766);
nor U1966 (N_1966,N_1723,N_1776);
or U1967 (N_1967,N_1798,N_1745);
xnor U1968 (N_1968,N_1672,N_1775);
and U1969 (N_1969,N_1636,N_1652);
and U1970 (N_1970,N_1620,N_1707);
nor U1971 (N_1971,N_1686,N_1741);
xor U1972 (N_1972,N_1725,N_1623);
nor U1973 (N_1973,N_1741,N_1646);
nand U1974 (N_1974,N_1683,N_1725);
nand U1975 (N_1975,N_1750,N_1646);
nor U1976 (N_1976,N_1748,N_1647);
xor U1977 (N_1977,N_1776,N_1685);
nand U1978 (N_1978,N_1752,N_1732);
xnor U1979 (N_1979,N_1664,N_1736);
or U1980 (N_1980,N_1777,N_1712);
nand U1981 (N_1981,N_1659,N_1695);
xor U1982 (N_1982,N_1741,N_1749);
nand U1983 (N_1983,N_1647,N_1634);
nor U1984 (N_1984,N_1719,N_1612);
nand U1985 (N_1985,N_1609,N_1707);
nor U1986 (N_1986,N_1646,N_1787);
or U1987 (N_1987,N_1796,N_1629);
nor U1988 (N_1988,N_1666,N_1796);
nand U1989 (N_1989,N_1765,N_1650);
and U1990 (N_1990,N_1797,N_1712);
nand U1991 (N_1991,N_1676,N_1744);
or U1992 (N_1992,N_1792,N_1739);
nor U1993 (N_1993,N_1773,N_1663);
and U1994 (N_1994,N_1723,N_1614);
nor U1995 (N_1995,N_1658,N_1689);
and U1996 (N_1996,N_1735,N_1611);
or U1997 (N_1997,N_1745,N_1794);
nor U1998 (N_1998,N_1710,N_1744);
nor U1999 (N_1999,N_1656,N_1739);
nor U2000 (N_2000,N_1951,N_1970);
and U2001 (N_2001,N_1899,N_1925);
nand U2002 (N_2002,N_1892,N_1927);
and U2003 (N_2003,N_1848,N_1859);
and U2004 (N_2004,N_1812,N_1871);
xnor U2005 (N_2005,N_1889,N_1864);
or U2006 (N_2006,N_1893,N_1847);
nor U2007 (N_2007,N_1860,N_1988);
or U2008 (N_2008,N_1833,N_1849);
and U2009 (N_2009,N_1972,N_1883);
nor U2010 (N_2010,N_1809,N_1828);
or U2011 (N_2011,N_1863,N_1855);
nor U2012 (N_2012,N_1983,N_1817);
nor U2013 (N_2013,N_1932,N_1999);
xnor U2014 (N_2014,N_1954,N_1955);
nand U2015 (N_2015,N_1894,N_1853);
xnor U2016 (N_2016,N_1857,N_1963);
and U2017 (N_2017,N_1827,N_1912);
nor U2018 (N_2018,N_1906,N_1978);
or U2019 (N_2019,N_1820,N_1982);
nand U2020 (N_2020,N_1844,N_1953);
or U2021 (N_2021,N_1800,N_1959);
xnor U2022 (N_2022,N_1845,N_1920);
or U2023 (N_2023,N_1815,N_1869);
xnor U2024 (N_2024,N_1938,N_1896);
nor U2025 (N_2025,N_1856,N_1923);
or U2026 (N_2026,N_1877,N_1985);
nor U2027 (N_2027,N_1830,N_1801);
nand U2028 (N_2028,N_1861,N_1885);
nor U2029 (N_2029,N_1980,N_1974);
xor U2030 (N_2030,N_1875,N_1836);
xor U2031 (N_2031,N_1891,N_1876);
and U2032 (N_2032,N_1942,N_1803);
xnor U2033 (N_2033,N_1916,N_1966);
or U2034 (N_2034,N_1890,N_1957);
nor U2035 (N_2035,N_1948,N_1979);
or U2036 (N_2036,N_1804,N_1986);
and U2037 (N_2037,N_1901,N_1882);
nand U2038 (N_2038,N_1850,N_1872);
nor U2039 (N_2039,N_1945,N_1989);
or U2040 (N_2040,N_1821,N_1858);
and U2041 (N_2041,N_1822,N_1840);
xnor U2042 (N_2042,N_1984,N_1825);
and U2043 (N_2043,N_1996,N_1919);
nand U2044 (N_2044,N_1843,N_1995);
xor U2045 (N_2045,N_1929,N_1903);
xor U2046 (N_2046,N_1941,N_1917);
nand U2047 (N_2047,N_1939,N_1926);
and U2048 (N_2048,N_1897,N_1818);
xor U2049 (N_2049,N_1922,N_1826);
xor U2050 (N_2050,N_1993,N_1943);
or U2051 (N_2051,N_1835,N_1905);
nand U2052 (N_2052,N_1937,N_1909);
nor U2053 (N_2053,N_1928,N_1958);
xnor U2054 (N_2054,N_1884,N_1965);
and U2055 (N_2055,N_1878,N_1839);
and U2056 (N_2056,N_1887,N_1910);
nand U2057 (N_2057,N_1831,N_1870);
nand U2058 (N_2058,N_1971,N_1908);
and U2059 (N_2059,N_1862,N_1935);
nor U2060 (N_2060,N_1832,N_1969);
xor U2061 (N_2061,N_1807,N_1900);
and U2062 (N_2062,N_1808,N_1911);
or U2063 (N_2063,N_1962,N_1838);
nand U2064 (N_2064,N_1829,N_1865);
or U2065 (N_2065,N_1898,N_1998);
and U2066 (N_2066,N_1805,N_1936);
and U2067 (N_2067,N_1886,N_1994);
or U2068 (N_2068,N_1921,N_1823);
xor U2069 (N_2069,N_1946,N_1924);
nand U2070 (N_2070,N_1879,N_1846);
nor U2071 (N_2071,N_1981,N_1888);
nand U2072 (N_2072,N_1913,N_1934);
nor U2073 (N_2073,N_1873,N_1866);
or U2074 (N_2074,N_1930,N_1907);
and U2075 (N_2075,N_1868,N_1904);
or U2076 (N_2076,N_1990,N_1960);
nand U2077 (N_2077,N_1854,N_1811);
and U2078 (N_2078,N_1947,N_1964);
nand U2079 (N_2079,N_1810,N_1976);
or U2080 (N_2080,N_1956,N_1874);
and U2081 (N_2081,N_1992,N_1813);
nor U2082 (N_2082,N_1881,N_1814);
or U2083 (N_2083,N_1952,N_1991);
nor U2084 (N_2084,N_1842,N_1997);
and U2085 (N_2085,N_1895,N_1819);
or U2086 (N_2086,N_1973,N_1816);
xnor U2087 (N_2087,N_1802,N_1968);
and U2088 (N_2088,N_1834,N_1915);
nand U2089 (N_2089,N_1851,N_1944);
or U2090 (N_2090,N_1987,N_1940);
xnor U2091 (N_2091,N_1902,N_1931);
xnor U2092 (N_2092,N_1806,N_1824);
or U2093 (N_2093,N_1837,N_1867);
nor U2094 (N_2094,N_1933,N_1975);
nor U2095 (N_2095,N_1950,N_1852);
or U2096 (N_2096,N_1880,N_1967);
nand U2097 (N_2097,N_1949,N_1918);
xor U2098 (N_2098,N_1977,N_1841);
or U2099 (N_2099,N_1961,N_1914);
nor U2100 (N_2100,N_1838,N_1957);
nand U2101 (N_2101,N_1861,N_1971);
or U2102 (N_2102,N_1972,N_1937);
and U2103 (N_2103,N_1870,N_1983);
or U2104 (N_2104,N_1853,N_1805);
xor U2105 (N_2105,N_1810,N_1920);
xnor U2106 (N_2106,N_1924,N_1872);
xnor U2107 (N_2107,N_1802,N_1974);
and U2108 (N_2108,N_1855,N_1954);
or U2109 (N_2109,N_1937,N_1928);
and U2110 (N_2110,N_1960,N_1912);
or U2111 (N_2111,N_1916,N_1808);
or U2112 (N_2112,N_1987,N_1885);
and U2113 (N_2113,N_1986,N_1819);
nor U2114 (N_2114,N_1956,N_1959);
nor U2115 (N_2115,N_1882,N_1978);
nor U2116 (N_2116,N_1881,N_1933);
and U2117 (N_2117,N_1964,N_1913);
and U2118 (N_2118,N_1959,N_1888);
nand U2119 (N_2119,N_1874,N_1919);
or U2120 (N_2120,N_1834,N_1957);
or U2121 (N_2121,N_1962,N_1973);
nor U2122 (N_2122,N_1825,N_1853);
nand U2123 (N_2123,N_1801,N_1855);
and U2124 (N_2124,N_1850,N_1914);
nor U2125 (N_2125,N_1926,N_1901);
or U2126 (N_2126,N_1901,N_1973);
and U2127 (N_2127,N_1983,N_1873);
nand U2128 (N_2128,N_1974,N_1891);
nand U2129 (N_2129,N_1800,N_1891);
and U2130 (N_2130,N_1972,N_1911);
nand U2131 (N_2131,N_1929,N_1863);
xnor U2132 (N_2132,N_1856,N_1945);
nor U2133 (N_2133,N_1946,N_1965);
nor U2134 (N_2134,N_1821,N_1814);
nor U2135 (N_2135,N_1885,N_1990);
nor U2136 (N_2136,N_1904,N_1981);
xor U2137 (N_2137,N_1856,N_1808);
and U2138 (N_2138,N_1925,N_1912);
xor U2139 (N_2139,N_1973,N_1910);
or U2140 (N_2140,N_1977,N_1871);
and U2141 (N_2141,N_1913,N_1801);
nor U2142 (N_2142,N_1946,N_1990);
xor U2143 (N_2143,N_1905,N_1864);
and U2144 (N_2144,N_1960,N_1807);
or U2145 (N_2145,N_1911,N_1836);
and U2146 (N_2146,N_1864,N_1829);
or U2147 (N_2147,N_1961,N_1874);
nand U2148 (N_2148,N_1905,N_1906);
nor U2149 (N_2149,N_1818,N_1928);
nor U2150 (N_2150,N_1883,N_1945);
and U2151 (N_2151,N_1830,N_1806);
nand U2152 (N_2152,N_1838,N_1827);
and U2153 (N_2153,N_1893,N_1950);
xnor U2154 (N_2154,N_1950,N_1836);
nor U2155 (N_2155,N_1971,N_1901);
and U2156 (N_2156,N_1987,N_1834);
or U2157 (N_2157,N_1901,N_1990);
nor U2158 (N_2158,N_1961,N_1856);
nand U2159 (N_2159,N_1830,N_1950);
nand U2160 (N_2160,N_1843,N_1801);
xor U2161 (N_2161,N_1874,N_1825);
or U2162 (N_2162,N_1835,N_1932);
nand U2163 (N_2163,N_1843,N_1973);
xor U2164 (N_2164,N_1974,N_1938);
or U2165 (N_2165,N_1930,N_1818);
and U2166 (N_2166,N_1989,N_1800);
or U2167 (N_2167,N_1857,N_1811);
xor U2168 (N_2168,N_1818,N_1977);
xnor U2169 (N_2169,N_1800,N_1896);
xnor U2170 (N_2170,N_1952,N_1809);
nor U2171 (N_2171,N_1876,N_1838);
nor U2172 (N_2172,N_1831,N_1859);
nand U2173 (N_2173,N_1937,N_1974);
and U2174 (N_2174,N_1881,N_1844);
nand U2175 (N_2175,N_1815,N_1825);
nor U2176 (N_2176,N_1932,N_1816);
xor U2177 (N_2177,N_1947,N_1837);
or U2178 (N_2178,N_1987,N_1903);
nand U2179 (N_2179,N_1964,N_1832);
xnor U2180 (N_2180,N_1863,N_1827);
xor U2181 (N_2181,N_1815,N_1953);
nor U2182 (N_2182,N_1861,N_1980);
and U2183 (N_2183,N_1863,N_1941);
xor U2184 (N_2184,N_1977,N_1835);
xnor U2185 (N_2185,N_1852,N_1856);
nand U2186 (N_2186,N_1873,N_1923);
nor U2187 (N_2187,N_1902,N_1855);
and U2188 (N_2188,N_1920,N_1824);
and U2189 (N_2189,N_1829,N_1870);
nor U2190 (N_2190,N_1995,N_1823);
xor U2191 (N_2191,N_1823,N_1889);
nand U2192 (N_2192,N_1845,N_1872);
or U2193 (N_2193,N_1956,N_1904);
and U2194 (N_2194,N_1869,N_1824);
nor U2195 (N_2195,N_1979,N_1900);
xnor U2196 (N_2196,N_1979,N_1803);
nor U2197 (N_2197,N_1815,N_1957);
and U2198 (N_2198,N_1819,N_1832);
or U2199 (N_2199,N_1881,N_1876);
and U2200 (N_2200,N_2158,N_2162);
xor U2201 (N_2201,N_2142,N_2067);
nor U2202 (N_2202,N_2066,N_2185);
nor U2203 (N_2203,N_2049,N_2004);
xor U2204 (N_2204,N_2083,N_2030);
xor U2205 (N_2205,N_2039,N_2051);
or U2206 (N_2206,N_2029,N_2034);
xnor U2207 (N_2207,N_2178,N_2168);
xor U2208 (N_2208,N_2044,N_2155);
or U2209 (N_2209,N_2194,N_2056);
nand U2210 (N_2210,N_2035,N_2015);
xor U2211 (N_2211,N_2046,N_2139);
nor U2212 (N_2212,N_2005,N_2058);
and U2213 (N_2213,N_2076,N_2082);
nor U2214 (N_2214,N_2060,N_2064);
nand U2215 (N_2215,N_2175,N_2053);
or U2216 (N_2216,N_2144,N_2013);
and U2217 (N_2217,N_2093,N_2106);
xnor U2218 (N_2218,N_2192,N_2000);
xnor U2219 (N_2219,N_2129,N_2100);
nand U2220 (N_2220,N_2117,N_2141);
and U2221 (N_2221,N_2102,N_2062);
nand U2222 (N_2222,N_2059,N_2161);
xnor U2223 (N_2223,N_2078,N_2176);
nand U2224 (N_2224,N_2113,N_2151);
nand U2225 (N_2225,N_2114,N_2198);
and U2226 (N_2226,N_2169,N_2024);
nand U2227 (N_2227,N_2080,N_2170);
nor U2228 (N_2228,N_2181,N_2027);
xnor U2229 (N_2229,N_2196,N_2009);
xor U2230 (N_2230,N_2197,N_2098);
and U2231 (N_2231,N_2130,N_2043);
xnor U2232 (N_2232,N_2026,N_2157);
or U2233 (N_2233,N_2074,N_2002);
and U2234 (N_2234,N_2111,N_2146);
nor U2235 (N_2235,N_2171,N_2095);
and U2236 (N_2236,N_2118,N_2077);
xor U2237 (N_2237,N_2092,N_2081);
or U2238 (N_2238,N_2164,N_2182);
xnor U2239 (N_2239,N_2068,N_2085);
nor U2240 (N_2240,N_2104,N_2133);
nand U2241 (N_2241,N_2089,N_2186);
or U2242 (N_2242,N_2001,N_2007);
nor U2243 (N_2243,N_2132,N_2097);
nor U2244 (N_2244,N_2127,N_2137);
xor U2245 (N_2245,N_2072,N_2031);
or U2246 (N_2246,N_2022,N_2070);
xnor U2247 (N_2247,N_2126,N_2011);
nor U2248 (N_2248,N_2017,N_2187);
nor U2249 (N_2249,N_2019,N_2055);
or U2250 (N_2250,N_2120,N_2195);
and U2251 (N_2251,N_2086,N_2087);
nor U2252 (N_2252,N_2071,N_2073);
nand U2253 (N_2253,N_2016,N_2173);
xnor U2254 (N_2254,N_2079,N_2033);
and U2255 (N_2255,N_2065,N_2138);
nand U2256 (N_2256,N_2160,N_2038);
nand U2257 (N_2257,N_2189,N_2048);
nand U2258 (N_2258,N_2145,N_2037);
or U2259 (N_2259,N_2149,N_2050);
nor U2260 (N_2260,N_2103,N_2003);
and U2261 (N_2261,N_2063,N_2099);
or U2262 (N_2262,N_2184,N_2183);
or U2263 (N_2263,N_2166,N_2172);
xor U2264 (N_2264,N_2040,N_2150);
nor U2265 (N_2265,N_2091,N_2084);
and U2266 (N_2266,N_2021,N_2052);
nor U2267 (N_2267,N_2167,N_2107);
xnor U2268 (N_2268,N_2075,N_2153);
or U2269 (N_2269,N_2032,N_2177);
nor U2270 (N_2270,N_2163,N_2193);
nand U2271 (N_2271,N_2054,N_2179);
nor U2272 (N_2272,N_2121,N_2174);
nor U2273 (N_2273,N_2131,N_2140);
or U2274 (N_2274,N_2136,N_2096);
or U2275 (N_2275,N_2191,N_2156);
and U2276 (N_2276,N_2057,N_2018);
and U2277 (N_2277,N_2110,N_2094);
or U2278 (N_2278,N_2147,N_2109);
xnor U2279 (N_2279,N_2006,N_2123);
and U2280 (N_2280,N_2045,N_2180);
or U2281 (N_2281,N_2042,N_2148);
nand U2282 (N_2282,N_2047,N_2199);
and U2283 (N_2283,N_2134,N_2088);
xnor U2284 (N_2284,N_2128,N_2152);
or U2285 (N_2285,N_2154,N_2124);
or U2286 (N_2286,N_2025,N_2122);
nand U2287 (N_2287,N_2143,N_2008);
xor U2288 (N_2288,N_2061,N_2036);
nand U2289 (N_2289,N_2108,N_2135);
nor U2290 (N_2290,N_2101,N_2116);
or U2291 (N_2291,N_2014,N_2159);
or U2292 (N_2292,N_2028,N_2012);
nand U2293 (N_2293,N_2069,N_2041);
and U2294 (N_2294,N_2020,N_2115);
xor U2295 (N_2295,N_2119,N_2188);
or U2296 (N_2296,N_2023,N_2190);
and U2297 (N_2297,N_2010,N_2112);
and U2298 (N_2298,N_2105,N_2125);
nor U2299 (N_2299,N_2165,N_2090);
or U2300 (N_2300,N_2044,N_2027);
xor U2301 (N_2301,N_2056,N_2148);
and U2302 (N_2302,N_2036,N_2183);
xnor U2303 (N_2303,N_2022,N_2046);
nand U2304 (N_2304,N_2185,N_2175);
xor U2305 (N_2305,N_2098,N_2103);
and U2306 (N_2306,N_2161,N_2184);
nor U2307 (N_2307,N_2016,N_2019);
nand U2308 (N_2308,N_2008,N_2169);
nand U2309 (N_2309,N_2121,N_2027);
or U2310 (N_2310,N_2022,N_2000);
nor U2311 (N_2311,N_2181,N_2124);
nor U2312 (N_2312,N_2010,N_2014);
nor U2313 (N_2313,N_2095,N_2130);
xor U2314 (N_2314,N_2136,N_2119);
or U2315 (N_2315,N_2111,N_2029);
xor U2316 (N_2316,N_2013,N_2104);
nand U2317 (N_2317,N_2081,N_2087);
or U2318 (N_2318,N_2160,N_2140);
or U2319 (N_2319,N_2068,N_2017);
or U2320 (N_2320,N_2101,N_2106);
nor U2321 (N_2321,N_2160,N_2166);
and U2322 (N_2322,N_2072,N_2000);
nand U2323 (N_2323,N_2025,N_2123);
xnor U2324 (N_2324,N_2030,N_2001);
xor U2325 (N_2325,N_2135,N_2192);
nor U2326 (N_2326,N_2037,N_2020);
nor U2327 (N_2327,N_2161,N_2033);
and U2328 (N_2328,N_2157,N_2162);
nor U2329 (N_2329,N_2123,N_2148);
nor U2330 (N_2330,N_2136,N_2090);
nor U2331 (N_2331,N_2184,N_2012);
nor U2332 (N_2332,N_2150,N_2165);
nand U2333 (N_2333,N_2117,N_2173);
xor U2334 (N_2334,N_2168,N_2028);
or U2335 (N_2335,N_2117,N_2120);
xor U2336 (N_2336,N_2179,N_2013);
nand U2337 (N_2337,N_2110,N_2195);
xnor U2338 (N_2338,N_2048,N_2045);
or U2339 (N_2339,N_2180,N_2070);
and U2340 (N_2340,N_2006,N_2199);
and U2341 (N_2341,N_2138,N_2191);
nand U2342 (N_2342,N_2174,N_2109);
and U2343 (N_2343,N_2152,N_2122);
nor U2344 (N_2344,N_2096,N_2126);
and U2345 (N_2345,N_2126,N_2127);
and U2346 (N_2346,N_2102,N_2073);
or U2347 (N_2347,N_2175,N_2032);
or U2348 (N_2348,N_2187,N_2070);
xnor U2349 (N_2349,N_2029,N_2069);
and U2350 (N_2350,N_2114,N_2090);
and U2351 (N_2351,N_2053,N_2064);
nor U2352 (N_2352,N_2181,N_2011);
nand U2353 (N_2353,N_2086,N_2114);
nor U2354 (N_2354,N_2018,N_2073);
nand U2355 (N_2355,N_2091,N_2199);
or U2356 (N_2356,N_2100,N_2050);
xnor U2357 (N_2357,N_2044,N_2110);
or U2358 (N_2358,N_2058,N_2052);
or U2359 (N_2359,N_2146,N_2049);
nor U2360 (N_2360,N_2032,N_2011);
nor U2361 (N_2361,N_2040,N_2105);
nor U2362 (N_2362,N_2180,N_2003);
xor U2363 (N_2363,N_2138,N_2024);
or U2364 (N_2364,N_2057,N_2194);
and U2365 (N_2365,N_2098,N_2044);
xor U2366 (N_2366,N_2135,N_2005);
nand U2367 (N_2367,N_2127,N_2111);
nand U2368 (N_2368,N_2022,N_2049);
and U2369 (N_2369,N_2139,N_2086);
or U2370 (N_2370,N_2028,N_2133);
nor U2371 (N_2371,N_2174,N_2020);
and U2372 (N_2372,N_2049,N_2137);
nand U2373 (N_2373,N_2174,N_2133);
xor U2374 (N_2374,N_2075,N_2057);
xnor U2375 (N_2375,N_2002,N_2004);
or U2376 (N_2376,N_2020,N_2165);
nor U2377 (N_2377,N_2102,N_2009);
nand U2378 (N_2378,N_2138,N_2167);
nand U2379 (N_2379,N_2104,N_2064);
and U2380 (N_2380,N_2160,N_2032);
or U2381 (N_2381,N_2073,N_2165);
xnor U2382 (N_2382,N_2062,N_2168);
xnor U2383 (N_2383,N_2170,N_2011);
nor U2384 (N_2384,N_2096,N_2058);
and U2385 (N_2385,N_2143,N_2148);
or U2386 (N_2386,N_2014,N_2060);
or U2387 (N_2387,N_2090,N_2096);
nor U2388 (N_2388,N_2165,N_2081);
xor U2389 (N_2389,N_2096,N_2067);
or U2390 (N_2390,N_2010,N_2066);
or U2391 (N_2391,N_2124,N_2017);
and U2392 (N_2392,N_2084,N_2050);
xnor U2393 (N_2393,N_2039,N_2043);
nand U2394 (N_2394,N_2039,N_2078);
nor U2395 (N_2395,N_2041,N_2115);
nor U2396 (N_2396,N_2084,N_2002);
or U2397 (N_2397,N_2014,N_2170);
or U2398 (N_2398,N_2160,N_2133);
and U2399 (N_2399,N_2093,N_2055);
nor U2400 (N_2400,N_2290,N_2324);
xnor U2401 (N_2401,N_2276,N_2389);
xor U2402 (N_2402,N_2213,N_2231);
nand U2403 (N_2403,N_2262,N_2329);
or U2404 (N_2404,N_2265,N_2327);
xor U2405 (N_2405,N_2310,N_2220);
or U2406 (N_2406,N_2342,N_2214);
xnor U2407 (N_2407,N_2201,N_2258);
xnor U2408 (N_2408,N_2367,N_2299);
or U2409 (N_2409,N_2234,N_2309);
and U2410 (N_2410,N_2316,N_2216);
nor U2411 (N_2411,N_2218,N_2243);
or U2412 (N_2412,N_2323,N_2311);
and U2413 (N_2413,N_2386,N_2289);
xnor U2414 (N_2414,N_2339,N_2259);
nand U2415 (N_2415,N_2352,N_2219);
or U2416 (N_2416,N_2224,N_2280);
or U2417 (N_2417,N_2306,N_2372);
xnor U2418 (N_2418,N_2206,N_2358);
and U2419 (N_2419,N_2221,N_2240);
and U2420 (N_2420,N_2254,N_2360);
or U2421 (N_2421,N_2350,N_2284);
nand U2422 (N_2422,N_2373,N_2287);
xnor U2423 (N_2423,N_2325,N_2361);
or U2424 (N_2424,N_2249,N_2236);
xnor U2425 (N_2425,N_2394,N_2272);
nor U2426 (N_2426,N_2237,N_2354);
xor U2427 (N_2427,N_2376,N_2229);
xnor U2428 (N_2428,N_2349,N_2378);
nand U2429 (N_2429,N_2371,N_2399);
nor U2430 (N_2430,N_2391,N_2283);
xor U2431 (N_2431,N_2331,N_2355);
and U2432 (N_2432,N_2314,N_2294);
nand U2433 (N_2433,N_2246,N_2322);
and U2434 (N_2434,N_2203,N_2281);
or U2435 (N_2435,N_2363,N_2307);
nand U2436 (N_2436,N_2387,N_2278);
xnor U2437 (N_2437,N_2225,N_2211);
nand U2438 (N_2438,N_2338,N_2270);
nor U2439 (N_2439,N_2321,N_2252);
nor U2440 (N_2440,N_2330,N_2318);
xor U2441 (N_2441,N_2359,N_2298);
nor U2442 (N_2442,N_2286,N_2362);
xnor U2443 (N_2443,N_2374,N_2343);
nand U2444 (N_2444,N_2257,N_2256);
nor U2445 (N_2445,N_2337,N_2244);
or U2446 (N_2446,N_2263,N_2313);
and U2447 (N_2447,N_2204,N_2296);
nor U2448 (N_2448,N_2304,N_2282);
xor U2449 (N_2449,N_2369,N_2388);
xnor U2450 (N_2450,N_2291,N_2266);
or U2451 (N_2451,N_2357,N_2348);
and U2452 (N_2452,N_2212,N_2390);
and U2453 (N_2453,N_2346,N_2381);
nand U2454 (N_2454,N_2293,N_2255);
xnor U2455 (N_2455,N_2353,N_2301);
nand U2456 (N_2456,N_2368,N_2217);
or U2457 (N_2457,N_2226,N_2279);
nand U2458 (N_2458,N_2334,N_2351);
and U2459 (N_2459,N_2300,N_2260);
nor U2460 (N_2460,N_2344,N_2332);
nor U2461 (N_2461,N_2379,N_2319);
nand U2462 (N_2462,N_2392,N_2210);
nand U2463 (N_2463,N_2317,N_2228);
nand U2464 (N_2464,N_2274,N_2275);
xnor U2465 (N_2465,N_2345,N_2297);
nand U2466 (N_2466,N_2207,N_2384);
or U2467 (N_2467,N_2380,N_2308);
nand U2468 (N_2468,N_2205,N_2326);
and U2469 (N_2469,N_2253,N_2365);
xor U2470 (N_2470,N_2232,N_2375);
xor U2471 (N_2471,N_2208,N_2285);
xnor U2472 (N_2472,N_2288,N_2340);
xnor U2473 (N_2473,N_2370,N_2328);
nor U2474 (N_2474,N_2242,N_2341);
xor U2475 (N_2475,N_2335,N_2312);
and U2476 (N_2476,N_2356,N_2238);
or U2477 (N_2477,N_2377,N_2267);
nand U2478 (N_2478,N_2333,N_2227);
or U2479 (N_2479,N_2302,N_2264);
xor U2480 (N_2480,N_2251,N_2295);
or U2481 (N_2481,N_2269,N_2239);
or U2482 (N_2482,N_2277,N_2347);
nand U2483 (N_2483,N_2396,N_2209);
nor U2484 (N_2484,N_2223,N_2261);
nor U2485 (N_2485,N_2235,N_2395);
nor U2486 (N_2486,N_2393,N_2222);
and U2487 (N_2487,N_2303,N_2383);
and U2488 (N_2488,N_2336,N_2273);
and U2489 (N_2489,N_2305,N_2215);
nor U2490 (N_2490,N_2320,N_2250);
nand U2491 (N_2491,N_2245,N_2233);
xor U2492 (N_2492,N_2200,N_2315);
nor U2493 (N_2493,N_2385,N_2397);
or U2494 (N_2494,N_2248,N_2271);
or U2495 (N_2495,N_2230,N_2292);
xnor U2496 (N_2496,N_2241,N_2398);
and U2497 (N_2497,N_2202,N_2268);
nand U2498 (N_2498,N_2364,N_2247);
xor U2499 (N_2499,N_2382,N_2366);
xnor U2500 (N_2500,N_2379,N_2334);
xnor U2501 (N_2501,N_2338,N_2209);
nor U2502 (N_2502,N_2346,N_2200);
nand U2503 (N_2503,N_2244,N_2335);
xor U2504 (N_2504,N_2299,N_2349);
and U2505 (N_2505,N_2213,N_2252);
and U2506 (N_2506,N_2336,N_2318);
and U2507 (N_2507,N_2214,N_2396);
or U2508 (N_2508,N_2366,N_2231);
or U2509 (N_2509,N_2285,N_2225);
nor U2510 (N_2510,N_2258,N_2237);
nand U2511 (N_2511,N_2351,N_2205);
xnor U2512 (N_2512,N_2395,N_2228);
nor U2513 (N_2513,N_2383,N_2391);
and U2514 (N_2514,N_2204,N_2205);
xnor U2515 (N_2515,N_2231,N_2206);
or U2516 (N_2516,N_2353,N_2298);
nand U2517 (N_2517,N_2394,N_2238);
nor U2518 (N_2518,N_2259,N_2301);
nor U2519 (N_2519,N_2304,N_2348);
nor U2520 (N_2520,N_2343,N_2334);
or U2521 (N_2521,N_2250,N_2296);
nand U2522 (N_2522,N_2242,N_2262);
xor U2523 (N_2523,N_2353,N_2215);
xnor U2524 (N_2524,N_2276,N_2214);
or U2525 (N_2525,N_2218,N_2351);
xnor U2526 (N_2526,N_2283,N_2275);
nand U2527 (N_2527,N_2316,N_2224);
or U2528 (N_2528,N_2377,N_2312);
or U2529 (N_2529,N_2360,N_2301);
nor U2530 (N_2530,N_2347,N_2271);
xnor U2531 (N_2531,N_2241,N_2252);
nand U2532 (N_2532,N_2300,N_2211);
or U2533 (N_2533,N_2288,N_2241);
nand U2534 (N_2534,N_2261,N_2207);
xnor U2535 (N_2535,N_2309,N_2205);
xnor U2536 (N_2536,N_2215,N_2278);
nor U2537 (N_2537,N_2229,N_2335);
and U2538 (N_2538,N_2254,N_2387);
or U2539 (N_2539,N_2372,N_2341);
xnor U2540 (N_2540,N_2219,N_2223);
nor U2541 (N_2541,N_2363,N_2369);
nor U2542 (N_2542,N_2348,N_2261);
or U2543 (N_2543,N_2382,N_2286);
nand U2544 (N_2544,N_2350,N_2224);
nor U2545 (N_2545,N_2372,N_2291);
or U2546 (N_2546,N_2349,N_2301);
xor U2547 (N_2547,N_2366,N_2260);
xor U2548 (N_2548,N_2376,N_2325);
and U2549 (N_2549,N_2276,N_2273);
nor U2550 (N_2550,N_2270,N_2369);
or U2551 (N_2551,N_2361,N_2336);
nor U2552 (N_2552,N_2291,N_2225);
nand U2553 (N_2553,N_2333,N_2366);
xor U2554 (N_2554,N_2334,N_2275);
xor U2555 (N_2555,N_2390,N_2358);
or U2556 (N_2556,N_2390,N_2326);
nand U2557 (N_2557,N_2347,N_2350);
or U2558 (N_2558,N_2227,N_2264);
nor U2559 (N_2559,N_2392,N_2207);
and U2560 (N_2560,N_2281,N_2398);
nor U2561 (N_2561,N_2334,N_2256);
and U2562 (N_2562,N_2330,N_2226);
and U2563 (N_2563,N_2386,N_2316);
xor U2564 (N_2564,N_2344,N_2317);
and U2565 (N_2565,N_2308,N_2245);
or U2566 (N_2566,N_2255,N_2307);
nor U2567 (N_2567,N_2308,N_2357);
nand U2568 (N_2568,N_2369,N_2348);
nor U2569 (N_2569,N_2378,N_2294);
nor U2570 (N_2570,N_2378,N_2205);
nor U2571 (N_2571,N_2263,N_2372);
nor U2572 (N_2572,N_2363,N_2375);
and U2573 (N_2573,N_2368,N_2235);
nand U2574 (N_2574,N_2273,N_2200);
or U2575 (N_2575,N_2368,N_2392);
xnor U2576 (N_2576,N_2222,N_2242);
xor U2577 (N_2577,N_2237,N_2350);
or U2578 (N_2578,N_2368,N_2365);
nor U2579 (N_2579,N_2247,N_2330);
xnor U2580 (N_2580,N_2356,N_2241);
xor U2581 (N_2581,N_2268,N_2308);
nand U2582 (N_2582,N_2247,N_2323);
xnor U2583 (N_2583,N_2266,N_2397);
or U2584 (N_2584,N_2396,N_2228);
xnor U2585 (N_2585,N_2356,N_2230);
nand U2586 (N_2586,N_2205,N_2250);
nand U2587 (N_2587,N_2202,N_2309);
xnor U2588 (N_2588,N_2289,N_2383);
nand U2589 (N_2589,N_2377,N_2232);
xor U2590 (N_2590,N_2313,N_2334);
and U2591 (N_2591,N_2243,N_2227);
or U2592 (N_2592,N_2261,N_2297);
or U2593 (N_2593,N_2281,N_2224);
and U2594 (N_2594,N_2263,N_2357);
or U2595 (N_2595,N_2229,N_2395);
and U2596 (N_2596,N_2328,N_2268);
nor U2597 (N_2597,N_2215,N_2311);
and U2598 (N_2598,N_2373,N_2363);
or U2599 (N_2599,N_2341,N_2378);
and U2600 (N_2600,N_2528,N_2437);
nand U2601 (N_2601,N_2511,N_2571);
xor U2602 (N_2602,N_2548,N_2584);
or U2603 (N_2603,N_2443,N_2538);
nand U2604 (N_2604,N_2568,N_2411);
nand U2605 (N_2605,N_2522,N_2462);
or U2606 (N_2606,N_2525,N_2553);
or U2607 (N_2607,N_2409,N_2434);
nand U2608 (N_2608,N_2527,N_2576);
and U2609 (N_2609,N_2408,N_2578);
and U2610 (N_2610,N_2467,N_2581);
nand U2611 (N_2611,N_2559,N_2587);
or U2612 (N_2612,N_2593,N_2509);
or U2613 (N_2613,N_2476,N_2418);
and U2614 (N_2614,N_2540,N_2585);
xor U2615 (N_2615,N_2543,N_2510);
nor U2616 (N_2616,N_2554,N_2499);
and U2617 (N_2617,N_2478,N_2465);
xor U2618 (N_2618,N_2452,N_2574);
or U2619 (N_2619,N_2401,N_2419);
xnor U2620 (N_2620,N_2454,N_2561);
nor U2621 (N_2621,N_2402,N_2557);
nor U2622 (N_2622,N_2479,N_2442);
xnor U2623 (N_2623,N_2506,N_2531);
nand U2624 (N_2624,N_2426,N_2507);
xor U2625 (N_2625,N_2451,N_2498);
nor U2626 (N_2626,N_2404,N_2450);
or U2627 (N_2627,N_2445,N_2589);
nor U2628 (N_2628,N_2466,N_2423);
xor U2629 (N_2629,N_2539,N_2513);
xor U2630 (N_2630,N_2551,N_2523);
and U2631 (N_2631,N_2432,N_2524);
nor U2632 (N_2632,N_2542,N_2471);
xor U2633 (N_2633,N_2563,N_2517);
nand U2634 (N_2634,N_2429,N_2458);
nor U2635 (N_2635,N_2449,N_2562);
and U2636 (N_2636,N_2470,N_2552);
xor U2637 (N_2637,N_2537,N_2516);
and U2638 (N_2638,N_2406,N_2438);
and U2639 (N_2639,N_2586,N_2564);
or U2640 (N_2640,N_2422,N_2530);
xor U2641 (N_2641,N_2541,N_2459);
or U2642 (N_2642,N_2424,N_2415);
or U2643 (N_2643,N_2456,N_2405);
and U2644 (N_2644,N_2484,N_2591);
xnor U2645 (N_2645,N_2472,N_2403);
nor U2646 (N_2646,N_2461,N_2446);
xnor U2647 (N_2647,N_2535,N_2504);
or U2648 (N_2648,N_2582,N_2428);
nor U2649 (N_2649,N_2491,N_2444);
xnor U2650 (N_2650,N_2529,N_2463);
nor U2651 (N_2651,N_2453,N_2549);
or U2652 (N_2652,N_2457,N_2421);
nand U2653 (N_2653,N_2569,N_2505);
nand U2654 (N_2654,N_2495,N_2448);
nand U2655 (N_2655,N_2514,N_2414);
nor U2656 (N_2656,N_2447,N_2433);
nand U2657 (N_2657,N_2469,N_2425);
or U2658 (N_2658,N_2580,N_2435);
nor U2659 (N_2659,N_2481,N_2420);
and U2660 (N_2660,N_2521,N_2489);
xnor U2661 (N_2661,N_2566,N_2413);
nor U2662 (N_2662,N_2407,N_2590);
nand U2663 (N_2663,N_2594,N_2595);
nand U2664 (N_2664,N_2497,N_2598);
or U2665 (N_2665,N_2441,N_2492);
or U2666 (N_2666,N_2485,N_2500);
or U2667 (N_2667,N_2494,N_2464);
nor U2668 (N_2668,N_2477,N_2460);
nand U2669 (N_2669,N_2502,N_2567);
nor U2670 (N_2670,N_2490,N_2534);
xor U2671 (N_2671,N_2592,N_2544);
or U2672 (N_2672,N_2496,N_2475);
nand U2673 (N_2673,N_2430,N_2588);
nor U2674 (N_2674,N_2455,N_2596);
or U2675 (N_2675,N_2488,N_2487);
or U2676 (N_2676,N_2572,N_2546);
nand U2677 (N_2677,N_2519,N_2431);
nor U2678 (N_2678,N_2482,N_2565);
and U2679 (N_2679,N_2573,N_2493);
xnor U2680 (N_2680,N_2550,N_2545);
nand U2681 (N_2681,N_2579,N_2558);
xor U2682 (N_2682,N_2555,N_2439);
or U2683 (N_2683,N_2577,N_2503);
or U2684 (N_2684,N_2512,N_2427);
nand U2685 (N_2685,N_2518,N_2412);
and U2686 (N_2686,N_2400,N_2570);
xor U2687 (N_2687,N_2508,N_2416);
nand U2688 (N_2688,N_2440,N_2480);
and U2689 (N_2689,N_2436,N_2526);
nor U2690 (N_2690,N_2486,N_2473);
and U2691 (N_2691,N_2597,N_2468);
xor U2692 (N_2692,N_2560,N_2599);
nand U2693 (N_2693,N_2547,N_2532);
or U2694 (N_2694,N_2583,N_2417);
nor U2695 (N_2695,N_2520,N_2575);
nand U2696 (N_2696,N_2483,N_2533);
xor U2697 (N_2697,N_2501,N_2556);
xor U2698 (N_2698,N_2474,N_2536);
nand U2699 (N_2699,N_2515,N_2410);
xor U2700 (N_2700,N_2484,N_2463);
nor U2701 (N_2701,N_2464,N_2531);
or U2702 (N_2702,N_2576,N_2459);
or U2703 (N_2703,N_2586,N_2540);
and U2704 (N_2704,N_2535,N_2531);
nand U2705 (N_2705,N_2509,N_2461);
xnor U2706 (N_2706,N_2587,N_2448);
and U2707 (N_2707,N_2416,N_2586);
nand U2708 (N_2708,N_2570,N_2561);
or U2709 (N_2709,N_2581,N_2512);
nor U2710 (N_2710,N_2448,N_2443);
nand U2711 (N_2711,N_2528,N_2401);
or U2712 (N_2712,N_2505,N_2513);
or U2713 (N_2713,N_2505,N_2428);
or U2714 (N_2714,N_2471,N_2548);
nand U2715 (N_2715,N_2445,N_2501);
xnor U2716 (N_2716,N_2537,N_2599);
xor U2717 (N_2717,N_2575,N_2582);
nand U2718 (N_2718,N_2452,N_2431);
nand U2719 (N_2719,N_2588,N_2531);
and U2720 (N_2720,N_2452,N_2505);
nand U2721 (N_2721,N_2494,N_2528);
nor U2722 (N_2722,N_2437,N_2501);
or U2723 (N_2723,N_2475,N_2470);
and U2724 (N_2724,N_2496,N_2474);
or U2725 (N_2725,N_2438,N_2540);
xnor U2726 (N_2726,N_2571,N_2585);
xor U2727 (N_2727,N_2532,N_2504);
nor U2728 (N_2728,N_2477,N_2474);
and U2729 (N_2729,N_2469,N_2446);
nand U2730 (N_2730,N_2412,N_2511);
or U2731 (N_2731,N_2549,N_2475);
or U2732 (N_2732,N_2486,N_2514);
nand U2733 (N_2733,N_2544,N_2431);
nand U2734 (N_2734,N_2431,N_2426);
nand U2735 (N_2735,N_2506,N_2453);
xor U2736 (N_2736,N_2595,N_2496);
and U2737 (N_2737,N_2498,N_2427);
nand U2738 (N_2738,N_2425,N_2432);
or U2739 (N_2739,N_2471,N_2497);
or U2740 (N_2740,N_2457,N_2415);
xor U2741 (N_2741,N_2411,N_2509);
nor U2742 (N_2742,N_2468,N_2494);
nor U2743 (N_2743,N_2475,N_2431);
and U2744 (N_2744,N_2543,N_2563);
or U2745 (N_2745,N_2526,N_2490);
nor U2746 (N_2746,N_2511,N_2402);
and U2747 (N_2747,N_2471,N_2596);
and U2748 (N_2748,N_2592,N_2545);
and U2749 (N_2749,N_2436,N_2518);
nand U2750 (N_2750,N_2447,N_2549);
and U2751 (N_2751,N_2542,N_2544);
nor U2752 (N_2752,N_2500,N_2421);
and U2753 (N_2753,N_2410,N_2536);
nor U2754 (N_2754,N_2550,N_2470);
xnor U2755 (N_2755,N_2471,N_2432);
nand U2756 (N_2756,N_2455,N_2493);
nand U2757 (N_2757,N_2580,N_2528);
nor U2758 (N_2758,N_2499,N_2539);
xor U2759 (N_2759,N_2564,N_2450);
nand U2760 (N_2760,N_2511,N_2582);
nand U2761 (N_2761,N_2533,N_2422);
or U2762 (N_2762,N_2598,N_2417);
or U2763 (N_2763,N_2593,N_2536);
nor U2764 (N_2764,N_2576,N_2443);
and U2765 (N_2765,N_2578,N_2488);
and U2766 (N_2766,N_2419,N_2507);
or U2767 (N_2767,N_2480,N_2547);
nor U2768 (N_2768,N_2497,N_2480);
or U2769 (N_2769,N_2584,N_2408);
and U2770 (N_2770,N_2416,N_2400);
or U2771 (N_2771,N_2581,N_2533);
xnor U2772 (N_2772,N_2448,N_2469);
xnor U2773 (N_2773,N_2441,N_2474);
or U2774 (N_2774,N_2509,N_2588);
xnor U2775 (N_2775,N_2442,N_2494);
or U2776 (N_2776,N_2485,N_2467);
nor U2777 (N_2777,N_2538,N_2431);
or U2778 (N_2778,N_2544,N_2565);
xor U2779 (N_2779,N_2429,N_2468);
and U2780 (N_2780,N_2560,N_2527);
and U2781 (N_2781,N_2490,N_2528);
and U2782 (N_2782,N_2574,N_2451);
or U2783 (N_2783,N_2481,N_2587);
nor U2784 (N_2784,N_2547,N_2417);
or U2785 (N_2785,N_2599,N_2413);
or U2786 (N_2786,N_2436,N_2450);
or U2787 (N_2787,N_2469,N_2519);
or U2788 (N_2788,N_2439,N_2411);
and U2789 (N_2789,N_2515,N_2486);
and U2790 (N_2790,N_2424,N_2500);
nand U2791 (N_2791,N_2592,N_2583);
or U2792 (N_2792,N_2543,N_2518);
xnor U2793 (N_2793,N_2507,N_2479);
and U2794 (N_2794,N_2544,N_2545);
nor U2795 (N_2795,N_2477,N_2458);
xnor U2796 (N_2796,N_2524,N_2493);
nand U2797 (N_2797,N_2592,N_2561);
xnor U2798 (N_2798,N_2435,N_2534);
and U2799 (N_2799,N_2585,N_2531);
nand U2800 (N_2800,N_2793,N_2645);
xnor U2801 (N_2801,N_2628,N_2634);
or U2802 (N_2802,N_2664,N_2659);
nor U2803 (N_2803,N_2684,N_2762);
and U2804 (N_2804,N_2785,N_2792);
or U2805 (N_2805,N_2739,N_2721);
xor U2806 (N_2806,N_2781,N_2641);
nor U2807 (N_2807,N_2661,N_2741);
xnor U2808 (N_2808,N_2644,N_2668);
nand U2809 (N_2809,N_2600,N_2643);
or U2810 (N_2810,N_2700,N_2677);
nor U2811 (N_2811,N_2795,N_2673);
or U2812 (N_2812,N_2611,N_2758);
nand U2813 (N_2813,N_2605,N_2743);
xnor U2814 (N_2814,N_2799,N_2618);
xnor U2815 (N_2815,N_2724,N_2732);
and U2816 (N_2816,N_2658,N_2748);
and U2817 (N_2817,N_2614,N_2697);
nor U2818 (N_2818,N_2728,N_2679);
or U2819 (N_2819,N_2610,N_2756);
or U2820 (N_2820,N_2609,N_2654);
nor U2821 (N_2821,N_2716,N_2760);
or U2822 (N_2822,N_2722,N_2776);
nor U2823 (N_2823,N_2685,N_2798);
and U2824 (N_2824,N_2742,N_2624);
or U2825 (N_2825,N_2759,N_2620);
or U2826 (N_2826,N_2660,N_2649);
xor U2827 (N_2827,N_2653,N_2681);
and U2828 (N_2828,N_2601,N_2630);
or U2829 (N_2829,N_2784,N_2692);
xor U2830 (N_2830,N_2791,N_2735);
or U2831 (N_2831,N_2655,N_2687);
xor U2832 (N_2832,N_2694,N_2637);
or U2833 (N_2833,N_2638,N_2733);
or U2834 (N_2834,N_2780,N_2767);
nor U2835 (N_2835,N_2725,N_2777);
and U2836 (N_2836,N_2744,N_2757);
nand U2837 (N_2837,N_2662,N_2730);
xnor U2838 (N_2838,N_2773,N_2670);
or U2839 (N_2839,N_2755,N_2640);
or U2840 (N_2840,N_2678,N_2752);
xor U2841 (N_2841,N_2627,N_2714);
nor U2842 (N_2842,N_2626,N_2604);
xor U2843 (N_2843,N_2676,N_2686);
xnor U2844 (N_2844,N_2667,N_2698);
nand U2845 (N_2845,N_2603,N_2656);
nand U2846 (N_2846,N_2726,N_2729);
xor U2847 (N_2847,N_2671,N_2608);
and U2848 (N_2848,N_2613,N_2727);
or U2849 (N_2849,N_2633,N_2717);
xor U2850 (N_2850,N_2736,N_2619);
nand U2851 (N_2851,N_2657,N_2769);
xnor U2852 (N_2852,N_2734,N_2771);
nor U2853 (N_2853,N_2650,N_2699);
xor U2854 (N_2854,N_2751,N_2674);
nor U2855 (N_2855,N_2647,N_2768);
and U2856 (N_2856,N_2711,N_2710);
nand U2857 (N_2857,N_2753,N_2616);
nand U2858 (N_2858,N_2754,N_2705);
or U2859 (N_2859,N_2715,N_2689);
xnor U2860 (N_2860,N_2690,N_2783);
nor U2861 (N_2861,N_2696,N_2693);
xor U2862 (N_2862,N_2788,N_2607);
nor U2863 (N_2863,N_2602,N_2629);
nor U2864 (N_2864,N_2625,N_2770);
and U2865 (N_2865,N_2720,N_2615);
xor U2866 (N_2866,N_2636,N_2761);
nand U2867 (N_2867,N_2790,N_2797);
nand U2868 (N_2868,N_2713,N_2680);
and U2869 (N_2869,N_2606,N_2709);
nor U2870 (N_2870,N_2731,N_2648);
and U2871 (N_2871,N_2622,N_2632);
or U2872 (N_2872,N_2688,N_2663);
xor U2873 (N_2873,N_2701,N_2639);
xnor U2874 (N_2874,N_2738,N_2621);
or U2875 (N_2875,N_2737,N_2750);
and U2876 (N_2876,N_2712,N_2703);
xnor U2877 (N_2877,N_2775,N_2612);
and U2878 (N_2878,N_2789,N_2651);
nor U2879 (N_2879,N_2746,N_2623);
and U2880 (N_2880,N_2772,N_2691);
nor U2881 (N_2881,N_2675,N_2766);
and U2882 (N_2882,N_2672,N_2707);
xor U2883 (N_2883,N_2794,N_2723);
or U2884 (N_2884,N_2635,N_2763);
nand U2885 (N_2885,N_2749,N_2782);
or U2886 (N_2886,N_2740,N_2719);
and U2887 (N_2887,N_2747,N_2745);
nand U2888 (N_2888,N_2666,N_2642);
and U2889 (N_2889,N_2764,N_2704);
nor U2890 (N_2890,N_2774,N_2718);
and U2891 (N_2891,N_2787,N_2646);
xor U2892 (N_2892,N_2708,N_2702);
or U2893 (N_2893,N_2682,N_2778);
or U2894 (N_2894,N_2652,N_2669);
nor U2895 (N_2895,N_2796,N_2706);
xnor U2896 (N_2896,N_2779,N_2765);
xnor U2897 (N_2897,N_2665,N_2631);
nor U2898 (N_2898,N_2617,N_2695);
or U2899 (N_2899,N_2786,N_2683);
or U2900 (N_2900,N_2650,N_2721);
xnor U2901 (N_2901,N_2652,N_2677);
or U2902 (N_2902,N_2600,N_2708);
nand U2903 (N_2903,N_2603,N_2714);
xnor U2904 (N_2904,N_2773,N_2744);
nor U2905 (N_2905,N_2699,N_2758);
or U2906 (N_2906,N_2707,N_2709);
or U2907 (N_2907,N_2652,N_2746);
xor U2908 (N_2908,N_2608,N_2733);
and U2909 (N_2909,N_2601,N_2712);
xnor U2910 (N_2910,N_2614,N_2689);
xnor U2911 (N_2911,N_2603,N_2792);
xor U2912 (N_2912,N_2612,N_2610);
nand U2913 (N_2913,N_2729,N_2625);
nand U2914 (N_2914,N_2674,N_2604);
and U2915 (N_2915,N_2603,N_2750);
xor U2916 (N_2916,N_2715,N_2605);
and U2917 (N_2917,N_2665,N_2638);
nor U2918 (N_2918,N_2799,N_2686);
xnor U2919 (N_2919,N_2778,N_2624);
or U2920 (N_2920,N_2790,N_2658);
nor U2921 (N_2921,N_2605,N_2717);
or U2922 (N_2922,N_2779,N_2730);
or U2923 (N_2923,N_2711,N_2641);
nor U2924 (N_2924,N_2750,N_2789);
xnor U2925 (N_2925,N_2712,N_2628);
or U2926 (N_2926,N_2637,N_2704);
or U2927 (N_2927,N_2745,N_2743);
xor U2928 (N_2928,N_2612,N_2763);
and U2929 (N_2929,N_2668,N_2760);
nand U2930 (N_2930,N_2725,N_2703);
or U2931 (N_2931,N_2788,N_2680);
xor U2932 (N_2932,N_2704,N_2788);
or U2933 (N_2933,N_2684,N_2666);
nand U2934 (N_2934,N_2743,N_2627);
nor U2935 (N_2935,N_2757,N_2762);
nor U2936 (N_2936,N_2674,N_2786);
nand U2937 (N_2937,N_2638,N_2623);
and U2938 (N_2938,N_2701,N_2605);
or U2939 (N_2939,N_2709,N_2608);
xor U2940 (N_2940,N_2710,N_2686);
nand U2941 (N_2941,N_2654,N_2644);
and U2942 (N_2942,N_2755,N_2764);
xnor U2943 (N_2943,N_2609,N_2718);
xor U2944 (N_2944,N_2718,N_2607);
or U2945 (N_2945,N_2696,N_2625);
and U2946 (N_2946,N_2751,N_2784);
and U2947 (N_2947,N_2640,N_2798);
and U2948 (N_2948,N_2768,N_2787);
nand U2949 (N_2949,N_2695,N_2608);
xnor U2950 (N_2950,N_2697,N_2738);
xor U2951 (N_2951,N_2783,N_2679);
nand U2952 (N_2952,N_2609,N_2705);
nor U2953 (N_2953,N_2781,N_2770);
xor U2954 (N_2954,N_2657,N_2716);
xnor U2955 (N_2955,N_2601,N_2603);
and U2956 (N_2956,N_2792,N_2793);
and U2957 (N_2957,N_2797,N_2771);
or U2958 (N_2958,N_2608,N_2622);
nand U2959 (N_2959,N_2759,N_2692);
and U2960 (N_2960,N_2681,N_2744);
or U2961 (N_2961,N_2673,N_2637);
or U2962 (N_2962,N_2715,N_2779);
xor U2963 (N_2963,N_2717,N_2797);
nand U2964 (N_2964,N_2705,N_2629);
xor U2965 (N_2965,N_2791,N_2624);
or U2966 (N_2966,N_2626,N_2668);
or U2967 (N_2967,N_2623,N_2709);
and U2968 (N_2968,N_2601,N_2719);
and U2969 (N_2969,N_2719,N_2613);
xor U2970 (N_2970,N_2610,N_2748);
or U2971 (N_2971,N_2784,N_2752);
and U2972 (N_2972,N_2749,N_2747);
nand U2973 (N_2973,N_2701,N_2633);
and U2974 (N_2974,N_2725,N_2651);
and U2975 (N_2975,N_2732,N_2741);
nor U2976 (N_2976,N_2799,N_2728);
xnor U2977 (N_2977,N_2630,N_2634);
or U2978 (N_2978,N_2635,N_2633);
nor U2979 (N_2979,N_2664,N_2687);
nor U2980 (N_2980,N_2609,N_2622);
nor U2981 (N_2981,N_2727,N_2797);
nor U2982 (N_2982,N_2676,N_2698);
and U2983 (N_2983,N_2657,N_2676);
or U2984 (N_2984,N_2744,N_2775);
or U2985 (N_2985,N_2729,N_2652);
or U2986 (N_2986,N_2666,N_2663);
xnor U2987 (N_2987,N_2729,N_2612);
xor U2988 (N_2988,N_2630,N_2754);
and U2989 (N_2989,N_2670,N_2625);
nand U2990 (N_2990,N_2640,N_2723);
nand U2991 (N_2991,N_2742,N_2685);
xor U2992 (N_2992,N_2720,N_2665);
or U2993 (N_2993,N_2764,N_2630);
and U2994 (N_2994,N_2779,N_2720);
xnor U2995 (N_2995,N_2623,N_2624);
nor U2996 (N_2996,N_2718,N_2700);
or U2997 (N_2997,N_2622,N_2728);
nand U2998 (N_2998,N_2729,N_2748);
nand U2999 (N_2999,N_2641,N_2793);
nor U3000 (N_3000,N_2969,N_2936);
or U3001 (N_3001,N_2951,N_2825);
nand U3002 (N_3002,N_2918,N_2865);
or U3003 (N_3003,N_2927,N_2888);
and U3004 (N_3004,N_2805,N_2988);
nand U3005 (N_3005,N_2948,N_2922);
nand U3006 (N_3006,N_2998,N_2989);
and U3007 (N_3007,N_2987,N_2923);
nor U3008 (N_3008,N_2855,N_2968);
nand U3009 (N_3009,N_2894,N_2934);
xor U3010 (N_3010,N_2991,N_2824);
or U3011 (N_3011,N_2812,N_2992);
nand U3012 (N_3012,N_2958,N_2952);
xnor U3013 (N_3013,N_2833,N_2841);
or U3014 (N_3014,N_2975,N_2947);
or U3015 (N_3015,N_2806,N_2950);
nand U3016 (N_3016,N_2878,N_2877);
nor U3017 (N_3017,N_2837,N_2827);
or U3018 (N_3018,N_2859,N_2884);
or U3019 (N_3019,N_2895,N_2817);
xor U3020 (N_3020,N_2974,N_2960);
xor U3021 (N_3021,N_2835,N_2816);
nand U3022 (N_3022,N_2866,N_2818);
nand U3023 (N_3023,N_2996,N_2813);
xnor U3024 (N_3024,N_2967,N_2857);
xnor U3025 (N_3025,N_2915,N_2963);
nor U3026 (N_3026,N_2905,N_2871);
or U3027 (N_3027,N_2867,N_2932);
or U3028 (N_3028,N_2800,N_2851);
nand U3029 (N_3029,N_2885,N_2807);
and U3030 (N_3030,N_2940,N_2848);
nand U3031 (N_3031,N_2902,N_2852);
nor U3032 (N_3032,N_2869,N_2803);
and U3033 (N_3033,N_2836,N_2946);
xor U3034 (N_3034,N_2929,N_2804);
nor U3035 (N_3035,N_2875,N_2868);
or U3036 (N_3036,N_2826,N_2994);
or U3037 (N_3037,N_2935,N_2928);
or U3038 (N_3038,N_2891,N_2986);
xnor U3039 (N_3039,N_2815,N_2930);
or U3040 (N_3040,N_2924,N_2844);
and U3041 (N_3041,N_2966,N_2858);
nand U3042 (N_3042,N_2962,N_2830);
nand U3043 (N_3043,N_2889,N_2901);
or U3044 (N_3044,N_2839,N_2912);
nand U3045 (N_3045,N_2876,N_2984);
xnor U3046 (N_3046,N_2870,N_2897);
xor U3047 (N_3047,N_2979,N_2890);
or U3048 (N_3048,N_2997,N_2913);
xnor U3049 (N_3049,N_2917,N_2823);
and U3050 (N_3050,N_2846,N_2971);
xnor U3051 (N_3051,N_2849,N_2945);
and U3052 (N_3052,N_2937,N_2909);
or U3053 (N_3053,N_2943,N_2821);
nand U3054 (N_3054,N_2903,N_2944);
xnor U3055 (N_3055,N_2842,N_2938);
xor U3056 (N_3056,N_2801,N_2972);
nor U3057 (N_3057,N_2896,N_2886);
nand U3058 (N_3058,N_2862,N_2955);
or U3059 (N_3059,N_2976,N_2808);
nor U3060 (N_3060,N_2985,N_2879);
nor U3061 (N_3061,N_2953,N_2925);
xnor U3062 (N_3062,N_2850,N_2983);
xor U3063 (N_3063,N_2882,N_2847);
nor U3064 (N_3064,N_2853,N_2904);
nor U3065 (N_3065,N_2961,N_2980);
or U3066 (N_3066,N_2977,N_2907);
nand U3067 (N_3067,N_2820,N_2829);
nor U3068 (N_3068,N_2995,N_2861);
nor U3069 (N_3069,N_2814,N_2811);
xor U3070 (N_3070,N_2910,N_2864);
nand U3071 (N_3071,N_2810,N_2957);
xor U3072 (N_3072,N_2819,N_2802);
or U3073 (N_3073,N_2834,N_2892);
nand U3074 (N_3074,N_2881,N_2911);
xor U3075 (N_3075,N_2874,N_2973);
xor U3076 (N_3076,N_2956,N_2838);
nand U3077 (N_3077,N_2873,N_2880);
nor U3078 (N_3078,N_2993,N_2900);
or U3079 (N_3079,N_2939,N_2970);
or U3080 (N_3080,N_2965,N_2831);
xor U3081 (N_3081,N_2920,N_2845);
nand U3082 (N_3082,N_2899,N_2914);
nand U3083 (N_3083,N_2964,N_2872);
and U3084 (N_3084,N_2982,N_2840);
and U3085 (N_3085,N_2822,N_2916);
nor U3086 (N_3086,N_2887,N_2854);
nor U3087 (N_3087,N_2921,N_2959);
nand U3088 (N_3088,N_2919,N_2893);
xnor U3089 (N_3089,N_2843,N_2978);
and U3090 (N_3090,N_2926,N_2856);
or U3091 (N_3091,N_2931,N_2954);
or U3092 (N_3092,N_2898,N_2933);
nand U3093 (N_3093,N_2941,N_2999);
nand U3094 (N_3094,N_2828,N_2832);
xor U3095 (N_3095,N_2863,N_2906);
xnor U3096 (N_3096,N_2942,N_2809);
and U3097 (N_3097,N_2949,N_2883);
nand U3098 (N_3098,N_2860,N_2990);
nand U3099 (N_3099,N_2981,N_2908);
nand U3100 (N_3100,N_2969,N_2959);
xor U3101 (N_3101,N_2996,N_2894);
nor U3102 (N_3102,N_2923,N_2972);
xor U3103 (N_3103,N_2970,N_2903);
nor U3104 (N_3104,N_2862,N_2881);
or U3105 (N_3105,N_2854,N_2901);
xor U3106 (N_3106,N_2857,N_2825);
nor U3107 (N_3107,N_2905,N_2940);
and U3108 (N_3108,N_2934,N_2856);
nand U3109 (N_3109,N_2950,N_2890);
nand U3110 (N_3110,N_2921,N_2989);
xor U3111 (N_3111,N_2907,N_2965);
nor U3112 (N_3112,N_2976,N_2946);
xor U3113 (N_3113,N_2959,N_2972);
or U3114 (N_3114,N_2921,N_2965);
xnor U3115 (N_3115,N_2915,N_2856);
xnor U3116 (N_3116,N_2825,N_2990);
or U3117 (N_3117,N_2806,N_2865);
nor U3118 (N_3118,N_2914,N_2947);
nor U3119 (N_3119,N_2998,N_2823);
nand U3120 (N_3120,N_2917,N_2804);
xnor U3121 (N_3121,N_2838,N_2968);
nor U3122 (N_3122,N_2939,N_2816);
and U3123 (N_3123,N_2955,N_2924);
xor U3124 (N_3124,N_2924,N_2887);
xor U3125 (N_3125,N_2929,N_2847);
and U3126 (N_3126,N_2940,N_2935);
nor U3127 (N_3127,N_2863,N_2956);
or U3128 (N_3128,N_2893,N_2825);
or U3129 (N_3129,N_2987,N_2952);
or U3130 (N_3130,N_2954,N_2879);
or U3131 (N_3131,N_2957,N_2804);
nor U3132 (N_3132,N_2957,N_2855);
nor U3133 (N_3133,N_2937,N_2904);
nand U3134 (N_3134,N_2966,N_2903);
xnor U3135 (N_3135,N_2932,N_2822);
and U3136 (N_3136,N_2846,N_2881);
nor U3137 (N_3137,N_2901,N_2982);
xnor U3138 (N_3138,N_2980,N_2865);
and U3139 (N_3139,N_2967,N_2929);
xor U3140 (N_3140,N_2953,N_2903);
or U3141 (N_3141,N_2973,N_2961);
xor U3142 (N_3142,N_2883,N_2817);
nand U3143 (N_3143,N_2902,N_2871);
nor U3144 (N_3144,N_2877,N_2870);
nor U3145 (N_3145,N_2837,N_2816);
nor U3146 (N_3146,N_2926,N_2997);
xnor U3147 (N_3147,N_2924,N_2903);
or U3148 (N_3148,N_2835,N_2962);
or U3149 (N_3149,N_2871,N_2878);
and U3150 (N_3150,N_2991,N_2868);
nor U3151 (N_3151,N_2870,N_2999);
or U3152 (N_3152,N_2957,N_2964);
and U3153 (N_3153,N_2843,N_2962);
and U3154 (N_3154,N_2816,N_2885);
nand U3155 (N_3155,N_2978,N_2839);
and U3156 (N_3156,N_2816,N_2824);
and U3157 (N_3157,N_2916,N_2989);
or U3158 (N_3158,N_2925,N_2802);
nor U3159 (N_3159,N_2990,N_2932);
and U3160 (N_3160,N_2959,N_2890);
nor U3161 (N_3161,N_2934,N_2956);
nand U3162 (N_3162,N_2970,N_2830);
or U3163 (N_3163,N_2999,N_2806);
nor U3164 (N_3164,N_2839,N_2865);
or U3165 (N_3165,N_2847,N_2987);
xor U3166 (N_3166,N_2926,N_2824);
or U3167 (N_3167,N_2823,N_2866);
and U3168 (N_3168,N_2874,N_2945);
or U3169 (N_3169,N_2815,N_2974);
or U3170 (N_3170,N_2822,N_2921);
xor U3171 (N_3171,N_2801,N_2899);
xnor U3172 (N_3172,N_2979,N_2902);
or U3173 (N_3173,N_2918,N_2810);
nor U3174 (N_3174,N_2869,N_2860);
or U3175 (N_3175,N_2909,N_2902);
xor U3176 (N_3176,N_2850,N_2937);
nand U3177 (N_3177,N_2847,N_2915);
nand U3178 (N_3178,N_2919,N_2836);
xnor U3179 (N_3179,N_2986,N_2820);
or U3180 (N_3180,N_2823,N_2909);
nand U3181 (N_3181,N_2905,N_2920);
and U3182 (N_3182,N_2965,N_2860);
xor U3183 (N_3183,N_2913,N_2936);
or U3184 (N_3184,N_2802,N_2956);
nor U3185 (N_3185,N_2914,N_2835);
or U3186 (N_3186,N_2882,N_2863);
or U3187 (N_3187,N_2954,N_2809);
xnor U3188 (N_3188,N_2928,N_2891);
xor U3189 (N_3189,N_2818,N_2998);
nand U3190 (N_3190,N_2808,N_2935);
xnor U3191 (N_3191,N_2802,N_2815);
xnor U3192 (N_3192,N_2990,N_2816);
and U3193 (N_3193,N_2839,N_2824);
or U3194 (N_3194,N_2930,N_2921);
or U3195 (N_3195,N_2898,N_2813);
nand U3196 (N_3196,N_2953,N_2872);
nand U3197 (N_3197,N_2958,N_2858);
nand U3198 (N_3198,N_2879,N_2902);
nor U3199 (N_3199,N_2934,N_2888);
nor U3200 (N_3200,N_3092,N_3007);
and U3201 (N_3201,N_3169,N_3000);
nor U3202 (N_3202,N_3143,N_3184);
xnor U3203 (N_3203,N_3193,N_3032);
or U3204 (N_3204,N_3062,N_3128);
or U3205 (N_3205,N_3106,N_3014);
and U3206 (N_3206,N_3085,N_3010);
or U3207 (N_3207,N_3081,N_3049);
xnor U3208 (N_3208,N_3102,N_3185);
or U3209 (N_3209,N_3186,N_3166);
nor U3210 (N_3210,N_3120,N_3150);
xor U3211 (N_3211,N_3151,N_3059);
or U3212 (N_3212,N_3117,N_3051);
xnor U3213 (N_3213,N_3132,N_3015);
nand U3214 (N_3214,N_3152,N_3172);
xor U3215 (N_3215,N_3027,N_3159);
and U3216 (N_3216,N_3191,N_3023);
nor U3217 (N_3217,N_3138,N_3013);
or U3218 (N_3218,N_3095,N_3149);
nor U3219 (N_3219,N_3100,N_3107);
xor U3220 (N_3220,N_3019,N_3034);
or U3221 (N_3221,N_3194,N_3112);
nor U3222 (N_3222,N_3134,N_3114);
and U3223 (N_3223,N_3137,N_3155);
nor U3224 (N_3224,N_3153,N_3125);
nor U3225 (N_3225,N_3060,N_3198);
nand U3226 (N_3226,N_3174,N_3113);
nor U3227 (N_3227,N_3181,N_3175);
nand U3228 (N_3228,N_3161,N_3024);
or U3229 (N_3229,N_3101,N_3182);
nand U3230 (N_3230,N_3074,N_3111);
nand U3231 (N_3231,N_3176,N_3131);
nand U3232 (N_3232,N_3030,N_3040);
nor U3233 (N_3233,N_3088,N_3077);
nor U3234 (N_3234,N_3164,N_3020);
or U3235 (N_3235,N_3009,N_3171);
nor U3236 (N_3236,N_3043,N_3170);
and U3237 (N_3237,N_3055,N_3006);
nor U3238 (N_3238,N_3173,N_3070);
and U3239 (N_3239,N_3105,N_3156);
and U3240 (N_3240,N_3039,N_3099);
and U3241 (N_3241,N_3069,N_3177);
and U3242 (N_3242,N_3179,N_3018);
xnor U3243 (N_3243,N_3035,N_3192);
nor U3244 (N_3244,N_3118,N_3086);
and U3245 (N_3245,N_3075,N_3076);
and U3246 (N_3246,N_3124,N_3168);
nor U3247 (N_3247,N_3056,N_3011);
xnor U3248 (N_3248,N_3083,N_3057);
and U3249 (N_3249,N_3073,N_3180);
nor U3250 (N_3250,N_3109,N_3133);
xnor U3251 (N_3251,N_3022,N_3157);
and U3252 (N_3252,N_3135,N_3044);
and U3253 (N_3253,N_3001,N_3126);
xnor U3254 (N_3254,N_3154,N_3045);
xor U3255 (N_3255,N_3091,N_3071);
and U3256 (N_3256,N_3190,N_3163);
xnor U3257 (N_3257,N_3122,N_3119);
and U3258 (N_3258,N_3089,N_3005);
and U3259 (N_3259,N_3054,N_3072);
nor U3260 (N_3260,N_3063,N_3110);
nand U3261 (N_3261,N_3065,N_3090);
nand U3262 (N_3262,N_3196,N_3042);
and U3263 (N_3263,N_3187,N_3053);
and U3264 (N_3264,N_3038,N_3004);
xor U3265 (N_3265,N_3158,N_3199);
nor U3266 (N_3266,N_3094,N_3016);
nand U3267 (N_3267,N_3178,N_3046);
and U3268 (N_3268,N_3021,N_3141);
or U3269 (N_3269,N_3130,N_3129);
and U3270 (N_3270,N_3116,N_3050);
or U3271 (N_3271,N_3115,N_3183);
nor U3272 (N_3272,N_3189,N_3123);
nor U3273 (N_3273,N_3025,N_3033);
and U3274 (N_3274,N_3002,N_3061);
xor U3275 (N_3275,N_3028,N_3140);
nand U3276 (N_3276,N_3003,N_3145);
and U3277 (N_3277,N_3047,N_3064);
xor U3278 (N_3278,N_3026,N_3012);
and U3279 (N_3279,N_3037,N_3160);
nand U3280 (N_3280,N_3029,N_3148);
nor U3281 (N_3281,N_3127,N_3144);
nor U3282 (N_3282,N_3188,N_3136);
nand U3283 (N_3283,N_3121,N_3066);
nand U3284 (N_3284,N_3078,N_3080);
nand U3285 (N_3285,N_3052,N_3104);
or U3286 (N_3286,N_3036,N_3097);
nand U3287 (N_3287,N_3167,N_3048);
and U3288 (N_3288,N_3147,N_3195);
or U3289 (N_3289,N_3096,N_3103);
xnor U3290 (N_3290,N_3084,N_3058);
nor U3291 (N_3291,N_3068,N_3142);
or U3292 (N_3292,N_3197,N_3008);
nand U3293 (N_3293,N_3139,N_3087);
and U3294 (N_3294,N_3146,N_3067);
and U3295 (N_3295,N_3162,N_3165);
and U3296 (N_3296,N_3017,N_3093);
and U3297 (N_3297,N_3079,N_3031);
xor U3298 (N_3298,N_3082,N_3108);
nor U3299 (N_3299,N_3041,N_3098);
nor U3300 (N_3300,N_3058,N_3185);
nor U3301 (N_3301,N_3099,N_3068);
nand U3302 (N_3302,N_3146,N_3071);
nor U3303 (N_3303,N_3092,N_3116);
and U3304 (N_3304,N_3098,N_3138);
xnor U3305 (N_3305,N_3058,N_3178);
nor U3306 (N_3306,N_3034,N_3147);
xnor U3307 (N_3307,N_3081,N_3091);
xnor U3308 (N_3308,N_3068,N_3131);
nand U3309 (N_3309,N_3185,N_3155);
or U3310 (N_3310,N_3151,N_3067);
xor U3311 (N_3311,N_3025,N_3179);
nor U3312 (N_3312,N_3159,N_3047);
nand U3313 (N_3313,N_3196,N_3028);
and U3314 (N_3314,N_3123,N_3182);
nand U3315 (N_3315,N_3015,N_3139);
nor U3316 (N_3316,N_3083,N_3151);
and U3317 (N_3317,N_3055,N_3082);
and U3318 (N_3318,N_3187,N_3004);
nand U3319 (N_3319,N_3172,N_3038);
or U3320 (N_3320,N_3149,N_3132);
or U3321 (N_3321,N_3184,N_3125);
and U3322 (N_3322,N_3180,N_3096);
nor U3323 (N_3323,N_3013,N_3079);
nand U3324 (N_3324,N_3028,N_3004);
and U3325 (N_3325,N_3106,N_3187);
or U3326 (N_3326,N_3073,N_3048);
xnor U3327 (N_3327,N_3065,N_3017);
and U3328 (N_3328,N_3114,N_3128);
nand U3329 (N_3329,N_3022,N_3152);
or U3330 (N_3330,N_3099,N_3058);
or U3331 (N_3331,N_3118,N_3073);
and U3332 (N_3332,N_3137,N_3039);
xor U3333 (N_3333,N_3169,N_3186);
nand U3334 (N_3334,N_3064,N_3105);
and U3335 (N_3335,N_3118,N_3185);
and U3336 (N_3336,N_3186,N_3151);
nor U3337 (N_3337,N_3081,N_3125);
nor U3338 (N_3338,N_3132,N_3014);
nor U3339 (N_3339,N_3183,N_3137);
or U3340 (N_3340,N_3088,N_3178);
xnor U3341 (N_3341,N_3005,N_3029);
or U3342 (N_3342,N_3158,N_3178);
and U3343 (N_3343,N_3142,N_3169);
xor U3344 (N_3344,N_3199,N_3129);
nor U3345 (N_3345,N_3180,N_3145);
nand U3346 (N_3346,N_3149,N_3191);
nor U3347 (N_3347,N_3167,N_3033);
xor U3348 (N_3348,N_3150,N_3001);
xnor U3349 (N_3349,N_3062,N_3018);
xor U3350 (N_3350,N_3043,N_3030);
nor U3351 (N_3351,N_3071,N_3136);
or U3352 (N_3352,N_3040,N_3087);
and U3353 (N_3353,N_3191,N_3013);
nor U3354 (N_3354,N_3175,N_3126);
or U3355 (N_3355,N_3093,N_3123);
and U3356 (N_3356,N_3127,N_3086);
nand U3357 (N_3357,N_3040,N_3061);
nor U3358 (N_3358,N_3139,N_3080);
and U3359 (N_3359,N_3021,N_3039);
and U3360 (N_3360,N_3177,N_3195);
xor U3361 (N_3361,N_3159,N_3034);
nand U3362 (N_3362,N_3104,N_3164);
nor U3363 (N_3363,N_3061,N_3153);
nand U3364 (N_3364,N_3095,N_3185);
nor U3365 (N_3365,N_3169,N_3097);
nor U3366 (N_3366,N_3194,N_3050);
xor U3367 (N_3367,N_3089,N_3122);
or U3368 (N_3368,N_3101,N_3113);
nor U3369 (N_3369,N_3047,N_3158);
and U3370 (N_3370,N_3189,N_3064);
nand U3371 (N_3371,N_3167,N_3008);
nor U3372 (N_3372,N_3173,N_3044);
or U3373 (N_3373,N_3129,N_3017);
xnor U3374 (N_3374,N_3164,N_3024);
nand U3375 (N_3375,N_3127,N_3184);
xor U3376 (N_3376,N_3197,N_3154);
and U3377 (N_3377,N_3029,N_3156);
or U3378 (N_3378,N_3093,N_3108);
or U3379 (N_3379,N_3089,N_3150);
xor U3380 (N_3380,N_3029,N_3119);
or U3381 (N_3381,N_3138,N_3088);
or U3382 (N_3382,N_3085,N_3060);
or U3383 (N_3383,N_3174,N_3146);
or U3384 (N_3384,N_3064,N_3081);
and U3385 (N_3385,N_3165,N_3013);
nand U3386 (N_3386,N_3198,N_3050);
and U3387 (N_3387,N_3100,N_3175);
nor U3388 (N_3388,N_3067,N_3186);
xnor U3389 (N_3389,N_3033,N_3173);
nand U3390 (N_3390,N_3137,N_3170);
xor U3391 (N_3391,N_3075,N_3095);
nand U3392 (N_3392,N_3181,N_3105);
and U3393 (N_3393,N_3023,N_3010);
nor U3394 (N_3394,N_3068,N_3020);
and U3395 (N_3395,N_3008,N_3021);
nand U3396 (N_3396,N_3145,N_3067);
and U3397 (N_3397,N_3192,N_3149);
and U3398 (N_3398,N_3058,N_3172);
or U3399 (N_3399,N_3070,N_3169);
and U3400 (N_3400,N_3324,N_3383);
or U3401 (N_3401,N_3313,N_3237);
nand U3402 (N_3402,N_3365,N_3216);
or U3403 (N_3403,N_3243,N_3359);
xor U3404 (N_3404,N_3375,N_3258);
nor U3405 (N_3405,N_3239,N_3298);
and U3406 (N_3406,N_3323,N_3384);
nand U3407 (N_3407,N_3262,N_3335);
nor U3408 (N_3408,N_3315,N_3208);
nor U3409 (N_3409,N_3334,N_3302);
or U3410 (N_3410,N_3235,N_3223);
xor U3411 (N_3411,N_3364,N_3367);
and U3412 (N_3412,N_3245,N_3215);
nand U3413 (N_3413,N_3331,N_3273);
and U3414 (N_3414,N_3321,N_3277);
nand U3415 (N_3415,N_3372,N_3203);
and U3416 (N_3416,N_3358,N_3309);
nor U3417 (N_3417,N_3211,N_3362);
and U3418 (N_3418,N_3387,N_3288);
nand U3419 (N_3419,N_3269,N_3221);
nand U3420 (N_3420,N_3395,N_3389);
and U3421 (N_3421,N_3308,N_3327);
and U3422 (N_3422,N_3396,N_3342);
and U3423 (N_3423,N_3380,N_3294);
nor U3424 (N_3424,N_3338,N_3339);
and U3425 (N_3425,N_3311,N_3265);
or U3426 (N_3426,N_3207,N_3213);
nand U3427 (N_3427,N_3398,N_3297);
and U3428 (N_3428,N_3206,N_3247);
or U3429 (N_3429,N_3290,N_3240);
xnor U3430 (N_3430,N_3345,N_3353);
or U3431 (N_3431,N_3317,N_3241);
or U3432 (N_3432,N_3248,N_3319);
or U3433 (N_3433,N_3219,N_3373);
xor U3434 (N_3434,N_3363,N_3326);
xnor U3435 (N_3435,N_3307,N_3312);
and U3436 (N_3436,N_3379,N_3322);
and U3437 (N_3437,N_3236,N_3299);
xnor U3438 (N_3438,N_3357,N_3356);
xor U3439 (N_3439,N_3336,N_3220);
or U3440 (N_3440,N_3200,N_3397);
xnor U3441 (N_3441,N_3230,N_3279);
nand U3442 (N_3442,N_3204,N_3244);
xor U3443 (N_3443,N_3314,N_3232);
nor U3444 (N_3444,N_3226,N_3305);
nand U3445 (N_3445,N_3284,N_3252);
and U3446 (N_3446,N_3275,N_3371);
nor U3447 (N_3447,N_3276,N_3257);
nor U3448 (N_3448,N_3361,N_3378);
xor U3449 (N_3449,N_3253,N_3306);
nand U3450 (N_3450,N_3388,N_3394);
nand U3451 (N_3451,N_3328,N_3251);
xor U3452 (N_3452,N_3280,N_3348);
nor U3453 (N_3453,N_3381,N_3391);
nand U3454 (N_3454,N_3346,N_3254);
xnor U3455 (N_3455,N_3201,N_3296);
or U3456 (N_3456,N_3289,N_3271);
nor U3457 (N_3457,N_3354,N_3374);
and U3458 (N_3458,N_3242,N_3368);
nand U3459 (N_3459,N_3218,N_3376);
nor U3460 (N_3460,N_3347,N_3349);
nand U3461 (N_3461,N_3343,N_3337);
xnor U3462 (N_3462,N_3225,N_3390);
xnor U3463 (N_3463,N_3274,N_3222);
nor U3464 (N_3464,N_3366,N_3259);
nor U3465 (N_3465,N_3256,N_3227);
or U3466 (N_3466,N_3217,N_3350);
and U3467 (N_3467,N_3304,N_3234);
nor U3468 (N_3468,N_3270,N_3263);
nor U3469 (N_3469,N_3281,N_3250);
and U3470 (N_3470,N_3231,N_3255);
nand U3471 (N_3471,N_3344,N_3249);
and U3472 (N_3472,N_3205,N_3295);
or U3473 (N_3473,N_3310,N_3260);
and U3474 (N_3474,N_3325,N_3210);
nand U3475 (N_3475,N_3369,N_3341);
nor U3476 (N_3476,N_3214,N_3209);
or U3477 (N_3477,N_3266,N_3340);
nand U3478 (N_3478,N_3330,N_3268);
and U3479 (N_3479,N_3351,N_3224);
xnor U3480 (N_3480,N_3292,N_3246);
nor U3481 (N_3481,N_3393,N_3386);
nor U3482 (N_3482,N_3360,N_3392);
or U3483 (N_3483,N_3332,N_3300);
or U3484 (N_3484,N_3282,N_3283);
or U3485 (N_3485,N_3287,N_3293);
nor U3486 (N_3486,N_3212,N_3318);
and U3487 (N_3487,N_3303,N_3285);
xor U3488 (N_3488,N_3228,N_3301);
and U3489 (N_3489,N_3238,N_3370);
nand U3490 (N_3490,N_3233,N_3355);
nor U3491 (N_3491,N_3377,N_3382);
nor U3492 (N_3492,N_3352,N_3399);
and U3493 (N_3493,N_3329,N_3316);
nand U3494 (N_3494,N_3278,N_3272);
nand U3495 (N_3495,N_3267,N_3286);
nor U3496 (N_3496,N_3261,N_3333);
or U3497 (N_3497,N_3229,N_3264);
or U3498 (N_3498,N_3202,N_3291);
xor U3499 (N_3499,N_3320,N_3385);
nor U3500 (N_3500,N_3240,N_3372);
or U3501 (N_3501,N_3238,N_3242);
xor U3502 (N_3502,N_3202,N_3284);
or U3503 (N_3503,N_3270,N_3348);
xnor U3504 (N_3504,N_3256,N_3339);
and U3505 (N_3505,N_3355,N_3397);
and U3506 (N_3506,N_3211,N_3229);
or U3507 (N_3507,N_3262,N_3395);
nor U3508 (N_3508,N_3231,N_3371);
and U3509 (N_3509,N_3311,N_3261);
nor U3510 (N_3510,N_3369,N_3348);
nor U3511 (N_3511,N_3361,N_3259);
nor U3512 (N_3512,N_3216,N_3302);
nand U3513 (N_3513,N_3265,N_3326);
xnor U3514 (N_3514,N_3348,N_3274);
or U3515 (N_3515,N_3310,N_3290);
nor U3516 (N_3516,N_3276,N_3208);
and U3517 (N_3517,N_3246,N_3211);
and U3518 (N_3518,N_3272,N_3352);
and U3519 (N_3519,N_3226,N_3392);
or U3520 (N_3520,N_3290,N_3348);
nand U3521 (N_3521,N_3366,N_3355);
nand U3522 (N_3522,N_3238,N_3223);
nor U3523 (N_3523,N_3229,N_3365);
xor U3524 (N_3524,N_3328,N_3397);
xnor U3525 (N_3525,N_3231,N_3399);
xnor U3526 (N_3526,N_3206,N_3382);
and U3527 (N_3527,N_3354,N_3241);
nand U3528 (N_3528,N_3315,N_3385);
or U3529 (N_3529,N_3346,N_3266);
nor U3530 (N_3530,N_3227,N_3281);
nor U3531 (N_3531,N_3220,N_3379);
or U3532 (N_3532,N_3233,N_3325);
and U3533 (N_3533,N_3290,N_3380);
xnor U3534 (N_3534,N_3358,N_3357);
nor U3535 (N_3535,N_3322,N_3350);
xor U3536 (N_3536,N_3333,N_3230);
nor U3537 (N_3537,N_3202,N_3330);
nor U3538 (N_3538,N_3336,N_3215);
nand U3539 (N_3539,N_3397,N_3250);
and U3540 (N_3540,N_3247,N_3305);
or U3541 (N_3541,N_3398,N_3224);
nor U3542 (N_3542,N_3211,N_3290);
or U3543 (N_3543,N_3345,N_3310);
and U3544 (N_3544,N_3329,N_3282);
xnor U3545 (N_3545,N_3340,N_3299);
xnor U3546 (N_3546,N_3367,N_3384);
xor U3547 (N_3547,N_3235,N_3312);
or U3548 (N_3548,N_3387,N_3211);
or U3549 (N_3549,N_3200,N_3215);
and U3550 (N_3550,N_3330,N_3266);
nor U3551 (N_3551,N_3310,N_3293);
nand U3552 (N_3552,N_3206,N_3361);
nor U3553 (N_3553,N_3240,N_3222);
or U3554 (N_3554,N_3310,N_3327);
nand U3555 (N_3555,N_3217,N_3356);
or U3556 (N_3556,N_3326,N_3250);
and U3557 (N_3557,N_3361,N_3258);
nand U3558 (N_3558,N_3304,N_3291);
nand U3559 (N_3559,N_3265,N_3284);
nor U3560 (N_3560,N_3226,N_3260);
xnor U3561 (N_3561,N_3325,N_3299);
xor U3562 (N_3562,N_3281,N_3206);
or U3563 (N_3563,N_3292,N_3307);
xnor U3564 (N_3564,N_3254,N_3376);
nand U3565 (N_3565,N_3299,N_3350);
nand U3566 (N_3566,N_3339,N_3266);
or U3567 (N_3567,N_3262,N_3344);
or U3568 (N_3568,N_3356,N_3243);
xor U3569 (N_3569,N_3365,N_3239);
or U3570 (N_3570,N_3276,N_3256);
and U3571 (N_3571,N_3213,N_3264);
and U3572 (N_3572,N_3300,N_3226);
nor U3573 (N_3573,N_3300,N_3287);
nor U3574 (N_3574,N_3352,N_3252);
nand U3575 (N_3575,N_3337,N_3210);
nor U3576 (N_3576,N_3258,N_3389);
or U3577 (N_3577,N_3274,N_3354);
nor U3578 (N_3578,N_3264,N_3381);
and U3579 (N_3579,N_3341,N_3367);
or U3580 (N_3580,N_3355,N_3375);
and U3581 (N_3581,N_3223,N_3299);
xnor U3582 (N_3582,N_3211,N_3210);
nor U3583 (N_3583,N_3325,N_3313);
nand U3584 (N_3584,N_3357,N_3373);
nand U3585 (N_3585,N_3309,N_3241);
nor U3586 (N_3586,N_3324,N_3254);
xor U3587 (N_3587,N_3314,N_3252);
or U3588 (N_3588,N_3313,N_3242);
nand U3589 (N_3589,N_3215,N_3251);
nor U3590 (N_3590,N_3267,N_3360);
nand U3591 (N_3591,N_3229,N_3353);
xor U3592 (N_3592,N_3322,N_3386);
xor U3593 (N_3593,N_3268,N_3396);
or U3594 (N_3594,N_3351,N_3388);
and U3595 (N_3595,N_3316,N_3229);
nor U3596 (N_3596,N_3257,N_3278);
xnor U3597 (N_3597,N_3396,N_3264);
nor U3598 (N_3598,N_3233,N_3240);
or U3599 (N_3599,N_3315,N_3218);
and U3600 (N_3600,N_3445,N_3558);
and U3601 (N_3601,N_3428,N_3535);
nand U3602 (N_3602,N_3473,N_3413);
or U3603 (N_3603,N_3463,N_3544);
nand U3604 (N_3604,N_3451,N_3454);
nor U3605 (N_3605,N_3580,N_3582);
xor U3606 (N_3606,N_3455,N_3512);
or U3607 (N_3607,N_3472,N_3407);
nand U3608 (N_3608,N_3575,N_3448);
or U3609 (N_3609,N_3539,N_3481);
or U3610 (N_3610,N_3443,N_3442);
nor U3611 (N_3611,N_3515,N_3487);
and U3612 (N_3612,N_3453,N_3457);
xor U3613 (N_3613,N_3595,N_3470);
nor U3614 (N_3614,N_3497,N_3495);
nor U3615 (N_3615,N_3412,N_3509);
nor U3616 (N_3616,N_3585,N_3446);
or U3617 (N_3617,N_3565,N_3519);
nor U3618 (N_3618,N_3459,N_3427);
and U3619 (N_3619,N_3500,N_3444);
or U3620 (N_3620,N_3400,N_3420);
xnor U3621 (N_3621,N_3489,N_3566);
nand U3622 (N_3622,N_3542,N_3559);
nand U3623 (N_3623,N_3402,N_3464);
and U3624 (N_3624,N_3468,N_3494);
or U3625 (N_3625,N_3404,N_3525);
nor U3626 (N_3626,N_3591,N_3552);
nor U3627 (N_3627,N_3488,N_3432);
xor U3628 (N_3628,N_3594,N_3460);
nand U3629 (N_3629,N_3556,N_3571);
or U3630 (N_3630,N_3521,N_3574);
nor U3631 (N_3631,N_3449,N_3549);
xnor U3632 (N_3632,N_3403,N_3490);
nor U3633 (N_3633,N_3541,N_3504);
and U3634 (N_3634,N_3540,N_3422);
or U3635 (N_3635,N_3408,N_3532);
nand U3636 (N_3636,N_3452,N_3456);
nand U3637 (N_3637,N_3598,N_3406);
nor U3638 (N_3638,N_3557,N_3416);
nand U3639 (N_3639,N_3531,N_3505);
nand U3640 (N_3640,N_3506,N_3530);
xnor U3641 (N_3641,N_3570,N_3496);
or U3642 (N_3642,N_3433,N_3499);
nand U3643 (N_3643,N_3415,N_3520);
nor U3644 (N_3644,N_3465,N_3438);
nor U3645 (N_3645,N_3480,N_3522);
or U3646 (N_3646,N_3462,N_3423);
nor U3647 (N_3647,N_3562,N_3476);
xor U3648 (N_3648,N_3529,N_3551);
or U3649 (N_3649,N_3498,N_3483);
nand U3650 (N_3650,N_3405,N_3418);
nand U3651 (N_3651,N_3550,N_3466);
nand U3652 (N_3652,N_3435,N_3471);
and U3653 (N_3653,N_3579,N_3461);
nand U3654 (N_3654,N_3482,N_3417);
and U3655 (N_3655,N_3501,N_3543);
xor U3656 (N_3656,N_3596,N_3584);
or U3657 (N_3657,N_3429,N_3436);
and U3658 (N_3658,N_3474,N_3564);
nor U3659 (N_3659,N_3511,N_3578);
and U3660 (N_3660,N_3524,N_3593);
nor U3661 (N_3661,N_3517,N_3587);
nand U3662 (N_3662,N_3586,N_3430);
xnor U3663 (N_3663,N_3437,N_3514);
xor U3664 (N_3664,N_3589,N_3560);
and U3665 (N_3665,N_3441,N_3507);
nand U3666 (N_3666,N_3590,N_3561);
nor U3667 (N_3667,N_3425,N_3410);
xor U3668 (N_3668,N_3475,N_3588);
xnor U3669 (N_3669,N_3518,N_3502);
or U3670 (N_3670,N_3583,N_3523);
or U3671 (N_3671,N_3548,N_3447);
nand U3672 (N_3672,N_3568,N_3577);
nor U3673 (N_3673,N_3478,N_3467);
or U3674 (N_3674,N_3411,N_3528);
nand U3675 (N_3675,N_3450,N_3414);
nand U3676 (N_3676,N_3426,N_3440);
or U3677 (N_3677,N_3439,N_3569);
or U3678 (N_3678,N_3592,N_3573);
nand U3679 (N_3679,N_3572,N_3485);
and U3680 (N_3680,N_3576,N_3563);
and U3681 (N_3681,N_3503,N_3484);
xor U3682 (N_3682,N_3508,N_3513);
nand U3683 (N_3683,N_3469,N_3545);
nor U3684 (N_3684,N_3527,N_3486);
and U3685 (N_3685,N_3538,N_3479);
xnor U3686 (N_3686,N_3493,N_3516);
xor U3687 (N_3687,N_3555,N_3421);
xnor U3688 (N_3688,N_3526,N_3510);
nand U3689 (N_3689,N_3401,N_3581);
nand U3690 (N_3690,N_3536,N_3477);
or U3691 (N_3691,N_3546,N_3424);
nor U3692 (N_3692,N_3458,N_3547);
nand U3693 (N_3693,N_3553,N_3599);
nand U3694 (N_3694,N_3491,N_3419);
xor U3695 (N_3695,N_3534,N_3554);
nand U3696 (N_3696,N_3409,N_3492);
nor U3697 (N_3697,N_3567,N_3434);
xnor U3698 (N_3698,N_3537,N_3431);
nor U3699 (N_3699,N_3533,N_3597);
or U3700 (N_3700,N_3572,N_3573);
or U3701 (N_3701,N_3527,N_3431);
xnor U3702 (N_3702,N_3420,N_3573);
nor U3703 (N_3703,N_3429,N_3572);
xor U3704 (N_3704,N_3497,N_3481);
nor U3705 (N_3705,N_3473,N_3583);
nand U3706 (N_3706,N_3404,N_3442);
or U3707 (N_3707,N_3523,N_3552);
nand U3708 (N_3708,N_3545,N_3567);
xor U3709 (N_3709,N_3534,N_3494);
or U3710 (N_3710,N_3424,N_3458);
nand U3711 (N_3711,N_3425,N_3511);
nor U3712 (N_3712,N_3518,N_3426);
or U3713 (N_3713,N_3507,N_3564);
xor U3714 (N_3714,N_3523,N_3500);
xnor U3715 (N_3715,N_3483,N_3407);
nor U3716 (N_3716,N_3503,N_3517);
or U3717 (N_3717,N_3412,N_3422);
or U3718 (N_3718,N_3488,N_3555);
nor U3719 (N_3719,N_3536,N_3552);
or U3720 (N_3720,N_3577,N_3456);
nand U3721 (N_3721,N_3581,N_3524);
and U3722 (N_3722,N_3535,N_3542);
or U3723 (N_3723,N_3503,N_3450);
nor U3724 (N_3724,N_3442,N_3590);
and U3725 (N_3725,N_3593,N_3586);
nand U3726 (N_3726,N_3473,N_3541);
nor U3727 (N_3727,N_3425,N_3547);
nand U3728 (N_3728,N_3585,N_3413);
xnor U3729 (N_3729,N_3570,N_3447);
xor U3730 (N_3730,N_3569,N_3510);
nor U3731 (N_3731,N_3400,N_3410);
nand U3732 (N_3732,N_3593,N_3599);
nand U3733 (N_3733,N_3420,N_3557);
nand U3734 (N_3734,N_3580,N_3418);
nor U3735 (N_3735,N_3420,N_3599);
nand U3736 (N_3736,N_3417,N_3401);
nor U3737 (N_3737,N_3534,N_3579);
and U3738 (N_3738,N_3475,N_3457);
or U3739 (N_3739,N_3497,N_3529);
xnor U3740 (N_3740,N_3480,N_3527);
nor U3741 (N_3741,N_3402,N_3478);
or U3742 (N_3742,N_3472,N_3591);
or U3743 (N_3743,N_3412,N_3591);
or U3744 (N_3744,N_3504,N_3571);
and U3745 (N_3745,N_3556,N_3500);
nor U3746 (N_3746,N_3404,N_3431);
and U3747 (N_3747,N_3427,N_3421);
nand U3748 (N_3748,N_3481,N_3507);
or U3749 (N_3749,N_3530,N_3509);
nor U3750 (N_3750,N_3429,N_3552);
nand U3751 (N_3751,N_3509,N_3514);
nor U3752 (N_3752,N_3578,N_3549);
or U3753 (N_3753,N_3477,N_3421);
nand U3754 (N_3754,N_3443,N_3516);
nand U3755 (N_3755,N_3558,N_3549);
nor U3756 (N_3756,N_3552,N_3497);
nand U3757 (N_3757,N_3470,N_3472);
xor U3758 (N_3758,N_3566,N_3508);
or U3759 (N_3759,N_3560,N_3583);
or U3760 (N_3760,N_3493,N_3501);
and U3761 (N_3761,N_3563,N_3559);
or U3762 (N_3762,N_3427,N_3483);
nand U3763 (N_3763,N_3595,N_3433);
xnor U3764 (N_3764,N_3499,N_3554);
nand U3765 (N_3765,N_3571,N_3489);
and U3766 (N_3766,N_3545,N_3563);
nand U3767 (N_3767,N_3477,N_3499);
xnor U3768 (N_3768,N_3593,N_3592);
nand U3769 (N_3769,N_3507,N_3416);
or U3770 (N_3770,N_3452,N_3560);
or U3771 (N_3771,N_3453,N_3545);
xnor U3772 (N_3772,N_3478,N_3525);
nor U3773 (N_3773,N_3554,N_3512);
nor U3774 (N_3774,N_3432,N_3479);
nor U3775 (N_3775,N_3544,N_3509);
nand U3776 (N_3776,N_3418,N_3522);
or U3777 (N_3777,N_3466,N_3442);
nand U3778 (N_3778,N_3405,N_3520);
or U3779 (N_3779,N_3491,N_3569);
and U3780 (N_3780,N_3567,N_3400);
and U3781 (N_3781,N_3501,N_3489);
or U3782 (N_3782,N_3571,N_3481);
nor U3783 (N_3783,N_3518,N_3415);
xnor U3784 (N_3784,N_3429,N_3594);
nand U3785 (N_3785,N_3556,N_3427);
xor U3786 (N_3786,N_3546,N_3554);
nor U3787 (N_3787,N_3459,N_3523);
nand U3788 (N_3788,N_3483,N_3491);
and U3789 (N_3789,N_3443,N_3490);
or U3790 (N_3790,N_3545,N_3566);
nand U3791 (N_3791,N_3554,N_3493);
and U3792 (N_3792,N_3426,N_3476);
or U3793 (N_3793,N_3480,N_3584);
nor U3794 (N_3794,N_3587,N_3541);
or U3795 (N_3795,N_3594,N_3595);
or U3796 (N_3796,N_3480,N_3503);
nor U3797 (N_3797,N_3596,N_3569);
or U3798 (N_3798,N_3589,N_3476);
nand U3799 (N_3799,N_3522,N_3443);
or U3800 (N_3800,N_3635,N_3787);
or U3801 (N_3801,N_3795,N_3649);
nand U3802 (N_3802,N_3713,N_3698);
or U3803 (N_3803,N_3615,N_3708);
or U3804 (N_3804,N_3656,N_3633);
nor U3805 (N_3805,N_3636,N_3648);
and U3806 (N_3806,N_3683,N_3764);
nand U3807 (N_3807,N_3645,N_3717);
and U3808 (N_3808,N_3791,N_3607);
and U3809 (N_3809,N_3673,N_3600);
nand U3810 (N_3810,N_3628,N_3680);
or U3811 (N_3811,N_3719,N_3729);
nand U3812 (N_3812,N_3634,N_3766);
nand U3813 (N_3813,N_3650,N_3785);
and U3814 (N_3814,N_3721,N_3726);
xor U3815 (N_3815,N_3614,N_3730);
and U3816 (N_3816,N_3706,N_3620);
or U3817 (N_3817,N_3627,N_3747);
or U3818 (N_3818,N_3704,N_3722);
and U3819 (N_3819,N_3754,N_3741);
and U3820 (N_3820,N_3731,N_3753);
or U3821 (N_3821,N_3782,N_3789);
xor U3822 (N_3822,N_3792,N_3779);
and U3823 (N_3823,N_3681,N_3701);
xor U3824 (N_3824,N_3765,N_3632);
nor U3825 (N_3825,N_3685,N_3646);
xor U3826 (N_3826,N_3703,N_3723);
xnor U3827 (N_3827,N_3748,N_3644);
xnor U3828 (N_3828,N_3696,N_3750);
xnor U3829 (N_3829,N_3734,N_3702);
and U3830 (N_3830,N_3638,N_3737);
xor U3831 (N_3831,N_3755,N_3629);
xnor U3832 (N_3832,N_3727,N_3712);
nor U3833 (N_3833,N_3616,N_3666);
or U3834 (N_3834,N_3661,N_3674);
nand U3835 (N_3835,N_3718,N_3767);
and U3836 (N_3836,N_3625,N_3602);
nand U3837 (N_3837,N_3679,N_3608);
and U3838 (N_3838,N_3793,N_3610);
or U3839 (N_3839,N_3763,N_3637);
xnor U3840 (N_3840,N_3746,N_3768);
nand U3841 (N_3841,N_3733,N_3735);
nand U3842 (N_3842,N_3690,N_3653);
or U3843 (N_3843,N_3740,N_3647);
nand U3844 (N_3844,N_3672,N_3669);
nand U3845 (N_3845,N_3752,N_3697);
nand U3846 (N_3846,N_3688,N_3682);
xnor U3847 (N_3847,N_3709,N_3714);
and U3848 (N_3848,N_3642,N_3770);
and U3849 (N_3849,N_3640,N_3694);
nor U3850 (N_3850,N_3799,N_3624);
nand U3851 (N_3851,N_3742,N_3758);
and U3852 (N_3852,N_3711,N_3715);
nand U3853 (N_3853,N_3759,N_3798);
or U3854 (N_3854,N_3777,N_3776);
nand U3855 (N_3855,N_3678,N_3728);
xnor U3856 (N_3856,N_3790,N_3736);
and U3857 (N_3857,N_3670,N_3738);
nand U3858 (N_3858,N_3655,N_3603);
xor U3859 (N_3859,N_3797,N_3716);
or U3860 (N_3860,N_3643,N_3664);
or U3861 (N_3861,N_3623,N_3732);
and U3862 (N_3862,N_3676,N_3760);
and U3863 (N_3863,N_3772,N_3699);
nor U3864 (N_3864,N_3675,N_3687);
and U3865 (N_3865,N_3775,N_3606);
nand U3866 (N_3866,N_3665,N_3684);
nand U3867 (N_3867,N_3619,N_3622);
nand U3868 (N_3868,N_3662,N_3778);
xnor U3869 (N_3869,N_3660,N_3631);
nand U3870 (N_3870,N_3700,N_3626);
nand U3871 (N_3871,N_3609,N_3693);
and U3872 (N_3872,N_3658,N_3668);
nor U3873 (N_3873,N_3686,N_3618);
nand U3874 (N_3874,N_3705,N_3677);
xnor U3875 (N_3875,N_3657,N_3761);
or U3876 (N_3876,N_3710,N_3651);
xor U3877 (N_3877,N_3663,N_3771);
nand U3878 (N_3878,N_3762,N_3691);
nand U3879 (N_3879,N_3654,N_3692);
xor U3880 (N_3880,N_3743,N_3601);
nor U3881 (N_3881,N_3613,N_3641);
nand U3882 (N_3882,N_3796,N_3786);
or U3883 (N_3883,N_3781,N_3749);
nand U3884 (N_3884,N_3780,N_3756);
nand U3885 (N_3885,N_3745,N_3788);
and U3886 (N_3886,N_3739,N_3774);
nor U3887 (N_3887,N_3671,N_3751);
xnor U3888 (N_3888,N_3744,N_3689);
and U3889 (N_3889,N_3794,N_3773);
xor U3890 (N_3890,N_3652,N_3757);
nor U3891 (N_3891,N_3769,N_3725);
and U3892 (N_3892,N_3621,N_3784);
and U3893 (N_3893,N_3659,N_3617);
or U3894 (N_3894,N_3720,N_3667);
nand U3895 (N_3895,N_3605,N_3612);
or U3896 (N_3896,N_3611,N_3724);
nor U3897 (N_3897,N_3783,N_3695);
nor U3898 (N_3898,N_3639,N_3707);
and U3899 (N_3899,N_3604,N_3630);
and U3900 (N_3900,N_3785,N_3687);
nor U3901 (N_3901,N_3661,N_3691);
nand U3902 (N_3902,N_3798,N_3691);
nor U3903 (N_3903,N_3787,N_3705);
xnor U3904 (N_3904,N_3628,N_3785);
or U3905 (N_3905,N_3604,N_3795);
nand U3906 (N_3906,N_3612,N_3720);
or U3907 (N_3907,N_3672,N_3635);
and U3908 (N_3908,N_3600,N_3714);
nand U3909 (N_3909,N_3748,N_3635);
xor U3910 (N_3910,N_3705,N_3755);
or U3911 (N_3911,N_3749,N_3740);
xnor U3912 (N_3912,N_3702,N_3710);
xnor U3913 (N_3913,N_3796,N_3709);
nand U3914 (N_3914,N_3736,N_3618);
nor U3915 (N_3915,N_3650,N_3699);
nor U3916 (N_3916,N_3659,N_3742);
nand U3917 (N_3917,N_3617,N_3767);
nand U3918 (N_3918,N_3775,N_3636);
nor U3919 (N_3919,N_3691,N_3718);
or U3920 (N_3920,N_3628,N_3748);
and U3921 (N_3921,N_3681,N_3732);
nor U3922 (N_3922,N_3718,N_3643);
and U3923 (N_3923,N_3724,N_3722);
and U3924 (N_3924,N_3672,N_3747);
and U3925 (N_3925,N_3706,N_3751);
and U3926 (N_3926,N_3646,N_3620);
and U3927 (N_3927,N_3627,N_3676);
nor U3928 (N_3928,N_3642,N_3613);
nand U3929 (N_3929,N_3707,N_3738);
nand U3930 (N_3930,N_3765,N_3741);
xor U3931 (N_3931,N_3735,N_3635);
or U3932 (N_3932,N_3601,N_3794);
nor U3933 (N_3933,N_3732,N_3790);
or U3934 (N_3934,N_3683,N_3775);
nand U3935 (N_3935,N_3620,N_3643);
nor U3936 (N_3936,N_3664,N_3739);
and U3937 (N_3937,N_3783,N_3769);
xor U3938 (N_3938,N_3745,N_3791);
nand U3939 (N_3939,N_3724,N_3677);
and U3940 (N_3940,N_3651,N_3737);
nand U3941 (N_3941,N_3695,N_3767);
nand U3942 (N_3942,N_3739,N_3648);
nor U3943 (N_3943,N_3760,N_3628);
or U3944 (N_3944,N_3727,N_3651);
and U3945 (N_3945,N_3604,N_3660);
or U3946 (N_3946,N_3734,N_3630);
or U3947 (N_3947,N_3791,N_3729);
nor U3948 (N_3948,N_3752,N_3757);
and U3949 (N_3949,N_3648,N_3743);
and U3950 (N_3950,N_3666,N_3641);
or U3951 (N_3951,N_3656,N_3744);
xor U3952 (N_3952,N_3602,N_3608);
or U3953 (N_3953,N_3698,N_3623);
and U3954 (N_3954,N_3607,N_3792);
nand U3955 (N_3955,N_3626,N_3676);
nor U3956 (N_3956,N_3624,N_3680);
nor U3957 (N_3957,N_3697,N_3773);
or U3958 (N_3958,N_3665,N_3696);
and U3959 (N_3959,N_3603,N_3721);
xnor U3960 (N_3960,N_3622,N_3605);
xnor U3961 (N_3961,N_3602,N_3794);
nand U3962 (N_3962,N_3739,N_3745);
or U3963 (N_3963,N_3637,N_3735);
nor U3964 (N_3964,N_3695,N_3724);
or U3965 (N_3965,N_3644,N_3641);
and U3966 (N_3966,N_3798,N_3728);
xor U3967 (N_3967,N_3606,N_3608);
nand U3968 (N_3968,N_3726,N_3641);
nand U3969 (N_3969,N_3739,N_3691);
nand U3970 (N_3970,N_3717,N_3718);
and U3971 (N_3971,N_3618,N_3630);
and U3972 (N_3972,N_3675,N_3692);
nand U3973 (N_3973,N_3754,N_3722);
xnor U3974 (N_3974,N_3750,N_3778);
nor U3975 (N_3975,N_3627,N_3713);
or U3976 (N_3976,N_3697,N_3651);
nor U3977 (N_3977,N_3646,N_3746);
nor U3978 (N_3978,N_3767,N_3779);
or U3979 (N_3979,N_3642,N_3732);
nor U3980 (N_3980,N_3600,N_3780);
and U3981 (N_3981,N_3656,N_3754);
nand U3982 (N_3982,N_3698,N_3742);
nor U3983 (N_3983,N_3779,N_3735);
nor U3984 (N_3984,N_3624,N_3750);
xor U3985 (N_3985,N_3750,N_3701);
xnor U3986 (N_3986,N_3643,N_3674);
xnor U3987 (N_3987,N_3706,N_3786);
and U3988 (N_3988,N_3656,N_3630);
or U3989 (N_3989,N_3737,N_3633);
and U3990 (N_3990,N_3737,N_3613);
xor U3991 (N_3991,N_3762,N_3779);
and U3992 (N_3992,N_3682,N_3750);
nor U3993 (N_3993,N_3779,N_3785);
and U3994 (N_3994,N_3775,N_3637);
nand U3995 (N_3995,N_3668,N_3652);
xor U3996 (N_3996,N_3675,N_3643);
or U3997 (N_3997,N_3731,N_3659);
nand U3998 (N_3998,N_3654,N_3703);
nand U3999 (N_3999,N_3785,N_3716);
and U4000 (N_4000,N_3982,N_3813);
nand U4001 (N_4001,N_3947,N_3826);
nand U4002 (N_4002,N_3925,N_3970);
and U4003 (N_4003,N_3894,N_3991);
nand U4004 (N_4004,N_3931,N_3888);
xnor U4005 (N_4005,N_3962,N_3956);
nand U4006 (N_4006,N_3915,N_3800);
and U4007 (N_4007,N_3876,N_3940);
nand U4008 (N_4008,N_3987,N_3859);
or U4009 (N_4009,N_3874,N_3938);
nand U4010 (N_4010,N_3990,N_3933);
or U4011 (N_4011,N_3966,N_3881);
nand U4012 (N_4012,N_3955,N_3952);
and U4013 (N_4013,N_3858,N_3946);
or U4014 (N_4014,N_3854,N_3944);
nand U4015 (N_4015,N_3864,N_3812);
xnor U4016 (N_4016,N_3939,N_3927);
nand U4017 (N_4017,N_3852,N_3849);
nand U4018 (N_4018,N_3880,N_3839);
and U4019 (N_4019,N_3937,N_3953);
nor U4020 (N_4020,N_3905,N_3995);
xor U4021 (N_4021,N_3992,N_3842);
nor U4022 (N_4022,N_3808,N_3890);
and U4023 (N_4023,N_3868,N_3855);
xnor U4024 (N_4024,N_3968,N_3950);
and U4025 (N_4025,N_3886,N_3814);
xnor U4026 (N_4026,N_3835,N_3872);
nand U4027 (N_4027,N_3932,N_3945);
nand U4028 (N_4028,N_3806,N_3900);
nor U4029 (N_4029,N_3830,N_3951);
and U4030 (N_4030,N_3924,N_3893);
and U4031 (N_4031,N_3973,N_3928);
xor U4032 (N_4032,N_3870,N_3838);
nor U4033 (N_4033,N_3909,N_3910);
xnor U4034 (N_4034,N_3977,N_3861);
nor U4035 (N_4035,N_3980,N_3862);
or U4036 (N_4036,N_3983,N_3804);
nand U4037 (N_4037,N_3887,N_3899);
nor U4038 (N_4038,N_3896,N_3914);
nor U4039 (N_4039,N_3892,N_3967);
and U4040 (N_4040,N_3949,N_3829);
nand U4041 (N_4041,N_3837,N_3803);
nand U4042 (N_4042,N_3822,N_3875);
xnor U4043 (N_4043,N_3972,N_3930);
nand U4044 (N_4044,N_3964,N_3817);
nor U4045 (N_4045,N_3853,N_3903);
xor U4046 (N_4046,N_3959,N_3845);
xor U4047 (N_4047,N_3936,N_3877);
or U4048 (N_4048,N_3878,N_3979);
xor U4049 (N_4049,N_3891,N_3923);
xor U4050 (N_4050,N_3828,N_3846);
xnor U4051 (N_4051,N_3848,N_3921);
nor U4052 (N_4052,N_3882,N_3901);
xnor U4053 (N_4053,N_3897,N_3907);
and U4054 (N_4054,N_3863,N_3867);
nor U4055 (N_4055,N_3856,N_3818);
xnor U4056 (N_4056,N_3801,N_3851);
and U4057 (N_4057,N_3988,N_3919);
xor U4058 (N_4058,N_3831,N_3918);
and U4059 (N_4059,N_3957,N_3833);
nand U4060 (N_4060,N_3963,N_3843);
nor U4061 (N_4061,N_3997,N_3815);
and U4062 (N_4062,N_3948,N_3998);
nor U4063 (N_4063,N_3895,N_3810);
xor U4064 (N_4064,N_3984,N_3840);
nand U4065 (N_4065,N_3994,N_3985);
and U4066 (N_4066,N_3844,N_3805);
nor U4067 (N_4067,N_3941,N_3871);
nand U4068 (N_4068,N_3847,N_3920);
and U4069 (N_4069,N_3943,N_3879);
xor U4070 (N_4070,N_3954,N_3821);
xor U4071 (N_4071,N_3935,N_3841);
and U4072 (N_4072,N_3993,N_3926);
nand U4073 (N_4073,N_3974,N_3999);
xnor U4074 (N_4074,N_3866,N_3965);
nor U4075 (N_4075,N_3827,N_3986);
xnor U4076 (N_4076,N_3917,N_3975);
and U4077 (N_4077,N_3884,N_3873);
xnor U4078 (N_4078,N_3857,N_3913);
nor U4079 (N_4079,N_3883,N_3869);
xor U4080 (N_4080,N_3929,N_3996);
nor U4081 (N_4081,N_3885,N_3811);
or U4082 (N_4082,N_3978,N_3809);
xnor U4083 (N_4083,N_3971,N_3904);
xor U4084 (N_4084,N_3834,N_3960);
nor U4085 (N_4085,N_3981,N_3989);
or U4086 (N_4086,N_3916,N_3961);
nand U4087 (N_4087,N_3976,N_3836);
or U4088 (N_4088,N_3911,N_3912);
xor U4089 (N_4089,N_3969,N_3908);
and U4090 (N_4090,N_3902,N_3802);
nand U4091 (N_4091,N_3819,N_3824);
or U4092 (N_4092,N_3889,N_3906);
and U4093 (N_4093,N_3922,N_3934);
nand U4094 (N_4094,N_3820,N_3865);
nor U4095 (N_4095,N_3832,N_3816);
or U4096 (N_4096,N_3898,N_3825);
and U4097 (N_4097,N_3860,N_3958);
nand U4098 (N_4098,N_3850,N_3823);
nor U4099 (N_4099,N_3807,N_3942);
nand U4100 (N_4100,N_3995,N_3829);
nor U4101 (N_4101,N_3826,N_3828);
and U4102 (N_4102,N_3857,N_3864);
nor U4103 (N_4103,N_3891,N_3878);
or U4104 (N_4104,N_3932,N_3837);
or U4105 (N_4105,N_3938,N_3898);
nand U4106 (N_4106,N_3897,N_3891);
and U4107 (N_4107,N_3943,N_3950);
xnor U4108 (N_4108,N_3829,N_3819);
nor U4109 (N_4109,N_3972,N_3994);
or U4110 (N_4110,N_3998,N_3989);
and U4111 (N_4111,N_3978,N_3931);
nand U4112 (N_4112,N_3836,N_3880);
and U4113 (N_4113,N_3897,N_3901);
and U4114 (N_4114,N_3901,N_3958);
or U4115 (N_4115,N_3984,N_3922);
and U4116 (N_4116,N_3974,N_3898);
xnor U4117 (N_4117,N_3925,N_3859);
or U4118 (N_4118,N_3810,N_3819);
or U4119 (N_4119,N_3817,N_3824);
or U4120 (N_4120,N_3890,N_3949);
and U4121 (N_4121,N_3817,N_3915);
and U4122 (N_4122,N_3986,N_3868);
nor U4123 (N_4123,N_3831,N_3965);
nor U4124 (N_4124,N_3833,N_3826);
xnor U4125 (N_4125,N_3906,N_3831);
xnor U4126 (N_4126,N_3828,N_3953);
and U4127 (N_4127,N_3894,N_3967);
nand U4128 (N_4128,N_3930,N_3814);
xor U4129 (N_4129,N_3991,N_3997);
or U4130 (N_4130,N_3862,N_3893);
and U4131 (N_4131,N_3854,N_3930);
nand U4132 (N_4132,N_3922,N_3999);
nand U4133 (N_4133,N_3971,N_3830);
xor U4134 (N_4134,N_3814,N_3862);
or U4135 (N_4135,N_3927,N_3862);
nor U4136 (N_4136,N_3866,N_3889);
xnor U4137 (N_4137,N_3806,N_3858);
nor U4138 (N_4138,N_3860,N_3881);
nor U4139 (N_4139,N_3902,N_3987);
and U4140 (N_4140,N_3917,N_3943);
and U4141 (N_4141,N_3979,N_3934);
or U4142 (N_4142,N_3831,N_3836);
nand U4143 (N_4143,N_3894,N_3825);
nand U4144 (N_4144,N_3946,N_3911);
nand U4145 (N_4145,N_3831,N_3845);
or U4146 (N_4146,N_3930,N_3890);
nand U4147 (N_4147,N_3946,N_3862);
or U4148 (N_4148,N_3923,N_3947);
or U4149 (N_4149,N_3958,N_3826);
nor U4150 (N_4150,N_3866,N_3914);
and U4151 (N_4151,N_3928,N_3957);
and U4152 (N_4152,N_3920,N_3834);
or U4153 (N_4153,N_3968,N_3934);
nand U4154 (N_4154,N_3997,N_3882);
or U4155 (N_4155,N_3817,N_3999);
xor U4156 (N_4156,N_3963,N_3921);
or U4157 (N_4157,N_3856,N_3882);
nor U4158 (N_4158,N_3896,N_3841);
nand U4159 (N_4159,N_3845,N_3975);
xnor U4160 (N_4160,N_3930,N_3981);
and U4161 (N_4161,N_3981,N_3904);
nor U4162 (N_4162,N_3850,N_3913);
nand U4163 (N_4163,N_3938,N_3897);
nand U4164 (N_4164,N_3915,N_3962);
and U4165 (N_4165,N_3863,N_3910);
xnor U4166 (N_4166,N_3951,N_3937);
nor U4167 (N_4167,N_3864,N_3950);
nand U4168 (N_4168,N_3802,N_3944);
xor U4169 (N_4169,N_3918,N_3807);
xor U4170 (N_4170,N_3986,N_3831);
nor U4171 (N_4171,N_3916,N_3966);
or U4172 (N_4172,N_3969,N_3899);
or U4173 (N_4173,N_3867,N_3883);
or U4174 (N_4174,N_3969,N_3805);
nor U4175 (N_4175,N_3839,N_3972);
nor U4176 (N_4176,N_3981,N_3869);
xor U4177 (N_4177,N_3833,N_3987);
xnor U4178 (N_4178,N_3853,N_3912);
nand U4179 (N_4179,N_3930,N_3856);
nand U4180 (N_4180,N_3855,N_3942);
or U4181 (N_4181,N_3917,N_3860);
xor U4182 (N_4182,N_3987,N_3929);
and U4183 (N_4183,N_3976,N_3933);
and U4184 (N_4184,N_3875,N_3833);
or U4185 (N_4185,N_3849,N_3866);
nor U4186 (N_4186,N_3882,N_3957);
or U4187 (N_4187,N_3806,N_3822);
xor U4188 (N_4188,N_3985,N_3978);
and U4189 (N_4189,N_3869,N_3995);
or U4190 (N_4190,N_3910,N_3921);
xor U4191 (N_4191,N_3809,N_3806);
nand U4192 (N_4192,N_3993,N_3945);
or U4193 (N_4193,N_3997,N_3870);
and U4194 (N_4194,N_3985,N_3819);
and U4195 (N_4195,N_3975,N_3849);
or U4196 (N_4196,N_3823,N_3975);
nor U4197 (N_4197,N_3814,N_3840);
nand U4198 (N_4198,N_3976,N_3912);
or U4199 (N_4199,N_3943,N_3819);
and U4200 (N_4200,N_4131,N_4171);
and U4201 (N_4201,N_4032,N_4096);
nand U4202 (N_4202,N_4078,N_4071);
nor U4203 (N_4203,N_4020,N_4007);
nand U4204 (N_4204,N_4187,N_4190);
xor U4205 (N_4205,N_4030,N_4045);
and U4206 (N_4206,N_4092,N_4022);
nor U4207 (N_4207,N_4063,N_4199);
and U4208 (N_4208,N_4049,N_4046);
and U4209 (N_4209,N_4181,N_4158);
and U4210 (N_4210,N_4028,N_4179);
or U4211 (N_4211,N_4129,N_4178);
nand U4212 (N_4212,N_4057,N_4068);
nand U4213 (N_4213,N_4060,N_4184);
xnor U4214 (N_4214,N_4036,N_4140);
xor U4215 (N_4215,N_4152,N_4002);
nor U4216 (N_4216,N_4198,N_4065);
xor U4217 (N_4217,N_4130,N_4144);
nand U4218 (N_4218,N_4070,N_4150);
and U4219 (N_4219,N_4112,N_4061);
or U4220 (N_4220,N_4091,N_4058);
or U4221 (N_4221,N_4004,N_4128);
xor U4222 (N_4222,N_4114,N_4080);
nand U4223 (N_4223,N_4133,N_4172);
or U4224 (N_4224,N_4116,N_4079);
or U4225 (N_4225,N_4182,N_4168);
and U4226 (N_4226,N_4165,N_4166);
and U4227 (N_4227,N_4113,N_4195);
nor U4228 (N_4228,N_4159,N_4154);
nor U4229 (N_4229,N_4126,N_4103);
xor U4230 (N_4230,N_4189,N_4107);
xnor U4231 (N_4231,N_4124,N_4164);
nor U4232 (N_4232,N_4034,N_4169);
nor U4233 (N_4233,N_4017,N_4157);
nand U4234 (N_4234,N_4014,N_4139);
xor U4235 (N_4235,N_4081,N_4136);
nor U4236 (N_4236,N_4194,N_4197);
xor U4237 (N_4237,N_4127,N_4191);
nand U4238 (N_4238,N_4023,N_4118);
or U4239 (N_4239,N_4084,N_4086);
or U4240 (N_4240,N_4097,N_4121);
nand U4241 (N_4241,N_4089,N_4073);
and U4242 (N_4242,N_4055,N_4110);
xnor U4243 (N_4243,N_4115,N_4038);
nor U4244 (N_4244,N_4082,N_4093);
xnor U4245 (N_4245,N_4037,N_4134);
xnor U4246 (N_4246,N_4012,N_4000);
nand U4247 (N_4247,N_4162,N_4156);
or U4248 (N_4248,N_4106,N_4109);
or U4249 (N_4249,N_4026,N_4008);
or U4250 (N_4250,N_4196,N_4027);
and U4251 (N_4251,N_4170,N_4183);
nor U4252 (N_4252,N_4153,N_4040);
nand U4253 (N_4253,N_4192,N_4174);
or U4254 (N_4254,N_4095,N_4039);
or U4255 (N_4255,N_4043,N_4031);
or U4256 (N_4256,N_4138,N_4054);
xnor U4257 (N_4257,N_4076,N_4019);
and U4258 (N_4258,N_4141,N_4016);
and U4259 (N_4259,N_4072,N_4108);
nor U4260 (N_4260,N_4143,N_4033);
nand U4261 (N_4261,N_4025,N_4119);
nand U4262 (N_4262,N_4044,N_4123);
and U4263 (N_4263,N_4132,N_4145);
nand U4264 (N_4264,N_4188,N_4125);
nand U4265 (N_4265,N_4161,N_4035);
nand U4266 (N_4266,N_4105,N_4104);
nand U4267 (N_4267,N_4135,N_4074);
nor U4268 (N_4268,N_4163,N_4180);
nor U4269 (N_4269,N_4160,N_4010);
and U4270 (N_4270,N_4018,N_4193);
and U4271 (N_4271,N_4024,N_4042);
or U4272 (N_4272,N_4186,N_4148);
or U4273 (N_4273,N_4021,N_4069);
nor U4274 (N_4274,N_4142,N_4006);
nand U4275 (N_4275,N_4075,N_4077);
and U4276 (N_4276,N_4117,N_4155);
and U4277 (N_4277,N_4064,N_4146);
or U4278 (N_4278,N_4062,N_4085);
nor U4279 (N_4279,N_4175,N_4011);
nand U4280 (N_4280,N_4098,N_4137);
nand U4281 (N_4281,N_4173,N_4090);
nand U4282 (N_4282,N_4167,N_4056);
nor U4283 (N_4283,N_4094,N_4041);
and U4284 (N_4284,N_4177,N_4088);
nor U4285 (N_4285,N_4013,N_4100);
or U4286 (N_4286,N_4151,N_4101);
or U4287 (N_4287,N_4059,N_4015);
nand U4288 (N_4288,N_4122,N_4005);
xor U4289 (N_4289,N_4185,N_4067);
and U4290 (N_4290,N_4120,N_4102);
or U4291 (N_4291,N_4176,N_4099);
and U4292 (N_4292,N_4009,N_4053);
or U4293 (N_4293,N_4029,N_4047);
and U4294 (N_4294,N_4050,N_4003);
nor U4295 (N_4295,N_4052,N_4111);
nand U4296 (N_4296,N_4048,N_4149);
or U4297 (N_4297,N_4083,N_4001);
xor U4298 (N_4298,N_4051,N_4087);
nor U4299 (N_4299,N_4147,N_4066);
and U4300 (N_4300,N_4057,N_4051);
nor U4301 (N_4301,N_4156,N_4006);
nor U4302 (N_4302,N_4082,N_4094);
nor U4303 (N_4303,N_4121,N_4140);
nor U4304 (N_4304,N_4141,N_4140);
or U4305 (N_4305,N_4157,N_4073);
or U4306 (N_4306,N_4188,N_4071);
or U4307 (N_4307,N_4191,N_4132);
or U4308 (N_4308,N_4032,N_4091);
or U4309 (N_4309,N_4008,N_4090);
nand U4310 (N_4310,N_4065,N_4194);
xor U4311 (N_4311,N_4170,N_4107);
and U4312 (N_4312,N_4130,N_4163);
xor U4313 (N_4313,N_4149,N_4095);
and U4314 (N_4314,N_4178,N_4116);
xor U4315 (N_4315,N_4198,N_4102);
xnor U4316 (N_4316,N_4125,N_4192);
or U4317 (N_4317,N_4023,N_4100);
xnor U4318 (N_4318,N_4198,N_4193);
xnor U4319 (N_4319,N_4180,N_4149);
nand U4320 (N_4320,N_4022,N_4191);
nand U4321 (N_4321,N_4196,N_4157);
and U4322 (N_4322,N_4080,N_4103);
and U4323 (N_4323,N_4161,N_4164);
and U4324 (N_4324,N_4032,N_4063);
nand U4325 (N_4325,N_4118,N_4031);
nand U4326 (N_4326,N_4013,N_4073);
nor U4327 (N_4327,N_4150,N_4196);
xor U4328 (N_4328,N_4163,N_4059);
nand U4329 (N_4329,N_4009,N_4077);
nor U4330 (N_4330,N_4105,N_4167);
nor U4331 (N_4331,N_4108,N_4050);
nand U4332 (N_4332,N_4172,N_4093);
or U4333 (N_4333,N_4103,N_4075);
nor U4334 (N_4334,N_4188,N_4092);
nor U4335 (N_4335,N_4192,N_4170);
xnor U4336 (N_4336,N_4098,N_4032);
xor U4337 (N_4337,N_4169,N_4150);
and U4338 (N_4338,N_4157,N_4104);
or U4339 (N_4339,N_4114,N_4097);
nor U4340 (N_4340,N_4094,N_4120);
nand U4341 (N_4341,N_4161,N_4033);
nor U4342 (N_4342,N_4022,N_4010);
or U4343 (N_4343,N_4043,N_4018);
xnor U4344 (N_4344,N_4025,N_4174);
and U4345 (N_4345,N_4012,N_4032);
nor U4346 (N_4346,N_4198,N_4087);
xnor U4347 (N_4347,N_4080,N_4054);
nand U4348 (N_4348,N_4175,N_4171);
and U4349 (N_4349,N_4007,N_4138);
xnor U4350 (N_4350,N_4119,N_4048);
or U4351 (N_4351,N_4059,N_4025);
and U4352 (N_4352,N_4004,N_4164);
nor U4353 (N_4353,N_4198,N_4034);
xor U4354 (N_4354,N_4126,N_4023);
nor U4355 (N_4355,N_4166,N_4022);
and U4356 (N_4356,N_4072,N_4070);
and U4357 (N_4357,N_4137,N_4125);
nand U4358 (N_4358,N_4058,N_4010);
nand U4359 (N_4359,N_4025,N_4079);
nor U4360 (N_4360,N_4098,N_4142);
nand U4361 (N_4361,N_4052,N_4135);
and U4362 (N_4362,N_4133,N_4159);
xnor U4363 (N_4363,N_4128,N_4131);
nor U4364 (N_4364,N_4048,N_4020);
and U4365 (N_4365,N_4088,N_4024);
xnor U4366 (N_4366,N_4063,N_4026);
xnor U4367 (N_4367,N_4102,N_4163);
nor U4368 (N_4368,N_4021,N_4063);
and U4369 (N_4369,N_4153,N_4127);
nor U4370 (N_4370,N_4175,N_4145);
nor U4371 (N_4371,N_4174,N_4133);
or U4372 (N_4372,N_4162,N_4096);
nor U4373 (N_4373,N_4145,N_4112);
or U4374 (N_4374,N_4026,N_4004);
or U4375 (N_4375,N_4078,N_4056);
or U4376 (N_4376,N_4137,N_4026);
xor U4377 (N_4377,N_4027,N_4148);
nor U4378 (N_4378,N_4007,N_4076);
xor U4379 (N_4379,N_4179,N_4019);
nand U4380 (N_4380,N_4149,N_4196);
and U4381 (N_4381,N_4088,N_4195);
nand U4382 (N_4382,N_4019,N_4015);
and U4383 (N_4383,N_4066,N_4110);
and U4384 (N_4384,N_4130,N_4176);
xnor U4385 (N_4385,N_4046,N_4133);
xnor U4386 (N_4386,N_4052,N_4186);
or U4387 (N_4387,N_4057,N_4134);
and U4388 (N_4388,N_4094,N_4150);
or U4389 (N_4389,N_4164,N_4057);
nor U4390 (N_4390,N_4177,N_4125);
or U4391 (N_4391,N_4107,N_4099);
or U4392 (N_4392,N_4003,N_4055);
nor U4393 (N_4393,N_4094,N_4163);
and U4394 (N_4394,N_4092,N_4196);
xnor U4395 (N_4395,N_4098,N_4105);
nand U4396 (N_4396,N_4103,N_4170);
nor U4397 (N_4397,N_4185,N_4184);
and U4398 (N_4398,N_4045,N_4072);
and U4399 (N_4399,N_4180,N_4045);
nand U4400 (N_4400,N_4263,N_4367);
xor U4401 (N_4401,N_4297,N_4287);
xnor U4402 (N_4402,N_4267,N_4343);
nor U4403 (N_4403,N_4331,N_4283);
and U4404 (N_4404,N_4219,N_4335);
nand U4405 (N_4405,N_4266,N_4216);
xor U4406 (N_4406,N_4278,N_4285);
xor U4407 (N_4407,N_4247,N_4346);
nor U4408 (N_4408,N_4383,N_4341);
nor U4409 (N_4409,N_4249,N_4371);
nor U4410 (N_4410,N_4228,N_4347);
xnor U4411 (N_4411,N_4350,N_4212);
xor U4412 (N_4412,N_4398,N_4245);
nor U4413 (N_4413,N_4234,N_4307);
xor U4414 (N_4414,N_4226,N_4254);
nand U4415 (N_4415,N_4381,N_4227);
xor U4416 (N_4416,N_4310,N_4319);
xor U4417 (N_4417,N_4220,N_4376);
nor U4418 (N_4418,N_4281,N_4391);
and U4419 (N_4419,N_4253,N_4360);
nor U4420 (N_4420,N_4200,N_4368);
nand U4421 (N_4421,N_4255,N_4204);
xor U4422 (N_4422,N_4277,N_4302);
nand U4423 (N_4423,N_4272,N_4221);
or U4424 (N_4424,N_4389,N_4311);
or U4425 (N_4425,N_4237,N_4316);
nor U4426 (N_4426,N_4375,N_4361);
nand U4427 (N_4427,N_4246,N_4329);
xor U4428 (N_4428,N_4348,N_4353);
xor U4429 (N_4429,N_4215,N_4290);
and U4430 (N_4430,N_4224,N_4313);
or U4431 (N_4431,N_4286,N_4328);
nor U4432 (N_4432,N_4233,N_4289);
xor U4433 (N_4433,N_4377,N_4356);
and U4434 (N_4434,N_4336,N_4251);
nand U4435 (N_4435,N_4238,N_4295);
nor U4436 (N_4436,N_4308,N_4303);
xnor U4437 (N_4437,N_4372,N_4355);
or U4438 (N_4438,N_4342,N_4292);
nand U4439 (N_4439,N_4270,N_4325);
and U4440 (N_4440,N_4378,N_4296);
or U4441 (N_4441,N_4257,N_4291);
and U4442 (N_4442,N_4240,N_4248);
nand U4443 (N_4443,N_4206,N_4385);
and U4444 (N_4444,N_4338,N_4304);
xor U4445 (N_4445,N_4274,N_4365);
xor U4446 (N_4446,N_4225,N_4396);
xnor U4447 (N_4447,N_4340,N_4264);
or U4448 (N_4448,N_4258,N_4305);
nand U4449 (N_4449,N_4201,N_4393);
xor U4450 (N_4450,N_4205,N_4299);
or U4451 (N_4451,N_4269,N_4217);
or U4452 (N_4452,N_4364,N_4236);
nand U4453 (N_4453,N_4298,N_4275);
xor U4454 (N_4454,N_4256,N_4394);
nand U4455 (N_4455,N_4207,N_4211);
nor U4456 (N_4456,N_4231,N_4386);
and U4457 (N_4457,N_4244,N_4312);
and U4458 (N_4458,N_4334,N_4326);
xor U4459 (N_4459,N_4242,N_4243);
and U4460 (N_4460,N_4314,N_4384);
nand U4461 (N_4461,N_4259,N_4324);
and U4462 (N_4462,N_4351,N_4323);
xnor U4463 (N_4463,N_4366,N_4229);
xnor U4464 (N_4464,N_4321,N_4306);
nand U4465 (N_4465,N_4260,N_4202);
xnor U4466 (N_4466,N_4210,N_4339);
nand U4467 (N_4467,N_4273,N_4239);
nor U4468 (N_4468,N_4363,N_4379);
xor U4469 (N_4469,N_4344,N_4279);
xnor U4470 (N_4470,N_4284,N_4374);
nand U4471 (N_4471,N_4399,N_4223);
nand U4472 (N_4472,N_4388,N_4230);
nor U4473 (N_4473,N_4349,N_4252);
or U4474 (N_4474,N_4333,N_4222);
or U4475 (N_4475,N_4213,N_4380);
and U4476 (N_4476,N_4352,N_4315);
xnor U4477 (N_4477,N_4276,N_4208);
nor U4478 (N_4478,N_4320,N_4203);
nand U4479 (N_4479,N_4358,N_4293);
or U4480 (N_4480,N_4271,N_4332);
or U4481 (N_4481,N_4280,N_4282);
nor U4482 (N_4482,N_4395,N_4359);
nor U4483 (N_4483,N_4261,N_4390);
nor U4484 (N_4484,N_4214,N_4397);
nand U4485 (N_4485,N_4209,N_4318);
nand U4486 (N_4486,N_4345,N_4235);
nor U4487 (N_4487,N_4250,N_4373);
xor U4488 (N_4488,N_4322,N_4262);
nor U4489 (N_4489,N_4268,N_4317);
nor U4490 (N_4490,N_4327,N_4387);
or U4491 (N_4491,N_4357,N_4370);
nand U4492 (N_4492,N_4232,N_4300);
xor U4493 (N_4493,N_4288,N_4309);
xor U4494 (N_4494,N_4265,N_4241);
nand U4495 (N_4495,N_4301,N_4362);
nor U4496 (N_4496,N_4330,N_4369);
nand U4497 (N_4497,N_4294,N_4337);
nand U4498 (N_4498,N_4218,N_4354);
nor U4499 (N_4499,N_4392,N_4382);
and U4500 (N_4500,N_4256,N_4250);
xnor U4501 (N_4501,N_4327,N_4272);
xor U4502 (N_4502,N_4240,N_4394);
or U4503 (N_4503,N_4380,N_4388);
xor U4504 (N_4504,N_4248,N_4362);
xor U4505 (N_4505,N_4357,N_4270);
nand U4506 (N_4506,N_4300,N_4307);
and U4507 (N_4507,N_4315,N_4383);
or U4508 (N_4508,N_4341,N_4276);
and U4509 (N_4509,N_4283,N_4251);
and U4510 (N_4510,N_4213,N_4356);
nand U4511 (N_4511,N_4305,N_4336);
or U4512 (N_4512,N_4299,N_4394);
nand U4513 (N_4513,N_4247,N_4363);
and U4514 (N_4514,N_4272,N_4258);
nor U4515 (N_4515,N_4257,N_4271);
xor U4516 (N_4516,N_4326,N_4287);
or U4517 (N_4517,N_4362,N_4217);
xor U4518 (N_4518,N_4308,N_4309);
nand U4519 (N_4519,N_4339,N_4285);
nand U4520 (N_4520,N_4386,N_4358);
or U4521 (N_4521,N_4386,N_4365);
or U4522 (N_4522,N_4260,N_4300);
nor U4523 (N_4523,N_4200,N_4399);
nor U4524 (N_4524,N_4271,N_4283);
and U4525 (N_4525,N_4237,N_4205);
nor U4526 (N_4526,N_4285,N_4236);
and U4527 (N_4527,N_4259,N_4392);
and U4528 (N_4528,N_4317,N_4255);
xor U4529 (N_4529,N_4313,N_4394);
nand U4530 (N_4530,N_4349,N_4261);
xor U4531 (N_4531,N_4360,N_4372);
xnor U4532 (N_4532,N_4295,N_4347);
or U4533 (N_4533,N_4347,N_4323);
nand U4534 (N_4534,N_4316,N_4211);
xor U4535 (N_4535,N_4275,N_4349);
xor U4536 (N_4536,N_4230,N_4268);
nor U4537 (N_4537,N_4258,N_4247);
or U4538 (N_4538,N_4208,N_4381);
nor U4539 (N_4539,N_4381,N_4275);
xor U4540 (N_4540,N_4328,N_4267);
nor U4541 (N_4541,N_4306,N_4217);
and U4542 (N_4542,N_4357,N_4356);
nor U4543 (N_4543,N_4388,N_4262);
and U4544 (N_4544,N_4314,N_4343);
nor U4545 (N_4545,N_4245,N_4290);
nor U4546 (N_4546,N_4354,N_4291);
xnor U4547 (N_4547,N_4386,N_4232);
and U4548 (N_4548,N_4264,N_4332);
nor U4549 (N_4549,N_4301,N_4264);
nand U4550 (N_4550,N_4253,N_4260);
nand U4551 (N_4551,N_4373,N_4224);
xor U4552 (N_4552,N_4352,N_4251);
or U4553 (N_4553,N_4243,N_4373);
and U4554 (N_4554,N_4282,N_4213);
and U4555 (N_4555,N_4207,N_4377);
nor U4556 (N_4556,N_4291,N_4317);
and U4557 (N_4557,N_4394,N_4321);
nor U4558 (N_4558,N_4219,N_4307);
and U4559 (N_4559,N_4296,N_4259);
nand U4560 (N_4560,N_4355,N_4309);
and U4561 (N_4561,N_4382,N_4386);
nand U4562 (N_4562,N_4262,N_4217);
nor U4563 (N_4563,N_4233,N_4204);
nor U4564 (N_4564,N_4394,N_4351);
and U4565 (N_4565,N_4242,N_4306);
xor U4566 (N_4566,N_4369,N_4351);
or U4567 (N_4567,N_4274,N_4270);
xor U4568 (N_4568,N_4371,N_4240);
nor U4569 (N_4569,N_4253,N_4390);
nor U4570 (N_4570,N_4326,N_4201);
nor U4571 (N_4571,N_4249,N_4352);
nor U4572 (N_4572,N_4321,N_4354);
or U4573 (N_4573,N_4353,N_4217);
nor U4574 (N_4574,N_4321,N_4206);
and U4575 (N_4575,N_4318,N_4203);
xnor U4576 (N_4576,N_4220,N_4331);
nor U4577 (N_4577,N_4373,N_4289);
nand U4578 (N_4578,N_4355,N_4316);
and U4579 (N_4579,N_4235,N_4260);
or U4580 (N_4580,N_4238,N_4347);
nor U4581 (N_4581,N_4212,N_4387);
nor U4582 (N_4582,N_4239,N_4206);
xor U4583 (N_4583,N_4228,N_4398);
or U4584 (N_4584,N_4268,N_4356);
or U4585 (N_4585,N_4216,N_4201);
and U4586 (N_4586,N_4313,N_4367);
and U4587 (N_4587,N_4242,N_4398);
nand U4588 (N_4588,N_4285,N_4397);
nand U4589 (N_4589,N_4396,N_4243);
or U4590 (N_4590,N_4207,N_4241);
nor U4591 (N_4591,N_4328,N_4268);
xnor U4592 (N_4592,N_4298,N_4212);
nor U4593 (N_4593,N_4230,N_4212);
and U4594 (N_4594,N_4283,N_4372);
and U4595 (N_4595,N_4274,N_4363);
xor U4596 (N_4596,N_4245,N_4222);
xor U4597 (N_4597,N_4204,N_4207);
or U4598 (N_4598,N_4343,N_4237);
xnor U4599 (N_4599,N_4334,N_4320);
nand U4600 (N_4600,N_4407,N_4595);
xor U4601 (N_4601,N_4451,N_4545);
and U4602 (N_4602,N_4598,N_4404);
and U4603 (N_4603,N_4454,N_4422);
xnor U4604 (N_4604,N_4476,N_4468);
or U4605 (N_4605,N_4449,N_4533);
nand U4606 (N_4606,N_4569,N_4535);
nand U4607 (N_4607,N_4578,N_4505);
xor U4608 (N_4608,N_4558,N_4499);
and U4609 (N_4609,N_4594,N_4571);
nor U4610 (N_4610,N_4534,N_4567);
nor U4611 (N_4611,N_4530,N_4450);
xor U4612 (N_4612,N_4587,N_4431);
nor U4613 (N_4613,N_4589,N_4428);
nand U4614 (N_4614,N_4596,N_4421);
nand U4615 (N_4615,N_4577,N_4480);
or U4616 (N_4616,N_4413,N_4478);
xnor U4617 (N_4617,N_4494,N_4455);
and U4618 (N_4618,N_4560,N_4457);
nor U4619 (N_4619,N_4460,N_4441);
or U4620 (N_4620,N_4590,N_4414);
or U4621 (N_4621,N_4511,N_4482);
and U4622 (N_4622,N_4588,N_4469);
nor U4623 (N_4623,N_4408,N_4492);
nor U4624 (N_4624,N_4464,N_4447);
and U4625 (N_4625,N_4437,N_4405);
xor U4626 (N_4626,N_4549,N_4527);
nor U4627 (N_4627,N_4430,N_4591);
xor U4628 (N_4628,N_4575,N_4537);
or U4629 (N_4629,N_4592,N_4593);
nand U4630 (N_4630,N_4419,N_4502);
nor U4631 (N_4631,N_4497,N_4446);
nand U4632 (N_4632,N_4445,N_4459);
and U4633 (N_4633,N_4532,N_4453);
xnor U4634 (N_4634,N_4461,N_4583);
or U4635 (N_4635,N_4529,N_4581);
and U4636 (N_4636,N_4495,N_4542);
and U4637 (N_4637,N_4540,N_4470);
nor U4638 (N_4638,N_4582,N_4429);
nand U4639 (N_4639,N_4481,N_4440);
and U4640 (N_4640,N_4501,N_4550);
or U4641 (N_4641,N_4515,N_4439);
and U4642 (N_4642,N_4516,N_4574);
xor U4643 (N_4643,N_4538,N_4425);
nor U4644 (N_4644,N_4400,N_4521);
nand U4645 (N_4645,N_4472,N_4564);
xor U4646 (N_4646,N_4547,N_4466);
xnor U4647 (N_4647,N_4543,N_4562);
and U4648 (N_4648,N_4403,N_4465);
nand U4649 (N_4649,N_4553,N_4536);
and U4650 (N_4650,N_4576,N_4416);
xor U4651 (N_4651,N_4504,N_4539);
xnor U4652 (N_4652,N_4573,N_4554);
xnor U4653 (N_4653,N_4556,N_4503);
and U4654 (N_4654,N_4493,N_4498);
xnor U4655 (N_4655,N_4597,N_4519);
xnor U4656 (N_4656,N_4496,N_4528);
nand U4657 (N_4657,N_4513,N_4420);
xnor U4658 (N_4658,N_4442,N_4525);
xor U4659 (N_4659,N_4426,N_4572);
nor U4660 (N_4660,N_4483,N_4585);
and U4661 (N_4661,N_4566,N_4415);
nor U4662 (N_4662,N_4402,N_4436);
or U4663 (N_4663,N_4412,N_4586);
xor U4664 (N_4664,N_4584,N_4488);
or U4665 (N_4665,N_4458,N_4444);
xnor U4666 (N_4666,N_4518,N_4435);
nand U4667 (N_4667,N_4401,N_4524);
or U4668 (N_4668,N_4520,N_4599);
nor U4669 (N_4669,N_4555,N_4552);
nand U4670 (N_4670,N_4490,N_4438);
nand U4671 (N_4671,N_4570,N_4448);
nand U4672 (N_4672,N_4563,N_4477);
xor U4673 (N_4673,N_4434,N_4418);
or U4674 (N_4674,N_4484,N_4508);
xor U4675 (N_4675,N_4486,N_4474);
or U4676 (N_4676,N_4541,N_4500);
xor U4677 (N_4677,N_4507,N_4557);
nand U4678 (N_4678,N_4423,N_4411);
nand U4679 (N_4679,N_4544,N_4509);
nor U4680 (N_4680,N_4456,N_4485);
nand U4681 (N_4681,N_4512,N_4565);
or U4682 (N_4682,N_4506,N_4463);
or U4683 (N_4683,N_4410,N_4443);
or U4684 (N_4684,N_4514,N_4432);
and U4685 (N_4685,N_4409,N_4523);
xor U4686 (N_4686,N_4471,N_4473);
xnor U4687 (N_4687,N_4546,N_4548);
xor U4688 (N_4688,N_4561,N_4462);
nand U4689 (N_4689,N_4551,N_4433);
and U4690 (N_4690,N_4475,N_4580);
or U4691 (N_4691,N_4531,N_4517);
nor U4692 (N_4692,N_4487,N_4568);
xor U4693 (N_4693,N_4491,N_4526);
nand U4694 (N_4694,N_4424,N_4522);
and U4695 (N_4695,N_4559,N_4452);
xor U4696 (N_4696,N_4510,N_4479);
nor U4697 (N_4697,N_4489,N_4467);
or U4698 (N_4698,N_4427,N_4579);
and U4699 (N_4699,N_4406,N_4417);
nand U4700 (N_4700,N_4481,N_4593);
nand U4701 (N_4701,N_4440,N_4463);
xor U4702 (N_4702,N_4538,N_4411);
and U4703 (N_4703,N_4400,N_4536);
or U4704 (N_4704,N_4596,N_4471);
or U4705 (N_4705,N_4444,N_4475);
nand U4706 (N_4706,N_4489,N_4554);
xnor U4707 (N_4707,N_4582,N_4518);
nor U4708 (N_4708,N_4484,N_4453);
or U4709 (N_4709,N_4556,N_4468);
or U4710 (N_4710,N_4515,N_4512);
nor U4711 (N_4711,N_4531,N_4536);
xnor U4712 (N_4712,N_4562,N_4432);
xor U4713 (N_4713,N_4597,N_4588);
nand U4714 (N_4714,N_4481,N_4405);
or U4715 (N_4715,N_4493,N_4423);
nor U4716 (N_4716,N_4412,N_4457);
and U4717 (N_4717,N_4488,N_4465);
and U4718 (N_4718,N_4570,N_4510);
xnor U4719 (N_4719,N_4458,N_4501);
xor U4720 (N_4720,N_4449,N_4522);
and U4721 (N_4721,N_4446,N_4439);
nand U4722 (N_4722,N_4534,N_4524);
or U4723 (N_4723,N_4553,N_4511);
xnor U4724 (N_4724,N_4439,N_4556);
nand U4725 (N_4725,N_4536,N_4462);
nor U4726 (N_4726,N_4428,N_4449);
nand U4727 (N_4727,N_4447,N_4400);
nand U4728 (N_4728,N_4454,N_4492);
and U4729 (N_4729,N_4528,N_4553);
xnor U4730 (N_4730,N_4593,N_4522);
nor U4731 (N_4731,N_4526,N_4469);
and U4732 (N_4732,N_4447,N_4414);
nand U4733 (N_4733,N_4584,N_4589);
nor U4734 (N_4734,N_4539,N_4583);
xor U4735 (N_4735,N_4533,N_4479);
or U4736 (N_4736,N_4579,N_4541);
nor U4737 (N_4737,N_4559,N_4557);
or U4738 (N_4738,N_4563,N_4428);
and U4739 (N_4739,N_4527,N_4533);
nand U4740 (N_4740,N_4478,N_4511);
xnor U4741 (N_4741,N_4423,N_4416);
nand U4742 (N_4742,N_4512,N_4550);
nand U4743 (N_4743,N_4583,N_4566);
xnor U4744 (N_4744,N_4576,N_4427);
nand U4745 (N_4745,N_4491,N_4481);
and U4746 (N_4746,N_4432,N_4570);
xor U4747 (N_4747,N_4476,N_4528);
and U4748 (N_4748,N_4408,N_4589);
xnor U4749 (N_4749,N_4441,N_4577);
xor U4750 (N_4750,N_4580,N_4405);
or U4751 (N_4751,N_4535,N_4476);
nand U4752 (N_4752,N_4511,N_4500);
and U4753 (N_4753,N_4497,N_4569);
and U4754 (N_4754,N_4406,N_4579);
nand U4755 (N_4755,N_4518,N_4545);
xnor U4756 (N_4756,N_4585,N_4492);
nor U4757 (N_4757,N_4505,N_4414);
and U4758 (N_4758,N_4474,N_4447);
nor U4759 (N_4759,N_4521,N_4589);
nor U4760 (N_4760,N_4596,N_4536);
and U4761 (N_4761,N_4468,N_4485);
xor U4762 (N_4762,N_4546,N_4571);
nor U4763 (N_4763,N_4475,N_4447);
and U4764 (N_4764,N_4478,N_4544);
nand U4765 (N_4765,N_4531,N_4417);
xnor U4766 (N_4766,N_4581,N_4557);
nor U4767 (N_4767,N_4599,N_4537);
or U4768 (N_4768,N_4591,N_4402);
nand U4769 (N_4769,N_4596,N_4576);
nor U4770 (N_4770,N_4553,N_4581);
xnor U4771 (N_4771,N_4549,N_4593);
xor U4772 (N_4772,N_4463,N_4559);
nand U4773 (N_4773,N_4578,N_4525);
nand U4774 (N_4774,N_4575,N_4496);
and U4775 (N_4775,N_4461,N_4400);
and U4776 (N_4776,N_4470,N_4408);
nor U4777 (N_4777,N_4463,N_4489);
or U4778 (N_4778,N_4485,N_4415);
and U4779 (N_4779,N_4530,N_4548);
or U4780 (N_4780,N_4474,N_4448);
nand U4781 (N_4781,N_4522,N_4486);
nand U4782 (N_4782,N_4430,N_4555);
or U4783 (N_4783,N_4502,N_4409);
nor U4784 (N_4784,N_4495,N_4559);
nand U4785 (N_4785,N_4402,N_4595);
xor U4786 (N_4786,N_4410,N_4478);
nand U4787 (N_4787,N_4438,N_4526);
nand U4788 (N_4788,N_4570,N_4433);
or U4789 (N_4789,N_4417,N_4578);
nand U4790 (N_4790,N_4470,N_4520);
nor U4791 (N_4791,N_4518,N_4446);
xor U4792 (N_4792,N_4542,N_4591);
nor U4793 (N_4793,N_4512,N_4587);
xor U4794 (N_4794,N_4506,N_4514);
and U4795 (N_4795,N_4441,N_4409);
and U4796 (N_4796,N_4485,N_4463);
and U4797 (N_4797,N_4537,N_4466);
xnor U4798 (N_4798,N_4548,N_4492);
nor U4799 (N_4799,N_4517,N_4530);
xnor U4800 (N_4800,N_4690,N_4774);
nand U4801 (N_4801,N_4799,N_4624);
and U4802 (N_4802,N_4603,N_4637);
nand U4803 (N_4803,N_4626,N_4663);
or U4804 (N_4804,N_4751,N_4667);
xnor U4805 (N_4805,N_4662,N_4730);
xnor U4806 (N_4806,N_4771,N_4610);
nor U4807 (N_4807,N_4783,N_4632);
nor U4808 (N_4808,N_4791,N_4782);
and U4809 (N_4809,N_4776,N_4617);
nor U4810 (N_4810,N_4772,N_4759);
nor U4811 (N_4811,N_4789,N_4634);
nor U4812 (N_4812,N_4723,N_4671);
xnor U4813 (N_4813,N_4682,N_4706);
xnor U4814 (N_4814,N_4696,N_4726);
nor U4815 (N_4815,N_4779,N_4633);
or U4816 (N_4816,N_4606,N_4658);
xor U4817 (N_4817,N_4630,N_4736);
nor U4818 (N_4818,N_4786,N_4677);
and U4819 (N_4819,N_4780,N_4763);
nor U4820 (N_4820,N_4672,N_4613);
nor U4821 (N_4821,N_4767,N_4729);
or U4822 (N_4822,N_4614,N_4695);
and U4823 (N_4823,N_4693,N_4708);
nand U4824 (N_4824,N_4732,N_4788);
nand U4825 (N_4825,N_4616,N_4704);
nor U4826 (N_4826,N_4722,N_4664);
and U4827 (N_4827,N_4714,N_4741);
and U4828 (N_4828,N_4660,N_4688);
xnor U4829 (N_4829,N_4620,N_4680);
nor U4830 (N_4830,N_4631,N_4675);
xor U4831 (N_4831,N_4777,N_4798);
nand U4832 (N_4832,N_4654,N_4647);
xor U4833 (N_4833,N_4792,N_4793);
xor U4834 (N_4834,N_4697,N_4773);
nand U4835 (N_4835,N_4754,N_4602);
and U4836 (N_4836,N_4689,N_4756);
nand U4837 (N_4837,N_4797,N_4661);
xnor U4838 (N_4838,N_4643,N_4629);
xnor U4839 (N_4839,N_4796,N_4712);
nor U4840 (N_4840,N_4687,N_4728);
nor U4841 (N_4841,N_4646,N_4642);
xor U4842 (N_4842,N_4638,N_4747);
nor U4843 (N_4843,N_4601,N_4657);
nand U4844 (N_4844,N_4619,N_4676);
and U4845 (N_4845,N_4775,N_4641);
or U4846 (N_4846,N_4769,N_4768);
xor U4847 (N_4847,N_4753,N_4758);
nand U4848 (N_4848,N_4618,N_4713);
and U4849 (N_4849,N_4717,N_4650);
nor U4850 (N_4850,N_4645,N_4757);
xnor U4851 (N_4851,N_4659,N_4770);
and U4852 (N_4852,N_4785,N_4605);
nor U4853 (N_4853,N_4720,N_4765);
and U4854 (N_4854,N_4694,N_4679);
nand U4855 (N_4855,N_4703,N_4738);
nand U4856 (N_4856,N_4653,N_4692);
xor U4857 (N_4857,N_4656,N_4790);
nand U4858 (N_4858,N_4673,N_4764);
or U4859 (N_4859,N_4752,N_4609);
and U4860 (N_4860,N_4625,N_4746);
or U4861 (N_4861,N_4795,N_4686);
or U4862 (N_4862,N_4719,N_4607);
xor U4863 (N_4863,N_4627,N_4685);
xor U4864 (N_4864,N_4784,N_4745);
nand U4865 (N_4865,N_4743,N_4702);
xnor U4866 (N_4866,N_4623,N_4781);
xnor U4867 (N_4867,N_4611,N_4621);
nand U4868 (N_4868,N_4698,N_4762);
or U4869 (N_4869,N_4651,N_4794);
nor U4870 (N_4870,N_4724,N_4665);
nand U4871 (N_4871,N_4640,N_4750);
and U4872 (N_4872,N_4669,N_4715);
xor U4873 (N_4873,N_4734,N_4612);
or U4874 (N_4874,N_4766,N_4749);
nand U4875 (N_4875,N_4716,N_4666);
xnor U4876 (N_4876,N_4733,N_4615);
xor U4877 (N_4877,N_4725,N_4684);
and U4878 (N_4878,N_4635,N_4721);
nand U4879 (N_4879,N_4622,N_4655);
or U4880 (N_4880,N_4760,N_4636);
or U4881 (N_4881,N_4710,N_4644);
xnor U4882 (N_4882,N_4648,N_4707);
or U4883 (N_4883,N_4639,N_4755);
nor U4884 (N_4884,N_4674,N_4740);
or U4885 (N_4885,N_4668,N_4737);
and U4886 (N_4886,N_4718,N_4731);
nor U4887 (N_4887,N_4705,N_4787);
or U4888 (N_4888,N_4699,N_4700);
xnor U4889 (N_4889,N_4735,N_4670);
nand U4890 (N_4890,N_4739,N_4709);
or U4891 (N_4891,N_4691,N_4778);
and U4892 (N_4892,N_4604,N_4681);
xnor U4893 (N_4893,N_4761,N_4678);
xor U4894 (N_4894,N_4742,N_4744);
nand U4895 (N_4895,N_4600,N_4701);
xor U4896 (N_4896,N_4649,N_4711);
nand U4897 (N_4897,N_4652,N_4608);
nor U4898 (N_4898,N_4628,N_4683);
and U4899 (N_4899,N_4748,N_4727);
nand U4900 (N_4900,N_4765,N_4700);
nor U4901 (N_4901,N_4611,N_4784);
nor U4902 (N_4902,N_4646,N_4645);
nand U4903 (N_4903,N_4725,N_4764);
nand U4904 (N_4904,N_4685,N_4676);
xnor U4905 (N_4905,N_4736,N_4760);
nand U4906 (N_4906,N_4676,N_4630);
nand U4907 (N_4907,N_4755,N_4722);
nor U4908 (N_4908,N_4606,N_4746);
and U4909 (N_4909,N_4656,N_4696);
or U4910 (N_4910,N_4720,N_4760);
or U4911 (N_4911,N_4630,N_4739);
and U4912 (N_4912,N_4627,N_4694);
or U4913 (N_4913,N_4680,N_4776);
or U4914 (N_4914,N_4767,N_4670);
nand U4915 (N_4915,N_4755,N_4717);
nand U4916 (N_4916,N_4797,N_4645);
nand U4917 (N_4917,N_4682,N_4739);
nand U4918 (N_4918,N_4745,N_4686);
and U4919 (N_4919,N_4792,N_4786);
nor U4920 (N_4920,N_4727,N_4771);
and U4921 (N_4921,N_4636,N_4695);
or U4922 (N_4922,N_4792,N_4624);
or U4923 (N_4923,N_4761,N_4693);
and U4924 (N_4924,N_4656,N_4703);
nand U4925 (N_4925,N_4665,N_4700);
nor U4926 (N_4926,N_4615,N_4708);
nor U4927 (N_4927,N_4651,N_4726);
and U4928 (N_4928,N_4621,N_4645);
nand U4929 (N_4929,N_4645,N_4728);
and U4930 (N_4930,N_4778,N_4675);
nand U4931 (N_4931,N_4633,N_4670);
or U4932 (N_4932,N_4785,N_4787);
xnor U4933 (N_4933,N_4792,N_4719);
xnor U4934 (N_4934,N_4734,N_4646);
nor U4935 (N_4935,N_4652,N_4765);
and U4936 (N_4936,N_4704,N_4731);
or U4937 (N_4937,N_4708,N_4773);
xnor U4938 (N_4938,N_4614,N_4697);
or U4939 (N_4939,N_4698,N_4723);
or U4940 (N_4940,N_4618,N_4789);
and U4941 (N_4941,N_4630,N_4619);
nor U4942 (N_4942,N_4731,N_4788);
xnor U4943 (N_4943,N_4682,N_4727);
nand U4944 (N_4944,N_4756,N_4608);
nand U4945 (N_4945,N_4717,N_4648);
nand U4946 (N_4946,N_4740,N_4671);
and U4947 (N_4947,N_4726,N_4670);
nand U4948 (N_4948,N_4752,N_4740);
or U4949 (N_4949,N_4745,N_4759);
or U4950 (N_4950,N_4612,N_4790);
nand U4951 (N_4951,N_4651,N_4775);
or U4952 (N_4952,N_4713,N_4644);
and U4953 (N_4953,N_4790,N_4630);
xnor U4954 (N_4954,N_4608,N_4643);
nor U4955 (N_4955,N_4746,N_4731);
nor U4956 (N_4956,N_4676,N_4799);
nor U4957 (N_4957,N_4766,N_4727);
nor U4958 (N_4958,N_4636,N_4657);
or U4959 (N_4959,N_4724,N_4703);
nor U4960 (N_4960,N_4632,N_4757);
and U4961 (N_4961,N_4636,N_4697);
nor U4962 (N_4962,N_4707,N_4705);
nor U4963 (N_4963,N_4772,N_4767);
xnor U4964 (N_4964,N_4772,N_4755);
nor U4965 (N_4965,N_4695,N_4660);
or U4966 (N_4966,N_4731,N_4712);
xnor U4967 (N_4967,N_4702,N_4706);
or U4968 (N_4968,N_4648,N_4635);
nor U4969 (N_4969,N_4665,N_4723);
xor U4970 (N_4970,N_4716,N_4658);
or U4971 (N_4971,N_4789,N_4637);
and U4972 (N_4972,N_4764,N_4601);
or U4973 (N_4973,N_4607,N_4675);
nand U4974 (N_4974,N_4706,N_4720);
or U4975 (N_4975,N_4795,N_4637);
nor U4976 (N_4976,N_4664,N_4787);
and U4977 (N_4977,N_4677,N_4615);
or U4978 (N_4978,N_4745,N_4742);
xnor U4979 (N_4979,N_4614,N_4625);
and U4980 (N_4980,N_4613,N_4782);
xor U4981 (N_4981,N_4716,N_4628);
and U4982 (N_4982,N_4746,N_4735);
and U4983 (N_4983,N_4782,N_4719);
nand U4984 (N_4984,N_4681,N_4608);
nor U4985 (N_4985,N_4724,N_4693);
xnor U4986 (N_4986,N_4790,N_4717);
nor U4987 (N_4987,N_4651,N_4797);
and U4988 (N_4988,N_4698,N_4704);
or U4989 (N_4989,N_4670,N_4792);
and U4990 (N_4990,N_4720,N_4781);
xnor U4991 (N_4991,N_4704,N_4674);
nand U4992 (N_4992,N_4687,N_4736);
xor U4993 (N_4993,N_4773,N_4775);
xor U4994 (N_4994,N_4695,N_4716);
nand U4995 (N_4995,N_4726,N_4644);
xnor U4996 (N_4996,N_4627,N_4659);
and U4997 (N_4997,N_4656,N_4761);
or U4998 (N_4998,N_4617,N_4778);
xor U4999 (N_4999,N_4655,N_4625);
and U5000 (N_5000,N_4846,N_4813);
and U5001 (N_5001,N_4832,N_4937);
or U5002 (N_5002,N_4910,N_4814);
and U5003 (N_5003,N_4938,N_4824);
nand U5004 (N_5004,N_4868,N_4927);
xor U5005 (N_5005,N_4969,N_4879);
xor U5006 (N_5006,N_4838,N_4958);
nand U5007 (N_5007,N_4944,N_4894);
and U5008 (N_5008,N_4989,N_4892);
or U5009 (N_5009,N_4970,N_4951);
and U5010 (N_5010,N_4851,N_4926);
nor U5011 (N_5011,N_4804,N_4901);
xor U5012 (N_5012,N_4835,N_4845);
nor U5013 (N_5013,N_4922,N_4872);
nand U5014 (N_5014,N_4850,N_4802);
nor U5015 (N_5015,N_4923,N_4945);
and U5016 (N_5016,N_4964,N_4997);
nor U5017 (N_5017,N_4909,N_4823);
or U5018 (N_5018,N_4856,N_4891);
and U5019 (N_5019,N_4866,N_4956);
nand U5020 (N_5020,N_4896,N_4864);
nand U5021 (N_5021,N_4943,N_4819);
or U5022 (N_5022,N_4820,N_4967);
nor U5023 (N_5023,N_4899,N_4890);
xor U5024 (N_5024,N_4809,N_4829);
and U5025 (N_5025,N_4998,N_4936);
or U5026 (N_5026,N_4827,N_4925);
nor U5027 (N_5027,N_4912,N_4844);
or U5028 (N_5028,N_4918,N_4875);
nand U5029 (N_5029,N_4911,N_4980);
nor U5030 (N_5030,N_4994,N_4990);
or U5031 (N_5031,N_4897,N_4984);
and U5032 (N_5032,N_4859,N_4807);
nor U5033 (N_5033,N_4975,N_4940);
nor U5034 (N_5034,N_4884,N_4839);
and U5035 (N_5035,N_4954,N_4916);
nor U5036 (N_5036,N_4905,N_4817);
xnor U5037 (N_5037,N_4948,N_4983);
nand U5038 (N_5038,N_4834,N_4867);
and U5039 (N_5039,N_4853,N_4836);
nand U5040 (N_5040,N_4955,N_4855);
or U5041 (N_5041,N_4881,N_4965);
or U5042 (N_5042,N_4914,N_4908);
xor U5043 (N_5043,N_4800,N_4935);
xnor U5044 (N_5044,N_4987,N_4822);
or U5045 (N_5045,N_4963,N_4842);
nand U5046 (N_5046,N_4885,N_4833);
or U5047 (N_5047,N_4886,N_4981);
or U5048 (N_5048,N_4883,N_4826);
xnor U5049 (N_5049,N_4862,N_4825);
nor U5050 (N_5050,N_4803,N_4861);
nand U5051 (N_5051,N_4888,N_4860);
or U5052 (N_5052,N_4929,N_4995);
nand U5053 (N_5053,N_4830,N_4960);
xor U5054 (N_5054,N_4934,N_4931);
and U5055 (N_5055,N_4808,N_4852);
or U5056 (N_5056,N_4977,N_4810);
and U5057 (N_5057,N_4873,N_4831);
or U5058 (N_5058,N_4928,N_4828);
or U5059 (N_5059,N_4816,N_4843);
and U5060 (N_5060,N_4917,N_4974);
xor U5061 (N_5061,N_4976,N_4882);
and U5062 (N_5062,N_4870,N_4930);
nor U5063 (N_5063,N_4993,N_4871);
and U5064 (N_5064,N_4887,N_4840);
and U5065 (N_5065,N_4973,N_4919);
xor U5066 (N_5066,N_4996,N_4847);
or U5067 (N_5067,N_4818,N_4992);
nand U5068 (N_5068,N_4821,N_4904);
nand U5069 (N_5069,N_4906,N_4986);
xnor U5070 (N_5070,N_4968,N_4915);
or U5071 (N_5071,N_4920,N_4982);
xor U5072 (N_5072,N_4950,N_4921);
nor U5073 (N_5073,N_4877,N_4913);
and U5074 (N_5074,N_4869,N_4893);
nor U5075 (N_5075,N_4952,N_4941);
xnor U5076 (N_5076,N_4900,N_4863);
nand U5077 (N_5077,N_4876,N_4895);
xor U5078 (N_5078,N_4957,N_4949);
or U5079 (N_5079,N_4801,N_4880);
xnor U5080 (N_5080,N_4959,N_4857);
nor U5081 (N_5081,N_4878,N_4946);
nand U5082 (N_5082,N_4966,N_4972);
nor U5083 (N_5083,N_4854,N_4837);
and U5084 (N_5084,N_4979,N_4812);
or U5085 (N_5085,N_4902,N_4815);
nor U5086 (N_5086,N_4999,N_4805);
or U5087 (N_5087,N_4933,N_4898);
nand U5088 (N_5088,N_4874,N_4841);
nand U5089 (N_5089,N_4961,N_4924);
nand U5090 (N_5090,N_4947,N_4848);
and U5091 (N_5091,N_4865,N_4991);
or U5092 (N_5092,N_4978,N_4988);
xor U5093 (N_5093,N_4858,N_4971);
xor U5094 (N_5094,N_4932,N_4939);
nor U5095 (N_5095,N_4953,N_4811);
or U5096 (N_5096,N_4907,N_4942);
or U5097 (N_5097,N_4962,N_4806);
nand U5098 (N_5098,N_4889,N_4985);
or U5099 (N_5099,N_4849,N_4903);
and U5100 (N_5100,N_4941,N_4845);
nand U5101 (N_5101,N_4921,N_4975);
and U5102 (N_5102,N_4900,N_4880);
or U5103 (N_5103,N_4953,N_4895);
xnor U5104 (N_5104,N_4867,N_4800);
or U5105 (N_5105,N_4801,N_4815);
nor U5106 (N_5106,N_4842,N_4806);
or U5107 (N_5107,N_4973,N_4915);
nand U5108 (N_5108,N_4813,N_4948);
nor U5109 (N_5109,N_4816,N_4908);
or U5110 (N_5110,N_4954,N_4928);
xnor U5111 (N_5111,N_4926,N_4882);
or U5112 (N_5112,N_4825,N_4801);
nand U5113 (N_5113,N_4955,N_4908);
nand U5114 (N_5114,N_4831,N_4986);
nor U5115 (N_5115,N_4934,N_4885);
xnor U5116 (N_5116,N_4841,N_4958);
and U5117 (N_5117,N_4874,N_4956);
and U5118 (N_5118,N_4976,N_4960);
xnor U5119 (N_5119,N_4949,N_4956);
or U5120 (N_5120,N_4865,N_4906);
xor U5121 (N_5121,N_4802,N_4845);
or U5122 (N_5122,N_4971,N_4959);
xnor U5123 (N_5123,N_4988,N_4937);
nand U5124 (N_5124,N_4862,N_4994);
or U5125 (N_5125,N_4969,N_4946);
nor U5126 (N_5126,N_4854,N_4924);
xor U5127 (N_5127,N_4981,N_4997);
or U5128 (N_5128,N_4960,N_4968);
or U5129 (N_5129,N_4962,N_4814);
or U5130 (N_5130,N_4839,N_4961);
and U5131 (N_5131,N_4949,N_4832);
and U5132 (N_5132,N_4886,N_4949);
and U5133 (N_5133,N_4839,N_4906);
xnor U5134 (N_5134,N_4863,N_4913);
and U5135 (N_5135,N_4902,N_4985);
nor U5136 (N_5136,N_4894,N_4920);
or U5137 (N_5137,N_4911,N_4872);
and U5138 (N_5138,N_4867,N_4812);
or U5139 (N_5139,N_4885,N_4828);
nand U5140 (N_5140,N_4956,N_4899);
xor U5141 (N_5141,N_4932,N_4809);
nand U5142 (N_5142,N_4803,N_4993);
or U5143 (N_5143,N_4935,N_4884);
or U5144 (N_5144,N_4947,N_4909);
nor U5145 (N_5145,N_4905,N_4947);
and U5146 (N_5146,N_4894,N_4851);
nand U5147 (N_5147,N_4915,N_4854);
xnor U5148 (N_5148,N_4981,N_4900);
xnor U5149 (N_5149,N_4853,N_4934);
nand U5150 (N_5150,N_4886,N_4941);
nor U5151 (N_5151,N_4994,N_4840);
nor U5152 (N_5152,N_4925,N_4902);
or U5153 (N_5153,N_4955,N_4944);
nand U5154 (N_5154,N_4873,N_4912);
nor U5155 (N_5155,N_4941,N_4972);
nor U5156 (N_5156,N_4861,N_4935);
nand U5157 (N_5157,N_4946,N_4897);
and U5158 (N_5158,N_4813,N_4912);
xor U5159 (N_5159,N_4888,N_4826);
nand U5160 (N_5160,N_4848,N_4847);
and U5161 (N_5161,N_4950,N_4887);
or U5162 (N_5162,N_4859,N_4950);
and U5163 (N_5163,N_4850,N_4824);
or U5164 (N_5164,N_4805,N_4849);
and U5165 (N_5165,N_4936,N_4803);
or U5166 (N_5166,N_4994,N_4969);
nor U5167 (N_5167,N_4819,N_4841);
or U5168 (N_5168,N_4991,N_4898);
nor U5169 (N_5169,N_4858,N_4805);
nor U5170 (N_5170,N_4901,N_4803);
nand U5171 (N_5171,N_4827,N_4877);
or U5172 (N_5172,N_4965,N_4952);
xor U5173 (N_5173,N_4959,N_4946);
nor U5174 (N_5174,N_4903,N_4883);
nor U5175 (N_5175,N_4840,N_4846);
xnor U5176 (N_5176,N_4916,N_4997);
nand U5177 (N_5177,N_4843,N_4916);
nor U5178 (N_5178,N_4845,N_4987);
nand U5179 (N_5179,N_4943,N_4849);
and U5180 (N_5180,N_4981,N_4994);
nand U5181 (N_5181,N_4939,N_4846);
or U5182 (N_5182,N_4846,N_4841);
or U5183 (N_5183,N_4976,N_4894);
and U5184 (N_5184,N_4990,N_4809);
xnor U5185 (N_5185,N_4942,N_4912);
and U5186 (N_5186,N_4901,N_4863);
nand U5187 (N_5187,N_4804,N_4831);
and U5188 (N_5188,N_4924,N_4818);
or U5189 (N_5189,N_4857,N_4813);
and U5190 (N_5190,N_4801,N_4831);
or U5191 (N_5191,N_4978,N_4948);
xor U5192 (N_5192,N_4937,N_4900);
nor U5193 (N_5193,N_4936,N_4900);
nor U5194 (N_5194,N_4886,N_4939);
nor U5195 (N_5195,N_4832,N_4910);
xor U5196 (N_5196,N_4934,N_4835);
nor U5197 (N_5197,N_4940,N_4927);
or U5198 (N_5198,N_4854,N_4861);
or U5199 (N_5199,N_4980,N_4998);
nor U5200 (N_5200,N_5165,N_5152);
and U5201 (N_5201,N_5069,N_5123);
nand U5202 (N_5202,N_5145,N_5048);
xor U5203 (N_5203,N_5157,N_5040);
xor U5204 (N_5204,N_5054,N_5044);
nand U5205 (N_5205,N_5004,N_5088);
xor U5206 (N_5206,N_5177,N_5128);
nor U5207 (N_5207,N_5050,N_5045);
nand U5208 (N_5208,N_5108,N_5019);
or U5209 (N_5209,N_5011,N_5194);
nand U5210 (N_5210,N_5083,N_5167);
xor U5211 (N_5211,N_5161,N_5066);
or U5212 (N_5212,N_5105,N_5084);
or U5213 (N_5213,N_5012,N_5160);
and U5214 (N_5214,N_5110,N_5116);
nor U5215 (N_5215,N_5133,N_5068);
or U5216 (N_5216,N_5016,N_5117);
nand U5217 (N_5217,N_5013,N_5008);
and U5218 (N_5218,N_5173,N_5111);
nor U5219 (N_5219,N_5005,N_5071);
nor U5220 (N_5220,N_5080,N_5026);
nor U5221 (N_5221,N_5073,N_5057);
and U5222 (N_5222,N_5086,N_5039);
nor U5223 (N_5223,N_5020,N_5169);
or U5224 (N_5224,N_5126,N_5132);
or U5225 (N_5225,N_5112,N_5082);
or U5226 (N_5226,N_5055,N_5154);
nand U5227 (N_5227,N_5017,N_5127);
nand U5228 (N_5228,N_5058,N_5076);
and U5229 (N_5229,N_5081,N_5085);
nor U5230 (N_5230,N_5174,N_5130);
and U5231 (N_5231,N_5183,N_5053);
and U5232 (N_5232,N_5035,N_5092);
nor U5233 (N_5233,N_5182,N_5185);
nand U5234 (N_5234,N_5029,N_5122);
nand U5235 (N_5235,N_5024,N_5023);
nor U5236 (N_5236,N_5119,N_5135);
xnor U5237 (N_5237,N_5078,N_5032);
nor U5238 (N_5238,N_5056,N_5146);
and U5239 (N_5239,N_5001,N_5179);
xnor U5240 (N_5240,N_5198,N_5060);
or U5241 (N_5241,N_5140,N_5103);
nand U5242 (N_5242,N_5137,N_5037);
and U5243 (N_5243,N_5094,N_5106);
nand U5244 (N_5244,N_5124,N_5079);
xnor U5245 (N_5245,N_5193,N_5155);
xor U5246 (N_5246,N_5100,N_5148);
nor U5247 (N_5247,N_5187,N_5028);
nand U5248 (N_5248,N_5150,N_5107);
nand U5249 (N_5249,N_5000,N_5136);
nor U5250 (N_5250,N_5034,N_5125);
xnor U5251 (N_5251,N_5170,N_5061);
and U5252 (N_5252,N_5180,N_5063);
nand U5253 (N_5253,N_5030,N_5093);
or U5254 (N_5254,N_5186,N_5134);
nor U5255 (N_5255,N_5062,N_5025);
or U5256 (N_5256,N_5049,N_5188);
nor U5257 (N_5257,N_5065,N_5118);
nor U5258 (N_5258,N_5052,N_5164);
xnor U5259 (N_5259,N_5087,N_5070);
nor U5260 (N_5260,N_5036,N_5131);
nor U5261 (N_5261,N_5089,N_5099);
or U5262 (N_5262,N_5181,N_5163);
nand U5263 (N_5263,N_5021,N_5144);
nand U5264 (N_5264,N_5149,N_5009);
nor U5265 (N_5265,N_5151,N_5172);
nand U5266 (N_5266,N_5038,N_5072);
nand U5267 (N_5267,N_5095,N_5033);
nor U5268 (N_5268,N_5147,N_5158);
nor U5269 (N_5269,N_5046,N_5102);
xor U5270 (N_5270,N_5113,N_5097);
nand U5271 (N_5271,N_5031,N_5143);
and U5272 (N_5272,N_5098,N_5014);
nand U5273 (N_5273,N_5153,N_5006);
or U5274 (N_5274,N_5109,N_5115);
nor U5275 (N_5275,N_5010,N_5042);
or U5276 (N_5276,N_5199,N_5190);
nand U5277 (N_5277,N_5007,N_5168);
and U5278 (N_5278,N_5139,N_5197);
nor U5279 (N_5279,N_5101,N_5015);
and U5280 (N_5280,N_5043,N_5002);
xnor U5281 (N_5281,N_5184,N_5192);
nor U5282 (N_5282,N_5178,N_5176);
and U5283 (N_5283,N_5196,N_5075);
or U5284 (N_5284,N_5141,N_5156);
or U5285 (N_5285,N_5077,N_5041);
and U5286 (N_5286,N_5027,N_5090);
nor U5287 (N_5287,N_5067,N_5104);
nand U5288 (N_5288,N_5129,N_5142);
nand U5289 (N_5289,N_5003,N_5121);
or U5290 (N_5290,N_5091,N_5166);
nand U5291 (N_5291,N_5175,N_5195);
and U5292 (N_5292,N_5191,N_5074);
nand U5293 (N_5293,N_5114,N_5096);
and U5294 (N_5294,N_5171,N_5051);
nand U5295 (N_5295,N_5189,N_5159);
or U5296 (N_5296,N_5047,N_5059);
xnor U5297 (N_5297,N_5064,N_5138);
and U5298 (N_5298,N_5022,N_5162);
and U5299 (N_5299,N_5120,N_5018);
xnor U5300 (N_5300,N_5130,N_5159);
nand U5301 (N_5301,N_5000,N_5077);
or U5302 (N_5302,N_5047,N_5193);
and U5303 (N_5303,N_5078,N_5086);
nand U5304 (N_5304,N_5055,N_5068);
nor U5305 (N_5305,N_5112,N_5199);
nor U5306 (N_5306,N_5173,N_5085);
or U5307 (N_5307,N_5137,N_5096);
or U5308 (N_5308,N_5121,N_5146);
nor U5309 (N_5309,N_5060,N_5073);
nor U5310 (N_5310,N_5107,N_5138);
nor U5311 (N_5311,N_5043,N_5106);
nand U5312 (N_5312,N_5137,N_5092);
nor U5313 (N_5313,N_5095,N_5129);
nand U5314 (N_5314,N_5030,N_5151);
nand U5315 (N_5315,N_5005,N_5077);
nor U5316 (N_5316,N_5146,N_5128);
nor U5317 (N_5317,N_5156,N_5018);
nand U5318 (N_5318,N_5174,N_5111);
nand U5319 (N_5319,N_5123,N_5180);
nand U5320 (N_5320,N_5106,N_5114);
xnor U5321 (N_5321,N_5016,N_5000);
nor U5322 (N_5322,N_5158,N_5097);
or U5323 (N_5323,N_5029,N_5143);
and U5324 (N_5324,N_5006,N_5163);
nor U5325 (N_5325,N_5191,N_5004);
nand U5326 (N_5326,N_5006,N_5162);
or U5327 (N_5327,N_5189,N_5116);
or U5328 (N_5328,N_5039,N_5156);
and U5329 (N_5329,N_5192,N_5165);
and U5330 (N_5330,N_5016,N_5115);
or U5331 (N_5331,N_5052,N_5114);
nand U5332 (N_5332,N_5022,N_5044);
nand U5333 (N_5333,N_5096,N_5103);
xnor U5334 (N_5334,N_5163,N_5100);
nand U5335 (N_5335,N_5107,N_5128);
nand U5336 (N_5336,N_5012,N_5193);
xor U5337 (N_5337,N_5000,N_5020);
and U5338 (N_5338,N_5192,N_5164);
nor U5339 (N_5339,N_5185,N_5079);
and U5340 (N_5340,N_5030,N_5197);
or U5341 (N_5341,N_5088,N_5103);
nor U5342 (N_5342,N_5095,N_5171);
or U5343 (N_5343,N_5045,N_5022);
or U5344 (N_5344,N_5044,N_5162);
or U5345 (N_5345,N_5083,N_5057);
nand U5346 (N_5346,N_5172,N_5020);
nand U5347 (N_5347,N_5130,N_5044);
xor U5348 (N_5348,N_5176,N_5033);
and U5349 (N_5349,N_5009,N_5158);
nand U5350 (N_5350,N_5059,N_5188);
and U5351 (N_5351,N_5133,N_5111);
nor U5352 (N_5352,N_5116,N_5030);
nor U5353 (N_5353,N_5181,N_5061);
nand U5354 (N_5354,N_5112,N_5027);
xor U5355 (N_5355,N_5176,N_5030);
or U5356 (N_5356,N_5195,N_5145);
or U5357 (N_5357,N_5077,N_5094);
and U5358 (N_5358,N_5152,N_5158);
nand U5359 (N_5359,N_5158,N_5055);
nand U5360 (N_5360,N_5173,N_5079);
xnor U5361 (N_5361,N_5154,N_5156);
and U5362 (N_5362,N_5069,N_5050);
xor U5363 (N_5363,N_5137,N_5097);
and U5364 (N_5364,N_5049,N_5035);
or U5365 (N_5365,N_5139,N_5028);
xnor U5366 (N_5366,N_5108,N_5189);
nor U5367 (N_5367,N_5006,N_5009);
xnor U5368 (N_5368,N_5067,N_5123);
and U5369 (N_5369,N_5093,N_5130);
and U5370 (N_5370,N_5106,N_5127);
xor U5371 (N_5371,N_5152,N_5009);
nor U5372 (N_5372,N_5007,N_5035);
nand U5373 (N_5373,N_5063,N_5090);
nand U5374 (N_5374,N_5087,N_5198);
nand U5375 (N_5375,N_5130,N_5170);
nor U5376 (N_5376,N_5058,N_5116);
nand U5377 (N_5377,N_5108,N_5149);
and U5378 (N_5378,N_5198,N_5050);
xnor U5379 (N_5379,N_5170,N_5137);
and U5380 (N_5380,N_5001,N_5009);
nand U5381 (N_5381,N_5042,N_5149);
and U5382 (N_5382,N_5165,N_5076);
or U5383 (N_5383,N_5080,N_5178);
nand U5384 (N_5384,N_5089,N_5072);
and U5385 (N_5385,N_5101,N_5053);
nand U5386 (N_5386,N_5067,N_5029);
xor U5387 (N_5387,N_5085,N_5113);
xor U5388 (N_5388,N_5056,N_5152);
and U5389 (N_5389,N_5078,N_5111);
xor U5390 (N_5390,N_5027,N_5073);
nor U5391 (N_5391,N_5159,N_5069);
nand U5392 (N_5392,N_5101,N_5092);
or U5393 (N_5393,N_5080,N_5170);
and U5394 (N_5394,N_5024,N_5123);
xor U5395 (N_5395,N_5183,N_5143);
or U5396 (N_5396,N_5146,N_5116);
or U5397 (N_5397,N_5164,N_5051);
nand U5398 (N_5398,N_5175,N_5164);
nor U5399 (N_5399,N_5139,N_5168);
nor U5400 (N_5400,N_5399,N_5309);
nor U5401 (N_5401,N_5234,N_5271);
and U5402 (N_5402,N_5252,N_5343);
and U5403 (N_5403,N_5257,N_5268);
nor U5404 (N_5404,N_5283,N_5344);
nor U5405 (N_5405,N_5236,N_5266);
xor U5406 (N_5406,N_5205,N_5259);
nand U5407 (N_5407,N_5241,N_5233);
nand U5408 (N_5408,N_5333,N_5210);
nor U5409 (N_5409,N_5287,N_5227);
or U5410 (N_5410,N_5381,N_5207);
xor U5411 (N_5411,N_5367,N_5388);
or U5412 (N_5412,N_5382,N_5330);
and U5413 (N_5413,N_5345,N_5229);
and U5414 (N_5414,N_5292,N_5261);
or U5415 (N_5415,N_5201,N_5384);
and U5416 (N_5416,N_5276,N_5238);
and U5417 (N_5417,N_5231,N_5264);
and U5418 (N_5418,N_5211,N_5249);
xnor U5419 (N_5419,N_5397,N_5281);
or U5420 (N_5420,N_5258,N_5293);
or U5421 (N_5421,N_5341,N_5306);
or U5422 (N_5422,N_5346,N_5393);
nor U5423 (N_5423,N_5314,N_5312);
xnor U5424 (N_5424,N_5379,N_5360);
and U5425 (N_5425,N_5365,N_5350);
and U5426 (N_5426,N_5377,N_5375);
nor U5427 (N_5427,N_5316,N_5349);
nand U5428 (N_5428,N_5369,N_5226);
nand U5429 (N_5429,N_5278,N_5364);
nand U5430 (N_5430,N_5300,N_5396);
xor U5431 (N_5431,N_5325,N_5298);
nor U5432 (N_5432,N_5255,N_5270);
nor U5433 (N_5433,N_5215,N_5395);
or U5434 (N_5434,N_5353,N_5222);
and U5435 (N_5435,N_5317,N_5336);
or U5436 (N_5436,N_5357,N_5260);
nand U5437 (N_5437,N_5262,N_5244);
or U5438 (N_5438,N_5319,N_5321);
nand U5439 (N_5439,N_5368,N_5214);
or U5440 (N_5440,N_5294,N_5256);
and U5441 (N_5441,N_5221,N_5303);
nand U5442 (N_5442,N_5323,N_5310);
nand U5443 (N_5443,N_5359,N_5254);
or U5444 (N_5444,N_5200,N_5340);
nor U5445 (N_5445,N_5206,N_5237);
nor U5446 (N_5446,N_5232,N_5263);
nor U5447 (N_5447,N_5394,N_5354);
nor U5448 (N_5448,N_5302,N_5253);
nor U5449 (N_5449,N_5362,N_5265);
nand U5450 (N_5450,N_5389,N_5304);
xor U5451 (N_5451,N_5387,N_5313);
nor U5452 (N_5452,N_5251,N_5398);
and U5453 (N_5453,N_5358,N_5390);
and U5454 (N_5454,N_5328,N_5248);
or U5455 (N_5455,N_5299,N_5216);
nand U5456 (N_5456,N_5352,N_5348);
or U5457 (N_5457,N_5275,N_5225);
or U5458 (N_5458,N_5296,N_5315);
nor U5459 (N_5459,N_5391,N_5272);
and U5460 (N_5460,N_5366,N_5335);
nor U5461 (N_5461,N_5242,N_5288);
nor U5462 (N_5462,N_5220,N_5213);
nor U5463 (N_5463,N_5361,N_5273);
xor U5464 (N_5464,N_5307,N_5223);
nand U5465 (N_5465,N_5279,N_5202);
or U5466 (N_5466,N_5356,N_5373);
nand U5467 (N_5467,N_5285,N_5370);
or U5468 (N_5468,N_5212,N_5332);
and U5469 (N_5469,N_5230,N_5308);
xor U5470 (N_5470,N_5282,N_5311);
or U5471 (N_5471,N_5372,N_5240);
nor U5472 (N_5472,N_5342,N_5267);
or U5473 (N_5473,N_5305,N_5385);
xor U5474 (N_5474,N_5245,N_5274);
nor U5475 (N_5475,N_5327,N_5326);
xnor U5476 (N_5476,N_5243,N_5269);
and U5477 (N_5477,N_5383,N_5291);
and U5478 (N_5478,N_5363,N_5277);
xnor U5479 (N_5479,N_5331,N_5218);
nor U5480 (N_5480,N_5355,N_5247);
and U5481 (N_5481,N_5320,N_5295);
or U5482 (N_5482,N_5339,N_5347);
nand U5483 (N_5483,N_5392,N_5224);
xnor U5484 (N_5484,N_5378,N_5351);
and U5485 (N_5485,N_5376,N_5209);
xnor U5486 (N_5486,N_5324,N_5386);
nand U5487 (N_5487,N_5322,N_5246);
or U5488 (N_5488,N_5338,N_5374);
or U5489 (N_5489,N_5337,N_5284);
nand U5490 (N_5490,N_5334,N_5250);
nor U5491 (N_5491,N_5371,N_5380);
nor U5492 (N_5492,N_5219,N_5280);
nand U5493 (N_5493,N_5297,N_5329);
nor U5494 (N_5494,N_5239,N_5204);
and U5495 (N_5495,N_5217,N_5208);
nor U5496 (N_5496,N_5235,N_5228);
nand U5497 (N_5497,N_5286,N_5301);
nor U5498 (N_5498,N_5318,N_5289);
nor U5499 (N_5499,N_5290,N_5203);
and U5500 (N_5500,N_5287,N_5325);
and U5501 (N_5501,N_5381,N_5316);
and U5502 (N_5502,N_5285,N_5227);
nand U5503 (N_5503,N_5305,N_5220);
or U5504 (N_5504,N_5286,N_5249);
nand U5505 (N_5505,N_5348,N_5345);
nor U5506 (N_5506,N_5242,N_5325);
or U5507 (N_5507,N_5251,N_5357);
nand U5508 (N_5508,N_5300,N_5318);
nor U5509 (N_5509,N_5277,N_5318);
nand U5510 (N_5510,N_5269,N_5234);
nor U5511 (N_5511,N_5399,N_5345);
or U5512 (N_5512,N_5212,N_5313);
nand U5513 (N_5513,N_5306,N_5248);
nand U5514 (N_5514,N_5245,N_5267);
nor U5515 (N_5515,N_5206,N_5264);
or U5516 (N_5516,N_5352,N_5217);
and U5517 (N_5517,N_5260,N_5340);
nand U5518 (N_5518,N_5251,N_5379);
or U5519 (N_5519,N_5332,N_5336);
and U5520 (N_5520,N_5392,N_5308);
and U5521 (N_5521,N_5398,N_5307);
xnor U5522 (N_5522,N_5266,N_5232);
nor U5523 (N_5523,N_5385,N_5346);
or U5524 (N_5524,N_5212,N_5323);
xor U5525 (N_5525,N_5254,N_5295);
and U5526 (N_5526,N_5367,N_5310);
nor U5527 (N_5527,N_5316,N_5323);
nand U5528 (N_5528,N_5315,N_5314);
nand U5529 (N_5529,N_5393,N_5298);
and U5530 (N_5530,N_5352,N_5376);
or U5531 (N_5531,N_5358,N_5247);
nand U5532 (N_5532,N_5382,N_5351);
and U5533 (N_5533,N_5336,N_5385);
nor U5534 (N_5534,N_5388,N_5313);
and U5535 (N_5535,N_5239,N_5368);
nor U5536 (N_5536,N_5278,N_5220);
nand U5537 (N_5537,N_5383,N_5257);
xnor U5538 (N_5538,N_5311,N_5370);
xor U5539 (N_5539,N_5384,N_5214);
xnor U5540 (N_5540,N_5280,N_5249);
and U5541 (N_5541,N_5331,N_5355);
and U5542 (N_5542,N_5263,N_5391);
and U5543 (N_5543,N_5227,N_5224);
nor U5544 (N_5544,N_5320,N_5359);
nand U5545 (N_5545,N_5369,N_5302);
nand U5546 (N_5546,N_5217,N_5273);
nor U5547 (N_5547,N_5228,N_5206);
nand U5548 (N_5548,N_5237,N_5394);
xnor U5549 (N_5549,N_5291,N_5278);
nor U5550 (N_5550,N_5250,N_5248);
or U5551 (N_5551,N_5320,N_5395);
xor U5552 (N_5552,N_5367,N_5357);
and U5553 (N_5553,N_5244,N_5307);
and U5554 (N_5554,N_5397,N_5241);
nand U5555 (N_5555,N_5283,N_5316);
xor U5556 (N_5556,N_5364,N_5248);
and U5557 (N_5557,N_5367,N_5312);
xnor U5558 (N_5558,N_5365,N_5325);
nor U5559 (N_5559,N_5262,N_5236);
xor U5560 (N_5560,N_5250,N_5246);
nor U5561 (N_5561,N_5333,N_5391);
or U5562 (N_5562,N_5261,N_5277);
nor U5563 (N_5563,N_5373,N_5300);
nor U5564 (N_5564,N_5355,N_5382);
nand U5565 (N_5565,N_5221,N_5373);
or U5566 (N_5566,N_5243,N_5290);
nor U5567 (N_5567,N_5372,N_5371);
or U5568 (N_5568,N_5309,N_5224);
nor U5569 (N_5569,N_5309,N_5230);
nand U5570 (N_5570,N_5221,N_5313);
and U5571 (N_5571,N_5294,N_5295);
and U5572 (N_5572,N_5287,N_5254);
nand U5573 (N_5573,N_5245,N_5248);
nand U5574 (N_5574,N_5298,N_5208);
or U5575 (N_5575,N_5304,N_5263);
xnor U5576 (N_5576,N_5389,N_5318);
xnor U5577 (N_5577,N_5393,N_5232);
nor U5578 (N_5578,N_5332,N_5291);
xor U5579 (N_5579,N_5268,N_5303);
or U5580 (N_5580,N_5355,N_5272);
xor U5581 (N_5581,N_5325,N_5217);
or U5582 (N_5582,N_5319,N_5324);
and U5583 (N_5583,N_5331,N_5377);
nor U5584 (N_5584,N_5396,N_5373);
nor U5585 (N_5585,N_5263,N_5202);
or U5586 (N_5586,N_5219,N_5331);
nand U5587 (N_5587,N_5396,N_5253);
nor U5588 (N_5588,N_5373,N_5292);
and U5589 (N_5589,N_5254,N_5354);
or U5590 (N_5590,N_5236,N_5268);
or U5591 (N_5591,N_5371,N_5310);
or U5592 (N_5592,N_5318,N_5325);
xor U5593 (N_5593,N_5272,N_5315);
xnor U5594 (N_5594,N_5271,N_5350);
and U5595 (N_5595,N_5226,N_5202);
or U5596 (N_5596,N_5235,N_5276);
nor U5597 (N_5597,N_5249,N_5338);
nor U5598 (N_5598,N_5342,N_5299);
nor U5599 (N_5599,N_5243,N_5384);
or U5600 (N_5600,N_5433,N_5575);
or U5601 (N_5601,N_5512,N_5565);
nand U5602 (N_5602,N_5448,N_5437);
nor U5603 (N_5603,N_5450,N_5486);
xor U5604 (N_5604,N_5556,N_5535);
or U5605 (N_5605,N_5434,N_5459);
nand U5606 (N_5606,N_5441,N_5520);
or U5607 (N_5607,N_5586,N_5558);
nand U5608 (N_5608,N_5514,N_5477);
nor U5609 (N_5609,N_5596,N_5528);
or U5610 (N_5610,N_5576,N_5403);
or U5611 (N_5611,N_5569,N_5530);
nor U5612 (N_5612,N_5513,N_5585);
xnor U5613 (N_5613,N_5534,N_5428);
nand U5614 (N_5614,N_5494,N_5589);
or U5615 (N_5615,N_5549,N_5551);
xnor U5616 (N_5616,N_5418,N_5489);
and U5617 (N_5617,N_5577,N_5402);
and U5618 (N_5618,N_5544,N_5538);
nor U5619 (N_5619,N_5469,N_5451);
xor U5620 (N_5620,N_5405,N_5499);
nor U5621 (N_5621,N_5473,N_5568);
xor U5622 (N_5622,N_5471,N_5597);
and U5623 (N_5623,N_5560,N_5567);
nor U5624 (N_5624,N_5498,N_5500);
nor U5625 (N_5625,N_5529,N_5474);
or U5626 (N_5626,N_5415,N_5493);
or U5627 (N_5627,N_5476,N_5484);
or U5628 (N_5628,N_5542,N_5546);
or U5629 (N_5629,N_5412,N_5482);
nand U5630 (N_5630,N_5419,N_5465);
nand U5631 (N_5631,N_5539,N_5436);
xnor U5632 (N_5632,N_5458,N_5481);
or U5633 (N_5633,N_5416,N_5464);
or U5634 (N_5634,N_5442,N_5492);
and U5635 (N_5635,N_5507,N_5570);
nand U5636 (N_5636,N_5488,N_5590);
nor U5637 (N_5637,N_5468,N_5566);
nand U5638 (N_5638,N_5525,N_5409);
nand U5639 (N_5639,N_5447,N_5445);
or U5640 (N_5640,N_5593,N_5502);
and U5641 (N_5641,N_5564,N_5592);
xnor U5642 (N_5642,N_5478,N_5540);
nand U5643 (N_5643,N_5490,N_5421);
nor U5644 (N_5644,N_5543,N_5518);
and U5645 (N_5645,N_5424,N_5410);
xor U5646 (N_5646,N_5532,N_5531);
xnor U5647 (N_5647,N_5425,N_5523);
nand U5648 (N_5648,N_5579,N_5594);
and U5649 (N_5649,N_5583,N_5557);
xnor U5650 (N_5650,N_5479,N_5444);
nand U5651 (N_5651,N_5470,N_5559);
nand U5652 (N_5652,N_5536,N_5460);
or U5653 (N_5653,N_5461,N_5504);
and U5654 (N_5654,N_5547,N_5526);
xnor U5655 (N_5655,N_5524,N_5561);
xnor U5656 (N_5656,N_5483,N_5407);
xor U5657 (N_5657,N_5519,N_5496);
xor U5658 (N_5658,N_5487,N_5521);
and U5659 (N_5659,N_5573,N_5527);
or U5660 (N_5660,N_5462,N_5509);
xor U5661 (N_5661,N_5422,N_5515);
and U5662 (N_5662,N_5495,N_5554);
or U5663 (N_5663,N_5435,N_5472);
and U5664 (N_5664,N_5430,N_5591);
nor U5665 (N_5665,N_5432,N_5506);
and U5666 (N_5666,N_5584,N_5588);
nand U5667 (N_5667,N_5427,N_5467);
nor U5668 (N_5668,N_5401,N_5562);
nand U5669 (N_5669,N_5548,N_5503);
xor U5670 (N_5670,N_5406,N_5533);
nor U5671 (N_5671,N_5413,N_5454);
xor U5672 (N_5672,N_5456,N_5537);
nand U5673 (N_5673,N_5563,N_5455);
or U5674 (N_5674,N_5587,N_5517);
or U5675 (N_5675,N_5582,N_5463);
or U5676 (N_5676,N_5580,N_5599);
xnor U5677 (N_5677,N_5446,N_5457);
or U5678 (N_5678,N_5511,N_5510);
xor U5679 (N_5679,N_5466,N_5501);
and U5680 (N_5680,N_5595,N_5443);
or U5681 (N_5681,N_5508,N_5552);
and U5682 (N_5682,N_5440,N_5426);
or U5683 (N_5683,N_5545,N_5404);
or U5684 (N_5684,N_5550,N_5572);
nor U5685 (N_5685,N_5429,N_5491);
nand U5686 (N_5686,N_5497,N_5581);
xor U5687 (N_5687,N_5516,N_5480);
and U5688 (N_5688,N_5485,N_5475);
and U5689 (N_5689,N_5555,N_5571);
nand U5690 (N_5690,N_5449,N_5452);
xor U5691 (N_5691,N_5505,N_5453);
or U5692 (N_5692,N_5578,N_5431);
xor U5693 (N_5693,N_5411,N_5417);
or U5694 (N_5694,N_5400,N_5598);
and U5695 (N_5695,N_5423,N_5522);
and U5696 (N_5696,N_5420,N_5408);
nand U5697 (N_5697,N_5553,N_5574);
xnor U5698 (N_5698,N_5414,N_5439);
nand U5699 (N_5699,N_5438,N_5541);
or U5700 (N_5700,N_5537,N_5515);
or U5701 (N_5701,N_5476,N_5414);
nor U5702 (N_5702,N_5512,N_5507);
xor U5703 (N_5703,N_5591,N_5403);
and U5704 (N_5704,N_5443,N_5402);
xnor U5705 (N_5705,N_5540,N_5502);
nor U5706 (N_5706,N_5433,N_5576);
xnor U5707 (N_5707,N_5585,N_5422);
nand U5708 (N_5708,N_5543,N_5508);
xor U5709 (N_5709,N_5474,N_5572);
nor U5710 (N_5710,N_5456,N_5528);
or U5711 (N_5711,N_5568,N_5583);
and U5712 (N_5712,N_5487,N_5426);
nor U5713 (N_5713,N_5543,N_5593);
or U5714 (N_5714,N_5420,N_5471);
nor U5715 (N_5715,N_5478,N_5419);
and U5716 (N_5716,N_5546,N_5534);
nor U5717 (N_5717,N_5576,N_5578);
nand U5718 (N_5718,N_5482,N_5417);
and U5719 (N_5719,N_5455,N_5460);
or U5720 (N_5720,N_5521,N_5528);
or U5721 (N_5721,N_5427,N_5449);
nand U5722 (N_5722,N_5542,N_5437);
nand U5723 (N_5723,N_5505,N_5462);
or U5724 (N_5724,N_5560,N_5475);
and U5725 (N_5725,N_5538,N_5551);
xor U5726 (N_5726,N_5489,N_5576);
nand U5727 (N_5727,N_5559,N_5520);
and U5728 (N_5728,N_5438,N_5407);
xnor U5729 (N_5729,N_5596,N_5549);
nor U5730 (N_5730,N_5582,N_5507);
xor U5731 (N_5731,N_5457,N_5422);
and U5732 (N_5732,N_5527,N_5406);
xor U5733 (N_5733,N_5405,N_5418);
xnor U5734 (N_5734,N_5490,N_5496);
or U5735 (N_5735,N_5453,N_5451);
or U5736 (N_5736,N_5495,N_5541);
nand U5737 (N_5737,N_5413,N_5540);
nor U5738 (N_5738,N_5412,N_5490);
nor U5739 (N_5739,N_5591,N_5459);
nand U5740 (N_5740,N_5579,N_5563);
and U5741 (N_5741,N_5512,N_5443);
xor U5742 (N_5742,N_5551,N_5413);
xnor U5743 (N_5743,N_5459,N_5525);
nand U5744 (N_5744,N_5422,N_5468);
nand U5745 (N_5745,N_5583,N_5425);
nand U5746 (N_5746,N_5575,N_5410);
nor U5747 (N_5747,N_5433,N_5473);
xor U5748 (N_5748,N_5537,N_5455);
or U5749 (N_5749,N_5484,N_5594);
nor U5750 (N_5750,N_5574,N_5443);
nor U5751 (N_5751,N_5400,N_5589);
nand U5752 (N_5752,N_5598,N_5506);
nand U5753 (N_5753,N_5519,N_5523);
or U5754 (N_5754,N_5453,N_5599);
nand U5755 (N_5755,N_5504,N_5485);
xnor U5756 (N_5756,N_5444,N_5402);
xor U5757 (N_5757,N_5414,N_5483);
xnor U5758 (N_5758,N_5450,N_5554);
xor U5759 (N_5759,N_5536,N_5515);
xnor U5760 (N_5760,N_5468,N_5477);
nand U5761 (N_5761,N_5549,N_5585);
and U5762 (N_5762,N_5488,N_5553);
or U5763 (N_5763,N_5411,N_5468);
and U5764 (N_5764,N_5478,N_5504);
and U5765 (N_5765,N_5486,N_5551);
nand U5766 (N_5766,N_5440,N_5483);
nand U5767 (N_5767,N_5582,N_5484);
nor U5768 (N_5768,N_5513,N_5418);
nor U5769 (N_5769,N_5596,N_5529);
nor U5770 (N_5770,N_5445,N_5585);
nand U5771 (N_5771,N_5463,N_5514);
and U5772 (N_5772,N_5587,N_5403);
and U5773 (N_5773,N_5557,N_5475);
nand U5774 (N_5774,N_5528,N_5565);
nor U5775 (N_5775,N_5597,N_5523);
nor U5776 (N_5776,N_5554,N_5598);
or U5777 (N_5777,N_5510,N_5400);
nand U5778 (N_5778,N_5476,N_5544);
nand U5779 (N_5779,N_5583,N_5581);
nor U5780 (N_5780,N_5598,N_5433);
nor U5781 (N_5781,N_5559,N_5586);
xor U5782 (N_5782,N_5497,N_5478);
and U5783 (N_5783,N_5502,N_5568);
nand U5784 (N_5784,N_5459,N_5503);
and U5785 (N_5785,N_5456,N_5482);
or U5786 (N_5786,N_5594,N_5493);
or U5787 (N_5787,N_5463,N_5500);
or U5788 (N_5788,N_5528,N_5552);
and U5789 (N_5789,N_5445,N_5579);
or U5790 (N_5790,N_5522,N_5470);
xor U5791 (N_5791,N_5592,N_5448);
nor U5792 (N_5792,N_5595,N_5554);
and U5793 (N_5793,N_5465,N_5456);
nand U5794 (N_5794,N_5514,N_5425);
xor U5795 (N_5795,N_5493,N_5543);
nand U5796 (N_5796,N_5443,N_5529);
nand U5797 (N_5797,N_5551,N_5474);
or U5798 (N_5798,N_5512,N_5524);
nor U5799 (N_5799,N_5468,N_5580);
or U5800 (N_5800,N_5781,N_5632);
or U5801 (N_5801,N_5699,N_5751);
nor U5802 (N_5802,N_5714,N_5766);
xor U5803 (N_5803,N_5637,N_5609);
and U5804 (N_5804,N_5791,N_5729);
nand U5805 (N_5805,N_5737,N_5630);
nor U5806 (N_5806,N_5635,N_5704);
nor U5807 (N_5807,N_5677,N_5755);
nor U5808 (N_5808,N_5733,N_5671);
nand U5809 (N_5809,N_5720,N_5735);
xnor U5810 (N_5810,N_5627,N_5612);
nor U5811 (N_5811,N_5744,N_5644);
nor U5812 (N_5812,N_5719,N_5701);
and U5813 (N_5813,N_5797,N_5680);
and U5814 (N_5814,N_5689,N_5741);
nand U5815 (N_5815,N_5652,N_5688);
or U5816 (N_5816,N_5665,N_5787);
xor U5817 (N_5817,N_5707,N_5711);
nor U5818 (N_5818,N_5758,N_5667);
xnor U5819 (N_5819,N_5777,N_5731);
and U5820 (N_5820,N_5788,N_5657);
or U5821 (N_5821,N_5601,N_5618);
nand U5822 (N_5822,N_5673,N_5708);
nor U5823 (N_5823,N_5659,N_5684);
and U5824 (N_5824,N_5681,N_5736);
and U5825 (N_5825,N_5760,N_5710);
xnor U5826 (N_5826,N_5639,N_5728);
xnor U5827 (N_5827,N_5694,N_5732);
and U5828 (N_5828,N_5700,N_5675);
nand U5829 (N_5829,N_5795,N_5793);
xor U5830 (N_5830,N_5726,N_5672);
or U5831 (N_5831,N_5628,N_5798);
nor U5832 (N_5832,N_5669,N_5705);
and U5833 (N_5833,N_5661,N_5757);
nand U5834 (N_5834,N_5603,N_5676);
nand U5835 (N_5835,N_5698,N_5656);
xnor U5836 (N_5836,N_5647,N_5654);
nor U5837 (N_5837,N_5625,N_5645);
or U5838 (N_5838,N_5713,N_5768);
nand U5839 (N_5839,N_5770,N_5646);
or U5840 (N_5840,N_5649,N_5622);
nand U5841 (N_5841,N_5611,N_5607);
and U5842 (N_5842,N_5750,N_5734);
or U5843 (N_5843,N_5642,N_5775);
xor U5844 (N_5844,N_5624,N_5638);
xnor U5845 (N_5845,N_5739,N_5730);
xnor U5846 (N_5846,N_5776,N_5602);
nand U5847 (N_5847,N_5702,N_5746);
xor U5848 (N_5848,N_5748,N_5716);
nor U5849 (N_5849,N_5670,N_5685);
xnor U5850 (N_5850,N_5650,N_5610);
or U5851 (N_5851,N_5686,N_5636);
nand U5852 (N_5852,N_5789,N_5754);
and U5853 (N_5853,N_5633,N_5703);
nor U5854 (N_5854,N_5648,N_5658);
nor U5855 (N_5855,N_5763,N_5779);
nand U5856 (N_5856,N_5774,N_5738);
xnor U5857 (N_5857,N_5778,N_5690);
xor U5858 (N_5858,N_5621,N_5653);
nand U5859 (N_5859,N_5682,N_5743);
xor U5860 (N_5860,N_5740,N_5606);
nand U5861 (N_5861,N_5693,N_5727);
or U5862 (N_5862,N_5742,N_5799);
and U5863 (N_5863,N_5722,N_5668);
and U5864 (N_5864,N_5785,N_5674);
xnor U5865 (N_5865,N_5641,N_5772);
or U5866 (N_5866,N_5780,N_5767);
xnor U5867 (N_5867,N_5664,N_5629);
or U5868 (N_5868,N_5761,N_5769);
and U5869 (N_5869,N_5753,N_5745);
or U5870 (N_5870,N_5717,N_5796);
nand U5871 (N_5871,N_5617,N_5786);
nor U5872 (N_5872,N_5655,N_5794);
xnor U5873 (N_5873,N_5695,N_5718);
nand U5874 (N_5874,N_5762,N_5616);
xnor U5875 (N_5875,N_5683,N_5604);
xor U5876 (N_5876,N_5631,N_5660);
nor U5877 (N_5877,N_5614,N_5662);
nor U5878 (N_5878,N_5608,N_5697);
nor U5879 (N_5879,N_5623,N_5619);
nor U5880 (N_5880,N_5782,N_5634);
xor U5881 (N_5881,N_5725,N_5691);
nand U5882 (N_5882,N_5626,N_5721);
and U5883 (N_5883,N_5752,N_5692);
and U5884 (N_5884,N_5783,N_5709);
nand U5885 (N_5885,N_5792,N_5640);
nor U5886 (N_5886,N_5651,N_5723);
xnor U5887 (N_5887,N_5615,N_5620);
xnor U5888 (N_5888,N_5747,N_5663);
xor U5889 (N_5889,N_5764,N_5687);
and U5890 (N_5890,N_5724,N_5605);
nand U5891 (N_5891,N_5712,N_5759);
xor U5892 (N_5892,N_5715,N_5771);
nand U5893 (N_5893,N_5678,N_5765);
or U5894 (N_5894,N_5706,N_5613);
nand U5895 (N_5895,N_5679,N_5749);
or U5896 (N_5896,N_5666,N_5756);
nand U5897 (N_5897,N_5784,N_5773);
or U5898 (N_5898,N_5696,N_5790);
nand U5899 (N_5899,N_5600,N_5643);
and U5900 (N_5900,N_5773,N_5677);
nor U5901 (N_5901,N_5690,N_5700);
xor U5902 (N_5902,N_5778,N_5783);
xnor U5903 (N_5903,N_5688,N_5657);
and U5904 (N_5904,N_5763,N_5797);
nor U5905 (N_5905,N_5746,N_5771);
and U5906 (N_5906,N_5623,N_5628);
and U5907 (N_5907,N_5758,N_5688);
xor U5908 (N_5908,N_5660,N_5618);
nor U5909 (N_5909,N_5673,N_5663);
nand U5910 (N_5910,N_5758,N_5725);
nor U5911 (N_5911,N_5769,N_5754);
nand U5912 (N_5912,N_5756,N_5697);
and U5913 (N_5913,N_5733,N_5783);
nor U5914 (N_5914,N_5738,N_5686);
or U5915 (N_5915,N_5710,N_5638);
or U5916 (N_5916,N_5601,N_5680);
or U5917 (N_5917,N_5721,N_5613);
nand U5918 (N_5918,N_5773,N_5728);
and U5919 (N_5919,N_5668,N_5760);
and U5920 (N_5920,N_5639,N_5787);
nand U5921 (N_5921,N_5773,N_5721);
nand U5922 (N_5922,N_5689,N_5788);
nand U5923 (N_5923,N_5764,N_5698);
or U5924 (N_5924,N_5795,N_5724);
xor U5925 (N_5925,N_5682,N_5755);
xor U5926 (N_5926,N_5709,N_5643);
xor U5927 (N_5927,N_5635,N_5769);
nor U5928 (N_5928,N_5767,N_5750);
xor U5929 (N_5929,N_5676,N_5661);
nand U5930 (N_5930,N_5632,N_5778);
or U5931 (N_5931,N_5700,N_5751);
nor U5932 (N_5932,N_5624,N_5778);
and U5933 (N_5933,N_5722,N_5794);
nor U5934 (N_5934,N_5631,N_5690);
or U5935 (N_5935,N_5692,N_5628);
and U5936 (N_5936,N_5679,N_5705);
nand U5937 (N_5937,N_5759,N_5652);
xor U5938 (N_5938,N_5660,N_5708);
nand U5939 (N_5939,N_5641,N_5798);
nor U5940 (N_5940,N_5794,N_5702);
or U5941 (N_5941,N_5646,N_5656);
nand U5942 (N_5942,N_5708,N_5754);
nand U5943 (N_5943,N_5625,N_5769);
and U5944 (N_5944,N_5648,N_5727);
nand U5945 (N_5945,N_5746,N_5638);
or U5946 (N_5946,N_5695,N_5677);
or U5947 (N_5947,N_5734,N_5665);
and U5948 (N_5948,N_5727,N_5720);
nand U5949 (N_5949,N_5763,N_5717);
nor U5950 (N_5950,N_5698,N_5798);
nor U5951 (N_5951,N_5642,N_5742);
nor U5952 (N_5952,N_5604,N_5750);
nor U5953 (N_5953,N_5720,N_5634);
nor U5954 (N_5954,N_5782,N_5757);
or U5955 (N_5955,N_5793,N_5624);
xnor U5956 (N_5956,N_5605,N_5642);
or U5957 (N_5957,N_5765,N_5703);
xnor U5958 (N_5958,N_5797,N_5736);
nor U5959 (N_5959,N_5666,N_5696);
xnor U5960 (N_5960,N_5644,N_5652);
nand U5961 (N_5961,N_5752,N_5621);
nor U5962 (N_5962,N_5645,N_5704);
xnor U5963 (N_5963,N_5769,N_5621);
nor U5964 (N_5964,N_5662,N_5640);
or U5965 (N_5965,N_5726,N_5703);
and U5966 (N_5966,N_5637,N_5728);
or U5967 (N_5967,N_5720,N_5797);
and U5968 (N_5968,N_5765,N_5782);
and U5969 (N_5969,N_5712,N_5605);
nor U5970 (N_5970,N_5738,N_5760);
nor U5971 (N_5971,N_5664,N_5738);
and U5972 (N_5972,N_5765,N_5676);
or U5973 (N_5973,N_5627,N_5677);
nor U5974 (N_5974,N_5781,N_5642);
nor U5975 (N_5975,N_5796,N_5708);
nand U5976 (N_5976,N_5711,N_5726);
nor U5977 (N_5977,N_5755,N_5604);
and U5978 (N_5978,N_5635,N_5787);
or U5979 (N_5979,N_5770,N_5728);
or U5980 (N_5980,N_5640,N_5695);
or U5981 (N_5981,N_5662,N_5740);
or U5982 (N_5982,N_5681,N_5799);
or U5983 (N_5983,N_5623,N_5624);
nor U5984 (N_5984,N_5793,N_5666);
nand U5985 (N_5985,N_5670,N_5757);
xor U5986 (N_5986,N_5601,N_5663);
nor U5987 (N_5987,N_5677,N_5762);
and U5988 (N_5988,N_5783,N_5630);
nand U5989 (N_5989,N_5657,N_5749);
nand U5990 (N_5990,N_5700,N_5659);
xor U5991 (N_5991,N_5668,N_5721);
nand U5992 (N_5992,N_5639,N_5767);
nor U5993 (N_5993,N_5638,N_5690);
nor U5994 (N_5994,N_5672,N_5676);
xor U5995 (N_5995,N_5731,N_5665);
nand U5996 (N_5996,N_5670,N_5708);
and U5997 (N_5997,N_5638,N_5615);
xor U5998 (N_5998,N_5713,N_5634);
or U5999 (N_5999,N_5608,N_5672);
nand U6000 (N_6000,N_5828,N_5820);
nand U6001 (N_6001,N_5829,N_5940);
and U6002 (N_6002,N_5914,N_5892);
nor U6003 (N_6003,N_5856,N_5858);
xnor U6004 (N_6004,N_5975,N_5826);
xor U6005 (N_6005,N_5827,N_5813);
nor U6006 (N_6006,N_5874,N_5850);
and U6007 (N_6007,N_5852,N_5970);
or U6008 (N_6008,N_5928,N_5901);
and U6009 (N_6009,N_5851,N_5802);
xnor U6010 (N_6010,N_5944,N_5977);
nand U6011 (N_6011,N_5877,N_5889);
or U6012 (N_6012,N_5902,N_5898);
or U6013 (N_6013,N_5987,N_5869);
and U6014 (N_6014,N_5997,N_5876);
and U6015 (N_6015,N_5918,N_5803);
nor U6016 (N_6016,N_5818,N_5971);
nor U6017 (N_6017,N_5915,N_5969);
or U6018 (N_6018,N_5837,N_5814);
and U6019 (N_6019,N_5998,N_5991);
and U6020 (N_6020,N_5861,N_5855);
nor U6021 (N_6021,N_5805,N_5839);
or U6022 (N_6022,N_5830,N_5848);
and U6023 (N_6023,N_5994,N_5859);
and U6024 (N_6024,N_5883,N_5941);
nor U6025 (N_6025,N_5894,N_5926);
and U6026 (N_6026,N_5983,N_5907);
xnor U6027 (N_6027,N_5811,N_5833);
nand U6028 (N_6028,N_5943,N_5909);
xor U6029 (N_6029,N_5937,N_5873);
or U6030 (N_6030,N_5862,N_5920);
nand U6031 (N_6031,N_5825,N_5962);
or U6032 (N_6032,N_5871,N_5906);
or U6033 (N_6033,N_5984,N_5932);
or U6034 (N_6034,N_5959,N_5957);
xor U6035 (N_6035,N_5887,N_5881);
xor U6036 (N_6036,N_5817,N_5973);
or U6037 (N_6037,N_5886,N_5964);
and U6038 (N_6038,N_5953,N_5936);
nor U6039 (N_6039,N_5917,N_5834);
xnor U6040 (N_6040,N_5913,N_5801);
xnor U6041 (N_6041,N_5812,N_5843);
xor U6042 (N_6042,N_5992,N_5868);
nand U6043 (N_6043,N_5946,N_5939);
xor U6044 (N_6044,N_5822,N_5916);
or U6045 (N_6045,N_5963,N_5844);
or U6046 (N_6046,N_5934,N_5900);
or U6047 (N_6047,N_5947,N_5808);
or U6048 (N_6048,N_5863,N_5821);
nor U6049 (N_6049,N_5896,N_5846);
and U6050 (N_6050,N_5985,N_5841);
xnor U6051 (N_6051,N_5870,N_5847);
or U6052 (N_6052,N_5804,N_5905);
xor U6053 (N_6053,N_5938,N_5930);
nand U6054 (N_6054,N_5935,N_5875);
nor U6055 (N_6055,N_5961,N_5911);
nand U6056 (N_6056,N_5922,N_5952);
xor U6057 (N_6057,N_5815,N_5979);
xor U6058 (N_6058,N_5835,N_5949);
nand U6059 (N_6059,N_5978,N_5897);
and U6060 (N_6060,N_5838,N_5824);
xnor U6061 (N_6061,N_5981,N_5965);
nand U6062 (N_6062,N_5831,N_5972);
and U6063 (N_6063,N_5809,N_5888);
nand U6064 (N_6064,N_5921,N_5995);
or U6065 (N_6065,N_5903,N_5951);
xnor U6066 (N_6066,N_5878,N_5958);
nor U6067 (N_6067,N_5895,N_5904);
xor U6068 (N_6068,N_5842,N_5866);
and U6069 (N_6069,N_5857,N_5982);
and U6070 (N_6070,N_5908,N_5819);
xnor U6071 (N_6071,N_5806,N_5960);
nand U6072 (N_6072,N_5840,N_5955);
or U6073 (N_6073,N_5925,N_5910);
nor U6074 (N_6074,N_5853,N_5891);
nand U6075 (N_6075,N_5807,N_5849);
xnor U6076 (N_6076,N_5948,N_5999);
and U6077 (N_6077,N_5810,N_5854);
and U6078 (N_6078,N_5988,N_5990);
and U6079 (N_6079,N_5950,N_5899);
nand U6080 (N_6080,N_5980,N_5880);
xor U6081 (N_6081,N_5816,N_5885);
nand U6082 (N_6082,N_5989,N_5974);
and U6083 (N_6083,N_5929,N_5872);
or U6084 (N_6084,N_5890,N_5996);
nor U6085 (N_6085,N_5968,N_5945);
and U6086 (N_6086,N_5823,N_5976);
xnor U6087 (N_6087,N_5832,N_5923);
xnor U6088 (N_6088,N_5800,N_5860);
nand U6089 (N_6089,N_5986,N_5845);
nand U6090 (N_6090,N_5884,N_5993);
xnor U6091 (N_6091,N_5942,N_5933);
and U6092 (N_6092,N_5912,N_5931);
or U6093 (N_6093,N_5882,N_5864);
nand U6094 (N_6094,N_5879,N_5919);
or U6095 (N_6095,N_5956,N_5867);
or U6096 (N_6096,N_5836,N_5927);
and U6097 (N_6097,N_5966,N_5865);
nand U6098 (N_6098,N_5924,N_5954);
and U6099 (N_6099,N_5893,N_5967);
and U6100 (N_6100,N_5894,N_5911);
xor U6101 (N_6101,N_5810,N_5953);
nor U6102 (N_6102,N_5855,N_5999);
xnor U6103 (N_6103,N_5811,N_5831);
nand U6104 (N_6104,N_5809,N_5863);
and U6105 (N_6105,N_5842,N_5803);
nor U6106 (N_6106,N_5905,N_5887);
nor U6107 (N_6107,N_5938,N_5991);
nand U6108 (N_6108,N_5920,N_5978);
nand U6109 (N_6109,N_5985,N_5878);
nor U6110 (N_6110,N_5862,N_5844);
nor U6111 (N_6111,N_5977,N_5830);
xnor U6112 (N_6112,N_5908,N_5909);
nor U6113 (N_6113,N_5946,N_5883);
nand U6114 (N_6114,N_5969,N_5911);
nand U6115 (N_6115,N_5952,N_5944);
nand U6116 (N_6116,N_5864,N_5827);
nand U6117 (N_6117,N_5941,N_5837);
or U6118 (N_6118,N_5827,N_5921);
nand U6119 (N_6119,N_5952,N_5801);
xnor U6120 (N_6120,N_5858,N_5903);
xnor U6121 (N_6121,N_5831,N_5841);
nand U6122 (N_6122,N_5983,N_5913);
nand U6123 (N_6123,N_5953,N_5918);
nand U6124 (N_6124,N_5966,N_5857);
nor U6125 (N_6125,N_5838,N_5809);
and U6126 (N_6126,N_5949,N_5801);
and U6127 (N_6127,N_5852,N_5873);
xor U6128 (N_6128,N_5917,N_5989);
or U6129 (N_6129,N_5921,N_5874);
nand U6130 (N_6130,N_5973,N_5919);
xor U6131 (N_6131,N_5989,N_5843);
nor U6132 (N_6132,N_5900,N_5838);
and U6133 (N_6133,N_5835,N_5921);
nand U6134 (N_6134,N_5807,N_5830);
nand U6135 (N_6135,N_5896,N_5830);
xnor U6136 (N_6136,N_5855,N_5996);
xor U6137 (N_6137,N_5861,N_5978);
or U6138 (N_6138,N_5940,N_5963);
xor U6139 (N_6139,N_5809,N_5941);
nor U6140 (N_6140,N_5808,N_5890);
nor U6141 (N_6141,N_5858,N_5948);
nand U6142 (N_6142,N_5930,N_5840);
nand U6143 (N_6143,N_5827,N_5846);
or U6144 (N_6144,N_5957,N_5918);
and U6145 (N_6145,N_5882,N_5990);
or U6146 (N_6146,N_5886,N_5981);
or U6147 (N_6147,N_5820,N_5945);
nand U6148 (N_6148,N_5811,N_5931);
and U6149 (N_6149,N_5925,N_5879);
and U6150 (N_6150,N_5949,N_5994);
and U6151 (N_6151,N_5855,N_5816);
nand U6152 (N_6152,N_5961,N_5975);
xor U6153 (N_6153,N_5980,N_5888);
nor U6154 (N_6154,N_5896,N_5867);
nor U6155 (N_6155,N_5863,N_5939);
xnor U6156 (N_6156,N_5953,N_5896);
and U6157 (N_6157,N_5850,N_5964);
and U6158 (N_6158,N_5939,N_5882);
or U6159 (N_6159,N_5996,N_5844);
xnor U6160 (N_6160,N_5949,N_5957);
nand U6161 (N_6161,N_5954,N_5989);
xnor U6162 (N_6162,N_5941,N_5907);
nand U6163 (N_6163,N_5897,N_5998);
nor U6164 (N_6164,N_5964,N_5845);
or U6165 (N_6165,N_5955,N_5902);
nand U6166 (N_6166,N_5970,N_5803);
xor U6167 (N_6167,N_5803,N_5810);
and U6168 (N_6168,N_5809,N_5983);
and U6169 (N_6169,N_5886,N_5824);
and U6170 (N_6170,N_5868,N_5840);
nor U6171 (N_6171,N_5805,N_5949);
xnor U6172 (N_6172,N_5859,N_5815);
and U6173 (N_6173,N_5809,N_5954);
nor U6174 (N_6174,N_5816,N_5910);
nand U6175 (N_6175,N_5805,N_5845);
and U6176 (N_6176,N_5891,N_5994);
nand U6177 (N_6177,N_5931,N_5958);
xor U6178 (N_6178,N_5843,N_5879);
or U6179 (N_6179,N_5865,N_5847);
nand U6180 (N_6180,N_5923,N_5834);
nand U6181 (N_6181,N_5991,N_5870);
and U6182 (N_6182,N_5970,N_5994);
xor U6183 (N_6183,N_5862,N_5892);
nand U6184 (N_6184,N_5811,N_5825);
and U6185 (N_6185,N_5874,N_5986);
nand U6186 (N_6186,N_5852,N_5910);
and U6187 (N_6187,N_5879,N_5946);
or U6188 (N_6188,N_5847,N_5896);
nor U6189 (N_6189,N_5973,N_5805);
nand U6190 (N_6190,N_5864,N_5922);
or U6191 (N_6191,N_5949,N_5862);
nand U6192 (N_6192,N_5933,N_5988);
xnor U6193 (N_6193,N_5880,N_5865);
nor U6194 (N_6194,N_5825,N_5849);
and U6195 (N_6195,N_5883,N_5866);
or U6196 (N_6196,N_5885,N_5872);
nor U6197 (N_6197,N_5990,N_5932);
or U6198 (N_6198,N_5835,N_5940);
and U6199 (N_6199,N_5805,N_5972);
nor U6200 (N_6200,N_6086,N_6158);
xnor U6201 (N_6201,N_6122,N_6106);
or U6202 (N_6202,N_6019,N_6075);
nand U6203 (N_6203,N_6185,N_6038);
and U6204 (N_6204,N_6176,N_6050);
and U6205 (N_6205,N_6067,N_6167);
nand U6206 (N_6206,N_6011,N_6026);
and U6207 (N_6207,N_6195,N_6047);
xor U6208 (N_6208,N_6058,N_6141);
xnor U6209 (N_6209,N_6193,N_6048);
nor U6210 (N_6210,N_6032,N_6118);
nor U6211 (N_6211,N_6124,N_6137);
xor U6212 (N_6212,N_6155,N_6018);
nor U6213 (N_6213,N_6049,N_6175);
xnor U6214 (N_6214,N_6017,N_6072);
or U6215 (N_6215,N_6186,N_6044);
and U6216 (N_6216,N_6103,N_6190);
and U6217 (N_6217,N_6116,N_6153);
xor U6218 (N_6218,N_6096,N_6088);
nand U6219 (N_6219,N_6097,N_6029);
and U6220 (N_6220,N_6008,N_6154);
xnor U6221 (N_6221,N_6066,N_6062);
or U6222 (N_6222,N_6108,N_6131);
or U6223 (N_6223,N_6087,N_6101);
nor U6224 (N_6224,N_6027,N_6129);
xnor U6225 (N_6225,N_6037,N_6083);
xnor U6226 (N_6226,N_6005,N_6120);
or U6227 (N_6227,N_6021,N_6149);
or U6228 (N_6228,N_6169,N_6188);
nand U6229 (N_6229,N_6171,N_6166);
and U6230 (N_6230,N_6045,N_6168);
and U6231 (N_6231,N_6043,N_6076);
nor U6232 (N_6232,N_6016,N_6023);
nand U6233 (N_6233,N_6015,N_6064);
nand U6234 (N_6234,N_6165,N_6100);
xnor U6235 (N_6235,N_6150,N_6152);
xor U6236 (N_6236,N_6157,N_6151);
xnor U6237 (N_6237,N_6055,N_6111);
and U6238 (N_6238,N_6069,N_6028);
or U6239 (N_6239,N_6107,N_6183);
xor U6240 (N_6240,N_6014,N_6148);
and U6241 (N_6241,N_6004,N_6054);
and U6242 (N_6242,N_6121,N_6179);
xnor U6243 (N_6243,N_6059,N_6102);
or U6244 (N_6244,N_6196,N_6147);
xnor U6245 (N_6245,N_6033,N_6079);
nor U6246 (N_6246,N_6132,N_6099);
xnor U6247 (N_6247,N_6110,N_6061);
or U6248 (N_6248,N_6022,N_6002);
nand U6249 (N_6249,N_6174,N_6143);
or U6250 (N_6250,N_6128,N_6010);
nor U6251 (N_6251,N_6080,N_6136);
or U6252 (N_6252,N_6056,N_6113);
nand U6253 (N_6253,N_6041,N_6142);
nor U6254 (N_6254,N_6051,N_6156);
xnor U6255 (N_6255,N_6130,N_6053);
nor U6256 (N_6256,N_6199,N_6123);
or U6257 (N_6257,N_6074,N_6036);
or U6258 (N_6258,N_6163,N_6119);
xnor U6259 (N_6259,N_6082,N_6104);
or U6260 (N_6260,N_6081,N_6138);
nor U6261 (N_6261,N_6125,N_6194);
or U6262 (N_6262,N_6115,N_6173);
nor U6263 (N_6263,N_6091,N_6063);
and U6264 (N_6264,N_6109,N_6024);
nor U6265 (N_6265,N_6057,N_6065);
nand U6266 (N_6266,N_6006,N_6139);
xor U6267 (N_6267,N_6007,N_6042);
nand U6268 (N_6268,N_6077,N_6133);
nand U6269 (N_6269,N_6025,N_6012);
nor U6270 (N_6270,N_6040,N_6162);
nor U6271 (N_6271,N_6034,N_6177);
nand U6272 (N_6272,N_6192,N_6180);
nor U6273 (N_6273,N_6178,N_6126);
and U6274 (N_6274,N_6117,N_6198);
xor U6275 (N_6275,N_6003,N_6046);
or U6276 (N_6276,N_6145,N_6084);
or U6277 (N_6277,N_6070,N_6078);
and U6278 (N_6278,N_6146,N_6094);
nor U6279 (N_6279,N_6085,N_6060);
xor U6280 (N_6280,N_6090,N_6140);
nand U6281 (N_6281,N_6170,N_6127);
xnor U6282 (N_6282,N_6052,N_6089);
nor U6283 (N_6283,N_6181,N_6035);
or U6284 (N_6284,N_6000,N_6039);
or U6285 (N_6285,N_6095,N_6182);
nand U6286 (N_6286,N_6114,N_6189);
nor U6287 (N_6287,N_6073,N_6093);
nand U6288 (N_6288,N_6071,N_6197);
or U6289 (N_6289,N_6161,N_6159);
or U6290 (N_6290,N_6001,N_6009);
xor U6291 (N_6291,N_6030,N_6144);
nor U6292 (N_6292,N_6020,N_6164);
xor U6293 (N_6293,N_6191,N_6134);
nor U6294 (N_6294,N_6172,N_6135);
nand U6295 (N_6295,N_6187,N_6068);
and U6296 (N_6296,N_6112,N_6031);
nor U6297 (N_6297,N_6184,N_6092);
or U6298 (N_6298,N_6013,N_6105);
xnor U6299 (N_6299,N_6098,N_6160);
and U6300 (N_6300,N_6147,N_6169);
xnor U6301 (N_6301,N_6076,N_6000);
nor U6302 (N_6302,N_6112,N_6156);
nor U6303 (N_6303,N_6027,N_6102);
nand U6304 (N_6304,N_6007,N_6117);
and U6305 (N_6305,N_6059,N_6127);
or U6306 (N_6306,N_6119,N_6098);
nor U6307 (N_6307,N_6059,N_6105);
nor U6308 (N_6308,N_6150,N_6015);
and U6309 (N_6309,N_6115,N_6006);
nor U6310 (N_6310,N_6172,N_6006);
nand U6311 (N_6311,N_6106,N_6164);
xor U6312 (N_6312,N_6064,N_6085);
and U6313 (N_6313,N_6194,N_6064);
or U6314 (N_6314,N_6173,N_6090);
and U6315 (N_6315,N_6155,N_6163);
or U6316 (N_6316,N_6135,N_6137);
and U6317 (N_6317,N_6092,N_6189);
and U6318 (N_6318,N_6141,N_6047);
nor U6319 (N_6319,N_6054,N_6140);
or U6320 (N_6320,N_6163,N_6117);
nor U6321 (N_6321,N_6198,N_6181);
nand U6322 (N_6322,N_6166,N_6120);
nand U6323 (N_6323,N_6059,N_6182);
xor U6324 (N_6324,N_6171,N_6194);
or U6325 (N_6325,N_6049,N_6020);
nor U6326 (N_6326,N_6180,N_6076);
and U6327 (N_6327,N_6199,N_6186);
and U6328 (N_6328,N_6114,N_6148);
nor U6329 (N_6329,N_6098,N_6122);
nand U6330 (N_6330,N_6028,N_6119);
nand U6331 (N_6331,N_6143,N_6081);
xnor U6332 (N_6332,N_6010,N_6155);
xor U6333 (N_6333,N_6110,N_6044);
nand U6334 (N_6334,N_6014,N_6100);
or U6335 (N_6335,N_6184,N_6198);
nor U6336 (N_6336,N_6138,N_6128);
xnor U6337 (N_6337,N_6167,N_6139);
xnor U6338 (N_6338,N_6001,N_6184);
nor U6339 (N_6339,N_6144,N_6160);
xor U6340 (N_6340,N_6068,N_6099);
and U6341 (N_6341,N_6098,N_6020);
nand U6342 (N_6342,N_6099,N_6186);
nand U6343 (N_6343,N_6021,N_6097);
nor U6344 (N_6344,N_6172,N_6119);
or U6345 (N_6345,N_6183,N_6109);
nor U6346 (N_6346,N_6148,N_6112);
or U6347 (N_6347,N_6166,N_6086);
nor U6348 (N_6348,N_6144,N_6099);
and U6349 (N_6349,N_6172,N_6116);
xor U6350 (N_6350,N_6195,N_6059);
xor U6351 (N_6351,N_6191,N_6166);
and U6352 (N_6352,N_6038,N_6042);
nor U6353 (N_6353,N_6075,N_6066);
nand U6354 (N_6354,N_6163,N_6128);
or U6355 (N_6355,N_6180,N_6025);
nor U6356 (N_6356,N_6104,N_6168);
and U6357 (N_6357,N_6050,N_6185);
nand U6358 (N_6358,N_6032,N_6128);
or U6359 (N_6359,N_6038,N_6015);
and U6360 (N_6360,N_6136,N_6098);
and U6361 (N_6361,N_6116,N_6012);
xnor U6362 (N_6362,N_6108,N_6177);
nor U6363 (N_6363,N_6029,N_6066);
nor U6364 (N_6364,N_6039,N_6063);
nor U6365 (N_6365,N_6149,N_6078);
nor U6366 (N_6366,N_6180,N_6046);
nand U6367 (N_6367,N_6046,N_6116);
nor U6368 (N_6368,N_6081,N_6053);
or U6369 (N_6369,N_6123,N_6157);
or U6370 (N_6370,N_6037,N_6090);
xnor U6371 (N_6371,N_6060,N_6189);
or U6372 (N_6372,N_6151,N_6066);
or U6373 (N_6373,N_6142,N_6055);
nand U6374 (N_6374,N_6131,N_6151);
nor U6375 (N_6375,N_6093,N_6072);
nor U6376 (N_6376,N_6024,N_6104);
or U6377 (N_6377,N_6066,N_6188);
and U6378 (N_6378,N_6134,N_6146);
and U6379 (N_6379,N_6145,N_6103);
nor U6380 (N_6380,N_6047,N_6197);
and U6381 (N_6381,N_6156,N_6017);
nor U6382 (N_6382,N_6126,N_6088);
and U6383 (N_6383,N_6023,N_6045);
and U6384 (N_6384,N_6187,N_6128);
nor U6385 (N_6385,N_6123,N_6158);
and U6386 (N_6386,N_6193,N_6098);
or U6387 (N_6387,N_6191,N_6111);
or U6388 (N_6388,N_6056,N_6000);
or U6389 (N_6389,N_6175,N_6199);
nand U6390 (N_6390,N_6083,N_6005);
nand U6391 (N_6391,N_6084,N_6099);
or U6392 (N_6392,N_6162,N_6012);
and U6393 (N_6393,N_6080,N_6011);
nand U6394 (N_6394,N_6163,N_6003);
nor U6395 (N_6395,N_6132,N_6117);
nor U6396 (N_6396,N_6025,N_6103);
and U6397 (N_6397,N_6078,N_6175);
nand U6398 (N_6398,N_6042,N_6010);
and U6399 (N_6399,N_6034,N_6141);
and U6400 (N_6400,N_6341,N_6357);
xnor U6401 (N_6401,N_6278,N_6237);
xor U6402 (N_6402,N_6218,N_6249);
nor U6403 (N_6403,N_6380,N_6202);
nand U6404 (N_6404,N_6304,N_6206);
and U6405 (N_6405,N_6224,N_6391);
nor U6406 (N_6406,N_6399,N_6299);
nand U6407 (N_6407,N_6372,N_6332);
or U6408 (N_6408,N_6253,N_6389);
and U6409 (N_6409,N_6352,N_6247);
xnor U6410 (N_6410,N_6209,N_6238);
nor U6411 (N_6411,N_6322,N_6207);
xor U6412 (N_6412,N_6330,N_6312);
nand U6413 (N_6413,N_6364,N_6254);
nand U6414 (N_6414,N_6388,N_6211);
or U6415 (N_6415,N_6212,N_6297);
or U6416 (N_6416,N_6284,N_6397);
nor U6417 (N_6417,N_6227,N_6320);
or U6418 (N_6418,N_6273,N_6325);
xnor U6419 (N_6419,N_6329,N_6272);
nor U6420 (N_6420,N_6353,N_6373);
or U6421 (N_6421,N_6266,N_6231);
xnor U6422 (N_6422,N_6354,N_6303);
nor U6423 (N_6423,N_6281,N_6392);
and U6424 (N_6424,N_6292,N_6245);
nand U6425 (N_6425,N_6323,N_6293);
xor U6426 (N_6426,N_6208,N_6366);
xor U6427 (N_6427,N_6302,N_6220);
nor U6428 (N_6428,N_6393,N_6213);
nand U6429 (N_6429,N_6290,N_6351);
or U6430 (N_6430,N_6205,N_6315);
or U6431 (N_6431,N_6216,N_6342);
nand U6432 (N_6432,N_6276,N_6313);
or U6433 (N_6433,N_6210,N_6260);
or U6434 (N_6434,N_6390,N_6338);
nor U6435 (N_6435,N_6318,N_6244);
and U6436 (N_6436,N_6333,N_6381);
nand U6437 (N_6437,N_6301,N_6204);
nand U6438 (N_6438,N_6239,N_6285);
nor U6439 (N_6439,N_6246,N_6267);
or U6440 (N_6440,N_6217,N_6326);
or U6441 (N_6441,N_6233,N_6280);
nand U6442 (N_6442,N_6374,N_6359);
nor U6443 (N_6443,N_6386,N_6378);
nand U6444 (N_6444,N_6257,N_6251);
nand U6445 (N_6445,N_6243,N_6258);
and U6446 (N_6446,N_6230,N_6379);
nand U6447 (N_6447,N_6309,N_6314);
xnor U6448 (N_6448,N_6382,N_6226);
nand U6449 (N_6449,N_6316,N_6360);
and U6450 (N_6450,N_6346,N_6328);
nor U6451 (N_6451,N_6248,N_6308);
xor U6452 (N_6452,N_6228,N_6368);
nand U6453 (N_6453,N_6305,N_6236);
or U6454 (N_6454,N_6363,N_6298);
or U6455 (N_6455,N_6370,N_6365);
xnor U6456 (N_6456,N_6340,N_6358);
or U6457 (N_6457,N_6222,N_6279);
xnor U6458 (N_6458,N_6283,N_6288);
xor U6459 (N_6459,N_6262,N_6271);
and U6460 (N_6460,N_6289,N_6232);
and U6461 (N_6461,N_6234,N_6261);
xor U6462 (N_6462,N_6270,N_6317);
nand U6463 (N_6463,N_6296,N_6367);
or U6464 (N_6464,N_6349,N_6294);
or U6465 (N_6465,N_6275,N_6331);
nor U6466 (N_6466,N_6229,N_6356);
or U6467 (N_6467,N_6215,N_6252);
nand U6468 (N_6468,N_6387,N_6263);
or U6469 (N_6469,N_6348,N_6344);
xnor U6470 (N_6470,N_6256,N_6334);
xor U6471 (N_6471,N_6335,N_6203);
nand U6472 (N_6472,N_6306,N_6336);
or U6473 (N_6473,N_6282,N_6327);
xnor U6474 (N_6474,N_6310,N_6240);
or U6475 (N_6475,N_6311,N_6339);
and U6476 (N_6476,N_6307,N_6200);
nor U6477 (N_6477,N_6268,N_6345);
xnor U6478 (N_6478,N_6235,N_6324);
or U6479 (N_6479,N_6250,N_6242);
nand U6480 (N_6480,N_6376,N_6377);
or U6481 (N_6481,N_6264,N_6396);
or U6482 (N_6482,N_6277,N_6295);
and U6483 (N_6483,N_6369,N_6225);
and U6484 (N_6484,N_6343,N_6385);
xor U6485 (N_6485,N_6395,N_6286);
or U6486 (N_6486,N_6214,N_6347);
nor U6487 (N_6487,N_6287,N_6291);
nor U6488 (N_6488,N_6384,N_6265);
xnor U6489 (N_6489,N_6274,N_6221);
and U6490 (N_6490,N_6319,N_6241);
nand U6491 (N_6491,N_6269,N_6383);
nor U6492 (N_6492,N_6394,N_6361);
or U6493 (N_6493,N_6337,N_6398);
xor U6494 (N_6494,N_6201,N_6255);
and U6495 (N_6495,N_6350,N_6219);
or U6496 (N_6496,N_6362,N_6371);
and U6497 (N_6497,N_6355,N_6300);
and U6498 (N_6498,N_6223,N_6375);
xnor U6499 (N_6499,N_6321,N_6259);
and U6500 (N_6500,N_6310,N_6208);
and U6501 (N_6501,N_6322,N_6217);
or U6502 (N_6502,N_6342,N_6245);
nor U6503 (N_6503,N_6249,N_6295);
nand U6504 (N_6504,N_6348,N_6281);
xnor U6505 (N_6505,N_6262,N_6229);
and U6506 (N_6506,N_6334,N_6286);
nand U6507 (N_6507,N_6279,N_6232);
nand U6508 (N_6508,N_6285,N_6328);
and U6509 (N_6509,N_6316,N_6347);
xnor U6510 (N_6510,N_6368,N_6375);
and U6511 (N_6511,N_6397,N_6342);
xnor U6512 (N_6512,N_6333,N_6377);
xnor U6513 (N_6513,N_6330,N_6276);
or U6514 (N_6514,N_6397,N_6308);
nand U6515 (N_6515,N_6364,N_6286);
nor U6516 (N_6516,N_6289,N_6290);
nand U6517 (N_6517,N_6268,N_6360);
nand U6518 (N_6518,N_6287,N_6330);
or U6519 (N_6519,N_6353,N_6244);
nor U6520 (N_6520,N_6210,N_6259);
or U6521 (N_6521,N_6398,N_6213);
or U6522 (N_6522,N_6278,N_6289);
nand U6523 (N_6523,N_6231,N_6398);
nor U6524 (N_6524,N_6333,N_6369);
xor U6525 (N_6525,N_6373,N_6292);
and U6526 (N_6526,N_6316,N_6251);
xnor U6527 (N_6527,N_6311,N_6244);
xor U6528 (N_6528,N_6326,N_6267);
nand U6529 (N_6529,N_6226,N_6333);
xor U6530 (N_6530,N_6218,N_6256);
or U6531 (N_6531,N_6269,N_6244);
xnor U6532 (N_6532,N_6289,N_6262);
or U6533 (N_6533,N_6272,N_6303);
or U6534 (N_6534,N_6236,N_6251);
nand U6535 (N_6535,N_6358,N_6222);
nand U6536 (N_6536,N_6302,N_6280);
and U6537 (N_6537,N_6245,N_6335);
and U6538 (N_6538,N_6255,N_6366);
xnor U6539 (N_6539,N_6211,N_6366);
xor U6540 (N_6540,N_6258,N_6284);
and U6541 (N_6541,N_6386,N_6307);
xnor U6542 (N_6542,N_6270,N_6284);
or U6543 (N_6543,N_6390,N_6302);
nor U6544 (N_6544,N_6277,N_6238);
xnor U6545 (N_6545,N_6340,N_6376);
and U6546 (N_6546,N_6330,N_6292);
nor U6547 (N_6547,N_6377,N_6201);
nor U6548 (N_6548,N_6204,N_6323);
xnor U6549 (N_6549,N_6289,N_6231);
and U6550 (N_6550,N_6200,N_6398);
and U6551 (N_6551,N_6399,N_6266);
xor U6552 (N_6552,N_6393,N_6274);
nor U6553 (N_6553,N_6306,N_6329);
or U6554 (N_6554,N_6306,N_6271);
xor U6555 (N_6555,N_6344,N_6389);
xnor U6556 (N_6556,N_6379,N_6361);
nor U6557 (N_6557,N_6342,N_6383);
and U6558 (N_6558,N_6216,N_6297);
nand U6559 (N_6559,N_6238,N_6348);
or U6560 (N_6560,N_6224,N_6292);
or U6561 (N_6561,N_6214,N_6228);
nand U6562 (N_6562,N_6371,N_6223);
nand U6563 (N_6563,N_6345,N_6227);
nand U6564 (N_6564,N_6319,N_6377);
nor U6565 (N_6565,N_6284,N_6301);
xor U6566 (N_6566,N_6262,N_6329);
xnor U6567 (N_6567,N_6370,N_6264);
nand U6568 (N_6568,N_6386,N_6370);
xor U6569 (N_6569,N_6298,N_6267);
nand U6570 (N_6570,N_6275,N_6381);
xor U6571 (N_6571,N_6340,N_6317);
and U6572 (N_6572,N_6299,N_6226);
xnor U6573 (N_6573,N_6355,N_6224);
nand U6574 (N_6574,N_6243,N_6328);
and U6575 (N_6575,N_6324,N_6209);
xnor U6576 (N_6576,N_6202,N_6351);
xnor U6577 (N_6577,N_6341,N_6350);
xor U6578 (N_6578,N_6362,N_6310);
nor U6579 (N_6579,N_6273,N_6316);
nor U6580 (N_6580,N_6259,N_6221);
or U6581 (N_6581,N_6349,N_6266);
and U6582 (N_6582,N_6378,N_6213);
or U6583 (N_6583,N_6277,N_6287);
and U6584 (N_6584,N_6242,N_6361);
xnor U6585 (N_6585,N_6253,N_6334);
and U6586 (N_6586,N_6331,N_6320);
nand U6587 (N_6587,N_6343,N_6243);
xor U6588 (N_6588,N_6303,N_6234);
xor U6589 (N_6589,N_6288,N_6272);
nand U6590 (N_6590,N_6342,N_6301);
nand U6591 (N_6591,N_6257,N_6372);
nand U6592 (N_6592,N_6219,N_6204);
or U6593 (N_6593,N_6362,N_6204);
nor U6594 (N_6594,N_6365,N_6263);
or U6595 (N_6595,N_6201,N_6258);
and U6596 (N_6596,N_6356,N_6370);
or U6597 (N_6597,N_6306,N_6393);
xor U6598 (N_6598,N_6249,N_6213);
or U6599 (N_6599,N_6205,N_6289);
nor U6600 (N_6600,N_6522,N_6448);
nor U6601 (N_6601,N_6575,N_6492);
xnor U6602 (N_6602,N_6535,N_6419);
xnor U6603 (N_6603,N_6439,N_6502);
xnor U6604 (N_6604,N_6475,N_6468);
xnor U6605 (N_6605,N_6525,N_6423);
or U6606 (N_6606,N_6563,N_6433);
xor U6607 (N_6607,N_6408,N_6561);
nor U6608 (N_6608,N_6596,N_6467);
or U6609 (N_6609,N_6430,N_6539);
or U6610 (N_6610,N_6519,N_6400);
and U6611 (N_6611,N_6573,N_6486);
nand U6612 (N_6612,N_6487,N_6526);
nand U6613 (N_6613,N_6454,N_6506);
xnor U6614 (N_6614,N_6427,N_6477);
xor U6615 (N_6615,N_6436,N_6424);
nand U6616 (N_6616,N_6559,N_6459);
nand U6617 (N_6617,N_6498,N_6579);
nor U6618 (N_6618,N_6517,N_6518);
nand U6619 (N_6619,N_6586,N_6413);
and U6620 (N_6620,N_6549,N_6570);
nand U6621 (N_6621,N_6493,N_6496);
xnor U6622 (N_6622,N_6440,N_6551);
nand U6623 (N_6623,N_6417,N_6510);
or U6624 (N_6624,N_6509,N_6420);
nand U6625 (N_6625,N_6404,N_6581);
xor U6626 (N_6626,N_6598,N_6558);
or U6627 (N_6627,N_6554,N_6547);
or U6628 (N_6628,N_6520,N_6577);
nand U6629 (N_6629,N_6421,N_6504);
or U6630 (N_6630,N_6499,N_6473);
nor U6631 (N_6631,N_6412,N_6515);
nor U6632 (N_6632,N_6500,N_6451);
xor U6633 (N_6633,N_6476,N_6401);
or U6634 (N_6634,N_6550,N_6490);
nand U6635 (N_6635,N_6453,N_6511);
and U6636 (N_6636,N_6501,N_6574);
or U6637 (N_6637,N_6489,N_6458);
nor U6638 (N_6638,N_6564,N_6548);
nand U6639 (N_6639,N_6508,N_6464);
xnor U6640 (N_6640,N_6481,N_6407);
xnor U6641 (N_6641,N_6572,N_6562);
and U6642 (N_6642,N_6514,N_6542);
nand U6643 (N_6643,N_6484,N_6443);
and U6644 (N_6644,N_6463,N_6403);
nand U6645 (N_6645,N_6576,N_6491);
nor U6646 (N_6646,N_6482,N_6405);
xnor U6647 (N_6647,N_6485,N_6461);
nor U6648 (N_6648,N_6435,N_6494);
nand U6649 (N_6649,N_6507,N_6534);
xnor U6650 (N_6650,N_6588,N_6533);
or U6651 (N_6651,N_6418,N_6471);
or U6652 (N_6652,N_6523,N_6536);
or U6653 (N_6653,N_6411,N_6546);
xor U6654 (N_6654,N_6474,N_6597);
xnor U6655 (N_6655,N_6479,N_6531);
xnor U6656 (N_6656,N_6585,N_6414);
nand U6657 (N_6657,N_6529,N_6465);
nand U6658 (N_6658,N_6444,N_6513);
nand U6659 (N_6659,N_6478,N_6582);
or U6660 (N_6660,N_6472,N_6469);
nor U6661 (N_6661,N_6512,N_6446);
nor U6662 (N_6662,N_6503,N_6555);
nand U6663 (N_6663,N_6599,N_6445);
or U6664 (N_6664,N_6545,N_6488);
and U6665 (N_6665,N_6455,N_6524);
xor U6666 (N_6666,N_6566,N_6415);
nand U6667 (N_6667,N_6544,N_6416);
nand U6668 (N_6668,N_6587,N_6593);
or U6669 (N_6669,N_6456,N_6470);
nor U6670 (N_6670,N_6429,N_6567);
and U6671 (N_6671,N_6556,N_6437);
nor U6672 (N_6672,N_6538,N_6528);
nor U6673 (N_6673,N_6442,N_6460);
xor U6674 (N_6674,N_6580,N_6590);
xor U6675 (N_6675,N_6541,N_6462);
or U6676 (N_6676,N_6527,N_6578);
nor U6677 (N_6677,N_6565,N_6426);
and U6678 (N_6678,N_6584,N_6422);
nor U6679 (N_6679,N_6591,N_6432);
xnor U6680 (N_6680,N_6466,N_6505);
xor U6681 (N_6681,N_6452,N_6543);
xor U6682 (N_6682,N_6530,N_6521);
nand U6683 (N_6683,N_6592,N_6583);
nand U6684 (N_6684,N_6450,N_6560);
or U6685 (N_6685,N_6425,N_6569);
nor U6686 (N_6686,N_6483,N_6409);
or U6687 (N_6687,N_6434,N_6589);
nor U6688 (N_6688,N_6441,N_6595);
or U6689 (N_6689,N_6553,N_6568);
or U6690 (N_6690,N_6428,N_6410);
nand U6691 (N_6691,N_6495,N_6449);
and U6692 (N_6692,N_6447,N_6540);
nand U6693 (N_6693,N_6532,N_6438);
or U6694 (N_6694,N_6431,N_6457);
or U6695 (N_6695,N_6516,N_6406);
nor U6696 (N_6696,N_6557,N_6571);
nand U6697 (N_6697,N_6552,N_6537);
xor U6698 (N_6698,N_6497,N_6594);
and U6699 (N_6699,N_6480,N_6402);
xnor U6700 (N_6700,N_6516,N_6401);
nand U6701 (N_6701,N_6556,N_6547);
xnor U6702 (N_6702,N_6454,N_6534);
and U6703 (N_6703,N_6598,N_6516);
nand U6704 (N_6704,N_6492,N_6412);
or U6705 (N_6705,N_6521,N_6499);
or U6706 (N_6706,N_6477,N_6523);
nand U6707 (N_6707,N_6550,N_6536);
xor U6708 (N_6708,N_6548,N_6598);
nand U6709 (N_6709,N_6450,N_6562);
or U6710 (N_6710,N_6503,N_6505);
and U6711 (N_6711,N_6492,N_6483);
xor U6712 (N_6712,N_6544,N_6557);
nor U6713 (N_6713,N_6428,N_6440);
nor U6714 (N_6714,N_6436,N_6544);
nor U6715 (N_6715,N_6464,N_6453);
or U6716 (N_6716,N_6410,N_6475);
or U6717 (N_6717,N_6553,N_6463);
nand U6718 (N_6718,N_6596,N_6422);
or U6719 (N_6719,N_6437,N_6541);
nor U6720 (N_6720,N_6490,N_6553);
and U6721 (N_6721,N_6407,N_6542);
and U6722 (N_6722,N_6508,N_6430);
nand U6723 (N_6723,N_6582,N_6567);
or U6724 (N_6724,N_6470,N_6411);
nand U6725 (N_6725,N_6535,N_6472);
xor U6726 (N_6726,N_6589,N_6468);
nor U6727 (N_6727,N_6461,N_6424);
nor U6728 (N_6728,N_6438,N_6504);
nor U6729 (N_6729,N_6490,N_6492);
xnor U6730 (N_6730,N_6536,N_6486);
and U6731 (N_6731,N_6436,N_6534);
or U6732 (N_6732,N_6499,N_6490);
xnor U6733 (N_6733,N_6540,N_6580);
nand U6734 (N_6734,N_6507,N_6549);
nor U6735 (N_6735,N_6426,N_6562);
xnor U6736 (N_6736,N_6591,N_6481);
xor U6737 (N_6737,N_6481,N_6440);
nand U6738 (N_6738,N_6565,N_6557);
nand U6739 (N_6739,N_6434,N_6499);
and U6740 (N_6740,N_6459,N_6462);
and U6741 (N_6741,N_6590,N_6523);
xnor U6742 (N_6742,N_6419,N_6557);
and U6743 (N_6743,N_6494,N_6444);
nor U6744 (N_6744,N_6530,N_6432);
nand U6745 (N_6745,N_6441,N_6461);
or U6746 (N_6746,N_6487,N_6422);
and U6747 (N_6747,N_6504,N_6521);
xor U6748 (N_6748,N_6440,N_6526);
or U6749 (N_6749,N_6423,N_6532);
or U6750 (N_6750,N_6403,N_6470);
and U6751 (N_6751,N_6581,N_6505);
xnor U6752 (N_6752,N_6485,N_6590);
nor U6753 (N_6753,N_6475,N_6561);
xnor U6754 (N_6754,N_6587,N_6585);
nor U6755 (N_6755,N_6583,N_6439);
and U6756 (N_6756,N_6559,N_6533);
and U6757 (N_6757,N_6448,N_6536);
nand U6758 (N_6758,N_6543,N_6442);
xor U6759 (N_6759,N_6495,N_6408);
nand U6760 (N_6760,N_6573,N_6474);
and U6761 (N_6761,N_6429,N_6468);
and U6762 (N_6762,N_6432,N_6535);
and U6763 (N_6763,N_6586,N_6482);
and U6764 (N_6764,N_6452,N_6528);
xor U6765 (N_6765,N_6574,N_6507);
xnor U6766 (N_6766,N_6442,N_6520);
and U6767 (N_6767,N_6473,N_6477);
xnor U6768 (N_6768,N_6556,N_6508);
or U6769 (N_6769,N_6482,N_6481);
or U6770 (N_6770,N_6455,N_6563);
and U6771 (N_6771,N_6495,N_6437);
nor U6772 (N_6772,N_6578,N_6492);
xnor U6773 (N_6773,N_6448,N_6529);
nand U6774 (N_6774,N_6572,N_6504);
and U6775 (N_6775,N_6477,N_6552);
or U6776 (N_6776,N_6581,N_6417);
and U6777 (N_6777,N_6595,N_6533);
nor U6778 (N_6778,N_6566,N_6511);
nor U6779 (N_6779,N_6576,N_6477);
and U6780 (N_6780,N_6498,N_6554);
and U6781 (N_6781,N_6552,N_6531);
nor U6782 (N_6782,N_6596,N_6454);
or U6783 (N_6783,N_6509,N_6470);
nor U6784 (N_6784,N_6521,N_6412);
nand U6785 (N_6785,N_6431,N_6520);
xor U6786 (N_6786,N_6401,N_6441);
nand U6787 (N_6787,N_6507,N_6466);
and U6788 (N_6788,N_6506,N_6546);
nor U6789 (N_6789,N_6555,N_6594);
and U6790 (N_6790,N_6525,N_6431);
or U6791 (N_6791,N_6492,N_6452);
nand U6792 (N_6792,N_6578,N_6482);
and U6793 (N_6793,N_6473,N_6479);
xnor U6794 (N_6794,N_6447,N_6518);
xor U6795 (N_6795,N_6484,N_6485);
nand U6796 (N_6796,N_6585,N_6567);
and U6797 (N_6797,N_6434,N_6521);
and U6798 (N_6798,N_6588,N_6537);
nor U6799 (N_6799,N_6544,N_6594);
and U6800 (N_6800,N_6670,N_6704);
and U6801 (N_6801,N_6657,N_6666);
xor U6802 (N_6802,N_6684,N_6787);
or U6803 (N_6803,N_6639,N_6634);
and U6804 (N_6804,N_6614,N_6782);
xor U6805 (N_6805,N_6613,N_6638);
nor U6806 (N_6806,N_6662,N_6604);
nand U6807 (N_6807,N_6734,N_6728);
xor U6808 (N_6808,N_6789,N_6742);
and U6809 (N_6809,N_6679,N_6785);
and U6810 (N_6810,N_6671,N_6744);
and U6811 (N_6811,N_6607,N_6699);
xor U6812 (N_6812,N_6667,N_6726);
nor U6813 (N_6813,N_6621,N_6755);
and U6814 (N_6814,N_6672,N_6658);
xnor U6815 (N_6815,N_6711,N_6625);
nand U6816 (N_6816,N_6641,N_6746);
nand U6817 (N_6817,N_6636,N_6761);
xor U6818 (N_6818,N_6643,N_6722);
nor U6819 (N_6819,N_6709,N_6732);
or U6820 (N_6820,N_6647,N_6717);
or U6821 (N_6821,N_6730,N_6741);
or U6822 (N_6822,N_6688,N_6630);
nor U6823 (N_6823,N_6617,N_6645);
nand U6824 (N_6824,N_6733,N_6780);
and U6825 (N_6825,N_6788,N_6767);
nor U6826 (N_6826,N_6655,N_6791);
and U6827 (N_6827,N_6677,N_6629);
or U6828 (N_6828,N_6695,N_6651);
or U6829 (N_6829,N_6784,N_6751);
or U6830 (N_6830,N_6686,N_6696);
nand U6831 (N_6831,N_6689,N_6764);
and U6832 (N_6832,N_6674,N_6714);
nand U6833 (N_6833,N_6762,N_6627);
and U6834 (N_6834,N_6713,N_6622);
nand U6835 (N_6835,N_6752,N_6631);
or U6836 (N_6836,N_6606,N_6637);
xor U6837 (N_6837,N_6757,N_6778);
and U6838 (N_6838,N_6793,N_6602);
xor U6839 (N_6839,N_6649,N_6760);
xor U6840 (N_6840,N_6668,N_6669);
nand U6841 (N_6841,N_6745,N_6646);
or U6842 (N_6842,N_6615,N_6790);
or U6843 (N_6843,N_6798,N_6619);
and U6844 (N_6844,N_6692,N_6756);
xnor U6845 (N_6845,N_6797,N_6792);
or U6846 (N_6846,N_6623,N_6683);
nor U6847 (N_6847,N_6700,N_6640);
xor U6848 (N_6848,N_6707,N_6766);
xor U6849 (N_6849,N_6690,N_6678);
and U6850 (N_6850,N_6654,N_6676);
nor U6851 (N_6851,N_6618,N_6706);
nor U6852 (N_6852,N_6719,N_6731);
nor U6853 (N_6853,N_6697,N_6691);
or U6854 (N_6854,N_6681,N_6773);
xor U6855 (N_6855,N_6694,N_6680);
nor U6856 (N_6856,N_6796,N_6776);
or U6857 (N_6857,N_6727,N_6608);
and U6858 (N_6858,N_6781,N_6601);
xor U6859 (N_6859,N_6783,N_6663);
and U6860 (N_6860,N_6770,N_6653);
and U6861 (N_6861,N_6652,N_6754);
or U6862 (N_6862,N_6650,N_6685);
nand U6863 (N_6863,N_6774,N_6611);
nand U6864 (N_6864,N_6673,N_6624);
nand U6865 (N_6865,N_6723,N_6605);
nor U6866 (N_6866,N_6600,N_6769);
nand U6867 (N_6867,N_6725,N_6738);
and U6868 (N_6868,N_6632,N_6644);
nand U6869 (N_6869,N_6633,N_6720);
and U6870 (N_6870,N_6698,N_6708);
or U6871 (N_6871,N_6701,N_6795);
xor U6872 (N_6872,N_6628,N_6665);
nand U6873 (N_6873,N_6777,N_6664);
xnor U6874 (N_6874,N_6703,N_6712);
and U6875 (N_6875,N_6724,N_6616);
or U6876 (N_6876,N_6771,N_6675);
or U6877 (N_6877,N_6735,N_6729);
xor U6878 (N_6878,N_6612,N_6743);
nand U6879 (N_6879,N_6779,N_6693);
or U6880 (N_6880,N_6642,N_6749);
nor U6881 (N_6881,N_6705,N_6721);
and U6882 (N_6882,N_6794,N_6661);
nand U6883 (N_6883,N_6659,N_6740);
nor U6884 (N_6884,N_6660,N_6772);
nor U6885 (N_6885,N_6648,N_6750);
nand U6886 (N_6886,N_6687,N_6716);
nor U6887 (N_6887,N_6758,N_6656);
nand U6888 (N_6888,N_6710,N_6765);
nand U6889 (N_6889,N_6747,N_6609);
xor U6890 (N_6890,N_6635,N_6753);
xor U6891 (N_6891,N_6799,N_6736);
and U6892 (N_6892,N_6603,N_6786);
or U6893 (N_6893,N_6610,N_6739);
nor U6894 (N_6894,N_6682,N_6702);
and U6895 (N_6895,N_6763,N_6737);
and U6896 (N_6896,N_6775,N_6715);
xor U6897 (N_6897,N_6626,N_6748);
nor U6898 (N_6898,N_6768,N_6759);
nor U6899 (N_6899,N_6718,N_6620);
and U6900 (N_6900,N_6705,N_6725);
nand U6901 (N_6901,N_6737,N_6749);
and U6902 (N_6902,N_6614,N_6721);
or U6903 (N_6903,N_6713,N_6644);
or U6904 (N_6904,N_6786,N_6732);
nor U6905 (N_6905,N_6735,N_6638);
nor U6906 (N_6906,N_6657,N_6707);
and U6907 (N_6907,N_6778,N_6613);
and U6908 (N_6908,N_6799,N_6658);
nor U6909 (N_6909,N_6777,N_6718);
nor U6910 (N_6910,N_6656,N_6743);
xnor U6911 (N_6911,N_6624,N_6697);
and U6912 (N_6912,N_6793,N_6678);
and U6913 (N_6913,N_6681,N_6741);
nand U6914 (N_6914,N_6717,N_6725);
and U6915 (N_6915,N_6779,N_6734);
xor U6916 (N_6916,N_6670,N_6706);
or U6917 (N_6917,N_6629,N_6687);
nand U6918 (N_6918,N_6636,N_6680);
nand U6919 (N_6919,N_6756,N_6699);
xor U6920 (N_6920,N_6679,N_6659);
xor U6921 (N_6921,N_6799,N_6727);
or U6922 (N_6922,N_6622,N_6769);
nand U6923 (N_6923,N_6720,N_6729);
nor U6924 (N_6924,N_6720,N_6606);
xor U6925 (N_6925,N_6654,N_6650);
or U6926 (N_6926,N_6624,N_6715);
nor U6927 (N_6927,N_6746,N_6727);
nand U6928 (N_6928,N_6720,N_6642);
nor U6929 (N_6929,N_6725,N_6768);
and U6930 (N_6930,N_6678,N_6718);
nand U6931 (N_6931,N_6766,N_6686);
xnor U6932 (N_6932,N_6661,N_6642);
and U6933 (N_6933,N_6602,N_6637);
xnor U6934 (N_6934,N_6754,N_6610);
nor U6935 (N_6935,N_6717,N_6643);
and U6936 (N_6936,N_6742,N_6688);
and U6937 (N_6937,N_6717,N_6675);
nor U6938 (N_6938,N_6666,N_6691);
or U6939 (N_6939,N_6750,N_6610);
or U6940 (N_6940,N_6699,N_6670);
and U6941 (N_6941,N_6617,N_6619);
and U6942 (N_6942,N_6622,N_6766);
nand U6943 (N_6943,N_6736,N_6723);
or U6944 (N_6944,N_6600,N_6781);
and U6945 (N_6945,N_6706,N_6627);
xnor U6946 (N_6946,N_6761,N_6606);
or U6947 (N_6947,N_6783,N_6758);
nand U6948 (N_6948,N_6744,N_6616);
or U6949 (N_6949,N_6789,N_6776);
nor U6950 (N_6950,N_6770,N_6704);
nor U6951 (N_6951,N_6799,N_6654);
xor U6952 (N_6952,N_6708,N_6729);
nor U6953 (N_6953,N_6769,N_6751);
and U6954 (N_6954,N_6676,N_6686);
or U6955 (N_6955,N_6633,N_6791);
or U6956 (N_6956,N_6711,N_6639);
and U6957 (N_6957,N_6635,N_6795);
or U6958 (N_6958,N_6624,N_6762);
nor U6959 (N_6959,N_6625,N_6752);
xnor U6960 (N_6960,N_6615,N_6722);
nand U6961 (N_6961,N_6690,N_6709);
xor U6962 (N_6962,N_6684,N_6664);
nor U6963 (N_6963,N_6797,N_6652);
or U6964 (N_6964,N_6643,N_6610);
nand U6965 (N_6965,N_6774,N_6794);
xor U6966 (N_6966,N_6727,N_6705);
or U6967 (N_6967,N_6619,N_6775);
and U6968 (N_6968,N_6796,N_6709);
xor U6969 (N_6969,N_6756,N_6635);
or U6970 (N_6970,N_6765,N_6733);
or U6971 (N_6971,N_6708,N_6613);
xnor U6972 (N_6972,N_6615,N_6629);
nand U6973 (N_6973,N_6723,N_6662);
xor U6974 (N_6974,N_6666,N_6663);
nand U6975 (N_6975,N_6611,N_6660);
nand U6976 (N_6976,N_6709,N_6676);
and U6977 (N_6977,N_6696,N_6681);
or U6978 (N_6978,N_6749,N_6791);
and U6979 (N_6979,N_6607,N_6763);
or U6980 (N_6980,N_6715,N_6744);
nand U6981 (N_6981,N_6622,N_6788);
nand U6982 (N_6982,N_6606,N_6744);
nand U6983 (N_6983,N_6614,N_6714);
nand U6984 (N_6984,N_6739,N_6737);
xnor U6985 (N_6985,N_6765,N_6624);
xnor U6986 (N_6986,N_6636,N_6774);
or U6987 (N_6987,N_6771,N_6788);
or U6988 (N_6988,N_6752,N_6674);
and U6989 (N_6989,N_6723,N_6799);
nand U6990 (N_6990,N_6713,N_6794);
nand U6991 (N_6991,N_6702,N_6724);
or U6992 (N_6992,N_6632,N_6693);
xnor U6993 (N_6993,N_6660,N_6627);
or U6994 (N_6994,N_6733,N_6701);
and U6995 (N_6995,N_6709,N_6760);
nand U6996 (N_6996,N_6644,N_6646);
xor U6997 (N_6997,N_6790,N_6773);
xor U6998 (N_6998,N_6697,N_6783);
nand U6999 (N_6999,N_6635,N_6614);
xnor U7000 (N_7000,N_6881,N_6857);
or U7001 (N_7001,N_6862,N_6885);
xor U7002 (N_7002,N_6930,N_6842);
nor U7003 (N_7003,N_6957,N_6899);
or U7004 (N_7004,N_6947,N_6819);
nand U7005 (N_7005,N_6886,N_6806);
and U7006 (N_7006,N_6867,N_6871);
nand U7007 (N_7007,N_6964,N_6802);
xor U7008 (N_7008,N_6945,N_6998);
xnor U7009 (N_7009,N_6993,N_6810);
or U7010 (N_7010,N_6876,N_6880);
xor U7011 (N_7011,N_6996,N_6887);
or U7012 (N_7012,N_6829,N_6851);
or U7013 (N_7013,N_6831,N_6959);
or U7014 (N_7014,N_6942,N_6852);
nor U7015 (N_7015,N_6997,N_6869);
and U7016 (N_7016,N_6977,N_6960);
nand U7017 (N_7017,N_6909,N_6934);
nand U7018 (N_7018,N_6937,N_6803);
and U7019 (N_7019,N_6999,N_6965);
nor U7020 (N_7020,N_6826,N_6863);
or U7021 (N_7021,N_6815,N_6870);
xnor U7022 (N_7022,N_6984,N_6895);
nand U7023 (N_7023,N_6972,N_6818);
or U7024 (N_7024,N_6839,N_6894);
xnor U7025 (N_7025,N_6950,N_6844);
xor U7026 (N_7026,N_6820,N_6986);
xor U7027 (N_7027,N_6836,N_6994);
or U7028 (N_7028,N_6898,N_6927);
or U7029 (N_7029,N_6875,N_6859);
or U7030 (N_7030,N_6854,N_6838);
xor U7031 (N_7031,N_6985,N_6834);
xnor U7032 (N_7032,N_6958,N_6878);
nand U7033 (N_7033,N_6808,N_6888);
xnor U7034 (N_7034,N_6801,N_6969);
or U7035 (N_7035,N_6981,N_6811);
nand U7036 (N_7036,N_6865,N_6827);
xor U7037 (N_7037,N_6916,N_6879);
and U7038 (N_7038,N_6989,N_6987);
xnor U7039 (N_7039,N_6856,N_6821);
and U7040 (N_7040,N_6861,N_6906);
and U7041 (N_7041,N_6953,N_6938);
and U7042 (N_7042,N_6873,N_6943);
xor U7043 (N_7043,N_6955,N_6817);
xor U7044 (N_7044,N_6828,N_6921);
nand U7045 (N_7045,N_6814,N_6872);
or U7046 (N_7046,N_6816,N_6979);
nand U7047 (N_7047,N_6841,N_6891);
nand U7048 (N_7048,N_6860,N_6813);
xor U7049 (N_7049,N_6931,N_6807);
or U7050 (N_7050,N_6833,N_6858);
nand U7051 (N_7051,N_6935,N_6874);
nor U7052 (N_7052,N_6883,N_6922);
or U7053 (N_7053,N_6825,N_6850);
nor U7054 (N_7054,N_6974,N_6903);
and U7055 (N_7055,N_6992,N_6968);
and U7056 (N_7056,N_6956,N_6849);
xor U7057 (N_7057,N_6915,N_6951);
or U7058 (N_7058,N_6902,N_6832);
and U7059 (N_7059,N_6936,N_6809);
xnor U7060 (N_7060,N_6966,N_6991);
and U7061 (N_7061,N_6884,N_6932);
and U7062 (N_7062,N_6864,N_6948);
nand U7063 (N_7063,N_6913,N_6954);
and U7064 (N_7064,N_6904,N_6963);
and U7065 (N_7065,N_6914,N_6892);
nand U7066 (N_7066,N_6900,N_6939);
and U7067 (N_7067,N_6975,N_6917);
nand U7068 (N_7068,N_6845,N_6933);
and U7069 (N_7069,N_6855,N_6853);
nor U7070 (N_7070,N_6990,N_6848);
nand U7071 (N_7071,N_6890,N_6868);
nand U7072 (N_7072,N_6800,N_6918);
nand U7073 (N_7073,N_6846,N_6982);
xor U7074 (N_7074,N_6812,N_6988);
xnor U7075 (N_7075,N_6843,N_6924);
xnor U7076 (N_7076,N_6912,N_6940);
or U7077 (N_7077,N_6971,N_6837);
nor U7078 (N_7078,N_6823,N_6976);
nand U7079 (N_7079,N_6978,N_6926);
nor U7080 (N_7080,N_6896,N_6928);
nand U7081 (N_7081,N_6866,N_6967);
or U7082 (N_7082,N_6889,N_6952);
or U7083 (N_7083,N_6847,N_6877);
nor U7084 (N_7084,N_6944,N_6835);
nand U7085 (N_7085,N_6983,N_6946);
xor U7086 (N_7086,N_6804,N_6805);
nand U7087 (N_7087,N_6882,N_6911);
and U7088 (N_7088,N_6907,N_6980);
or U7089 (N_7089,N_6925,N_6923);
and U7090 (N_7090,N_6919,N_6961);
nor U7091 (N_7091,N_6897,N_6824);
xnor U7092 (N_7092,N_6970,N_6995);
nor U7093 (N_7093,N_6840,N_6901);
and U7094 (N_7094,N_6905,N_6941);
and U7095 (N_7095,N_6893,N_6830);
nor U7096 (N_7096,N_6973,N_6908);
or U7097 (N_7097,N_6910,N_6929);
or U7098 (N_7098,N_6822,N_6949);
nor U7099 (N_7099,N_6920,N_6962);
xnor U7100 (N_7100,N_6892,N_6967);
nor U7101 (N_7101,N_6962,N_6963);
nand U7102 (N_7102,N_6973,N_6910);
or U7103 (N_7103,N_6982,N_6868);
and U7104 (N_7104,N_6994,N_6924);
or U7105 (N_7105,N_6970,N_6845);
xor U7106 (N_7106,N_6986,N_6901);
nor U7107 (N_7107,N_6901,N_6858);
and U7108 (N_7108,N_6938,N_6827);
nor U7109 (N_7109,N_6850,N_6981);
or U7110 (N_7110,N_6909,N_6964);
nand U7111 (N_7111,N_6919,N_6953);
nand U7112 (N_7112,N_6844,N_6909);
nand U7113 (N_7113,N_6826,N_6979);
xnor U7114 (N_7114,N_6900,N_6971);
or U7115 (N_7115,N_6989,N_6992);
and U7116 (N_7116,N_6959,N_6906);
or U7117 (N_7117,N_6915,N_6887);
or U7118 (N_7118,N_6859,N_6877);
or U7119 (N_7119,N_6915,N_6972);
or U7120 (N_7120,N_6955,N_6889);
nor U7121 (N_7121,N_6901,N_6929);
nor U7122 (N_7122,N_6841,N_6802);
xor U7123 (N_7123,N_6949,N_6973);
or U7124 (N_7124,N_6932,N_6970);
xnor U7125 (N_7125,N_6849,N_6931);
nand U7126 (N_7126,N_6902,N_6934);
and U7127 (N_7127,N_6866,N_6924);
or U7128 (N_7128,N_6869,N_6933);
nand U7129 (N_7129,N_6953,N_6997);
or U7130 (N_7130,N_6810,N_6970);
and U7131 (N_7131,N_6933,N_6822);
and U7132 (N_7132,N_6950,N_6956);
or U7133 (N_7133,N_6911,N_6972);
xnor U7134 (N_7134,N_6983,N_6849);
or U7135 (N_7135,N_6931,N_6860);
xor U7136 (N_7136,N_6997,N_6803);
and U7137 (N_7137,N_6889,N_6933);
xnor U7138 (N_7138,N_6919,N_6879);
and U7139 (N_7139,N_6945,N_6876);
and U7140 (N_7140,N_6947,N_6863);
or U7141 (N_7141,N_6971,N_6889);
nand U7142 (N_7142,N_6881,N_6923);
nor U7143 (N_7143,N_6878,N_6862);
nand U7144 (N_7144,N_6985,N_6814);
nor U7145 (N_7145,N_6947,N_6873);
nor U7146 (N_7146,N_6980,N_6831);
and U7147 (N_7147,N_6823,N_6960);
or U7148 (N_7148,N_6826,N_6985);
nand U7149 (N_7149,N_6895,N_6914);
nand U7150 (N_7150,N_6934,N_6968);
nand U7151 (N_7151,N_6957,N_6833);
xor U7152 (N_7152,N_6950,N_6809);
or U7153 (N_7153,N_6981,N_6873);
and U7154 (N_7154,N_6802,N_6860);
and U7155 (N_7155,N_6877,N_6993);
nor U7156 (N_7156,N_6889,N_6847);
or U7157 (N_7157,N_6837,N_6861);
nor U7158 (N_7158,N_6940,N_6877);
or U7159 (N_7159,N_6953,N_6859);
and U7160 (N_7160,N_6827,N_6999);
nor U7161 (N_7161,N_6970,N_6920);
and U7162 (N_7162,N_6967,N_6815);
xor U7163 (N_7163,N_6896,N_6952);
xnor U7164 (N_7164,N_6974,N_6976);
and U7165 (N_7165,N_6945,N_6944);
xnor U7166 (N_7166,N_6952,N_6848);
nor U7167 (N_7167,N_6918,N_6989);
xor U7168 (N_7168,N_6969,N_6830);
and U7169 (N_7169,N_6966,N_6919);
nand U7170 (N_7170,N_6941,N_6982);
xnor U7171 (N_7171,N_6942,N_6880);
or U7172 (N_7172,N_6993,N_6852);
or U7173 (N_7173,N_6959,N_6964);
nand U7174 (N_7174,N_6850,N_6878);
xnor U7175 (N_7175,N_6812,N_6854);
xor U7176 (N_7176,N_6831,N_6948);
nor U7177 (N_7177,N_6971,N_6919);
xor U7178 (N_7178,N_6916,N_6999);
and U7179 (N_7179,N_6977,N_6914);
nor U7180 (N_7180,N_6814,N_6976);
or U7181 (N_7181,N_6886,N_6880);
xnor U7182 (N_7182,N_6907,N_6821);
nor U7183 (N_7183,N_6992,N_6993);
nand U7184 (N_7184,N_6970,N_6876);
or U7185 (N_7185,N_6949,N_6967);
nand U7186 (N_7186,N_6901,N_6833);
and U7187 (N_7187,N_6800,N_6902);
nor U7188 (N_7188,N_6886,N_6875);
or U7189 (N_7189,N_6894,N_6891);
nand U7190 (N_7190,N_6853,N_6959);
and U7191 (N_7191,N_6800,N_6846);
and U7192 (N_7192,N_6866,N_6983);
nor U7193 (N_7193,N_6941,N_6892);
nand U7194 (N_7194,N_6897,N_6902);
or U7195 (N_7195,N_6865,N_6806);
or U7196 (N_7196,N_6865,N_6918);
nor U7197 (N_7197,N_6816,N_6845);
nand U7198 (N_7198,N_6959,N_6811);
and U7199 (N_7199,N_6948,N_6910);
and U7200 (N_7200,N_7109,N_7103);
or U7201 (N_7201,N_7177,N_7152);
or U7202 (N_7202,N_7126,N_7059);
xnor U7203 (N_7203,N_7197,N_7023);
xnor U7204 (N_7204,N_7085,N_7193);
and U7205 (N_7205,N_7089,N_7105);
nand U7206 (N_7206,N_7112,N_7020);
and U7207 (N_7207,N_7130,N_7119);
nand U7208 (N_7208,N_7036,N_7117);
nand U7209 (N_7209,N_7047,N_7082);
or U7210 (N_7210,N_7066,N_7192);
and U7211 (N_7211,N_7118,N_7196);
nand U7212 (N_7212,N_7166,N_7004);
nand U7213 (N_7213,N_7186,N_7090);
nand U7214 (N_7214,N_7151,N_7058);
xor U7215 (N_7215,N_7108,N_7191);
nand U7216 (N_7216,N_7184,N_7178);
and U7217 (N_7217,N_7144,N_7024);
xor U7218 (N_7218,N_7054,N_7037);
nand U7219 (N_7219,N_7150,N_7172);
and U7220 (N_7220,N_7040,N_7005);
or U7221 (N_7221,N_7043,N_7171);
nor U7222 (N_7222,N_7042,N_7012);
nor U7223 (N_7223,N_7064,N_7159);
or U7224 (N_7224,N_7104,N_7003);
and U7225 (N_7225,N_7070,N_7162);
nor U7226 (N_7226,N_7149,N_7068);
or U7227 (N_7227,N_7028,N_7124);
nand U7228 (N_7228,N_7121,N_7132);
nand U7229 (N_7229,N_7136,N_7049);
nor U7230 (N_7230,N_7014,N_7022);
nor U7231 (N_7231,N_7176,N_7111);
xnor U7232 (N_7232,N_7065,N_7088);
nand U7233 (N_7233,N_7038,N_7034);
or U7234 (N_7234,N_7060,N_7195);
nor U7235 (N_7235,N_7135,N_7129);
or U7236 (N_7236,N_7185,N_7148);
nor U7237 (N_7237,N_7086,N_7181);
nor U7238 (N_7238,N_7173,N_7045);
nor U7239 (N_7239,N_7075,N_7027);
nor U7240 (N_7240,N_7120,N_7073);
nand U7241 (N_7241,N_7077,N_7194);
or U7242 (N_7242,N_7039,N_7025);
or U7243 (N_7243,N_7067,N_7099);
xnor U7244 (N_7244,N_7098,N_7153);
nand U7245 (N_7245,N_7123,N_7008);
xnor U7246 (N_7246,N_7163,N_7096);
nand U7247 (N_7247,N_7134,N_7026);
xor U7248 (N_7248,N_7174,N_7106);
nor U7249 (N_7249,N_7019,N_7076);
and U7250 (N_7250,N_7102,N_7001);
xor U7251 (N_7251,N_7107,N_7128);
xor U7252 (N_7252,N_7133,N_7030);
or U7253 (N_7253,N_7157,N_7018);
or U7254 (N_7254,N_7180,N_7013);
or U7255 (N_7255,N_7011,N_7168);
nor U7256 (N_7256,N_7188,N_7198);
xnor U7257 (N_7257,N_7115,N_7048);
or U7258 (N_7258,N_7140,N_7155);
nor U7259 (N_7259,N_7170,N_7138);
nand U7260 (N_7260,N_7044,N_7071);
or U7261 (N_7261,N_7051,N_7057);
and U7262 (N_7262,N_7156,N_7079);
xnor U7263 (N_7263,N_7035,N_7052);
nor U7264 (N_7264,N_7053,N_7182);
nand U7265 (N_7265,N_7160,N_7093);
and U7266 (N_7266,N_7031,N_7017);
nor U7267 (N_7267,N_7046,N_7183);
nand U7268 (N_7268,N_7116,N_7101);
or U7269 (N_7269,N_7000,N_7063);
xnor U7270 (N_7270,N_7110,N_7010);
xor U7271 (N_7271,N_7164,N_7167);
and U7272 (N_7272,N_7199,N_7145);
and U7273 (N_7273,N_7083,N_7095);
nand U7274 (N_7274,N_7032,N_7056);
nand U7275 (N_7275,N_7154,N_7141);
xor U7276 (N_7276,N_7021,N_7069);
nor U7277 (N_7277,N_7143,N_7080);
and U7278 (N_7278,N_7114,N_7165);
and U7279 (N_7279,N_7087,N_7041);
nor U7280 (N_7280,N_7007,N_7055);
nand U7281 (N_7281,N_7146,N_7158);
nor U7282 (N_7282,N_7072,N_7091);
and U7283 (N_7283,N_7006,N_7084);
nand U7284 (N_7284,N_7029,N_7127);
nand U7285 (N_7285,N_7139,N_7189);
nor U7286 (N_7286,N_7094,N_7147);
nor U7287 (N_7287,N_7097,N_7175);
nand U7288 (N_7288,N_7002,N_7100);
nand U7289 (N_7289,N_7074,N_7016);
xnor U7290 (N_7290,N_7061,N_7009);
xnor U7291 (N_7291,N_7137,N_7161);
xnor U7292 (N_7292,N_7015,N_7142);
nand U7293 (N_7293,N_7125,N_7092);
nor U7294 (N_7294,N_7062,N_7078);
nor U7295 (N_7295,N_7050,N_7190);
nor U7296 (N_7296,N_7179,N_7113);
xnor U7297 (N_7297,N_7187,N_7169);
xor U7298 (N_7298,N_7131,N_7033);
nor U7299 (N_7299,N_7081,N_7122);
xnor U7300 (N_7300,N_7045,N_7030);
or U7301 (N_7301,N_7195,N_7026);
xnor U7302 (N_7302,N_7161,N_7009);
or U7303 (N_7303,N_7034,N_7060);
nor U7304 (N_7304,N_7133,N_7052);
nand U7305 (N_7305,N_7149,N_7057);
xnor U7306 (N_7306,N_7045,N_7177);
nand U7307 (N_7307,N_7104,N_7087);
nand U7308 (N_7308,N_7038,N_7177);
nand U7309 (N_7309,N_7078,N_7166);
xor U7310 (N_7310,N_7083,N_7188);
nand U7311 (N_7311,N_7031,N_7064);
nand U7312 (N_7312,N_7103,N_7008);
or U7313 (N_7313,N_7099,N_7005);
xor U7314 (N_7314,N_7170,N_7020);
xnor U7315 (N_7315,N_7069,N_7172);
nor U7316 (N_7316,N_7176,N_7063);
or U7317 (N_7317,N_7121,N_7143);
and U7318 (N_7318,N_7052,N_7154);
nand U7319 (N_7319,N_7077,N_7030);
nor U7320 (N_7320,N_7138,N_7181);
and U7321 (N_7321,N_7049,N_7011);
nand U7322 (N_7322,N_7117,N_7065);
or U7323 (N_7323,N_7128,N_7005);
nand U7324 (N_7324,N_7085,N_7166);
nand U7325 (N_7325,N_7003,N_7025);
or U7326 (N_7326,N_7030,N_7066);
and U7327 (N_7327,N_7091,N_7013);
nand U7328 (N_7328,N_7035,N_7074);
and U7329 (N_7329,N_7132,N_7051);
nor U7330 (N_7330,N_7120,N_7162);
nor U7331 (N_7331,N_7178,N_7030);
nand U7332 (N_7332,N_7196,N_7113);
nand U7333 (N_7333,N_7141,N_7058);
and U7334 (N_7334,N_7165,N_7146);
and U7335 (N_7335,N_7153,N_7043);
nor U7336 (N_7336,N_7064,N_7197);
or U7337 (N_7337,N_7161,N_7164);
or U7338 (N_7338,N_7007,N_7134);
nor U7339 (N_7339,N_7036,N_7158);
and U7340 (N_7340,N_7179,N_7047);
and U7341 (N_7341,N_7118,N_7143);
or U7342 (N_7342,N_7010,N_7082);
xor U7343 (N_7343,N_7063,N_7068);
nor U7344 (N_7344,N_7140,N_7061);
nor U7345 (N_7345,N_7104,N_7155);
xor U7346 (N_7346,N_7065,N_7135);
nand U7347 (N_7347,N_7129,N_7198);
nand U7348 (N_7348,N_7159,N_7104);
nor U7349 (N_7349,N_7116,N_7194);
nor U7350 (N_7350,N_7178,N_7181);
xor U7351 (N_7351,N_7061,N_7074);
xnor U7352 (N_7352,N_7113,N_7103);
nand U7353 (N_7353,N_7146,N_7183);
xor U7354 (N_7354,N_7102,N_7134);
xnor U7355 (N_7355,N_7127,N_7155);
nor U7356 (N_7356,N_7157,N_7068);
or U7357 (N_7357,N_7193,N_7019);
nor U7358 (N_7358,N_7027,N_7192);
xnor U7359 (N_7359,N_7073,N_7137);
xor U7360 (N_7360,N_7018,N_7015);
and U7361 (N_7361,N_7179,N_7197);
or U7362 (N_7362,N_7054,N_7073);
xnor U7363 (N_7363,N_7153,N_7191);
or U7364 (N_7364,N_7177,N_7046);
or U7365 (N_7365,N_7122,N_7191);
nand U7366 (N_7366,N_7038,N_7187);
or U7367 (N_7367,N_7078,N_7114);
or U7368 (N_7368,N_7187,N_7115);
xnor U7369 (N_7369,N_7100,N_7028);
nand U7370 (N_7370,N_7174,N_7140);
nor U7371 (N_7371,N_7007,N_7173);
or U7372 (N_7372,N_7189,N_7118);
nand U7373 (N_7373,N_7024,N_7010);
nor U7374 (N_7374,N_7080,N_7113);
nand U7375 (N_7375,N_7031,N_7139);
xnor U7376 (N_7376,N_7007,N_7164);
and U7377 (N_7377,N_7168,N_7192);
nor U7378 (N_7378,N_7092,N_7039);
and U7379 (N_7379,N_7178,N_7036);
xnor U7380 (N_7380,N_7096,N_7149);
nand U7381 (N_7381,N_7013,N_7160);
or U7382 (N_7382,N_7037,N_7150);
xnor U7383 (N_7383,N_7190,N_7183);
and U7384 (N_7384,N_7184,N_7150);
xnor U7385 (N_7385,N_7176,N_7046);
or U7386 (N_7386,N_7040,N_7139);
and U7387 (N_7387,N_7095,N_7133);
and U7388 (N_7388,N_7048,N_7146);
nor U7389 (N_7389,N_7036,N_7153);
nor U7390 (N_7390,N_7188,N_7107);
xor U7391 (N_7391,N_7068,N_7123);
xnor U7392 (N_7392,N_7079,N_7173);
nor U7393 (N_7393,N_7005,N_7019);
nand U7394 (N_7394,N_7168,N_7021);
and U7395 (N_7395,N_7132,N_7126);
and U7396 (N_7396,N_7123,N_7119);
and U7397 (N_7397,N_7197,N_7106);
and U7398 (N_7398,N_7145,N_7126);
and U7399 (N_7399,N_7148,N_7038);
nand U7400 (N_7400,N_7366,N_7329);
xor U7401 (N_7401,N_7229,N_7263);
or U7402 (N_7402,N_7292,N_7361);
xor U7403 (N_7403,N_7286,N_7240);
and U7404 (N_7404,N_7255,N_7321);
xor U7405 (N_7405,N_7338,N_7244);
or U7406 (N_7406,N_7352,N_7228);
xor U7407 (N_7407,N_7267,N_7290);
xnor U7408 (N_7408,N_7394,N_7353);
xor U7409 (N_7409,N_7325,N_7223);
or U7410 (N_7410,N_7318,N_7306);
or U7411 (N_7411,N_7310,N_7380);
and U7412 (N_7412,N_7373,N_7268);
nand U7413 (N_7413,N_7265,N_7397);
nor U7414 (N_7414,N_7235,N_7371);
or U7415 (N_7415,N_7249,N_7294);
and U7416 (N_7416,N_7216,N_7337);
nor U7417 (N_7417,N_7354,N_7279);
and U7418 (N_7418,N_7341,N_7232);
xnor U7419 (N_7419,N_7204,N_7365);
and U7420 (N_7420,N_7209,N_7266);
nand U7421 (N_7421,N_7214,N_7393);
and U7422 (N_7422,N_7340,N_7347);
and U7423 (N_7423,N_7360,N_7331);
and U7424 (N_7424,N_7211,N_7330);
or U7425 (N_7425,N_7308,N_7281);
and U7426 (N_7426,N_7355,N_7233);
xnor U7427 (N_7427,N_7298,N_7309);
or U7428 (N_7428,N_7243,N_7297);
or U7429 (N_7429,N_7395,N_7379);
or U7430 (N_7430,N_7377,N_7324);
or U7431 (N_7431,N_7391,N_7358);
or U7432 (N_7432,N_7274,N_7207);
nand U7433 (N_7433,N_7250,N_7284);
nor U7434 (N_7434,N_7317,N_7328);
and U7435 (N_7435,N_7372,N_7200);
and U7436 (N_7436,N_7220,N_7319);
nor U7437 (N_7437,N_7231,N_7208);
xnor U7438 (N_7438,N_7261,N_7367);
xor U7439 (N_7439,N_7362,N_7217);
and U7440 (N_7440,N_7224,N_7332);
nor U7441 (N_7441,N_7226,N_7376);
and U7442 (N_7442,N_7398,N_7282);
xnor U7443 (N_7443,N_7323,N_7369);
or U7444 (N_7444,N_7262,N_7205);
nand U7445 (N_7445,N_7264,N_7320);
and U7446 (N_7446,N_7385,N_7234);
and U7447 (N_7447,N_7335,N_7212);
nor U7448 (N_7448,N_7272,N_7288);
or U7449 (N_7449,N_7351,N_7237);
or U7450 (N_7450,N_7384,N_7390);
and U7451 (N_7451,N_7239,N_7247);
or U7452 (N_7452,N_7370,N_7386);
xor U7453 (N_7453,N_7219,N_7291);
or U7454 (N_7454,N_7210,N_7333);
or U7455 (N_7455,N_7368,N_7202);
nor U7456 (N_7456,N_7388,N_7381);
and U7457 (N_7457,N_7270,N_7221);
or U7458 (N_7458,N_7280,N_7311);
nand U7459 (N_7459,N_7387,N_7343);
or U7460 (N_7460,N_7301,N_7382);
and U7461 (N_7461,N_7383,N_7322);
nor U7462 (N_7462,N_7246,N_7271);
or U7463 (N_7463,N_7345,N_7314);
xnor U7464 (N_7464,N_7206,N_7278);
nor U7465 (N_7465,N_7227,N_7349);
or U7466 (N_7466,N_7269,N_7396);
and U7467 (N_7467,N_7275,N_7339);
or U7468 (N_7468,N_7222,N_7359);
nand U7469 (N_7469,N_7277,N_7389);
or U7470 (N_7470,N_7248,N_7312);
or U7471 (N_7471,N_7399,N_7378);
and U7472 (N_7472,N_7350,N_7299);
and U7473 (N_7473,N_7225,N_7215);
xor U7474 (N_7474,N_7342,N_7236);
nand U7475 (N_7475,N_7392,N_7364);
or U7476 (N_7476,N_7287,N_7257);
nor U7477 (N_7477,N_7285,N_7241);
nor U7478 (N_7478,N_7316,N_7313);
nor U7479 (N_7479,N_7295,N_7276);
xor U7480 (N_7480,N_7327,N_7256);
nor U7481 (N_7481,N_7300,N_7303);
or U7482 (N_7482,N_7230,N_7203);
xnor U7483 (N_7483,N_7346,N_7334);
nor U7484 (N_7484,N_7289,N_7336);
or U7485 (N_7485,N_7259,N_7307);
xor U7486 (N_7486,N_7357,N_7326);
and U7487 (N_7487,N_7296,N_7348);
or U7488 (N_7488,N_7356,N_7315);
nand U7489 (N_7489,N_7213,N_7242);
or U7490 (N_7490,N_7245,N_7302);
and U7491 (N_7491,N_7283,N_7344);
nor U7492 (N_7492,N_7304,N_7258);
nor U7493 (N_7493,N_7305,N_7254);
xor U7494 (N_7494,N_7252,N_7375);
or U7495 (N_7495,N_7293,N_7260);
nand U7496 (N_7496,N_7253,N_7201);
or U7497 (N_7497,N_7218,N_7363);
nand U7498 (N_7498,N_7251,N_7238);
xnor U7499 (N_7499,N_7374,N_7273);
nor U7500 (N_7500,N_7234,N_7224);
nor U7501 (N_7501,N_7318,N_7352);
xnor U7502 (N_7502,N_7243,N_7346);
or U7503 (N_7503,N_7236,N_7223);
nand U7504 (N_7504,N_7214,N_7272);
or U7505 (N_7505,N_7396,N_7238);
or U7506 (N_7506,N_7390,N_7354);
xor U7507 (N_7507,N_7210,N_7239);
xor U7508 (N_7508,N_7234,N_7274);
and U7509 (N_7509,N_7264,N_7350);
nor U7510 (N_7510,N_7299,N_7273);
xnor U7511 (N_7511,N_7235,N_7360);
and U7512 (N_7512,N_7276,N_7366);
and U7513 (N_7513,N_7228,N_7218);
and U7514 (N_7514,N_7323,N_7229);
or U7515 (N_7515,N_7280,N_7214);
and U7516 (N_7516,N_7287,N_7269);
nor U7517 (N_7517,N_7204,N_7360);
xnor U7518 (N_7518,N_7246,N_7303);
xor U7519 (N_7519,N_7305,N_7204);
nand U7520 (N_7520,N_7255,N_7268);
or U7521 (N_7521,N_7376,N_7267);
or U7522 (N_7522,N_7355,N_7336);
xnor U7523 (N_7523,N_7391,N_7213);
nand U7524 (N_7524,N_7309,N_7280);
xor U7525 (N_7525,N_7276,N_7328);
or U7526 (N_7526,N_7300,N_7296);
and U7527 (N_7527,N_7398,N_7397);
or U7528 (N_7528,N_7376,N_7224);
or U7529 (N_7529,N_7357,N_7340);
nor U7530 (N_7530,N_7345,N_7273);
nor U7531 (N_7531,N_7249,N_7247);
xor U7532 (N_7532,N_7365,N_7287);
nor U7533 (N_7533,N_7297,N_7228);
and U7534 (N_7534,N_7295,N_7275);
xnor U7535 (N_7535,N_7355,N_7392);
xnor U7536 (N_7536,N_7331,N_7396);
xor U7537 (N_7537,N_7334,N_7289);
and U7538 (N_7538,N_7242,N_7221);
nand U7539 (N_7539,N_7290,N_7215);
nor U7540 (N_7540,N_7339,N_7377);
or U7541 (N_7541,N_7376,N_7269);
or U7542 (N_7542,N_7365,N_7356);
and U7543 (N_7543,N_7275,N_7340);
xor U7544 (N_7544,N_7298,N_7235);
nor U7545 (N_7545,N_7298,N_7308);
xor U7546 (N_7546,N_7218,N_7237);
xor U7547 (N_7547,N_7220,N_7358);
nor U7548 (N_7548,N_7200,N_7358);
and U7549 (N_7549,N_7229,N_7370);
and U7550 (N_7550,N_7352,N_7280);
xor U7551 (N_7551,N_7389,N_7261);
xnor U7552 (N_7552,N_7231,N_7355);
xnor U7553 (N_7553,N_7345,N_7230);
xor U7554 (N_7554,N_7227,N_7396);
nand U7555 (N_7555,N_7359,N_7393);
xnor U7556 (N_7556,N_7231,N_7249);
or U7557 (N_7557,N_7293,N_7305);
xnor U7558 (N_7558,N_7277,N_7394);
and U7559 (N_7559,N_7247,N_7200);
nor U7560 (N_7560,N_7225,N_7234);
nor U7561 (N_7561,N_7277,N_7311);
and U7562 (N_7562,N_7392,N_7337);
and U7563 (N_7563,N_7203,N_7228);
or U7564 (N_7564,N_7224,N_7392);
and U7565 (N_7565,N_7384,N_7296);
nand U7566 (N_7566,N_7250,N_7338);
nand U7567 (N_7567,N_7390,N_7300);
nand U7568 (N_7568,N_7369,N_7309);
xnor U7569 (N_7569,N_7264,N_7274);
xor U7570 (N_7570,N_7299,N_7265);
and U7571 (N_7571,N_7274,N_7239);
nor U7572 (N_7572,N_7206,N_7378);
and U7573 (N_7573,N_7220,N_7311);
and U7574 (N_7574,N_7212,N_7290);
nand U7575 (N_7575,N_7398,N_7309);
xnor U7576 (N_7576,N_7382,N_7391);
nor U7577 (N_7577,N_7237,N_7347);
or U7578 (N_7578,N_7353,N_7366);
and U7579 (N_7579,N_7252,N_7311);
xor U7580 (N_7580,N_7301,N_7224);
or U7581 (N_7581,N_7253,N_7304);
nor U7582 (N_7582,N_7259,N_7302);
nor U7583 (N_7583,N_7371,N_7276);
and U7584 (N_7584,N_7222,N_7339);
nor U7585 (N_7585,N_7290,N_7202);
or U7586 (N_7586,N_7242,N_7254);
xnor U7587 (N_7587,N_7233,N_7296);
and U7588 (N_7588,N_7291,N_7363);
nor U7589 (N_7589,N_7271,N_7368);
xnor U7590 (N_7590,N_7226,N_7207);
or U7591 (N_7591,N_7345,N_7386);
and U7592 (N_7592,N_7222,N_7386);
and U7593 (N_7593,N_7383,N_7307);
xor U7594 (N_7594,N_7280,N_7322);
xor U7595 (N_7595,N_7247,N_7341);
or U7596 (N_7596,N_7250,N_7393);
or U7597 (N_7597,N_7321,N_7359);
nand U7598 (N_7598,N_7250,N_7303);
or U7599 (N_7599,N_7261,N_7331);
nor U7600 (N_7600,N_7550,N_7438);
and U7601 (N_7601,N_7406,N_7512);
nor U7602 (N_7602,N_7556,N_7429);
xor U7603 (N_7603,N_7530,N_7452);
nand U7604 (N_7604,N_7595,N_7469);
nand U7605 (N_7605,N_7569,N_7422);
nand U7606 (N_7606,N_7566,N_7497);
or U7607 (N_7607,N_7509,N_7526);
nor U7608 (N_7608,N_7475,N_7579);
and U7609 (N_7609,N_7544,N_7415);
xnor U7610 (N_7610,N_7405,N_7403);
nor U7611 (N_7611,N_7559,N_7477);
or U7612 (N_7612,N_7454,N_7560);
nor U7613 (N_7613,N_7424,N_7464);
nand U7614 (N_7614,N_7553,N_7525);
or U7615 (N_7615,N_7439,N_7590);
or U7616 (N_7616,N_7598,N_7571);
or U7617 (N_7617,N_7490,N_7541);
nand U7618 (N_7618,N_7599,N_7478);
or U7619 (N_7619,N_7486,N_7518);
and U7620 (N_7620,N_7427,N_7433);
and U7621 (N_7621,N_7507,N_7549);
nand U7622 (N_7622,N_7574,N_7471);
nand U7623 (N_7623,N_7521,N_7539);
nor U7624 (N_7624,N_7505,N_7476);
nor U7625 (N_7625,N_7536,N_7514);
or U7626 (N_7626,N_7445,N_7594);
xnor U7627 (N_7627,N_7470,N_7558);
and U7628 (N_7628,N_7561,N_7565);
xnor U7629 (N_7629,N_7576,N_7531);
or U7630 (N_7630,N_7513,N_7451);
xnor U7631 (N_7631,N_7472,N_7582);
xor U7632 (N_7632,N_7435,N_7436);
xor U7633 (N_7633,N_7463,N_7444);
and U7634 (N_7634,N_7428,N_7409);
nand U7635 (N_7635,N_7504,N_7401);
and U7636 (N_7636,N_7410,N_7519);
xnor U7637 (N_7637,N_7557,N_7473);
nand U7638 (N_7638,N_7546,N_7495);
and U7639 (N_7639,N_7593,N_7529);
or U7640 (N_7640,N_7527,N_7468);
and U7641 (N_7641,N_7533,N_7440);
and U7642 (N_7642,N_7404,N_7426);
nor U7643 (N_7643,N_7414,N_7573);
xnor U7644 (N_7644,N_7417,N_7425);
nor U7645 (N_7645,N_7508,N_7583);
nor U7646 (N_7646,N_7570,N_7537);
nand U7647 (N_7647,N_7596,N_7562);
and U7648 (N_7648,N_7547,N_7466);
nand U7649 (N_7649,N_7450,N_7413);
or U7650 (N_7650,N_7586,N_7487);
nand U7651 (N_7651,N_7510,N_7453);
or U7652 (N_7652,N_7480,N_7578);
xor U7653 (N_7653,N_7502,N_7483);
and U7654 (N_7654,N_7515,N_7492);
nor U7655 (N_7655,N_7589,N_7555);
and U7656 (N_7656,N_7479,N_7551);
xnor U7657 (N_7657,N_7462,N_7460);
nand U7658 (N_7658,N_7542,N_7457);
or U7659 (N_7659,N_7482,N_7431);
xor U7660 (N_7660,N_7437,N_7420);
nor U7661 (N_7661,N_7461,N_7434);
or U7662 (N_7662,N_7488,N_7493);
xnor U7663 (N_7663,N_7489,N_7554);
or U7664 (N_7664,N_7443,N_7584);
nor U7665 (N_7665,N_7506,N_7499);
nand U7666 (N_7666,N_7592,N_7575);
and U7667 (N_7667,N_7484,N_7432);
or U7668 (N_7668,N_7418,N_7442);
nor U7669 (N_7669,N_7441,N_7552);
nand U7670 (N_7670,N_7408,N_7567);
and U7671 (N_7671,N_7416,N_7459);
nand U7672 (N_7672,N_7524,N_7516);
xor U7673 (N_7673,N_7449,N_7458);
xor U7674 (N_7674,N_7503,N_7446);
nor U7675 (N_7675,N_7522,N_7501);
and U7676 (N_7676,N_7520,N_7467);
or U7677 (N_7677,N_7581,N_7485);
or U7678 (N_7678,N_7448,N_7494);
nor U7679 (N_7679,N_7548,N_7419);
nor U7680 (N_7680,N_7421,N_7423);
nand U7681 (N_7681,N_7538,N_7474);
nand U7682 (N_7682,N_7577,N_7540);
nand U7683 (N_7683,N_7534,N_7580);
nand U7684 (N_7684,N_7587,N_7532);
and U7685 (N_7685,N_7568,N_7412);
nand U7686 (N_7686,N_7407,N_7597);
and U7687 (N_7687,N_7402,N_7585);
and U7688 (N_7688,N_7496,N_7543);
nor U7689 (N_7689,N_7511,N_7517);
xor U7690 (N_7690,N_7400,N_7500);
xor U7691 (N_7691,N_7465,N_7411);
or U7692 (N_7692,N_7545,N_7564);
xnor U7693 (N_7693,N_7498,N_7528);
and U7694 (N_7694,N_7481,N_7572);
xnor U7695 (N_7695,N_7563,N_7535);
xor U7696 (N_7696,N_7447,N_7456);
nand U7697 (N_7697,N_7455,N_7491);
nand U7698 (N_7698,N_7588,N_7523);
or U7699 (N_7699,N_7591,N_7430);
nand U7700 (N_7700,N_7469,N_7428);
xor U7701 (N_7701,N_7506,N_7413);
or U7702 (N_7702,N_7426,N_7414);
nor U7703 (N_7703,N_7457,N_7406);
nor U7704 (N_7704,N_7597,N_7518);
nand U7705 (N_7705,N_7505,N_7475);
nor U7706 (N_7706,N_7427,N_7462);
or U7707 (N_7707,N_7435,N_7504);
nor U7708 (N_7708,N_7438,N_7498);
nor U7709 (N_7709,N_7539,N_7504);
or U7710 (N_7710,N_7465,N_7400);
nand U7711 (N_7711,N_7405,N_7460);
xnor U7712 (N_7712,N_7529,N_7583);
nor U7713 (N_7713,N_7403,N_7525);
xnor U7714 (N_7714,N_7583,N_7591);
nand U7715 (N_7715,N_7568,N_7519);
and U7716 (N_7716,N_7500,N_7586);
nand U7717 (N_7717,N_7590,N_7522);
xnor U7718 (N_7718,N_7511,N_7495);
and U7719 (N_7719,N_7506,N_7555);
xnor U7720 (N_7720,N_7497,N_7561);
and U7721 (N_7721,N_7584,N_7592);
nand U7722 (N_7722,N_7541,N_7527);
and U7723 (N_7723,N_7497,N_7494);
xnor U7724 (N_7724,N_7468,N_7508);
and U7725 (N_7725,N_7576,N_7490);
xor U7726 (N_7726,N_7476,N_7518);
or U7727 (N_7727,N_7576,N_7456);
nor U7728 (N_7728,N_7567,N_7498);
xnor U7729 (N_7729,N_7436,N_7560);
or U7730 (N_7730,N_7494,N_7498);
nor U7731 (N_7731,N_7573,N_7501);
nand U7732 (N_7732,N_7570,N_7555);
nor U7733 (N_7733,N_7483,N_7407);
and U7734 (N_7734,N_7589,N_7471);
or U7735 (N_7735,N_7561,N_7406);
nor U7736 (N_7736,N_7443,N_7577);
or U7737 (N_7737,N_7507,N_7449);
nand U7738 (N_7738,N_7435,N_7599);
or U7739 (N_7739,N_7545,N_7423);
and U7740 (N_7740,N_7456,N_7572);
nand U7741 (N_7741,N_7509,N_7460);
or U7742 (N_7742,N_7560,N_7559);
nor U7743 (N_7743,N_7410,N_7422);
or U7744 (N_7744,N_7406,N_7505);
nor U7745 (N_7745,N_7411,N_7444);
nand U7746 (N_7746,N_7569,N_7576);
xnor U7747 (N_7747,N_7477,N_7446);
and U7748 (N_7748,N_7518,N_7514);
or U7749 (N_7749,N_7549,N_7442);
or U7750 (N_7750,N_7566,N_7537);
nand U7751 (N_7751,N_7428,N_7532);
or U7752 (N_7752,N_7542,N_7551);
xor U7753 (N_7753,N_7526,N_7530);
or U7754 (N_7754,N_7400,N_7476);
and U7755 (N_7755,N_7462,N_7454);
nand U7756 (N_7756,N_7465,N_7599);
xor U7757 (N_7757,N_7478,N_7476);
and U7758 (N_7758,N_7539,N_7536);
nor U7759 (N_7759,N_7457,N_7446);
and U7760 (N_7760,N_7458,N_7514);
and U7761 (N_7761,N_7560,N_7432);
and U7762 (N_7762,N_7469,N_7575);
nor U7763 (N_7763,N_7401,N_7464);
nand U7764 (N_7764,N_7545,N_7569);
nand U7765 (N_7765,N_7425,N_7590);
or U7766 (N_7766,N_7420,N_7433);
or U7767 (N_7767,N_7499,N_7511);
nand U7768 (N_7768,N_7555,N_7451);
xnor U7769 (N_7769,N_7490,N_7524);
nor U7770 (N_7770,N_7481,N_7508);
nor U7771 (N_7771,N_7590,N_7400);
nor U7772 (N_7772,N_7419,N_7497);
nor U7773 (N_7773,N_7596,N_7452);
or U7774 (N_7774,N_7423,N_7457);
or U7775 (N_7775,N_7589,N_7515);
and U7776 (N_7776,N_7493,N_7557);
nor U7777 (N_7777,N_7447,N_7551);
nand U7778 (N_7778,N_7420,N_7534);
xor U7779 (N_7779,N_7556,N_7458);
nor U7780 (N_7780,N_7574,N_7598);
or U7781 (N_7781,N_7418,N_7505);
and U7782 (N_7782,N_7520,N_7412);
or U7783 (N_7783,N_7463,N_7441);
and U7784 (N_7784,N_7587,N_7419);
xor U7785 (N_7785,N_7527,N_7459);
and U7786 (N_7786,N_7420,N_7590);
xnor U7787 (N_7787,N_7452,N_7420);
nand U7788 (N_7788,N_7524,N_7481);
nand U7789 (N_7789,N_7483,N_7589);
nand U7790 (N_7790,N_7583,N_7517);
or U7791 (N_7791,N_7508,N_7517);
nor U7792 (N_7792,N_7521,N_7431);
nor U7793 (N_7793,N_7436,N_7462);
xnor U7794 (N_7794,N_7545,N_7594);
or U7795 (N_7795,N_7564,N_7563);
nand U7796 (N_7796,N_7557,N_7556);
and U7797 (N_7797,N_7483,N_7471);
nor U7798 (N_7798,N_7449,N_7450);
xnor U7799 (N_7799,N_7552,N_7530);
nand U7800 (N_7800,N_7676,N_7626);
or U7801 (N_7801,N_7672,N_7712);
xor U7802 (N_7802,N_7754,N_7720);
xor U7803 (N_7803,N_7644,N_7699);
or U7804 (N_7804,N_7619,N_7737);
and U7805 (N_7805,N_7746,N_7731);
nand U7806 (N_7806,N_7793,N_7664);
or U7807 (N_7807,N_7740,N_7601);
and U7808 (N_7808,N_7656,N_7735);
xor U7809 (N_7809,N_7722,N_7756);
or U7810 (N_7810,N_7642,N_7772);
and U7811 (N_7811,N_7715,N_7782);
nand U7812 (N_7812,N_7713,N_7692);
nand U7813 (N_7813,N_7663,N_7788);
xnor U7814 (N_7814,N_7653,N_7693);
xor U7815 (N_7815,N_7657,N_7795);
and U7816 (N_7816,N_7602,N_7797);
and U7817 (N_7817,N_7688,N_7751);
or U7818 (N_7818,N_7783,N_7671);
and U7819 (N_7819,N_7697,N_7690);
nor U7820 (N_7820,N_7798,N_7670);
or U7821 (N_7821,N_7762,N_7630);
nor U7822 (N_7822,N_7714,N_7617);
xor U7823 (N_7823,N_7682,N_7615);
or U7824 (N_7824,N_7659,N_7652);
nand U7825 (N_7825,N_7632,N_7607);
nand U7826 (N_7826,N_7736,N_7681);
nand U7827 (N_7827,N_7745,N_7799);
nor U7828 (N_7828,N_7662,N_7766);
nor U7829 (N_7829,N_7640,N_7605);
or U7830 (N_7830,N_7684,N_7748);
xnor U7831 (N_7831,N_7734,N_7753);
xor U7832 (N_7832,N_7708,N_7628);
and U7833 (N_7833,N_7709,N_7743);
or U7834 (N_7834,N_7667,N_7647);
or U7835 (N_7835,N_7616,N_7780);
or U7836 (N_7836,N_7608,N_7711);
nand U7837 (N_7837,N_7622,N_7779);
and U7838 (N_7838,N_7778,N_7765);
nand U7839 (N_7839,N_7604,N_7627);
nor U7840 (N_7840,N_7658,N_7629);
nand U7841 (N_7841,N_7763,N_7638);
xor U7842 (N_7842,N_7755,N_7654);
nand U7843 (N_7843,N_7635,N_7660);
xnor U7844 (N_7844,N_7789,N_7678);
and U7845 (N_7845,N_7606,N_7669);
nand U7846 (N_7846,N_7760,N_7691);
or U7847 (N_7847,N_7600,N_7695);
and U7848 (N_7848,N_7764,N_7674);
and U7849 (N_7849,N_7687,N_7680);
nor U7850 (N_7850,N_7796,N_7651);
nor U7851 (N_7851,N_7750,N_7634);
or U7852 (N_7852,N_7646,N_7718);
xor U7853 (N_7853,N_7759,N_7752);
xor U7854 (N_7854,N_7790,N_7698);
nor U7855 (N_7855,N_7757,N_7641);
nand U7856 (N_7856,N_7694,N_7618);
or U7857 (N_7857,N_7744,N_7785);
nor U7858 (N_7858,N_7701,N_7729);
nor U7859 (N_7859,N_7761,N_7794);
and U7860 (N_7860,N_7774,N_7706);
or U7861 (N_7861,N_7721,N_7775);
and U7862 (N_7862,N_7683,N_7770);
or U7863 (N_7863,N_7727,N_7631);
or U7864 (N_7864,N_7771,N_7747);
xor U7865 (N_7865,N_7686,N_7645);
or U7866 (N_7866,N_7633,N_7643);
xor U7867 (N_7867,N_7625,N_7639);
and U7868 (N_7868,N_7685,N_7777);
and U7869 (N_7869,N_7749,N_7666);
xor U7870 (N_7870,N_7610,N_7741);
nor U7871 (N_7871,N_7636,N_7784);
and U7872 (N_7872,N_7738,N_7621);
or U7873 (N_7873,N_7702,N_7603);
nor U7874 (N_7874,N_7689,N_7769);
nand U7875 (N_7875,N_7637,N_7733);
nand U7876 (N_7876,N_7707,N_7661);
xor U7877 (N_7877,N_7624,N_7730);
xnor U7878 (N_7878,N_7705,N_7673);
and U7879 (N_7879,N_7649,N_7716);
xnor U7880 (N_7880,N_7696,N_7675);
nand U7881 (N_7881,N_7723,N_7700);
nand U7882 (N_7882,N_7791,N_7725);
nor U7883 (N_7883,N_7739,N_7710);
or U7884 (N_7884,N_7728,N_7665);
or U7885 (N_7885,N_7773,N_7742);
nand U7886 (N_7886,N_7623,N_7768);
nor U7887 (N_7887,N_7758,N_7655);
nor U7888 (N_7888,N_7703,N_7620);
nand U7889 (N_7889,N_7668,N_7609);
nand U7890 (N_7890,N_7613,N_7677);
nand U7891 (N_7891,N_7679,N_7732);
or U7892 (N_7892,N_7614,N_7787);
xor U7893 (N_7893,N_7792,N_7650);
xnor U7894 (N_7894,N_7719,N_7704);
nor U7895 (N_7895,N_7767,N_7717);
or U7896 (N_7896,N_7648,N_7776);
or U7897 (N_7897,N_7786,N_7724);
xor U7898 (N_7898,N_7612,N_7726);
xor U7899 (N_7899,N_7611,N_7781);
nand U7900 (N_7900,N_7727,N_7661);
and U7901 (N_7901,N_7723,N_7702);
and U7902 (N_7902,N_7771,N_7640);
nand U7903 (N_7903,N_7746,N_7678);
xnor U7904 (N_7904,N_7713,N_7656);
or U7905 (N_7905,N_7745,N_7739);
or U7906 (N_7906,N_7635,N_7683);
or U7907 (N_7907,N_7745,N_7736);
nand U7908 (N_7908,N_7662,N_7741);
xor U7909 (N_7909,N_7751,N_7658);
and U7910 (N_7910,N_7720,N_7602);
nor U7911 (N_7911,N_7760,N_7659);
or U7912 (N_7912,N_7733,N_7795);
xnor U7913 (N_7913,N_7799,N_7719);
nand U7914 (N_7914,N_7628,N_7618);
xnor U7915 (N_7915,N_7706,N_7783);
or U7916 (N_7916,N_7657,N_7641);
or U7917 (N_7917,N_7603,N_7622);
or U7918 (N_7918,N_7719,N_7698);
nand U7919 (N_7919,N_7692,N_7739);
xnor U7920 (N_7920,N_7615,N_7725);
or U7921 (N_7921,N_7685,N_7726);
or U7922 (N_7922,N_7728,N_7746);
and U7923 (N_7923,N_7644,N_7603);
nor U7924 (N_7924,N_7656,N_7682);
nand U7925 (N_7925,N_7728,N_7657);
nor U7926 (N_7926,N_7764,N_7648);
and U7927 (N_7927,N_7622,N_7770);
and U7928 (N_7928,N_7738,N_7677);
and U7929 (N_7929,N_7637,N_7611);
and U7930 (N_7930,N_7757,N_7769);
and U7931 (N_7931,N_7651,N_7606);
xnor U7932 (N_7932,N_7666,N_7625);
xor U7933 (N_7933,N_7699,N_7746);
nand U7934 (N_7934,N_7786,N_7600);
or U7935 (N_7935,N_7601,N_7795);
nor U7936 (N_7936,N_7750,N_7757);
nand U7937 (N_7937,N_7647,N_7731);
or U7938 (N_7938,N_7649,N_7796);
or U7939 (N_7939,N_7782,N_7696);
and U7940 (N_7940,N_7631,N_7624);
xnor U7941 (N_7941,N_7769,N_7742);
xor U7942 (N_7942,N_7799,N_7764);
and U7943 (N_7943,N_7690,N_7724);
nand U7944 (N_7944,N_7679,N_7786);
nand U7945 (N_7945,N_7781,N_7653);
nand U7946 (N_7946,N_7645,N_7622);
or U7947 (N_7947,N_7660,N_7735);
and U7948 (N_7948,N_7761,N_7747);
or U7949 (N_7949,N_7615,N_7739);
xnor U7950 (N_7950,N_7631,N_7671);
or U7951 (N_7951,N_7744,N_7731);
or U7952 (N_7952,N_7752,N_7756);
and U7953 (N_7953,N_7730,N_7638);
nand U7954 (N_7954,N_7615,N_7778);
or U7955 (N_7955,N_7653,N_7734);
nor U7956 (N_7956,N_7707,N_7728);
or U7957 (N_7957,N_7646,N_7724);
nand U7958 (N_7958,N_7719,N_7759);
nor U7959 (N_7959,N_7736,N_7609);
or U7960 (N_7960,N_7659,N_7736);
and U7961 (N_7961,N_7769,N_7674);
and U7962 (N_7962,N_7720,N_7792);
nor U7963 (N_7963,N_7610,N_7614);
xor U7964 (N_7964,N_7776,N_7603);
and U7965 (N_7965,N_7629,N_7702);
and U7966 (N_7966,N_7668,N_7633);
and U7967 (N_7967,N_7724,N_7706);
or U7968 (N_7968,N_7700,N_7681);
xnor U7969 (N_7969,N_7678,N_7683);
and U7970 (N_7970,N_7685,N_7796);
xnor U7971 (N_7971,N_7600,N_7617);
and U7972 (N_7972,N_7617,N_7674);
nor U7973 (N_7973,N_7725,N_7754);
or U7974 (N_7974,N_7607,N_7751);
nand U7975 (N_7975,N_7746,N_7619);
and U7976 (N_7976,N_7637,N_7687);
xnor U7977 (N_7977,N_7706,N_7645);
xnor U7978 (N_7978,N_7740,N_7766);
nor U7979 (N_7979,N_7728,N_7785);
xnor U7980 (N_7980,N_7719,N_7600);
nor U7981 (N_7981,N_7719,N_7751);
xnor U7982 (N_7982,N_7633,N_7779);
nand U7983 (N_7983,N_7630,N_7601);
nor U7984 (N_7984,N_7743,N_7733);
nand U7985 (N_7985,N_7644,N_7623);
or U7986 (N_7986,N_7699,N_7602);
and U7987 (N_7987,N_7613,N_7626);
or U7988 (N_7988,N_7705,N_7706);
and U7989 (N_7989,N_7603,N_7715);
nor U7990 (N_7990,N_7632,N_7646);
nor U7991 (N_7991,N_7727,N_7685);
nand U7992 (N_7992,N_7732,N_7683);
nor U7993 (N_7993,N_7627,N_7713);
nand U7994 (N_7994,N_7798,N_7751);
xnor U7995 (N_7995,N_7711,N_7689);
nand U7996 (N_7996,N_7635,N_7666);
xor U7997 (N_7997,N_7620,N_7702);
nand U7998 (N_7998,N_7782,N_7667);
nor U7999 (N_7999,N_7681,N_7744);
or U8000 (N_8000,N_7977,N_7983);
or U8001 (N_8001,N_7838,N_7944);
or U8002 (N_8002,N_7900,N_7876);
nor U8003 (N_8003,N_7802,N_7884);
xor U8004 (N_8004,N_7930,N_7870);
or U8005 (N_8005,N_7835,N_7975);
and U8006 (N_8006,N_7879,N_7901);
nand U8007 (N_8007,N_7817,N_7910);
nor U8008 (N_8008,N_7887,N_7927);
xnor U8009 (N_8009,N_7994,N_7890);
xor U8010 (N_8010,N_7940,N_7912);
nor U8011 (N_8011,N_7866,N_7963);
nor U8012 (N_8012,N_7855,N_7850);
nand U8013 (N_8013,N_7925,N_7996);
or U8014 (N_8014,N_7857,N_7934);
or U8015 (N_8015,N_7923,N_7935);
or U8016 (N_8016,N_7916,N_7859);
xor U8017 (N_8017,N_7810,N_7952);
xor U8018 (N_8018,N_7949,N_7874);
nand U8019 (N_8019,N_7897,N_7959);
or U8020 (N_8020,N_7929,N_7973);
and U8021 (N_8021,N_7978,N_7896);
and U8022 (N_8022,N_7889,N_7974);
xnor U8023 (N_8023,N_7836,N_7869);
xnor U8024 (N_8024,N_7989,N_7988);
or U8025 (N_8025,N_7800,N_7811);
or U8026 (N_8026,N_7843,N_7803);
nor U8027 (N_8027,N_7998,N_7909);
nor U8028 (N_8028,N_7950,N_7954);
nand U8029 (N_8029,N_7840,N_7953);
nor U8030 (N_8030,N_7958,N_7863);
nand U8031 (N_8031,N_7945,N_7961);
nand U8032 (N_8032,N_7902,N_7951);
nor U8033 (N_8033,N_7914,N_7827);
nand U8034 (N_8034,N_7832,N_7856);
nand U8035 (N_8035,N_7861,N_7862);
nor U8036 (N_8036,N_7967,N_7853);
xnor U8037 (N_8037,N_7875,N_7839);
xor U8038 (N_8038,N_7928,N_7830);
nand U8039 (N_8039,N_7898,N_7819);
nor U8040 (N_8040,N_7968,N_7846);
nor U8041 (N_8041,N_7960,N_7980);
nor U8042 (N_8042,N_7931,N_7812);
and U8043 (N_8043,N_7904,N_7921);
and U8044 (N_8044,N_7885,N_7985);
and U8045 (N_8045,N_7997,N_7993);
xnor U8046 (N_8046,N_7878,N_7882);
or U8047 (N_8047,N_7947,N_7824);
or U8048 (N_8048,N_7906,N_7871);
nand U8049 (N_8049,N_7886,N_7880);
or U8050 (N_8050,N_7804,N_7917);
or U8051 (N_8051,N_7933,N_7814);
xnor U8052 (N_8052,N_7922,N_7825);
or U8053 (N_8053,N_7913,N_7976);
xor U8054 (N_8054,N_7979,N_7971);
nor U8055 (N_8055,N_7864,N_7820);
and U8056 (N_8056,N_7808,N_7895);
and U8057 (N_8057,N_7932,N_7962);
and U8058 (N_8058,N_7833,N_7970);
xor U8059 (N_8059,N_7867,N_7848);
and U8060 (N_8060,N_7822,N_7946);
nor U8061 (N_8061,N_7956,N_7965);
xnor U8062 (N_8062,N_7926,N_7821);
and U8063 (N_8063,N_7823,N_7941);
and U8064 (N_8064,N_7992,N_7999);
or U8065 (N_8065,N_7888,N_7984);
and U8066 (N_8066,N_7936,N_7943);
nor U8067 (N_8067,N_7868,N_7986);
and U8068 (N_8068,N_7828,N_7990);
and U8069 (N_8069,N_7908,N_7842);
and U8070 (N_8070,N_7894,N_7873);
nor U8071 (N_8071,N_7877,N_7806);
nor U8072 (N_8072,N_7851,N_7981);
and U8073 (N_8073,N_7815,N_7987);
or U8074 (N_8074,N_7911,N_7858);
xor U8075 (N_8075,N_7816,N_7849);
nor U8076 (N_8076,N_7899,N_7891);
nor U8077 (N_8077,N_7964,N_7847);
xor U8078 (N_8078,N_7826,N_7915);
and U8079 (N_8079,N_7918,N_7924);
nand U8080 (N_8080,N_7893,N_7905);
or U8081 (N_8081,N_7845,N_7865);
nor U8082 (N_8082,N_7837,N_7966);
xnor U8083 (N_8083,N_7805,N_7948);
xor U8084 (N_8084,N_7807,N_7903);
and U8085 (N_8085,N_7938,N_7969);
nor U8086 (N_8086,N_7831,N_7957);
nor U8087 (N_8087,N_7982,N_7991);
and U8088 (N_8088,N_7881,N_7841);
xnor U8089 (N_8089,N_7955,N_7829);
nor U8090 (N_8090,N_7939,N_7852);
nor U8091 (N_8091,N_7995,N_7834);
nor U8092 (N_8092,N_7919,N_7818);
xor U8093 (N_8093,N_7872,N_7813);
nand U8094 (N_8094,N_7942,N_7809);
nor U8095 (N_8095,N_7920,N_7844);
nand U8096 (N_8096,N_7907,N_7801);
and U8097 (N_8097,N_7972,N_7860);
and U8098 (N_8098,N_7937,N_7883);
nand U8099 (N_8099,N_7854,N_7892);
nand U8100 (N_8100,N_7915,N_7991);
xor U8101 (N_8101,N_7915,N_7840);
xor U8102 (N_8102,N_7826,N_7894);
xor U8103 (N_8103,N_7872,N_7853);
or U8104 (N_8104,N_7960,N_7818);
and U8105 (N_8105,N_7972,N_7808);
and U8106 (N_8106,N_7903,N_7878);
xnor U8107 (N_8107,N_7944,N_7847);
and U8108 (N_8108,N_7953,N_7932);
nand U8109 (N_8109,N_7977,N_7924);
and U8110 (N_8110,N_7934,N_7820);
and U8111 (N_8111,N_7923,N_7946);
nand U8112 (N_8112,N_7928,N_7901);
and U8113 (N_8113,N_7970,N_7899);
xnor U8114 (N_8114,N_7995,N_7878);
xor U8115 (N_8115,N_7895,N_7903);
nand U8116 (N_8116,N_7853,N_7984);
nand U8117 (N_8117,N_7951,N_7866);
or U8118 (N_8118,N_7934,N_7970);
and U8119 (N_8119,N_7866,N_7995);
nor U8120 (N_8120,N_7866,N_7800);
xnor U8121 (N_8121,N_7946,N_7949);
or U8122 (N_8122,N_7867,N_7954);
or U8123 (N_8123,N_7998,N_7828);
nor U8124 (N_8124,N_7910,N_7808);
and U8125 (N_8125,N_7923,N_7998);
or U8126 (N_8126,N_7964,N_7926);
nand U8127 (N_8127,N_7982,N_7987);
nor U8128 (N_8128,N_7887,N_7861);
nor U8129 (N_8129,N_7950,N_7837);
nor U8130 (N_8130,N_7858,N_7977);
xor U8131 (N_8131,N_7990,N_7844);
and U8132 (N_8132,N_7817,N_7835);
nor U8133 (N_8133,N_7986,N_7930);
and U8134 (N_8134,N_7942,N_7913);
xor U8135 (N_8135,N_7821,N_7800);
nor U8136 (N_8136,N_7852,N_7867);
or U8137 (N_8137,N_7934,N_7942);
nand U8138 (N_8138,N_7953,N_7956);
and U8139 (N_8139,N_7824,N_7874);
nor U8140 (N_8140,N_7871,N_7898);
nor U8141 (N_8141,N_7878,N_7894);
xor U8142 (N_8142,N_7909,N_7927);
xor U8143 (N_8143,N_7906,N_7933);
xnor U8144 (N_8144,N_7981,N_7974);
or U8145 (N_8145,N_7879,N_7825);
and U8146 (N_8146,N_7950,N_7841);
nand U8147 (N_8147,N_7958,N_7894);
nor U8148 (N_8148,N_7953,N_7834);
xor U8149 (N_8149,N_7834,N_7860);
nor U8150 (N_8150,N_7939,N_7981);
or U8151 (N_8151,N_7889,N_7818);
nor U8152 (N_8152,N_7876,N_7819);
and U8153 (N_8153,N_7854,N_7898);
nand U8154 (N_8154,N_7999,N_7903);
xnor U8155 (N_8155,N_7841,N_7921);
nand U8156 (N_8156,N_7911,N_7870);
or U8157 (N_8157,N_7902,N_7991);
nor U8158 (N_8158,N_7999,N_7836);
and U8159 (N_8159,N_7971,N_7966);
and U8160 (N_8160,N_7847,N_7814);
or U8161 (N_8161,N_7904,N_7913);
nand U8162 (N_8162,N_7846,N_7955);
nor U8163 (N_8163,N_7859,N_7902);
or U8164 (N_8164,N_7800,N_7877);
nand U8165 (N_8165,N_7823,N_7876);
nor U8166 (N_8166,N_7850,N_7830);
nor U8167 (N_8167,N_7884,N_7811);
or U8168 (N_8168,N_7892,N_7963);
and U8169 (N_8169,N_7931,N_7937);
nand U8170 (N_8170,N_7869,N_7938);
and U8171 (N_8171,N_7912,N_7833);
or U8172 (N_8172,N_7966,N_7902);
nor U8173 (N_8173,N_7901,N_7984);
and U8174 (N_8174,N_7961,N_7812);
nand U8175 (N_8175,N_7847,N_7893);
xnor U8176 (N_8176,N_7897,N_7913);
nor U8177 (N_8177,N_7904,N_7985);
or U8178 (N_8178,N_7942,N_7886);
or U8179 (N_8179,N_7802,N_7891);
and U8180 (N_8180,N_7965,N_7845);
xnor U8181 (N_8181,N_7894,N_7875);
xor U8182 (N_8182,N_7886,N_7867);
or U8183 (N_8183,N_7901,N_7897);
nor U8184 (N_8184,N_7834,N_7917);
xnor U8185 (N_8185,N_7935,N_7997);
and U8186 (N_8186,N_7882,N_7879);
and U8187 (N_8187,N_7814,N_7875);
nand U8188 (N_8188,N_7941,N_7889);
or U8189 (N_8189,N_7832,N_7896);
or U8190 (N_8190,N_7876,N_7962);
or U8191 (N_8191,N_7935,N_7874);
nand U8192 (N_8192,N_7972,N_7919);
nor U8193 (N_8193,N_7854,N_7951);
and U8194 (N_8194,N_7801,N_7954);
nor U8195 (N_8195,N_7817,N_7822);
or U8196 (N_8196,N_7947,N_7831);
xor U8197 (N_8197,N_7889,N_7828);
and U8198 (N_8198,N_7824,N_7800);
xor U8199 (N_8199,N_7927,N_7939);
nand U8200 (N_8200,N_8100,N_8063);
xnor U8201 (N_8201,N_8066,N_8157);
nor U8202 (N_8202,N_8046,N_8134);
xor U8203 (N_8203,N_8081,N_8142);
or U8204 (N_8204,N_8003,N_8088);
or U8205 (N_8205,N_8035,N_8159);
and U8206 (N_8206,N_8069,N_8004);
or U8207 (N_8207,N_8094,N_8020);
xnor U8208 (N_8208,N_8008,N_8022);
xor U8209 (N_8209,N_8018,N_8045);
and U8210 (N_8210,N_8122,N_8039);
or U8211 (N_8211,N_8087,N_8176);
nor U8212 (N_8212,N_8034,N_8080);
xor U8213 (N_8213,N_8179,N_8047);
nand U8214 (N_8214,N_8058,N_8108);
xnor U8215 (N_8215,N_8148,N_8114);
or U8216 (N_8216,N_8167,N_8196);
nand U8217 (N_8217,N_8186,N_8064);
or U8218 (N_8218,N_8185,N_8151);
and U8219 (N_8219,N_8191,N_8060);
xnor U8220 (N_8220,N_8120,N_8197);
nor U8221 (N_8221,N_8101,N_8001);
nor U8222 (N_8222,N_8077,N_8127);
nand U8223 (N_8223,N_8011,N_8175);
or U8224 (N_8224,N_8147,N_8014);
and U8225 (N_8225,N_8017,N_8160);
xnor U8226 (N_8226,N_8051,N_8109);
or U8227 (N_8227,N_8059,N_8164);
or U8228 (N_8228,N_8118,N_8023);
nand U8229 (N_8229,N_8139,N_8103);
nand U8230 (N_8230,N_8005,N_8061);
or U8231 (N_8231,N_8161,N_8082);
and U8232 (N_8232,N_8187,N_8123);
xor U8233 (N_8233,N_8140,N_8054);
nor U8234 (N_8234,N_8053,N_8162);
nand U8235 (N_8235,N_8062,N_8195);
or U8236 (N_8236,N_8068,N_8188);
or U8237 (N_8237,N_8007,N_8036);
nor U8238 (N_8238,N_8073,N_8032);
and U8239 (N_8239,N_8026,N_8070);
xor U8240 (N_8240,N_8093,N_8130);
nand U8241 (N_8241,N_8010,N_8178);
or U8242 (N_8242,N_8121,N_8021);
nor U8243 (N_8243,N_8099,N_8057);
xor U8244 (N_8244,N_8075,N_8155);
and U8245 (N_8245,N_8015,N_8166);
nand U8246 (N_8246,N_8016,N_8171);
and U8247 (N_8247,N_8193,N_8030);
or U8248 (N_8248,N_8145,N_8044);
nor U8249 (N_8249,N_8144,N_8091);
or U8250 (N_8250,N_8071,N_8141);
nand U8251 (N_8251,N_8084,N_8183);
xor U8252 (N_8252,N_8174,N_8168);
nand U8253 (N_8253,N_8050,N_8138);
or U8254 (N_8254,N_8095,N_8156);
or U8255 (N_8255,N_8189,N_8042);
nand U8256 (N_8256,N_8025,N_8079);
nand U8257 (N_8257,N_8043,N_8110);
nand U8258 (N_8258,N_8096,N_8158);
and U8259 (N_8259,N_8078,N_8124);
or U8260 (N_8260,N_8119,N_8169);
or U8261 (N_8261,N_8040,N_8028);
xnor U8262 (N_8262,N_8177,N_8131);
nor U8263 (N_8263,N_8170,N_8086);
nand U8264 (N_8264,N_8019,N_8146);
or U8265 (N_8265,N_8048,N_8098);
nor U8266 (N_8266,N_8085,N_8113);
nor U8267 (N_8267,N_8083,N_8037);
and U8268 (N_8268,N_8194,N_8106);
xor U8269 (N_8269,N_8067,N_8190);
or U8270 (N_8270,N_8027,N_8182);
and U8271 (N_8271,N_8136,N_8024);
and U8272 (N_8272,N_8065,N_8107);
nand U8273 (N_8273,N_8089,N_8104);
or U8274 (N_8274,N_8143,N_8002);
or U8275 (N_8275,N_8149,N_8135);
nand U8276 (N_8276,N_8115,N_8013);
or U8277 (N_8277,N_8125,N_8097);
and U8278 (N_8278,N_8116,N_8126);
nand U8279 (N_8279,N_8192,N_8092);
and U8280 (N_8280,N_8128,N_8076);
and U8281 (N_8281,N_8111,N_8012);
or U8282 (N_8282,N_8041,N_8009);
nor U8283 (N_8283,N_8033,N_8000);
and U8284 (N_8284,N_8112,N_8006);
xnor U8285 (N_8285,N_8199,N_8133);
and U8286 (N_8286,N_8055,N_8137);
or U8287 (N_8287,N_8105,N_8198);
and U8288 (N_8288,N_8038,N_8117);
xor U8289 (N_8289,N_8172,N_8165);
xnor U8290 (N_8290,N_8180,N_8074);
or U8291 (N_8291,N_8181,N_8184);
xor U8292 (N_8292,N_8056,N_8052);
and U8293 (N_8293,N_8163,N_8150);
xor U8294 (N_8294,N_8031,N_8102);
nor U8295 (N_8295,N_8173,N_8049);
nor U8296 (N_8296,N_8152,N_8072);
xor U8297 (N_8297,N_8154,N_8153);
nor U8298 (N_8298,N_8090,N_8132);
and U8299 (N_8299,N_8029,N_8129);
nor U8300 (N_8300,N_8068,N_8195);
or U8301 (N_8301,N_8144,N_8116);
nor U8302 (N_8302,N_8009,N_8092);
nor U8303 (N_8303,N_8172,N_8057);
xor U8304 (N_8304,N_8105,N_8003);
or U8305 (N_8305,N_8159,N_8185);
nand U8306 (N_8306,N_8003,N_8002);
nor U8307 (N_8307,N_8085,N_8048);
nor U8308 (N_8308,N_8041,N_8180);
nand U8309 (N_8309,N_8025,N_8182);
xor U8310 (N_8310,N_8050,N_8162);
nand U8311 (N_8311,N_8108,N_8183);
xnor U8312 (N_8312,N_8018,N_8149);
nor U8313 (N_8313,N_8054,N_8195);
and U8314 (N_8314,N_8110,N_8034);
or U8315 (N_8315,N_8115,N_8032);
or U8316 (N_8316,N_8015,N_8033);
xnor U8317 (N_8317,N_8192,N_8130);
xnor U8318 (N_8318,N_8024,N_8043);
nand U8319 (N_8319,N_8094,N_8071);
xor U8320 (N_8320,N_8028,N_8162);
nor U8321 (N_8321,N_8140,N_8184);
nand U8322 (N_8322,N_8183,N_8160);
nor U8323 (N_8323,N_8048,N_8145);
xor U8324 (N_8324,N_8088,N_8197);
and U8325 (N_8325,N_8198,N_8166);
and U8326 (N_8326,N_8040,N_8161);
nor U8327 (N_8327,N_8183,N_8167);
or U8328 (N_8328,N_8079,N_8158);
or U8329 (N_8329,N_8100,N_8030);
nand U8330 (N_8330,N_8077,N_8017);
nor U8331 (N_8331,N_8105,N_8093);
or U8332 (N_8332,N_8148,N_8158);
and U8333 (N_8333,N_8096,N_8017);
nand U8334 (N_8334,N_8072,N_8198);
nand U8335 (N_8335,N_8165,N_8157);
nand U8336 (N_8336,N_8088,N_8040);
nor U8337 (N_8337,N_8054,N_8076);
and U8338 (N_8338,N_8192,N_8015);
and U8339 (N_8339,N_8161,N_8182);
and U8340 (N_8340,N_8166,N_8101);
nor U8341 (N_8341,N_8104,N_8102);
nor U8342 (N_8342,N_8093,N_8181);
or U8343 (N_8343,N_8102,N_8198);
nand U8344 (N_8344,N_8048,N_8190);
nand U8345 (N_8345,N_8002,N_8184);
xor U8346 (N_8346,N_8189,N_8106);
and U8347 (N_8347,N_8156,N_8097);
nor U8348 (N_8348,N_8060,N_8112);
nand U8349 (N_8349,N_8181,N_8177);
or U8350 (N_8350,N_8143,N_8029);
or U8351 (N_8351,N_8095,N_8090);
nand U8352 (N_8352,N_8063,N_8193);
and U8353 (N_8353,N_8116,N_8060);
xnor U8354 (N_8354,N_8072,N_8134);
xnor U8355 (N_8355,N_8066,N_8150);
or U8356 (N_8356,N_8002,N_8083);
and U8357 (N_8357,N_8156,N_8078);
or U8358 (N_8358,N_8090,N_8138);
nand U8359 (N_8359,N_8134,N_8198);
or U8360 (N_8360,N_8118,N_8151);
nor U8361 (N_8361,N_8180,N_8106);
nand U8362 (N_8362,N_8181,N_8037);
nand U8363 (N_8363,N_8184,N_8094);
nor U8364 (N_8364,N_8191,N_8148);
or U8365 (N_8365,N_8119,N_8096);
and U8366 (N_8366,N_8183,N_8002);
xnor U8367 (N_8367,N_8074,N_8121);
or U8368 (N_8368,N_8159,N_8093);
or U8369 (N_8369,N_8167,N_8058);
and U8370 (N_8370,N_8114,N_8134);
nor U8371 (N_8371,N_8085,N_8194);
and U8372 (N_8372,N_8027,N_8141);
nand U8373 (N_8373,N_8179,N_8184);
nor U8374 (N_8374,N_8055,N_8124);
xor U8375 (N_8375,N_8121,N_8110);
or U8376 (N_8376,N_8073,N_8157);
and U8377 (N_8377,N_8148,N_8179);
or U8378 (N_8378,N_8040,N_8195);
and U8379 (N_8379,N_8195,N_8053);
nor U8380 (N_8380,N_8192,N_8071);
nor U8381 (N_8381,N_8190,N_8110);
nor U8382 (N_8382,N_8003,N_8018);
or U8383 (N_8383,N_8029,N_8149);
xnor U8384 (N_8384,N_8032,N_8104);
xnor U8385 (N_8385,N_8179,N_8098);
and U8386 (N_8386,N_8026,N_8008);
and U8387 (N_8387,N_8024,N_8174);
xnor U8388 (N_8388,N_8026,N_8181);
or U8389 (N_8389,N_8071,N_8185);
xnor U8390 (N_8390,N_8111,N_8135);
and U8391 (N_8391,N_8024,N_8153);
xor U8392 (N_8392,N_8033,N_8195);
or U8393 (N_8393,N_8066,N_8065);
nand U8394 (N_8394,N_8111,N_8136);
xor U8395 (N_8395,N_8182,N_8197);
and U8396 (N_8396,N_8002,N_8082);
nor U8397 (N_8397,N_8005,N_8153);
or U8398 (N_8398,N_8142,N_8199);
or U8399 (N_8399,N_8120,N_8041);
nor U8400 (N_8400,N_8346,N_8316);
and U8401 (N_8401,N_8341,N_8280);
xor U8402 (N_8402,N_8345,N_8373);
nand U8403 (N_8403,N_8229,N_8201);
or U8404 (N_8404,N_8392,N_8340);
or U8405 (N_8405,N_8378,N_8384);
nand U8406 (N_8406,N_8352,N_8317);
xor U8407 (N_8407,N_8302,N_8292);
nand U8408 (N_8408,N_8290,N_8236);
xnor U8409 (N_8409,N_8295,N_8315);
nand U8410 (N_8410,N_8283,N_8233);
nand U8411 (N_8411,N_8342,N_8337);
or U8412 (N_8412,N_8370,N_8354);
or U8413 (N_8413,N_8360,N_8227);
or U8414 (N_8414,N_8329,N_8322);
nor U8415 (N_8415,N_8278,N_8323);
xor U8416 (N_8416,N_8257,N_8299);
nand U8417 (N_8417,N_8301,N_8297);
and U8418 (N_8418,N_8399,N_8205);
or U8419 (N_8419,N_8335,N_8330);
nor U8420 (N_8420,N_8397,N_8394);
xor U8421 (N_8421,N_8287,N_8222);
or U8422 (N_8422,N_8310,N_8237);
and U8423 (N_8423,N_8367,N_8389);
or U8424 (N_8424,N_8303,N_8253);
nor U8425 (N_8425,N_8348,N_8324);
xnor U8426 (N_8426,N_8379,N_8272);
xnor U8427 (N_8427,N_8234,N_8251);
nand U8428 (N_8428,N_8262,N_8261);
nor U8429 (N_8429,N_8286,N_8217);
nand U8430 (N_8430,N_8291,N_8239);
nor U8431 (N_8431,N_8393,N_8339);
and U8432 (N_8432,N_8318,N_8336);
nand U8433 (N_8433,N_8380,N_8264);
nand U8434 (N_8434,N_8351,N_8396);
nand U8435 (N_8435,N_8349,N_8238);
and U8436 (N_8436,N_8383,N_8288);
or U8437 (N_8437,N_8395,N_8304);
xnor U8438 (N_8438,N_8377,N_8214);
and U8439 (N_8439,N_8271,N_8333);
xnor U8440 (N_8440,N_8281,N_8265);
xnor U8441 (N_8441,N_8343,N_8248);
xor U8442 (N_8442,N_8366,N_8215);
or U8443 (N_8443,N_8307,N_8213);
nand U8444 (N_8444,N_8279,N_8244);
nor U8445 (N_8445,N_8321,N_8332);
and U8446 (N_8446,N_8277,N_8259);
nand U8447 (N_8447,N_8356,N_8296);
and U8448 (N_8448,N_8359,N_8344);
nor U8449 (N_8449,N_8243,N_8365);
nor U8450 (N_8450,N_8350,N_8211);
nor U8451 (N_8451,N_8230,N_8221);
nor U8452 (N_8452,N_8391,N_8282);
and U8453 (N_8453,N_8212,N_8362);
or U8454 (N_8454,N_8347,N_8293);
nand U8455 (N_8455,N_8328,N_8206);
nor U8456 (N_8456,N_8326,N_8270);
nand U8457 (N_8457,N_8255,N_8249);
or U8458 (N_8458,N_8358,N_8273);
or U8459 (N_8459,N_8285,N_8325);
nor U8460 (N_8460,N_8247,N_8269);
or U8461 (N_8461,N_8202,N_8266);
or U8462 (N_8462,N_8240,N_8388);
or U8463 (N_8463,N_8241,N_8220);
nor U8464 (N_8464,N_8294,N_8235);
and U8465 (N_8465,N_8331,N_8312);
nand U8466 (N_8466,N_8226,N_8254);
or U8467 (N_8467,N_8232,N_8387);
or U8468 (N_8468,N_8245,N_8225);
nor U8469 (N_8469,N_8231,N_8313);
nor U8470 (N_8470,N_8275,N_8203);
nor U8471 (N_8471,N_8372,N_8258);
or U8472 (N_8472,N_8308,N_8228);
xnor U8473 (N_8473,N_8224,N_8267);
xor U8474 (N_8474,N_8371,N_8361);
and U8475 (N_8475,N_8207,N_8306);
or U8476 (N_8476,N_8376,N_8256);
xor U8477 (N_8477,N_8320,N_8338);
and U8478 (N_8478,N_8305,N_8390);
nor U8479 (N_8479,N_8219,N_8210);
nand U8480 (N_8480,N_8375,N_8398);
xor U8481 (N_8481,N_8309,N_8289);
or U8482 (N_8482,N_8334,N_8268);
nor U8483 (N_8483,N_8216,N_8357);
nor U8484 (N_8484,N_8223,N_8386);
nand U8485 (N_8485,N_8385,N_8208);
and U8486 (N_8486,N_8327,N_8369);
and U8487 (N_8487,N_8276,N_8252);
nand U8488 (N_8488,N_8298,N_8274);
nor U8489 (N_8489,N_8300,N_8374);
nand U8490 (N_8490,N_8263,N_8246);
and U8491 (N_8491,N_8218,N_8260);
or U8492 (N_8492,N_8355,N_8314);
nand U8493 (N_8493,N_8319,N_8353);
and U8494 (N_8494,N_8204,N_8381);
nor U8495 (N_8495,N_8209,N_8200);
xor U8496 (N_8496,N_8364,N_8363);
or U8497 (N_8497,N_8382,N_8311);
xnor U8498 (N_8498,N_8368,N_8284);
xnor U8499 (N_8499,N_8250,N_8242);
and U8500 (N_8500,N_8218,N_8217);
nor U8501 (N_8501,N_8223,N_8306);
xor U8502 (N_8502,N_8275,N_8313);
nor U8503 (N_8503,N_8242,N_8246);
nor U8504 (N_8504,N_8346,N_8304);
nor U8505 (N_8505,N_8252,N_8220);
nor U8506 (N_8506,N_8241,N_8269);
or U8507 (N_8507,N_8224,N_8275);
nor U8508 (N_8508,N_8354,N_8294);
nand U8509 (N_8509,N_8225,N_8259);
and U8510 (N_8510,N_8386,N_8305);
or U8511 (N_8511,N_8353,N_8366);
nor U8512 (N_8512,N_8223,N_8283);
xnor U8513 (N_8513,N_8380,N_8276);
nor U8514 (N_8514,N_8294,N_8360);
or U8515 (N_8515,N_8339,N_8284);
nor U8516 (N_8516,N_8396,N_8303);
nor U8517 (N_8517,N_8314,N_8320);
nor U8518 (N_8518,N_8368,N_8236);
or U8519 (N_8519,N_8367,N_8396);
nor U8520 (N_8520,N_8273,N_8356);
xor U8521 (N_8521,N_8256,N_8379);
nand U8522 (N_8522,N_8281,N_8350);
nand U8523 (N_8523,N_8296,N_8329);
nor U8524 (N_8524,N_8235,N_8338);
or U8525 (N_8525,N_8218,N_8234);
and U8526 (N_8526,N_8349,N_8324);
or U8527 (N_8527,N_8264,N_8340);
nand U8528 (N_8528,N_8250,N_8300);
nand U8529 (N_8529,N_8292,N_8340);
or U8530 (N_8530,N_8265,N_8396);
nand U8531 (N_8531,N_8201,N_8389);
and U8532 (N_8532,N_8315,N_8225);
nor U8533 (N_8533,N_8265,N_8212);
xor U8534 (N_8534,N_8251,N_8252);
and U8535 (N_8535,N_8352,N_8357);
and U8536 (N_8536,N_8221,N_8217);
or U8537 (N_8537,N_8317,N_8286);
or U8538 (N_8538,N_8296,N_8266);
nand U8539 (N_8539,N_8247,N_8337);
or U8540 (N_8540,N_8309,N_8285);
or U8541 (N_8541,N_8238,N_8270);
and U8542 (N_8542,N_8338,N_8315);
nand U8543 (N_8543,N_8257,N_8374);
nor U8544 (N_8544,N_8248,N_8351);
and U8545 (N_8545,N_8224,N_8337);
nand U8546 (N_8546,N_8326,N_8329);
or U8547 (N_8547,N_8252,N_8259);
nor U8548 (N_8548,N_8296,N_8229);
and U8549 (N_8549,N_8219,N_8207);
or U8550 (N_8550,N_8359,N_8230);
nand U8551 (N_8551,N_8333,N_8370);
or U8552 (N_8552,N_8328,N_8263);
xnor U8553 (N_8553,N_8308,N_8399);
xnor U8554 (N_8554,N_8364,N_8315);
nand U8555 (N_8555,N_8385,N_8366);
or U8556 (N_8556,N_8237,N_8366);
nand U8557 (N_8557,N_8322,N_8248);
and U8558 (N_8558,N_8275,N_8381);
nand U8559 (N_8559,N_8338,N_8357);
or U8560 (N_8560,N_8335,N_8391);
nand U8561 (N_8561,N_8356,N_8263);
xnor U8562 (N_8562,N_8365,N_8298);
or U8563 (N_8563,N_8354,N_8248);
nand U8564 (N_8564,N_8397,N_8287);
nand U8565 (N_8565,N_8269,N_8369);
and U8566 (N_8566,N_8304,N_8384);
nor U8567 (N_8567,N_8226,N_8259);
xnor U8568 (N_8568,N_8287,N_8221);
xor U8569 (N_8569,N_8237,N_8374);
nor U8570 (N_8570,N_8340,N_8341);
and U8571 (N_8571,N_8335,N_8268);
xor U8572 (N_8572,N_8206,N_8360);
nor U8573 (N_8573,N_8322,N_8275);
nand U8574 (N_8574,N_8208,N_8353);
nand U8575 (N_8575,N_8358,N_8384);
nor U8576 (N_8576,N_8331,N_8397);
or U8577 (N_8577,N_8342,N_8269);
nor U8578 (N_8578,N_8352,N_8214);
nor U8579 (N_8579,N_8276,N_8321);
or U8580 (N_8580,N_8368,N_8270);
xnor U8581 (N_8581,N_8362,N_8322);
xor U8582 (N_8582,N_8374,N_8358);
xor U8583 (N_8583,N_8338,N_8229);
xor U8584 (N_8584,N_8365,N_8277);
xor U8585 (N_8585,N_8235,N_8344);
and U8586 (N_8586,N_8210,N_8267);
or U8587 (N_8587,N_8204,N_8219);
nor U8588 (N_8588,N_8240,N_8239);
or U8589 (N_8589,N_8297,N_8326);
nor U8590 (N_8590,N_8383,N_8264);
or U8591 (N_8591,N_8365,N_8387);
and U8592 (N_8592,N_8380,N_8295);
xor U8593 (N_8593,N_8267,N_8312);
or U8594 (N_8594,N_8201,N_8288);
nor U8595 (N_8595,N_8239,N_8382);
xnor U8596 (N_8596,N_8368,N_8202);
nor U8597 (N_8597,N_8324,N_8357);
xnor U8598 (N_8598,N_8311,N_8302);
nor U8599 (N_8599,N_8356,N_8291);
nand U8600 (N_8600,N_8551,N_8469);
xor U8601 (N_8601,N_8425,N_8460);
or U8602 (N_8602,N_8466,N_8567);
or U8603 (N_8603,N_8413,N_8497);
or U8604 (N_8604,N_8417,N_8562);
and U8605 (N_8605,N_8522,N_8412);
xnor U8606 (N_8606,N_8570,N_8426);
and U8607 (N_8607,N_8490,N_8411);
or U8608 (N_8608,N_8442,N_8408);
xor U8609 (N_8609,N_8509,N_8564);
or U8610 (N_8610,N_8597,N_8448);
nor U8611 (N_8611,N_8540,N_8410);
and U8612 (N_8612,N_8557,N_8505);
xnor U8613 (N_8613,N_8534,N_8471);
nor U8614 (N_8614,N_8544,N_8599);
or U8615 (N_8615,N_8496,N_8571);
xnor U8616 (N_8616,N_8431,N_8456);
nand U8617 (N_8617,N_8553,N_8515);
nand U8618 (N_8618,N_8424,N_8483);
or U8619 (N_8619,N_8578,N_8545);
and U8620 (N_8620,N_8576,N_8434);
nor U8621 (N_8621,N_8559,N_8439);
nor U8622 (N_8622,N_8577,N_8519);
or U8623 (N_8623,N_8558,N_8445);
or U8624 (N_8624,N_8430,N_8579);
and U8625 (N_8625,N_8446,N_8414);
or U8626 (N_8626,N_8504,N_8407);
and U8627 (N_8627,N_8594,N_8563);
xnor U8628 (N_8628,N_8533,N_8512);
and U8629 (N_8629,N_8472,N_8555);
nor U8630 (N_8630,N_8421,N_8473);
nand U8631 (N_8631,N_8574,N_8569);
or U8632 (N_8632,N_8548,N_8423);
nor U8633 (N_8633,N_8476,N_8573);
nor U8634 (N_8634,N_8531,N_8590);
xnor U8635 (N_8635,N_8420,N_8532);
and U8636 (N_8636,N_8543,N_8575);
or U8637 (N_8637,N_8595,N_8494);
nand U8638 (N_8638,N_8463,N_8582);
xor U8639 (N_8639,N_8539,N_8556);
nand U8640 (N_8640,N_8542,N_8524);
or U8641 (N_8641,N_8457,N_8580);
nor U8642 (N_8642,N_8514,N_8478);
or U8643 (N_8643,N_8429,N_8596);
nor U8644 (N_8644,N_8440,N_8458);
or U8645 (N_8645,N_8529,N_8589);
nor U8646 (N_8646,N_8453,N_8493);
nand U8647 (N_8647,N_8501,N_8526);
and U8648 (N_8648,N_8550,N_8527);
or U8649 (N_8649,N_8403,N_8565);
and U8650 (N_8650,N_8485,N_8549);
nand U8651 (N_8651,N_8450,N_8554);
and U8652 (N_8652,N_8419,N_8462);
and U8653 (N_8653,N_8481,N_8518);
xor U8654 (N_8654,N_8464,N_8468);
nand U8655 (N_8655,N_8435,N_8588);
xnor U8656 (N_8656,N_8523,N_8441);
nand U8657 (N_8657,N_8491,N_8593);
xnor U8658 (N_8658,N_8428,N_8418);
or U8659 (N_8659,N_8443,N_8492);
and U8660 (N_8660,N_8475,N_8547);
and U8661 (N_8661,N_8535,N_8400);
or U8662 (N_8662,N_8467,N_8487);
xor U8663 (N_8663,N_8516,N_8499);
or U8664 (N_8664,N_8479,N_8538);
or U8665 (N_8665,N_8585,N_8454);
nand U8666 (N_8666,N_8511,N_8572);
nor U8667 (N_8667,N_8508,N_8488);
or U8668 (N_8668,N_8525,N_8452);
nand U8669 (N_8669,N_8506,N_8402);
and U8670 (N_8670,N_8586,N_8474);
xnor U8671 (N_8671,N_8500,N_8432);
or U8672 (N_8672,N_8484,N_8447);
xnor U8673 (N_8673,N_8530,N_8401);
nor U8674 (N_8674,N_8502,N_8489);
xnor U8675 (N_8675,N_8480,N_8438);
nand U8676 (N_8676,N_8536,N_8404);
nand U8677 (N_8677,N_8409,N_8507);
nand U8678 (N_8678,N_8433,N_8498);
nor U8679 (N_8679,N_8477,N_8405);
and U8680 (N_8680,N_8406,N_8455);
and U8681 (N_8681,N_8465,N_8470);
nand U8682 (N_8682,N_8459,N_8510);
nand U8683 (N_8683,N_8560,N_8427);
and U8684 (N_8684,N_8561,N_8486);
nor U8685 (N_8685,N_8546,N_8581);
and U8686 (N_8686,N_8591,N_8598);
or U8687 (N_8687,N_8587,N_8449);
nand U8688 (N_8688,N_8584,N_8436);
or U8689 (N_8689,N_8444,N_8541);
or U8690 (N_8690,N_8521,N_8513);
or U8691 (N_8691,N_8583,N_8503);
nand U8692 (N_8692,N_8537,N_8451);
and U8693 (N_8693,N_8568,N_8552);
xor U8694 (N_8694,N_8416,N_8422);
or U8695 (N_8695,N_8528,N_8520);
xor U8696 (N_8696,N_8566,N_8517);
xor U8697 (N_8697,N_8482,N_8415);
xnor U8698 (N_8698,N_8461,N_8592);
nand U8699 (N_8699,N_8495,N_8437);
nor U8700 (N_8700,N_8402,N_8523);
nand U8701 (N_8701,N_8499,N_8435);
nor U8702 (N_8702,N_8562,N_8555);
xnor U8703 (N_8703,N_8411,N_8451);
xor U8704 (N_8704,N_8507,N_8553);
nand U8705 (N_8705,N_8547,N_8477);
nand U8706 (N_8706,N_8545,N_8468);
or U8707 (N_8707,N_8579,N_8580);
xor U8708 (N_8708,N_8437,N_8499);
nand U8709 (N_8709,N_8573,N_8436);
xnor U8710 (N_8710,N_8534,N_8554);
nand U8711 (N_8711,N_8411,N_8477);
and U8712 (N_8712,N_8527,N_8458);
xor U8713 (N_8713,N_8596,N_8494);
and U8714 (N_8714,N_8539,N_8413);
and U8715 (N_8715,N_8472,N_8413);
xor U8716 (N_8716,N_8473,N_8470);
xnor U8717 (N_8717,N_8487,N_8566);
xnor U8718 (N_8718,N_8522,N_8559);
xnor U8719 (N_8719,N_8497,N_8480);
and U8720 (N_8720,N_8568,N_8434);
nor U8721 (N_8721,N_8571,N_8414);
nand U8722 (N_8722,N_8568,N_8419);
nand U8723 (N_8723,N_8546,N_8501);
nor U8724 (N_8724,N_8504,N_8412);
nand U8725 (N_8725,N_8548,N_8534);
or U8726 (N_8726,N_8588,N_8551);
xor U8727 (N_8727,N_8498,N_8596);
or U8728 (N_8728,N_8486,N_8587);
nand U8729 (N_8729,N_8497,N_8404);
xor U8730 (N_8730,N_8539,N_8478);
nand U8731 (N_8731,N_8566,N_8588);
nand U8732 (N_8732,N_8417,N_8423);
and U8733 (N_8733,N_8519,N_8440);
or U8734 (N_8734,N_8552,N_8537);
xor U8735 (N_8735,N_8502,N_8408);
nor U8736 (N_8736,N_8508,N_8535);
nand U8737 (N_8737,N_8487,N_8461);
or U8738 (N_8738,N_8567,N_8491);
and U8739 (N_8739,N_8493,N_8527);
and U8740 (N_8740,N_8483,N_8571);
and U8741 (N_8741,N_8587,N_8457);
xnor U8742 (N_8742,N_8457,N_8504);
nor U8743 (N_8743,N_8588,N_8445);
nand U8744 (N_8744,N_8435,N_8578);
nand U8745 (N_8745,N_8485,N_8459);
and U8746 (N_8746,N_8430,N_8497);
and U8747 (N_8747,N_8590,N_8557);
and U8748 (N_8748,N_8458,N_8529);
and U8749 (N_8749,N_8597,N_8495);
and U8750 (N_8750,N_8503,N_8466);
xor U8751 (N_8751,N_8533,N_8592);
and U8752 (N_8752,N_8400,N_8455);
or U8753 (N_8753,N_8497,N_8597);
nor U8754 (N_8754,N_8427,N_8502);
nor U8755 (N_8755,N_8529,N_8420);
xor U8756 (N_8756,N_8436,N_8458);
or U8757 (N_8757,N_8566,N_8533);
and U8758 (N_8758,N_8471,N_8473);
nor U8759 (N_8759,N_8445,N_8524);
nor U8760 (N_8760,N_8474,N_8572);
nor U8761 (N_8761,N_8570,N_8592);
nor U8762 (N_8762,N_8405,N_8529);
and U8763 (N_8763,N_8536,N_8417);
or U8764 (N_8764,N_8425,N_8471);
nand U8765 (N_8765,N_8458,N_8500);
xnor U8766 (N_8766,N_8448,N_8529);
nor U8767 (N_8767,N_8544,N_8518);
or U8768 (N_8768,N_8415,N_8449);
xnor U8769 (N_8769,N_8428,N_8439);
nand U8770 (N_8770,N_8406,N_8470);
and U8771 (N_8771,N_8514,N_8424);
nand U8772 (N_8772,N_8504,N_8467);
and U8773 (N_8773,N_8525,N_8559);
nor U8774 (N_8774,N_8519,N_8564);
or U8775 (N_8775,N_8448,N_8524);
xor U8776 (N_8776,N_8460,N_8539);
and U8777 (N_8777,N_8566,N_8401);
and U8778 (N_8778,N_8546,N_8598);
or U8779 (N_8779,N_8414,N_8559);
nor U8780 (N_8780,N_8542,N_8482);
or U8781 (N_8781,N_8515,N_8471);
xor U8782 (N_8782,N_8536,N_8405);
nor U8783 (N_8783,N_8598,N_8564);
xnor U8784 (N_8784,N_8526,N_8541);
or U8785 (N_8785,N_8544,N_8562);
nand U8786 (N_8786,N_8493,N_8455);
or U8787 (N_8787,N_8517,N_8411);
and U8788 (N_8788,N_8509,N_8581);
xnor U8789 (N_8789,N_8597,N_8505);
and U8790 (N_8790,N_8413,N_8419);
or U8791 (N_8791,N_8403,N_8539);
nor U8792 (N_8792,N_8437,N_8405);
xnor U8793 (N_8793,N_8409,N_8577);
nand U8794 (N_8794,N_8529,N_8488);
and U8795 (N_8795,N_8560,N_8475);
and U8796 (N_8796,N_8518,N_8409);
and U8797 (N_8797,N_8437,N_8598);
nor U8798 (N_8798,N_8409,N_8441);
nor U8799 (N_8799,N_8415,N_8423);
or U8800 (N_8800,N_8707,N_8774);
and U8801 (N_8801,N_8659,N_8605);
or U8802 (N_8802,N_8777,N_8733);
xnor U8803 (N_8803,N_8682,N_8652);
nand U8804 (N_8804,N_8677,N_8622);
xnor U8805 (N_8805,N_8785,N_8759);
nor U8806 (N_8806,N_8726,N_8630);
xnor U8807 (N_8807,N_8765,N_8638);
nor U8808 (N_8808,N_8668,N_8639);
nor U8809 (N_8809,N_8631,N_8650);
and U8810 (N_8810,N_8629,N_8767);
xnor U8811 (N_8811,N_8715,N_8628);
nor U8812 (N_8812,N_8753,N_8794);
nand U8813 (N_8813,N_8646,N_8713);
xor U8814 (N_8814,N_8618,N_8632);
nand U8815 (N_8815,N_8776,N_8613);
and U8816 (N_8816,N_8704,N_8658);
and U8817 (N_8817,N_8625,N_8661);
and U8818 (N_8818,N_8616,N_8705);
and U8819 (N_8819,N_8731,N_8708);
nand U8820 (N_8820,N_8697,N_8643);
nor U8821 (N_8821,N_8608,N_8626);
or U8822 (N_8822,N_8790,N_8745);
nand U8823 (N_8823,N_8746,N_8734);
xor U8824 (N_8824,N_8645,N_8681);
nand U8825 (N_8825,N_8676,N_8662);
or U8826 (N_8826,N_8684,N_8665);
nor U8827 (N_8827,N_8673,N_8700);
xor U8828 (N_8828,N_8642,N_8620);
or U8829 (N_8829,N_8671,N_8792);
nor U8830 (N_8830,N_8768,N_8739);
or U8831 (N_8831,N_8685,N_8761);
nand U8832 (N_8832,N_8722,N_8773);
nor U8833 (N_8833,N_8667,N_8771);
xnor U8834 (N_8834,N_8669,N_8600);
and U8835 (N_8835,N_8711,N_8649);
nand U8836 (N_8836,N_8793,N_8747);
or U8837 (N_8837,N_8751,N_8604);
xor U8838 (N_8838,N_8760,N_8772);
nand U8839 (N_8839,N_8743,N_8607);
nand U8840 (N_8840,N_8648,N_8735);
nand U8841 (N_8841,N_8758,N_8742);
nor U8842 (N_8842,N_8691,N_8741);
nand U8843 (N_8843,N_8627,N_8687);
and U8844 (N_8844,N_8728,N_8709);
or U8845 (N_8845,N_8624,N_8752);
xor U8846 (N_8846,N_8729,N_8783);
xor U8847 (N_8847,N_8717,N_8663);
nor U8848 (N_8848,N_8779,N_8688);
xor U8849 (N_8849,N_8797,N_8634);
or U8850 (N_8850,N_8699,N_8701);
xnor U8851 (N_8851,N_8763,N_8764);
and U8852 (N_8852,N_8689,N_8748);
nor U8853 (N_8853,N_8617,N_8621);
or U8854 (N_8854,N_8635,N_8703);
xnor U8855 (N_8855,N_8675,N_8791);
and U8856 (N_8856,N_8723,N_8798);
xnor U8857 (N_8857,N_8784,N_8611);
nand U8858 (N_8858,N_8660,N_8712);
nand U8859 (N_8859,N_8690,N_8683);
nand U8860 (N_8860,N_8637,N_8636);
xor U8861 (N_8861,N_8795,N_8680);
nand U8862 (N_8862,N_8615,N_8702);
and U8863 (N_8863,N_8653,N_8692);
and U8864 (N_8864,N_8640,N_8606);
or U8865 (N_8865,N_8725,N_8782);
xor U8866 (N_8866,N_8651,N_8756);
nand U8867 (N_8867,N_8738,N_8693);
and U8868 (N_8868,N_8786,N_8749);
xnor U8869 (N_8869,N_8789,N_8770);
xnor U8870 (N_8870,N_8720,N_8737);
nor U8871 (N_8871,N_8672,N_8710);
nor U8872 (N_8872,N_8778,N_8647);
and U8873 (N_8873,N_8740,N_8769);
xor U8874 (N_8874,N_8766,N_8623);
xnor U8875 (N_8875,N_8619,N_8657);
xnor U8876 (N_8876,N_8670,N_8732);
nor U8877 (N_8877,N_8655,N_8609);
or U8878 (N_8878,N_8614,N_8679);
and U8879 (N_8879,N_8744,N_8666);
nand U8880 (N_8880,N_8602,N_8654);
nand U8881 (N_8881,N_8674,N_8721);
xnor U8882 (N_8882,N_8694,N_8762);
nand U8883 (N_8883,N_8781,N_8601);
nand U8884 (N_8884,N_8787,N_8633);
and U8885 (N_8885,N_8750,N_8612);
nor U8886 (N_8886,N_8780,N_8754);
nand U8887 (N_8887,N_8714,N_8719);
xor U8888 (N_8888,N_8788,N_8796);
or U8889 (N_8889,N_8644,N_8736);
xor U8890 (N_8890,N_8724,N_8695);
or U8891 (N_8891,N_8664,N_8678);
nor U8892 (N_8892,N_8706,N_8641);
xor U8893 (N_8893,N_8775,N_8656);
or U8894 (N_8894,N_8730,N_8757);
and U8895 (N_8895,N_8755,N_8718);
or U8896 (N_8896,N_8696,N_8727);
and U8897 (N_8897,N_8603,N_8686);
nand U8898 (N_8898,N_8610,N_8716);
and U8899 (N_8899,N_8799,N_8698);
nand U8900 (N_8900,N_8614,N_8700);
nand U8901 (N_8901,N_8619,N_8763);
or U8902 (N_8902,N_8798,N_8685);
nor U8903 (N_8903,N_8782,N_8785);
and U8904 (N_8904,N_8680,N_8764);
and U8905 (N_8905,N_8682,N_8681);
nand U8906 (N_8906,N_8750,N_8786);
nand U8907 (N_8907,N_8612,N_8704);
nor U8908 (N_8908,N_8799,N_8768);
nor U8909 (N_8909,N_8678,N_8762);
or U8910 (N_8910,N_8790,N_8661);
xnor U8911 (N_8911,N_8785,N_8734);
or U8912 (N_8912,N_8650,N_8645);
nand U8913 (N_8913,N_8614,N_8793);
or U8914 (N_8914,N_8651,N_8661);
or U8915 (N_8915,N_8757,N_8705);
nand U8916 (N_8916,N_8757,N_8738);
xnor U8917 (N_8917,N_8734,N_8765);
xor U8918 (N_8918,N_8784,N_8723);
xor U8919 (N_8919,N_8671,N_8786);
nand U8920 (N_8920,N_8796,N_8600);
and U8921 (N_8921,N_8725,N_8649);
or U8922 (N_8922,N_8769,N_8659);
nor U8923 (N_8923,N_8677,N_8629);
nor U8924 (N_8924,N_8612,N_8628);
xnor U8925 (N_8925,N_8604,N_8646);
xor U8926 (N_8926,N_8679,N_8670);
xor U8927 (N_8927,N_8700,N_8610);
nor U8928 (N_8928,N_8617,N_8773);
nand U8929 (N_8929,N_8778,N_8766);
xnor U8930 (N_8930,N_8636,N_8778);
nor U8931 (N_8931,N_8632,N_8713);
xnor U8932 (N_8932,N_8634,N_8780);
nand U8933 (N_8933,N_8624,N_8780);
xor U8934 (N_8934,N_8644,N_8647);
and U8935 (N_8935,N_8786,N_8748);
nor U8936 (N_8936,N_8781,N_8683);
nand U8937 (N_8937,N_8749,N_8637);
or U8938 (N_8938,N_8652,N_8726);
or U8939 (N_8939,N_8783,N_8636);
nor U8940 (N_8940,N_8776,N_8700);
and U8941 (N_8941,N_8666,N_8796);
and U8942 (N_8942,N_8612,N_8792);
nor U8943 (N_8943,N_8740,N_8692);
or U8944 (N_8944,N_8630,N_8602);
xnor U8945 (N_8945,N_8718,N_8633);
or U8946 (N_8946,N_8681,N_8629);
or U8947 (N_8947,N_8682,N_8615);
xor U8948 (N_8948,N_8647,N_8673);
nand U8949 (N_8949,N_8705,N_8752);
and U8950 (N_8950,N_8788,N_8620);
xor U8951 (N_8951,N_8767,N_8603);
nor U8952 (N_8952,N_8611,N_8666);
nor U8953 (N_8953,N_8659,N_8691);
nand U8954 (N_8954,N_8620,N_8688);
xnor U8955 (N_8955,N_8635,N_8620);
xor U8956 (N_8956,N_8661,N_8628);
or U8957 (N_8957,N_8700,N_8668);
nor U8958 (N_8958,N_8655,N_8691);
xnor U8959 (N_8959,N_8735,N_8728);
nor U8960 (N_8960,N_8608,N_8770);
xnor U8961 (N_8961,N_8682,N_8767);
and U8962 (N_8962,N_8771,N_8711);
or U8963 (N_8963,N_8651,N_8709);
and U8964 (N_8964,N_8719,N_8789);
nor U8965 (N_8965,N_8621,N_8772);
nand U8966 (N_8966,N_8758,N_8720);
nand U8967 (N_8967,N_8690,N_8658);
nand U8968 (N_8968,N_8752,N_8762);
and U8969 (N_8969,N_8762,N_8723);
or U8970 (N_8970,N_8639,N_8704);
xor U8971 (N_8971,N_8706,N_8623);
or U8972 (N_8972,N_8742,N_8683);
and U8973 (N_8973,N_8735,N_8745);
or U8974 (N_8974,N_8647,N_8797);
or U8975 (N_8975,N_8784,N_8624);
and U8976 (N_8976,N_8720,N_8662);
xnor U8977 (N_8977,N_8642,N_8794);
nor U8978 (N_8978,N_8635,N_8735);
xnor U8979 (N_8979,N_8763,N_8606);
or U8980 (N_8980,N_8656,N_8784);
xnor U8981 (N_8981,N_8692,N_8651);
nand U8982 (N_8982,N_8785,N_8698);
nor U8983 (N_8983,N_8613,N_8601);
xor U8984 (N_8984,N_8618,N_8608);
or U8985 (N_8985,N_8699,N_8717);
and U8986 (N_8986,N_8748,N_8706);
or U8987 (N_8987,N_8748,N_8608);
nor U8988 (N_8988,N_8615,N_8706);
or U8989 (N_8989,N_8631,N_8768);
xnor U8990 (N_8990,N_8602,N_8604);
and U8991 (N_8991,N_8759,N_8732);
nand U8992 (N_8992,N_8750,N_8648);
xor U8993 (N_8993,N_8685,N_8691);
or U8994 (N_8994,N_8647,N_8630);
nor U8995 (N_8995,N_8763,N_8780);
nor U8996 (N_8996,N_8744,N_8785);
nand U8997 (N_8997,N_8679,N_8757);
nor U8998 (N_8998,N_8679,N_8638);
xor U8999 (N_8999,N_8719,N_8793);
and U9000 (N_9000,N_8858,N_8890);
or U9001 (N_9001,N_8830,N_8979);
xnor U9002 (N_9002,N_8859,N_8918);
and U9003 (N_9003,N_8849,N_8880);
xnor U9004 (N_9004,N_8927,N_8995);
nand U9005 (N_9005,N_8833,N_8982);
nor U9006 (N_9006,N_8812,N_8990);
or U9007 (N_9007,N_8948,N_8856);
xnor U9008 (N_9008,N_8840,N_8896);
xor U9009 (N_9009,N_8884,N_8981);
and U9010 (N_9010,N_8914,N_8824);
nand U9011 (N_9011,N_8956,N_8816);
or U9012 (N_9012,N_8877,N_8898);
nor U9013 (N_9013,N_8901,N_8854);
xor U9014 (N_9014,N_8944,N_8800);
or U9015 (N_9015,N_8875,N_8998);
nor U9016 (N_9016,N_8984,N_8946);
nand U9017 (N_9017,N_8966,N_8973);
or U9018 (N_9018,N_8878,N_8822);
and U9019 (N_9019,N_8953,N_8845);
and U9020 (N_9020,N_8920,N_8974);
xnor U9021 (N_9021,N_8819,N_8969);
or U9022 (N_9022,N_8806,N_8965);
nor U9023 (N_9023,N_8980,N_8887);
xor U9024 (N_9024,N_8831,N_8915);
or U9025 (N_9025,N_8983,N_8860);
nor U9026 (N_9026,N_8805,N_8975);
and U9027 (N_9027,N_8910,N_8809);
xor U9028 (N_9028,N_8818,N_8913);
and U9029 (N_9029,N_8971,N_8977);
and U9030 (N_9030,N_8852,N_8931);
nor U9031 (N_9031,N_8850,N_8970);
xnor U9032 (N_9032,N_8954,N_8874);
and U9033 (N_9033,N_8903,N_8814);
xnor U9034 (N_9034,N_8879,N_8959);
and U9035 (N_9035,N_8897,N_8928);
nor U9036 (N_9036,N_8976,N_8817);
xor U9037 (N_9037,N_8828,N_8941);
or U9038 (N_9038,N_8904,N_8855);
xor U9039 (N_9039,N_8912,N_8906);
xor U9040 (N_9040,N_8865,N_8943);
or U9041 (N_9041,N_8821,N_8844);
xnor U9042 (N_9042,N_8846,N_8967);
nor U9043 (N_9043,N_8803,N_8909);
nor U9044 (N_9044,N_8908,N_8924);
or U9045 (N_9045,N_8891,N_8911);
or U9046 (N_9046,N_8992,N_8815);
nand U9047 (N_9047,N_8832,N_8994);
and U9048 (N_9048,N_8950,N_8867);
and U9049 (N_9049,N_8861,N_8945);
or U9050 (N_9050,N_8963,N_8837);
nand U9051 (N_9051,N_8813,N_8864);
xnor U9052 (N_9052,N_8876,N_8881);
nor U9053 (N_9053,N_8820,N_8999);
nor U9054 (N_9054,N_8951,N_8839);
nand U9055 (N_9055,N_8873,N_8936);
nor U9056 (N_9056,N_8826,N_8989);
xor U9057 (N_9057,N_8968,N_8929);
xor U9058 (N_9058,N_8905,N_8834);
nand U9059 (N_9059,N_8886,N_8802);
nor U9060 (N_9060,N_8848,N_8957);
nand U9061 (N_9061,N_8825,N_8986);
or U9062 (N_9062,N_8917,N_8838);
nor U9063 (N_9063,N_8921,N_8811);
nand U9064 (N_9064,N_8960,N_8807);
nand U9065 (N_9065,N_8853,N_8902);
nand U9066 (N_9066,N_8894,N_8949);
nor U9067 (N_9067,N_8939,N_8985);
nand U9068 (N_9068,N_8841,N_8938);
nand U9069 (N_9069,N_8892,N_8857);
xor U9070 (N_9070,N_8978,N_8862);
nor U9071 (N_9071,N_8997,N_8958);
nor U9072 (N_9072,N_8863,N_8827);
and U9073 (N_9073,N_8810,N_8882);
xor U9074 (N_9074,N_8842,N_8889);
or U9075 (N_9075,N_8932,N_8919);
nand U9076 (N_9076,N_8930,N_8829);
or U9077 (N_9077,N_8934,N_8972);
and U9078 (N_9078,N_8993,N_8899);
nor U9079 (N_9079,N_8942,N_8962);
xor U9080 (N_9080,N_8922,N_8869);
or U9081 (N_9081,N_8916,N_8900);
or U9082 (N_9082,N_8988,N_8835);
nand U9083 (N_9083,N_8893,N_8925);
nand U9084 (N_9084,N_8952,N_8868);
xnor U9085 (N_9085,N_8801,N_8937);
and U9086 (N_9086,N_8885,N_8866);
xnor U9087 (N_9087,N_8964,N_8895);
and U9088 (N_9088,N_8935,N_8947);
or U9089 (N_9089,N_8872,N_8870);
nand U9090 (N_9090,N_8961,N_8823);
nor U9091 (N_9091,N_8836,N_8923);
nand U9092 (N_9092,N_8888,N_8996);
nor U9093 (N_9093,N_8883,N_8926);
and U9094 (N_9094,N_8843,N_8847);
or U9095 (N_9095,N_8955,N_8907);
nor U9096 (N_9096,N_8933,N_8987);
or U9097 (N_9097,N_8991,N_8851);
and U9098 (N_9098,N_8871,N_8804);
and U9099 (N_9099,N_8808,N_8940);
or U9100 (N_9100,N_8961,N_8854);
or U9101 (N_9101,N_8895,N_8941);
nand U9102 (N_9102,N_8974,N_8913);
and U9103 (N_9103,N_8987,N_8962);
or U9104 (N_9104,N_8852,N_8912);
nand U9105 (N_9105,N_8979,N_8840);
xor U9106 (N_9106,N_8938,N_8931);
nor U9107 (N_9107,N_8993,N_8931);
xor U9108 (N_9108,N_8837,N_8819);
xnor U9109 (N_9109,N_8903,N_8906);
and U9110 (N_9110,N_8820,N_8864);
or U9111 (N_9111,N_8833,N_8964);
and U9112 (N_9112,N_8914,N_8872);
and U9113 (N_9113,N_8967,N_8974);
or U9114 (N_9114,N_8996,N_8954);
nand U9115 (N_9115,N_8980,N_8851);
nand U9116 (N_9116,N_8851,N_8861);
or U9117 (N_9117,N_8805,N_8828);
xnor U9118 (N_9118,N_8806,N_8911);
nor U9119 (N_9119,N_8877,N_8981);
and U9120 (N_9120,N_8806,N_8866);
nor U9121 (N_9121,N_8848,N_8883);
and U9122 (N_9122,N_8885,N_8908);
xor U9123 (N_9123,N_8903,N_8851);
and U9124 (N_9124,N_8812,N_8923);
nand U9125 (N_9125,N_8901,N_8860);
or U9126 (N_9126,N_8967,N_8952);
nand U9127 (N_9127,N_8814,N_8928);
or U9128 (N_9128,N_8829,N_8890);
nor U9129 (N_9129,N_8853,N_8891);
or U9130 (N_9130,N_8942,N_8813);
or U9131 (N_9131,N_8892,N_8984);
and U9132 (N_9132,N_8961,N_8913);
nor U9133 (N_9133,N_8899,N_8893);
nor U9134 (N_9134,N_8898,N_8815);
nor U9135 (N_9135,N_8895,N_8988);
and U9136 (N_9136,N_8842,N_8986);
and U9137 (N_9137,N_8850,N_8917);
nor U9138 (N_9138,N_8828,N_8950);
xnor U9139 (N_9139,N_8920,N_8928);
and U9140 (N_9140,N_8960,N_8930);
nor U9141 (N_9141,N_8950,N_8847);
xor U9142 (N_9142,N_8878,N_8980);
or U9143 (N_9143,N_8959,N_8966);
nor U9144 (N_9144,N_8991,N_8848);
and U9145 (N_9145,N_8996,N_8922);
nand U9146 (N_9146,N_8971,N_8844);
nor U9147 (N_9147,N_8821,N_8957);
and U9148 (N_9148,N_8900,N_8821);
xnor U9149 (N_9149,N_8967,N_8937);
xnor U9150 (N_9150,N_8871,N_8813);
and U9151 (N_9151,N_8878,N_8927);
and U9152 (N_9152,N_8909,N_8981);
or U9153 (N_9153,N_8909,N_8894);
and U9154 (N_9154,N_8999,N_8945);
and U9155 (N_9155,N_8989,N_8925);
nand U9156 (N_9156,N_8904,N_8999);
nor U9157 (N_9157,N_8935,N_8985);
xor U9158 (N_9158,N_8902,N_8942);
xnor U9159 (N_9159,N_8949,N_8904);
nor U9160 (N_9160,N_8920,N_8987);
nor U9161 (N_9161,N_8829,N_8939);
or U9162 (N_9162,N_8863,N_8858);
and U9163 (N_9163,N_8896,N_8975);
or U9164 (N_9164,N_8944,N_8846);
nand U9165 (N_9165,N_8995,N_8802);
xor U9166 (N_9166,N_8944,N_8913);
nor U9167 (N_9167,N_8936,N_8810);
nand U9168 (N_9168,N_8959,N_8895);
or U9169 (N_9169,N_8810,N_8927);
and U9170 (N_9170,N_8989,N_8877);
nand U9171 (N_9171,N_8901,N_8973);
nor U9172 (N_9172,N_8834,N_8977);
nand U9173 (N_9173,N_8935,N_8895);
nor U9174 (N_9174,N_8966,N_8910);
or U9175 (N_9175,N_8988,N_8842);
or U9176 (N_9176,N_8916,N_8830);
and U9177 (N_9177,N_8865,N_8846);
or U9178 (N_9178,N_8832,N_8820);
and U9179 (N_9179,N_8834,N_8851);
nor U9180 (N_9180,N_8806,N_8878);
nor U9181 (N_9181,N_8914,N_8848);
and U9182 (N_9182,N_8822,N_8883);
or U9183 (N_9183,N_8806,N_8971);
and U9184 (N_9184,N_8856,N_8907);
nand U9185 (N_9185,N_8991,N_8821);
nor U9186 (N_9186,N_8800,N_8885);
xnor U9187 (N_9187,N_8863,N_8959);
and U9188 (N_9188,N_8957,N_8985);
nor U9189 (N_9189,N_8951,N_8960);
nor U9190 (N_9190,N_8908,N_8982);
nand U9191 (N_9191,N_8939,N_8867);
nand U9192 (N_9192,N_8875,N_8823);
and U9193 (N_9193,N_8899,N_8917);
xor U9194 (N_9194,N_8896,N_8869);
and U9195 (N_9195,N_8814,N_8945);
nor U9196 (N_9196,N_8862,N_8919);
xnor U9197 (N_9197,N_8965,N_8966);
xnor U9198 (N_9198,N_8905,N_8985);
or U9199 (N_9199,N_8960,N_8974);
or U9200 (N_9200,N_9033,N_9144);
nand U9201 (N_9201,N_9092,N_9022);
and U9202 (N_9202,N_9163,N_9130);
or U9203 (N_9203,N_9042,N_9061);
xnor U9204 (N_9204,N_9174,N_9002);
and U9205 (N_9205,N_9156,N_9068);
nor U9206 (N_9206,N_9082,N_9176);
or U9207 (N_9207,N_9106,N_9089);
xnor U9208 (N_9208,N_9105,N_9003);
xnor U9209 (N_9209,N_9189,N_9053);
xor U9210 (N_9210,N_9087,N_9031);
or U9211 (N_9211,N_9046,N_9147);
or U9212 (N_9212,N_9184,N_9050);
or U9213 (N_9213,N_9039,N_9146);
or U9214 (N_9214,N_9152,N_9102);
nor U9215 (N_9215,N_9067,N_9186);
and U9216 (N_9216,N_9076,N_9109);
nand U9217 (N_9217,N_9014,N_9045);
xnor U9218 (N_9218,N_9162,N_9027);
nor U9219 (N_9219,N_9173,N_9141);
nand U9220 (N_9220,N_9083,N_9063);
xor U9221 (N_9221,N_9161,N_9080);
or U9222 (N_9222,N_9058,N_9047);
nor U9223 (N_9223,N_9167,N_9123);
or U9224 (N_9224,N_9037,N_9016);
or U9225 (N_9225,N_9006,N_9113);
or U9226 (N_9226,N_9172,N_9137);
nand U9227 (N_9227,N_9054,N_9199);
xnor U9228 (N_9228,N_9023,N_9028);
and U9229 (N_9229,N_9185,N_9029);
nor U9230 (N_9230,N_9191,N_9049);
nor U9231 (N_9231,N_9011,N_9094);
nand U9232 (N_9232,N_9013,N_9090);
or U9233 (N_9233,N_9060,N_9164);
nor U9234 (N_9234,N_9085,N_9040);
and U9235 (N_9235,N_9001,N_9120);
nor U9236 (N_9236,N_9078,N_9150);
and U9237 (N_9237,N_9032,N_9066);
nor U9238 (N_9238,N_9157,N_9151);
nand U9239 (N_9239,N_9115,N_9128);
xor U9240 (N_9240,N_9038,N_9117);
xnor U9241 (N_9241,N_9129,N_9169);
nand U9242 (N_9242,N_9035,N_9025);
xor U9243 (N_9243,N_9114,N_9072);
nor U9244 (N_9244,N_9136,N_9148);
or U9245 (N_9245,N_9075,N_9119);
and U9246 (N_9246,N_9064,N_9183);
or U9247 (N_9247,N_9097,N_9197);
nor U9248 (N_9248,N_9194,N_9187);
xor U9249 (N_9249,N_9122,N_9099);
nor U9250 (N_9250,N_9056,N_9166);
nor U9251 (N_9251,N_9158,N_9101);
xor U9252 (N_9252,N_9112,N_9143);
or U9253 (N_9253,N_9175,N_9015);
nand U9254 (N_9254,N_9160,N_9057);
and U9255 (N_9255,N_9052,N_9145);
nand U9256 (N_9256,N_9134,N_9103);
nand U9257 (N_9257,N_9195,N_9008);
nand U9258 (N_9258,N_9104,N_9000);
xor U9259 (N_9259,N_9084,N_9044);
or U9260 (N_9260,N_9073,N_9181);
xor U9261 (N_9261,N_9138,N_9041);
or U9262 (N_9262,N_9024,N_9121);
xor U9263 (N_9263,N_9048,N_9100);
or U9264 (N_9264,N_9124,N_9065);
xor U9265 (N_9265,N_9142,N_9055);
nor U9266 (N_9266,N_9132,N_9180);
nor U9267 (N_9267,N_9153,N_9098);
and U9268 (N_9268,N_9093,N_9071);
or U9269 (N_9269,N_9192,N_9178);
xnor U9270 (N_9270,N_9140,N_9111);
xnor U9271 (N_9271,N_9179,N_9107);
nor U9272 (N_9272,N_9043,N_9170);
or U9273 (N_9273,N_9086,N_9118);
and U9274 (N_9274,N_9020,N_9133);
xnor U9275 (N_9275,N_9182,N_9159);
nor U9276 (N_9276,N_9193,N_9018);
and U9277 (N_9277,N_9004,N_9110);
nand U9278 (N_9278,N_9081,N_9139);
nand U9279 (N_9279,N_9009,N_9088);
nor U9280 (N_9280,N_9188,N_9062);
and U9281 (N_9281,N_9171,N_9127);
xnor U9282 (N_9282,N_9095,N_9125);
xor U9283 (N_9283,N_9165,N_9012);
nor U9284 (N_9284,N_9108,N_9135);
nor U9285 (N_9285,N_9154,N_9096);
or U9286 (N_9286,N_9196,N_9190);
or U9287 (N_9287,N_9051,N_9059);
nor U9288 (N_9288,N_9198,N_9074);
xor U9289 (N_9289,N_9168,N_9026);
nor U9290 (N_9290,N_9126,N_9079);
or U9291 (N_9291,N_9019,N_9069);
nor U9292 (N_9292,N_9077,N_9021);
xor U9293 (N_9293,N_9005,N_9091);
nor U9294 (N_9294,N_9030,N_9155);
nor U9295 (N_9295,N_9116,N_9177);
nand U9296 (N_9296,N_9034,N_9036);
and U9297 (N_9297,N_9010,N_9131);
or U9298 (N_9298,N_9149,N_9070);
nand U9299 (N_9299,N_9017,N_9007);
and U9300 (N_9300,N_9109,N_9197);
or U9301 (N_9301,N_9071,N_9118);
xnor U9302 (N_9302,N_9076,N_9057);
xor U9303 (N_9303,N_9129,N_9193);
and U9304 (N_9304,N_9152,N_9176);
nor U9305 (N_9305,N_9130,N_9133);
and U9306 (N_9306,N_9037,N_9033);
nand U9307 (N_9307,N_9081,N_9050);
and U9308 (N_9308,N_9158,N_9030);
or U9309 (N_9309,N_9143,N_9125);
nor U9310 (N_9310,N_9124,N_9191);
xnor U9311 (N_9311,N_9062,N_9091);
xor U9312 (N_9312,N_9197,N_9174);
xor U9313 (N_9313,N_9050,N_9020);
xor U9314 (N_9314,N_9046,N_9141);
nor U9315 (N_9315,N_9110,N_9050);
or U9316 (N_9316,N_9142,N_9049);
nor U9317 (N_9317,N_9107,N_9102);
and U9318 (N_9318,N_9071,N_9144);
xnor U9319 (N_9319,N_9089,N_9100);
xnor U9320 (N_9320,N_9059,N_9124);
xor U9321 (N_9321,N_9012,N_9123);
nand U9322 (N_9322,N_9133,N_9177);
xor U9323 (N_9323,N_9016,N_9102);
or U9324 (N_9324,N_9036,N_9038);
nand U9325 (N_9325,N_9008,N_9062);
and U9326 (N_9326,N_9033,N_9065);
and U9327 (N_9327,N_9016,N_9076);
or U9328 (N_9328,N_9006,N_9040);
nand U9329 (N_9329,N_9168,N_9174);
xor U9330 (N_9330,N_9187,N_9038);
xnor U9331 (N_9331,N_9095,N_9026);
or U9332 (N_9332,N_9167,N_9133);
and U9333 (N_9333,N_9051,N_9027);
or U9334 (N_9334,N_9054,N_9180);
and U9335 (N_9335,N_9010,N_9008);
and U9336 (N_9336,N_9134,N_9157);
xor U9337 (N_9337,N_9002,N_9088);
nand U9338 (N_9338,N_9028,N_9141);
nand U9339 (N_9339,N_9060,N_9008);
or U9340 (N_9340,N_9101,N_9153);
xnor U9341 (N_9341,N_9177,N_9095);
or U9342 (N_9342,N_9105,N_9053);
nor U9343 (N_9343,N_9114,N_9067);
and U9344 (N_9344,N_9085,N_9084);
and U9345 (N_9345,N_9007,N_9013);
xnor U9346 (N_9346,N_9191,N_9021);
and U9347 (N_9347,N_9028,N_9123);
nand U9348 (N_9348,N_9139,N_9000);
nand U9349 (N_9349,N_9132,N_9103);
and U9350 (N_9350,N_9161,N_9101);
or U9351 (N_9351,N_9019,N_9030);
or U9352 (N_9352,N_9021,N_9007);
or U9353 (N_9353,N_9071,N_9127);
nor U9354 (N_9354,N_9081,N_9051);
xor U9355 (N_9355,N_9071,N_9113);
nor U9356 (N_9356,N_9176,N_9146);
nor U9357 (N_9357,N_9005,N_9152);
and U9358 (N_9358,N_9130,N_9019);
and U9359 (N_9359,N_9094,N_9139);
and U9360 (N_9360,N_9001,N_9054);
nor U9361 (N_9361,N_9005,N_9129);
xnor U9362 (N_9362,N_9026,N_9023);
xnor U9363 (N_9363,N_9056,N_9185);
nor U9364 (N_9364,N_9159,N_9064);
nand U9365 (N_9365,N_9079,N_9088);
nand U9366 (N_9366,N_9064,N_9182);
xnor U9367 (N_9367,N_9043,N_9006);
nand U9368 (N_9368,N_9015,N_9157);
nand U9369 (N_9369,N_9099,N_9128);
and U9370 (N_9370,N_9081,N_9003);
or U9371 (N_9371,N_9126,N_9180);
xor U9372 (N_9372,N_9176,N_9129);
or U9373 (N_9373,N_9183,N_9020);
xor U9374 (N_9374,N_9016,N_9071);
nand U9375 (N_9375,N_9072,N_9167);
xnor U9376 (N_9376,N_9169,N_9034);
nor U9377 (N_9377,N_9150,N_9195);
and U9378 (N_9378,N_9169,N_9114);
nand U9379 (N_9379,N_9118,N_9079);
or U9380 (N_9380,N_9173,N_9191);
and U9381 (N_9381,N_9084,N_9014);
or U9382 (N_9382,N_9166,N_9168);
nand U9383 (N_9383,N_9150,N_9183);
nor U9384 (N_9384,N_9146,N_9026);
xor U9385 (N_9385,N_9111,N_9018);
nor U9386 (N_9386,N_9057,N_9111);
xor U9387 (N_9387,N_9110,N_9076);
nand U9388 (N_9388,N_9153,N_9163);
or U9389 (N_9389,N_9166,N_9140);
xnor U9390 (N_9390,N_9176,N_9133);
nor U9391 (N_9391,N_9190,N_9037);
and U9392 (N_9392,N_9114,N_9016);
nand U9393 (N_9393,N_9088,N_9077);
and U9394 (N_9394,N_9172,N_9125);
nand U9395 (N_9395,N_9041,N_9156);
nor U9396 (N_9396,N_9133,N_9188);
nand U9397 (N_9397,N_9131,N_9180);
xor U9398 (N_9398,N_9161,N_9077);
nor U9399 (N_9399,N_9165,N_9022);
nor U9400 (N_9400,N_9201,N_9280);
xnor U9401 (N_9401,N_9220,N_9230);
or U9402 (N_9402,N_9233,N_9305);
nand U9403 (N_9403,N_9269,N_9355);
xor U9404 (N_9404,N_9332,N_9366);
or U9405 (N_9405,N_9255,N_9313);
nor U9406 (N_9406,N_9397,N_9270);
and U9407 (N_9407,N_9381,N_9302);
nand U9408 (N_9408,N_9390,N_9253);
nor U9409 (N_9409,N_9227,N_9214);
xor U9410 (N_9410,N_9247,N_9337);
nor U9411 (N_9411,N_9356,N_9380);
xnor U9412 (N_9412,N_9203,N_9311);
or U9413 (N_9413,N_9234,N_9232);
nand U9414 (N_9414,N_9245,N_9238);
nor U9415 (N_9415,N_9357,N_9229);
and U9416 (N_9416,N_9271,N_9360);
and U9417 (N_9417,N_9386,N_9239);
nand U9418 (N_9418,N_9364,N_9316);
or U9419 (N_9419,N_9301,N_9263);
xnor U9420 (N_9420,N_9336,N_9249);
nor U9421 (N_9421,N_9359,N_9382);
nand U9422 (N_9422,N_9369,N_9211);
or U9423 (N_9423,N_9399,N_9254);
nand U9424 (N_9424,N_9290,N_9308);
nand U9425 (N_9425,N_9373,N_9235);
or U9426 (N_9426,N_9218,N_9210);
nand U9427 (N_9427,N_9378,N_9289);
nor U9428 (N_9428,N_9391,N_9326);
xnor U9429 (N_9429,N_9347,N_9292);
nor U9430 (N_9430,N_9307,N_9324);
and U9431 (N_9431,N_9212,N_9368);
nor U9432 (N_9432,N_9200,N_9328);
and U9433 (N_9433,N_9206,N_9228);
or U9434 (N_9434,N_9398,N_9310);
or U9435 (N_9435,N_9272,N_9246);
nor U9436 (N_9436,N_9265,N_9361);
or U9437 (N_9437,N_9330,N_9352);
nand U9438 (N_9438,N_9275,N_9259);
or U9439 (N_9439,N_9241,N_9341);
nand U9440 (N_9440,N_9348,N_9394);
and U9441 (N_9441,N_9297,N_9262);
nand U9442 (N_9442,N_9375,N_9374);
xor U9443 (N_9443,N_9251,N_9343);
xnor U9444 (N_9444,N_9379,N_9388);
xor U9445 (N_9445,N_9231,N_9358);
and U9446 (N_9446,N_9294,N_9257);
nor U9447 (N_9447,N_9282,N_9268);
and U9448 (N_9448,N_9303,N_9248);
nor U9449 (N_9449,N_9350,N_9383);
and U9450 (N_9450,N_9395,N_9365);
nand U9451 (N_9451,N_9309,N_9338);
or U9452 (N_9452,N_9258,N_9242);
or U9453 (N_9453,N_9319,N_9296);
and U9454 (N_9454,N_9276,N_9216);
xnor U9455 (N_9455,N_9340,N_9204);
xnor U9456 (N_9456,N_9312,N_9353);
nor U9457 (N_9457,N_9278,N_9277);
nand U9458 (N_9458,N_9349,N_9329);
and U9459 (N_9459,N_9215,N_9287);
or U9460 (N_9460,N_9222,N_9252);
xor U9461 (N_9461,N_9226,N_9284);
xor U9462 (N_9462,N_9260,N_9315);
xor U9463 (N_9463,N_9208,N_9376);
xor U9464 (N_9464,N_9327,N_9320);
xnor U9465 (N_9465,N_9205,N_9384);
nor U9466 (N_9466,N_9261,N_9293);
and U9467 (N_9467,N_9244,N_9371);
and U9468 (N_9468,N_9213,N_9281);
and U9469 (N_9469,N_9342,N_9331);
nor U9470 (N_9470,N_9354,N_9219);
nor U9471 (N_9471,N_9345,N_9236);
and U9472 (N_9472,N_9298,N_9240);
xor U9473 (N_9473,N_9237,N_9291);
xor U9474 (N_9474,N_9334,N_9372);
and U9475 (N_9475,N_9225,N_9267);
nor U9476 (N_9476,N_9264,N_9223);
nand U9477 (N_9477,N_9250,N_9325);
and U9478 (N_9478,N_9221,N_9243);
nor U9479 (N_9479,N_9318,N_9317);
nor U9480 (N_9480,N_9224,N_9344);
xor U9481 (N_9481,N_9266,N_9295);
xor U9482 (N_9482,N_9209,N_9362);
or U9483 (N_9483,N_9256,N_9387);
nor U9484 (N_9484,N_9202,N_9339);
nor U9485 (N_9485,N_9385,N_9333);
and U9486 (N_9486,N_9279,N_9351);
or U9487 (N_9487,N_9367,N_9363);
nand U9488 (N_9488,N_9314,N_9286);
xnor U9489 (N_9489,N_9389,N_9283);
or U9490 (N_9490,N_9370,N_9285);
and U9491 (N_9491,N_9377,N_9392);
nor U9492 (N_9492,N_9306,N_9393);
xnor U9493 (N_9493,N_9300,N_9323);
nor U9494 (N_9494,N_9207,N_9288);
nand U9495 (N_9495,N_9274,N_9346);
and U9496 (N_9496,N_9322,N_9217);
and U9497 (N_9497,N_9396,N_9321);
nor U9498 (N_9498,N_9304,N_9335);
xnor U9499 (N_9499,N_9299,N_9273);
nor U9500 (N_9500,N_9345,N_9377);
xnor U9501 (N_9501,N_9232,N_9251);
or U9502 (N_9502,N_9294,N_9360);
or U9503 (N_9503,N_9374,N_9354);
nor U9504 (N_9504,N_9298,N_9373);
and U9505 (N_9505,N_9231,N_9213);
nor U9506 (N_9506,N_9342,N_9289);
xor U9507 (N_9507,N_9315,N_9376);
nand U9508 (N_9508,N_9282,N_9284);
nand U9509 (N_9509,N_9225,N_9270);
nand U9510 (N_9510,N_9216,N_9275);
xnor U9511 (N_9511,N_9251,N_9273);
nor U9512 (N_9512,N_9338,N_9275);
xor U9513 (N_9513,N_9376,N_9351);
nor U9514 (N_9514,N_9205,N_9212);
nor U9515 (N_9515,N_9358,N_9276);
nor U9516 (N_9516,N_9392,N_9289);
nor U9517 (N_9517,N_9343,N_9227);
xor U9518 (N_9518,N_9370,N_9343);
nand U9519 (N_9519,N_9368,N_9216);
or U9520 (N_9520,N_9210,N_9255);
or U9521 (N_9521,N_9383,N_9352);
xor U9522 (N_9522,N_9236,N_9319);
or U9523 (N_9523,N_9389,N_9328);
or U9524 (N_9524,N_9237,N_9282);
and U9525 (N_9525,N_9227,N_9248);
or U9526 (N_9526,N_9236,N_9315);
nand U9527 (N_9527,N_9394,N_9392);
and U9528 (N_9528,N_9216,N_9285);
and U9529 (N_9529,N_9279,N_9365);
and U9530 (N_9530,N_9279,N_9355);
nor U9531 (N_9531,N_9396,N_9274);
nor U9532 (N_9532,N_9336,N_9392);
nand U9533 (N_9533,N_9265,N_9350);
xor U9534 (N_9534,N_9213,N_9247);
or U9535 (N_9535,N_9277,N_9369);
xnor U9536 (N_9536,N_9234,N_9384);
nor U9537 (N_9537,N_9225,N_9254);
or U9538 (N_9538,N_9217,N_9219);
xor U9539 (N_9539,N_9392,N_9226);
and U9540 (N_9540,N_9398,N_9345);
nand U9541 (N_9541,N_9303,N_9317);
nor U9542 (N_9542,N_9261,N_9376);
and U9543 (N_9543,N_9287,N_9286);
nand U9544 (N_9544,N_9299,N_9200);
and U9545 (N_9545,N_9322,N_9319);
nand U9546 (N_9546,N_9398,N_9233);
nand U9547 (N_9547,N_9358,N_9293);
and U9548 (N_9548,N_9277,N_9376);
nor U9549 (N_9549,N_9275,N_9298);
or U9550 (N_9550,N_9357,N_9262);
xnor U9551 (N_9551,N_9329,N_9276);
or U9552 (N_9552,N_9216,N_9312);
or U9553 (N_9553,N_9373,N_9348);
xor U9554 (N_9554,N_9356,N_9200);
nor U9555 (N_9555,N_9371,N_9393);
or U9556 (N_9556,N_9370,N_9331);
xor U9557 (N_9557,N_9334,N_9263);
nand U9558 (N_9558,N_9388,N_9292);
nand U9559 (N_9559,N_9325,N_9200);
nor U9560 (N_9560,N_9358,N_9213);
nand U9561 (N_9561,N_9310,N_9338);
nor U9562 (N_9562,N_9353,N_9318);
xor U9563 (N_9563,N_9360,N_9245);
nand U9564 (N_9564,N_9276,N_9327);
and U9565 (N_9565,N_9208,N_9219);
nand U9566 (N_9566,N_9255,N_9253);
nand U9567 (N_9567,N_9297,N_9261);
and U9568 (N_9568,N_9312,N_9231);
and U9569 (N_9569,N_9376,N_9286);
and U9570 (N_9570,N_9365,N_9360);
nor U9571 (N_9571,N_9292,N_9378);
and U9572 (N_9572,N_9254,N_9333);
and U9573 (N_9573,N_9357,N_9282);
or U9574 (N_9574,N_9333,N_9381);
and U9575 (N_9575,N_9248,N_9335);
and U9576 (N_9576,N_9309,N_9283);
or U9577 (N_9577,N_9393,N_9229);
nor U9578 (N_9578,N_9381,N_9363);
xnor U9579 (N_9579,N_9276,N_9364);
and U9580 (N_9580,N_9256,N_9211);
and U9581 (N_9581,N_9275,N_9283);
or U9582 (N_9582,N_9352,N_9328);
and U9583 (N_9583,N_9350,N_9201);
xnor U9584 (N_9584,N_9259,N_9361);
or U9585 (N_9585,N_9352,N_9323);
nand U9586 (N_9586,N_9233,N_9378);
xnor U9587 (N_9587,N_9357,N_9396);
nor U9588 (N_9588,N_9331,N_9355);
nor U9589 (N_9589,N_9216,N_9396);
xnor U9590 (N_9590,N_9284,N_9241);
nor U9591 (N_9591,N_9390,N_9354);
and U9592 (N_9592,N_9386,N_9343);
xor U9593 (N_9593,N_9317,N_9362);
nor U9594 (N_9594,N_9239,N_9214);
or U9595 (N_9595,N_9344,N_9294);
nor U9596 (N_9596,N_9242,N_9327);
nor U9597 (N_9597,N_9338,N_9251);
nor U9598 (N_9598,N_9211,N_9290);
and U9599 (N_9599,N_9265,N_9295);
nand U9600 (N_9600,N_9577,N_9596);
or U9601 (N_9601,N_9564,N_9405);
nor U9602 (N_9602,N_9569,N_9479);
xnor U9603 (N_9603,N_9400,N_9553);
nor U9604 (N_9604,N_9548,N_9470);
and U9605 (N_9605,N_9535,N_9526);
nor U9606 (N_9606,N_9512,N_9586);
xor U9607 (N_9607,N_9509,N_9568);
xor U9608 (N_9608,N_9552,N_9446);
and U9609 (N_9609,N_9562,N_9412);
nand U9610 (N_9610,N_9591,N_9524);
and U9611 (N_9611,N_9543,N_9421);
and U9612 (N_9612,N_9460,N_9403);
xor U9613 (N_9613,N_9461,N_9589);
and U9614 (N_9614,N_9522,N_9554);
or U9615 (N_9615,N_9532,N_9468);
or U9616 (N_9616,N_9527,N_9525);
nor U9617 (N_9617,N_9503,N_9563);
xor U9618 (N_9618,N_9587,N_9549);
nor U9619 (N_9619,N_9423,N_9481);
xnor U9620 (N_9620,N_9440,N_9570);
or U9621 (N_9621,N_9567,N_9437);
nor U9622 (N_9622,N_9447,N_9558);
nor U9623 (N_9623,N_9555,N_9443);
nor U9624 (N_9624,N_9414,N_9534);
or U9625 (N_9625,N_9599,N_9530);
nand U9626 (N_9626,N_9420,N_9478);
and U9627 (N_9627,N_9542,N_9444);
nor U9628 (N_9628,N_9445,N_9408);
or U9629 (N_9629,N_9401,N_9545);
nor U9630 (N_9630,N_9463,N_9594);
or U9631 (N_9631,N_9514,N_9583);
xnor U9632 (N_9632,N_9546,N_9458);
nor U9633 (N_9633,N_9550,N_9584);
or U9634 (N_9634,N_9469,N_9511);
and U9635 (N_9635,N_9531,N_9588);
nor U9636 (N_9636,N_9472,N_9415);
nand U9637 (N_9637,N_9510,N_9572);
or U9638 (N_9638,N_9457,N_9474);
nand U9639 (N_9639,N_9560,N_9404);
or U9640 (N_9640,N_9465,N_9565);
and U9641 (N_9641,N_9559,N_9533);
nand U9642 (N_9642,N_9536,N_9467);
nor U9643 (N_9643,N_9482,N_9590);
nand U9644 (N_9644,N_9430,N_9402);
or U9645 (N_9645,N_9449,N_9574);
or U9646 (N_9646,N_9413,N_9561);
nand U9647 (N_9647,N_9480,N_9433);
xnor U9648 (N_9648,N_9450,N_9556);
nand U9649 (N_9649,N_9496,N_9505);
nor U9650 (N_9650,N_9487,N_9455);
and U9651 (N_9651,N_9418,N_9452);
or U9652 (N_9652,N_9571,N_9442);
and U9653 (N_9653,N_9491,N_9406);
or U9654 (N_9654,N_9597,N_9429);
nand U9655 (N_9655,N_9477,N_9432);
or U9656 (N_9656,N_9581,N_9436);
nor U9657 (N_9657,N_9579,N_9488);
or U9658 (N_9658,N_9409,N_9498);
xnor U9659 (N_9659,N_9504,N_9434);
xor U9660 (N_9660,N_9501,N_9464);
xnor U9661 (N_9661,N_9598,N_9416);
and U9662 (N_9662,N_9502,N_9476);
nand U9663 (N_9663,N_9507,N_9438);
and U9664 (N_9664,N_9493,N_9489);
nor U9665 (N_9665,N_9528,N_9483);
nand U9666 (N_9666,N_9427,N_9519);
xnor U9667 (N_9667,N_9499,N_9544);
or U9668 (N_9668,N_9431,N_9454);
nand U9669 (N_9669,N_9518,N_9486);
and U9670 (N_9670,N_9497,N_9576);
or U9671 (N_9671,N_9557,N_9453);
xor U9672 (N_9672,N_9494,N_9537);
xor U9673 (N_9673,N_9538,N_9466);
xnor U9674 (N_9674,N_9539,N_9515);
or U9675 (N_9675,N_9541,N_9417);
nor U9676 (N_9676,N_9513,N_9475);
or U9677 (N_9677,N_9439,N_9566);
or U9678 (N_9678,N_9523,N_9540);
xor U9679 (N_9679,N_9441,N_9506);
or U9680 (N_9680,N_9573,N_9435);
xnor U9681 (N_9681,N_9448,N_9516);
nand U9682 (N_9682,N_9422,N_9428);
or U9683 (N_9683,N_9508,N_9547);
nor U9684 (N_9684,N_9520,N_9473);
xnor U9685 (N_9685,N_9593,N_9551);
xor U9686 (N_9686,N_9462,N_9456);
xor U9687 (N_9687,N_9582,N_9424);
and U9688 (N_9688,N_9500,N_9521);
nor U9689 (N_9689,N_9451,N_9411);
nor U9690 (N_9690,N_9410,N_9484);
nor U9691 (N_9691,N_9595,N_9585);
and U9692 (N_9692,N_9407,N_9471);
xnor U9693 (N_9693,N_9575,N_9529);
or U9694 (N_9694,N_9580,N_9419);
or U9695 (N_9695,N_9578,N_9492);
or U9696 (N_9696,N_9592,N_9459);
nand U9697 (N_9697,N_9490,N_9485);
xnor U9698 (N_9698,N_9426,N_9517);
xor U9699 (N_9699,N_9495,N_9425);
xnor U9700 (N_9700,N_9558,N_9511);
nand U9701 (N_9701,N_9457,N_9525);
or U9702 (N_9702,N_9531,N_9560);
nor U9703 (N_9703,N_9593,N_9541);
or U9704 (N_9704,N_9418,N_9436);
or U9705 (N_9705,N_9537,N_9544);
and U9706 (N_9706,N_9438,N_9409);
or U9707 (N_9707,N_9498,N_9530);
xnor U9708 (N_9708,N_9416,N_9551);
or U9709 (N_9709,N_9530,N_9474);
or U9710 (N_9710,N_9407,N_9578);
xnor U9711 (N_9711,N_9428,N_9408);
xor U9712 (N_9712,N_9512,N_9414);
or U9713 (N_9713,N_9419,N_9437);
nand U9714 (N_9714,N_9512,N_9554);
xnor U9715 (N_9715,N_9582,N_9564);
xnor U9716 (N_9716,N_9425,N_9465);
xor U9717 (N_9717,N_9461,N_9498);
nor U9718 (N_9718,N_9503,N_9591);
and U9719 (N_9719,N_9487,N_9477);
xnor U9720 (N_9720,N_9417,N_9513);
and U9721 (N_9721,N_9413,N_9401);
or U9722 (N_9722,N_9402,N_9554);
or U9723 (N_9723,N_9452,N_9463);
nor U9724 (N_9724,N_9489,N_9446);
xor U9725 (N_9725,N_9447,N_9445);
and U9726 (N_9726,N_9569,N_9544);
xnor U9727 (N_9727,N_9450,N_9473);
nor U9728 (N_9728,N_9489,N_9455);
nand U9729 (N_9729,N_9486,N_9445);
and U9730 (N_9730,N_9449,N_9472);
or U9731 (N_9731,N_9440,N_9446);
nor U9732 (N_9732,N_9578,N_9469);
nor U9733 (N_9733,N_9410,N_9486);
nand U9734 (N_9734,N_9491,N_9566);
xnor U9735 (N_9735,N_9429,N_9450);
and U9736 (N_9736,N_9466,N_9471);
xnor U9737 (N_9737,N_9417,N_9499);
xnor U9738 (N_9738,N_9466,N_9448);
or U9739 (N_9739,N_9494,N_9487);
nor U9740 (N_9740,N_9479,N_9522);
xnor U9741 (N_9741,N_9496,N_9459);
nor U9742 (N_9742,N_9465,N_9511);
and U9743 (N_9743,N_9463,N_9541);
nand U9744 (N_9744,N_9487,N_9570);
nor U9745 (N_9745,N_9480,N_9512);
and U9746 (N_9746,N_9408,N_9542);
xor U9747 (N_9747,N_9468,N_9478);
or U9748 (N_9748,N_9535,N_9545);
nand U9749 (N_9749,N_9495,N_9451);
nand U9750 (N_9750,N_9409,N_9467);
or U9751 (N_9751,N_9499,N_9478);
and U9752 (N_9752,N_9588,N_9473);
or U9753 (N_9753,N_9458,N_9575);
xnor U9754 (N_9754,N_9469,N_9415);
and U9755 (N_9755,N_9571,N_9545);
or U9756 (N_9756,N_9547,N_9410);
nand U9757 (N_9757,N_9507,N_9451);
and U9758 (N_9758,N_9484,N_9516);
nand U9759 (N_9759,N_9595,N_9555);
nand U9760 (N_9760,N_9435,N_9554);
xor U9761 (N_9761,N_9473,N_9430);
or U9762 (N_9762,N_9491,N_9526);
and U9763 (N_9763,N_9490,N_9461);
or U9764 (N_9764,N_9589,N_9487);
xor U9765 (N_9765,N_9501,N_9502);
nor U9766 (N_9766,N_9538,N_9462);
or U9767 (N_9767,N_9581,N_9494);
nand U9768 (N_9768,N_9412,N_9590);
or U9769 (N_9769,N_9524,N_9449);
and U9770 (N_9770,N_9425,N_9555);
nand U9771 (N_9771,N_9591,N_9523);
xnor U9772 (N_9772,N_9403,N_9587);
and U9773 (N_9773,N_9557,N_9487);
and U9774 (N_9774,N_9518,N_9458);
nor U9775 (N_9775,N_9422,N_9460);
nor U9776 (N_9776,N_9483,N_9510);
xor U9777 (N_9777,N_9494,N_9577);
nor U9778 (N_9778,N_9436,N_9469);
or U9779 (N_9779,N_9418,N_9583);
or U9780 (N_9780,N_9560,N_9552);
or U9781 (N_9781,N_9558,N_9416);
and U9782 (N_9782,N_9522,N_9533);
and U9783 (N_9783,N_9542,N_9534);
nand U9784 (N_9784,N_9517,N_9579);
nor U9785 (N_9785,N_9491,N_9592);
and U9786 (N_9786,N_9401,N_9523);
or U9787 (N_9787,N_9436,N_9568);
or U9788 (N_9788,N_9502,N_9516);
xor U9789 (N_9789,N_9451,N_9491);
and U9790 (N_9790,N_9539,N_9414);
or U9791 (N_9791,N_9411,N_9576);
xor U9792 (N_9792,N_9530,N_9457);
nand U9793 (N_9793,N_9576,N_9420);
nor U9794 (N_9794,N_9414,N_9473);
xnor U9795 (N_9795,N_9450,N_9420);
and U9796 (N_9796,N_9528,N_9503);
or U9797 (N_9797,N_9593,N_9523);
and U9798 (N_9798,N_9577,N_9434);
nand U9799 (N_9799,N_9447,N_9475);
xnor U9800 (N_9800,N_9726,N_9648);
nor U9801 (N_9801,N_9624,N_9701);
nand U9802 (N_9802,N_9778,N_9621);
nand U9803 (N_9803,N_9661,N_9714);
nor U9804 (N_9804,N_9659,N_9706);
nor U9805 (N_9805,N_9623,N_9657);
and U9806 (N_9806,N_9777,N_9737);
nor U9807 (N_9807,N_9782,N_9727);
nor U9808 (N_9808,N_9733,N_9679);
and U9809 (N_9809,N_9795,N_9616);
or U9810 (N_9810,N_9700,N_9710);
and U9811 (N_9811,N_9754,N_9681);
nor U9812 (N_9812,N_9652,N_9758);
and U9813 (N_9813,N_9673,N_9677);
or U9814 (N_9814,N_9744,N_9745);
or U9815 (N_9815,N_9746,N_9761);
and U9816 (N_9816,N_9609,N_9707);
nand U9817 (N_9817,N_9667,N_9721);
nand U9818 (N_9818,N_9762,N_9763);
or U9819 (N_9819,N_9760,N_9725);
nand U9820 (N_9820,N_9772,N_9783);
nand U9821 (N_9821,N_9645,N_9632);
or U9822 (N_9822,N_9653,N_9643);
nor U9823 (N_9823,N_9757,N_9613);
and U9824 (N_9824,N_9708,N_9791);
xor U9825 (N_9825,N_9743,N_9713);
nand U9826 (N_9826,N_9704,N_9784);
or U9827 (N_9827,N_9687,N_9719);
nor U9828 (N_9828,N_9690,N_9739);
and U9829 (N_9829,N_9734,N_9693);
or U9830 (N_9830,N_9751,N_9773);
xor U9831 (N_9831,N_9634,N_9697);
or U9832 (N_9832,N_9639,N_9664);
or U9833 (N_9833,N_9793,N_9781);
and U9834 (N_9834,N_9640,N_9615);
nand U9835 (N_9835,N_9668,N_9633);
xor U9836 (N_9836,N_9626,N_9741);
nand U9837 (N_9837,N_9790,N_9675);
nand U9838 (N_9838,N_9750,N_9684);
nand U9839 (N_9839,N_9711,N_9604);
nor U9840 (N_9840,N_9646,N_9798);
nor U9841 (N_9841,N_9601,N_9663);
or U9842 (N_9842,N_9605,N_9769);
xnor U9843 (N_9843,N_9674,N_9665);
or U9844 (N_9844,N_9644,N_9670);
nand U9845 (N_9845,N_9678,N_9655);
nor U9846 (N_9846,N_9768,N_9635);
nor U9847 (N_9847,N_9729,N_9617);
or U9848 (N_9848,N_9703,N_9686);
xor U9849 (N_9849,N_9636,N_9694);
nand U9850 (N_9850,N_9669,N_9740);
nand U9851 (N_9851,N_9662,N_9614);
or U9852 (N_9852,N_9787,N_9622);
nand U9853 (N_9853,N_9767,N_9785);
and U9854 (N_9854,N_9619,N_9628);
nor U9855 (N_9855,N_9649,N_9759);
nand U9856 (N_9856,N_9683,N_9748);
or U9857 (N_9857,N_9776,N_9606);
or U9858 (N_9858,N_9647,N_9738);
xor U9859 (N_9859,N_9797,N_9756);
or U9860 (N_9860,N_9625,N_9642);
nand U9861 (N_9861,N_9731,N_9608);
and U9862 (N_9862,N_9792,N_9692);
and U9863 (N_9863,N_9765,N_9660);
and U9864 (N_9864,N_9732,N_9771);
xor U9865 (N_9865,N_9728,N_9724);
or U9866 (N_9866,N_9717,N_9709);
nand U9867 (N_9867,N_9650,N_9629);
and U9868 (N_9868,N_9658,N_9656);
and U9869 (N_9869,N_9752,N_9774);
nand U9870 (N_9870,N_9796,N_9651);
xor U9871 (N_9871,N_9695,N_9766);
xor U9872 (N_9872,N_9672,N_9638);
or U9873 (N_9873,N_9631,N_9666);
or U9874 (N_9874,N_9794,N_9627);
nand U9875 (N_9875,N_9775,N_9723);
xor U9876 (N_9876,N_9720,N_9730);
nand U9877 (N_9877,N_9780,N_9696);
and U9878 (N_9878,N_9689,N_9654);
xor U9879 (N_9879,N_9749,N_9718);
or U9880 (N_9880,N_9680,N_9671);
or U9881 (N_9881,N_9600,N_9712);
nand U9882 (N_9882,N_9607,N_9789);
and U9883 (N_9883,N_9685,N_9612);
nor U9884 (N_9884,N_9691,N_9641);
or U9885 (N_9885,N_9799,N_9637);
nor U9886 (N_9886,N_9702,N_9716);
or U9887 (N_9887,N_9676,N_9779);
or U9888 (N_9888,N_9786,N_9602);
xor U9889 (N_9889,N_9620,N_9742);
and U9890 (N_9890,N_9788,N_9698);
xnor U9891 (N_9891,N_9755,N_9715);
nor U9892 (N_9892,N_9736,N_9682);
xor U9893 (N_9893,N_9764,N_9753);
nand U9894 (N_9894,N_9735,N_9770);
or U9895 (N_9895,N_9611,N_9603);
or U9896 (N_9896,N_9722,N_9688);
or U9897 (N_9897,N_9699,N_9618);
nor U9898 (N_9898,N_9747,N_9705);
and U9899 (N_9899,N_9630,N_9610);
and U9900 (N_9900,N_9763,N_9666);
xnor U9901 (N_9901,N_9698,N_9783);
xor U9902 (N_9902,N_9657,N_9695);
nand U9903 (N_9903,N_9724,N_9620);
xnor U9904 (N_9904,N_9747,N_9765);
and U9905 (N_9905,N_9614,N_9751);
or U9906 (N_9906,N_9692,N_9619);
or U9907 (N_9907,N_9709,N_9791);
or U9908 (N_9908,N_9786,N_9752);
xor U9909 (N_9909,N_9758,N_9743);
xnor U9910 (N_9910,N_9735,N_9753);
and U9911 (N_9911,N_9729,N_9783);
and U9912 (N_9912,N_9663,N_9786);
nand U9913 (N_9913,N_9752,N_9681);
xor U9914 (N_9914,N_9766,N_9691);
and U9915 (N_9915,N_9648,N_9627);
nand U9916 (N_9916,N_9770,N_9780);
nor U9917 (N_9917,N_9755,N_9757);
xor U9918 (N_9918,N_9728,N_9606);
xnor U9919 (N_9919,N_9788,N_9639);
xor U9920 (N_9920,N_9644,N_9708);
nor U9921 (N_9921,N_9724,N_9679);
nor U9922 (N_9922,N_9766,N_9647);
or U9923 (N_9923,N_9753,N_9607);
and U9924 (N_9924,N_9623,N_9699);
xor U9925 (N_9925,N_9670,N_9631);
and U9926 (N_9926,N_9631,N_9638);
xnor U9927 (N_9927,N_9751,N_9608);
nor U9928 (N_9928,N_9638,N_9683);
nor U9929 (N_9929,N_9727,N_9669);
and U9930 (N_9930,N_9664,N_9792);
and U9931 (N_9931,N_9758,N_9633);
nand U9932 (N_9932,N_9654,N_9668);
nand U9933 (N_9933,N_9779,N_9621);
nand U9934 (N_9934,N_9679,N_9749);
and U9935 (N_9935,N_9672,N_9714);
or U9936 (N_9936,N_9687,N_9680);
nand U9937 (N_9937,N_9778,N_9689);
and U9938 (N_9938,N_9670,N_9615);
nand U9939 (N_9939,N_9620,N_9643);
nand U9940 (N_9940,N_9658,N_9666);
xnor U9941 (N_9941,N_9603,N_9789);
nand U9942 (N_9942,N_9730,N_9768);
and U9943 (N_9943,N_9767,N_9701);
xnor U9944 (N_9944,N_9616,N_9695);
nor U9945 (N_9945,N_9668,N_9690);
and U9946 (N_9946,N_9694,N_9728);
nand U9947 (N_9947,N_9693,N_9629);
and U9948 (N_9948,N_9789,N_9618);
nand U9949 (N_9949,N_9792,N_9667);
and U9950 (N_9950,N_9714,N_9799);
nor U9951 (N_9951,N_9669,N_9732);
xor U9952 (N_9952,N_9753,N_9793);
and U9953 (N_9953,N_9670,N_9713);
and U9954 (N_9954,N_9631,N_9759);
and U9955 (N_9955,N_9787,N_9617);
nor U9956 (N_9956,N_9775,N_9653);
nand U9957 (N_9957,N_9787,N_9615);
or U9958 (N_9958,N_9709,N_9664);
and U9959 (N_9959,N_9680,N_9604);
xor U9960 (N_9960,N_9665,N_9731);
nor U9961 (N_9961,N_9704,N_9716);
or U9962 (N_9962,N_9768,N_9700);
and U9963 (N_9963,N_9790,N_9735);
nor U9964 (N_9964,N_9703,N_9637);
nand U9965 (N_9965,N_9731,N_9793);
or U9966 (N_9966,N_9718,N_9795);
and U9967 (N_9967,N_9680,N_9697);
xor U9968 (N_9968,N_9792,N_9609);
nor U9969 (N_9969,N_9713,N_9632);
xnor U9970 (N_9970,N_9695,N_9723);
nand U9971 (N_9971,N_9796,N_9618);
and U9972 (N_9972,N_9710,N_9686);
nand U9973 (N_9973,N_9720,N_9668);
and U9974 (N_9974,N_9711,N_9724);
nand U9975 (N_9975,N_9747,N_9722);
nor U9976 (N_9976,N_9734,N_9708);
nand U9977 (N_9977,N_9790,N_9706);
and U9978 (N_9978,N_9639,N_9601);
or U9979 (N_9979,N_9641,N_9628);
or U9980 (N_9980,N_9731,N_9729);
nor U9981 (N_9981,N_9661,N_9793);
nor U9982 (N_9982,N_9607,N_9750);
or U9983 (N_9983,N_9692,N_9704);
xor U9984 (N_9984,N_9662,N_9621);
and U9985 (N_9985,N_9743,N_9737);
nand U9986 (N_9986,N_9644,N_9676);
and U9987 (N_9987,N_9683,N_9670);
nor U9988 (N_9988,N_9600,N_9789);
xor U9989 (N_9989,N_9768,N_9655);
and U9990 (N_9990,N_9601,N_9734);
and U9991 (N_9991,N_9729,N_9648);
nor U9992 (N_9992,N_9636,N_9683);
or U9993 (N_9993,N_9787,N_9605);
and U9994 (N_9994,N_9617,N_9725);
nand U9995 (N_9995,N_9620,N_9700);
and U9996 (N_9996,N_9790,N_9753);
nor U9997 (N_9997,N_9602,N_9614);
nor U9998 (N_9998,N_9778,N_9633);
nand U9999 (N_9999,N_9766,N_9782);
and U10000 (N_10000,N_9883,N_9930);
nand U10001 (N_10001,N_9898,N_9899);
xnor U10002 (N_10002,N_9901,N_9892);
nor U10003 (N_10003,N_9902,N_9880);
xnor U10004 (N_10004,N_9807,N_9992);
and U10005 (N_10005,N_9873,N_9900);
nand U10006 (N_10006,N_9998,N_9826);
nor U10007 (N_10007,N_9856,N_9920);
nand U10008 (N_10008,N_9805,N_9868);
or U10009 (N_10009,N_9957,N_9859);
or U10010 (N_10010,N_9939,N_9876);
and U10011 (N_10011,N_9905,N_9976);
or U10012 (N_10012,N_9829,N_9843);
nand U10013 (N_10013,N_9879,N_9926);
xnor U10014 (N_10014,N_9889,N_9855);
and U10015 (N_10015,N_9913,N_9987);
and U10016 (N_10016,N_9935,N_9921);
or U10017 (N_10017,N_9980,N_9949);
or U10018 (N_10018,N_9986,N_9941);
xnor U10019 (N_10019,N_9842,N_9997);
xnor U10020 (N_10020,N_9929,N_9928);
nor U10021 (N_10021,N_9955,N_9831);
nor U10022 (N_10022,N_9828,N_9847);
or U10023 (N_10023,N_9836,N_9864);
nor U10024 (N_10024,N_9870,N_9852);
xor U10025 (N_10025,N_9890,N_9991);
nor U10026 (N_10026,N_9824,N_9954);
nand U10027 (N_10027,N_9952,N_9869);
xor U10028 (N_10028,N_9802,N_9906);
and U10029 (N_10029,N_9912,N_9819);
nor U10030 (N_10030,N_9993,N_9881);
nor U10031 (N_10031,N_9996,N_9968);
nor U10032 (N_10032,N_9896,N_9950);
xor U10033 (N_10033,N_9959,N_9885);
or U10034 (N_10034,N_9811,N_9841);
and U10035 (N_10035,N_9973,N_9882);
nor U10036 (N_10036,N_9853,N_9851);
or U10037 (N_10037,N_9985,N_9867);
and U10038 (N_10038,N_9972,N_9922);
xor U10039 (N_10039,N_9812,N_9931);
or U10040 (N_10040,N_9917,N_9801);
nand U10041 (N_10041,N_9871,N_9914);
and U10042 (N_10042,N_9903,N_9895);
and U10043 (N_10043,N_9887,N_9800);
nand U10044 (N_10044,N_9933,N_9814);
and U10045 (N_10045,N_9809,N_9817);
nand U10046 (N_10046,N_9951,N_9848);
or U10047 (N_10047,N_9907,N_9983);
nor U10048 (N_10048,N_9915,N_9988);
nand U10049 (N_10049,N_9823,N_9821);
xnor U10050 (N_10050,N_9813,N_9863);
xor U10051 (N_10051,N_9924,N_9978);
nand U10052 (N_10052,N_9891,N_9904);
or U10053 (N_10053,N_9875,N_9844);
and U10054 (N_10054,N_9846,N_9936);
and U10055 (N_10055,N_9865,N_9984);
xnor U10056 (N_10056,N_9925,N_9832);
xor U10057 (N_10057,N_9893,N_9818);
nor U10058 (N_10058,N_9849,N_9910);
and U10059 (N_10059,N_9944,N_9969);
nand U10060 (N_10060,N_9861,N_9872);
or U10061 (N_10061,N_9945,N_9977);
nor U10062 (N_10062,N_9961,N_9909);
nor U10063 (N_10063,N_9990,N_9975);
or U10064 (N_10064,N_9816,N_9974);
and U10065 (N_10065,N_9923,N_9989);
xor U10066 (N_10066,N_9884,N_9850);
and U10067 (N_10067,N_9845,N_9894);
and U10068 (N_10068,N_9854,N_9981);
or U10069 (N_10069,N_9916,N_9964);
or U10070 (N_10070,N_9970,N_9934);
or U10071 (N_10071,N_9803,N_9956);
nor U10072 (N_10072,N_9938,N_9810);
nand U10073 (N_10073,N_9808,N_9948);
and U10074 (N_10074,N_9966,N_9837);
nor U10075 (N_10075,N_9835,N_9953);
or U10076 (N_10076,N_9815,N_9962);
xnor U10077 (N_10077,N_9862,N_9874);
xor U10078 (N_10078,N_9927,N_9833);
or U10079 (N_10079,N_9866,N_9888);
or U10080 (N_10080,N_9999,N_9967);
nor U10081 (N_10081,N_9908,N_9979);
nor U10082 (N_10082,N_9806,N_9940);
or U10083 (N_10083,N_9825,N_9860);
nand U10084 (N_10084,N_9830,N_9918);
nor U10085 (N_10085,N_9958,N_9982);
nand U10086 (N_10086,N_9804,N_9877);
nand U10087 (N_10087,N_9937,N_9897);
and U10088 (N_10088,N_9942,N_9947);
nor U10089 (N_10089,N_9960,N_9838);
or U10090 (N_10090,N_9827,N_9963);
or U10091 (N_10091,N_9994,N_9858);
and U10092 (N_10092,N_9943,N_9839);
nand U10093 (N_10093,N_9878,N_9946);
or U10094 (N_10094,N_9919,N_9834);
nand U10095 (N_10095,N_9932,N_9820);
nor U10096 (N_10096,N_9857,N_9822);
xor U10097 (N_10097,N_9886,N_9995);
nand U10098 (N_10098,N_9911,N_9971);
and U10099 (N_10099,N_9965,N_9840);
nor U10100 (N_10100,N_9927,N_9891);
or U10101 (N_10101,N_9846,N_9972);
xnor U10102 (N_10102,N_9905,N_9858);
nand U10103 (N_10103,N_9938,N_9933);
xnor U10104 (N_10104,N_9929,N_9866);
xnor U10105 (N_10105,N_9948,N_9933);
nor U10106 (N_10106,N_9879,N_9935);
xor U10107 (N_10107,N_9971,N_9885);
xnor U10108 (N_10108,N_9993,N_9811);
and U10109 (N_10109,N_9914,N_9891);
or U10110 (N_10110,N_9988,N_9829);
and U10111 (N_10111,N_9942,N_9842);
nor U10112 (N_10112,N_9986,N_9810);
xor U10113 (N_10113,N_9912,N_9906);
nor U10114 (N_10114,N_9873,N_9893);
xor U10115 (N_10115,N_9926,N_9880);
or U10116 (N_10116,N_9928,N_9800);
xnor U10117 (N_10117,N_9963,N_9967);
xor U10118 (N_10118,N_9838,N_9902);
nand U10119 (N_10119,N_9873,N_9854);
nand U10120 (N_10120,N_9905,N_9861);
or U10121 (N_10121,N_9828,N_9940);
and U10122 (N_10122,N_9848,N_9930);
nand U10123 (N_10123,N_9984,N_9917);
xor U10124 (N_10124,N_9952,N_9941);
or U10125 (N_10125,N_9932,N_9850);
xor U10126 (N_10126,N_9865,N_9959);
nor U10127 (N_10127,N_9994,N_9998);
xor U10128 (N_10128,N_9901,N_9849);
xor U10129 (N_10129,N_9884,N_9894);
nand U10130 (N_10130,N_9900,N_9954);
or U10131 (N_10131,N_9951,N_9908);
nand U10132 (N_10132,N_9977,N_9954);
and U10133 (N_10133,N_9948,N_9995);
xnor U10134 (N_10134,N_9904,N_9907);
xor U10135 (N_10135,N_9871,N_9877);
xnor U10136 (N_10136,N_9963,N_9845);
nand U10137 (N_10137,N_9885,N_9937);
nor U10138 (N_10138,N_9859,N_9977);
nand U10139 (N_10139,N_9833,N_9845);
nor U10140 (N_10140,N_9861,N_9845);
or U10141 (N_10141,N_9829,N_9876);
or U10142 (N_10142,N_9833,N_9810);
nor U10143 (N_10143,N_9946,N_9891);
and U10144 (N_10144,N_9813,N_9906);
xor U10145 (N_10145,N_9875,N_9917);
xor U10146 (N_10146,N_9833,N_9976);
nor U10147 (N_10147,N_9911,N_9830);
xor U10148 (N_10148,N_9846,N_9899);
xor U10149 (N_10149,N_9988,N_9996);
nand U10150 (N_10150,N_9831,N_9959);
xnor U10151 (N_10151,N_9913,N_9859);
nor U10152 (N_10152,N_9902,N_9998);
nand U10153 (N_10153,N_9892,N_9923);
xor U10154 (N_10154,N_9885,N_9852);
or U10155 (N_10155,N_9936,N_9944);
and U10156 (N_10156,N_9997,N_9937);
nor U10157 (N_10157,N_9991,N_9904);
or U10158 (N_10158,N_9985,N_9868);
or U10159 (N_10159,N_9907,N_9848);
xor U10160 (N_10160,N_9883,N_9854);
and U10161 (N_10161,N_9908,N_9904);
nand U10162 (N_10162,N_9801,N_9898);
nor U10163 (N_10163,N_9830,N_9843);
nor U10164 (N_10164,N_9834,N_9902);
or U10165 (N_10165,N_9914,N_9963);
xnor U10166 (N_10166,N_9845,N_9801);
or U10167 (N_10167,N_9971,N_9848);
or U10168 (N_10168,N_9931,N_9923);
nor U10169 (N_10169,N_9891,N_9886);
xor U10170 (N_10170,N_9816,N_9873);
xnor U10171 (N_10171,N_9935,N_9869);
xnor U10172 (N_10172,N_9884,N_9948);
xnor U10173 (N_10173,N_9921,N_9909);
nor U10174 (N_10174,N_9996,N_9975);
xnor U10175 (N_10175,N_9810,N_9901);
or U10176 (N_10176,N_9870,N_9874);
xnor U10177 (N_10177,N_9979,N_9999);
nor U10178 (N_10178,N_9845,N_9981);
xor U10179 (N_10179,N_9820,N_9934);
nor U10180 (N_10180,N_9994,N_9838);
nand U10181 (N_10181,N_9801,N_9987);
or U10182 (N_10182,N_9931,N_9911);
or U10183 (N_10183,N_9874,N_9820);
nand U10184 (N_10184,N_9937,N_9936);
or U10185 (N_10185,N_9890,N_9845);
or U10186 (N_10186,N_9971,N_9931);
and U10187 (N_10187,N_9911,N_9921);
nand U10188 (N_10188,N_9857,N_9873);
nand U10189 (N_10189,N_9900,N_9966);
or U10190 (N_10190,N_9838,N_9898);
xnor U10191 (N_10191,N_9903,N_9802);
nor U10192 (N_10192,N_9823,N_9900);
nor U10193 (N_10193,N_9928,N_9997);
or U10194 (N_10194,N_9861,N_9934);
xnor U10195 (N_10195,N_9871,N_9873);
and U10196 (N_10196,N_9834,N_9882);
and U10197 (N_10197,N_9822,N_9919);
xor U10198 (N_10198,N_9893,N_9896);
xnor U10199 (N_10199,N_9819,N_9870);
and U10200 (N_10200,N_10156,N_10071);
xnor U10201 (N_10201,N_10177,N_10110);
xnor U10202 (N_10202,N_10093,N_10180);
and U10203 (N_10203,N_10175,N_10066);
nor U10204 (N_10204,N_10128,N_10152);
nand U10205 (N_10205,N_10002,N_10191);
nor U10206 (N_10206,N_10131,N_10115);
nand U10207 (N_10207,N_10084,N_10146);
or U10208 (N_10208,N_10104,N_10012);
and U10209 (N_10209,N_10140,N_10057);
nand U10210 (N_10210,N_10113,N_10196);
nor U10211 (N_10211,N_10042,N_10036);
and U10212 (N_10212,N_10044,N_10194);
xnor U10213 (N_10213,N_10018,N_10137);
or U10214 (N_10214,N_10145,N_10070);
xnor U10215 (N_10215,N_10157,N_10000);
nand U10216 (N_10216,N_10091,N_10103);
or U10217 (N_10217,N_10123,N_10199);
nor U10218 (N_10218,N_10179,N_10045);
nor U10219 (N_10219,N_10166,N_10190);
nor U10220 (N_10220,N_10171,N_10051);
nand U10221 (N_10221,N_10170,N_10069);
nor U10222 (N_10222,N_10035,N_10095);
or U10223 (N_10223,N_10024,N_10129);
and U10224 (N_10224,N_10038,N_10081);
or U10225 (N_10225,N_10004,N_10118);
nor U10226 (N_10226,N_10072,N_10155);
xor U10227 (N_10227,N_10039,N_10074);
or U10228 (N_10228,N_10100,N_10169);
nor U10229 (N_10229,N_10099,N_10174);
and U10230 (N_10230,N_10183,N_10067);
nand U10231 (N_10231,N_10089,N_10014);
xor U10232 (N_10232,N_10101,N_10083);
or U10233 (N_10233,N_10043,N_10154);
and U10234 (N_10234,N_10168,N_10141);
nor U10235 (N_10235,N_10165,N_10078);
xor U10236 (N_10236,N_10122,N_10173);
or U10237 (N_10237,N_10047,N_10003);
and U10238 (N_10238,N_10037,N_10094);
or U10239 (N_10239,N_10021,N_10050);
nor U10240 (N_10240,N_10148,N_10046);
and U10241 (N_10241,N_10181,N_10015);
and U10242 (N_10242,N_10108,N_10164);
and U10243 (N_10243,N_10007,N_10030);
and U10244 (N_10244,N_10106,N_10151);
nand U10245 (N_10245,N_10025,N_10011);
nor U10246 (N_10246,N_10060,N_10052);
nor U10247 (N_10247,N_10127,N_10197);
nor U10248 (N_10248,N_10090,N_10096);
and U10249 (N_10249,N_10133,N_10054);
xor U10250 (N_10250,N_10193,N_10126);
nor U10251 (N_10251,N_10041,N_10049);
nor U10252 (N_10252,N_10098,N_10028);
or U10253 (N_10253,N_10111,N_10013);
xor U10254 (N_10254,N_10023,N_10121);
or U10255 (N_10255,N_10105,N_10107);
nor U10256 (N_10256,N_10097,N_10144);
or U10257 (N_10257,N_10195,N_10027);
nor U10258 (N_10258,N_10082,N_10001);
and U10259 (N_10259,N_10068,N_10092);
xor U10260 (N_10260,N_10172,N_10119);
and U10261 (N_10261,N_10150,N_10117);
nand U10262 (N_10262,N_10153,N_10147);
and U10263 (N_10263,N_10125,N_10130);
nand U10264 (N_10264,N_10142,N_10182);
or U10265 (N_10265,N_10124,N_10186);
nor U10266 (N_10266,N_10010,N_10178);
or U10267 (N_10267,N_10059,N_10160);
and U10268 (N_10268,N_10022,N_10187);
or U10269 (N_10269,N_10132,N_10159);
and U10270 (N_10270,N_10031,N_10167);
or U10271 (N_10271,N_10020,N_10029);
or U10272 (N_10272,N_10076,N_10189);
nand U10273 (N_10273,N_10114,N_10065);
and U10274 (N_10274,N_10188,N_10026);
nor U10275 (N_10275,N_10079,N_10176);
and U10276 (N_10276,N_10143,N_10063);
xor U10277 (N_10277,N_10138,N_10058);
nor U10278 (N_10278,N_10185,N_10088);
or U10279 (N_10279,N_10009,N_10184);
xor U10280 (N_10280,N_10161,N_10073);
nor U10281 (N_10281,N_10149,N_10087);
xor U10282 (N_10282,N_10017,N_10075);
nor U10283 (N_10283,N_10086,N_10158);
nand U10284 (N_10284,N_10008,N_10134);
or U10285 (N_10285,N_10080,N_10062);
nor U10286 (N_10286,N_10109,N_10198);
or U10287 (N_10287,N_10061,N_10033);
nand U10288 (N_10288,N_10102,N_10040);
or U10289 (N_10289,N_10077,N_10034);
nand U10290 (N_10290,N_10005,N_10136);
and U10291 (N_10291,N_10053,N_10139);
nand U10292 (N_10292,N_10135,N_10048);
or U10293 (N_10293,N_10019,N_10162);
nor U10294 (N_10294,N_10064,N_10032);
nand U10295 (N_10295,N_10006,N_10112);
and U10296 (N_10296,N_10085,N_10192);
nor U10297 (N_10297,N_10163,N_10120);
xor U10298 (N_10298,N_10016,N_10116);
and U10299 (N_10299,N_10055,N_10056);
nor U10300 (N_10300,N_10045,N_10090);
nand U10301 (N_10301,N_10073,N_10074);
nand U10302 (N_10302,N_10167,N_10153);
and U10303 (N_10303,N_10042,N_10008);
or U10304 (N_10304,N_10151,N_10170);
nor U10305 (N_10305,N_10160,N_10095);
and U10306 (N_10306,N_10137,N_10005);
nor U10307 (N_10307,N_10034,N_10102);
and U10308 (N_10308,N_10174,N_10131);
nand U10309 (N_10309,N_10012,N_10121);
nand U10310 (N_10310,N_10119,N_10102);
nand U10311 (N_10311,N_10067,N_10104);
nor U10312 (N_10312,N_10159,N_10070);
nor U10313 (N_10313,N_10177,N_10053);
nand U10314 (N_10314,N_10041,N_10036);
xor U10315 (N_10315,N_10041,N_10096);
nor U10316 (N_10316,N_10191,N_10102);
xor U10317 (N_10317,N_10164,N_10172);
nand U10318 (N_10318,N_10103,N_10058);
and U10319 (N_10319,N_10005,N_10058);
xnor U10320 (N_10320,N_10071,N_10139);
nand U10321 (N_10321,N_10155,N_10196);
nand U10322 (N_10322,N_10165,N_10190);
xnor U10323 (N_10323,N_10131,N_10166);
nor U10324 (N_10324,N_10189,N_10042);
nand U10325 (N_10325,N_10060,N_10079);
nor U10326 (N_10326,N_10009,N_10144);
nor U10327 (N_10327,N_10113,N_10160);
nand U10328 (N_10328,N_10117,N_10077);
and U10329 (N_10329,N_10166,N_10123);
or U10330 (N_10330,N_10047,N_10139);
xnor U10331 (N_10331,N_10180,N_10147);
or U10332 (N_10332,N_10061,N_10167);
xor U10333 (N_10333,N_10141,N_10065);
nor U10334 (N_10334,N_10095,N_10138);
nor U10335 (N_10335,N_10014,N_10105);
nor U10336 (N_10336,N_10039,N_10087);
xnor U10337 (N_10337,N_10126,N_10092);
nand U10338 (N_10338,N_10086,N_10140);
nand U10339 (N_10339,N_10094,N_10177);
nand U10340 (N_10340,N_10031,N_10035);
or U10341 (N_10341,N_10070,N_10188);
nand U10342 (N_10342,N_10128,N_10022);
nor U10343 (N_10343,N_10170,N_10185);
nor U10344 (N_10344,N_10034,N_10149);
nand U10345 (N_10345,N_10033,N_10186);
and U10346 (N_10346,N_10061,N_10014);
nor U10347 (N_10347,N_10132,N_10099);
nor U10348 (N_10348,N_10193,N_10090);
nor U10349 (N_10349,N_10177,N_10054);
nand U10350 (N_10350,N_10023,N_10165);
nor U10351 (N_10351,N_10148,N_10080);
xor U10352 (N_10352,N_10019,N_10072);
nor U10353 (N_10353,N_10022,N_10148);
nand U10354 (N_10354,N_10037,N_10176);
nor U10355 (N_10355,N_10045,N_10087);
nand U10356 (N_10356,N_10105,N_10168);
xor U10357 (N_10357,N_10056,N_10169);
xnor U10358 (N_10358,N_10126,N_10042);
nand U10359 (N_10359,N_10006,N_10077);
xor U10360 (N_10360,N_10165,N_10093);
and U10361 (N_10361,N_10072,N_10179);
and U10362 (N_10362,N_10134,N_10146);
nand U10363 (N_10363,N_10185,N_10097);
and U10364 (N_10364,N_10176,N_10084);
nor U10365 (N_10365,N_10109,N_10075);
xnor U10366 (N_10366,N_10105,N_10009);
nand U10367 (N_10367,N_10121,N_10187);
xor U10368 (N_10368,N_10063,N_10197);
nor U10369 (N_10369,N_10075,N_10091);
or U10370 (N_10370,N_10001,N_10125);
or U10371 (N_10371,N_10053,N_10187);
xnor U10372 (N_10372,N_10066,N_10075);
nand U10373 (N_10373,N_10087,N_10085);
or U10374 (N_10374,N_10043,N_10052);
xor U10375 (N_10375,N_10146,N_10077);
nor U10376 (N_10376,N_10074,N_10125);
nor U10377 (N_10377,N_10187,N_10127);
nor U10378 (N_10378,N_10058,N_10116);
nand U10379 (N_10379,N_10197,N_10084);
or U10380 (N_10380,N_10157,N_10073);
xor U10381 (N_10381,N_10013,N_10095);
or U10382 (N_10382,N_10186,N_10118);
xor U10383 (N_10383,N_10194,N_10042);
nor U10384 (N_10384,N_10021,N_10096);
nor U10385 (N_10385,N_10189,N_10095);
nor U10386 (N_10386,N_10051,N_10079);
or U10387 (N_10387,N_10071,N_10056);
and U10388 (N_10388,N_10022,N_10157);
and U10389 (N_10389,N_10072,N_10006);
xor U10390 (N_10390,N_10014,N_10128);
nand U10391 (N_10391,N_10070,N_10148);
and U10392 (N_10392,N_10082,N_10171);
nor U10393 (N_10393,N_10147,N_10041);
or U10394 (N_10394,N_10189,N_10133);
xor U10395 (N_10395,N_10115,N_10096);
or U10396 (N_10396,N_10059,N_10128);
xnor U10397 (N_10397,N_10182,N_10086);
nand U10398 (N_10398,N_10108,N_10187);
xnor U10399 (N_10399,N_10093,N_10153);
or U10400 (N_10400,N_10202,N_10285);
nand U10401 (N_10401,N_10396,N_10360);
nand U10402 (N_10402,N_10370,N_10327);
and U10403 (N_10403,N_10217,N_10314);
nand U10404 (N_10404,N_10302,N_10204);
xnor U10405 (N_10405,N_10381,N_10395);
or U10406 (N_10406,N_10319,N_10211);
nand U10407 (N_10407,N_10260,N_10247);
xnor U10408 (N_10408,N_10226,N_10358);
nand U10409 (N_10409,N_10265,N_10359);
or U10410 (N_10410,N_10398,N_10235);
and U10411 (N_10411,N_10289,N_10266);
xor U10412 (N_10412,N_10207,N_10344);
xor U10413 (N_10413,N_10333,N_10248);
or U10414 (N_10414,N_10384,N_10349);
xor U10415 (N_10415,N_10342,N_10251);
and U10416 (N_10416,N_10318,N_10250);
nor U10417 (N_10417,N_10297,N_10218);
and U10418 (N_10418,N_10225,N_10375);
nor U10419 (N_10419,N_10267,N_10240);
and U10420 (N_10420,N_10364,N_10346);
or U10421 (N_10421,N_10334,N_10223);
xor U10422 (N_10422,N_10389,N_10283);
nor U10423 (N_10423,N_10227,N_10306);
nor U10424 (N_10424,N_10234,N_10237);
and U10425 (N_10425,N_10343,N_10254);
or U10426 (N_10426,N_10230,N_10262);
or U10427 (N_10427,N_10373,N_10268);
nor U10428 (N_10428,N_10313,N_10249);
nor U10429 (N_10429,N_10321,N_10326);
or U10430 (N_10430,N_10372,N_10238);
and U10431 (N_10431,N_10216,N_10214);
and U10432 (N_10432,N_10284,N_10350);
xnor U10433 (N_10433,N_10331,N_10257);
xor U10434 (N_10434,N_10355,N_10387);
xor U10435 (N_10435,N_10304,N_10246);
xor U10436 (N_10436,N_10368,N_10203);
and U10437 (N_10437,N_10374,N_10366);
and U10438 (N_10438,N_10392,N_10229);
nor U10439 (N_10439,N_10224,N_10328);
nand U10440 (N_10440,N_10341,N_10354);
and U10441 (N_10441,N_10290,N_10213);
and U10442 (N_10442,N_10258,N_10339);
or U10443 (N_10443,N_10336,N_10200);
nand U10444 (N_10444,N_10288,N_10309);
xnor U10445 (N_10445,N_10365,N_10206);
and U10446 (N_10446,N_10210,N_10394);
nand U10447 (N_10447,N_10340,N_10239);
nand U10448 (N_10448,N_10303,N_10241);
nor U10449 (N_10449,N_10294,N_10263);
nand U10450 (N_10450,N_10243,N_10363);
xnor U10451 (N_10451,N_10277,N_10305);
nor U10452 (N_10452,N_10264,N_10293);
xor U10453 (N_10453,N_10222,N_10219);
xnor U10454 (N_10454,N_10242,N_10311);
or U10455 (N_10455,N_10338,N_10201);
nor U10456 (N_10456,N_10380,N_10208);
nand U10457 (N_10457,N_10244,N_10332);
nand U10458 (N_10458,N_10352,N_10287);
xnor U10459 (N_10459,N_10324,N_10255);
nor U10460 (N_10460,N_10393,N_10378);
xor U10461 (N_10461,N_10212,N_10231);
nor U10462 (N_10462,N_10296,N_10356);
and U10463 (N_10463,N_10233,N_10232);
nor U10464 (N_10464,N_10269,N_10348);
or U10465 (N_10465,N_10329,N_10298);
xnor U10466 (N_10466,N_10376,N_10275);
nand U10467 (N_10467,N_10220,N_10276);
or U10468 (N_10468,N_10347,N_10310);
nor U10469 (N_10469,N_10337,N_10335);
and U10470 (N_10470,N_10386,N_10369);
or U10471 (N_10471,N_10322,N_10377);
nor U10472 (N_10472,N_10279,N_10252);
nor U10473 (N_10473,N_10273,N_10228);
xor U10474 (N_10474,N_10357,N_10280);
or U10475 (N_10475,N_10286,N_10317);
and U10476 (N_10476,N_10312,N_10300);
nor U10477 (N_10477,N_10282,N_10270);
or U10478 (N_10478,N_10351,N_10253);
and U10479 (N_10479,N_10245,N_10299);
or U10480 (N_10480,N_10209,N_10397);
nand U10481 (N_10481,N_10353,N_10390);
xor U10482 (N_10482,N_10362,N_10307);
nand U10483 (N_10483,N_10301,N_10308);
and U10484 (N_10484,N_10236,N_10323);
and U10485 (N_10485,N_10382,N_10259);
nor U10486 (N_10486,N_10345,N_10371);
or U10487 (N_10487,N_10399,N_10325);
or U10488 (N_10488,N_10391,N_10330);
xor U10489 (N_10489,N_10361,N_10205);
and U10490 (N_10490,N_10385,N_10367);
nor U10491 (N_10491,N_10315,N_10320);
or U10492 (N_10492,N_10383,N_10388);
nor U10493 (N_10493,N_10292,N_10281);
nand U10494 (N_10494,N_10221,N_10316);
nor U10495 (N_10495,N_10278,N_10291);
and U10496 (N_10496,N_10261,N_10271);
or U10497 (N_10497,N_10295,N_10256);
and U10498 (N_10498,N_10272,N_10379);
and U10499 (N_10499,N_10215,N_10274);
nor U10500 (N_10500,N_10214,N_10340);
or U10501 (N_10501,N_10227,N_10347);
nor U10502 (N_10502,N_10287,N_10208);
nor U10503 (N_10503,N_10367,N_10257);
xnor U10504 (N_10504,N_10288,N_10252);
and U10505 (N_10505,N_10324,N_10242);
and U10506 (N_10506,N_10373,N_10365);
and U10507 (N_10507,N_10265,N_10276);
and U10508 (N_10508,N_10350,N_10293);
nor U10509 (N_10509,N_10231,N_10213);
and U10510 (N_10510,N_10264,N_10221);
and U10511 (N_10511,N_10338,N_10300);
xor U10512 (N_10512,N_10257,N_10323);
and U10513 (N_10513,N_10211,N_10313);
nand U10514 (N_10514,N_10378,N_10260);
and U10515 (N_10515,N_10375,N_10269);
or U10516 (N_10516,N_10373,N_10287);
or U10517 (N_10517,N_10231,N_10322);
nand U10518 (N_10518,N_10318,N_10313);
or U10519 (N_10519,N_10313,N_10279);
or U10520 (N_10520,N_10365,N_10377);
xor U10521 (N_10521,N_10368,N_10357);
or U10522 (N_10522,N_10351,N_10340);
nand U10523 (N_10523,N_10316,N_10360);
and U10524 (N_10524,N_10379,N_10251);
nor U10525 (N_10525,N_10292,N_10364);
and U10526 (N_10526,N_10324,N_10214);
xnor U10527 (N_10527,N_10326,N_10267);
nand U10528 (N_10528,N_10382,N_10355);
nor U10529 (N_10529,N_10216,N_10263);
xor U10530 (N_10530,N_10230,N_10317);
or U10531 (N_10531,N_10397,N_10355);
or U10532 (N_10532,N_10267,N_10359);
and U10533 (N_10533,N_10394,N_10341);
or U10534 (N_10534,N_10233,N_10236);
nor U10535 (N_10535,N_10214,N_10206);
xnor U10536 (N_10536,N_10241,N_10285);
nand U10537 (N_10537,N_10351,N_10381);
xor U10538 (N_10538,N_10341,N_10207);
xor U10539 (N_10539,N_10286,N_10292);
or U10540 (N_10540,N_10264,N_10208);
nor U10541 (N_10541,N_10375,N_10312);
and U10542 (N_10542,N_10246,N_10309);
or U10543 (N_10543,N_10224,N_10398);
nor U10544 (N_10544,N_10236,N_10309);
xnor U10545 (N_10545,N_10368,N_10318);
and U10546 (N_10546,N_10285,N_10286);
nor U10547 (N_10547,N_10270,N_10370);
xnor U10548 (N_10548,N_10341,N_10333);
xnor U10549 (N_10549,N_10306,N_10225);
or U10550 (N_10550,N_10367,N_10218);
or U10551 (N_10551,N_10385,N_10352);
xor U10552 (N_10552,N_10274,N_10384);
and U10553 (N_10553,N_10315,N_10370);
xnor U10554 (N_10554,N_10258,N_10383);
or U10555 (N_10555,N_10381,N_10350);
or U10556 (N_10556,N_10305,N_10355);
or U10557 (N_10557,N_10272,N_10254);
and U10558 (N_10558,N_10205,N_10299);
nor U10559 (N_10559,N_10290,N_10303);
and U10560 (N_10560,N_10396,N_10242);
and U10561 (N_10561,N_10300,N_10215);
and U10562 (N_10562,N_10226,N_10396);
and U10563 (N_10563,N_10295,N_10294);
nor U10564 (N_10564,N_10383,N_10398);
nand U10565 (N_10565,N_10357,N_10217);
nand U10566 (N_10566,N_10324,N_10206);
nor U10567 (N_10567,N_10373,N_10294);
nor U10568 (N_10568,N_10392,N_10254);
nand U10569 (N_10569,N_10213,N_10361);
nor U10570 (N_10570,N_10260,N_10269);
or U10571 (N_10571,N_10398,N_10374);
nor U10572 (N_10572,N_10365,N_10343);
xor U10573 (N_10573,N_10377,N_10314);
and U10574 (N_10574,N_10389,N_10258);
and U10575 (N_10575,N_10222,N_10271);
xnor U10576 (N_10576,N_10290,N_10294);
nand U10577 (N_10577,N_10332,N_10272);
or U10578 (N_10578,N_10278,N_10264);
and U10579 (N_10579,N_10352,N_10275);
or U10580 (N_10580,N_10301,N_10268);
or U10581 (N_10581,N_10374,N_10209);
and U10582 (N_10582,N_10321,N_10222);
nor U10583 (N_10583,N_10214,N_10256);
or U10584 (N_10584,N_10233,N_10231);
xnor U10585 (N_10585,N_10286,N_10245);
or U10586 (N_10586,N_10287,N_10353);
or U10587 (N_10587,N_10217,N_10308);
xnor U10588 (N_10588,N_10223,N_10372);
nor U10589 (N_10589,N_10369,N_10288);
nand U10590 (N_10590,N_10382,N_10308);
nor U10591 (N_10591,N_10209,N_10345);
or U10592 (N_10592,N_10364,N_10283);
nand U10593 (N_10593,N_10274,N_10229);
or U10594 (N_10594,N_10393,N_10318);
nor U10595 (N_10595,N_10312,N_10204);
xor U10596 (N_10596,N_10390,N_10209);
and U10597 (N_10597,N_10247,N_10392);
nor U10598 (N_10598,N_10208,N_10396);
nand U10599 (N_10599,N_10248,N_10349);
nor U10600 (N_10600,N_10590,N_10523);
xor U10601 (N_10601,N_10505,N_10465);
xor U10602 (N_10602,N_10563,N_10527);
nor U10603 (N_10603,N_10475,N_10440);
or U10604 (N_10604,N_10506,N_10410);
nand U10605 (N_10605,N_10513,N_10538);
xnor U10606 (N_10606,N_10420,N_10443);
and U10607 (N_10607,N_10496,N_10498);
nor U10608 (N_10608,N_10437,N_10482);
or U10609 (N_10609,N_10509,N_10514);
nor U10610 (N_10610,N_10466,N_10403);
nand U10611 (N_10611,N_10419,N_10494);
xnor U10612 (N_10612,N_10438,N_10500);
and U10613 (N_10613,N_10452,N_10512);
xnor U10614 (N_10614,N_10483,N_10454);
nor U10615 (N_10615,N_10400,N_10521);
nand U10616 (N_10616,N_10518,N_10432);
nor U10617 (N_10617,N_10537,N_10455);
nor U10618 (N_10618,N_10427,N_10592);
or U10619 (N_10619,N_10453,N_10479);
nand U10620 (N_10620,N_10543,N_10407);
nand U10621 (N_10621,N_10591,N_10486);
and U10622 (N_10622,N_10573,N_10507);
nand U10623 (N_10623,N_10584,N_10426);
and U10624 (N_10624,N_10583,N_10560);
nor U10625 (N_10625,N_10588,N_10520);
or U10626 (N_10626,N_10476,N_10579);
and U10627 (N_10627,N_10534,N_10596);
nor U10628 (N_10628,N_10567,N_10499);
and U10629 (N_10629,N_10472,N_10481);
or U10630 (N_10630,N_10416,N_10434);
or U10631 (N_10631,N_10593,N_10546);
xnor U10632 (N_10632,N_10492,N_10459);
xnor U10633 (N_10633,N_10471,N_10460);
nor U10634 (N_10634,N_10418,N_10478);
xnor U10635 (N_10635,N_10473,N_10408);
or U10636 (N_10636,N_10539,N_10467);
nor U10637 (N_10637,N_10450,N_10547);
and U10638 (N_10638,N_10424,N_10530);
xor U10639 (N_10639,N_10544,N_10417);
and U10640 (N_10640,N_10557,N_10595);
nor U10641 (N_10641,N_10491,N_10565);
nand U10642 (N_10642,N_10429,N_10413);
nand U10643 (N_10643,N_10526,N_10597);
xnor U10644 (N_10644,N_10501,N_10566);
and U10645 (N_10645,N_10462,N_10562);
nor U10646 (N_10646,N_10423,N_10422);
nor U10647 (N_10647,N_10594,N_10581);
or U10648 (N_10648,N_10540,N_10556);
xnor U10649 (N_10649,N_10541,N_10405);
or U10650 (N_10650,N_10582,N_10587);
and U10651 (N_10651,N_10570,N_10542);
nand U10652 (N_10652,N_10517,N_10532);
nand U10653 (N_10653,N_10571,N_10490);
or U10654 (N_10654,N_10474,N_10554);
or U10655 (N_10655,N_10524,N_10431);
xnor U10656 (N_10656,N_10522,N_10525);
xor U10657 (N_10657,N_10568,N_10444);
xnor U10658 (N_10658,N_10430,N_10575);
xnor U10659 (N_10659,N_10464,N_10421);
nand U10660 (N_10660,N_10445,N_10458);
or U10661 (N_10661,N_10489,N_10436);
and U10662 (N_10662,N_10558,N_10577);
or U10663 (N_10663,N_10519,N_10493);
or U10664 (N_10664,N_10545,N_10516);
and U10665 (N_10665,N_10533,N_10457);
nand U10666 (N_10666,N_10511,N_10503);
nor U10667 (N_10667,N_10409,N_10548);
nor U10668 (N_10668,N_10470,N_10572);
xor U10669 (N_10669,N_10551,N_10515);
and U10670 (N_10670,N_10433,N_10497);
and U10671 (N_10671,N_10586,N_10552);
nand U10672 (N_10672,N_10488,N_10529);
nor U10673 (N_10673,N_10549,N_10480);
xnor U10674 (N_10674,N_10463,N_10448);
xnor U10675 (N_10675,N_10484,N_10406);
nand U10676 (N_10676,N_10502,N_10477);
xnor U10677 (N_10677,N_10447,N_10439);
nand U10678 (N_10678,N_10415,N_10535);
or U10679 (N_10679,N_10411,N_10441);
and U10680 (N_10680,N_10485,N_10461);
and U10681 (N_10681,N_10574,N_10508);
xnor U10682 (N_10682,N_10559,N_10561);
and U10683 (N_10683,N_10469,N_10531);
and U10684 (N_10684,N_10589,N_10528);
and U10685 (N_10685,N_10425,N_10536);
xor U10686 (N_10686,N_10504,N_10569);
or U10687 (N_10687,N_10495,N_10555);
and U10688 (N_10688,N_10401,N_10446);
and U10689 (N_10689,N_10553,N_10428);
and U10690 (N_10690,N_10578,N_10585);
or U10691 (N_10691,N_10414,N_10412);
xnor U10692 (N_10692,N_10451,N_10510);
and U10693 (N_10693,N_10435,N_10580);
xnor U10694 (N_10694,N_10404,N_10550);
nor U10695 (N_10695,N_10402,N_10576);
and U10696 (N_10696,N_10564,N_10487);
or U10697 (N_10697,N_10442,N_10449);
and U10698 (N_10698,N_10599,N_10456);
xor U10699 (N_10699,N_10468,N_10598);
or U10700 (N_10700,N_10463,N_10560);
nor U10701 (N_10701,N_10418,N_10552);
xor U10702 (N_10702,N_10533,N_10572);
xor U10703 (N_10703,N_10464,N_10507);
or U10704 (N_10704,N_10409,N_10459);
and U10705 (N_10705,N_10481,N_10412);
xnor U10706 (N_10706,N_10537,N_10418);
xnor U10707 (N_10707,N_10453,N_10529);
or U10708 (N_10708,N_10569,N_10484);
and U10709 (N_10709,N_10466,N_10409);
and U10710 (N_10710,N_10513,N_10584);
or U10711 (N_10711,N_10574,N_10415);
nor U10712 (N_10712,N_10529,N_10566);
and U10713 (N_10713,N_10423,N_10549);
and U10714 (N_10714,N_10581,N_10480);
xor U10715 (N_10715,N_10553,N_10557);
nor U10716 (N_10716,N_10427,N_10475);
or U10717 (N_10717,N_10589,N_10543);
and U10718 (N_10718,N_10591,N_10433);
xor U10719 (N_10719,N_10456,N_10446);
nor U10720 (N_10720,N_10469,N_10485);
xor U10721 (N_10721,N_10483,N_10569);
nor U10722 (N_10722,N_10599,N_10410);
or U10723 (N_10723,N_10563,N_10420);
xnor U10724 (N_10724,N_10589,N_10529);
nand U10725 (N_10725,N_10485,N_10483);
xnor U10726 (N_10726,N_10427,N_10455);
nand U10727 (N_10727,N_10408,N_10470);
nand U10728 (N_10728,N_10456,N_10463);
xor U10729 (N_10729,N_10452,N_10540);
nand U10730 (N_10730,N_10499,N_10482);
nor U10731 (N_10731,N_10414,N_10442);
xnor U10732 (N_10732,N_10566,N_10430);
nor U10733 (N_10733,N_10525,N_10596);
or U10734 (N_10734,N_10516,N_10413);
nand U10735 (N_10735,N_10576,N_10534);
nand U10736 (N_10736,N_10592,N_10538);
and U10737 (N_10737,N_10442,N_10475);
nor U10738 (N_10738,N_10458,N_10439);
and U10739 (N_10739,N_10433,N_10574);
xor U10740 (N_10740,N_10547,N_10471);
nor U10741 (N_10741,N_10495,N_10546);
xor U10742 (N_10742,N_10435,N_10544);
nand U10743 (N_10743,N_10523,N_10591);
nor U10744 (N_10744,N_10433,N_10496);
nand U10745 (N_10745,N_10463,N_10567);
or U10746 (N_10746,N_10519,N_10543);
xor U10747 (N_10747,N_10527,N_10531);
or U10748 (N_10748,N_10453,N_10592);
and U10749 (N_10749,N_10524,N_10475);
nand U10750 (N_10750,N_10552,N_10477);
or U10751 (N_10751,N_10431,N_10498);
xor U10752 (N_10752,N_10437,N_10435);
or U10753 (N_10753,N_10417,N_10535);
nand U10754 (N_10754,N_10416,N_10410);
and U10755 (N_10755,N_10417,N_10577);
nor U10756 (N_10756,N_10502,N_10512);
xor U10757 (N_10757,N_10404,N_10512);
and U10758 (N_10758,N_10550,N_10536);
xor U10759 (N_10759,N_10455,N_10419);
nor U10760 (N_10760,N_10435,N_10541);
or U10761 (N_10761,N_10426,N_10524);
or U10762 (N_10762,N_10468,N_10477);
xor U10763 (N_10763,N_10455,N_10501);
nor U10764 (N_10764,N_10435,N_10458);
nand U10765 (N_10765,N_10568,N_10518);
and U10766 (N_10766,N_10511,N_10401);
nand U10767 (N_10767,N_10491,N_10461);
nor U10768 (N_10768,N_10475,N_10456);
nor U10769 (N_10769,N_10467,N_10546);
xnor U10770 (N_10770,N_10472,N_10418);
or U10771 (N_10771,N_10428,N_10576);
nor U10772 (N_10772,N_10573,N_10471);
xor U10773 (N_10773,N_10453,N_10428);
xor U10774 (N_10774,N_10596,N_10566);
and U10775 (N_10775,N_10591,N_10555);
xor U10776 (N_10776,N_10520,N_10404);
nand U10777 (N_10777,N_10549,N_10430);
xnor U10778 (N_10778,N_10543,N_10420);
or U10779 (N_10779,N_10552,N_10553);
nand U10780 (N_10780,N_10550,N_10460);
or U10781 (N_10781,N_10576,N_10506);
nand U10782 (N_10782,N_10499,N_10498);
and U10783 (N_10783,N_10522,N_10419);
or U10784 (N_10784,N_10416,N_10539);
or U10785 (N_10785,N_10558,N_10487);
nor U10786 (N_10786,N_10586,N_10444);
xnor U10787 (N_10787,N_10546,N_10520);
nand U10788 (N_10788,N_10569,N_10527);
or U10789 (N_10789,N_10485,N_10562);
or U10790 (N_10790,N_10528,N_10464);
xor U10791 (N_10791,N_10442,N_10588);
and U10792 (N_10792,N_10555,N_10528);
xor U10793 (N_10793,N_10484,N_10480);
nor U10794 (N_10794,N_10519,N_10469);
or U10795 (N_10795,N_10491,N_10459);
nand U10796 (N_10796,N_10470,N_10458);
xnor U10797 (N_10797,N_10590,N_10573);
nor U10798 (N_10798,N_10561,N_10500);
nand U10799 (N_10799,N_10564,N_10473);
and U10800 (N_10800,N_10668,N_10604);
nor U10801 (N_10801,N_10729,N_10742);
and U10802 (N_10802,N_10623,N_10730);
and U10803 (N_10803,N_10703,N_10645);
or U10804 (N_10804,N_10601,N_10677);
and U10805 (N_10805,N_10624,N_10636);
xnor U10806 (N_10806,N_10760,N_10776);
or U10807 (N_10807,N_10631,N_10753);
nand U10808 (N_10808,N_10646,N_10744);
nand U10809 (N_10809,N_10625,N_10612);
nor U10810 (N_10810,N_10772,N_10672);
and U10811 (N_10811,N_10643,N_10711);
nand U10812 (N_10812,N_10722,N_10695);
nor U10813 (N_10813,N_10712,N_10725);
xor U10814 (N_10814,N_10609,N_10774);
nor U10815 (N_10815,N_10699,N_10716);
xor U10816 (N_10816,N_10727,N_10691);
and U10817 (N_10817,N_10634,N_10673);
nor U10818 (N_10818,N_10787,N_10683);
nor U10819 (N_10819,N_10632,N_10629);
or U10820 (N_10820,N_10641,N_10667);
and U10821 (N_10821,N_10686,N_10766);
xor U10822 (N_10822,N_10687,N_10737);
or U10823 (N_10823,N_10637,N_10782);
and U10824 (N_10824,N_10701,N_10786);
xnor U10825 (N_10825,N_10795,N_10713);
or U10826 (N_10826,N_10728,N_10648);
xnor U10827 (N_10827,N_10676,N_10666);
and U10828 (N_10828,N_10778,N_10622);
nand U10829 (N_10829,N_10651,N_10628);
nor U10830 (N_10830,N_10626,N_10747);
nor U10831 (N_10831,N_10617,N_10662);
xnor U10832 (N_10832,N_10756,N_10783);
or U10833 (N_10833,N_10755,N_10680);
nand U10834 (N_10834,N_10619,N_10799);
and U10835 (N_10835,N_10752,N_10758);
nor U10836 (N_10836,N_10750,N_10740);
nor U10837 (N_10837,N_10706,N_10763);
and U10838 (N_10838,N_10773,N_10769);
and U10839 (N_10839,N_10764,N_10649);
xor U10840 (N_10840,N_10674,N_10647);
nand U10841 (N_10841,N_10743,N_10603);
xnor U10842 (N_10842,N_10745,N_10704);
xnor U10843 (N_10843,N_10663,N_10638);
nor U10844 (N_10844,N_10633,N_10656);
nor U10845 (N_10845,N_10717,N_10757);
xor U10846 (N_10846,N_10694,N_10768);
xor U10847 (N_10847,N_10709,N_10610);
nand U10848 (N_10848,N_10790,N_10739);
xnor U10849 (N_10849,N_10690,N_10736);
and U10850 (N_10850,N_10784,N_10738);
nor U10851 (N_10851,N_10788,N_10779);
nor U10852 (N_10852,N_10731,N_10765);
and U10853 (N_10853,N_10707,N_10658);
and U10854 (N_10854,N_10660,N_10798);
or U10855 (N_10855,N_10705,N_10607);
nor U10856 (N_10856,N_10661,N_10692);
nand U10857 (N_10857,N_10767,N_10762);
and U10858 (N_10858,N_10771,N_10741);
xor U10859 (N_10859,N_10777,N_10749);
xnor U10860 (N_10860,N_10642,N_10723);
xor U10861 (N_10861,N_10791,N_10652);
nand U10862 (N_10862,N_10785,N_10748);
xnor U10863 (N_10863,N_10689,N_10697);
nand U10864 (N_10864,N_10781,N_10608);
nor U10865 (N_10865,N_10630,N_10770);
nand U10866 (N_10866,N_10669,N_10684);
xor U10867 (N_10867,N_10675,N_10635);
nand U10868 (N_10868,N_10754,N_10746);
and U10869 (N_10869,N_10644,N_10797);
xnor U10870 (N_10870,N_10715,N_10794);
or U10871 (N_10871,N_10724,N_10655);
and U10872 (N_10872,N_10780,N_10679);
nand U10873 (N_10873,N_10613,N_10714);
and U10874 (N_10874,N_10735,N_10650);
nor U10875 (N_10875,N_10702,N_10696);
or U10876 (N_10876,N_10659,N_10606);
or U10877 (N_10877,N_10733,N_10627);
or U10878 (N_10878,N_10751,N_10732);
nor U10879 (N_10879,N_10614,N_10670);
nand U10880 (N_10880,N_10718,N_10600);
nor U10881 (N_10881,N_10685,N_10621);
nor U10882 (N_10882,N_10796,N_10793);
nand U10883 (N_10883,N_10602,N_10726);
and U10884 (N_10884,N_10688,N_10639);
or U10885 (N_10885,N_10721,N_10710);
nand U10886 (N_10886,N_10789,N_10700);
and U10887 (N_10887,N_10759,N_10654);
xnor U10888 (N_10888,N_10640,N_10681);
or U10889 (N_10889,N_10618,N_10720);
xnor U10890 (N_10890,N_10611,N_10761);
xnor U10891 (N_10891,N_10775,N_10671);
and U10892 (N_10892,N_10719,N_10698);
or U10893 (N_10893,N_10615,N_10605);
and U10894 (N_10894,N_10792,N_10664);
and U10895 (N_10895,N_10665,N_10693);
nor U10896 (N_10896,N_10616,N_10682);
nand U10897 (N_10897,N_10708,N_10734);
and U10898 (N_10898,N_10653,N_10620);
and U10899 (N_10899,N_10678,N_10657);
or U10900 (N_10900,N_10788,N_10787);
or U10901 (N_10901,N_10676,N_10723);
or U10902 (N_10902,N_10754,N_10786);
nor U10903 (N_10903,N_10727,N_10626);
and U10904 (N_10904,N_10728,N_10747);
and U10905 (N_10905,N_10623,N_10626);
xnor U10906 (N_10906,N_10692,N_10707);
nor U10907 (N_10907,N_10724,N_10697);
and U10908 (N_10908,N_10608,N_10650);
and U10909 (N_10909,N_10748,N_10681);
nand U10910 (N_10910,N_10727,N_10689);
and U10911 (N_10911,N_10687,N_10602);
xor U10912 (N_10912,N_10733,N_10659);
and U10913 (N_10913,N_10748,N_10769);
nor U10914 (N_10914,N_10636,N_10775);
nand U10915 (N_10915,N_10746,N_10799);
or U10916 (N_10916,N_10677,N_10655);
or U10917 (N_10917,N_10622,N_10626);
nand U10918 (N_10918,N_10745,N_10665);
xor U10919 (N_10919,N_10791,N_10625);
xnor U10920 (N_10920,N_10754,N_10698);
and U10921 (N_10921,N_10659,N_10765);
nor U10922 (N_10922,N_10740,N_10706);
or U10923 (N_10923,N_10702,N_10706);
nor U10924 (N_10924,N_10715,N_10623);
nor U10925 (N_10925,N_10714,N_10759);
xor U10926 (N_10926,N_10724,N_10756);
xnor U10927 (N_10927,N_10768,N_10704);
and U10928 (N_10928,N_10748,N_10796);
nand U10929 (N_10929,N_10623,N_10718);
xnor U10930 (N_10930,N_10752,N_10661);
nand U10931 (N_10931,N_10677,N_10753);
nor U10932 (N_10932,N_10622,N_10701);
xnor U10933 (N_10933,N_10785,N_10660);
nor U10934 (N_10934,N_10777,N_10760);
nand U10935 (N_10935,N_10707,N_10630);
and U10936 (N_10936,N_10737,N_10761);
xnor U10937 (N_10937,N_10699,N_10705);
xnor U10938 (N_10938,N_10733,N_10717);
nand U10939 (N_10939,N_10674,N_10659);
xnor U10940 (N_10940,N_10731,N_10662);
or U10941 (N_10941,N_10634,N_10676);
and U10942 (N_10942,N_10727,N_10664);
and U10943 (N_10943,N_10755,N_10659);
xor U10944 (N_10944,N_10767,N_10665);
nor U10945 (N_10945,N_10759,N_10627);
nand U10946 (N_10946,N_10712,N_10698);
and U10947 (N_10947,N_10685,N_10624);
nor U10948 (N_10948,N_10722,N_10697);
nor U10949 (N_10949,N_10610,N_10726);
or U10950 (N_10950,N_10747,N_10697);
or U10951 (N_10951,N_10621,N_10651);
or U10952 (N_10952,N_10783,N_10623);
or U10953 (N_10953,N_10601,N_10766);
or U10954 (N_10954,N_10758,N_10611);
or U10955 (N_10955,N_10677,N_10754);
nor U10956 (N_10956,N_10706,N_10690);
or U10957 (N_10957,N_10684,N_10765);
xor U10958 (N_10958,N_10704,N_10700);
xnor U10959 (N_10959,N_10695,N_10737);
nor U10960 (N_10960,N_10673,N_10605);
nand U10961 (N_10961,N_10797,N_10689);
nor U10962 (N_10962,N_10793,N_10661);
xor U10963 (N_10963,N_10641,N_10717);
nand U10964 (N_10964,N_10626,N_10697);
xnor U10965 (N_10965,N_10694,N_10761);
or U10966 (N_10966,N_10789,N_10705);
nand U10967 (N_10967,N_10751,N_10692);
nor U10968 (N_10968,N_10643,N_10734);
or U10969 (N_10969,N_10627,N_10798);
nand U10970 (N_10970,N_10661,N_10654);
or U10971 (N_10971,N_10609,N_10750);
nand U10972 (N_10972,N_10781,N_10729);
nand U10973 (N_10973,N_10683,N_10705);
xor U10974 (N_10974,N_10691,N_10712);
nand U10975 (N_10975,N_10754,N_10799);
nor U10976 (N_10976,N_10775,N_10687);
and U10977 (N_10977,N_10703,N_10676);
xnor U10978 (N_10978,N_10772,N_10793);
or U10979 (N_10979,N_10665,N_10638);
xor U10980 (N_10980,N_10695,N_10701);
nand U10981 (N_10981,N_10760,N_10602);
and U10982 (N_10982,N_10667,N_10759);
or U10983 (N_10983,N_10639,N_10724);
xnor U10984 (N_10984,N_10602,N_10728);
or U10985 (N_10985,N_10647,N_10702);
nor U10986 (N_10986,N_10648,N_10715);
nand U10987 (N_10987,N_10737,N_10739);
nand U10988 (N_10988,N_10707,N_10625);
nand U10989 (N_10989,N_10792,N_10736);
and U10990 (N_10990,N_10617,N_10668);
and U10991 (N_10991,N_10792,N_10758);
nor U10992 (N_10992,N_10707,N_10682);
and U10993 (N_10993,N_10673,N_10782);
xor U10994 (N_10994,N_10628,N_10647);
or U10995 (N_10995,N_10624,N_10765);
nand U10996 (N_10996,N_10766,N_10616);
nand U10997 (N_10997,N_10787,N_10759);
nand U10998 (N_10998,N_10629,N_10754);
or U10999 (N_10999,N_10767,N_10639);
or U11000 (N_11000,N_10876,N_10910);
nand U11001 (N_11001,N_10951,N_10939);
and U11002 (N_11002,N_10818,N_10877);
nor U11003 (N_11003,N_10954,N_10855);
or U11004 (N_11004,N_10973,N_10995);
nor U11005 (N_11005,N_10839,N_10865);
nor U11006 (N_11006,N_10874,N_10958);
nand U11007 (N_11007,N_10940,N_10947);
and U11008 (N_11008,N_10926,N_10920);
and U11009 (N_11009,N_10864,N_10967);
nor U11010 (N_11010,N_10938,N_10982);
or U11011 (N_11011,N_10956,N_10979);
xor U11012 (N_11012,N_10883,N_10928);
nand U11013 (N_11013,N_10837,N_10870);
and U11014 (N_11014,N_10831,N_10988);
nand U11015 (N_11015,N_10853,N_10812);
nand U11016 (N_11016,N_10856,N_10801);
xnor U11017 (N_11017,N_10963,N_10850);
nor U11018 (N_11018,N_10994,N_10971);
or U11019 (N_11019,N_10843,N_10948);
nor U11020 (N_11020,N_10822,N_10815);
nand U11021 (N_11021,N_10983,N_10900);
nand U11022 (N_11022,N_10820,N_10888);
and U11023 (N_11023,N_10860,N_10962);
nor U11024 (N_11024,N_10932,N_10990);
nor U11025 (N_11025,N_10969,N_10887);
xnor U11026 (N_11026,N_10827,N_10895);
and U11027 (N_11027,N_10993,N_10985);
xnor U11028 (N_11028,N_10965,N_10824);
nor U11029 (N_11029,N_10921,N_10832);
nor U11030 (N_11030,N_10817,N_10809);
nand U11031 (N_11031,N_10924,N_10886);
or U11032 (N_11032,N_10929,N_10978);
xnor U11033 (N_11033,N_10851,N_10849);
xor U11034 (N_11034,N_10804,N_10945);
nor U11035 (N_11035,N_10953,N_10922);
or U11036 (N_11036,N_10814,N_10959);
and U11037 (N_11037,N_10961,N_10835);
and U11038 (N_11038,N_10896,N_10943);
nand U11039 (N_11039,N_10999,N_10976);
xor U11040 (N_11040,N_10934,N_10970);
and U11041 (N_11041,N_10936,N_10975);
xor U11042 (N_11042,N_10918,N_10879);
and U11043 (N_11043,N_10881,N_10977);
xnor U11044 (N_11044,N_10813,N_10841);
nor U11045 (N_11045,N_10937,N_10889);
nand U11046 (N_11046,N_10885,N_10955);
nor U11047 (N_11047,N_10823,N_10904);
nand U11048 (N_11048,N_10878,N_10927);
xor U11049 (N_11049,N_10981,N_10840);
nor U11050 (N_11050,N_10807,N_10834);
or U11051 (N_11051,N_10846,N_10857);
and U11052 (N_11052,N_10964,N_10906);
nand U11053 (N_11053,N_10960,N_10919);
nand U11054 (N_11054,N_10861,N_10903);
or U11055 (N_11055,N_10862,N_10838);
nor U11056 (N_11056,N_10829,N_10825);
or U11057 (N_11057,N_10806,N_10941);
or U11058 (N_11058,N_10957,N_10873);
and U11059 (N_11059,N_10884,N_10996);
or U11060 (N_11060,N_10803,N_10845);
nand U11061 (N_11061,N_10933,N_10826);
nand U11062 (N_11062,N_10998,N_10897);
xnor U11063 (N_11063,N_10871,N_10819);
xor U11064 (N_11064,N_10950,N_10952);
or U11065 (N_11065,N_10987,N_10890);
nand U11066 (N_11066,N_10913,N_10935);
and U11067 (N_11067,N_10867,N_10863);
nor U11068 (N_11068,N_10946,N_10836);
nand U11069 (N_11069,N_10875,N_10833);
and U11070 (N_11070,N_10872,N_10830);
and U11071 (N_11071,N_10848,N_10917);
xnor U11072 (N_11072,N_10923,N_10800);
and U11073 (N_11073,N_10925,N_10898);
and U11074 (N_11074,N_10907,N_10931);
or U11075 (N_11075,N_10802,N_10816);
and U11076 (N_11076,N_10880,N_10909);
or U11077 (N_11077,N_10810,N_10852);
or U11078 (N_11078,N_10858,N_10902);
xor U11079 (N_11079,N_10901,N_10908);
nand U11080 (N_11080,N_10869,N_10894);
and U11081 (N_11081,N_10811,N_10984);
nor U11082 (N_11082,N_10821,N_10966);
and U11083 (N_11083,N_10844,N_10997);
xor U11084 (N_11084,N_10893,N_10914);
and U11085 (N_11085,N_10944,N_10882);
nand U11086 (N_11086,N_10828,N_10989);
nand U11087 (N_11087,N_10974,N_10986);
xor U11088 (N_11088,N_10911,N_10968);
nand U11089 (N_11089,N_10942,N_10992);
nor U11090 (N_11090,N_10916,N_10972);
and U11091 (N_11091,N_10930,N_10859);
nand U11092 (N_11092,N_10912,N_10991);
nand U11093 (N_11093,N_10868,N_10949);
xor U11094 (N_11094,N_10854,N_10847);
nor U11095 (N_11095,N_10808,N_10805);
nor U11096 (N_11096,N_10899,N_10915);
xnor U11097 (N_11097,N_10891,N_10866);
or U11098 (N_11098,N_10905,N_10842);
nor U11099 (N_11099,N_10892,N_10980);
xor U11100 (N_11100,N_10845,N_10935);
nand U11101 (N_11101,N_10825,N_10899);
nand U11102 (N_11102,N_10948,N_10821);
nor U11103 (N_11103,N_10856,N_10937);
or U11104 (N_11104,N_10829,N_10813);
nand U11105 (N_11105,N_10907,N_10969);
and U11106 (N_11106,N_10952,N_10968);
nor U11107 (N_11107,N_10946,N_10834);
nor U11108 (N_11108,N_10855,N_10997);
xor U11109 (N_11109,N_10850,N_10920);
and U11110 (N_11110,N_10954,N_10850);
and U11111 (N_11111,N_10802,N_10930);
nand U11112 (N_11112,N_10987,N_10886);
nor U11113 (N_11113,N_10918,N_10954);
nor U11114 (N_11114,N_10817,N_10858);
xnor U11115 (N_11115,N_10951,N_10967);
or U11116 (N_11116,N_10860,N_10822);
xor U11117 (N_11117,N_10899,N_10913);
nand U11118 (N_11118,N_10850,N_10801);
or U11119 (N_11119,N_10961,N_10996);
nand U11120 (N_11120,N_10884,N_10807);
nor U11121 (N_11121,N_10926,N_10857);
and U11122 (N_11122,N_10958,N_10831);
and U11123 (N_11123,N_10903,N_10985);
and U11124 (N_11124,N_10894,N_10830);
nand U11125 (N_11125,N_10941,N_10809);
nor U11126 (N_11126,N_10941,N_10854);
nor U11127 (N_11127,N_10851,N_10951);
nor U11128 (N_11128,N_10905,N_10820);
or U11129 (N_11129,N_10930,N_10958);
and U11130 (N_11130,N_10904,N_10817);
or U11131 (N_11131,N_10955,N_10883);
nand U11132 (N_11132,N_10841,N_10932);
nand U11133 (N_11133,N_10934,N_10987);
or U11134 (N_11134,N_10832,N_10872);
nand U11135 (N_11135,N_10986,N_10975);
or U11136 (N_11136,N_10955,N_10800);
nor U11137 (N_11137,N_10965,N_10892);
and U11138 (N_11138,N_10968,N_10874);
nand U11139 (N_11139,N_10851,N_10995);
and U11140 (N_11140,N_10964,N_10919);
xnor U11141 (N_11141,N_10814,N_10836);
xor U11142 (N_11142,N_10858,N_10892);
nand U11143 (N_11143,N_10845,N_10817);
nand U11144 (N_11144,N_10866,N_10837);
xnor U11145 (N_11145,N_10861,N_10870);
nand U11146 (N_11146,N_10957,N_10975);
nand U11147 (N_11147,N_10999,N_10817);
nor U11148 (N_11148,N_10819,N_10800);
nand U11149 (N_11149,N_10910,N_10843);
or U11150 (N_11150,N_10845,N_10911);
or U11151 (N_11151,N_10805,N_10924);
nor U11152 (N_11152,N_10911,N_10866);
and U11153 (N_11153,N_10868,N_10893);
xnor U11154 (N_11154,N_10909,N_10913);
nand U11155 (N_11155,N_10979,N_10967);
and U11156 (N_11156,N_10961,N_10848);
nor U11157 (N_11157,N_10816,N_10935);
xnor U11158 (N_11158,N_10897,N_10859);
or U11159 (N_11159,N_10882,N_10996);
nor U11160 (N_11160,N_10967,N_10989);
nand U11161 (N_11161,N_10901,N_10818);
and U11162 (N_11162,N_10978,N_10891);
nor U11163 (N_11163,N_10881,N_10833);
xor U11164 (N_11164,N_10815,N_10823);
nand U11165 (N_11165,N_10944,N_10914);
or U11166 (N_11166,N_10808,N_10821);
xor U11167 (N_11167,N_10955,N_10983);
or U11168 (N_11168,N_10991,N_10903);
and U11169 (N_11169,N_10900,N_10889);
nor U11170 (N_11170,N_10895,N_10946);
and U11171 (N_11171,N_10973,N_10919);
or U11172 (N_11172,N_10801,N_10820);
nor U11173 (N_11173,N_10883,N_10898);
nor U11174 (N_11174,N_10914,N_10983);
nand U11175 (N_11175,N_10823,N_10950);
nand U11176 (N_11176,N_10846,N_10972);
xor U11177 (N_11177,N_10988,N_10920);
and U11178 (N_11178,N_10815,N_10920);
nor U11179 (N_11179,N_10840,N_10987);
or U11180 (N_11180,N_10988,N_10999);
nor U11181 (N_11181,N_10844,N_10939);
nand U11182 (N_11182,N_10830,N_10882);
nand U11183 (N_11183,N_10859,N_10800);
and U11184 (N_11184,N_10808,N_10907);
nor U11185 (N_11185,N_10817,N_10807);
xor U11186 (N_11186,N_10810,N_10893);
xor U11187 (N_11187,N_10899,N_10971);
or U11188 (N_11188,N_10899,N_10874);
and U11189 (N_11189,N_10944,N_10814);
nand U11190 (N_11190,N_10877,N_10914);
and U11191 (N_11191,N_10961,N_10883);
or U11192 (N_11192,N_10851,N_10971);
or U11193 (N_11193,N_10958,N_10962);
and U11194 (N_11194,N_10815,N_10911);
xnor U11195 (N_11195,N_10882,N_10801);
xor U11196 (N_11196,N_10991,N_10804);
xor U11197 (N_11197,N_10820,N_10941);
nor U11198 (N_11198,N_10864,N_10963);
or U11199 (N_11199,N_10955,N_10893);
and U11200 (N_11200,N_11035,N_11136);
nor U11201 (N_11201,N_11193,N_11062);
nand U11202 (N_11202,N_11078,N_11155);
xnor U11203 (N_11203,N_11099,N_11080);
and U11204 (N_11204,N_11024,N_11060);
xor U11205 (N_11205,N_11145,N_11076);
nand U11206 (N_11206,N_11146,N_11142);
nor U11207 (N_11207,N_11166,N_11088);
nand U11208 (N_11208,N_11064,N_11017);
and U11209 (N_11209,N_11175,N_11137);
nor U11210 (N_11210,N_11037,N_11039);
or U11211 (N_11211,N_11028,N_11143);
nand U11212 (N_11212,N_11161,N_11114);
xor U11213 (N_11213,N_11052,N_11069);
nor U11214 (N_11214,N_11048,N_11007);
nand U11215 (N_11215,N_11051,N_11125);
nand U11216 (N_11216,N_11185,N_11092);
and U11217 (N_11217,N_11027,N_11004);
xnor U11218 (N_11218,N_11077,N_11176);
nand U11219 (N_11219,N_11107,N_11187);
xor U11220 (N_11220,N_11041,N_11101);
nor U11221 (N_11221,N_11119,N_11124);
or U11222 (N_11222,N_11083,N_11163);
xor U11223 (N_11223,N_11116,N_11192);
and U11224 (N_11224,N_11105,N_11094);
nor U11225 (N_11225,N_11082,N_11063);
nand U11226 (N_11226,N_11043,N_11065);
nand U11227 (N_11227,N_11093,N_11072);
xor U11228 (N_11228,N_11046,N_11188);
nand U11229 (N_11229,N_11170,N_11144);
nor U11230 (N_11230,N_11133,N_11001);
and U11231 (N_11231,N_11122,N_11067);
and U11232 (N_11232,N_11014,N_11130);
xnor U11233 (N_11233,N_11073,N_11047);
nor U11234 (N_11234,N_11061,N_11159);
or U11235 (N_11235,N_11059,N_11167);
or U11236 (N_11236,N_11070,N_11013);
xnor U11237 (N_11237,N_11154,N_11045);
nor U11238 (N_11238,N_11085,N_11050);
xnor U11239 (N_11239,N_11174,N_11126);
and U11240 (N_11240,N_11008,N_11058);
or U11241 (N_11241,N_11178,N_11110);
or U11242 (N_11242,N_11010,N_11148);
xnor U11243 (N_11243,N_11079,N_11115);
or U11244 (N_11244,N_11030,N_11168);
or U11245 (N_11245,N_11102,N_11003);
or U11246 (N_11246,N_11016,N_11151);
nand U11247 (N_11247,N_11029,N_11180);
and U11248 (N_11248,N_11123,N_11135);
xnor U11249 (N_11249,N_11086,N_11177);
or U11250 (N_11250,N_11087,N_11111);
nand U11251 (N_11251,N_11054,N_11040);
or U11252 (N_11252,N_11131,N_11056);
xnor U11253 (N_11253,N_11173,N_11129);
nor U11254 (N_11254,N_11150,N_11036);
nor U11255 (N_11255,N_11127,N_11128);
nor U11256 (N_11256,N_11165,N_11186);
or U11257 (N_11257,N_11147,N_11183);
nand U11258 (N_11258,N_11112,N_11171);
and U11259 (N_11259,N_11162,N_11021);
and U11260 (N_11260,N_11108,N_11172);
and U11261 (N_11261,N_11199,N_11197);
and U11262 (N_11262,N_11002,N_11113);
and U11263 (N_11263,N_11194,N_11149);
and U11264 (N_11264,N_11139,N_11023);
or U11265 (N_11265,N_11015,N_11089);
nor U11266 (N_11266,N_11057,N_11009);
nand U11267 (N_11267,N_11032,N_11179);
or U11268 (N_11268,N_11121,N_11025);
nor U11269 (N_11269,N_11000,N_11097);
or U11270 (N_11270,N_11081,N_11095);
or U11271 (N_11271,N_11138,N_11134);
and U11272 (N_11272,N_11038,N_11006);
and U11273 (N_11273,N_11049,N_11091);
nand U11274 (N_11274,N_11164,N_11169);
nand U11275 (N_11275,N_11053,N_11132);
xor U11276 (N_11276,N_11157,N_11153);
xnor U11277 (N_11277,N_11100,N_11019);
xnor U11278 (N_11278,N_11189,N_11141);
xnor U11279 (N_11279,N_11117,N_11022);
and U11280 (N_11280,N_11104,N_11042);
xor U11281 (N_11281,N_11074,N_11106);
and U11282 (N_11282,N_11034,N_11195);
nand U11283 (N_11283,N_11190,N_11031);
nand U11284 (N_11284,N_11075,N_11071);
and U11285 (N_11285,N_11012,N_11191);
and U11286 (N_11286,N_11011,N_11118);
or U11287 (N_11287,N_11152,N_11160);
and U11288 (N_11288,N_11184,N_11005);
and U11289 (N_11289,N_11196,N_11158);
xnor U11290 (N_11290,N_11044,N_11103);
nor U11291 (N_11291,N_11020,N_11098);
xnor U11292 (N_11292,N_11018,N_11026);
nor U11293 (N_11293,N_11120,N_11182);
nand U11294 (N_11294,N_11140,N_11156);
or U11295 (N_11295,N_11090,N_11055);
or U11296 (N_11296,N_11066,N_11198);
or U11297 (N_11297,N_11096,N_11033);
xnor U11298 (N_11298,N_11181,N_11109);
xnor U11299 (N_11299,N_11068,N_11084);
xor U11300 (N_11300,N_11044,N_11084);
nand U11301 (N_11301,N_11094,N_11041);
nor U11302 (N_11302,N_11038,N_11123);
nor U11303 (N_11303,N_11077,N_11064);
nor U11304 (N_11304,N_11029,N_11113);
nor U11305 (N_11305,N_11072,N_11083);
nand U11306 (N_11306,N_11019,N_11146);
nand U11307 (N_11307,N_11044,N_11138);
xor U11308 (N_11308,N_11078,N_11150);
or U11309 (N_11309,N_11181,N_11015);
and U11310 (N_11310,N_11145,N_11132);
or U11311 (N_11311,N_11019,N_11010);
nand U11312 (N_11312,N_11154,N_11024);
xor U11313 (N_11313,N_11139,N_11077);
and U11314 (N_11314,N_11004,N_11062);
xnor U11315 (N_11315,N_11136,N_11189);
xnor U11316 (N_11316,N_11162,N_11112);
and U11317 (N_11317,N_11126,N_11155);
and U11318 (N_11318,N_11076,N_11102);
xor U11319 (N_11319,N_11150,N_11155);
xor U11320 (N_11320,N_11087,N_11192);
or U11321 (N_11321,N_11010,N_11150);
xor U11322 (N_11322,N_11169,N_11114);
and U11323 (N_11323,N_11037,N_11051);
and U11324 (N_11324,N_11138,N_11005);
xnor U11325 (N_11325,N_11122,N_11111);
nand U11326 (N_11326,N_11187,N_11071);
nor U11327 (N_11327,N_11025,N_11053);
or U11328 (N_11328,N_11034,N_11002);
or U11329 (N_11329,N_11103,N_11048);
nor U11330 (N_11330,N_11103,N_11004);
nor U11331 (N_11331,N_11026,N_11044);
nand U11332 (N_11332,N_11021,N_11140);
nor U11333 (N_11333,N_11016,N_11162);
nor U11334 (N_11334,N_11101,N_11075);
and U11335 (N_11335,N_11043,N_11126);
and U11336 (N_11336,N_11140,N_11010);
xor U11337 (N_11337,N_11075,N_11111);
xor U11338 (N_11338,N_11111,N_11092);
xnor U11339 (N_11339,N_11198,N_11134);
xnor U11340 (N_11340,N_11066,N_11068);
nand U11341 (N_11341,N_11085,N_11059);
xor U11342 (N_11342,N_11116,N_11171);
nor U11343 (N_11343,N_11065,N_11041);
or U11344 (N_11344,N_11166,N_11034);
nor U11345 (N_11345,N_11108,N_11103);
and U11346 (N_11346,N_11041,N_11090);
and U11347 (N_11347,N_11114,N_11087);
nor U11348 (N_11348,N_11172,N_11049);
xor U11349 (N_11349,N_11084,N_11147);
or U11350 (N_11350,N_11173,N_11106);
or U11351 (N_11351,N_11050,N_11127);
or U11352 (N_11352,N_11012,N_11158);
or U11353 (N_11353,N_11003,N_11098);
xor U11354 (N_11354,N_11060,N_11012);
nor U11355 (N_11355,N_11026,N_11053);
nor U11356 (N_11356,N_11136,N_11139);
or U11357 (N_11357,N_11024,N_11018);
nand U11358 (N_11358,N_11151,N_11079);
xor U11359 (N_11359,N_11167,N_11039);
and U11360 (N_11360,N_11019,N_11183);
and U11361 (N_11361,N_11111,N_11120);
nand U11362 (N_11362,N_11109,N_11069);
nor U11363 (N_11363,N_11089,N_11014);
or U11364 (N_11364,N_11099,N_11024);
xor U11365 (N_11365,N_11015,N_11085);
nand U11366 (N_11366,N_11167,N_11135);
xnor U11367 (N_11367,N_11197,N_11027);
and U11368 (N_11368,N_11112,N_11142);
and U11369 (N_11369,N_11190,N_11126);
nor U11370 (N_11370,N_11072,N_11050);
nor U11371 (N_11371,N_11199,N_11180);
nor U11372 (N_11372,N_11193,N_11033);
xor U11373 (N_11373,N_11056,N_11115);
nor U11374 (N_11374,N_11144,N_11027);
xor U11375 (N_11375,N_11124,N_11039);
nor U11376 (N_11376,N_11004,N_11021);
or U11377 (N_11377,N_11022,N_11134);
xnor U11378 (N_11378,N_11152,N_11093);
or U11379 (N_11379,N_11054,N_11167);
xor U11380 (N_11380,N_11186,N_11069);
xnor U11381 (N_11381,N_11052,N_11025);
and U11382 (N_11382,N_11103,N_11119);
and U11383 (N_11383,N_11093,N_11170);
and U11384 (N_11384,N_11194,N_11181);
nand U11385 (N_11385,N_11168,N_11163);
nand U11386 (N_11386,N_11178,N_11101);
and U11387 (N_11387,N_11198,N_11186);
and U11388 (N_11388,N_11034,N_11180);
xor U11389 (N_11389,N_11148,N_11028);
and U11390 (N_11390,N_11125,N_11004);
nor U11391 (N_11391,N_11170,N_11118);
or U11392 (N_11392,N_11009,N_11090);
nand U11393 (N_11393,N_11021,N_11101);
or U11394 (N_11394,N_11154,N_11040);
or U11395 (N_11395,N_11118,N_11143);
nand U11396 (N_11396,N_11046,N_11088);
nand U11397 (N_11397,N_11172,N_11148);
or U11398 (N_11398,N_11089,N_11057);
or U11399 (N_11399,N_11099,N_11015);
xor U11400 (N_11400,N_11361,N_11393);
nand U11401 (N_11401,N_11386,N_11286);
nor U11402 (N_11402,N_11292,N_11347);
and U11403 (N_11403,N_11256,N_11360);
nand U11404 (N_11404,N_11259,N_11341);
nor U11405 (N_11405,N_11253,N_11217);
nand U11406 (N_11406,N_11282,N_11306);
xor U11407 (N_11407,N_11260,N_11235);
xor U11408 (N_11408,N_11350,N_11241);
nand U11409 (N_11409,N_11240,N_11381);
or U11410 (N_11410,N_11336,N_11303);
xnor U11411 (N_11411,N_11375,N_11296);
and U11412 (N_11412,N_11294,N_11378);
xnor U11413 (N_11413,N_11279,N_11211);
xor U11414 (N_11414,N_11273,N_11288);
or U11415 (N_11415,N_11221,N_11359);
nand U11416 (N_11416,N_11210,N_11280);
and U11417 (N_11417,N_11356,N_11213);
nor U11418 (N_11418,N_11325,N_11377);
xor U11419 (N_11419,N_11388,N_11307);
or U11420 (N_11420,N_11236,N_11340);
nand U11421 (N_11421,N_11209,N_11371);
or U11422 (N_11422,N_11365,N_11281);
or U11423 (N_11423,N_11216,N_11278);
nor U11424 (N_11424,N_11249,N_11284);
nor U11425 (N_11425,N_11215,N_11298);
nor U11426 (N_11426,N_11372,N_11364);
nand U11427 (N_11427,N_11353,N_11232);
xnor U11428 (N_11428,N_11313,N_11200);
nand U11429 (N_11429,N_11342,N_11276);
and U11430 (N_11430,N_11206,N_11223);
xor U11431 (N_11431,N_11351,N_11320);
and U11432 (N_11432,N_11255,N_11376);
xor U11433 (N_11433,N_11308,N_11326);
nand U11434 (N_11434,N_11318,N_11335);
nor U11435 (N_11435,N_11315,N_11290);
xor U11436 (N_11436,N_11390,N_11330);
or U11437 (N_11437,N_11258,N_11266);
xor U11438 (N_11438,N_11310,N_11245);
nor U11439 (N_11439,N_11251,N_11287);
and U11440 (N_11440,N_11323,N_11369);
and U11441 (N_11441,N_11384,N_11225);
xnor U11442 (N_11442,N_11385,N_11202);
and U11443 (N_11443,N_11319,N_11379);
or U11444 (N_11444,N_11231,N_11366);
nand U11445 (N_11445,N_11222,N_11337);
nor U11446 (N_11446,N_11274,N_11218);
or U11447 (N_11447,N_11305,N_11238);
or U11448 (N_11448,N_11208,N_11264);
or U11449 (N_11449,N_11399,N_11397);
nor U11450 (N_11450,N_11345,N_11301);
xor U11451 (N_11451,N_11242,N_11243);
nor U11452 (N_11452,N_11237,N_11270);
xnor U11453 (N_11453,N_11297,N_11394);
nand U11454 (N_11454,N_11387,N_11229);
nor U11455 (N_11455,N_11391,N_11374);
xnor U11456 (N_11456,N_11309,N_11267);
nand U11457 (N_11457,N_11214,N_11254);
nand U11458 (N_11458,N_11263,N_11327);
nand U11459 (N_11459,N_11220,N_11212);
nor U11460 (N_11460,N_11205,N_11349);
nand U11461 (N_11461,N_11333,N_11291);
nor U11462 (N_11462,N_11227,N_11275);
xnor U11463 (N_11463,N_11239,N_11244);
or U11464 (N_11464,N_11373,N_11314);
nand U11465 (N_11465,N_11396,N_11334);
nor U11466 (N_11466,N_11317,N_11271);
nor U11467 (N_11467,N_11201,N_11219);
or U11468 (N_11468,N_11261,N_11207);
nor U11469 (N_11469,N_11324,N_11382);
nand U11470 (N_11470,N_11289,N_11269);
xnor U11471 (N_11471,N_11304,N_11344);
nand U11472 (N_11472,N_11203,N_11250);
nand U11473 (N_11473,N_11247,N_11362);
or U11474 (N_11474,N_11300,N_11338);
xor U11475 (N_11475,N_11257,N_11228);
nor U11476 (N_11476,N_11368,N_11346);
and U11477 (N_11477,N_11265,N_11252);
nor U11478 (N_11478,N_11230,N_11262);
or U11479 (N_11479,N_11358,N_11383);
nor U11480 (N_11480,N_11299,N_11339);
or U11481 (N_11481,N_11380,N_11348);
xor U11482 (N_11482,N_11224,N_11295);
and U11483 (N_11483,N_11248,N_11355);
xor U11484 (N_11484,N_11322,N_11392);
nand U11485 (N_11485,N_11321,N_11398);
nor U11486 (N_11486,N_11389,N_11283);
nand U11487 (N_11487,N_11285,N_11302);
or U11488 (N_11488,N_11352,N_11246);
nor U11489 (N_11489,N_11328,N_11316);
xnor U11490 (N_11490,N_11357,N_11332);
or U11491 (N_11491,N_11395,N_11370);
and U11492 (N_11492,N_11226,N_11311);
xnor U11493 (N_11493,N_11354,N_11268);
xnor U11494 (N_11494,N_11234,N_11329);
nor U11495 (N_11495,N_11312,N_11272);
xor U11496 (N_11496,N_11293,N_11343);
nor U11497 (N_11497,N_11331,N_11277);
nand U11498 (N_11498,N_11233,N_11363);
or U11499 (N_11499,N_11204,N_11367);
nor U11500 (N_11500,N_11256,N_11238);
xor U11501 (N_11501,N_11305,N_11302);
xnor U11502 (N_11502,N_11336,N_11276);
and U11503 (N_11503,N_11322,N_11328);
and U11504 (N_11504,N_11211,N_11234);
nand U11505 (N_11505,N_11268,N_11386);
xnor U11506 (N_11506,N_11368,N_11347);
or U11507 (N_11507,N_11219,N_11373);
nand U11508 (N_11508,N_11222,N_11381);
xnor U11509 (N_11509,N_11391,N_11236);
and U11510 (N_11510,N_11307,N_11396);
nor U11511 (N_11511,N_11260,N_11245);
nand U11512 (N_11512,N_11234,N_11268);
and U11513 (N_11513,N_11284,N_11323);
nand U11514 (N_11514,N_11221,N_11237);
nand U11515 (N_11515,N_11367,N_11345);
nor U11516 (N_11516,N_11298,N_11263);
nor U11517 (N_11517,N_11266,N_11361);
or U11518 (N_11518,N_11316,N_11272);
or U11519 (N_11519,N_11238,N_11268);
and U11520 (N_11520,N_11278,N_11220);
and U11521 (N_11521,N_11388,N_11291);
xor U11522 (N_11522,N_11261,N_11235);
or U11523 (N_11523,N_11279,N_11301);
xnor U11524 (N_11524,N_11270,N_11241);
nand U11525 (N_11525,N_11380,N_11280);
nor U11526 (N_11526,N_11339,N_11381);
xor U11527 (N_11527,N_11395,N_11369);
and U11528 (N_11528,N_11376,N_11214);
or U11529 (N_11529,N_11286,N_11271);
or U11530 (N_11530,N_11364,N_11279);
xnor U11531 (N_11531,N_11309,N_11381);
or U11532 (N_11532,N_11356,N_11375);
or U11533 (N_11533,N_11331,N_11254);
and U11534 (N_11534,N_11396,N_11286);
nand U11535 (N_11535,N_11205,N_11249);
xnor U11536 (N_11536,N_11260,N_11350);
and U11537 (N_11537,N_11327,N_11239);
or U11538 (N_11538,N_11360,N_11236);
nor U11539 (N_11539,N_11288,N_11213);
nand U11540 (N_11540,N_11299,N_11376);
xor U11541 (N_11541,N_11289,N_11327);
nor U11542 (N_11542,N_11227,N_11206);
or U11543 (N_11543,N_11241,N_11318);
nor U11544 (N_11544,N_11306,N_11366);
xnor U11545 (N_11545,N_11331,N_11212);
and U11546 (N_11546,N_11247,N_11380);
nand U11547 (N_11547,N_11365,N_11392);
xor U11548 (N_11548,N_11315,N_11366);
and U11549 (N_11549,N_11224,N_11213);
xor U11550 (N_11550,N_11231,N_11392);
nor U11551 (N_11551,N_11291,N_11263);
nand U11552 (N_11552,N_11212,N_11261);
or U11553 (N_11553,N_11335,N_11282);
and U11554 (N_11554,N_11255,N_11232);
or U11555 (N_11555,N_11220,N_11394);
xor U11556 (N_11556,N_11224,N_11360);
xor U11557 (N_11557,N_11257,N_11372);
nand U11558 (N_11558,N_11251,N_11228);
or U11559 (N_11559,N_11232,N_11235);
or U11560 (N_11560,N_11285,N_11391);
and U11561 (N_11561,N_11304,N_11352);
nor U11562 (N_11562,N_11259,N_11246);
and U11563 (N_11563,N_11308,N_11247);
xnor U11564 (N_11564,N_11308,N_11246);
xnor U11565 (N_11565,N_11234,N_11250);
xnor U11566 (N_11566,N_11241,N_11323);
xor U11567 (N_11567,N_11248,N_11239);
xnor U11568 (N_11568,N_11300,N_11250);
nand U11569 (N_11569,N_11247,N_11343);
nand U11570 (N_11570,N_11277,N_11337);
xor U11571 (N_11571,N_11284,N_11234);
and U11572 (N_11572,N_11244,N_11233);
nor U11573 (N_11573,N_11267,N_11269);
or U11574 (N_11574,N_11264,N_11258);
or U11575 (N_11575,N_11290,N_11322);
and U11576 (N_11576,N_11291,N_11298);
nor U11577 (N_11577,N_11246,N_11379);
xor U11578 (N_11578,N_11391,N_11211);
nand U11579 (N_11579,N_11334,N_11228);
nand U11580 (N_11580,N_11262,N_11255);
or U11581 (N_11581,N_11339,N_11325);
nand U11582 (N_11582,N_11299,N_11288);
nand U11583 (N_11583,N_11283,N_11364);
nand U11584 (N_11584,N_11312,N_11243);
xnor U11585 (N_11585,N_11200,N_11263);
xor U11586 (N_11586,N_11205,N_11283);
xor U11587 (N_11587,N_11307,N_11301);
nand U11588 (N_11588,N_11384,N_11243);
nor U11589 (N_11589,N_11245,N_11334);
or U11590 (N_11590,N_11371,N_11286);
or U11591 (N_11591,N_11346,N_11356);
nand U11592 (N_11592,N_11222,N_11335);
or U11593 (N_11593,N_11234,N_11275);
nand U11594 (N_11594,N_11344,N_11303);
nand U11595 (N_11595,N_11262,N_11210);
and U11596 (N_11596,N_11338,N_11381);
or U11597 (N_11597,N_11203,N_11284);
or U11598 (N_11598,N_11394,N_11347);
nor U11599 (N_11599,N_11297,N_11350);
or U11600 (N_11600,N_11445,N_11576);
or U11601 (N_11601,N_11526,N_11435);
and U11602 (N_11602,N_11592,N_11582);
nor U11603 (N_11603,N_11413,N_11595);
xnor U11604 (N_11604,N_11579,N_11523);
or U11605 (N_11605,N_11454,N_11598);
xnor U11606 (N_11606,N_11492,N_11418);
nor U11607 (N_11607,N_11476,N_11572);
nor U11608 (N_11608,N_11486,N_11457);
nor U11609 (N_11609,N_11458,N_11519);
xnor U11610 (N_11610,N_11412,N_11470);
and U11611 (N_11611,N_11522,N_11439);
nand U11612 (N_11612,N_11567,N_11585);
or U11613 (N_11613,N_11527,N_11540);
nor U11614 (N_11614,N_11436,N_11544);
nand U11615 (N_11615,N_11449,N_11531);
or U11616 (N_11616,N_11483,N_11501);
or U11617 (N_11617,N_11403,N_11533);
nand U11618 (N_11618,N_11584,N_11546);
or U11619 (N_11619,N_11485,N_11562);
and U11620 (N_11620,N_11547,N_11437);
xor U11621 (N_11621,N_11524,N_11409);
or U11622 (N_11622,N_11539,N_11575);
or U11623 (N_11623,N_11462,N_11477);
or U11624 (N_11624,N_11565,N_11407);
nor U11625 (N_11625,N_11441,N_11591);
xnor U11626 (N_11626,N_11472,N_11488);
xor U11627 (N_11627,N_11507,N_11559);
nor U11628 (N_11628,N_11447,N_11528);
and U11629 (N_11629,N_11543,N_11459);
nor U11630 (N_11630,N_11594,N_11564);
xor U11631 (N_11631,N_11479,N_11534);
nor U11632 (N_11632,N_11471,N_11597);
and U11633 (N_11633,N_11513,N_11495);
or U11634 (N_11634,N_11431,N_11506);
xnor U11635 (N_11635,N_11434,N_11566);
or U11636 (N_11636,N_11429,N_11573);
nor U11637 (N_11637,N_11535,N_11463);
nor U11638 (N_11638,N_11411,N_11550);
nand U11639 (N_11639,N_11590,N_11424);
nor U11640 (N_11640,N_11503,N_11549);
nand U11641 (N_11641,N_11551,N_11474);
or U11642 (N_11642,N_11490,N_11465);
and U11643 (N_11643,N_11475,N_11599);
or U11644 (N_11644,N_11442,N_11410);
xor U11645 (N_11645,N_11473,N_11538);
xnor U11646 (N_11646,N_11560,N_11421);
xor U11647 (N_11647,N_11510,N_11419);
nand U11648 (N_11648,N_11545,N_11593);
nand U11649 (N_11649,N_11499,N_11433);
nand U11650 (N_11650,N_11541,N_11496);
nor U11651 (N_11651,N_11512,N_11516);
and U11652 (N_11652,N_11466,N_11481);
or U11653 (N_11653,N_11570,N_11468);
nand U11654 (N_11654,N_11569,N_11583);
xor U11655 (N_11655,N_11461,N_11518);
and U11656 (N_11656,N_11525,N_11498);
nor U11657 (N_11657,N_11405,N_11430);
or U11658 (N_11658,N_11558,N_11581);
xor U11659 (N_11659,N_11505,N_11408);
nand U11660 (N_11660,N_11511,N_11440);
nand U11661 (N_11661,N_11467,N_11456);
xnor U11662 (N_11662,N_11552,N_11432);
nor U11663 (N_11663,N_11554,N_11548);
or U11664 (N_11664,N_11482,N_11469);
and U11665 (N_11665,N_11464,N_11571);
and U11666 (N_11666,N_11423,N_11553);
or U11667 (N_11667,N_11452,N_11530);
and U11668 (N_11668,N_11406,N_11416);
or U11669 (N_11669,N_11497,N_11460);
nor U11670 (N_11670,N_11508,N_11450);
xor U11671 (N_11671,N_11537,N_11577);
xnor U11672 (N_11672,N_11420,N_11444);
xor U11673 (N_11673,N_11509,N_11517);
nor U11674 (N_11674,N_11400,N_11532);
xor U11675 (N_11675,N_11453,N_11451);
xor U11676 (N_11676,N_11568,N_11493);
and U11677 (N_11677,N_11448,N_11402);
nor U11678 (N_11678,N_11529,N_11489);
and U11679 (N_11679,N_11589,N_11438);
nor U11680 (N_11680,N_11484,N_11487);
xor U11681 (N_11681,N_11427,N_11563);
nand U11682 (N_11682,N_11491,N_11426);
and U11683 (N_11683,N_11494,N_11561);
and U11684 (N_11684,N_11514,N_11521);
xor U11685 (N_11685,N_11455,N_11443);
and U11686 (N_11686,N_11580,N_11500);
or U11687 (N_11687,N_11588,N_11596);
or U11688 (N_11688,N_11555,N_11414);
nor U11689 (N_11689,N_11578,N_11415);
xor U11690 (N_11690,N_11504,N_11446);
or U11691 (N_11691,N_11557,N_11428);
or U11692 (N_11692,N_11422,N_11542);
nand U11693 (N_11693,N_11586,N_11574);
nand U11694 (N_11694,N_11417,N_11401);
xnor U11695 (N_11695,N_11556,N_11520);
nand U11696 (N_11696,N_11404,N_11587);
nand U11697 (N_11697,N_11502,N_11536);
nor U11698 (N_11698,N_11425,N_11515);
and U11699 (N_11699,N_11478,N_11480);
nand U11700 (N_11700,N_11472,N_11504);
or U11701 (N_11701,N_11563,N_11494);
and U11702 (N_11702,N_11557,N_11443);
nand U11703 (N_11703,N_11435,N_11479);
and U11704 (N_11704,N_11453,N_11484);
xnor U11705 (N_11705,N_11480,N_11449);
or U11706 (N_11706,N_11403,N_11432);
xor U11707 (N_11707,N_11455,N_11429);
or U11708 (N_11708,N_11427,N_11575);
or U11709 (N_11709,N_11495,N_11509);
nand U11710 (N_11710,N_11493,N_11494);
xnor U11711 (N_11711,N_11586,N_11464);
and U11712 (N_11712,N_11418,N_11588);
xor U11713 (N_11713,N_11516,N_11440);
or U11714 (N_11714,N_11597,N_11480);
and U11715 (N_11715,N_11578,N_11472);
nor U11716 (N_11716,N_11431,N_11501);
or U11717 (N_11717,N_11492,N_11585);
and U11718 (N_11718,N_11478,N_11584);
and U11719 (N_11719,N_11475,N_11474);
and U11720 (N_11720,N_11553,N_11460);
nor U11721 (N_11721,N_11429,N_11486);
nor U11722 (N_11722,N_11467,N_11503);
nand U11723 (N_11723,N_11423,N_11434);
xnor U11724 (N_11724,N_11411,N_11487);
or U11725 (N_11725,N_11427,N_11504);
nand U11726 (N_11726,N_11509,N_11472);
nand U11727 (N_11727,N_11449,N_11485);
and U11728 (N_11728,N_11540,N_11566);
nor U11729 (N_11729,N_11450,N_11563);
and U11730 (N_11730,N_11470,N_11557);
and U11731 (N_11731,N_11497,N_11556);
nor U11732 (N_11732,N_11455,N_11541);
and U11733 (N_11733,N_11478,N_11486);
nand U11734 (N_11734,N_11403,N_11561);
and U11735 (N_11735,N_11557,N_11595);
xor U11736 (N_11736,N_11470,N_11561);
and U11737 (N_11737,N_11441,N_11418);
or U11738 (N_11738,N_11400,N_11485);
and U11739 (N_11739,N_11524,N_11416);
and U11740 (N_11740,N_11477,N_11564);
xnor U11741 (N_11741,N_11517,N_11531);
nor U11742 (N_11742,N_11567,N_11572);
nor U11743 (N_11743,N_11487,N_11586);
or U11744 (N_11744,N_11595,N_11424);
xor U11745 (N_11745,N_11524,N_11461);
or U11746 (N_11746,N_11515,N_11414);
nand U11747 (N_11747,N_11479,N_11525);
or U11748 (N_11748,N_11548,N_11531);
nor U11749 (N_11749,N_11455,N_11433);
xor U11750 (N_11750,N_11540,N_11541);
nor U11751 (N_11751,N_11588,N_11595);
nand U11752 (N_11752,N_11427,N_11572);
nand U11753 (N_11753,N_11587,N_11407);
or U11754 (N_11754,N_11486,N_11430);
and U11755 (N_11755,N_11565,N_11527);
xnor U11756 (N_11756,N_11568,N_11505);
and U11757 (N_11757,N_11538,N_11492);
nand U11758 (N_11758,N_11477,N_11412);
nor U11759 (N_11759,N_11443,N_11441);
xor U11760 (N_11760,N_11553,N_11402);
or U11761 (N_11761,N_11472,N_11564);
nor U11762 (N_11762,N_11506,N_11583);
nand U11763 (N_11763,N_11495,N_11455);
xor U11764 (N_11764,N_11455,N_11479);
xnor U11765 (N_11765,N_11532,N_11411);
or U11766 (N_11766,N_11529,N_11536);
or U11767 (N_11767,N_11531,N_11448);
nand U11768 (N_11768,N_11496,N_11513);
nor U11769 (N_11769,N_11569,N_11577);
nor U11770 (N_11770,N_11512,N_11541);
nor U11771 (N_11771,N_11490,N_11556);
nand U11772 (N_11772,N_11465,N_11470);
xnor U11773 (N_11773,N_11544,N_11580);
or U11774 (N_11774,N_11443,N_11461);
or U11775 (N_11775,N_11599,N_11554);
xnor U11776 (N_11776,N_11483,N_11455);
nor U11777 (N_11777,N_11540,N_11551);
nor U11778 (N_11778,N_11588,N_11598);
nand U11779 (N_11779,N_11595,N_11554);
nor U11780 (N_11780,N_11401,N_11466);
nand U11781 (N_11781,N_11559,N_11541);
nand U11782 (N_11782,N_11460,N_11569);
nor U11783 (N_11783,N_11404,N_11581);
and U11784 (N_11784,N_11409,N_11430);
or U11785 (N_11785,N_11525,N_11516);
nor U11786 (N_11786,N_11453,N_11498);
xnor U11787 (N_11787,N_11402,N_11472);
nand U11788 (N_11788,N_11465,N_11486);
nand U11789 (N_11789,N_11548,N_11461);
nand U11790 (N_11790,N_11557,N_11484);
and U11791 (N_11791,N_11508,N_11461);
nand U11792 (N_11792,N_11419,N_11554);
nor U11793 (N_11793,N_11515,N_11484);
nand U11794 (N_11794,N_11465,N_11505);
xor U11795 (N_11795,N_11538,N_11470);
xor U11796 (N_11796,N_11521,N_11528);
and U11797 (N_11797,N_11508,N_11556);
and U11798 (N_11798,N_11472,N_11556);
nand U11799 (N_11799,N_11479,N_11420);
nor U11800 (N_11800,N_11760,N_11645);
nand U11801 (N_11801,N_11790,N_11796);
xnor U11802 (N_11802,N_11666,N_11723);
nor U11803 (N_11803,N_11747,N_11683);
xnor U11804 (N_11804,N_11636,N_11756);
nor U11805 (N_11805,N_11719,N_11694);
nand U11806 (N_11806,N_11651,N_11758);
and U11807 (N_11807,N_11707,N_11622);
nand U11808 (N_11808,N_11712,N_11721);
nor U11809 (N_11809,N_11684,N_11686);
nand U11810 (N_11810,N_11662,N_11609);
nand U11811 (N_11811,N_11687,N_11616);
nand U11812 (N_11812,N_11613,N_11744);
nor U11813 (N_11813,N_11799,N_11665);
or U11814 (N_11814,N_11634,N_11675);
nand U11815 (N_11815,N_11720,N_11786);
nor U11816 (N_11816,N_11788,N_11695);
nand U11817 (N_11817,N_11601,N_11604);
xnor U11818 (N_11818,N_11745,N_11726);
nor U11819 (N_11819,N_11728,N_11681);
nand U11820 (N_11820,N_11737,N_11739);
and U11821 (N_11821,N_11753,N_11668);
and U11822 (N_11822,N_11653,N_11759);
and U11823 (N_11823,N_11638,N_11690);
and U11824 (N_11824,N_11671,N_11669);
or U11825 (N_11825,N_11658,N_11659);
nor U11826 (N_11826,N_11794,N_11632);
nor U11827 (N_11827,N_11688,N_11764);
nor U11828 (N_11828,N_11614,N_11680);
or U11829 (N_11829,N_11674,N_11773);
or U11830 (N_11830,N_11623,N_11702);
nand U11831 (N_11831,N_11761,N_11615);
or U11832 (N_11832,N_11672,N_11742);
nand U11833 (N_11833,N_11693,N_11648);
nor U11834 (N_11834,N_11787,N_11682);
and U11835 (N_11835,N_11768,N_11673);
nand U11836 (N_11836,N_11780,N_11631);
nand U11837 (N_11837,N_11637,N_11706);
nand U11838 (N_11838,N_11733,N_11661);
and U11839 (N_11839,N_11797,N_11704);
nor U11840 (N_11840,N_11600,N_11646);
and U11841 (N_11841,N_11722,N_11779);
or U11842 (N_11842,N_11696,N_11718);
nand U11843 (N_11843,N_11767,N_11713);
xor U11844 (N_11844,N_11677,N_11743);
nand U11845 (N_11845,N_11748,N_11617);
nand U11846 (N_11846,N_11778,N_11732);
or U11847 (N_11847,N_11627,N_11765);
nand U11848 (N_11848,N_11749,N_11620);
xor U11849 (N_11849,N_11624,N_11716);
xnor U11850 (N_11850,N_11628,N_11736);
xor U11851 (N_11851,N_11642,N_11678);
and U11852 (N_11852,N_11660,N_11751);
nor U11853 (N_11853,N_11689,N_11698);
or U11854 (N_11854,N_11781,N_11782);
nor U11855 (N_11855,N_11750,N_11776);
nor U11856 (N_11856,N_11643,N_11650);
and U11857 (N_11857,N_11606,N_11731);
nor U11858 (N_11858,N_11644,N_11783);
xor U11859 (N_11859,N_11798,N_11766);
and U11860 (N_11860,N_11676,N_11785);
xnor U11861 (N_11861,N_11639,N_11626);
nand U11862 (N_11862,N_11618,N_11649);
and U11863 (N_11863,N_11667,N_11777);
or U11864 (N_11864,N_11755,N_11709);
nand U11865 (N_11865,N_11629,N_11770);
xor U11866 (N_11866,N_11714,N_11602);
nand U11867 (N_11867,N_11738,N_11697);
nor U11868 (N_11868,N_11611,N_11652);
xnor U11869 (N_11869,N_11717,N_11699);
and U11870 (N_11870,N_11656,N_11774);
nand U11871 (N_11871,N_11663,N_11740);
xnor U11872 (N_11872,N_11710,N_11730);
nand U11873 (N_11873,N_11692,N_11610);
xor U11874 (N_11874,N_11795,N_11685);
xnor U11875 (N_11875,N_11734,N_11705);
xor U11876 (N_11876,N_11746,N_11700);
nand U11877 (N_11877,N_11727,N_11654);
and U11878 (N_11878,N_11625,N_11612);
nand U11879 (N_11879,N_11752,N_11715);
nand U11880 (N_11880,N_11703,N_11605);
xnor U11881 (N_11881,N_11641,N_11793);
or U11882 (N_11882,N_11711,N_11691);
or U11883 (N_11883,N_11608,N_11619);
nor U11884 (N_11884,N_11708,N_11679);
xnor U11885 (N_11885,N_11769,N_11635);
xor U11886 (N_11886,N_11757,N_11724);
nor U11887 (N_11887,N_11657,N_11784);
and U11888 (N_11888,N_11633,N_11607);
or U11889 (N_11889,N_11789,N_11763);
nor U11890 (N_11890,N_11792,N_11725);
xor U11891 (N_11891,N_11762,N_11664);
xnor U11892 (N_11892,N_11791,N_11735);
nor U11893 (N_11893,N_11647,N_11621);
and U11894 (N_11894,N_11772,N_11630);
nand U11895 (N_11895,N_11771,N_11741);
and U11896 (N_11896,N_11640,N_11775);
nor U11897 (N_11897,N_11701,N_11754);
and U11898 (N_11898,N_11729,N_11655);
nand U11899 (N_11899,N_11670,N_11603);
nor U11900 (N_11900,N_11706,N_11772);
xnor U11901 (N_11901,N_11699,N_11789);
nand U11902 (N_11902,N_11710,N_11613);
xor U11903 (N_11903,N_11797,N_11795);
xnor U11904 (N_11904,N_11625,N_11774);
nor U11905 (N_11905,N_11699,N_11741);
nand U11906 (N_11906,N_11704,N_11632);
nand U11907 (N_11907,N_11692,N_11731);
nand U11908 (N_11908,N_11694,N_11737);
nor U11909 (N_11909,N_11754,N_11668);
nand U11910 (N_11910,N_11716,N_11623);
nor U11911 (N_11911,N_11761,N_11707);
or U11912 (N_11912,N_11700,N_11627);
xor U11913 (N_11913,N_11708,N_11643);
xor U11914 (N_11914,N_11788,N_11628);
nand U11915 (N_11915,N_11714,N_11665);
or U11916 (N_11916,N_11659,N_11656);
or U11917 (N_11917,N_11791,N_11797);
nand U11918 (N_11918,N_11620,N_11601);
nand U11919 (N_11919,N_11683,N_11664);
and U11920 (N_11920,N_11758,N_11775);
xnor U11921 (N_11921,N_11643,N_11791);
nand U11922 (N_11922,N_11745,N_11637);
xor U11923 (N_11923,N_11694,N_11629);
xor U11924 (N_11924,N_11692,N_11658);
or U11925 (N_11925,N_11615,N_11793);
or U11926 (N_11926,N_11723,N_11784);
nor U11927 (N_11927,N_11654,N_11645);
nand U11928 (N_11928,N_11775,N_11613);
xor U11929 (N_11929,N_11603,N_11695);
or U11930 (N_11930,N_11636,N_11715);
xor U11931 (N_11931,N_11619,N_11615);
nor U11932 (N_11932,N_11733,N_11783);
or U11933 (N_11933,N_11687,N_11778);
and U11934 (N_11934,N_11688,N_11623);
or U11935 (N_11935,N_11669,N_11642);
nor U11936 (N_11936,N_11615,N_11643);
nand U11937 (N_11937,N_11749,N_11781);
or U11938 (N_11938,N_11689,N_11628);
nand U11939 (N_11939,N_11794,N_11743);
nand U11940 (N_11940,N_11616,N_11633);
nor U11941 (N_11941,N_11650,N_11780);
nor U11942 (N_11942,N_11638,N_11662);
or U11943 (N_11943,N_11652,N_11746);
nand U11944 (N_11944,N_11742,N_11632);
nor U11945 (N_11945,N_11684,N_11688);
xor U11946 (N_11946,N_11711,N_11739);
nor U11947 (N_11947,N_11793,N_11772);
and U11948 (N_11948,N_11778,N_11639);
or U11949 (N_11949,N_11673,N_11601);
and U11950 (N_11950,N_11779,N_11754);
xnor U11951 (N_11951,N_11701,N_11643);
and U11952 (N_11952,N_11793,N_11636);
or U11953 (N_11953,N_11617,N_11747);
and U11954 (N_11954,N_11798,N_11786);
nor U11955 (N_11955,N_11799,N_11747);
xnor U11956 (N_11956,N_11663,N_11644);
nor U11957 (N_11957,N_11628,N_11793);
nor U11958 (N_11958,N_11655,N_11760);
nand U11959 (N_11959,N_11691,N_11728);
nor U11960 (N_11960,N_11702,N_11789);
xnor U11961 (N_11961,N_11691,N_11793);
nor U11962 (N_11962,N_11780,N_11749);
nor U11963 (N_11963,N_11666,N_11792);
and U11964 (N_11964,N_11736,N_11763);
xor U11965 (N_11965,N_11781,N_11684);
or U11966 (N_11966,N_11659,N_11687);
nand U11967 (N_11967,N_11758,N_11682);
xor U11968 (N_11968,N_11781,N_11692);
or U11969 (N_11969,N_11710,N_11695);
or U11970 (N_11970,N_11741,N_11715);
and U11971 (N_11971,N_11623,N_11625);
nor U11972 (N_11972,N_11649,N_11614);
xor U11973 (N_11973,N_11680,N_11741);
nand U11974 (N_11974,N_11754,N_11603);
xor U11975 (N_11975,N_11737,N_11731);
nand U11976 (N_11976,N_11653,N_11651);
or U11977 (N_11977,N_11712,N_11701);
and U11978 (N_11978,N_11607,N_11785);
xor U11979 (N_11979,N_11705,N_11616);
nand U11980 (N_11980,N_11792,N_11771);
nand U11981 (N_11981,N_11618,N_11660);
nand U11982 (N_11982,N_11624,N_11651);
xnor U11983 (N_11983,N_11749,N_11642);
nand U11984 (N_11984,N_11640,N_11753);
and U11985 (N_11985,N_11738,N_11601);
and U11986 (N_11986,N_11705,N_11642);
nand U11987 (N_11987,N_11772,N_11667);
nand U11988 (N_11988,N_11780,N_11621);
or U11989 (N_11989,N_11795,N_11638);
xnor U11990 (N_11990,N_11691,N_11694);
or U11991 (N_11991,N_11716,N_11630);
xor U11992 (N_11992,N_11710,N_11610);
or U11993 (N_11993,N_11624,N_11718);
xnor U11994 (N_11994,N_11791,N_11777);
or U11995 (N_11995,N_11691,N_11710);
nor U11996 (N_11996,N_11627,N_11782);
xnor U11997 (N_11997,N_11637,N_11623);
or U11998 (N_11998,N_11639,N_11710);
nor U11999 (N_11999,N_11647,N_11684);
xor U12000 (N_12000,N_11866,N_11978);
nor U12001 (N_12001,N_11805,N_11895);
and U12002 (N_12002,N_11951,N_11896);
nand U12003 (N_12003,N_11920,N_11986);
nor U12004 (N_12004,N_11946,N_11898);
and U12005 (N_12005,N_11862,N_11891);
or U12006 (N_12006,N_11999,N_11808);
and U12007 (N_12007,N_11987,N_11817);
nor U12008 (N_12008,N_11965,N_11988);
nor U12009 (N_12009,N_11809,N_11838);
and U12010 (N_12010,N_11997,N_11923);
and U12011 (N_12011,N_11868,N_11875);
nor U12012 (N_12012,N_11913,N_11959);
nor U12013 (N_12013,N_11921,N_11881);
nand U12014 (N_12014,N_11833,N_11827);
nand U12015 (N_12015,N_11812,N_11856);
or U12016 (N_12016,N_11874,N_11929);
nand U12017 (N_12017,N_11907,N_11815);
and U12018 (N_12018,N_11937,N_11814);
nor U12019 (N_12019,N_11905,N_11962);
and U12020 (N_12020,N_11983,N_11925);
and U12021 (N_12021,N_11903,N_11943);
and U12022 (N_12022,N_11841,N_11956);
and U12023 (N_12023,N_11870,N_11961);
nor U12024 (N_12024,N_11900,N_11849);
and U12025 (N_12025,N_11919,N_11975);
or U12026 (N_12026,N_11971,N_11974);
and U12027 (N_12027,N_11911,N_11835);
and U12028 (N_12028,N_11947,N_11816);
and U12029 (N_12029,N_11878,N_11801);
nand U12030 (N_12030,N_11939,N_11928);
nor U12031 (N_12031,N_11982,N_11940);
and U12032 (N_12032,N_11877,N_11955);
nor U12033 (N_12033,N_11932,N_11984);
or U12034 (N_12034,N_11897,N_11885);
nand U12035 (N_12035,N_11848,N_11800);
nor U12036 (N_12036,N_11996,N_11845);
or U12037 (N_12037,N_11821,N_11926);
or U12038 (N_12038,N_11843,N_11853);
or U12039 (N_12039,N_11938,N_11882);
nor U12040 (N_12040,N_11976,N_11852);
xor U12041 (N_12041,N_11886,N_11910);
and U12042 (N_12042,N_11872,N_11917);
nor U12043 (N_12043,N_11831,N_11859);
or U12044 (N_12044,N_11930,N_11847);
nand U12045 (N_12045,N_11850,N_11989);
or U12046 (N_12046,N_11820,N_11924);
nor U12047 (N_12047,N_11963,N_11966);
and U12048 (N_12048,N_11941,N_11828);
and U12049 (N_12049,N_11980,N_11804);
nand U12050 (N_12050,N_11889,N_11837);
nor U12051 (N_12051,N_11927,N_11888);
nand U12052 (N_12052,N_11811,N_11918);
nor U12053 (N_12053,N_11873,N_11969);
and U12054 (N_12054,N_11880,N_11855);
xor U12055 (N_12055,N_11899,N_11964);
nor U12056 (N_12056,N_11842,N_11883);
nand U12057 (N_12057,N_11960,N_11942);
or U12058 (N_12058,N_11884,N_11807);
nand U12059 (N_12059,N_11931,N_11892);
nor U12060 (N_12060,N_11967,N_11981);
nand U12061 (N_12061,N_11819,N_11936);
nand U12062 (N_12062,N_11934,N_11972);
nand U12063 (N_12063,N_11826,N_11912);
or U12064 (N_12064,N_11863,N_11968);
nor U12065 (N_12065,N_11832,N_11970);
xnor U12066 (N_12066,N_11858,N_11864);
or U12067 (N_12067,N_11901,N_11952);
nor U12068 (N_12068,N_11893,N_11949);
and U12069 (N_12069,N_11958,N_11876);
or U12070 (N_12070,N_11829,N_11890);
nand U12071 (N_12071,N_11806,N_11979);
or U12072 (N_12072,N_11825,N_11953);
or U12073 (N_12073,N_11908,N_11813);
xnor U12074 (N_12074,N_11865,N_11857);
nand U12075 (N_12075,N_11973,N_11945);
xor U12076 (N_12076,N_11948,N_11935);
or U12077 (N_12077,N_11957,N_11802);
or U12078 (N_12078,N_11810,N_11902);
and U12079 (N_12079,N_11985,N_11922);
nor U12080 (N_12080,N_11995,N_11887);
nand U12081 (N_12081,N_11909,N_11914);
or U12082 (N_12082,N_11822,N_11830);
nand U12083 (N_12083,N_11991,N_11916);
or U12084 (N_12084,N_11836,N_11992);
xor U12085 (N_12085,N_11834,N_11854);
and U12086 (N_12086,N_11803,N_11867);
nor U12087 (N_12087,N_11906,N_11861);
xnor U12088 (N_12088,N_11839,N_11894);
xor U12089 (N_12089,N_11851,N_11844);
nand U12090 (N_12090,N_11818,N_11904);
or U12091 (N_12091,N_11840,N_11860);
nor U12092 (N_12092,N_11824,N_11823);
nand U12093 (N_12093,N_11879,N_11954);
nor U12094 (N_12094,N_11993,N_11915);
nand U12095 (N_12095,N_11871,N_11846);
and U12096 (N_12096,N_11944,N_11977);
xor U12097 (N_12097,N_11869,N_11933);
or U12098 (N_12098,N_11994,N_11950);
nor U12099 (N_12099,N_11998,N_11990);
nor U12100 (N_12100,N_11888,N_11897);
xor U12101 (N_12101,N_11839,N_11987);
nand U12102 (N_12102,N_11917,N_11951);
or U12103 (N_12103,N_11942,N_11919);
nor U12104 (N_12104,N_11824,N_11809);
and U12105 (N_12105,N_11869,N_11874);
nand U12106 (N_12106,N_11991,N_11842);
and U12107 (N_12107,N_11988,N_11887);
and U12108 (N_12108,N_11942,N_11902);
and U12109 (N_12109,N_11926,N_11847);
and U12110 (N_12110,N_11916,N_11974);
and U12111 (N_12111,N_11976,N_11928);
nor U12112 (N_12112,N_11951,N_11900);
or U12113 (N_12113,N_11852,N_11985);
and U12114 (N_12114,N_11981,N_11987);
or U12115 (N_12115,N_11872,N_11843);
or U12116 (N_12116,N_11868,N_11890);
nor U12117 (N_12117,N_11803,N_11875);
nand U12118 (N_12118,N_11951,N_11869);
nand U12119 (N_12119,N_11848,N_11940);
or U12120 (N_12120,N_11905,N_11843);
nand U12121 (N_12121,N_11990,N_11919);
and U12122 (N_12122,N_11999,N_11895);
nor U12123 (N_12123,N_11981,N_11917);
xor U12124 (N_12124,N_11967,N_11847);
and U12125 (N_12125,N_11857,N_11812);
and U12126 (N_12126,N_11821,N_11951);
xor U12127 (N_12127,N_11867,N_11968);
xnor U12128 (N_12128,N_11913,N_11988);
or U12129 (N_12129,N_11847,N_11987);
or U12130 (N_12130,N_11879,N_11801);
nor U12131 (N_12131,N_11911,N_11878);
xnor U12132 (N_12132,N_11967,N_11815);
xor U12133 (N_12133,N_11865,N_11968);
and U12134 (N_12134,N_11930,N_11898);
xor U12135 (N_12135,N_11851,N_11969);
nand U12136 (N_12136,N_11832,N_11955);
or U12137 (N_12137,N_11893,N_11971);
and U12138 (N_12138,N_11874,N_11916);
xnor U12139 (N_12139,N_11944,N_11893);
or U12140 (N_12140,N_11856,N_11895);
or U12141 (N_12141,N_11956,N_11877);
or U12142 (N_12142,N_11847,N_11981);
and U12143 (N_12143,N_11922,N_11950);
and U12144 (N_12144,N_11802,N_11950);
nor U12145 (N_12145,N_11964,N_11987);
and U12146 (N_12146,N_11982,N_11844);
or U12147 (N_12147,N_11932,N_11809);
xnor U12148 (N_12148,N_11993,N_11884);
xnor U12149 (N_12149,N_11881,N_11975);
and U12150 (N_12150,N_11971,N_11848);
or U12151 (N_12151,N_11932,N_11893);
and U12152 (N_12152,N_11827,N_11971);
and U12153 (N_12153,N_11900,N_11914);
nor U12154 (N_12154,N_11914,N_11917);
xor U12155 (N_12155,N_11864,N_11854);
and U12156 (N_12156,N_11823,N_11806);
and U12157 (N_12157,N_11985,N_11946);
or U12158 (N_12158,N_11803,N_11947);
and U12159 (N_12159,N_11904,N_11837);
nand U12160 (N_12160,N_11885,N_11945);
xnor U12161 (N_12161,N_11986,N_11927);
and U12162 (N_12162,N_11911,N_11822);
nand U12163 (N_12163,N_11943,N_11891);
xor U12164 (N_12164,N_11895,N_11845);
and U12165 (N_12165,N_11818,N_11807);
nand U12166 (N_12166,N_11969,N_11940);
or U12167 (N_12167,N_11945,N_11934);
nand U12168 (N_12168,N_11807,N_11921);
nand U12169 (N_12169,N_11856,N_11838);
xor U12170 (N_12170,N_11997,N_11804);
nor U12171 (N_12171,N_11893,N_11870);
nand U12172 (N_12172,N_11939,N_11998);
xnor U12173 (N_12173,N_11868,N_11904);
and U12174 (N_12174,N_11825,N_11827);
and U12175 (N_12175,N_11823,N_11897);
nand U12176 (N_12176,N_11861,N_11899);
or U12177 (N_12177,N_11892,N_11935);
nor U12178 (N_12178,N_11801,N_11865);
xor U12179 (N_12179,N_11838,N_11841);
and U12180 (N_12180,N_11966,N_11981);
nand U12181 (N_12181,N_11840,N_11963);
xor U12182 (N_12182,N_11920,N_11848);
nor U12183 (N_12183,N_11929,N_11889);
or U12184 (N_12184,N_11927,N_11892);
and U12185 (N_12185,N_11875,N_11843);
nand U12186 (N_12186,N_11816,N_11905);
or U12187 (N_12187,N_11937,N_11824);
and U12188 (N_12188,N_11876,N_11806);
nor U12189 (N_12189,N_11941,N_11864);
xor U12190 (N_12190,N_11891,N_11887);
or U12191 (N_12191,N_11840,N_11834);
xnor U12192 (N_12192,N_11827,N_11829);
nand U12193 (N_12193,N_11838,N_11881);
or U12194 (N_12194,N_11942,N_11830);
nand U12195 (N_12195,N_11880,N_11831);
nor U12196 (N_12196,N_11829,N_11997);
nor U12197 (N_12197,N_11853,N_11915);
nor U12198 (N_12198,N_11821,N_11937);
xor U12199 (N_12199,N_11974,N_11982);
xor U12200 (N_12200,N_12010,N_12083);
nand U12201 (N_12201,N_12086,N_12152);
or U12202 (N_12202,N_12077,N_12003);
or U12203 (N_12203,N_12111,N_12139);
nand U12204 (N_12204,N_12035,N_12093);
nand U12205 (N_12205,N_12098,N_12020);
nand U12206 (N_12206,N_12120,N_12079);
xnor U12207 (N_12207,N_12121,N_12102);
nand U12208 (N_12208,N_12017,N_12150);
xnor U12209 (N_12209,N_12054,N_12162);
xor U12210 (N_12210,N_12199,N_12067);
nand U12211 (N_12211,N_12059,N_12024);
or U12212 (N_12212,N_12005,N_12151);
and U12213 (N_12213,N_12049,N_12160);
and U12214 (N_12214,N_12131,N_12084);
xnor U12215 (N_12215,N_12047,N_12088);
and U12216 (N_12216,N_12155,N_12008);
or U12217 (N_12217,N_12133,N_12068);
xor U12218 (N_12218,N_12195,N_12104);
or U12219 (N_12219,N_12148,N_12128);
and U12220 (N_12220,N_12082,N_12075);
and U12221 (N_12221,N_12180,N_12168);
xnor U12222 (N_12222,N_12112,N_12033);
or U12223 (N_12223,N_12137,N_12187);
nand U12224 (N_12224,N_12129,N_12080);
and U12225 (N_12225,N_12081,N_12193);
or U12226 (N_12226,N_12127,N_12073);
nor U12227 (N_12227,N_12040,N_12135);
nand U12228 (N_12228,N_12028,N_12132);
and U12229 (N_12229,N_12190,N_12048);
nand U12230 (N_12230,N_12140,N_12026);
xnor U12231 (N_12231,N_12101,N_12114);
nor U12232 (N_12232,N_12058,N_12146);
nand U12233 (N_12233,N_12034,N_12175);
nand U12234 (N_12234,N_12108,N_12167);
xnor U12235 (N_12235,N_12041,N_12012);
nand U12236 (N_12236,N_12069,N_12092);
nor U12237 (N_12237,N_12061,N_12060);
nand U12238 (N_12238,N_12094,N_12030);
or U12239 (N_12239,N_12043,N_12057);
or U12240 (N_12240,N_12134,N_12182);
or U12241 (N_12241,N_12161,N_12087);
xor U12242 (N_12242,N_12066,N_12025);
nand U12243 (N_12243,N_12157,N_12042);
or U12244 (N_12244,N_12116,N_12095);
nor U12245 (N_12245,N_12109,N_12100);
or U12246 (N_12246,N_12145,N_12021);
nor U12247 (N_12247,N_12013,N_12178);
nand U12248 (N_12248,N_12007,N_12044);
nor U12249 (N_12249,N_12027,N_12181);
nand U12250 (N_12250,N_12141,N_12019);
and U12251 (N_12251,N_12176,N_12183);
or U12252 (N_12252,N_12110,N_12117);
nor U12253 (N_12253,N_12179,N_12016);
nor U12254 (N_12254,N_12072,N_12062);
or U12255 (N_12255,N_12053,N_12001);
nor U12256 (N_12256,N_12136,N_12125);
and U12257 (N_12257,N_12031,N_12159);
nor U12258 (N_12258,N_12188,N_12197);
xnor U12259 (N_12259,N_12039,N_12038);
and U12260 (N_12260,N_12126,N_12052);
nor U12261 (N_12261,N_12163,N_12189);
nor U12262 (N_12262,N_12147,N_12011);
and U12263 (N_12263,N_12124,N_12085);
nand U12264 (N_12264,N_12165,N_12154);
or U12265 (N_12265,N_12130,N_12196);
xnor U12266 (N_12266,N_12036,N_12169);
nand U12267 (N_12267,N_12091,N_12064);
nor U12268 (N_12268,N_12023,N_12096);
xnor U12269 (N_12269,N_12050,N_12123);
xor U12270 (N_12270,N_12122,N_12097);
and U12271 (N_12271,N_12090,N_12004);
xnor U12272 (N_12272,N_12006,N_12078);
or U12273 (N_12273,N_12143,N_12149);
xnor U12274 (N_12274,N_12099,N_12173);
or U12275 (N_12275,N_12118,N_12037);
xor U12276 (N_12276,N_12051,N_12065);
and U12277 (N_12277,N_12174,N_12103);
or U12278 (N_12278,N_12171,N_12071);
and U12279 (N_12279,N_12089,N_12009);
nor U12280 (N_12280,N_12113,N_12115);
and U12281 (N_12281,N_12002,N_12166);
or U12282 (N_12282,N_12185,N_12032);
or U12283 (N_12283,N_12074,N_12194);
xnor U12284 (N_12284,N_12177,N_12184);
and U12285 (N_12285,N_12198,N_12045);
or U12286 (N_12286,N_12170,N_12144);
nand U12287 (N_12287,N_12063,N_12172);
and U12288 (N_12288,N_12156,N_12055);
and U12289 (N_12289,N_12022,N_12076);
and U12290 (N_12290,N_12119,N_12164);
or U12291 (N_12291,N_12158,N_12070);
xnor U12292 (N_12292,N_12106,N_12191);
and U12293 (N_12293,N_12105,N_12046);
nand U12294 (N_12294,N_12018,N_12153);
nor U12295 (N_12295,N_12014,N_12000);
or U12296 (N_12296,N_12192,N_12142);
and U12297 (N_12297,N_12107,N_12029);
nor U12298 (N_12298,N_12138,N_12186);
xnor U12299 (N_12299,N_12015,N_12056);
and U12300 (N_12300,N_12004,N_12052);
and U12301 (N_12301,N_12198,N_12065);
nor U12302 (N_12302,N_12149,N_12012);
nand U12303 (N_12303,N_12104,N_12138);
nand U12304 (N_12304,N_12023,N_12069);
and U12305 (N_12305,N_12113,N_12093);
nor U12306 (N_12306,N_12055,N_12163);
nor U12307 (N_12307,N_12096,N_12127);
and U12308 (N_12308,N_12016,N_12109);
and U12309 (N_12309,N_12127,N_12008);
xor U12310 (N_12310,N_12184,N_12193);
xnor U12311 (N_12311,N_12149,N_12162);
nand U12312 (N_12312,N_12119,N_12099);
and U12313 (N_12313,N_12182,N_12022);
nand U12314 (N_12314,N_12047,N_12129);
xnor U12315 (N_12315,N_12141,N_12126);
xor U12316 (N_12316,N_12143,N_12080);
nand U12317 (N_12317,N_12114,N_12039);
nor U12318 (N_12318,N_12188,N_12147);
nor U12319 (N_12319,N_12093,N_12166);
nand U12320 (N_12320,N_12135,N_12016);
and U12321 (N_12321,N_12193,N_12114);
nand U12322 (N_12322,N_12197,N_12107);
nor U12323 (N_12323,N_12061,N_12088);
and U12324 (N_12324,N_12157,N_12067);
or U12325 (N_12325,N_12024,N_12152);
nand U12326 (N_12326,N_12042,N_12088);
nor U12327 (N_12327,N_12107,N_12121);
nor U12328 (N_12328,N_12181,N_12071);
or U12329 (N_12329,N_12023,N_12137);
and U12330 (N_12330,N_12097,N_12148);
xor U12331 (N_12331,N_12077,N_12004);
nand U12332 (N_12332,N_12156,N_12090);
or U12333 (N_12333,N_12109,N_12195);
or U12334 (N_12334,N_12113,N_12089);
or U12335 (N_12335,N_12061,N_12040);
xnor U12336 (N_12336,N_12024,N_12038);
nor U12337 (N_12337,N_12027,N_12149);
nor U12338 (N_12338,N_12043,N_12069);
xor U12339 (N_12339,N_12099,N_12192);
or U12340 (N_12340,N_12054,N_12181);
or U12341 (N_12341,N_12000,N_12087);
nand U12342 (N_12342,N_12107,N_12028);
xor U12343 (N_12343,N_12010,N_12003);
and U12344 (N_12344,N_12000,N_12187);
or U12345 (N_12345,N_12000,N_12004);
xnor U12346 (N_12346,N_12084,N_12106);
xnor U12347 (N_12347,N_12152,N_12167);
nor U12348 (N_12348,N_12115,N_12028);
xnor U12349 (N_12349,N_12073,N_12060);
nor U12350 (N_12350,N_12026,N_12005);
xnor U12351 (N_12351,N_12013,N_12038);
or U12352 (N_12352,N_12011,N_12171);
nor U12353 (N_12353,N_12014,N_12166);
or U12354 (N_12354,N_12111,N_12045);
and U12355 (N_12355,N_12044,N_12118);
nand U12356 (N_12356,N_12005,N_12190);
or U12357 (N_12357,N_12188,N_12168);
nand U12358 (N_12358,N_12014,N_12003);
or U12359 (N_12359,N_12086,N_12112);
xnor U12360 (N_12360,N_12178,N_12175);
xnor U12361 (N_12361,N_12181,N_12024);
nor U12362 (N_12362,N_12094,N_12078);
and U12363 (N_12363,N_12069,N_12004);
or U12364 (N_12364,N_12079,N_12189);
nand U12365 (N_12365,N_12105,N_12057);
nor U12366 (N_12366,N_12045,N_12098);
or U12367 (N_12367,N_12038,N_12163);
and U12368 (N_12368,N_12176,N_12032);
xor U12369 (N_12369,N_12139,N_12085);
xnor U12370 (N_12370,N_12020,N_12003);
nor U12371 (N_12371,N_12145,N_12050);
nor U12372 (N_12372,N_12177,N_12044);
or U12373 (N_12373,N_12171,N_12076);
nand U12374 (N_12374,N_12186,N_12106);
nand U12375 (N_12375,N_12102,N_12023);
or U12376 (N_12376,N_12012,N_12115);
nor U12377 (N_12377,N_12115,N_12010);
and U12378 (N_12378,N_12086,N_12055);
xor U12379 (N_12379,N_12029,N_12055);
and U12380 (N_12380,N_12058,N_12134);
nand U12381 (N_12381,N_12185,N_12167);
or U12382 (N_12382,N_12068,N_12107);
and U12383 (N_12383,N_12137,N_12018);
nand U12384 (N_12384,N_12028,N_12053);
nor U12385 (N_12385,N_12136,N_12186);
and U12386 (N_12386,N_12184,N_12188);
or U12387 (N_12387,N_12038,N_12084);
or U12388 (N_12388,N_12088,N_12129);
xor U12389 (N_12389,N_12120,N_12193);
nor U12390 (N_12390,N_12043,N_12197);
or U12391 (N_12391,N_12192,N_12065);
nor U12392 (N_12392,N_12083,N_12099);
and U12393 (N_12393,N_12099,N_12197);
nor U12394 (N_12394,N_12103,N_12049);
xnor U12395 (N_12395,N_12181,N_12127);
xor U12396 (N_12396,N_12189,N_12129);
nand U12397 (N_12397,N_12197,N_12050);
nor U12398 (N_12398,N_12052,N_12085);
nor U12399 (N_12399,N_12075,N_12091);
or U12400 (N_12400,N_12327,N_12287);
and U12401 (N_12401,N_12253,N_12236);
and U12402 (N_12402,N_12232,N_12319);
xnor U12403 (N_12403,N_12302,N_12233);
nor U12404 (N_12404,N_12258,N_12346);
xnor U12405 (N_12405,N_12215,N_12390);
or U12406 (N_12406,N_12248,N_12340);
nand U12407 (N_12407,N_12342,N_12268);
nand U12408 (N_12408,N_12266,N_12255);
xor U12409 (N_12409,N_12359,N_12353);
and U12410 (N_12410,N_12247,N_12269);
nor U12411 (N_12411,N_12219,N_12238);
nor U12412 (N_12412,N_12358,N_12355);
or U12413 (N_12413,N_12237,N_12365);
nand U12414 (N_12414,N_12254,N_12283);
or U12415 (N_12415,N_12304,N_12343);
nand U12416 (N_12416,N_12231,N_12347);
xnor U12417 (N_12417,N_12203,N_12307);
and U12418 (N_12418,N_12244,N_12210);
xor U12419 (N_12419,N_12202,N_12354);
xnor U12420 (N_12420,N_12261,N_12386);
and U12421 (N_12421,N_12399,N_12218);
or U12422 (N_12422,N_12364,N_12290);
nor U12423 (N_12423,N_12381,N_12387);
nand U12424 (N_12424,N_12378,N_12265);
and U12425 (N_12425,N_12291,N_12344);
nor U12426 (N_12426,N_12338,N_12326);
nor U12427 (N_12427,N_12242,N_12382);
or U12428 (N_12428,N_12309,N_12250);
nor U12429 (N_12429,N_12259,N_12288);
nand U12430 (N_12430,N_12267,N_12249);
xor U12431 (N_12431,N_12278,N_12229);
nand U12432 (N_12432,N_12368,N_12377);
xor U12433 (N_12433,N_12213,N_12351);
or U12434 (N_12434,N_12257,N_12306);
or U12435 (N_12435,N_12356,N_12339);
nor U12436 (N_12436,N_12212,N_12375);
nand U12437 (N_12437,N_12240,N_12311);
or U12438 (N_12438,N_12363,N_12332);
nand U12439 (N_12439,N_12333,N_12209);
nor U12440 (N_12440,N_12388,N_12262);
or U12441 (N_12441,N_12222,N_12221);
nand U12442 (N_12442,N_12362,N_12398);
xor U12443 (N_12443,N_12371,N_12337);
nand U12444 (N_12444,N_12389,N_12227);
or U12445 (N_12445,N_12372,N_12397);
or U12446 (N_12446,N_12366,N_12297);
and U12447 (N_12447,N_12360,N_12211);
xnor U12448 (N_12448,N_12384,N_12361);
nor U12449 (N_12449,N_12315,N_12301);
nand U12450 (N_12450,N_12289,N_12251);
nor U12451 (N_12451,N_12349,N_12282);
xnor U12452 (N_12452,N_12243,N_12330);
xnor U12453 (N_12453,N_12220,N_12200);
nor U12454 (N_12454,N_12226,N_12313);
and U12455 (N_12455,N_12252,N_12274);
nor U12456 (N_12456,N_12341,N_12273);
nand U12457 (N_12457,N_12246,N_12345);
or U12458 (N_12458,N_12321,N_12383);
and U12459 (N_12459,N_12271,N_12348);
nand U12460 (N_12460,N_12208,N_12239);
nor U12461 (N_12461,N_12277,N_12336);
or U12462 (N_12462,N_12393,N_12207);
nor U12463 (N_12463,N_12334,N_12296);
nand U12464 (N_12464,N_12316,N_12325);
nand U12465 (N_12465,N_12217,N_12352);
nand U12466 (N_12466,N_12394,N_12357);
xnor U12467 (N_12467,N_12395,N_12206);
and U12468 (N_12468,N_12308,N_12317);
nor U12469 (N_12469,N_12216,N_12392);
nand U12470 (N_12470,N_12225,N_12369);
nor U12471 (N_12471,N_12380,N_12241);
or U12472 (N_12472,N_12367,N_12204);
and U12473 (N_12473,N_12328,N_12331);
or U12474 (N_12474,N_12303,N_12305);
nor U12475 (N_12475,N_12294,N_12295);
and U12476 (N_12476,N_12300,N_12385);
and U12477 (N_12477,N_12391,N_12284);
or U12478 (N_12478,N_12276,N_12299);
or U12479 (N_12479,N_12279,N_12350);
xor U12480 (N_12480,N_12298,N_12245);
nor U12481 (N_12481,N_12376,N_12374);
xor U12482 (N_12482,N_12264,N_12312);
or U12483 (N_12483,N_12230,N_12263);
nor U12484 (N_12484,N_12310,N_12275);
nand U12485 (N_12485,N_12324,N_12318);
and U12486 (N_12486,N_12234,N_12280);
nor U12487 (N_12487,N_12224,N_12292);
nand U12488 (N_12488,N_12396,N_12323);
or U12489 (N_12489,N_12272,N_12270);
nand U12490 (N_12490,N_12329,N_12320);
nand U12491 (N_12491,N_12256,N_12205);
and U12492 (N_12492,N_12228,N_12293);
xor U12493 (N_12493,N_12214,N_12286);
and U12494 (N_12494,N_12335,N_12379);
or U12495 (N_12495,N_12235,N_12281);
or U12496 (N_12496,N_12201,N_12322);
and U12497 (N_12497,N_12260,N_12223);
or U12498 (N_12498,N_12285,N_12370);
or U12499 (N_12499,N_12314,N_12373);
xor U12500 (N_12500,N_12268,N_12374);
or U12501 (N_12501,N_12374,N_12275);
or U12502 (N_12502,N_12397,N_12248);
nor U12503 (N_12503,N_12348,N_12291);
nand U12504 (N_12504,N_12241,N_12341);
and U12505 (N_12505,N_12302,N_12332);
xor U12506 (N_12506,N_12337,N_12259);
and U12507 (N_12507,N_12295,N_12327);
or U12508 (N_12508,N_12252,N_12347);
and U12509 (N_12509,N_12326,N_12291);
xnor U12510 (N_12510,N_12232,N_12243);
xnor U12511 (N_12511,N_12316,N_12395);
nor U12512 (N_12512,N_12329,N_12351);
xor U12513 (N_12513,N_12336,N_12363);
and U12514 (N_12514,N_12201,N_12293);
xor U12515 (N_12515,N_12255,N_12367);
nand U12516 (N_12516,N_12353,N_12334);
nand U12517 (N_12517,N_12211,N_12381);
nor U12518 (N_12518,N_12294,N_12375);
and U12519 (N_12519,N_12391,N_12210);
xor U12520 (N_12520,N_12281,N_12364);
or U12521 (N_12521,N_12258,N_12328);
and U12522 (N_12522,N_12343,N_12262);
nand U12523 (N_12523,N_12306,N_12272);
nor U12524 (N_12524,N_12233,N_12294);
and U12525 (N_12525,N_12208,N_12219);
xnor U12526 (N_12526,N_12337,N_12291);
xnor U12527 (N_12527,N_12206,N_12393);
nand U12528 (N_12528,N_12229,N_12351);
or U12529 (N_12529,N_12301,N_12283);
and U12530 (N_12530,N_12366,N_12375);
nor U12531 (N_12531,N_12253,N_12224);
or U12532 (N_12532,N_12280,N_12244);
nor U12533 (N_12533,N_12381,N_12236);
nor U12534 (N_12534,N_12305,N_12273);
or U12535 (N_12535,N_12372,N_12292);
nor U12536 (N_12536,N_12371,N_12231);
nand U12537 (N_12537,N_12333,N_12383);
nor U12538 (N_12538,N_12313,N_12383);
nand U12539 (N_12539,N_12342,N_12217);
nand U12540 (N_12540,N_12323,N_12381);
nor U12541 (N_12541,N_12375,N_12395);
or U12542 (N_12542,N_12242,N_12324);
or U12543 (N_12543,N_12232,N_12397);
and U12544 (N_12544,N_12277,N_12282);
and U12545 (N_12545,N_12350,N_12392);
nor U12546 (N_12546,N_12229,N_12399);
nor U12547 (N_12547,N_12383,N_12343);
xnor U12548 (N_12548,N_12359,N_12344);
or U12549 (N_12549,N_12266,N_12214);
nor U12550 (N_12550,N_12258,N_12232);
xnor U12551 (N_12551,N_12294,N_12378);
nor U12552 (N_12552,N_12398,N_12365);
xnor U12553 (N_12553,N_12374,N_12380);
nand U12554 (N_12554,N_12226,N_12340);
xnor U12555 (N_12555,N_12367,N_12374);
xnor U12556 (N_12556,N_12356,N_12210);
xor U12557 (N_12557,N_12308,N_12358);
xor U12558 (N_12558,N_12344,N_12380);
nand U12559 (N_12559,N_12331,N_12394);
and U12560 (N_12560,N_12373,N_12397);
or U12561 (N_12561,N_12306,N_12376);
and U12562 (N_12562,N_12269,N_12273);
nor U12563 (N_12563,N_12371,N_12286);
nand U12564 (N_12564,N_12389,N_12360);
nor U12565 (N_12565,N_12265,N_12337);
nor U12566 (N_12566,N_12217,N_12363);
or U12567 (N_12567,N_12399,N_12339);
or U12568 (N_12568,N_12305,N_12274);
nand U12569 (N_12569,N_12397,N_12390);
and U12570 (N_12570,N_12237,N_12363);
nor U12571 (N_12571,N_12343,N_12233);
nand U12572 (N_12572,N_12375,N_12390);
or U12573 (N_12573,N_12292,N_12332);
or U12574 (N_12574,N_12221,N_12310);
or U12575 (N_12575,N_12396,N_12215);
or U12576 (N_12576,N_12255,N_12204);
and U12577 (N_12577,N_12391,N_12396);
and U12578 (N_12578,N_12275,N_12279);
and U12579 (N_12579,N_12377,N_12239);
nand U12580 (N_12580,N_12307,N_12320);
and U12581 (N_12581,N_12261,N_12256);
xnor U12582 (N_12582,N_12284,N_12282);
xor U12583 (N_12583,N_12386,N_12384);
or U12584 (N_12584,N_12362,N_12298);
and U12585 (N_12585,N_12218,N_12268);
nor U12586 (N_12586,N_12285,N_12255);
nor U12587 (N_12587,N_12264,N_12317);
and U12588 (N_12588,N_12382,N_12273);
or U12589 (N_12589,N_12383,N_12277);
and U12590 (N_12590,N_12242,N_12279);
nor U12591 (N_12591,N_12347,N_12212);
nand U12592 (N_12592,N_12245,N_12374);
nand U12593 (N_12593,N_12320,N_12222);
xnor U12594 (N_12594,N_12386,N_12238);
and U12595 (N_12595,N_12224,N_12269);
nor U12596 (N_12596,N_12231,N_12283);
or U12597 (N_12597,N_12205,N_12362);
xor U12598 (N_12598,N_12238,N_12286);
or U12599 (N_12599,N_12317,N_12382);
and U12600 (N_12600,N_12433,N_12472);
xnor U12601 (N_12601,N_12483,N_12575);
nor U12602 (N_12602,N_12453,N_12541);
or U12603 (N_12603,N_12495,N_12535);
and U12604 (N_12604,N_12486,N_12493);
or U12605 (N_12605,N_12475,N_12415);
xnor U12606 (N_12606,N_12410,N_12594);
xor U12607 (N_12607,N_12544,N_12446);
and U12608 (N_12608,N_12401,N_12517);
nor U12609 (N_12609,N_12492,N_12542);
and U12610 (N_12610,N_12507,N_12585);
xnor U12611 (N_12611,N_12509,N_12598);
and U12612 (N_12612,N_12487,N_12559);
nand U12613 (N_12613,N_12568,N_12500);
or U12614 (N_12614,N_12471,N_12422);
nor U12615 (N_12615,N_12451,N_12463);
and U12616 (N_12616,N_12587,N_12409);
xnor U12617 (N_12617,N_12571,N_12527);
and U12618 (N_12618,N_12537,N_12403);
nand U12619 (N_12619,N_12424,N_12512);
xnor U12620 (N_12620,N_12489,N_12404);
nor U12621 (N_12621,N_12498,N_12482);
nor U12622 (N_12622,N_12469,N_12581);
xnor U12623 (N_12623,N_12513,N_12519);
or U12624 (N_12624,N_12461,N_12560);
or U12625 (N_12625,N_12494,N_12408);
and U12626 (N_12626,N_12421,N_12556);
and U12627 (N_12627,N_12413,N_12439);
and U12628 (N_12628,N_12515,N_12456);
nor U12629 (N_12629,N_12427,N_12430);
nand U12630 (N_12630,N_12460,N_12431);
or U12631 (N_12631,N_12450,N_12502);
nor U12632 (N_12632,N_12457,N_12429);
or U12633 (N_12633,N_12562,N_12582);
nor U12634 (N_12634,N_12593,N_12438);
and U12635 (N_12635,N_12503,N_12538);
and U12636 (N_12636,N_12442,N_12553);
nand U12637 (N_12637,N_12576,N_12584);
nor U12638 (N_12638,N_12434,N_12435);
nand U12639 (N_12639,N_12530,N_12583);
xor U12640 (N_12640,N_12449,N_12477);
xnor U12641 (N_12641,N_12595,N_12533);
xnor U12642 (N_12642,N_12443,N_12579);
nor U12643 (N_12643,N_12545,N_12468);
nor U12644 (N_12644,N_12557,N_12566);
xor U12645 (N_12645,N_12470,N_12567);
and U12646 (N_12646,N_12417,N_12580);
nand U12647 (N_12647,N_12528,N_12501);
nand U12648 (N_12648,N_12574,N_12428);
or U12649 (N_12649,N_12529,N_12478);
or U12650 (N_12650,N_12518,N_12534);
and U12651 (N_12651,N_12485,N_12554);
nor U12652 (N_12652,N_12532,N_12570);
and U12653 (N_12653,N_12547,N_12592);
nor U12654 (N_12654,N_12569,N_12526);
nand U12655 (N_12655,N_12578,N_12491);
and U12656 (N_12656,N_12552,N_12536);
or U12657 (N_12657,N_12406,N_12437);
xor U12658 (N_12658,N_12546,N_12504);
nand U12659 (N_12659,N_12467,N_12419);
xor U12660 (N_12660,N_12590,N_12531);
or U12661 (N_12661,N_12555,N_12405);
nor U12662 (N_12662,N_12420,N_12514);
nor U12663 (N_12663,N_12597,N_12550);
nor U12664 (N_12664,N_12473,N_12448);
and U12665 (N_12665,N_12572,N_12496);
and U12666 (N_12666,N_12400,N_12589);
or U12667 (N_12667,N_12563,N_12490);
nand U12668 (N_12668,N_12520,N_12522);
nand U12669 (N_12669,N_12436,N_12479);
nand U12670 (N_12670,N_12425,N_12497);
nand U12671 (N_12671,N_12418,N_12412);
and U12672 (N_12672,N_12599,N_12573);
nor U12673 (N_12673,N_12480,N_12426);
xor U12674 (N_12674,N_12510,N_12516);
and U12675 (N_12675,N_12474,N_12577);
and U12676 (N_12676,N_12445,N_12481);
or U12677 (N_12677,N_12524,N_12505);
nor U12678 (N_12678,N_12499,N_12506);
and U12679 (N_12679,N_12447,N_12596);
xnor U12680 (N_12680,N_12511,N_12551);
xnor U12681 (N_12681,N_12539,N_12525);
nor U12682 (N_12682,N_12564,N_12432);
or U12683 (N_12683,N_12459,N_12591);
xnor U12684 (N_12684,N_12484,N_12462);
or U12685 (N_12685,N_12588,N_12407);
nand U12686 (N_12686,N_12586,N_12423);
nor U12687 (N_12687,N_12416,N_12543);
nand U12688 (N_12688,N_12488,N_12521);
xnor U12689 (N_12689,N_12466,N_12549);
nand U12690 (N_12690,N_12411,N_12454);
xnor U12691 (N_12691,N_12465,N_12414);
nand U12692 (N_12692,N_12440,N_12548);
xor U12693 (N_12693,N_12464,N_12455);
and U12694 (N_12694,N_12458,N_12444);
xor U12695 (N_12695,N_12508,N_12561);
or U12696 (N_12696,N_12441,N_12476);
nand U12697 (N_12697,N_12402,N_12452);
xnor U12698 (N_12698,N_12565,N_12558);
and U12699 (N_12699,N_12523,N_12540);
xor U12700 (N_12700,N_12449,N_12479);
or U12701 (N_12701,N_12404,N_12448);
and U12702 (N_12702,N_12484,N_12416);
or U12703 (N_12703,N_12589,N_12436);
and U12704 (N_12704,N_12485,N_12572);
and U12705 (N_12705,N_12472,N_12528);
nor U12706 (N_12706,N_12580,N_12455);
or U12707 (N_12707,N_12465,N_12482);
nand U12708 (N_12708,N_12589,N_12427);
nor U12709 (N_12709,N_12485,N_12596);
xor U12710 (N_12710,N_12576,N_12572);
xor U12711 (N_12711,N_12442,N_12561);
nor U12712 (N_12712,N_12417,N_12455);
xnor U12713 (N_12713,N_12573,N_12511);
nand U12714 (N_12714,N_12407,N_12565);
or U12715 (N_12715,N_12523,N_12563);
nor U12716 (N_12716,N_12546,N_12577);
nand U12717 (N_12717,N_12463,N_12563);
and U12718 (N_12718,N_12519,N_12428);
nor U12719 (N_12719,N_12481,N_12495);
or U12720 (N_12720,N_12598,N_12474);
nand U12721 (N_12721,N_12592,N_12452);
nand U12722 (N_12722,N_12574,N_12526);
nor U12723 (N_12723,N_12494,N_12466);
and U12724 (N_12724,N_12496,N_12436);
nand U12725 (N_12725,N_12439,N_12482);
or U12726 (N_12726,N_12547,N_12448);
xor U12727 (N_12727,N_12561,N_12458);
xor U12728 (N_12728,N_12525,N_12592);
and U12729 (N_12729,N_12569,N_12586);
nor U12730 (N_12730,N_12578,N_12425);
and U12731 (N_12731,N_12403,N_12412);
nor U12732 (N_12732,N_12489,N_12525);
and U12733 (N_12733,N_12526,N_12512);
or U12734 (N_12734,N_12578,N_12493);
xnor U12735 (N_12735,N_12405,N_12579);
and U12736 (N_12736,N_12419,N_12468);
or U12737 (N_12737,N_12409,N_12488);
nand U12738 (N_12738,N_12599,N_12409);
nand U12739 (N_12739,N_12515,N_12449);
xor U12740 (N_12740,N_12566,N_12479);
xor U12741 (N_12741,N_12457,N_12483);
or U12742 (N_12742,N_12520,N_12566);
or U12743 (N_12743,N_12591,N_12596);
and U12744 (N_12744,N_12515,N_12400);
nor U12745 (N_12745,N_12401,N_12522);
or U12746 (N_12746,N_12539,N_12506);
or U12747 (N_12747,N_12589,N_12534);
and U12748 (N_12748,N_12415,N_12462);
and U12749 (N_12749,N_12584,N_12410);
xor U12750 (N_12750,N_12510,N_12421);
nor U12751 (N_12751,N_12559,N_12459);
xnor U12752 (N_12752,N_12411,N_12453);
nand U12753 (N_12753,N_12468,N_12572);
nor U12754 (N_12754,N_12553,N_12487);
xnor U12755 (N_12755,N_12531,N_12566);
and U12756 (N_12756,N_12598,N_12569);
nor U12757 (N_12757,N_12410,N_12434);
or U12758 (N_12758,N_12532,N_12597);
or U12759 (N_12759,N_12562,N_12492);
and U12760 (N_12760,N_12535,N_12429);
and U12761 (N_12761,N_12516,N_12571);
xor U12762 (N_12762,N_12482,N_12409);
and U12763 (N_12763,N_12533,N_12527);
nand U12764 (N_12764,N_12480,N_12447);
and U12765 (N_12765,N_12558,N_12504);
or U12766 (N_12766,N_12494,N_12510);
nor U12767 (N_12767,N_12598,N_12455);
nor U12768 (N_12768,N_12458,N_12588);
nor U12769 (N_12769,N_12589,N_12531);
nand U12770 (N_12770,N_12481,N_12564);
nor U12771 (N_12771,N_12558,N_12463);
nand U12772 (N_12772,N_12558,N_12401);
nand U12773 (N_12773,N_12460,N_12413);
xnor U12774 (N_12774,N_12488,N_12414);
xor U12775 (N_12775,N_12528,N_12551);
nor U12776 (N_12776,N_12528,N_12511);
and U12777 (N_12777,N_12563,N_12488);
xnor U12778 (N_12778,N_12593,N_12404);
nand U12779 (N_12779,N_12418,N_12528);
and U12780 (N_12780,N_12423,N_12578);
or U12781 (N_12781,N_12575,N_12563);
xor U12782 (N_12782,N_12468,N_12590);
nor U12783 (N_12783,N_12435,N_12460);
and U12784 (N_12784,N_12471,N_12538);
nand U12785 (N_12785,N_12457,N_12465);
and U12786 (N_12786,N_12404,N_12434);
nand U12787 (N_12787,N_12520,N_12486);
xor U12788 (N_12788,N_12595,N_12567);
xnor U12789 (N_12789,N_12462,N_12584);
and U12790 (N_12790,N_12401,N_12470);
or U12791 (N_12791,N_12501,N_12473);
nor U12792 (N_12792,N_12447,N_12460);
xnor U12793 (N_12793,N_12525,N_12406);
nor U12794 (N_12794,N_12407,N_12494);
xor U12795 (N_12795,N_12476,N_12506);
or U12796 (N_12796,N_12497,N_12407);
and U12797 (N_12797,N_12421,N_12502);
nor U12798 (N_12798,N_12404,N_12421);
or U12799 (N_12799,N_12467,N_12589);
nor U12800 (N_12800,N_12781,N_12753);
and U12801 (N_12801,N_12640,N_12755);
or U12802 (N_12802,N_12698,N_12691);
nor U12803 (N_12803,N_12706,N_12602);
and U12804 (N_12804,N_12618,N_12692);
and U12805 (N_12805,N_12757,N_12702);
and U12806 (N_12806,N_12601,N_12688);
xnor U12807 (N_12807,N_12600,N_12758);
or U12808 (N_12808,N_12678,N_12682);
xnor U12809 (N_12809,N_12625,N_12690);
or U12810 (N_12810,N_12783,N_12773);
xor U12811 (N_12811,N_12627,N_12761);
xor U12812 (N_12812,N_12684,N_12654);
and U12813 (N_12813,N_12655,N_12778);
nand U12814 (N_12814,N_12703,N_12637);
nor U12815 (N_12815,N_12718,N_12669);
nand U12816 (N_12816,N_12624,N_12786);
and U12817 (N_12817,N_12708,N_12769);
nand U12818 (N_12818,N_12653,N_12792);
nand U12819 (N_12819,N_12738,N_12610);
and U12820 (N_12820,N_12799,N_12686);
nand U12821 (N_12821,N_12659,N_12707);
nand U12822 (N_12822,N_12651,N_12789);
nand U12823 (N_12823,N_12794,N_12607);
nand U12824 (N_12824,N_12784,N_12603);
or U12825 (N_12825,N_12623,N_12733);
nor U12826 (N_12826,N_12726,N_12736);
or U12827 (N_12827,N_12614,N_12720);
nor U12828 (N_12828,N_12643,N_12683);
or U12829 (N_12829,N_12656,N_12797);
nand U12830 (N_12830,N_12664,N_12670);
nor U12831 (N_12831,N_12700,N_12609);
nand U12832 (N_12832,N_12652,N_12729);
nand U12833 (N_12833,N_12663,N_12742);
and U12834 (N_12834,N_12766,N_12631);
and U12835 (N_12835,N_12730,N_12611);
and U12836 (N_12836,N_12696,N_12775);
nor U12837 (N_12837,N_12677,N_12679);
or U12838 (N_12838,N_12795,N_12605);
and U12839 (N_12839,N_12645,N_12616);
xor U12840 (N_12840,N_12763,N_12648);
and U12841 (N_12841,N_12734,N_12728);
or U12842 (N_12842,N_12737,N_12777);
nand U12843 (N_12843,N_12715,N_12796);
and U12844 (N_12844,N_12768,N_12639);
nor U12845 (N_12845,N_12608,N_12642);
or U12846 (N_12846,N_12619,N_12701);
nand U12847 (N_12847,N_12740,N_12617);
nand U12848 (N_12848,N_12687,N_12672);
or U12849 (N_12849,N_12722,N_12732);
or U12850 (N_12850,N_12725,N_12746);
or U12851 (N_12851,N_12704,N_12661);
nand U12852 (N_12852,N_12699,N_12731);
nor U12853 (N_12853,N_12749,N_12622);
nand U12854 (N_12854,N_12748,N_12615);
or U12855 (N_12855,N_12739,N_12780);
xnor U12856 (N_12856,N_12710,N_12790);
nor U12857 (N_12857,N_12717,N_12693);
nand U12858 (N_12858,N_12675,N_12716);
or U12859 (N_12859,N_12657,N_12628);
xor U12860 (N_12860,N_12666,N_12750);
and U12861 (N_12861,N_12697,N_12764);
and U12862 (N_12862,N_12668,N_12667);
xnor U12863 (N_12863,N_12641,N_12662);
and U12864 (N_12864,N_12646,N_12647);
xnor U12865 (N_12865,N_12685,N_12660);
or U12866 (N_12866,N_12612,N_12771);
or U12867 (N_12867,N_12712,N_12759);
and U12868 (N_12868,N_12689,N_12779);
nor U12869 (N_12869,N_12798,N_12694);
nand U12870 (N_12870,N_12630,N_12752);
or U12871 (N_12871,N_12724,N_12606);
xnor U12872 (N_12872,N_12695,N_12681);
or U12873 (N_12873,N_12629,N_12649);
or U12874 (N_12874,N_12671,N_12711);
nand U12875 (N_12875,N_12638,N_12674);
and U12876 (N_12876,N_12791,N_12634);
and U12877 (N_12877,N_12604,N_12727);
xor U12878 (N_12878,N_12621,N_12787);
xnor U12879 (N_12879,N_12658,N_12770);
nand U12880 (N_12880,N_12762,N_12747);
and U12881 (N_12881,N_12741,N_12644);
and U12882 (N_12882,N_12676,N_12709);
nor U12883 (N_12883,N_12714,N_12765);
nor U12884 (N_12884,N_12756,N_12782);
nand U12885 (N_12885,N_12620,N_12723);
and U12886 (N_12886,N_12680,N_12760);
or U12887 (N_12887,N_12719,N_12705);
or U12888 (N_12888,N_12767,N_12626);
nand U12889 (N_12889,N_12776,N_12744);
xor U12890 (N_12890,N_12721,N_12743);
or U12891 (N_12891,N_12754,N_12751);
and U12892 (N_12892,N_12673,N_12632);
and U12893 (N_12893,N_12785,N_12774);
or U12894 (N_12894,N_12735,N_12772);
nand U12895 (N_12895,N_12650,N_12793);
nand U12896 (N_12896,N_12613,N_12635);
nor U12897 (N_12897,N_12788,N_12745);
nor U12898 (N_12898,N_12713,N_12636);
xnor U12899 (N_12899,N_12633,N_12665);
xor U12900 (N_12900,N_12746,N_12645);
and U12901 (N_12901,N_12791,N_12785);
or U12902 (N_12902,N_12789,N_12765);
xor U12903 (N_12903,N_12672,N_12621);
nor U12904 (N_12904,N_12787,N_12608);
xor U12905 (N_12905,N_12773,N_12623);
nor U12906 (N_12906,N_12642,N_12785);
or U12907 (N_12907,N_12624,N_12633);
and U12908 (N_12908,N_12735,N_12650);
or U12909 (N_12909,N_12730,N_12777);
nor U12910 (N_12910,N_12649,N_12624);
or U12911 (N_12911,N_12695,N_12608);
or U12912 (N_12912,N_12619,N_12721);
or U12913 (N_12913,N_12732,N_12726);
nor U12914 (N_12914,N_12704,N_12792);
or U12915 (N_12915,N_12718,N_12639);
and U12916 (N_12916,N_12704,N_12731);
xnor U12917 (N_12917,N_12664,N_12653);
or U12918 (N_12918,N_12702,N_12749);
and U12919 (N_12919,N_12714,N_12792);
and U12920 (N_12920,N_12752,N_12779);
nand U12921 (N_12921,N_12617,N_12732);
or U12922 (N_12922,N_12698,N_12773);
or U12923 (N_12923,N_12683,N_12662);
nand U12924 (N_12924,N_12792,N_12633);
nand U12925 (N_12925,N_12782,N_12679);
xnor U12926 (N_12926,N_12729,N_12603);
and U12927 (N_12927,N_12782,N_12649);
nor U12928 (N_12928,N_12634,N_12643);
xnor U12929 (N_12929,N_12685,N_12692);
or U12930 (N_12930,N_12775,N_12753);
nand U12931 (N_12931,N_12678,N_12747);
xnor U12932 (N_12932,N_12683,N_12640);
and U12933 (N_12933,N_12747,N_12751);
xnor U12934 (N_12934,N_12680,N_12708);
and U12935 (N_12935,N_12694,N_12777);
or U12936 (N_12936,N_12670,N_12795);
or U12937 (N_12937,N_12658,N_12700);
and U12938 (N_12938,N_12728,N_12769);
or U12939 (N_12939,N_12623,N_12724);
nor U12940 (N_12940,N_12626,N_12709);
nand U12941 (N_12941,N_12746,N_12630);
nand U12942 (N_12942,N_12641,N_12769);
nand U12943 (N_12943,N_12670,N_12657);
and U12944 (N_12944,N_12691,N_12677);
xor U12945 (N_12945,N_12796,N_12627);
nor U12946 (N_12946,N_12605,N_12732);
nand U12947 (N_12947,N_12671,N_12739);
or U12948 (N_12948,N_12780,N_12673);
or U12949 (N_12949,N_12648,N_12668);
xor U12950 (N_12950,N_12665,N_12760);
xor U12951 (N_12951,N_12765,N_12777);
and U12952 (N_12952,N_12781,N_12663);
nand U12953 (N_12953,N_12751,N_12668);
and U12954 (N_12954,N_12647,N_12657);
xor U12955 (N_12955,N_12663,N_12624);
and U12956 (N_12956,N_12743,N_12648);
nand U12957 (N_12957,N_12757,N_12753);
or U12958 (N_12958,N_12762,N_12779);
xor U12959 (N_12959,N_12749,N_12632);
nand U12960 (N_12960,N_12767,N_12617);
nor U12961 (N_12961,N_12663,N_12669);
nor U12962 (N_12962,N_12609,N_12677);
nand U12963 (N_12963,N_12779,N_12661);
or U12964 (N_12964,N_12690,N_12631);
nand U12965 (N_12965,N_12677,N_12681);
nor U12966 (N_12966,N_12676,N_12683);
xnor U12967 (N_12967,N_12646,N_12780);
nor U12968 (N_12968,N_12731,N_12632);
nand U12969 (N_12969,N_12692,N_12769);
nor U12970 (N_12970,N_12621,N_12767);
and U12971 (N_12971,N_12780,N_12644);
xnor U12972 (N_12972,N_12648,N_12782);
nand U12973 (N_12973,N_12624,N_12660);
xor U12974 (N_12974,N_12673,N_12634);
nor U12975 (N_12975,N_12637,N_12719);
nand U12976 (N_12976,N_12756,N_12727);
and U12977 (N_12977,N_12773,N_12789);
xnor U12978 (N_12978,N_12686,N_12638);
xnor U12979 (N_12979,N_12792,N_12782);
nor U12980 (N_12980,N_12623,N_12622);
or U12981 (N_12981,N_12762,N_12773);
or U12982 (N_12982,N_12600,N_12721);
nand U12983 (N_12983,N_12685,N_12625);
or U12984 (N_12984,N_12792,N_12793);
and U12985 (N_12985,N_12726,N_12609);
nand U12986 (N_12986,N_12710,N_12659);
nor U12987 (N_12987,N_12705,N_12780);
nor U12988 (N_12988,N_12702,N_12786);
nand U12989 (N_12989,N_12729,N_12629);
xor U12990 (N_12990,N_12705,N_12749);
nor U12991 (N_12991,N_12797,N_12655);
and U12992 (N_12992,N_12619,N_12639);
nor U12993 (N_12993,N_12650,N_12750);
nand U12994 (N_12994,N_12628,N_12782);
and U12995 (N_12995,N_12710,N_12772);
and U12996 (N_12996,N_12639,N_12791);
nand U12997 (N_12997,N_12771,N_12699);
nand U12998 (N_12998,N_12617,N_12709);
nand U12999 (N_12999,N_12610,N_12789);
xnor U13000 (N_13000,N_12881,N_12825);
nor U13001 (N_13001,N_12806,N_12901);
xor U13002 (N_13002,N_12814,N_12935);
xnor U13003 (N_13003,N_12990,N_12829);
and U13004 (N_13004,N_12998,N_12858);
or U13005 (N_13005,N_12955,N_12986);
xor U13006 (N_13006,N_12804,N_12960);
xor U13007 (N_13007,N_12981,N_12803);
nor U13008 (N_13008,N_12802,N_12912);
and U13009 (N_13009,N_12915,N_12866);
nor U13010 (N_13010,N_12900,N_12840);
nor U13011 (N_13011,N_12819,N_12953);
nand U13012 (N_13012,N_12879,N_12907);
and U13013 (N_13013,N_12834,N_12911);
and U13014 (N_13014,N_12952,N_12966);
and U13015 (N_13015,N_12841,N_12941);
nor U13016 (N_13016,N_12848,N_12877);
and U13017 (N_13017,N_12930,N_12861);
and U13018 (N_13018,N_12882,N_12983);
nor U13019 (N_13019,N_12893,N_12887);
xnor U13020 (N_13020,N_12818,N_12862);
nor U13021 (N_13021,N_12926,N_12922);
xnor U13022 (N_13022,N_12820,N_12962);
and U13023 (N_13023,N_12849,N_12967);
or U13024 (N_13024,N_12874,N_12944);
nand U13025 (N_13025,N_12826,N_12931);
or U13026 (N_13026,N_12857,N_12869);
and U13027 (N_13027,N_12934,N_12868);
nand U13028 (N_13028,N_12894,N_12828);
xor U13029 (N_13029,N_12816,N_12871);
nor U13030 (N_13030,N_12957,N_12830);
xor U13031 (N_13031,N_12860,N_12845);
or U13032 (N_13032,N_12973,N_12899);
xnor U13033 (N_13033,N_12995,N_12815);
xnor U13034 (N_13034,N_12932,N_12927);
and U13035 (N_13035,N_12898,N_12936);
and U13036 (N_13036,N_12925,N_12961);
or U13037 (N_13037,N_12831,N_12942);
nor U13038 (N_13038,N_12821,N_12836);
xor U13039 (N_13039,N_12916,N_12940);
nand U13040 (N_13040,N_12801,N_12959);
nand U13041 (N_13041,N_12867,N_12933);
nor U13042 (N_13042,N_12993,N_12949);
or U13043 (N_13043,N_12856,N_12888);
xor U13044 (N_13044,N_12977,N_12805);
nand U13045 (N_13045,N_12904,N_12895);
xor U13046 (N_13046,N_12937,N_12905);
nor U13047 (N_13047,N_12914,N_12880);
nand U13048 (N_13048,N_12883,N_12903);
nand U13049 (N_13049,N_12808,N_12992);
nand U13050 (N_13050,N_12996,N_12850);
nor U13051 (N_13051,N_12999,N_12978);
or U13052 (N_13052,N_12946,N_12884);
xnor U13053 (N_13053,N_12913,N_12918);
or U13054 (N_13054,N_12950,N_12800);
nand U13055 (N_13055,N_12994,N_12833);
nor U13056 (N_13056,N_12902,N_12908);
nand U13057 (N_13057,N_12964,N_12954);
xor U13058 (N_13058,N_12919,N_12975);
xnor U13059 (N_13059,N_12811,N_12958);
xor U13060 (N_13060,N_12985,N_12832);
nor U13061 (N_13061,N_12863,N_12854);
or U13062 (N_13062,N_12963,N_12917);
and U13063 (N_13063,N_12890,N_12965);
xnor U13064 (N_13064,N_12980,N_12943);
nand U13065 (N_13065,N_12870,N_12948);
or U13066 (N_13066,N_12974,N_12824);
and U13067 (N_13067,N_12989,N_12873);
nor U13068 (N_13068,N_12921,N_12971);
nand U13069 (N_13069,N_12807,N_12976);
and U13070 (N_13070,N_12891,N_12865);
nand U13071 (N_13071,N_12817,N_12979);
xnor U13072 (N_13072,N_12875,N_12988);
xnor U13073 (N_13073,N_12972,N_12982);
xnor U13074 (N_13074,N_12835,N_12909);
and U13075 (N_13075,N_12906,N_12843);
nor U13076 (N_13076,N_12844,N_12984);
nand U13077 (N_13077,N_12939,N_12889);
or U13078 (N_13078,N_12896,N_12837);
and U13079 (N_13079,N_12823,N_12842);
or U13080 (N_13080,N_12855,N_12872);
xnor U13081 (N_13081,N_12924,N_12827);
xnor U13082 (N_13082,N_12991,N_12853);
nor U13083 (N_13083,N_12897,N_12812);
nand U13084 (N_13084,N_12928,N_12847);
or U13085 (N_13085,N_12838,N_12910);
nor U13086 (N_13086,N_12809,N_12969);
nand U13087 (N_13087,N_12846,N_12864);
xnor U13088 (N_13088,N_12892,N_12878);
xor U13089 (N_13089,N_12920,N_12859);
xor U13090 (N_13090,N_12839,N_12987);
and U13091 (N_13091,N_12970,N_12852);
or U13092 (N_13092,N_12956,N_12876);
and U13093 (N_13093,N_12947,N_12938);
xor U13094 (N_13094,N_12886,N_12885);
xnor U13095 (N_13095,N_12951,N_12813);
nand U13096 (N_13096,N_12997,N_12822);
xnor U13097 (N_13097,N_12923,N_12945);
nand U13098 (N_13098,N_12851,N_12810);
nor U13099 (N_13099,N_12968,N_12929);
and U13100 (N_13100,N_12916,N_12928);
nor U13101 (N_13101,N_12808,N_12908);
nand U13102 (N_13102,N_12871,N_12931);
nand U13103 (N_13103,N_12814,N_12930);
xor U13104 (N_13104,N_12853,N_12872);
and U13105 (N_13105,N_12932,N_12847);
nand U13106 (N_13106,N_12808,N_12862);
or U13107 (N_13107,N_12933,N_12861);
xnor U13108 (N_13108,N_12810,N_12910);
and U13109 (N_13109,N_12951,N_12954);
and U13110 (N_13110,N_12813,N_12839);
and U13111 (N_13111,N_12820,N_12801);
nor U13112 (N_13112,N_12945,N_12835);
or U13113 (N_13113,N_12809,N_12974);
or U13114 (N_13114,N_12960,N_12832);
nand U13115 (N_13115,N_12939,N_12917);
and U13116 (N_13116,N_12941,N_12950);
xnor U13117 (N_13117,N_12974,N_12910);
xnor U13118 (N_13118,N_12917,N_12893);
and U13119 (N_13119,N_12847,N_12897);
and U13120 (N_13120,N_12931,N_12951);
and U13121 (N_13121,N_12814,N_12827);
nand U13122 (N_13122,N_12923,N_12800);
xnor U13123 (N_13123,N_12867,N_12850);
xor U13124 (N_13124,N_12931,N_12834);
or U13125 (N_13125,N_12929,N_12941);
or U13126 (N_13126,N_12946,N_12968);
nand U13127 (N_13127,N_12850,N_12874);
xnor U13128 (N_13128,N_12996,N_12872);
nor U13129 (N_13129,N_12816,N_12824);
nor U13130 (N_13130,N_12955,N_12942);
or U13131 (N_13131,N_12892,N_12964);
xor U13132 (N_13132,N_12828,N_12811);
nor U13133 (N_13133,N_12970,N_12915);
nor U13134 (N_13134,N_12848,N_12972);
and U13135 (N_13135,N_12837,N_12997);
nand U13136 (N_13136,N_12839,N_12921);
nand U13137 (N_13137,N_12999,N_12948);
xnor U13138 (N_13138,N_12858,N_12977);
and U13139 (N_13139,N_12957,N_12893);
and U13140 (N_13140,N_12896,N_12814);
and U13141 (N_13141,N_12835,N_12947);
and U13142 (N_13142,N_12928,N_12819);
and U13143 (N_13143,N_12906,N_12929);
nand U13144 (N_13144,N_12972,N_12835);
or U13145 (N_13145,N_12829,N_12822);
and U13146 (N_13146,N_12882,N_12912);
nor U13147 (N_13147,N_12813,N_12972);
or U13148 (N_13148,N_12992,N_12880);
xnor U13149 (N_13149,N_12803,N_12999);
nor U13150 (N_13150,N_12825,N_12908);
nand U13151 (N_13151,N_12977,N_12916);
nor U13152 (N_13152,N_12940,N_12842);
xor U13153 (N_13153,N_12967,N_12842);
nand U13154 (N_13154,N_12992,N_12984);
nor U13155 (N_13155,N_12856,N_12811);
or U13156 (N_13156,N_12922,N_12821);
and U13157 (N_13157,N_12893,N_12881);
xnor U13158 (N_13158,N_12882,N_12929);
xor U13159 (N_13159,N_12979,N_12846);
or U13160 (N_13160,N_12808,N_12833);
and U13161 (N_13161,N_12955,N_12982);
or U13162 (N_13162,N_12834,N_12889);
xor U13163 (N_13163,N_12930,N_12902);
nor U13164 (N_13164,N_12899,N_12802);
nor U13165 (N_13165,N_12900,N_12989);
or U13166 (N_13166,N_12818,N_12852);
nor U13167 (N_13167,N_12964,N_12878);
xnor U13168 (N_13168,N_12927,N_12909);
or U13169 (N_13169,N_12822,N_12925);
and U13170 (N_13170,N_12972,N_12829);
or U13171 (N_13171,N_12954,N_12918);
xor U13172 (N_13172,N_12938,N_12904);
xnor U13173 (N_13173,N_12865,N_12898);
nand U13174 (N_13174,N_12857,N_12814);
nand U13175 (N_13175,N_12973,N_12812);
or U13176 (N_13176,N_12888,N_12900);
xor U13177 (N_13177,N_12826,N_12998);
nand U13178 (N_13178,N_12984,N_12807);
nor U13179 (N_13179,N_12863,N_12878);
and U13180 (N_13180,N_12992,N_12827);
nand U13181 (N_13181,N_12937,N_12993);
and U13182 (N_13182,N_12975,N_12973);
xor U13183 (N_13183,N_12834,N_12846);
xnor U13184 (N_13184,N_12824,N_12994);
and U13185 (N_13185,N_12817,N_12812);
and U13186 (N_13186,N_12948,N_12862);
nor U13187 (N_13187,N_12919,N_12930);
or U13188 (N_13188,N_12995,N_12996);
nor U13189 (N_13189,N_12847,N_12971);
nor U13190 (N_13190,N_12929,N_12936);
or U13191 (N_13191,N_12865,N_12838);
nand U13192 (N_13192,N_12918,N_12803);
xnor U13193 (N_13193,N_12960,N_12944);
nand U13194 (N_13194,N_12823,N_12930);
nand U13195 (N_13195,N_12849,N_12924);
nor U13196 (N_13196,N_12920,N_12844);
and U13197 (N_13197,N_12931,N_12906);
or U13198 (N_13198,N_12875,N_12873);
nand U13199 (N_13199,N_12938,N_12908);
and U13200 (N_13200,N_13032,N_13131);
nor U13201 (N_13201,N_13098,N_13156);
xnor U13202 (N_13202,N_13025,N_13014);
or U13203 (N_13203,N_13018,N_13091);
nor U13204 (N_13204,N_13102,N_13082);
or U13205 (N_13205,N_13045,N_13072);
xor U13206 (N_13206,N_13002,N_13012);
and U13207 (N_13207,N_13041,N_13024);
and U13208 (N_13208,N_13171,N_13095);
nor U13209 (N_13209,N_13114,N_13175);
nor U13210 (N_13210,N_13015,N_13123);
nand U13211 (N_13211,N_13051,N_13009);
or U13212 (N_13212,N_13159,N_13142);
nand U13213 (N_13213,N_13000,N_13145);
or U13214 (N_13214,N_13126,N_13003);
xor U13215 (N_13215,N_13099,N_13147);
and U13216 (N_13216,N_13083,N_13075);
or U13217 (N_13217,N_13093,N_13193);
and U13218 (N_13218,N_13143,N_13121);
nand U13219 (N_13219,N_13031,N_13042);
and U13220 (N_13220,N_13013,N_13162);
nand U13221 (N_13221,N_13058,N_13027);
or U13222 (N_13222,N_13150,N_13155);
and U13223 (N_13223,N_13053,N_13017);
nor U13224 (N_13224,N_13029,N_13070);
nor U13225 (N_13225,N_13004,N_13116);
nor U13226 (N_13226,N_13074,N_13113);
and U13227 (N_13227,N_13065,N_13157);
nor U13228 (N_13228,N_13179,N_13184);
nand U13229 (N_13229,N_13194,N_13103);
or U13230 (N_13230,N_13039,N_13063);
nor U13231 (N_13231,N_13117,N_13006);
nor U13232 (N_13232,N_13188,N_13108);
and U13233 (N_13233,N_13059,N_13010);
and U13234 (N_13234,N_13137,N_13097);
and U13235 (N_13235,N_13043,N_13005);
or U13236 (N_13236,N_13183,N_13192);
nor U13237 (N_13237,N_13189,N_13119);
or U13238 (N_13238,N_13177,N_13066);
and U13239 (N_13239,N_13067,N_13166);
nand U13240 (N_13240,N_13105,N_13073);
and U13241 (N_13241,N_13081,N_13084);
and U13242 (N_13242,N_13094,N_13057);
xor U13243 (N_13243,N_13125,N_13139);
or U13244 (N_13244,N_13047,N_13158);
nor U13245 (N_13245,N_13050,N_13185);
xnor U13246 (N_13246,N_13169,N_13138);
nand U13247 (N_13247,N_13187,N_13181);
nor U13248 (N_13248,N_13174,N_13148);
and U13249 (N_13249,N_13182,N_13052);
or U13250 (N_13250,N_13037,N_13046);
xnor U13251 (N_13251,N_13186,N_13011);
xnor U13252 (N_13252,N_13089,N_13136);
or U13253 (N_13253,N_13100,N_13023);
xnor U13254 (N_13254,N_13118,N_13160);
nor U13255 (N_13255,N_13104,N_13176);
xnor U13256 (N_13256,N_13168,N_13151);
xor U13257 (N_13257,N_13085,N_13054);
nor U13258 (N_13258,N_13195,N_13008);
nor U13259 (N_13259,N_13115,N_13064);
nand U13260 (N_13260,N_13061,N_13180);
nand U13261 (N_13261,N_13164,N_13172);
nand U13262 (N_13262,N_13049,N_13132);
nor U13263 (N_13263,N_13129,N_13001);
xor U13264 (N_13264,N_13106,N_13130);
and U13265 (N_13265,N_13196,N_13178);
nand U13266 (N_13266,N_13096,N_13197);
nor U13267 (N_13267,N_13034,N_13110);
xor U13268 (N_13268,N_13133,N_13144);
xor U13269 (N_13269,N_13109,N_13190);
nor U13270 (N_13270,N_13153,N_13198);
and U13271 (N_13271,N_13048,N_13086);
nand U13272 (N_13272,N_13079,N_13088);
nand U13273 (N_13273,N_13026,N_13120);
xnor U13274 (N_13274,N_13135,N_13068);
nor U13275 (N_13275,N_13127,N_13161);
and U13276 (N_13276,N_13101,N_13019);
xor U13277 (N_13277,N_13199,N_13141);
xor U13278 (N_13278,N_13122,N_13112);
xor U13279 (N_13279,N_13124,N_13022);
nor U13280 (N_13280,N_13044,N_13055);
nor U13281 (N_13281,N_13191,N_13111);
and U13282 (N_13282,N_13040,N_13035);
nand U13283 (N_13283,N_13071,N_13146);
and U13284 (N_13284,N_13007,N_13078);
xnor U13285 (N_13285,N_13092,N_13163);
xor U13286 (N_13286,N_13021,N_13090);
and U13287 (N_13287,N_13016,N_13165);
nand U13288 (N_13288,N_13173,N_13062);
xnor U13289 (N_13289,N_13036,N_13060);
and U13290 (N_13290,N_13076,N_13056);
nor U13291 (N_13291,N_13149,N_13069);
nor U13292 (N_13292,N_13033,N_13140);
and U13293 (N_13293,N_13080,N_13038);
nand U13294 (N_13294,N_13087,N_13167);
and U13295 (N_13295,N_13128,N_13077);
and U13296 (N_13296,N_13030,N_13107);
and U13297 (N_13297,N_13020,N_13028);
xor U13298 (N_13298,N_13152,N_13170);
and U13299 (N_13299,N_13134,N_13154);
xor U13300 (N_13300,N_13174,N_13166);
and U13301 (N_13301,N_13180,N_13155);
nor U13302 (N_13302,N_13170,N_13171);
or U13303 (N_13303,N_13025,N_13104);
nand U13304 (N_13304,N_13183,N_13086);
nor U13305 (N_13305,N_13167,N_13062);
nor U13306 (N_13306,N_13110,N_13044);
and U13307 (N_13307,N_13090,N_13052);
nand U13308 (N_13308,N_13068,N_13048);
and U13309 (N_13309,N_13107,N_13174);
xnor U13310 (N_13310,N_13171,N_13111);
and U13311 (N_13311,N_13000,N_13156);
nand U13312 (N_13312,N_13100,N_13132);
and U13313 (N_13313,N_13026,N_13162);
or U13314 (N_13314,N_13186,N_13142);
xnor U13315 (N_13315,N_13059,N_13114);
or U13316 (N_13316,N_13049,N_13010);
and U13317 (N_13317,N_13026,N_13128);
and U13318 (N_13318,N_13073,N_13035);
nor U13319 (N_13319,N_13062,N_13003);
xnor U13320 (N_13320,N_13143,N_13117);
or U13321 (N_13321,N_13099,N_13098);
and U13322 (N_13322,N_13031,N_13094);
and U13323 (N_13323,N_13199,N_13147);
and U13324 (N_13324,N_13091,N_13180);
or U13325 (N_13325,N_13067,N_13042);
and U13326 (N_13326,N_13061,N_13093);
nand U13327 (N_13327,N_13071,N_13067);
and U13328 (N_13328,N_13059,N_13005);
nor U13329 (N_13329,N_13152,N_13182);
nand U13330 (N_13330,N_13175,N_13098);
xor U13331 (N_13331,N_13182,N_13082);
nand U13332 (N_13332,N_13105,N_13021);
and U13333 (N_13333,N_13150,N_13089);
nand U13334 (N_13334,N_13100,N_13120);
nor U13335 (N_13335,N_13130,N_13085);
nand U13336 (N_13336,N_13053,N_13057);
or U13337 (N_13337,N_13186,N_13059);
nor U13338 (N_13338,N_13008,N_13163);
or U13339 (N_13339,N_13069,N_13141);
nor U13340 (N_13340,N_13139,N_13062);
xnor U13341 (N_13341,N_13175,N_13095);
nand U13342 (N_13342,N_13102,N_13084);
or U13343 (N_13343,N_13001,N_13152);
and U13344 (N_13344,N_13057,N_13093);
and U13345 (N_13345,N_13199,N_13183);
nor U13346 (N_13346,N_13038,N_13128);
nor U13347 (N_13347,N_13076,N_13064);
xor U13348 (N_13348,N_13114,N_13149);
and U13349 (N_13349,N_13123,N_13086);
nor U13350 (N_13350,N_13096,N_13098);
nor U13351 (N_13351,N_13072,N_13196);
or U13352 (N_13352,N_13041,N_13015);
or U13353 (N_13353,N_13077,N_13159);
nand U13354 (N_13354,N_13071,N_13138);
and U13355 (N_13355,N_13171,N_13056);
xor U13356 (N_13356,N_13103,N_13179);
and U13357 (N_13357,N_13129,N_13063);
nand U13358 (N_13358,N_13056,N_13058);
and U13359 (N_13359,N_13074,N_13138);
xnor U13360 (N_13360,N_13156,N_13066);
nand U13361 (N_13361,N_13132,N_13034);
and U13362 (N_13362,N_13171,N_13180);
and U13363 (N_13363,N_13134,N_13053);
nand U13364 (N_13364,N_13158,N_13130);
and U13365 (N_13365,N_13092,N_13157);
nor U13366 (N_13366,N_13004,N_13028);
nand U13367 (N_13367,N_13187,N_13025);
and U13368 (N_13368,N_13116,N_13175);
nand U13369 (N_13369,N_13115,N_13178);
and U13370 (N_13370,N_13036,N_13165);
nor U13371 (N_13371,N_13142,N_13126);
and U13372 (N_13372,N_13030,N_13164);
nor U13373 (N_13373,N_13016,N_13038);
or U13374 (N_13374,N_13113,N_13175);
nor U13375 (N_13375,N_13171,N_13060);
xor U13376 (N_13376,N_13144,N_13004);
and U13377 (N_13377,N_13179,N_13186);
and U13378 (N_13378,N_13186,N_13138);
xor U13379 (N_13379,N_13039,N_13137);
xor U13380 (N_13380,N_13117,N_13137);
and U13381 (N_13381,N_13184,N_13069);
and U13382 (N_13382,N_13115,N_13008);
nor U13383 (N_13383,N_13177,N_13086);
nor U13384 (N_13384,N_13052,N_13072);
nor U13385 (N_13385,N_13148,N_13193);
nor U13386 (N_13386,N_13037,N_13141);
and U13387 (N_13387,N_13064,N_13198);
or U13388 (N_13388,N_13008,N_13037);
or U13389 (N_13389,N_13030,N_13141);
nor U13390 (N_13390,N_13003,N_13154);
or U13391 (N_13391,N_13102,N_13128);
nand U13392 (N_13392,N_13038,N_13004);
or U13393 (N_13393,N_13055,N_13079);
xnor U13394 (N_13394,N_13010,N_13102);
nor U13395 (N_13395,N_13081,N_13057);
xor U13396 (N_13396,N_13183,N_13112);
nor U13397 (N_13397,N_13190,N_13188);
nand U13398 (N_13398,N_13193,N_13117);
and U13399 (N_13399,N_13077,N_13009);
and U13400 (N_13400,N_13364,N_13229);
xnor U13401 (N_13401,N_13264,N_13284);
nor U13402 (N_13402,N_13317,N_13215);
or U13403 (N_13403,N_13203,N_13230);
and U13404 (N_13404,N_13385,N_13245);
nor U13405 (N_13405,N_13321,N_13318);
or U13406 (N_13406,N_13362,N_13337);
or U13407 (N_13407,N_13239,N_13236);
nor U13408 (N_13408,N_13292,N_13212);
nand U13409 (N_13409,N_13383,N_13240);
nand U13410 (N_13410,N_13251,N_13228);
xor U13411 (N_13411,N_13387,N_13370);
nand U13412 (N_13412,N_13344,N_13270);
or U13413 (N_13413,N_13269,N_13331);
xnor U13414 (N_13414,N_13329,N_13361);
and U13415 (N_13415,N_13297,N_13231);
nand U13416 (N_13416,N_13375,N_13306);
and U13417 (N_13417,N_13369,N_13273);
and U13418 (N_13418,N_13341,N_13382);
or U13419 (N_13419,N_13290,N_13340);
nor U13420 (N_13420,N_13254,N_13350);
nand U13421 (N_13421,N_13255,N_13305);
nor U13422 (N_13422,N_13399,N_13267);
nor U13423 (N_13423,N_13276,N_13288);
or U13424 (N_13424,N_13293,N_13384);
nor U13425 (N_13425,N_13334,N_13304);
or U13426 (N_13426,N_13286,N_13338);
xnor U13427 (N_13427,N_13394,N_13398);
xor U13428 (N_13428,N_13249,N_13241);
xnor U13429 (N_13429,N_13295,N_13223);
and U13430 (N_13430,N_13280,N_13393);
and U13431 (N_13431,N_13376,N_13265);
nor U13432 (N_13432,N_13257,N_13386);
nor U13433 (N_13433,N_13396,N_13388);
nand U13434 (N_13434,N_13234,N_13221);
nor U13435 (N_13435,N_13374,N_13314);
nand U13436 (N_13436,N_13253,N_13200);
or U13437 (N_13437,N_13335,N_13237);
nor U13438 (N_13438,N_13354,N_13258);
nor U13439 (N_13439,N_13353,N_13323);
or U13440 (N_13440,N_13242,N_13207);
and U13441 (N_13441,N_13302,N_13325);
nand U13442 (N_13442,N_13328,N_13281);
nor U13443 (N_13443,N_13220,N_13345);
nor U13444 (N_13444,N_13360,N_13232);
nand U13445 (N_13445,N_13282,N_13308);
and U13446 (N_13446,N_13377,N_13392);
and U13447 (N_13447,N_13209,N_13256);
nor U13448 (N_13448,N_13247,N_13205);
nand U13449 (N_13449,N_13227,N_13271);
or U13450 (N_13450,N_13274,N_13378);
or U13451 (N_13451,N_13252,N_13372);
xor U13452 (N_13452,N_13349,N_13355);
xor U13453 (N_13453,N_13332,N_13397);
xor U13454 (N_13454,N_13246,N_13285);
or U13455 (N_13455,N_13366,N_13298);
or U13456 (N_13456,N_13358,N_13300);
xnor U13457 (N_13457,N_13216,N_13336);
nor U13458 (N_13458,N_13356,N_13311);
or U13459 (N_13459,N_13206,N_13294);
and U13460 (N_13460,N_13275,N_13390);
nand U13461 (N_13461,N_13208,N_13243);
or U13462 (N_13462,N_13233,N_13333);
nand U13463 (N_13463,N_13266,N_13214);
xor U13464 (N_13464,N_13248,N_13277);
or U13465 (N_13465,N_13201,N_13299);
and U13466 (N_13466,N_13368,N_13222);
and U13467 (N_13467,N_13316,N_13309);
xor U13468 (N_13468,N_13301,N_13389);
nor U13469 (N_13469,N_13307,N_13296);
or U13470 (N_13470,N_13313,N_13315);
and U13471 (N_13471,N_13278,N_13367);
and U13472 (N_13472,N_13226,N_13204);
xor U13473 (N_13473,N_13263,N_13289);
and U13474 (N_13474,N_13224,N_13244);
nand U13475 (N_13475,N_13381,N_13268);
xor U13476 (N_13476,N_13272,N_13351);
nand U13477 (N_13477,N_13373,N_13217);
xor U13478 (N_13478,N_13202,N_13283);
and U13479 (N_13479,N_13347,N_13346);
and U13480 (N_13480,N_13303,N_13395);
xnor U13481 (N_13481,N_13262,N_13322);
or U13482 (N_13482,N_13259,N_13210);
and U13483 (N_13483,N_13213,N_13348);
or U13484 (N_13484,N_13339,N_13219);
or U13485 (N_13485,N_13279,N_13238);
nand U13486 (N_13486,N_13357,N_13291);
and U13487 (N_13487,N_13327,N_13250);
nand U13488 (N_13488,N_13235,N_13312);
or U13489 (N_13489,N_13287,N_13319);
and U13490 (N_13490,N_13343,N_13310);
and U13491 (N_13491,N_13365,N_13342);
nor U13492 (N_13492,N_13330,N_13371);
or U13493 (N_13493,N_13380,N_13211);
xnor U13494 (N_13494,N_13218,N_13359);
and U13495 (N_13495,N_13320,N_13260);
nand U13496 (N_13496,N_13363,N_13225);
xnor U13497 (N_13497,N_13391,N_13352);
nor U13498 (N_13498,N_13379,N_13324);
xor U13499 (N_13499,N_13261,N_13326);
nand U13500 (N_13500,N_13238,N_13209);
or U13501 (N_13501,N_13229,N_13379);
nand U13502 (N_13502,N_13280,N_13258);
and U13503 (N_13503,N_13348,N_13390);
or U13504 (N_13504,N_13226,N_13314);
nand U13505 (N_13505,N_13307,N_13286);
or U13506 (N_13506,N_13231,N_13381);
nand U13507 (N_13507,N_13239,N_13251);
nand U13508 (N_13508,N_13342,N_13270);
and U13509 (N_13509,N_13258,N_13235);
xnor U13510 (N_13510,N_13313,N_13210);
xnor U13511 (N_13511,N_13276,N_13336);
nor U13512 (N_13512,N_13294,N_13287);
or U13513 (N_13513,N_13235,N_13297);
xnor U13514 (N_13514,N_13274,N_13375);
xor U13515 (N_13515,N_13226,N_13240);
nand U13516 (N_13516,N_13391,N_13389);
and U13517 (N_13517,N_13395,N_13289);
xnor U13518 (N_13518,N_13267,N_13252);
and U13519 (N_13519,N_13360,N_13398);
nand U13520 (N_13520,N_13372,N_13212);
nand U13521 (N_13521,N_13275,N_13397);
nor U13522 (N_13522,N_13346,N_13398);
and U13523 (N_13523,N_13382,N_13258);
nand U13524 (N_13524,N_13357,N_13252);
or U13525 (N_13525,N_13268,N_13223);
or U13526 (N_13526,N_13222,N_13353);
nor U13527 (N_13527,N_13214,N_13309);
or U13528 (N_13528,N_13206,N_13309);
and U13529 (N_13529,N_13232,N_13251);
or U13530 (N_13530,N_13275,N_13203);
or U13531 (N_13531,N_13246,N_13308);
and U13532 (N_13532,N_13215,N_13345);
nor U13533 (N_13533,N_13251,N_13300);
xnor U13534 (N_13534,N_13336,N_13289);
or U13535 (N_13535,N_13391,N_13331);
or U13536 (N_13536,N_13380,N_13210);
xor U13537 (N_13537,N_13236,N_13293);
nor U13538 (N_13538,N_13305,N_13258);
and U13539 (N_13539,N_13338,N_13242);
nor U13540 (N_13540,N_13275,N_13286);
xor U13541 (N_13541,N_13391,N_13222);
nor U13542 (N_13542,N_13247,N_13308);
nor U13543 (N_13543,N_13332,N_13316);
xor U13544 (N_13544,N_13255,N_13257);
nor U13545 (N_13545,N_13246,N_13248);
nand U13546 (N_13546,N_13367,N_13222);
xor U13547 (N_13547,N_13348,N_13242);
nor U13548 (N_13548,N_13346,N_13307);
nor U13549 (N_13549,N_13308,N_13208);
and U13550 (N_13550,N_13284,N_13305);
xor U13551 (N_13551,N_13261,N_13300);
nor U13552 (N_13552,N_13331,N_13316);
xnor U13553 (N_13553,N_13270,N_13210);
or U13554 (N_13554,N_13227,N_13252);
xnor U13555 (N_13555,N_13399,N_13300);
xnor U13556 (N_13556,N_13396,N_13236);
nand U13557 (N_13557,N_13290,N_13272);
nand U13558 (N_13558,N_13257,N_13323);
nand U13559 (N_13559,N_13354,N_13255);
or U13560 (N_13560,N_13205,N_13312);
or U13561 (N_13561,N_13367,N_13223);
nand U13562 (N_13562,N_13394,N_13261);
or U13563 (N_13563,N_13261,N_13228);
xnor U13564 (N_13564,N_13349,N_13321);
nand U13565 (N_13565,N_13245,N_13282);
or U13566 (N_13566,N_13240,N_13232);
nor U13567 (N_13567,N_13292,N_13254);
nor U13568 (N_13568,N_13365,N_13390);
and U13569 (N_13569,N_13351,N_13363);
nand U13570 (N_13570,N_13303,N_13216);
or U13571 (N_13571,N_13382,N_13367);
or U13572 (N_13572,N_13284,N_13365);
nand U13573 (N_13573,N_13363,N_13320);
or U13574 (N_13574,N_13320,N_13241);
nor U13575 (N_13575,N_13305,N_13384);
nand U13576 (N_13576,N_13287,N_13358);
xor U13577 (N_13577,N_13309,N_13325);
nand U13578 (N_13578,N_13311,N_13393);
nand U13579 (N_13579,N_13318,N_13326);
and U13580 (N_13580,N_13308,N_13256);
nor U13581 (N_13581,N_13378,N_13364);
or U13582 (N_13582,N_13265,N_13369);
xnor U13583 (N_13583,N_13369,N_13232);
and U13584 (N_13584,N_13363,N_13204);
nor U13585 (N_13585,N_13227,N_13248);
nor U13586 (N_13586,N_13397,N_13297);
nor U13587 (N_13587,N_13255,N_13224);
nand U13588 (N_13588,N_13374,N_13264);
or U13589 (N_13589,N_13225,N_13325);
and U13590 (N_13590,N_13220,N_13344);
nand U13591 (N_13591,N_13277,N_13349);
nor U13592 (N_13592,N_13208,N_13281);
or U13593 (N_13593,N_13362,N_13386);
and U13594 (N_13594,N_13209,N_13325);
nor U13595 (N_13595,N_13336,N_13226);
xnor U13596 (N_13596,N_13277,N_13282);
and U13597 (N_13597,N_13204,N_13331);
and U13598 (N_13598,N_13234,N_13343);
nand U13599 (N_13599,N_13322,N_13349);
nand U13600 (N_13600,N_13596,N_13400);
xor U13601 (N_13601,N_13487,N_13585);
nor U13602 (N_13602,N_13434,N_13404);
and U13603 (N_13603,N_13423,N_13550);
xor U13604 (N_13604,N_13538,N_13582);
nand U13605 (N_13605,N_13593,N_13542);
and U13606 (N_13606,N_13403,N_13548);
nand U13607 (N_13607,N_13561,N_13444);
or U13608 (N_13608,N_13409,N_13569);
nand U13609 (N_13609,N_13599,N_13432);
and U13610 (N_13610,N_13498,N_13454);
nand U13611 (N_13611,N_13420,N_13483);
nand U13612 (N_13612,N_13429,N_13441);
xnor U13613 (N_13613,N_13562,N_13502);
xor U13614 (N_13614,N_13430,N_13508);
or U13615 (N_13615,N_13473,N_13459);
nor U13616 (N_13616,N_13504,N_13500);
or U13617 (N_13617,N_13571,N_13486);
nand U13618 (N_13618,N_13476,N_13405);
nor U13619 (N_13619,N_13477,N_13590);
and U13620 (N_13620,N_13478,N_13517);
xnor U13621 (N_13621,N_13540,N_13474);
nor U13622 (N_13622,N_13446,N_13453);
xnor U13623 (N_13623,N_13445,N_13412);
nor U13624 (N_13624,N_13470,N_13431);
nand U13625 (N_13625,N_13584,N_13523);
nor U13626 (N_13626,N_13497,N_13480);
or U13627 (N_13627,N_13521,N_13435);
or U13628 (N_13628,N_13595,N_13428);
nand U13629 (N_13629,N_13531,N_13463);
and U13630 (N_13630,N_13577,N_13547);
xor U13631 (N_13631,N_13576,N_13570);
nand U13632 (N_13632,N_13482,N_13511);
or U13633 (N_13633,N_13578,N_13575);
nand U13634 (N_13634,N_13493,N_13415);
nand U13635 (N_13635,N_13447,N_13501);
xor U13636 (N_13636,N_13565,N_13568);
nand U13637 (N_13637,N_13560,N_13559);
or U13638 (N_13638,N_13468,N_13591);
nand U13639 (N_13639,N_13455,N_13489);
or U13640 (N_13640,N_13552,N_13522);
nand U13641 (N_13641,N_13472,N_13573);
and U13642 (N_13642,N_13416,N_13436);
xnor U13643 (N_13643,N_13481,N_13564);
and U13644 (N_13644,N_13469,N_13563);
and U13645 (N_13645,N_13479,N_13530);
xnor U13646 (N_13646,N_13541,N_13592);
nor U13647 (N_13647,N_13425,N_13583);
nand U13648 (N_13648,N_13465,N_13555);
xnor U13649 (N_13649,N_13402,N_13491);
or U13650 (N_13650,N_13461,N_13515);
nor U13651 (N_13651,N_13527,N_13533);
nor U13652 (N_13652,N_13495,N_13534);
or U13653 (N_13653,N_13572,N_13551);
nand U13654 (N_13654,N_13554,N_13464);
nand U13655 (N_13655,N_13443,N_13507);
nor U13656 (N_13656,N_13456,N_13410);
xnor U13657 (N_13657,N_13485,N_13520);
nor U13658 (N_13658,N_13494,N_13427);
nor U13659 (N_13659,N_13411,N_13496);
nand U13660 (N_13660,N_13450,N_13537);
and U13661 (N_13661,N_13525,N_13549);
nand U13662 (N_13662,N_13490,N_13509);
nor U13663 (N_13663,N_13524,N_13598);
or U13664 (N_13664,N_13516,N_13518);
nor U13665 (N_13665,N_13579,N_13492);
nor U13666 (N_13666,N_13407,N_13536);
or U13667 (N_13667,N_13586,N_13544);
nand U13668 (N_13668,N_13421,N_13514);
and U13669 (N_13669,N_13546,N_13528);
and U13670 (N_13670,N_13581,N_13557);
xor U13671 (N_13671,N_13597,N_13401);
xor U13672 (N_13672,N_13457,N_13566);
xnor U13673 (N_13673,N_13535,N_13466);
xor U13674 (N_13674,N_13589,N_13408);
nand U13675 (N_13675,N_13422,N_13574);
nand U13676 (N_13676,N_13499,N_13558);
xor U13677 (N_13677,N_13567,N_13440);
nand U13678 (N_13678,N_13418,N_13471);
nand U13679 (N_13679,N_13594,N_13451);
or U13680 (N_13680,N_13462,N_13529);
nor U13681 (N_13681,N_13460,N_13458);
nand U13682 (N_13682,N_13510,N_13503);
xor U13683 (N_13683,N_13513,N_13413);
xor U13684 (N_13684,N_13406,N_13448);
nor U13685 (N_13685,N_13475,N_13419);
or U13686 (N_13686,N_13433,N_13484);
and U13687 (N_13687,N_13426,N_13532);
or U13688 (N_13688,N_13545,N_13556);
xor U13689 (N_13689,N_13452,N_13588);
nor U13690 (N_13690,N_13505,N_13424);
and U13691 (N_13691,N_13437,N_13587);
and U13692 (N_13692,N_13512,N_13442);
and U13693 (N_13693,N_13417,N_13539);
nand U13694 (N_13694,N_13543,N_13506);
nor U13695 (N_13695,N_13467,N_13488);
or U13696 (N_13696,N_13519,N_13553);
nor U13697 (N_13697,N_13439,N_13580);
xor U13698 (N_13698,N_13526,N_13414);
or U13699 (N_13699,N_13449,N_13438);
xnor U13700 (N_13700,N_13599,N_13532);
or U13701 (N_13701,N_13415,N_13471);
and U13702 (N_13702,N_13562,N_13578);
nand U13703 (N_13703,N_13491,N_13487);
and U13704 (N_13704,N_13590,N_13464);
nand U13705 (N_13705,N_13401,N_13446);
nor U13706 (N_13706,N_13530,N_13424);
xnor U13707 (N_13707,N_13541,N_13452);
nor U13708 (N_13708,N_13425,N_13512);
and U13709 (N_13709,N_13405,N_13487);
xnor U13710 (N_13710,N_13439,N_13536);
nor U13711 (N_13711,N_13465,N_13476);
or U13712 (N_13712,N_13414,N_13534);
nand U13713 (N_13713,N_13482,N_13447);
and U13714 (N_13714,N_13570,N_13425);
nand U13715 (N_13715,N_13544,N_13582);
nand U13716 (N_13716,N_13427,N_13404);
nor U13717 (N_13717,N_13460,N_13581);
or U13718 (N_13718,N_13453,N_13516);
xor U13719 (N_13719,N_13562,N_13508);
or U13720 (N_13720,N_13574,N_13464);
or U13721 (N_13721,N_13530,N_13501);
nand U13722 (N_13722,N_13544,N_13588);
xnor U13723 (N_13723,N_13440,N_13582);
and U13724 (N_13724,N_13517,N_13578);
or U13725 (N_13725,N_13483,N_13434);
or U13726 (N_13726,N_13580,N_13549);
nor U13727 (N_13727,N_13455,N_13425);
or U13728 (N_13728,N_13473,N_13513);
nand U13729 (N_13729,N_13475,N_13597);
nor U13730 (N_13730,N_13438,N_13555);
or U13731 (N_13731,N_13416,N_13415);
and U13732 (N_13732,N_13421,N_13518);
nand U13733 (N_13733,N_13531,N_13410);
nand U13734 (N_13734,N_13524,N_13447);
nor U13735 (N_13735,N_13405,N_13564);
nor U13736 (N_13736,N_13459,N_13599);
or U13737 (N_13737,N_13551,N_13534);
or U13738 (N_13738,N_13442,N_13410);
or U13739 (N_13739,N_13594,N_13479);
or U13740 (N_13740,N_13468,N_13400);
nor U13741 (N_13741,N_13475,N_13415);
nand U13742 (N_13742,N_13420,N_13469);
nor U13743 (N_13743,N_13564,N_13403);
or U13744 (N_13744,N_13592,N_13428);
nand U13745 (N_13745,N_13470,N_13500);
xor U13746 (N_13746,N_13464,N_13567);
nand U13747 (N_13747,N_13461,N_13525);
nand U13748 (N_13748,N_13557,N_13442);
and U13749 (N_13749,N_13472,N_13513);
or U13750 (N_13750,N_13587,N_13417);
xor U13751 (N_13751,N_13546,N_13447);
and U13752 (N_13752,N_13437,N_13498);
nor U13753 (N_13753,N_13516,N_13595);
and U13754 (N_13754,N_13507,N_13470);
or U13755 (N_13755,N_13402,N_13483);
and U13756 (N_13756,N_13421,N_13440);
nor U13757 (N_13757,N_13467,N_13402);
or U13758 (N_13758,N_13516,N_13527);
and U13759 (N_13759,N_13573,N_13566);
nor U13760 (N_13760,N_13595,N_13517);
or U13761 (N_13761,N_13597,N_13559);
and U13762 (N_13762,N_13442,N_13526);
or U13763 (N_13763,N_13418,N_13512);
or U13764 (N_13764,N_13407,N_13414);
nor U13765 (N_13765,N_13596,N_13552);
xor U13766 (N_13766,N_13591,N_13578);
nor U13767 (N_13767,N_13569,N_13550);
nand U13768 (N_13768,N_13439,N_13503);
and U13769 (N_13769,N_13597,N_13571);
xnor U13770 (N_13770,N_13534,N_13588);
and U13771 (N_13771,N_13523,N_13565);
nor U13772 (N_13772,N_13441,N_13403);
nand U13773 (N_13773,N_13548,N_13583);
nand U13774 (N_13774,N_13464,N_13480);
nor U13775 (N_13775,N_13560,N_13581);
nor U13776 (N_13776,N_13573,N_13538);
or U13777 (N_13777,N_13460,N_13507);
nor U13778 (N_13778,N_13435,N_13529);
nor U13779 (N_13779,N_13525,N_13448);
xnor U13780 (N_13780,N_13463,N_13464);
or U13781 (N_13781,N_13451,N_13568);
and U13782 (N_13782,N_13475,N_13448);
or U13783 (N_13783,N_13401,N_13545);
nor U13784 (N_13784,N_13465,N_13420);
nor U13785 (N_13785,N_13584,N_13472);
and U13786 (N_13786,N_13579,N_13462);
and U13787 (N_13787,N_13411,N_13536);
nor U13788 (N_13788,N_13470,N_13545);
and U13789 (N_13789,N_13586,N_13419);
or U13790 (N_13790,N_13555,N_13527);
xor U13791 (N_13791,N_13407,N_13540);
nor U13792 (N_13792,N_13484,N_13489);
or U13793 (N_13793,N_13489,N_13594);
or U13794 (N_13794,N_13576,N_13512);
xnor U13795 (N_13795,N_13556,N_13473);
nor U13796 (N_13796,N_13433,N_13440);
nor U13797 (N_13797,N_13559,N_13450);
xnor U13798 (N_13798,N_13430,N_13403);
xnor U13799 (N_13799,N_13530,N_13435);
xnor U13800 (N_13800,N_13698,N_13726);
or U13801 (N_13801,N_13658,N_13770);
xor U13802 (N_13802,N_13661,N_13614);
nand U13803 (N_13803,N_13624,N_13704);
and U13804 (N_13804,N_13749,N_13687);
and U13805 (N_13805,N_13662,N_13689);
and U13806 (N_13806,N_13609,N_13620);
or U13807 (N_13807,N_13743,N_13762);
nand U13808 (N_13808,N_13722,N_13744);
nand U13809 (N_13809,N_13653,N_13767);
or U13810 (N_13810,N_13669,N_13768);
and U13811 (N_13811,N_13606,N_13707);
or U13812 (N_13812,N_13626,N_13633);
nand U13813 (N_13813,N_13725,N_13637);
or U13814 (N_13814,N_13763,N_13772);
nand U13815 (N_13815,N_13607,N_13643);
nand U13816 (N_13816,N_13747,N_13769);
or U13817 (N_13817,N_13655,N_13636);
and U13818 (N_13818,N_13667,N_13730);
nand U13819 (N_13819,N_13791,N_13714);
and U13820 (N_13820,N_13660,N_13797);
nor U13821 (N_13821,N_13746,N_13638);
or U13822 (N_13822,N_13649,N_13748);
nor U13823 (N_13823,N_13779,N_13732);
or U13824 (N_13824,N_13654,N_13647);
xor U13825 (N_13825,N_13682,N_13799);
xor U13826 (N_13826,N_13758,N_13639);
nand U13827 (N_13827,N_13645,N_13603);
and U13828 (N_13828,N_13793,N_13776);
nand U13829 (N_13829,N_13604,N_13712);
xnor U13830 (N_13830,N_13617,N_13677);
or U13831 (N_13831,N_13668,N_13690);
or U13832 (N_13832,N_13724,N_13720);
or U13833 (N_13833,N_13740,N_13723);
nor U13834 (N_13834,N_13728,N_13782);
xnor U13835 (N_13835,N_13641,N_13702);
xor U13836 (N_13836,N_13703,N_13798);
nor U13837 (N_13837,N_13678,N_13775);
nor U13838 (N_13838,N_13651,N_13789);
nand U13839 (N_13839,N_13680,N_13737);
nor U13840 (N_13840,N_13771,N_13627);
nand U13841 (N_13841,N_13623,N_13686);
nor U13842 (N_13842,N_13628,N_13709);
nand U13843 (N_13843,N_13759,N_13729);
or U13844 (N_13844,N_13656,N_13630);
and U13845 (N_13845,N_13664,N_13670);
or U13846 (N_13846,N_13688,N_13773);
xnor U13847 (N_13847,N_13784,N_13706);
nor U13848 (N_13848,N_13665,N_13684);
or U13849 (N_13849,N_13629,N_13766);
nand U13850 (N_13850,N_13650,N_13632);
or U13851 (N_13851,N_13781,N_13674);
xnor U13852 (N_13852,N_13774,N_13696);
and U13853 (N_13853,N_13635,N_13701);
and U13854 (N_13854,N_13676,N_13608);
nor U13855 (N_13855,N_13765,N_13700);
nand U13856 (N_13856,N_13794,N_13716);
nor U13857 (N_13857,N_13754,N_13710);
or U13858 (N_13858,N_13646,N_13659);
and U13859 (N_13859,N_13634,N_13652);
or U13860 (N_13860,N_13605,N_13741);
nand U13861 (N_13861,N_13760,N_13622);
or U13862 (N_13862,N_13751,N_13672);
nand U13863 (N_13863,N_13691,N_13601);
nand U13864 (N_13864,N_13618,N_13619);
xnor U13865 (N_13865,N_13752,N_13734);
nand U13866 (N_13866,N_13764,N_13699);
xor U13867 (N_13867,N_13785,N_13621);
nand U13868 (N_13868,N_13761,N_13692);
nor U13869 (N_13869,N_13657,N_13612);
and U13870 (N_13870,N_13695,N_13648);
nor U13871 (N_13871,N_13640,N_13790);
xor U13872 (N_13872,N_13625,N_13739);
xnor U13873 (N_13873,N_13671,N_13611);
and U13874 (N_13874,N_13733,N_13600);
nor U13875 (N_13875,N_13780,N_13717);
and U13876 (N_13876,N_13792,N_13738);
xor U13877 (N_13877,N_13745,N_13750);
nor U13878 (N_13878,N_13788,N_13679);
nand U13879 (N_13879,N_13718,N_13719);
nor U13880 (N_13880,N_13783,N_13777);
nand U13881 (N_13881,N_13711,N_13715);
or U13882 (N_13882,N_13778,N_13673);
nand U13883 (N_13883,N_13685,N_13755);
nor U13884 (N_13884,N_13795,N_13757);
nor U13885 (N_13885,N_13731,N_13683);
or U13886 (N_13886,N_13610,N_13693);
or U13887 (N_13887,N_13796,N_13786);
or U13888 (N_13888,N_13756,N_13705);
or U13889 (N_13889,N_13713,N_13616);
xor U13890 (N_13890,N_13708,N_13694);
nand U13891 (N_13891,N_13721,N_13697);
nor U13892 (N_13892,N_13642,N_13742);
xor U13893 (N_13893,N_13753,N_13735);
and U13894 (N_13894,N_13602,N_13666);
xor U13895 (N_13895,N_13615,N_13675);
and U13896 (N_13896,N_13736,N_13631);
nand U13897 (N_13897,N_13787,N_13644);
xor U13898 (N_13898,N_13613,N_13727);
or U13899 (N_13899,N_13681,N_13663);
nand U13900 (N_13900,N_13688,N_13601);
nor U13901 (N_13901,N_13698,N_13623);
nand U13902 (N_13902,N_13665,N_13701);
nor U13903 (N_13903,N_13708,N_13665);
and U13904 (N_13904,N_13713,N_13680);
and U13905 (N_13905,N_13778,N_13711);
or U13906 (N_13906,N_13730,N_13755);
and U13907 (N_13907,N_13660,N_13754);
or U13908 (N_13908,N_13762,N_13746);
nand U13909 (N_13909,N_13691,N_13668);
nand U13910 (N_13910,N_13624,N_13764);
and U13911 (N_13911,N_13630,N_13712);
and U13912 (N_13912,N_13730,N_13642);
xor U13913 (N_13913,N_13791,N_13660);
or U13914 (N_13914,N_13695,N_13688);
and U13915 (N_13915,N_13623,N_13601);
and U13916 (N_13916,N_13671,N_13663);
or U13917 (N_13917,N_13707,N_13779);
xnor U13918 (N_13918,N_13787,N_13759);
nand U13919 (N_13919,N_13607,N_13644);
nor U13920 (N_13920,N_13741,N_13786);
xnor U13921 (N_13921,N_13657,N_13635);
nor U13922 (N_13922,N_13634,N_13789);
and U13923 (N_13923,N_13743,N_13757);
xnor U13924 (N_13924,N_13676,N_13750);
xnor U13925 (N_13925,N_13644,N_13715);
xnor U13926 (N_13926,N_13687,N_13615);
or U13927 (N_13927,N_13720,N_13625);
xnor U13928 (N_13928,N_13725,N_13645);
or U13929 (N_13929,N_13611,N_13758);
nor U13930 (N_13930,N_13791,N_13673);
nand U13931 (N_13931,N_13633,N_13788);
and U13932 (N_13932,N_13644,N_13762);
or U13933 (N_13933,N_13637,N_13681);
nand U13934 (N_13934,N_13782,N_13620);
and U13935 (N_13935,N_13777,N_13637);
or U13936 (N_13936,N_13696,N_13622);
nor U13937 (N_13937,N_13635,N_13659);
xnor U13938 (N_13938,N_13735,N_13691);
nand U13939 (N_13939,N_13729,N_13781);
and U13940 (N_13940,N_13769,N_13765);
nor U13941 (N_13941,N_13693,N_13680);
xnor U13942 (N_13942,N_13756,N_13645);
nand U13943 (N_13943,N_13759,N_13629);
nand U13944 (N_13944,N_13770,N_13739);
nand U13945 (N_13945,N_13689,N_13724);
and U13946 (N_13946,N_13648,N_13799);
or U13947 (N_13947,N_13679,N_13616);
nand U13948 (N_13948,N_13684,N_13681);
nand U13949 (N_13949,N_13736,N_13695);
or U13950 (N_13950,N_13798,N_13615);
or U13951 (N_13951,N_13778,N_13729);
and U13952 (N_13952,N_13646,N_13779);
xor U13953 (N_13953,N_13699,N_13794);
nor U13954 (N_13954,N_13685,N_13703);
nor U13955 (N_13955,N_13765,N_13643);
nand U13956 (N_13956,N_13624,N_13693);
xor U13957 (N_13957,N_13784,N_13642);
xnor U13958 (N_13958,N_13605,N_13676);
and U13959 (N_13959,N_13633,N_13733);
or U13960 (N_13960,N_13739,N_13720);
nor U13961 (N_13961,N_13739,N_13634);
xnor U13962 (N_13962,N_13605,N_13744);
xnor U13963 (N_13963,N_13694,N_13666);
or U13964 (N_13964,N_13767,N_13718);
nor U13965 (N_13965,N_13666,N_13751);
xnor U13966 (N_13966,N_13601,N_13714);
or U13967 (N_13967,N_13668,N_13744);
nor U13968 (N_13968,N_13653,N_13624);
or U13969 (N_13969,N_13690,N_13763);
nor U13970 (N_13970,N_13729,N_13725);
nor U13971 (N_13971,N_13770,N_13745);
or U13972 (N_13972,N_13675,N_13639);
xor U13973 (N_13973,N_13679,N_13685);
or U13974 (N_13974,N_13756,N_13602);
nor U13975 (N_13975,N_13695,N_13616);
nand U13976 (N_13976,N_13791,N_13662);
nor U13977 (N_13977,N_13654,N_13642);
xnor U13978 (N_13978,N_13697,N_13718);
xor U13979 (N_13979,N_13651,N_13695);
or U13980 (N_13980,N_13678,N_13740);
nand U13981 (N_13981,N_13768,N_13631);
xnor U13982 (N_13982,N_13685,N_13652);
or U13983 (N_13983,N_13784,N_13723);
nand U13984 (N_13984,N_13773,N_13735);
nand U13985 (N_13985,N_13739,N_13702);
and U13986 (N_13986,N_13672,N_13727);
nor U13987 (N_13987,N_13630,N_13620);
and U13988 (N_13988,N_13725,N_13642);
nand U13989 (N_13989,N_13652,N_13754);
or U13990 (N_13990,N_13717,N_13772);
or U13991 (N_13991,N_13766,N_13641);
and U13992 (N_13992,N_13691,N_13634);
nand U13993 (N_13993,N_13700,N_13724);
xor U13994 (N_13994,N_13788,N_13684);
and U13995 (N_13995,N_13738,N_13784);
xnor U13996 (N_13996,N_13671,N_13748);
xor U13997 (N_13997,N_13622,N_13691);
or U13998 (N_13998,N_13695,N_13701);
or U13999 (N_13999,N_13611,N_13763);
xor U14000 (N_14000,N_13957,N_13872);
and U14001 (N_14001,N_13803,N_13920);
and U14002 (N_14002,N_13989,N_13999);
and U14003 (N_14003,N_13990,N_13810);
nor U14004 (N_14004,N_13862,N_13868);
xor U14005 (N_14005,N_13801,N_13972);
nand U14006 (N_14006,N_13958,N_13848);
nand U14007 (N_14007,N_13996,N_13968);
and U14008 (N_14008,N_13973,N_13829);
nand U14009 (N_14009,N_13870,N_13952);
and U14010 (N_14010,N_13809,N_13910);
nand U14011 (N_14011,N_13974,N_13885);
and U14012 (N_14012,N_13914,N_13962);
and U14013 (N_14013,N_13867,N_13964);
nor U14014 (N_14014,N_13844,N_13992);
xor U14015 (N_14015,N_13811,N_13971);
nor U14016 (N_14016,N_13942,N_13921);
nand U14017 (N_14017,N_13976,N_13800);
or U14018 (N_14018,N_13877,N_13986);
and U14019 (N_14019,N_13951,N_13836);
or U14020 (N_14020,N_13997,N_13837);
xnor U14021 (N_14021,N_13915,N_13939);
nor U14022 (N_14022,N_13938,N_13859);
or U14023 (N_14023,N_13961,N_13948);
and U14024 (N_14024,N_13852,N_13869);
or U14025 (N_14025,N_13984,N_13988);
or U14026 (N_14026,N_13830,N_13846);
or U14027 (N_14027,N_13955,N_13930);
and U14028 (N_14028,N_13928,N_13860);
or U14029 (N_14029,N_13900,N_13816);
or U14030 (N_14030,N_13980,N_13815);
xor U14031 (N_14031,N_13937,N_13923);
nand U14032 (N_14032,N_13904,N_13833);
and U14033 (N_14033,N_13929,N_13981);
xnor U14034 (N_14034,N_13845,N_13805);
nor U14035 (N_14035,N_13857,N_13880);
nand U14036 (N_14036,N_13934,N_13975);
or U14037 (N_14037,N_13926,N_13995);
xnor U14038 (N_14038,N_13849,N_13970);
or U14039 (N_14039,N_13899,N_13806);
and U14040 (N_14040,N_13819,N_13977);
nand U14041 (N_14041,N_13853,N_13932);
or U14042 (N_14042,N_13898,N_13931);
xnor U14043 (N_14043,N_13893,N_13828);
nand U14044 (N_14044,N_13843,N_13812);
and U14045 (N_14045,N_13823,N_13891);
xor U14046 (N_14046,N_13919,N_13922);
and U14047 (N_14047,N_13993,N_13822);
or U14048 (N_14048,N_13960,N_13905);
or U14049 (N_14049,N_13936,N_13979);
nor U14050 (N_14050,N_13945,N_13876);
and U14051 (N_14051,N_13894,N_13892);
xor U14052 (N_14052,N_13835,N_13953);
nor U14053 (N_14053,N_13879,N_13987);
nand U14054 (N_14054,N_13943,N_13983);
nor U14055 (N_14055,N_13969,N_13839);
nand U14056 (N_14056,N_13924,N_13890);
xor U14057 (N_14057,N_13933,N_13826);
xor U14058 (N_14058,N_13861,N_13820);
nor U14059 (N_14059,N_13991,N_13950);
nor U14060 (N_14060,N_13827,N_13918);
and U14061 (N_14061,N_13818,N_13956);
xnor U14062 (N_14062,N_13927,N_13998);
and U14063 (N_14063,N_13886,N_13832);
xor U14064 (N_14064,N_13874,N_13831);
and U14065 (N_14065,N_13947,N_13944);
or U14066 (N_14066,N_13871,N_13949);
or U14067 (N_14067,N_13912,N_13881);
or U14068 (N_14068,N_13908,N_13911);
or U14069 (N_14069,N_13935,N_13834);
and U14070 (N_14070,N_13946,N_13873);
or U14071 (N_14071,N_13994,N_13907);
or U14072 (N_14072,N_13856,N_13913);
xor U14073 (N_14073,N_13917,N_13840);
nand U14074 (N_14074,N_13909,N_13889);
or U14075 (N_14075,N_13850,N_13825);
and U14076 (N_14076,N_13883,N_13821);
nand U14077 (N_14077,N_13851,N_13941);
or U14078 (N_14078,N_13884,N_13863);
nor U14079 (N_14079,N_13804,N_13940);
and U14080 (N_14080,N_13966,N_13978);
or U14081 (N_14081,N_13982,N_13967);
nor U14082 (N_14082,N_13813,N_13965);
and U14083 (N_14083,N_13817,N_13985);
or U14084 (N_14084,N_13897,N_13864);
nor U14085 (N_14085,N_13808,N_13895);
and U14086 (N_14086,N_13802,N_13847);
nor U14087 (N_14087,N_13882,N_13896);
or U14088 (N_14088,N_13858,N_13824);
or U14089 (N_14089,N_13901,N_13842);
and U14090 (N_14090,N_13903,N_13925);
and U14091 (N_14091,N_13841,N_13902);
xnor U14092 (N_14092,N_13855,N_13838);
nor U14093 (N_14093,N_13865,N_13959);
xnor U14094 (N_14094,N_13807,N_13916);
or U14095 (N_14095,N_13854,N_13875);
xor U14096 (N_14096,N_13906,N_13954);
xor U14097 (N_14097,N_13963,N_13888);
or U14098 (N_14098,N_13878,N_13866);
and U14099 (N_14099,N_13814,N_13887);
and U14100 (N_14100,N_13912,N_13907);
nor U14101 (N_14101,N_13894,N_13945);
xor U14102 (N_14102,N_13977,N_13835);
nor U14103 (N_14103,N_13892,N_13820);
xor U14104 (N_14104,N_13950,N_13820);
nor U14105 (N_14105,N_13804,N_13926);
nand U14106 (N_14106,N_13856,N_13881);
xor U14107 (N_14107,N_13855,N_13984);
xnor U14108 (N_14108,N_13936,N_13894);
nor U14109 (N_14109,N_13896,N_13836);
xnor U14110 (N_14110,N_13935,N_13830);
or U14111 (N_14111,N_13960,N_13994);
or U14112 (N_14112,N_13920,N_13965);
nand U14113 (N_14113,N_13865,N_13988);
nor U14114 (N_14114,N_13960,N_13946);
xor U14115 (N_14115,N_13820,N_13836);
nor U14116 (N_14116,N_13806,N_13821);
and U14117 (N_14117,N_13902,N_13855);
or U14118 (N_14118,N_13897,N_13992);
nor U14119 (N_14119,N_13997,N_13928);
or U14120 (N_14120,N_13932,N_13925);
nor U14121 (N_14121,N_13986,N_13855);
or U14122 (N_14122,N_13873,N_13958);
xor U14123 (N_14123,N_13916,N_13989);
nor U14124 (N_14124,N_13882,N_13990);
or U14125 (N_14125,N_13837,N_13943);
and U14126 (N_14126,N_13916,N_13991);
xor U14127 (N_14127,N_13839,N_13979);
and U14128 (N_14128,N_13808,N_13978);
nor U14129 (N_14129,N_13801,N_13911);
or U14130 (N_14130,N_13822,N_13825);
nor U14131 (N_14131,N_13962,N_13823);
xnor U14132 (N_14132,N_13860,N_13983);
xnor U14133 (N_14133,N_13881,N_13823);
nor U14134 (N_14134,N_13948,N_13815);
xnor U14135 (N_14135,N_13900,N_13918);
or U14136 (N_14136,N_13902,N_13957);
nand U14137 (N_14137,N_13976,N_13970);
nand U14138 (N_14138,N_13855,N_13817);
or U14139 (N_14139,N_13848,N_13938);
and U14140 (N_14140,N_13817,N_13847);
and U14141 (N_14141,N_13864,N_13858);
or U14142 (N_14142,N_13816,N_13956);
and U14143 (N_14143,N_13837,N_13834);
nand U14144 (N_14144,N_13931,N_13888);
nor U14145 (N_14145,N_13910,N_13828);
and U14146 (N_14146,N_13942,N_13955);
nor U14147 (N_14147,N_13813,N_13886);
xnor U14148 (N_14148,N_13919,N_13938);
and U14149 (N_14149,N_13912,N_13980);
nand U14150 (N_14150,N_13973,N_13811);
xnor U14151 (N_14151,N_13852,N_13880);
nand U14152 (N_14152,N_13846,N_13843);
nor U14153 (N_14153,N_13950,N_13807);
and U14154 (N_14154,N_13975,N_13821);
nor U14155 (N_14155,N_13824,N_13903);
nor U14156 (N_14156,N_13852,N_13942);
and U14157 (N_14157,N_13838,N_13950);
or U14158 (N_14158,N_13830,N_13882);
nand U14159 (N_14159,N_13848,N_13867);
and U14160 (N_14160,N_13856,N_13808);
nor U14161 (N_14161,N_13941,N_13976);
nand U14162 (N_14162,N_13983,N_13874);
or U14163 (N_14163,N_13961,N_13860);
xor U14164 (N_14164,N_13884,N_13822);
or U14165 (N_14165,N_13827,N_13969);
and U14166 (N_14166,N_13981,N_13932);
and U14167 (N_14167,N_13826,N_13908);
xnor U14168 (N_14168,N_13905,N_13868);
and U14169 (N_14169,N_13982,N_13992);
nand U14170 (N_14170,N_13991,N_13868);
nand U14171 (N_14171,N_13959,N_13882);
nand U14172 (N_14172,N_13848,N_13984);
nor U14173 (N_14173,N_13863,N_13818);
nand U14174 (N_14174,N_13866,N_13958);
and U14175 (N_14175,N_13936,N_13954);
nor U14176 (N_14176,N_13904,N_13993);
and U14177 (N_14177,N_13848,N_13995);
nand U14178 (N_14178,N_13936,N_13927);
and U14179 (N_14179,N_13921,N_13815);
and U14180 (N_14180,N_13982,N_13904);
or U14181 (N_14181,N_13828,N_13930);
nor U14182 (N_14182,N_13863,N_13845);
nor U14183 (N_14183,N_13918,N_13920);
xnor U14184 (N_14184,N_13969,N_13926);
nand U14185 (N_14185,N_13861,N_13858);
xor U14186 (N_14186,N_13920,N_13987);
nor U14187 (N_14187,N_13958,N_13882);
nand U14188 (N_14188,N_13835,N_13820);
xor U14189 (N_14189,N_13954,N_13951);
or U14190 (N_14190,N_13853,N_13983);
xor U14191 (N_14191,N_13860,N_13999);
and U14192 (N_14192,N_13998,N_13960);
nor U14193 (N_14193,N_13969,N_13803);
nor U14194 (N_14194,N_13922,N_13807);
nand U14195 (N_14195,N_13933,N_13815);
nor U14196 (N_14196,N_13828,N_13954);
or U14197 (N_14197,N_13895,N_13975);
nand U14198 (N_14198,N_13970,N_13860);
nand U14199 (N_14199,N_13855,N_13919);
xnor U14200 (N_14200,N_14158,N_14014);
or U14201 (N_14201,N_14010,N_14113);
xnor U14202 (N_14202,N_14072,N_14027);
or U14203 (N_14203,N_14116,N_14132);
and U14204 (N_14204,N_14109,N_14172);
and U14205 (N_14205,N_14056,N_14050);
xnor U14206 (N_14206,N_14197,N_14075);
xnor U14207 (N_14207,N_14142,N_14126);
nand U14208 (N_14208,N_14133,N_14193);
xor U14209 (N_14209,N_14022,N_14054);
xnor U14210 (N_14210,N_14057,N_14139);
nand U14211 (N_14211,N_14097,N_14157);
or U14212 (N_14212,N_14006,N_14161);
or U14213 (N_14213,N_14195,N_14007);
xnor U14214 (N_14214,N_14160,N_14173);
xnor U14215 (N_14215,N_14005,N_14047);
nor U14216 (N_14216,N_14138,N_14037);
xnor U14217 (N_14217,N_14020,N_14012);
xnor U14218 (N_14218,N_14147,N_14189);
nand U14219 (N_14219,N_14123,N_14001);
nand U14220 (N_14220,N_14103,N_14021);
nor U14221 (N_14221,N_14099,N_14073);
and U14222 (N_14222,N_14024,N_14082);
xor U14223 (N_14223,N_14069,N_14090);
xnor U14224 (N_14224,N_14034,N_14141);
nor U14225 (N_14225,N_14135,N_14087);
xor U14226 (N_14226,N_14119,N_14129);
and U14227 (N_14227,N_14148,N_14033);
or U14228 (N_14228,N_14115,N_14081);
and U14229 (N_14229,N_14002,N_14185);
nand U14230 (N_14230,N_14016,N_14156);
nand U14231 (N_14231,N_14196,N_14124);
xor U14232 (N_14232,N_14180,N_14111);
nand U14233 (N_14233,N_14074,N_14077);
nor U14234 (N_14234,N_14044,N_14192);
xnor U14235 (N_14235,N_14046,N_14182);
nor U14236 (N_14236,N_14166,N_14036);
or U14237 (N_14237,N_14155,N_14025);
xnor U14238 (N_14238,N_14093,N_14003);
nand U14239 (N_14239,N_14162,N_14144);
or U14240 (N_14240,N_14145,N_14096);
and U14241 (N_14241,N_14055,N_14105);
or U14242 (N_14242,N_14004,N_14177);
nand U14243 (N_14243,N_14110,N_14108);
nand U14244 (N_14244,N_14104,N_14154);
nand U14245 (N_14245,N_14017,N_14136);
nand U14246 (N_14246,N_14052,N_14152);
nand U14247 (N_14247,N_14041,N_14187);
xnor U14248 (N_14248,N_14053,N_14153);
nor U14249 (N_14249,N_14190,N_14080);
and U14250 (N_14250,N_14076,N_14030);
xor U14251 (N_14251,N_14092,N_14070);
or U14252 (N_14252,N_14163,N_14100);
nand U14253 (N_14253,N_14101,N_14184);
nor U14254 (N_14254,N_14062,N_14065);
xor U14255 (N_14255,N_14137,N_14178);
or U14256 (N_14256,N_14088,N_14031);
or U14257 (N_14257,N_14015,N_14067);
xnor U14258 (N_14258,N_14168,N_14169);
nor U14259 (N_14259,N_14049,N_14029);
nand U14260 (N_14260,N_14112,N_14086);
or U14261 (N_14261,N_14085,N_14198);
or U14262 (N_14262,N_14117,N_14174);
or U14263 (N_14263,N_14134,N_14051);
xnor U14264 (N_14264,N_14127,N_14165);
and U14265 (N_14265,N_14060,N_14023);
xnor U14266 (N_14266,N_14159,N_14120);
xor U14267 (N_14267,N_14058,N_14179);
and U14268 (N_14268,N_14183,N_14008);
nor U14269 (N_14269,N_14083,N_14170);
nor U14270 (N_14270,N_14151,N_14164);
or U14271 (N_14271,N_14194,N_14045);
nor U14272 (N_14272,N_14107,N_14019);
nand U14273 (N_14273,N_14094,N_14114);
and U14274 (N_14274,N_14118,N_14130);
nand U14275 (N_14275,N_14048,N_14128);
and U14276 (N_14276,N_14167,N_14098);
and U14277 (N_14277,N_14181,N_14125);
or U14278 (N_14278,N_14018,N_14039);
xnor U14279 (N_14279,N_14106,N_14071);
xor U14280 (N_14280,N_14102,N_14011);
nand U14281 (N_14281,N_14043,N_14061);
and U14282 (N_14282,N_14091,N_14143);
xor U14283 (N_14283,N_14186,N_14078);
or U14284 (N_14284,N_14191,N_14064);
nor U14285 (N_14285,N_14089,N_14084);
nor U14286 (N_14286,N_14095,N_14068);
or U14287 (N_14287,N_14063,N_14032);
xor U14288 (N_14288,N_14038,N_14013);
nand U14289 (N_14289,N_14042,N_14122);
xor U14290 (N_14290,N_14188,N_14150);
and U14291 (N_14291,N_14059,N_14140);
nor U14292 (N_14292,N_14066,N_14079);
xor U14293 (N_14293,N_14146,N_14028);
xnor U14294 (N_14294,N_14175,N_14131);
xnor U14295 (N_14295,N_14121,N_14026);
xnor U14296 (N_14296,N_14176,N_14009);
nand U14297 (N_14297,N_14040,N_14171);
and U14298 (N_14298,N_14199,N_14000);
xor U14299 (N_14299,N_14035,N_14149);
nand U14300 (N_14300,N_14043,N_14109);
nor U14301 (N_14301,N_14144,N_14177);
nor U14302 (N_14302,N_14108,N_14058);
nor U14303 (N_14303,N_14165,N_14097);
and U14304 (N_14304,N_14088,N_14008);
and U14305 (N_14305,N_14079,N_14022);
nor U14306 (N_14306,N_14181,N_14121);
and U14307 (N_14307,N_14070,N_14154);
xor U14308 (N_14308,N_14128,N_14107);
and U14309 (N_14309,N_14046,N_14131);
nand U14310 (N_14310,N_14148,N_14155);
or U14311 (N_14311,N_14135,N_14050);
and U14312 (N_14312,N_14080,N_14051);
nand U14313 (N_14313,N_14180,N_14166);
or U14314 (N_14314,N_14146,N_14071);
xnor U14315 (N_14315,N_14001,N_14002);
nand U14316 (N_14316,N_14017,N_14188);
xor U14317 (N_14317,N_14136,N_14144);
xor U14318 (N_14318,N_14019,N_14157);
xnor U14319 (N_14319,N_14014,N_14199);
nor U14320 (N_14320,N_14040,N_14155);
or U14321 (N_14321,N_14056,N_14130);
or U14322 (N_14322,N_14037,N_14118);
xor U14323 (N_14323,N_14058,N_14154);
or U14324 (N_14324,N_14018,N_14143);
and U14325 (N_14325,N_14078,N_14053);
xnor U14326 (N_14326,N_14086,N_14033);
or U14327 (N_14327,N_14189,N_14116);
xor U14328 (N_14328,N_14022,N_14136);
and U14329 (N_14329,N_14084,N_14198);
xnor U14330 (N_14330,N_14114,N_14124);
and U14331 (N_14331,N_14175,N_14092);
xor U14332 (N_14332,N_14065,N_14040);
and U14333 (N_14333,N_14097,N_14051);
and U14334 (N_14334,N_14102,N_14020);
nand U14335 (N_14335,N_14120,N_14118);
xor U14336 (N_14336,N_14117,N_14145);
nor U14337 (N_14337,N_14030,N_14164);
nand U14338 (N_14338,N_14183,N_14177);
and U14339 (N_14339,N_14198,N_14176);
xor U14340 (N_14340,N_14112,N_14166);
xor U14341 (N_14341,N_14164,N_14043);
and U14342 (N_14342,N_14191,N_14040);
nor U14343 (N_14343,N_14017,N_14071);
and U14344 (N_14344,N_14197,N_14029);
or U14345 (N_14345,N_14093,N_14021);
xnor U14346 (N_14346,N_14141,N_14010);
and U14347 (N_14347,N_14119,N_14006);
and U14348 (N_14348,N_14053,N_14076);
nand U14349 (N_14349,N_14112,N_14063);
xnor U14350 (N_14350,N_14074,N_14185);
and U14351 (N_14351,N_14036,N_14100);
xor U14352 (N_14352,N_14103,N_14185);
nor U14353 (N_14353,N_14096,N_14008);
or U14354 (N_14354,N_14139,N_14103);
or U14355 (N_14355,N_14110,N_14118);
nand U14356 (N_14356,N_14170,N_14156);
xnor U14357 (N_14357,N_14100,N_14025);
or U14358 (N_14358,N_14183,N_14028);
nor U14359 (N_14359,N_14094,N_14132);
nor U14360 (N_14360,N_14083,N_14012);
and U14361 (N_14361,N_14036,N_14149);
nand U14362 (N_14362,N_14073,N_14080);
and U14363 (N_14363,N_14180,N_14014);
nor U14364 (N_14364,N_14055,N_14081);
nand U14365 (N_14365,N_14156,N_14072);
and U14366 (N_14366,N_14103,N_14014);
nand U14367 (N_14367,N_14039,N_14173);
xor U14368 (N_14368,N_14011,N_14052);
nor U14369 (N_14369,N_14128,N_14105);
nand U14370 (N_14370,N_14029,N_14159);
or U14371 (N_14371,N_14198,N_14145);
nand U14372 (N_14372,N_14085,N_14059);
nand U14373 (N_14373,N_14070,N_14188);
xor U14374 (N_14374,N_14050,N_14125);
or U14375 (N_14375,N_14014,N_14024);
nor U14376 (N_14376,N_14143,N_14067);
and U14377 (N_14377,N_14066,N_14088);
and U14378 (N_14378,N_14103,N_14146);
or U14379 (N_14379,N_14182,N_14124);
nand U14380 (N_14380,N_14172,N_14034);
and U14381 (N_14381,N_14012,N_14142);
xnor U14382 (N_14382,N_14113,N_14045);
nand U14383 (N_14383,N_14083,N_14050);
or U14384 (N_14384,N_14074,N_14052);
xnor U14385 (N_14385,N_14119,N_14111);
and U14386 (N_14386,N_14040,N_14000);
nor U14387 (N_14387,N_14141,N_14186);
nor U14388 (N_14388,N_14091,N_14164);
or U14389 (N_14389,N_14068,N_14035);
nand U14390 (N_14390,N_14000,N_14024);
xor U14391 (N_14391,N_14094,N_14166);
and U14392 (N_14392,N_14014,N_14108);
nand U14393 (N_14393,N_14059,N_14196);
and U14394 (N_14394,N_14189,N_14107);
nand U14395 (N_14395,N_14184,N_14180);
nand U14396 (N_14396,N_14048,N_14087);
xor U14397 (N_14397,N_14039,N_14007);
and U14398 (N_14398,N_14054,N_14006);
and U14399 (N_14399,N_14177,N_14038);
nor U14400 (N_14400,N_14222,N_14237);
nor U14401 (N_14401,N_14301,N_14224);
nand U14402 (N_14402,N_14343,N_14209);
xnor U14403 (N_14403,N_14316,N_14255);
or U14404 (N_14404,N_14382,N_14306);
xor U14405 (N_14405,N_14305,N_14366);
nor U14406 (N_14406,N_14216,N_14335);
xnor U14407 (N_14407,N_14205,N_14259);
or U14408 (N_14408,N_14353,N_14210);
and U14409 (N_14409,N_14326,N_14318);
nand U14410 (N_14410,N_14311,N_14321);
xor U14411 (N_14411,N_14283,N_14264);
nor U14412 (N_14412,N_14394,N_14315);
and U14413 (N_14413,N_14284,N_14274);
xnor U14414 (N_14414,N_14341,N_14363);
nand U14415 (N_14415,N_14355,N_14360);
xor U14416 (N_14416,N_14374,N_14225);
or U14417 (N_14417,N_14215,N_14281);
nand U14418 (N_14418,N_14376,N_14300);
nand U14419 (N_14419,N_14386,N_14320);
or U14420 (N_14420,N_14354,N_14368);
and U14421 (N_14421,N_14344,N_14277);
xor U14422 (N_14422,N_14314,N_14358);
nand U14423 (N_14423,N_14251,N_14203);
xor U14424 (N_14424,N_14325,N_14240);
nor U14425 (N_14425,N_14218,N_14339);
nand U14426 (N_14426,N_14295,N_14357);
nand U14427 (N_14427,N_14219,N_14313);
or U14428 (N_14428,N_14310,N_14282);
xnor U14429 (N_14429,N_14389,N_14383);
nor U14430 (N_14430,N_14324,N_14345);
and U14431 (N_14431,N_14211,N_14204);
nand U14432 (N_14432,N_14245,N_14390);
nor U14433 (N_14433,N_14279,N_14262);
nor U14434 (N_14434,N_14228,N_14242);
nand U14435 (N_14435,N_14296,N_14328);
and U14436 (N_14436,N_14348,N_14246);
or U14437 (N_14437,N_14258,N_14298);
nor U14438 (N_14438,N_14292,N_14346);
nand U14439 (N_14439,N_14280,N_14332);
and U14440 (N_14440,N_14372,N_14220);
nor U14441 (N_14441,N_14369,N_14388);
and U14442 (N_14442,N_14391,N_14365);
nor U14443 (N_14443,N_14331,N_14289);
or U14444 (N_14444,N_14254,N_14392);
and U14445 (N_14445,N_14230,N_14309);
or U14446 (N_14446,N_14260,N_14217);
and U14447 (N_14447,N_14263,N_14380);
nand U14448 (N_14448,N_14303,N_14304);
nor U14449 (N_14449,N_14385,N_14234);
nand U14450 (N_14450,N_14239,N_14285);
nor U14451 (N_14451,N_14256,N_14379);
nand U14452 (N_14452,N_14213,N_14227);
and U14453 (N_14453,N_14247,N_14398);
or U14454 (N_14454,N_14327,N_14378);
xnor U14455 (N_14455,N_14275,N_14208);
or U14456 (N_14456,N_14322,N_14384);
nand U14457 (N_14457,N_14393,N_14317);
xor U14458 (N_14458,N_14200,N_14356);
and U14459 (N_14459,N_14248,N_14334);
and U14460 (N_14460,N_14359,N_14336);
nor U14461 (N_14461,N_14362,N_14257);
and U14462 (N_14462,N_14267,N_14207);
xnor U14463 (N_14463,N_14319,N_14243);
xnor U14464 (N_14464,N_14290,N_14202);
xor U14465 (N_14465,N_14381,N_14342);
and U14466 (N_14466,N_14308,N_14370);
xor U14467 (N_14467,N_14395,N_14250);
or U14468 (N_14468,N_14252,N_14312);
xnor U14469 (N_14469,N_14232,N_14288);
and U14470 (N_14470,N_14337,N_14291);
nand U14471 (N_14471,N_14399,N_14396);
and U14472 (N_14472,N_14397,N_14201);
nor U14473 (N_14473,N_14361,N_14278);
and U14474 (N_14474,N_14329,N_14330);
or U14475 (N_14475,N_14377,N_14235);
and U14476 (N_14476,N_14233,N_14231);
and U14477 (N_14477,N_14351,N_14387);
or U14478 (N_14478,N_14249,N_14236);
nand U14479 (N_14479,N_14273,N_14244);
nand U14480 (N_14480,N_14340,N_14261);
or U14481 (N_14481,N_14287,N_14272);
and U14482 (N_14482,N_14221,N_14212);
and U14483 (N_14483,N_14286,N_14350);
nor U14484 (N_14484,N_14367,N_14338);
nand U14485 (N_14485,N_14347,N_14294);
and U14486 (N_14486,N_14293,N_14302);
xnor U14487 (N_14487,N_14333,N_14375);
xor U14488 (N_14488,N_14253,N_14276);
nand U14489 (N_14489,N_14373,N_14352);
and U14490 (N_14490,N_14271,N_14226);
and U14491 (N_14491,N_14269,N_14223);
and U14492 (N_14492,N_14268,N_14323);
xnor U14493 (N_14493,N_14206,N_14229);
or U14494 (N_14494,N_14270,N_14307);
and U14495 (N_14495,N_14265,N_14364);
and U14496 (N_14496,N_14238,N_14241);
or U14497 (N_14497,N_14214,N_14299);
or U14498 (N_14498,N_14349,N_14297);
and U14499 (N_14499,N_14266,N_14371);
and U14500 (N_14500,N_14200,N_14333);
and U14501 (N_14501,N_14373,N_14264);
nand U14502 (N_14502,N_14295,N_14240);
nand U14503 (N_14503,N_14357,N_14324);
nor U14504 (N_14504,N_14279,N_14352);
xnor U14505 (N_14505,N_14259,N_14275);
nor U14506 (N_14506,N_14233,N_14234);
or U14507 (N_14507,N_14236,N_14393);
or U14508 (N_14508,N_14362,N_14304);
xnor U14509 (N_14509,N_14303,N_14215);
and U14510 (N_14510,N_14238,N_14376);
nand U14511 (N_14511,N_14225,N_14304);
xor U14512 (N_14512,N_14345,N_14287);
or U14513 (N_14513,N_14332,N_14266);
nand U14514 (N_14514,N_14394,N_14368);
and U14515 (N_14515,N_14217,N_14319);
nor U14516 (N_14516,N_14213,N_14334);
nand U14517 (N_14517,N_14335,N_14295);
and U14518 (N_14518,N_14318,N_14386);
and U14519 (N_14519,N_14339,N_14262);
xnor U14520 (N_14520,N_14230,N_14243);
nor U14521 (N_14521,N_14226,N_14259);
or U14522 (N_14522,N_14259,N_14245);
nor U14523 (N_14523,N_14341,N_14336);
or U14524 (N_14524,N_14232,N_14382);
xnor U14525 (N_14525,N_14251,N_14333);
xnor U14526 (N_14526,N_14397,N_14382);
nor U14527 (N_14527,N_14275,N_14301);
nor U14528 (N_14528,N_14278,N_14282);
xor U14529 (N_14529,N_14341,N_14284);
nor U14530 (N_14530,N_14385,N_14257);
xnor U14531 (N_14531,N_14296,N_14203);
nor U14532 (N_14532,N_14208,N_14395);
nand U14533 (N_14533,N_14307,N_14281);
or U14534 (N_14534,N_14310,N_14225);
xor U14535 (N_14535,N_14340,N_14302);
or U14536 (N_14536,N_14372,N_14204);
xor U14537 (N_14537,N_14302,N_14347);
and U14538 (N_14538,N_14236,N_14260);
or U14539 (N_14539,N_14367,N_14239);
xor U14540 (N_14540,N_14289,N_14374);
and U14541 (N_14541,N_14274,N_14281);
and U14542 (N_14542,N_14300,N_14267);
and U14543 (N_14543,N_14362,N_14386);
xor U14544 (N_14544,N_14372,N_14295);
and U14545 (N_14545,N_14206,N_14278);
nand U14546 (N_14546,N_14298,N_14268);
nand U14547 (N_14547,N_14314,N_14210);
xnor U14548 (N_14548,N_14358,N_14340);
nor U14549 (N_14549,N_14279,N_14361);
nor U14550 (N_14550,N_14388,N_14246);
nor U14551 (N_14551,N_14340,N_14319);
nor U14552 (N_14552,N_14362,N_14233);
or U14553 (N_14553,N_14222,N_14364);
and U14554 (N_14554,N_14313,N_14357);
and U14555 (N_14555,N_14363,N_14356);
nor U14556 (N_14556,N_14204,N_14373);
xor U14557 (N_14557,N_14299,N_14216);
and U14558 (N_14558,N_14343,N_14341);
xnor U14559 (N_14559,N_14227,N_14383);
xnor U14560 (N_14560,N_14330,N_14294);
xnor U14561 (N_14561,N_14369,N_14206);
nand U14562 (N_14562,N_14307,N_14207);
xnor U14563 (N_14563,N_14297,N_14261);
and U14564 (N_14564,N_14312,N_14359);
or U14565 (N_14565,N_14375,N_14307);
nand U14566 (N_14566,N_14320,N_14207);
and U14567 (N_14567,N_14281,N_14280);
nor U14568 (N_14568,N_14265,N_14201);
nor U14569 (N_14569,N_14234,N_14394);
or U14570 (N_14570,N_14301,N_14230);
xnor U14571 (N_14571,N_14262,N_14355);
nor U14572 (N_14572,N_14294,N_14242);
nor U14573 (N_14573,N_14251,N_14397);
xor U14574 (N_14574,N_14254,N_14238);
and U14575 (N_14575,N_14251,N_14394);
and U14576 (N_14576,N_14231,N_14291);
and U14577 (N_14577,N_14275,N_14382);
xor U14578 (N_14578,N_14263,N_14232);
nor U14579 (N_14579,N_14347,N_14210);
nand U14580 (N_14580,N_14201,N_14363);
or U14581 (N_14581,N_14205,N_14214);
or U14582 (N_14582,N_14232,N_14372);
nand U14583 (N_14583,N_14368,N_14222);
or U14584 (N_14584,N_14347,N_14357);
nor U14585 (N_14585,N_14318,N_14281);
nand U14586 (N_14586,N_14307,N_14212);
or U14587 (N_14587,N_14324,N_14248);
or U14588 (N_14588,N_14306,N_14260);
or U14589 (N_14589,N_14368,N_14345);
and U14590 (N_14590,N_14242,N_14335);
nand U14591 (N_14591,N_14209,N_14230);
nor U14592 (N_14592,N_14205,N_14375);
xor U14593 (N_14593,N_14204,N_14399);
xor U14594 (N_14594,N_14316,N_14256);
nor U14595 (N_14595,N_14306,N_14302);
nand U14596 (N_14596,N_14221,N_14283);
nand U14597 (N_14597,N_14373,N_14291);
nand U14598 (N_14598,N_14234,N_14255);
nand U14599 (N_14599,N_14366,N_14319);
or U14600 (N_14600,N_14433,N_14485);
xnor U14601 (N_14601,N_14528,N_14505);
nor U14602 (N_14602,N_14561,N_14453);
xnor U14603 (N_14603,N_14513,N_14437);
nand U14604 (N_14604,N_14546,N_14571);
nand U14605 (N_14605,N_14471,N_14401);
nor U14606 (N_14606,N_14483,N_14515);
xor U14607 (N_14607,N_14527,N_14415);
or U14608 (N_14608,N_14411,N_14523);
or U14609 (N_14609,N_14574,N_14590);
xor U14610 (N_14610,N_14412,N_14583);
or U14611 (N_14611,N_14495,N_14491);
nand U14612 (N_14612,N_14566,N_14425);
and U14613 (N_14613,N_14484,N_14497);
xnor U14614 (N_14614,N_14479,N_14441);
or U14615 (N_14615,N_14499,N_14461);
or U14616 (N_14616,N_14598,N_14439);
nand U14617 (N_14617,N_14444,N_14406);
nand U14618 (N_14618,N_14562,N_14500);
nand U14619 (N_14619,N_14510,N_14476);
or U14620 (N_14620,N_14543,N_14522);
or U14621 (N_14621,N_14596,N_14554);
nand U14622 (N_14622,N_14516,N_14558);
xor U14623 (N_14623,N_14477,N_14587);
and U14624 (N_14624,N_14487,N_14502);
nor U14625 (N_14625,N_14424,N_14430);
nor U14626 (N_14626,N_14573,N_14560);
and U14627 (N_14627,N_14525,N_14409);
and U14628 (N_14628,N_14580,N_14595);
xnor U14629 (N_14629,N_14427,N_14530);
nand U14630 (N_14630,N_14504,N_14532);
or U14631 (N_14631,N_14593,N_14576);
xnor U14632 (N_14632,N_14570,N_14478);
nand U14633 (N_14633,N_14402,N_14416);
xnor U14634 (N_14634,N_14531,N_14462);
nand U14635 (N_14635,N_14470,N_14592);
nor U14636 (N_14636,N_14534,N_14553);
and U14637 (N_14637,N_14454,N_14432);
xor U14638 (N_14638,N_14434,N_14493);
or U14639 (N_14639,N_14535,N_14448);
nand U14640 (N_14640,N_14506,N_14517);
nand U14641 (N_14641,N_14465,N_14551);
or U14642 (N_14642,N_14422,N_14468);
or U14643 (N_14643,N_14450,N_14557);
nand U14644 (N_14644,N_14539,N_14521);
nand U14645 (N_14645,N_14526,N_14435);
nand U14646 (N_14646,N_14445,N_14418);
xor U14647 (N_14647,N_14466,N_14508);
nor U14648 (N_14648,N_14537,N_14542);
nand U14649 (N_14649,N_14579,N_14536);
or U14650 (N_14650,N_14544,N_14581);
nand U14651 (N_14651,N_14519,N_14586);
xor U14652 (N_14652,N_14423,N_14452);
or U14653 (N_14653,N_14456,N_14559);
and U14654 (N_14654,N_14458,N_14467);
xnor U14655 (N_14655,N_14463,N_14589);
and U14656 (N_14656,N_14563,N_14572);
xor U14657 (N_14657,N_14496,N_14457);
or U14658 (N_14658,N_14529,N_14431);
nand U14659 (N_14659,N_14541,N_14509);
or U14660 (N_14660,N_14520,N_14464);
or U14661 (N_14661,N_14414,N_14408);
nor U14662 (N_14662,N_14400,N_14577);
nor U14663 (N_14663,N_14486,N_14555);
nand U14664 (N_14664,N_14417,N_14489);
and U14665 (N_14665,N_14507,N_14429);
nand U14666 (N_14666,N_14455,N_14449);
nor U14667 (N_14667,N_14443,N_14419);
nand U14668 (N_14668,N_14421,N_14472);
nand U14669 (N_14669,N_14550,N_14498);
nor U14670 (N_14670,N_14503,N_14459);
or U14671 (N_14671,N_14492,N_14490);
and U14672 (N_14672,N_14488,N_14407);
and U14673 (N_14673,N_14568,N_14569);
nand U14674 (N_14674,N_14547,N_14545);
nand U14675 (N_14675,N_14548,N_14480);
and U14676 (N_14676,N_14460,N_14575);
xnor U14677 (N_14677,N_14451,N_14440);
xor U14678 (N_14678,N_14428,N_14420);
nor U14679 (N_14679,N_14533,N_14549);
nand U14680 (N_14680,N_14501,N_14594);
or U14681 (N_14681,N_14514,N_14404);
nor U14682 (N_14682,N_14538,N_14403);
xnor U14683 (N_14683,N_14556,N_14481);
or U14684 (N_14684,N_14426,N_14540);
nor U14685 (N_14685,N_14469,N_14591);
nor U14686 (N_14686,N_14564,N_14410);
nor U14687 (N_14687,N_14446,N_14552);
and U14688 (N_14688,N_14578,N_14405);
nand U14689 (N_14689,N_14582,N_14567);
nand U14690 (N_14690,N_14512,N_14442);
or U14691 (N_14691,N_14524,N_14413);
nand U14692 (N_14692,N_14585,N_14511);
or U14693 (N_14693,N_14588,N_14518);
and U14694 (N_14694,N_14494,N_14584);
xnor U14695 (N_14695,N_14565,N_14597);
nand U14696 (N_14696,N_14447,N_14473);
and U14697 (N_14697,N_14599,N_14436);
nor U14698 (N_14698,N_14482,N_14438);
xnor U14699 (N_14699,N_14474,N_14475);
xor U14700 (N_14700,N_14474,N_14591);
or U14701 (N_14701,N_14592,N_14541);
nand U14702 (N_14702,N_14447,N_14584);
nand U14703 (N_14703,N_14578,N_14402);
or U14704 (N_14704,N_14581,N_14576);
xnor U14705 (N_14705,N_14450,N_14526);
nand U14706 (N_14706,N_14498,N_14589);
nor U14707 (N_14707,N_14455,N_14485);
nand U14708 (N_14708,N_14491,N_14594);
xnor U14709 (N_14709,N_14410,N_14561);
xnor U14710 (N_14710,N_14496,N_14435);
nor U14711 (N_14711,N_14432,N_14496);
nor U14712 (N_14712,N_14409,N_14422);
nor U14713 (N_14713,N_14515,N_14552);
xnor U14714 (N_14714,N_14475,N_14530);
nand U14715 (N_14715,N_14525,N_14551);
and U14716 (N_14716,N_14569,N_14431);
or U14717 (N_14717,N_14559,N_14449);
nand U14718 (N_14718,N_14550,N_14515);
nand U14719 (N_14719,N_14417,N_14533);
and U14720 (N_14720,N_14412,N_14478);
and U14721 (N_14721,N_14560,N_14487);
and U14722 (N_14722,N_14448,N_14451);
nor U14723 (N_14723,N_14596,N_14495);
or U14724 (N_14724,N_14524,N_14560);
or U14725 (N_14725,N_14575,N_14462);
nor U14726 (N_14726,N_14485,N_14419);
nand U14727 (N_14727,N_14576,N_14455);
and U14728 (N_14728,N_14442,N_14595);
and U14729 (N_14729,N_14577,N_14503);
or U14730 (N_14730,N_14405,N_14563);
nor U14731 (N_14731,N_14503,N_14573);
nand U14732 (N_14732,N_14561,N_14509);
nor U14733 (N_14733,N_14417,N_14488);
nand U14734 (N_14734,N_14447,N_14598);
nand U14735 (N_14735,N_14534,N_14479);
nor U14736 (N_14736,N_14539,N_14404);
nand U14737 (N_14737,N_14457,N_14476);
nand U14738 (N_14738,N_14402,N_14484);
or U14739 (N_14739,N_14595,N_14517);
xnor U14740 (N_14740,N_14462,N_14583);
or U14741 (N_14741,N_14461,N_14429);
xnor U14742 (N_14742,N_14574,N_14579);
or U14743 (N_14743,N_14583,N_14499);
and U14744 (N_14744,N_14405,N_14417);
or U14745 (N_14745,N_14597,N_14547);
and U14746 (N_14746,N_14516,N_14513);
nor U14747 (N_14747,N_14575,N_14465);
nor U14748 (N_14748,N_14459,N_14479);
and U14749 (N_14749,N_14424,N_14488);
and U14750 (N_14750,N_14473,N_14518);
nor U14751 (N_14751,N_14595,N_14570);
nand U14752 (N_14752,N_14503,N_14487);
and U14753 (N_14753,N_14484,N_14524);
xnor U14754 (N_14754,N_14518,N_14500);
xnor U14755 (N_14755,N_14542,N_14479);
xnor U14756 (N_14756,N_14479,N_14466);
xor U14757 (N_14757,N_14582,N_14590);
nand U14758 (N_14758,N_14418,N_14502);
nor U14759 (N_14759,N_14540,N_14457);
nor U14760 (N_14760,N_14467,N_14575);
nor U14761 (N_14761,N_14573,N_14461);
nor U14762 (N_14762,N_14564,N_14503);
and U14763 (N_14763,N_14403,N_14517);
nand U14764 (N_14764,N_14543,N_14593);
nor U14765 (N_14765,N_14504,N_14516);
nand U14766 (N_14766,N_14518,N_14522);
xor U14767 (N_14767,N_14434,N_14484);
nor U14768 (N_14768,N_14519,N_14578);
nor U14769 (N_14769,N_14462,N_14436);
and U14770 (N_14770,N_14473,N_14568);
nor U14771 (N_14771,N_14419,N_14407);
nand U14772 (N_14772,N_14470,N_14496);
or U14773 (N_14773,N_14571,N_14489);
xnor U14774 (N_14774,N_14566,N_14501);
xnor U14775 (N_14775,N_14510,N_14594);
nor U14776 (N_14776,N_14491,N_14528);
nand U14777 (N_14777,N_14464,N_14413);
or U14778 (N_14778,N_14405,N_14471);
nor U14779 (N_14779,N_14481,N_14577);
nor U14780 (N_14780,N_14444,N_14587);
nor U14781 (N_14781,N_14528,N_14468);
nor U14782 (N_14782,N_14486,N_14495);
nand U14783 (N_14783,N_14466,N_14435);
nor U14784 (N_14784,N_14529,N_14563);
and U14785 (N_14785,N_14519,N_14580);
or U14786 (N_14786,N_14571,N_14493);
or U14787 (N_14787,N_14422,N_14406);
nand U14788 (N_14788,N_14402,N_14507);
and U14789 (N_14789,N_14531,N_14519);
xnor U14790 (N_14790,N_14589,N_14427);
or U14791 (N_14791,N_14490,N_14439);
and U14792 (N_14792,N_14512,N_14538);
and U14793 (N_14793,N_14556,N_14484);
nor U14794 (N_14794,N_14586,N_14531);
or U14795 (N_14795,N_14445,N_14524);
nor U14796 (N_14796,N_14481,N_14584);
nor U14797 (N_14797,N_14561,N_14514);
xor U14798 (N_14798,N_14574,N_14561);
and U14799 (N_14799,N_14579,N_14549);
nand U14800 (N_14800,N_14737,N_14685);
or U14801 (N_14801,N_14771,N_14778);
xor U14802 (N_14802,N_14707,N_14687);
xor U14803 (N_14803,N_14752,N_14795);
or U14804 (N_14804,N_14789,N_14772);
nor U14805 (N_14805,N_14726,N_14730);
xnor U14806 (N_14806,N_14723,N_14613);
xnor U14807 (N_14807,N_14641,N_14649);
or U14808 (N_14808,N_14756,N_14762);
and U14809 (N_14809,N_14692,N_14798);
or U14810 (N_14810,N_14635,N_14663);
and U14811 (N_14811,N_14677,N_14769);
and U14812 (N_14812,N_14767,N_14793);
or U14813 (N_14813,N_14765,N_14655);
or U14814 (N_14814,N_14788,N_14693);
nand U14815 (N_14815,N_14624,N_14782);
nor U14816 (N_14816,N_14748,N_14619);
or U14817 (N_14817,N_14700,N_14689);
nor U14818 (N_14818,N_14733,N_14740);
nand U14819 (N_14819,N_14751,N_14761);
and U14820 (N_14820,N_14732,N_14658);
and U14821 (N_14821,N_14754,N_14775);
and U14822 (N_14822,N_14786,N_14713);
nand U14823 (N_14823,N_14695,N_14736);
xor U14824 (N_14824,N_14637,N_14631);
nand U14825 (N_14825,N_14717,N_14675);
nor U14826 (N_14826,N_14640,N_14626);
nor U14827 (N_14827,N_14780,N_14605);
nand U14828 (N_14828,N_14682,N_14719);
xor U14829 (N_14829,N_14758,N_14671);
xor U14830 (N_14830,N_14623,N_14622);
nand U14831 (N_14831,N_14670,N_14665);
or U14832 (N_14832,N_14743,N_14648);
nor U14833 (N_14833,N_14790,N_14755);
nor U14834 (N_14834,N_14629,N_14796);
xor U14835 (N_14835,N_14638,N_14759);
or U14836 (N_14836,N_14760,N_14698);
xnor U14837 (N_14837,N_14628,N_14673);
nor U14838 (N_14838,N_14714,N_14776);
xnor U14839 (N_14839,N_14634,N_14794);
xor U14840 (N_14840,N_14781,N_14630);
nand U14841 (N_14841,N_14712,N_14651);
and U14842 (N_14842,N_14676,N_14787);
nand U14843 (N_14843,N_14618,N_14627);
or U14844 (N_14844,N_14610,N_14791);
nand U14845 (N_14845,N_14686,N_14683);
xor U14846 (N_14846,N_14600,N_14617);
xnor U14847 (N_14847,N_14615,N_14728);
nand U14848 (N_14848,N_14734,N_14702);
nand U14849 (N_14849,N_14753,N_14645);
nand U14850 (N_14850,N_14715,N_14738);
or U14851 (N_14851,N_14768,N_14770);
xnor U14852 (N_14852,N_14666,N_14729);
xor U14853 (N_14853,N_14691,N_14625);
and U14854 (N_14854,N_14757,N_14697);
xor U14855 (N_14855,N_14709,N_14611);
and U14856 (N_14856,N_14703,N_14750);
or U14857 (N_14857,N_14799,N_14764);
nand U14858 (N_14858,N_14797,N_14746);
xor U14859 (N_14859,N_14735,N_14642);
nor U14860 (N_14860,N_14609,N_14745);
nand U14861 (N_14861,N_14603,N_14679);
or U14862 (N_14862,N_14783,N_14701);
nor U14863 (N_14863,N_14784,N_14654);
or U14864 (N_14864,N_14664,N_14653);
nand U14865 (N_14865,N_14668,N_14711);
nor U14866 (N_14866,N_14646,N_14774);
xnor U14867 (N_14867,N_14644,N_14601);
or U14868 (N_14868,N_14727,N_14620);
or U14869 (N_14869,N_14792,N_14747);
xor U14870 (N_14870,N_14680,N_14696);
nor U14871 (N_14871,N_14636,N_14633);
nor U14872 (N_14872,N_14694,N_14725);
or U14873 (N_14873,N_14699,N_14766);
or U14874 (N_14874,N_14744,N_14721);
or U14875 (N_14875,N_14785,N_14674);
or U14876 (N_14876,N_14705,N_14614);
xnor U14877 (N_14877,N_14662,N_14643);
xnor U14878 (N_14878,N_14716,N_14657);
and U14879 (N_14879,N_14612,N_14604);
nor U14880 (N_14880,N_14739,N_14602);
or U14881 (N_14881,N_14706,N_14621);
nor U14882 (N_14882,N_14741,N_14656);
nand U14883 (N_14883,N_14777,N_14684);
and U14884 (N_14884,N_14678,N_14690);
nand U14885 (N_14885,N_14606,N_14607);
or U14886 (N_14886,N_14632,N_14763);
nor U14887 (N_14887,N_14688,N_14773);
and U14888 (N_14888,N_14704,N_14710);
xnor U14889 (N_14889,N_14661,N_14681);
and U14890 (N_14890,N_14650,N_14749);
or U14891 (N_14891,N_14669,N_14708);
nand U14892 (N_14892,N_14718,N_14647);
nand U14893 (N_14893,N_14639,N_14779);
and U14894 (N_14894,N_14724,N_14616);
nor U14895 (N_14895,N_14652,N_14659);
and U14896 (N_14896,N_14731,N_14742);
xnor U14897 (N_14897,N_14667,N_14672);
or U14898 (N_14898,N_14660,N_14722);
xnor U14899 (N_14899,N_14608,N_14720);
nand U14900 (N_14900,N_14678,N_14617);
xor U14901 (N_14901,N_14717,N_14661);
nor U14902 (N_14902,N_14694,N_14758);
xor U14903 (N_14903,N_14611,N_14616);
xnor U14904 (N_14904,N_14764,N_14672);
and U14905 (N_14905,N_14787,N_14693);
xnor U14906 (N_14906,N_14635,N_14672);
xor U14907 (N_14907,N_14663,N_14692);
xor U14908 (N_14908,N_14606,N_14742);
xor U14909 (N_14909,N_14734,N_14761);
nand U14910 (N_14910,N_14737,N_14762);
xnor U14911 (N_14911,N_14615,N_14661);
nor U14912 (N_14912,N_14773,N_14738);
nor U14913 (N_14913,N_14790,N_14608);
nand U14914 (N_14914,N_14615,N_14775);
xor U14915 (N_14915,N_14621,N_14705);
nand U14916 (N_14916,N_14769,N_14742);
and U14917 (N_14917,N_14730,N_14663);
nor U14918 (N_14918,N_14634,N_14605);
nor U14919 (N_14919,N_14757,N_14794);
nand U14920 (N_14920,N_14604,N_14762);
or U14921 (N_14921,N_14693,N_14735);
or U14922 (N_14922,N_14655,N_14605);
nor U14923 (N_14923,N_14789,N_14703);
nor U14924 (N_14924,N_14718,N_14772);
and U14925 (N_14925,N_14659,N_14603);
and U14926 (N_14926,N_14752,N_14768);
nor U14927 (N_14927,N_14743,N_14727);
xor U14928 (N_14928,N_14706,N_14664);
xor U14929 (N_14929,N_14649,N_14792);
xor U14930 (N_14930,N_14665,N_14675);
xor U14931 (N_14931,N_14766,N_14658);
nor U14932 (N_14932,N_14615,N_14749);
xor U14933 (N_14933,N_14794,N_14605);
nand U14934 (N_14934,N_14685,N_14794);
nand U14935 (N_14935,N_14611,N_14694);
nand U14936 (N_14936,N_14645,N_14626);
or U14937 (N_14937,N_14719,N_14691);
and U14938 (N_14938,N_14682,N_14699);
xnor U14939 (N_14939,N_14602,N_14717);
xor U14940 (N_14940,N_14755,N_14752);
nor U14941 (N_14941,N_14659,N_14729);
nor U14942 (N_14942,N_14680,N_14752);
and U14943 (N_14943,N_14780,N_14772);
xnor U14944 (N_14944,N_14624,N_14668);
and U14945 (N_14945,N_14708,N_14726);
or U14946 (N_14946,N_14689,N_14653);
and U14947 (N_14947,N_14685,N_14647);
or U14948 (N_14948,N_14761,N_14721);
or U14949 (N_14949,N_14725,N_14711);
or U14950 (N_14950,N_14682,N_14689);
nand U14951 (N_14951,N_14600,N_14723);
and U14952 (N_14952,N_14746,N_14655);
and U14953 (N_14953,N_14782,N_14774);
nor U14954 (N_14954,N_14716,N_14663);
and U14955 (N_14955,N_14706,N_14730);
and U14956 (N_14956,N_14657,N_14769);
nor U14957 (N_14957,N_14724,N_14646);
xnor U14958 (N_14958,N_14719,N_14684);
nand U14959 (N_14959,N_14732,N_14775);
nand U14960 (N_14960,N_14698,N_14726);
nor U14961 (N_14961,N_14644,N_14751);
nand U14962 (N_14962,N_14667,N_14674);
nor U14963 (N_14963,N_14632,N_14620);
and U14964 (N_14964,N_14620,N_14720);
or U14965 (N_14965,N_14667,N_14631);
or U14966 (N_14966,N_14655,N_14619);
nor U14967 (N_14967,N_14798,N_14653);
nor U14968 (N_14968,N_14662,N_14798);
nor U14969 (N_14969,N_14740,N_14729);
xor U14970 (N_14970,N_14752,N_14602);
xor U14971 (N_14971,N_14785,N_14629);
and U14972 (N_14972,N_14645,N_14649);
xnor U14973 (N_14973,N_14633,N_14745);
xor U14974 (N_14974,N_14707,N_14641);
or U14975 (N_14975,N_14711,N_14646);
nand U14976 (N_14976,N_14696,N_14747);
or U14977 (N_14977,N_14785,N_14615);
and U14978 (N_14978,N_14675,N_14763);
nand U14979 (N_14979,N_14755,N_14608);
and U14980 (N_14980,N_14625,N_14717);
or U14981 (N_14981,N_14673,N_14767);
or U14982 (N_14982,N_14702,N_14641);
or U14983 (N_14983,N_14642,N_14611);
nand U14984 (N_14984,N_14654,N_14699);
nand U14985 (N_14985,N_14766,N_14799);
nand U14986 (N_14986,N_14753,N_14668);
and U14987 (N_14987,N_14752,N_14709);
and U14988 (N_14988,N_14617,N_14615);
nand U14989 (N_14989,N_14744,N_14733);
nor U14990 (N_14990,N_14777,N_14754);
nor U14991 (N_14991,N_14635,N_14634);
and U14992 (N_14992,N_14732,N_14667);
nand U14993 (N_14993,N_14606,N_14617);
nor U14994 (N_14994,N_14735,N_14730);
nor U14995 (N_14995,N_14751,N_14750);
nor U14996 (N_14996,N_14604,N_14640);
nor U14997 (N_14997,N_14776,N_14752);
nor U14998 (N_14998,N_14616,N_14600);
or U14999 (N_14999,N_14789,N_14701);
nand UO_0 (O_0,N_14910,N_14930);
nor UO_1 (O_1,N_14827,N_14839);
nand UO_2 (O_2,N_14819,N_14817);
and UO_3 (O_3,N_14886,N_14836);
nand UO_4 (O_4,N_14983,N_14824);
nor UO_5 (O_5,N_14865,N_14904);
nand UO_6 (O_6,N_14866,N_14869);
and UO_7 (O_7,N_14849,N_14897);
xnor UO_8 (O_8,N_14860,N_14960);
or UO_9 (O_9,N_14932,N_14846);
xor UO_10 (O_10,N_14894,N_14812);
and UO_11 (O_11,N_14864,N_14959);
and UO_12 (O_12,N_14908,N_14898);
nand UO_13 (O_13,N_14835,N_14803);
xor UO_14 (O_14,N_14945,N_14918);
nor UO_15 (O_15,N_14831,N_14950);
nor UO_16 (O_16,N_14858,N_14970);
nand UO_17 (O_17,N_14820,N_14913);
xor UO_18 (O_18,N_14916,N_14911);
xnor UO_19 (O_19,N_14991,N_14892);
and UO_20 (O_20,N_14906,N_14879);
or UO_21 (O_21,N_14999,N_14828);
nor UO_22 (O_22,N_14901,N_14893);
xor UO_23 (O_23,N_14997,N_14889);
xnor UO_24 (O_24,N_14914,N_14810);
nor UO_25 (O_25,N_14905,N_14829);
xor UO_26 (O_26,N_14938,N_14811);
nand UO_27 (O_27,N_14826,N_14925);
nand UO_28 (O_28,N_14816,N_14888);
nand UO_29 (O_29,N_14882,N_14856);
nand UO_30 (O_30,N_14834,N_14937);
nor UO_31 (O_31,N_14854,N_14963);
and UO_32 (O_32,N_14994,N_14955);
nor UO_33 (O_33,N_14890,N_14808);
xnor UO_34 (O_34,N_14915,N_14952);
nand UO_35 (O_35,N_14832,N_14992);
or UO_36 (O_36,N_14953,N_14806);
and UO_37 (O_37,N_14948,N_14917);
nor UO_38 (O_38,N_14941,N_14919);
or UO_39 (O_39,N_14976,N_14927);
and UO_40 (O_40,N_14958,N_14800);
or UO_41 (O_41,N_14875,N_14968);
nand UO_42 (O_42,N_14821,N_14802);
and UO_43 (O_43,N_14857,N_14928);
nand UO_44 (O_44,N_14880,N_14801);
xnor UO_45 (O_45,N_14934,N_14982);
nand UO_46 (O_46,N_14840,N_14986);
nor UO_47 (O_47,N_14838,N_14896);
nor UO_48 (O_48,N_14951,N_14837);
nand UO_49 (O_49,N_14907,N_14987);
nor UO_50 (O_50,N_14845,N_14964);
nand UO_51 (O_51,N_14926,N_14990);
nand UO_52 (O_52,N_14962,N_14931);
nand UO_53 (O_53,N_14965,N_14853);
or UO_54 (O_54,N_14924,N_14844);
xnor UO_55 (O_55,N_14949,N_14985);
nor UO_56 (O_56,N_14935,N_14872);
and UO_57 (O_57,N_14996,N_14979);
and UO_58 (O_58,N_14807,N_14900);
xnor UO_59 (O_59,N_14881,N_14943);
nor UO_60 (O_60,N_14862,N_14946);
and UO_61 (O_61,N_14944,N_14841);
or UO_62 (O_62,N_14850,N_14984);
or UO_63 (O_63,N_14877,N_14973);
xor UO_64 (O_64,N_14902,N_14921);
nor UO_65 (O_65,N_14922,N_14874);
xnor UO_66 (O_66,N_14929,N_14891);
and UO_67 (O_67,N_14966,N_14895);
and UO_68 (O_68,N_14939,N_14995);
nand UO_69 (O_69,N_14912,N_14868);
nand UO_70 (O_70,N_14967,N_14822);
nand UO_71 (O_71,N_14814,N_14855);
and UO_72 (O_72,N_14847,N_14947);
or UO_73 (O_73,N_14936,N_14848);
or UO_74 (O_74,N_14954,N_14873);
and UO_75 (O_75,N_14956,N_14833);
and UO_76 (O_76,N_14842,N_14989);
xnor UO_77 (O_77,N_14978,N_14899);
nor UO_78 (O_78,N_14867,N_14969);
xor UO_79 (O_79,N_14813,N_14818);
nand UO_80 (O_80,N_14843,N_14870);
or UO_81 (O_81,N_14971,N_14815);
or UO_82 (O_82,N_14961,N_14923);
xnor UO_83 (O_83,N_14993,N_14975);
or UO_84 (O_84,N_14980,N_14885);
and UO_85 (O_85,N_14977,N_14940);
or UO_86 (O_86,N_14852,N_14861);
and UO_87 (O_87,N_14859,N_14957);
or UO_88 (O_88,N_14851,N_14876);
nor UO_89 (O_89,N_14974,N_14909);
and UO_90 (O_90,N_14805,N_14998);
nor UO_91 (O_91,N_14804,N_14942);
nand UO_92 (O_92,N_14809,N_14883);
nand UO_93 (O_93,N_14863,N_14933);
nor UO_94 (O_94,N_14887,N_14988);
nand UO_95 (O_95,N_14871,N_14825);
xor UO_96 (O_96,N_14823,N_14878);
nor UO_97 (O_97,N_14903,N_14981);
or UO_98 (O_98,N_14972,N_14884);
nand UO_99 (O_99,N_14920,N_14830);
xor UO_100 (O_100,N_14802,N_14939);
nand UO_101 (O_101,N_14957,N_14892);
nor UO_102 (O_102,N_14971,N_14869);
or UO_103 (O_103,N_14887,N_14909);
nand UO_104 (O_104,N_14965,N_14865);
and UO_105 (O_105,N_14800,N_14829);
xnor UO_106 (O_106,N_14879,N_14996);
and UO_107 (O_107,N_14885,N_14899);
nand UO_108 (O_108,N_14912,N_14827);
and UO_109 (O_109,N_14887,N_14879);
or UO_110 (O_110,N_14881,N_14841);
and UO_111 (O_111,N_14903,N_14839);
nor UO_112 (O_112,N_14988,N_14840);
and UO_113 (O_113,N_14941,N_14824);
and UO_114 (O_114,N_14897,N_14950);
nor UO_115 (O_115,N_14954,N_14971);
nor UO_116 (O_116,N_14834,N_14801);
nand UO_117 (O_117,N_14968,N_14839);
or UO_118 (O_118,N_14810,N_14963);
xor UO_119 (O_119,N_14982,N_14825);
nor UO_120 (O_120,N_14928,N_14830);
nand UO_121 (O_121,N_14905,N_14960);
nor UO_122 (O_122,N_14852,N_14948);
xnor UO_123 (O_123,N_14818,N_14852);
nand UO_124 (O_124,N_14979,N_14956);
and UO_125 (O_125,N_14967,N_14993);
or UO_126 (O_126,N_14972,N_14869);
nor UO_127 (O_127,N_14837,N_14910);
or UO_128 (O_128,N_14818,N_14902);
and UO_129 (O_129,N_14894,N_14912);
nor UO_130 (O_130,N_14823,N_14902);
nand UO_131 (O_131,N_14811,N_14845);
nand UO_132 (O_132,N_14912,N_14859);
or UO_133 (O_133,N_14934,N_14967);
xnor UO_134 (O_134,N_14842,N_14971);
and UO_135 (O_135,N_14928,N_14903);
xnor UO_136 (O_136,N_14977,N_14844);
xnor UO_137 (O_137,N_14976,N_14900);
nor UO_138 (O_138,N_14996,N_14976);
or UO_139 (O_139,N_14935,N_14924);
xnor UO_140 (O_140,N_14831,N_14974);
xor UO_141 (O_141,N_14992,N_14872);
and UO_142 (O_142,N_14825,N_14909);
nand UO_143 (O_143,N_14892,N_14922);
xnor UO_144 (O_144,N_14865,N_14839);
nor UO_145 (O_145,N_14887,N_14889);
xnor UO_146 (O_146,N_14837,N_14998);
or UO_147 (O_147,N_14802,N_14840);
and UO_148 (O_148,N_14994,N_14975);
xor UO_149 (O_149,N_14912,N_14968);
nor UO_150 (O_150,N_14933,N_14807);
or UO_151 (O_151,N_14842,N_14868);
xnor UO_152 (O_152,N_14894,N_14927);
xnor UO_153 (O_153,N_14890,N_14982);
or UO_154 (O_154,N_14882,N_14961);
or UO_155 (O_155,N_14920,N_14897);
nor UO_156 (O_156,N_14848,N_14885);
and UO_157 (O_157,N_14927,N_14928);
and UO_158 (O_158,N_14925,N_14994);
xnor UO_159 (O_159,N_14979,N_14910);
and UO_160 (O_160,N_14993,N_14977);
nor UO_161 (O_161,N_14813,N_14987);
nor UO_162 (O_162,N_14977,N_14806);
nor UO_163 (O_163,N_14903,N_14812);
nand UO_164 (O_164,N_14910,N_14882);
and UO_165 (O_165,N_14864,N_14926);
nand UO_166 (O_166,N_14884,N_14837);
or UO_167 (O_167,N_14919,N_14882);
or UO_168 (O_168,N_14819,N_14970);
and UO_169 (O_169,N_14932,N_14892);
xnor UO_170 (O_170,N_14918,N_14844);
xor UO_171 (O_171,N_14997,N_14985);
and UO_172 (O_172,N_14823,N_14849);
and UO_173 (O_173,N_14807,N_14988);
and UO_174 (O_174,N_14818,N_14890);
nor UO_175 (O_175,N_14988,N_14928);
and UO_176 (O_176,N_14809,N_14942);
nand UO_177 (O_177,N_14908,N_14998);
xor UO_178 (O_178,N_14983,N_14839);
nand UO_179 (O_179,N_14952,N_14867);
and UO_180 (O_180,N_14916,N_14932);
nor UO_181 (O_181,N_14960,N_14820);
nand UO_182 (O_182,N_14816,N_14957);
nor UO_183 (O_183,N_14978,N_14910);
nand UO_184 (O_184,N_14936,N_14866);
xor UO_185 (O_185,N_14914,N_14994);
nand UO_186 (O_186,N_14908,N_14991);
and UO_187 (O_187,N_14886,N_14899);
nand UO_188 (O_188,N_14956,N_14968);
xor UO_189 (O_189,N_14996,N_14844);
xnor UO_190 (O_190,N_14959,N_14992);
xnor UO_191 (O_191,N_14972,N_14845);
and UO_192 (O_192,N_14974,N_14860);
and UO_193 (O_193,N_14977,N_14963);
and UO_194 (O_194,N_14882,N_14849);
nor UO_195 (O_195,N_14820,N_14877);
nor UO_196 (O_196,N_14834,N_14869);
xor UO_197 (O_197,N_14814,N_14905);
and UO_198 (O_198,N_14824,N_14947);
nand UO_199 (O_199,N_14906,N_14841);
or UO_200 (O_200,N_14893,N_14843);
and UO_201 (O_201,N_14944,N_14939);
and UO_202 (O_202,N_14882,N_14869);
nand UO_203 (O_203,N_14917,N_14998);
or UO_204 (O_204,N_14995,N_14929);
nand UO_205 (O_205,N_14861,N_14986);
or UO_206 (O_206,N_14917,N_14972);
xor UO_207 (O_207,N_14800,N_14821);
nor UO_208 (O_208,N_14908,N_14826);
nor UO_209 (O_209,N_14891,N_14997);
nor UO_210 (O_210,N_14806,N_14881);
xnor UO_211 (O_211,N_14864,N_14977);
nor UO_212 (O_212,N_14841,N_14928);
or UO_213 (O_213,N_14960,N_14990);
or UO_214 (O_214,N_14841,N_14978);
nand UO_215 (O_215,N_14992,N_14914);
xnor UO_216 (O_216,N_14983,N_14978);
and UO_217 (O_217,N_14958,N_14862);
xnor UO_218 (O_218,N_14888,N_14896);
or UO_219 (O_219,N_14851,N_14945);
xnor UO_220 (O_220,N_14833,N_14981);
and UO_221 (O_221,N_14845,N_14812);
xnor UO_222 (O_222,N_14800,N_14910);
nor UO_223 (O_223,N_14936,N_14940);
xnor UO_224 (O_224,N_14817,N_14940);
nor UO_225 (O_225,N_14829,N_14907);
xor UO_226 (O_226,N_14969,N_14881);
and UO_227 (O_227,N_14895,N_14943);
nand UO_228 (O_228,N_14843,N_14966);
and UO_229 (O_229,N_14990,N_14934);
or UO_230 (O_230,N_14829,N_14854);
or UO_231 (O_231,N_14804,N_14847);
nand UO_232 (O_232,N_14885,N_14934);
xnor UO_233 (O_233,N_14968,N_14892);
nand UO_234 (O_234,N_14974,N_14847);
xnor UO_235 (O_235,N_14991,N_14918);
nand UO_236 (O_236,N_14842,N_14970);
or UO_237 (O_237,N_14820,N_14867);
nor UO_238 (O_238,N_14975,N_14806);
and UO_239 (O_239,N_14876,N_14832);
or UO_240 (O_240,N_14856,N_14808);
nor UO_241 (O_241,N_14973,N_14863);
and UO_242 (O_242,N_14891,N_14961);
nand UO_243 (O_243,N_14909,N_14970);
or UO_244 (O_244,N_14910,N_14852);
nor UO_245 (O_245,N_14837,N_14926);
xor UO_246 (O_246,N_14885,N_14861);
or UO_247 (O_247,N_14984,N_14803);
and UO_248 (O_248,N_14819,N_14975);
nor UO_249 (O_249,N_14994,N_14980);
nand UO_250 (O_250,N_14885,N_14828);
nand UO_251 (O_251,N_14953,N_14934);
xor UO_252 (O_252,N_14803,N_14944);
nor UO_253 (O_253,N_14805,N_14824);
nand UO_254 (O_254,N_14861,N_14997);
nor UO_255 (O_255,N_14968,N_14896);
nor UO_256 (O_256,N_14974,N_14940);
and UO_257 (O_257,N_14988,N_14885);
xor UO_258 (O_258,N_14839,N_14915);
and UO_259 (O_259,N_14847,N_14988);
and UO_260 (O_260,N_14958,N_14823);
xnor UO_261 (O_261,N_14971,N_14966);
nand UO_262 (O_262,N_14909,N_14947);
or UO_263 (O_263,N_14939,N_14977);
or UO_264 (O_264,N_14917,N_14982);
and UO_265 (O_265,N_14897,N_14993);
nand UO_266 (O_266,N_14880,N_14850);
nand UO_267 (O_267,N_14977,N_14829);
xnor UO_268 (O_268,N_14887,N_14985);
or UO_269 (O_269,N_14921,N_14896);
nor UO_270 (O_270,N_14992,N_14895);
xor UO_271 (O_271,N_14829,N_14970);
xnor UO_272 (O_272,N_14947,N_14901);
nand UO_273 (O_273,N_14999,N_14817);
xnor UO_274 (O_274,N_14883,N_14829);
nor UO_275 (O_275,N_14973,N_14883);
and UO_276 (O_276,N_14831,N_14844);
nand UO_277 (O_277,N_14879,N_14907);
xnor UO_278 (O_278,N_14949,N_14921);
xnor UO_279 (O_279,N_14922,N_14859);
xnor UO_280 (O_280,N_14950,N_14953);
and UO_281 (O_281,N_14878,N_14922);
and UO_282 (O_282,N_14950,N_14810);
nor UO_283 (O_283,N_14917,N_14971);
xnor UO_284 (O_284,N_14916,N_14966);
or UO_285 (O_285,N_14893,N_14933);
or UO_286 (O_286,N_14960,N_14826);
xor UO_287 (O_287,N_14945,N_14943);
nand UO_288 (O_288,N_14955,N_14841);
nand UO_289 (O_289,N_14885,N_14879);
nand UO_290 (O_290,N_14887,N_14977);
nor UO_291 (O_291,N_14887,N_14883);
xor UO_292 (O_292,N_14834,N_14974);
xor UO_293 (O_293,N_14938,N_14989);
nor UO_294 (O_294,N_14847,N_14894);
and UO_295 (O_295,N_14959,N_14941);
nor UO_296 (O_296,N_14987,N_14982);
xor UO_297 (O_297,N_14978,N_14839);
or UO_298 (O_298,N_14876,N_14999);
nor UO_299 (O_299,N_14957,N_14875);
and UO_300 (O_300,N_14835,N_14890);
and UO_301 (O_301,N_14866,N_14933);
or UO_302 (O_302,N_14848,N_14938);
nor UO_303 (O_303,N_14984,N_14939);
nor UO_304 (O_304,N_14920,N_14982);
nand UO_305 (O_305,N_14808,N_14914);
nor UO_306 (O_306,N_14995,N_14801);
nand UO_307 (O_307,N_14982,N_14966);
and UO_308 (O_308,N_14834,N_14807);
nor UO_309 (O_309,N_14859,N_14960);
and UO_310 (O_310,N_14938,N_14969);
nor UO_311 (O_311,N_14984,N_14988);
and UO_312 (O_312,N_14943,N_14927);
or UO_313 (O_313,N_14919,N_14964);
nand UO_314 (O_314,N_14905,N_14835);
and UO_315 (O_315,N_14838,N_14992);
nor UO_316 (O_316,N_14996,N_14823);
xnor UO_317 (O_317,N_14923,N_14894);
xnor UO_318 (O_318,N_14978,N_14840);
nand UO_319 (O_319,N_14830,N_14855);
nand UO_320 (O_320,N_14811,N_14805);
and UO_321 (O_321,N_14967,N_14825);
nand UO_322 (O_322,N_14874,N_14928);
nor UO_323 (O_323,N_14826,N_14933);
nor UO_324 (O_324,N_14976,N_14809);
nor UO_325 (O_325,N_14827,N_14877);
nor UO_326 (O_326,N_14887,N_14933);
and UO_327 (O_327,N_14870,N_14982);
and UO_328 (O_328,N_14958,N_14967);
or UO_329 (O_329,N_14823,N_14992);
xnor UO_330 (O_330,N_14987,N_14927);
nor UO_331 (O_331,N_14864,N_14933);
nor UO_332 (O_332,N_14814,N_14903);
nand UO_333 (O_333,N_14999,N_14863);
nor UO_334 (O_334,N_14844,N_14809);
xor UO_335 (O_335,N_14807,N_14920);
or UO_336 (O_336,N_14870,N_14929);
or UO_337 (O_337,N_14959,N_14889);
and UO_338 (O_338,N_14995,N_14950);
and UO_339 (O_339,N_14834,N_14961);
nor UO_340 (O_340,N_14917,N_14888);
and UO_341 (O_341,N_14948,N_14812);
and UO_342 (O_342,N_14971,N_14947);
and UO_343 (O_343,N_14902,N_14957);
xnor UO_344 (O_344,N_14909,N_14874);
and UO_345 (O_345,N_14840,N_14854);
and UO_346 (O_346,N_14869,N_14900);
and UO_347 (O_347,N_14978,N_14825);
nand UO_348 (O_348,N_14978,N_14897);
and UO_349 (O_349,N_14915,N_14921);
nor UO_350 (O_350,N_14939,N_14947);
or UO_351 (O_351,N_14937,N_14934);
nor UO_352 (O_352,N_14928,N_14858);
or UO_353 (O_353,N_14950,N_14890);
and UO_354 (O_354,N_14900,N_14923);
nand UO_355 (O_355,N_14979,N_14922);
nor UO_356 (O_356,N_14829,N_14817);
nand UO_357 (O_357,N_14969,N_14843);
xnor UO_358 (O_358,N_14986,N_14999);
or UO_359 (O_359,N_14935,N_14966);
and UO_360 (O_360,N_14930,N_14878);
xor UO_361 (O_361,N_14907,N_14848);
nor UO_362 (O_362,N_14827,N_14944);
nand UO_363 (O_363,N_14920,N_14898);
nor UO_364 (O_364,N_14939,N_14836);
xor UO_365 (O_365,N_14997,N_14866);
nand UO_366 (O_366,N_14824,N_14914);
nand UO_367 (O_367,N_14875,N_14857);
or UO_368 (O_368,N_14895,N_14909);
xnor UO_369 (O_369,N_14984,N_14813);
and UO_370 (O_370,N_14950,N_14940);
nand UO_371 (O_371,N_14957,N_14806);
and UO_372 (O_372,N_14880,N_14959);
and UO_373 (O_373,N_14808,N_14828);
nand UO_374 (O_374,N_14821,N_14838);
nand UO_375 (O_375,N_14863,N_14936);
and UO_376 (O_376,N_14819,N_14918);
or UO_377 (O_377,N_14912,N_14945);
or UO_378 (O_378,N_14883,N_14934);
nand UO_379 (O_379,N_14881,N_14964);
xor UO_380 (O_380,N_14927,N_14992);
xnor UO_381 (O_381,N_14976,N_14986);
and UO_382 (O_382,N_14883,N_14879);
and UO_383 (O_383,N_14903,N_14939);
xnor UO_384 (O_384,N_14952,N_14854);
or UO_385 (O_385,N_14936,N_14899);
nor UO_386 (O_386,N_14987,N_14884);
nand UO_387 (O_387,N_14883,N_14820);
and UO_388 (O_388,N_14814,N_14899);
nor UO_389 (O_389,N_14927,N_14999);
and UO_390 (O_390,N_14940,N_14997);
or UO_391 (O_391,N_14962,N_14997);
nor UO_392 (O_392,N_14996,N_14812);
or UO_393 (O_393,N_14870,N_14932);
and UO_394 (O_394,N_14859,N_14969);
xnor UO_395 (O_395,N_14832,N_14838);
or UO_396 (O_396,N_14900,N_14879);
xnor UO_397 (O_397,N_14865,N_14853);
nand UO_398 (O_398,N_14828,N_14803);
nor UO_399 (O_399,N_14943,N_14838);
xor UO_400 (O_400,N_14847,N_14814);
and UO_401 (O_401,N_14910,N_14805);
nand UO_402 (O_402,N_14986,N_14947);
or UO_403 (O_403,N_14927,N_14901);
or UO_404 (O_404,N_14856,N_14825);
nand UO_405 (O_405,N_14960,N_14809);
or UO_406 (O_406,N_14943,N_14869);
and UO_407 (O_407,N_14856,N_14928);
or UO_408 (O_408,N_14970,N_14868);
and UO_409 (O_409,N_14994,N_14942);
and UO_410 (O_410,N_14917,N_14963);
xnor UO_411 (O_411,N_14914,N_14925);
and UO_412 (O_412,N_14815,N_14906);
xnor UO_413 (O_413,N_14933,N_14917);
xor UO_414 (O_414,N_14871,N_14907);
nand UO_415 (O_415,N_14883,N_14956);
xor UO_416 (O_416,N_14932,N_14929);
nor UO_417 (O_417,N_14978,N_14962);
nor UO_418 (O_418,N_14863,N_14902);
nand UO_419 (O_419,N_14864,N_14820);
or UO_420 (O_420,N_14822,N_14950);
or UO_421 (O_421,N_14902,N_14913);
and UO_422 (O_422,N_14913,N_14933);
nand UO_423 (O_423,N_14827,N_14913);
and UO_424 (O_424,N_14853,N_14876);
or UO_425 (O_425,N_14863,N_14835);
or UO_426 (O_426,N_14904,N_14851);
and UO_427 (O_427,N_14907,N_14966);
nand UO_428 (O_428,N_14987,N_14812);
nor UO_429 (O_429,N_14876,N_14946);
xor UO_430 (O_430,N_14937,N_14826);
and UO_431 (O_431,N_14922,N_14942);
or UO_432 (O_432,N_14838,N_14855);
or UO_433 (O_433,N_14916,N_14931);
or UO_434 (O_434,N_14846,N_14830);
xor UO_435 (O_435,N_14952,N_14853);
or UO_436 (O_436,N_14820,N_14995);
or UO_437 (O_437,N_14983,N_14961);
nand UO_438 (O_438,N_14833,N_14878);
and UO_439 (O_439,N_14982,N_14835);
xor UO_440 (O_440,N_14972,N_14945);
and UO_441 (O_441,N_14871,N_14870);
and UO_442 (O_442,N_14960,N_14850);
xor UO_443 (O_443,N_14869,N_14844);
nor UO_444 (O_444,N_14972,N_14995);
xor UO_445 (O_445,N_14879,N_14874);
and UO_446 (O_446,N_14892,N_14848);
and UO_447 (O_447,N_14955,N_14917);
xnor UO_448 (O_448,N_14960,N_14972);
or UO_449 (O_449,N_14929,N_14939);
or UO_450 (O_450,N_14994,N_14991);
xor UO_451 (O_451,N_14945,N_14843);
and UO_452 (O_452,N_14903,N_14884);
and UO_453 (O_453,N_14883,N_14968);
xor UO_454 (O_454,N_14900,N_14858);
nor UO_455 (O_455,N_14886,N_14853);
and UO_456 (O_456,N_14991,N_14812);
nor UO_457 (O_457,N_14897,N_14812);
and UO_458 (O_458,N_14875,N_14962);
xnor UO_459 (O_459,N_14840,N_14889);
xor UO_460 (O_460,N_14893,N_14900);
and UO_461 (O_461,N_14975,N_14842);
nor UO_462 (O_462,N_14931,N_14827);
xnor UO_463 (O_463,N_14874,N_14847);
nand UO_464 (O_464,N_14977,N_14943);
xnor UO_465 (O_465,N_14992,N_14980);
xor UO_466 (O_466,N_14937,N_14912);
xor UO_467 (O_467,N_14919,N_14813);
and UO_468 (O_468,N_14858,N_14808);
or UO_469 (O_469,N_14819,N_14876);
nor UO_470 (O_470,N_14858,N_14957);
or UO_471 (O_471,N_14830,N_14950);
nand UO_472 (O_472,N_14814,N_14929);
nor UO_473 (O_473,N_14824,N_14921);
nor UO_474 (O_474,N_14966,N_14823);
xnor UO_475 (O_475,N_14848,N_14935);
xnor UO_476 (O_476,N_14909,N_14905);
xor UO_477 (O_477,N_14824,N_14968);
nor UO_478 (O_478,N_14925,N_14923);
nor UO_479 (O_479,N_14855,N_14898);
or UO_480 (O_480,N_14953,N_14803);
and UO_481 (O_481,N_14897,N_14971);
and UO_482 (O_482,N_14921,N_14928);
and UO_483 (O_483,N_14992,N_14824);
xnor UO_484 (O_484,N_14859,N_14963);
nand UO_485 (O_485,N_14949,N_14868);
xnor UO_486 (O_486,N_14880,N_14916);
xor UO_487 (O_487,N_14922,N_14831);
or UO_488 (O_488,N_14828,N_14913);
or UO_489 (O_489,N_14964,N_14884);
nor UO_490 (O_490,N_14997,N_14948);
xnor UO_491 (O_491,N_14959,N_14930);
xor UO_492 (O_492,N_14979,N_14974);
nand UO_493 (O_493,N_14839,N_14984);
or UO_494 (O_494,N_14984,N_14849);
and UO_495 (O_495,N_14899,N_14824);
nor UO_496 (O_496,N_14894,N_14827);
and UO_497 (O_497,N_14845,N_14947);
nand UO_498 (O_498,N_14911,N_14987);
or UO_499 (O_499,N_14888,N_14897);
nor UO_500 (O_500,N_14883,N_14815);
xnor UO_501 (O_501,N_14928,N_14812);
nand UO_502 (O_502,N_14914,N_14811);
or UO_503 (O_503,N_14944,N_14949);
nor UO_504 (O_504,N_14922,N_14958);
xnor UO_505 (O_505,N_14944,N_14899);
or UO_506 (O_506,N_14988,N_14879);
nor UO_507 (O_507,N_14818,N_14870);
and UO_508 (O_508,N_14882,N_14896);
or UO_509 (O_509,N_14897,N_14807);
nand UO_510 (O_510,N_14912,N_14879);
or UO_511 (O_511,N_14881,N_14994);
xor UO_512 (O_512,N_14914,N_14958);
nor UO_513 (O_513,N_14988,N_14904);
and UO_514 (O_514,N_14892,N_14819);
xnor UO_515 (O_515,N_14967,N_14828);
nand UO_516 (O_516,N_14821,N_14873);
nor UO_517 (O_517,N_14939,N_14820);
or UO_518 (O_518,N_14873,N_14989);
or UO_519 (O_519,N_14856,N_14994);
xor UO_520 (O_520,N_14819,N_14878);
xor UO_521 (O_521,N_14825,N_14850);
and UO_522 (O_522,N_14861,N_14907);
nor UO_523 (O_523,N_14906,N_14824);
and UO_524 (O_524,N_14926,N_14936);
and UO_525 (O_525,N_14817,N_14935);
nor UO_526 (O_526,N_14809,N_14852);
nand UO_527 (O_527,N_14892,N_14944);
or UO_528 (O_528,N_14965,N_14806);
nand UO_529 (O_529,N_14931,N_14856);
nor UO_530 (O_530,N_14809,N_14982);
nand UO_531 (O_531,N_14973,N_14962);
xnor UO_532 (O_532,N_14803,N_14938);
nand UO_533 (O_533,N_14885,N_14994);
xnor UO_534 (O_534,N_14946,N_14812);
nand UO_535 (O_535,N_14899,N_14911);
xnor UO_536 (O_536,N_14853,N_14947);
xnor UO_537 (O_537,N_14932,N_14958);
and UO_538 (O_538,N_14992,N_14965);
nand UO_539 (O_539,N_14942,N_14980);
nor UO_540 (O_540,N_14994,N_14930);
nand UO_541 (O_541,N_14960,N_14808);
and UO_542 (O_542,N_14898,N_14865);
nor UO_543 (O_543,N_14829,N_14998);
xor UO_544 (O_544,N_14810,N_14858);
xnor UO_545 (O_545,N_14930,N_14970);
or UO_546 (O_546,N_14931,N_14970);
xnor UO_547 (O_547,N_14932,N_14994);
nand UO_548 (O_548,N_14879,N_14823);
xor UO_549 (O_549,N_14826,N_14898);
nor UO_550 (O_550,N_14868,N_14941);
or UO_551 (O_551,N_14897,N_14865);
xor UO_552 (O_552,N_14835,N_14974);
or UO_553 (O_553,N_14965,N_14915);
xor UO_554 (O_554,N_14994,N_14844);
and UO_555 (O_555,N_14867,N_14917);
or UO_556 (O_556,N_14994,N_14819);
xor UO_557 (O_557,N_14933,N_14827);
and UO_558 (O_558,N_14827,N_14999);
nor UO_559 (O_559,N_14828,N_14928);
or UO_560 (O_560,N_14977,N_14862);
and UO_561 (O_561,N_14898,N_14951);
or UO_562 (O_562,N_14846,N_14800);
xnor UO_563 (O_563,N_14964,N_14863);
or UO_564 (O_564,N_14807,N_14829);
or UO_565 (O_565,N_14832,N_14988);
nand UO_566 (O_566,N_14983,N_14828);
xor UO_567 (O_567,N_14869,N_14984);
or UO_568 (O_568,N_14908,N_14817);
or UO_569 (O_569,N_14857,N_14943);
nand UO_570 (O_570,N_14911,N_14863);
nand UO_571 (O_571,N_14835,N_14882);
nor UO_572 (O_572,N_14884,N_14973);
and UO_573 (O_573,N_14815,N_14981);
nand UO_574 (O_574,N_14983,N_14823);
and UO_575 (O_575,N_14883,N_14988);
nand UO_576 (O_576,N_14950,N_14867);
xor UO_577 (O_577,N_14928,N_14936);
xor UO_578 (O_578,N_14830,N_14887);
and UO_579 (O_579,N_14944,N_14872);
nand UO_580 (O_580,N_14858,N_14987);
nor UO_581 (O_581,N_14982,N_14922);
xnor UO_582 (O_582,N_14952,N_14809);
nand UO_583 (O_583,N_14989,N_14909);
xor UO_584 (O_584,N_14946,N_14838);
and UO_585 (O_585,N_14887,N_14859);
nand UO_586 (O_586,N_14866,N_14962);
and UO_587 (O_587,N_14931,N_14926);
and UO_588 (O_588,N_14986,N_14978);
nor UO_589 (O_589,N_14807,N_14956);
xor UO_590 (O_590,N_14838,N_14930);
and UO_591 (O_591,N_14996,N_14852);
and UO_592 (O_592,N_14980,N_14954);
xor UO_593 (O_593,N_14989,N_14980);
nand UO_594 (O_594,N_14859,N_14954);
nand UO_595 (O_595,N_14892,N_14876);
nand UO_596 (O_596,N_14861,N_14804);
xnor UO_597 (O_597,N_14920,N_14922);
or UO_598 (O_598,N_14806,N_14888);
nor UO_599 (O_599,N_14886,N_14943);
and UO_600 (O_600,N_14830,N_14939);
xor UO_601 (O_601,N_14959,N_14836);
nand UO_602 (O_602,N_14831,N_14837);
and UO_603 (O_603,N_14983,N_14856);
or UO_604 (O_604,N_14824,N_14858);
nor UO_605 (O_605,N_14830,N_14910);
or UO_606 (O_606,N_14820,N_14822);
nand UO_607 (O_607,N_14864,N_14985);
or UO_608 (O_608,N_14946,N_14920);
nor UO_609 (O_609,N_14867,N_14825);
xnor UO_610 (O_610,N_14880,N_14999);
nor UO_611 (O_611,N_14800,N_14885);
nor UO_612 (O_612,N_14907,N_14878);
and UO_613 (O_613,N_14877,N_14974);
or UO_614 (O_614,N_14953,N_14811);
xnor UO_615 (O_615,N_14920,N_14998);
and UO_616 (O_616,N_14993,N_14899);
xnor UO_617 (O_617,N_14899,N_14893);
or UO_618 (O_618,N_14881,N_14877);
xnor UO_619 (O_619,N_14826,N_14915);
nand UO_620 (O_620,N_14805,N_14940);
or UO_621 (O_621,N_14854,N_14817);
or UO_622 (O_622,N_14943,N_14926);
and UO_623 (O_623,N_14996,N_14832);
or UO_624 (O_624,N_14991,N_14841);
nand UO_625 (O_625,N_14956,N_14846);
nor UO_626 (O_626,N_14986,N_14932);
or UO_627 (O_627,N_14825,N_14810);
xnor UO_628 (O_628,N_14906,N_14986);
and UO_629 (O_629,N_14993,N_14803);
nor UO_630 (O_630,N_14821,N_14919);
nor UO_631 (O_631,N_14898,N_14965);
nand UO_632 (O_632,N_14812,N_14939);
xor UO_633 (O_633,N_14887,N_14993);
xnor UO_634 (O_634,N_14829,N_14818);
nor UO_635 (O_635,N_14933,N_14837);
nor UO_636 (O_636,N_14965,N_14918);
nand UO_637 (O_637,N_14878,N_14886);
nor UO_638 (O_638,N_14985,N_14807);
and UO_639 (O_639,N_14932,N_14871);
and UO_640 (O_640,N_14915,N_14877);
nor UO_641 (O_641,N_14903,N_14904);
and UO_642 (O_642,N_14881,N_14980);
nor UO_643 (O_643,N_14965,N_14954);
nor UO_644 (O_644,N_14992,N_14958);
or UO_645 (O_645,N_14999,N_14963);
xor UO_646 (O_646,N_14883,N_14913);
and UO_647 (O_647,N_14889,N_14995);
nor UO_648 (O_648,N_14821,N_14998);
and UO_649 (O_649,N_14868,N_14950);
nor UO_650 (O_650,N_14996,N_14860);
or UO_651 (O_651,N_14898,N_14871);
nor UO_652 (O_652,N_14998,N_14817);
nand UO_653 (O_653,N_14836,N_14910);
nand UO_654 (O_654,N_14953,N_14835);
or UO_655 (O_655,N_14963,N_14967);
nand UO_656 (O_656,N_14911,N_14993);
and UO_657 (O_657,N_14951,N_14832);
xnor UO_658 (O_658,N_14937,N_14914);
nand UO_659 (O_659,N_14882,N_14970);
nor UO_660 (O_660,N_14869,N_14968);
and UO_661 (O_661,N_14936,N_14855);
nor UO_662 (O_662,N_14849,N_14894);
and UO_663 (O_663,N_14987,N_14939);
nand UO_664 (O_664,N_14801,N_14909);
or UO_665 (O_665,N_14820,N_14842);
xor UO_666 (O_666,N_14886,N_14837);
nand UO_667 (O_667,N_14987,N_14899);
or UO_668 (O_668,N_14880,N_14885);
and UO_669 (O_669,N_14994,N_14936);
xor UO_670 (O_670,N_14891,N_14955);
and UO_671 (O_671,N_14904,N_14956);
nor UO_672 (O_672,N_14949,N_14858);
and UO_673 (O_673,N_14955,N_14893);
xnor UO_674 (O_674,N_14819,N_14824);
nand UO_675 (O_675,N_14928,N_14986);
nor UO_676 (O_676,N_14907,N_14995);
nand UO_677 (O_677,N_14981,N_14923);
xor UO_678 (O_678,N_14983,N_14894);
and UO_679 (O_679,N_14902,N_14989);
and UO_680 (O_680,N_14836,N_14987);
nand UO_681 (O_681,N_14992,N_14943);
and UO_682 (O_682,N_14982,N_14990);
and UO_683 (O_683,N_14853,N_14926);
and UO_684 (O_684,N_14843,N_14869);
xnor UO_685 (O_685,N_14948,N_14813);
nor UO_686 (O_686,N_14808,N_14947);
nor UO_687 (O_687,N_14930,N_14867);
and UO_688 (O_688,N_14889,N_14856);
or UO_689 (O_689,N_14829,N_14900);
xnor UO_690 (O_690,N_14994,N_14943);
nor UO_691 (O_691,N_14910,N_14802);
or UO_692 (O_692,N_14902,N_14960);
nor UO_693 (O_693,N_14828,N_14912);
or UO_694 (O_694,N_14991,N_14961);
and UO_695 (O_695,N_14896,N_14919);
and UO_696 (O_696,N_14962,N_14803);
nand UO_697 (O_697,N_14904,N_14813);
or UO_698 (O_698,N_14966,N_14970);
and UO_699 (O_699,N_14993,N_14973);
xor UO_700 (O_700,N_14877,N_14953);
or UO_701 (O_701,N_14820,N_14908);
nand UO_702 (O_702,N_14860,N_14972);
and UO_703 (O_703,N_14894,N_14915);
nor UO_704 (O_704,N_14935,N_14840);
or UO_705 (O_705,N_14907,N_14805);
and UO_706 (O_706,N_14866,N_14988);
and UO_707 (O_707,N_14856,N_14854);
nand UO_708 (O_708,N_14912,N_14942);
nand UO_709 (O_709,N_14881,N_14861);
nor UO_710 (O_710,N_14861,N_14806);
or UO_711 (O_711,N_14819,N_14959);
nor UO_712 (O_712,N_14890,N_14860);
nor UO_713 (O_713,N_14919,N_14890);
and UO_714 (O_714,N_14830,N_14821);
nor UO_715 (O_715,N_14943,N_14915);
and UO_716 (O_716,N_14977,N_14812);
nor UO_717 (O_717,N_14819,N_14865);
nor UO_718 (O_718,N_14851,N_14992);
xnor UO_719 (O_719,N_14894,N_14832);
xnor UO_720 (O_720,N_14860,N_14841);
nor UO_721 (O_721,N_14929,N_14872);
xor UO_722 (O_722,N_14969,N_14979);
and UO_723 (O_723,N_14990,N_14915);
and UO_724 (O_724,N_14817,N_14902);
and UO_725 (O_725,N_14822,N_14900);
nand UO_726 (O_726,N_14826,N_14829);
or UO_727 (O_727,N_14855,N_14948);
and UO_728 (O_728,N_14973,N_14852);
nand UO_729 (O_729,N_14930,N_14804);
or UO_730 (O_730,N_14956,N_14907);
nor UO_731 (O_731,N_14962,N_14840);
and UO_732 (O_732,N_14934,N_14876);
and UO_733 (O_733,N_14836,N_14829);
or UO_734 (O_734,N_14905,N_14956);
nand UO_735 (O_735,N_14995,N_14844);
xor UO_736 (O_736,N_14869,N_14806);
xnor UO_737 (O_737,N_14951,N_14996);
nand UO_738 (O_738,N_14800,N_14834);
nor UO_739 (O_739,N_14863,N_14893);
and UO_740 (O_740,N_14850,N_14895);
nor UO_741 (O_741,N_14987,N_14898);
and UO_742 (O_742,N_14828,N_14910);
xnor UO_743 (O_743,N_14819,N_14919);
and UO_744 (O_744,N_14806,N_14945);
xor UO_745 (O_745,N_14971,N_14809);
xnor UO_746 (O_746,N_14880,N_14924);
and UO_747 (O_747,N_14867,N_14830);
and UO_748 (O_748,N_14867,N_14810);
and UO_749 (O_749,N_14846,N_14972);
or UO_750 (O_750,N_14832,N_14835);
and UO_751 (O_751,N_14885,N_14876);
nor UO_752 (O_752,N_14807,N_14866);
nand UO_753 (O_753,N_14907,N_14880);
nand UO_754 (O_754,N_14827,N_14951);
nand UO_755 (O_755,N_14943,N_14965);
nand UO_756 (O_756,N_14961,N_14811);
nor UO_757 (O_757,N_14919,N_14960);
xnor UO_758 (O_758,N_14882,N_14991);
or UO_759 (O_759,N_14979,N_14900);
or UO_760 (O_760,N_14992,N_14825);
xnor UO_761 (O_761,N_14845,N_14813);
nand UO_762 (O_762,N_14937,N_14855);
or UO_763 (O_763,N_14829,N_14902);
xor UO_764 (O_764,N_14842,N_14826);
nor UO_765 (O_765,N_14849,N_14886);
nor UO_766 (O_766,N_14835,N_14987);
nor UO_767 (O_767,N_14848,N_14800);
nor UO_768 (O_768,N_14945,N_14884);
nand UO_769 (O_769,N_14946,N_14961);
or UO_770 (O_770,N_14898,N_14882);
or UO_771 (O_771,N_14959,N_14925);
nor UO_772 (O_772,N_14917,N_14988);
nand UO_773 (O_773,N_14938,N_14861);
xor UO_774 (O_774,N_14837,N_14806);
and UO_775 (O_775,N_14814,N_14819);
nand UO_776 (O_776,N_14927,N_14929);
nor UO_777 (O_777,N_14969,N_14915);
or UO_778 (O_778,N_14802,N_14960);
nand UO_779 (O_779,N_14863,N_14886);
xnor UO_780 (O_780,N_14954,N_14947);
nor UO_781 (O_781,N_14844,N_14842);
and UO_782 (O_782,N_14808,N_14973);
nor UO_783 (O_783,N_14826,N_14873);
and UO_784 (O_784,N_14893,N_14924);
xor UO_785 (O_785,N_14895,N_14875);
xor UO_786 (O_786,N_14929,N_14852);
xnor UO_787 (O_787,N_14999,N_14896);
nor UO_788 (O_788,N_14915,N_14853);
xor UO_789 (O_789,N_14975,N_14946);
nand UO_790 (O_790,N_14973,N_14976);
xor UO_791 (O_791,N_14839,N_14905);
xor UO_792 (O_792,N_14818,N_14816);
or UO_793 (O_793,N_14984,N_14815);
or UO_794 (O_794,N_14910,N_14960);
nand UO_795 (O_795,N_14891,N_14909);
nor UO_796 (O_796,N_14944,N_14806);
or UO_797 (O_797,N_14920,N_14894);
nand UO_798 (O_798,N_14975,N_14950);
or UO_799 (O_799,N_14970,N_14805);
nand UO_800 (O_800,N_14925,N_14986);
nand UO_801 (O_801,N_14947,N_14848);
nor UO_802 (O_802,N_14980,N_14818);
nand UO_803 (O_803,N_14961,N_14997);
nor UO_804 (O_804,N_14960,N_14945);
xor UO_805 (O_805,N_14874,N_14819);
xor UO_806 (O_806,N_14850,N_14872);
nand UO_807 (O_807,N_14973,N_14820);
or UO_808 (O_808,N_14971,N_14957);
or UO_809 (O_809,N_14988,N_14905);
xor UO_810 (O_810,N_14924,N_14915);
xnor UO_811 (O_811,N_14998,N_14831);
or UO_812 (O_812,N_14890,N_14841);
xor UO_813 (O_813,N_14802,N_14819);
or UO_814 (O_814,N_14875,N_14987);
xor UO_815 (O_815,N_14827,N_14882);
nor UO_816 (O_816,N_14886,N_14844);
nand UO_817 (O_817,N_14926,N_14991);
or UO_818 (O_818,N_14802,N_14847);
or UO_819 (O_819,N_14911,N_14982);
and UO_820 (O_820,N_14960,N_14856);
nand UO_821 (O_821,N_14904,N_14930);
or UO_822 (O_822,N_14958,N_14859);
xnor UO_823 (O_823,N_14936,N_14859);
nand UO_824 (O_824,N_14919,N_14814);
and UO_825 (O_825,N_14918,N_14860);
or UO_826 (O_826,N_14900,N_14943);
and UO_827 (O_827,N_14828,N_14821);
nor UO_828 (O_828,N_14958,N_14885);
or UO_829 (O_829,N_14964,N_14902);
nor UO_830 (O_830,N_14985,N_14844);
xnor UO_831 (O_831,N_14965,N_14928);
and UO_832 (O_832,N_14951,N_14807);
and UO_833 (O_833,N_14877,N_14817);
xor UO_834 (O_834,N_14958,N_14993);
nor UO_835 (O_835,N_14924,N_14847);
nand UO_836 (O_836,N_14833,N_14828);
nand UO_837 (O_837,N_14931,N_14963);
nand UO_838 (O_838,N_14801,N_14882);
nand UO_839 (O_839,N_14921,N_14941);
nor UO_840 (O_840,N_14912,N_14887);
or UO_841 (O_841,N_14927,N_14994);
or UO_842 (O_842,N_14906,N_14887);
and UO_843 (O_843,N_14806,N_14969);
or UO_844 (O_844,N_14804,N_14829);
nand UO_845 (O_845,N_14886,N_14962);
or UO_846 (O_846,N_14983,N_14966);
or UO_847 (O_847,N_14981,N_14950);
or UO_848 (O_848,N_14853,N_14882);
nand UO_849 (O_849,N_14988,N_14920);
and UO_850 (O_850,N_14931,N_14875);
nand UO_851 (O_851,N_14894,N_14999);
or UO_852 (O_852,N_14919,N_14999);
nor UO_853 (O_853,N_14976,N_14974);
nand UO_854 (O_854,N_14856,N_14918);
nand UO_855 (O_855,N_14886,N_14893);
and UO_856 (O_856,N_14842,N_14929);
nor UO_857 (O_857,N_14936,N_14844);
and UO_858 (O_858,N_14807,N_14919);
nand UO_859 (O_859,N_14956,N_14917);
and UO_860 (O_860,N_14971,N_14906);
xor UO_861 (O_861,N_14839,N_14889);
nor UO_862 (O_862,N_14952,N_14805);
or UO_863 (O_863,N_14834,N_14888);
xor UO_864 (O_864,N_14932,N_14991);
or UO_865 (O_865,N_14842,N_14907);
or UO_866 (O_866,N_14993,N_14896);
nand UO_867 (O_867,N_14943,N_14947);
or UO_868 (O_868,N_14980,N_14844);
and UO_869 (O_869,N_14919,N_14901);
or UO_870 (O_870,N_14940,N_14831);
xor UO_871 (O_871,N_14993,N_14865);
and UO_872 (O_872,N_14988,N_14871);
or UO_873 (O_873,N_14954,N_14914);
or UO_874 (O_874,N_14858,N_14941);
and UO_875 (O_875,N_14837,N_14991);
nor UO_876 (O_876,N_14941,N_14820);
nor UO_877 (O_877,N_14821,N_14868);
nand UO_878 (O_878,N_14843,N_14990);
nand UO_879 (O_879,N_14889,N_14805);
and UO_880 (O_880,N_14968,N_14960);
nand UO_881 (O_881,N_14809,N_14994);
nor UO_882 (O_882,N_14947,N_14869);
or UO_883 (O_883,N_14978,N_14816);
nand UO_884 (O_884,N_14987,N_14890);
nor UO_885 (O_885,N_14814,N_14853);
and UO_886 (O_886,N_14895,N_14817);
and UO_887 (O_887,N_14917,N_14944);
or UO_888 (O_888,N_14945,N_14848);
nand UO_889 (O_889,N_14852,N_14897);
xor UO_890 (O_890,N_14933,N_14809);
nand UO_891 (O_891,N_14936,N_14811);
nor UO_892 (O_892,N_14929,N_14961);
nand UO_893 (O_893,N_14943,N_14854);
and UO_894 (O_894,N_14917,N_14824);
nand UO_895 (O_895,N_14841,N_14989);
nor UO_896 (O_896,N_14906,N_14812);
or UO_897 (O_897,N_14805,N_14839);
or UO_898 (O_898,N_14919,N_14881);
and UO_899 (O_899,N_14893,N_14906);
nor UO_900 (O_900,N_14969,N_14876);
nand UO_901 (O_901,N_14873,N_14913);
or UO_902 (O_902,N_14826,N_14827);
xor UO_903 (O_903,N_14920,N_14829);
nand UO_904 (O_904,N_14890,N_14907);
or UO_905 (O_905,N_14942,N_14959);
or UO_906 (O_906,N_14897,N_14995);
nor UO_907 (O_907,N_14836,N_14888);
xnor UO_908 (O_908,N_14958,N_14820);
nand UO_909 (O_909,N_14894,N_14958);
nand UO_910 (O_910,N_14811,N_14947);
xnor UO_911 (O_911,N_14976,N_14888);
nand UO_912 (O_912,N_14901,N_14938);
and UO_913 (O_913,N_14861,N_14812);
nand UO_914 (O_914,N_14832,N_14810);
nand UO_915 (O_915,N_14983,N_14893);
nor UO_916 (O_916,N_14815,N_14816);
nor UO_917 (O_917,N_14851,N_14917);
and UO_918 (O_918,N_14807,N_14822);
nor UO_919 (O_919,N_14940,N_14836);
nor UO_920 (O_920,N_14945,N_14877);
xnor UO_921 (O_921,N_14968,N_14846);
and UO_922 (O_922,N_14923,N_14835);
and UO_923 (O_923,N_14938,N_14801);
or UO_924 (O_924,N_14872,N_14902);
nand UO_925 (O_925,N_14849,N_14996);
nor UO_926 (O_926,N_14927,N_14925);
xnor UO_927 (O_927,N_14817,N_14973);
or UO_928 (O_928,N_14980,N_14801);
or UO_929 (O_929,N_14801,N_14993);
nand UO_930 (O_930,N_14875,N_14816);
or UO_931 (O_931,N_14827,N_14812);
nor UO_932 (O_932,N_14918,N_14956);
xnor UO_933 (O_933,N_14862,N_14920);
xnor UO_934 (O_934,N_14926,N_14824);
nor UO_935 (O_935,N_14851,N_14852);
nand UO_936 (O_936,N_14897,N_14879);
nand UO_937 (O_937,N_14836,N_14805);
nand UO_938 (O_938,N_14955,N_14832);
or UO_939 (O_939,N_14967,N_14920);
nor UO_940 (O_940,N_14871,N_14950);
nand UO_941 (O_941,N_14965,N_14870);
or UO_942 (O_942,N_14908,N_14885);
xnor UO_943 (O_943,N_14843,N_14858);
nand UO_944 (O_944,N_14825,N_14844);
and UO_945 (O_945,N_14886,N_14981);
xnor UO_946 (O_946,N_14917,N_14976);
nor UO_947 (O_947,N_14854,N_14993);
or UO_948 (O_948,N_14944,N_14947);
or UO_949 (O_949,N_14959,N_14966);
nand UO_950 (O_950,N_14850,N_14904);
nand UO_951 (O_951,N_14880,N_14891);
nor UO_952 (O_952,N_14836,N_14889);
and UO_953 (O_953,N_14990,N_14849);
and UO_954 (O_954,N_14803,N_14954);
xor UO_955 (O_955,N_14927,N_14932);
nor UO_956 (O_956,N_14977,N_14975);
or UO_957 (O_957,N_14802,N_14940);
nand UO_958 (O_958,N_14826,N_14992);
xnor UO_959 (O_959,N_14848,N_14942);
nand UO_960 (O_960,N_14873,N_14927);
xor UO_961 (O_961,N_14931,N_14986);
nand UO_962 (O_962,N_14822,N_14934);
nand UO_963 (O_963,N_14849,N_14930);
xnor UO_964 (O_964,N_14951,N_14959);
nand UO_965 (O_965,N_14806,N_14862);
nor UO_966 (O_966,N_14853,N_14828);
nand UO_967 (O_967,N_14873,N_14984);
and UO_968 (O_968,N_14910,N_14801);
nand UO_969 (O_969,N_14986,N_14913);
and UO_970 (O_970,N_14819,N_14886);
and UO_971 (O_971,N_14871,N_14925);
xnor UO_972 (O_972,N_14899,N_14974);
nor UO_973 (O_973,N_14933,N_14843);
xor UO_974 (O_974,N_14851,N_14813);
or UO_975 (O_975,N_14900,N_14842);
xor UO_976 (O_976,N_14889,N_14825);
or UO_977 (O_977,N_14963,N_14985);
nand UO_978 (O_978,N_14970,N_14985);
nand UO_979 (O_979,N_14939,N_14931);
or UO_980 (O_980,N_14953,N_14838);
xor UO_981 (O_981,N_14982,N_14970);
nor UO_982 (O_982,N_14912,N_14951);
nand UO_983 (O_983,N_14853,N_14889);
nand UO_984 (O_984,N_14970,N_14937);
nor UO_985 (O_985,N_14966,N_14816);
nand UO_986 (O_986,N_14826,N_14830);
and UO_987 (O_987,N_14871,N_14803);
or UO_988 (O_988,N_14987,N_14959);
nand UO_989 (O_989,N_14900,N_14932);
nor UO_990 (O_990,N_14934,N_14994);
and UO_991 (O_991,N_14823,N_14847);
nor UO_992 (O_992,N_14866,N_14983);
nand UO_993 (O_993,N_14935,N_14980);
or UO_994 (O_994,N_14875,N_14844);
or UO_995 (O_995,N_14912,N_14927);
xnor UO_996 (O_996,N_14963,N_14914);
or UO_997 (O_997,N_14978,N_14997);
or UO_998 (O_998,N_14997,N_14933);
and UO_999 (O_999,N_14887,N_14971);
xnor UO_1000 (O_1000,N_14897,N_14985);
nand UO_1001 (O_1001,N_14821,N_14970);
and UO_1002 (O_1002,N_14879,N_14878);
nor UO_1003 (O_1003,N_14835,N_14888);
xor UO_1004 (O_1004,N_14813,N_14837);
and UO_1005 (O_1005,N_14828,N_14973);
and UO_1006 (O_1006,N_14983,N_14915);
and UO_1007 (O_1007,N_14884,N_14984);
and UO_1008 (O_1008,N_14945,N_14955);
nor UO_1009 (O_1009,N_14808,N_14834);
nor UO_1010 (O_1010,N_14991,N_14944);
and UO_1011 (O_1011,N_14990,N_14831);
and UO_1012 (O_1012,N_14890,N_14894);
and UO_1013 (O_1013,N_14944,N_14861);
xnor UO_1014 (O_1014,N_14990,N_14807);
and UO_1015 (O_1015,N_14889,N_14872);
nor UO_1016 (O_1016,N_14810,N_14939);
or UO_1017 (O_1017,N_14966,N_14899);
nor UO_1018 (O_1018,N_14951,N_14990);
nand UO_1019 (O_1019,N_14976,N_14818);
xnor UO_1020 (O_1020,N_14886,N_14828);
or UO_1021 (O_1021,N_14849,N_14809);
nor UO_1022 (O_1022,N_14870,N_14981);
xor UO_1023 (O_1023,N_14935,N_14892);
or UO_1024 (O_1024,N_14916,N_14963);
xor UO_1025 (O_1025,N_14871,N_14912);
xnor UO_1026 (O_1026,N_14963,N_14839);
nor UO_1027 (O_1027,N_14850,N_14907);
nand UO_1028 (O_1028,N_14877,N_14968);
nor UO_1029 (O_1029,N_14855,N_14910);
nor UO_1030 (O_1030,N_14861,N_14993);
or UO_1031 (O_1031,N_14853,N_14850);
or UO_1032 (O_1032,N_14948,N_14913);
or UO_1033 (O_1033,N_14935,N_14812);
nand UO_1034 (O_1034,N_14847,N_14916);
or UO_1035 (O_1035,N_14866,N_14878);
and UO_1036 (O_1036,N_14877,N_14869);
and UO_1037 (O_1037,N_14800,N_14971);
nand UO_1038 (O_1038,N_14862,N_14870);
nand UO_1039 (O_1039,N_14962,N_14869);
or UO_1040 (O_1040,N_14908,N_14945);
nor UO_1041 (O_1041,N_14948,N_14889);
nand UO_1042 (O_1042,N_14839,N_14940);
nor UO_1043 (O_1043,N_14922,N_14936);
nor UO_1044 (O_1044,N_14836,N_14856);
or UO_1045 (O_1045,N_14888,N_14825);
and UO_1046 (O_1046,N_14892,N_14969);
nor UO_1047 (O_1047,N_14919,N_14930);
and UO_1048 (O_1048,N_14843,N_14850);
or UO_1049 (O_1049,N_14913,N_14917);
or UO_1050 (O_1050,N_14810,N_14815);
xor UO_1051 (O_1051,N_14909,N_14828);
nand UO_1052 (O_1052,N_14868,N_14994);
and UO_1053 (O_1053,N_14887,N_14827);
xnor UO_1054 (O_1054,N_14962,N_14809);
or UO_1055 (O_1055,N_14952,N_14888);
nor UO_1056 (O_1056,N_14932,N_14965);
xor UO_1057 (O_1057,N_14803,N_14840);
nor UO_1058 (O_1058,N_14907,N_14810);
xor UO_1059 (O_1059,N_14982,N_14841);
xor UO_1060 (O_1060,N_14901,N_14973);
nand UO_1061 (O_1061,N_14931,N_14981);
and UO_1062 (O_1062,N_14916,N_14897);
xor UO_1063 (O_1063,N_14820,N_14896);
or UO_1064 (O_1064,N_14943,N_14865);
or UO_1065 (O_1065,N_14997,N_14897);
or UO_1066 (O_1066,N_14852,N_14923);
xnor UO_1067 (O_1067,N_14804,N_14973);
nand UO_1068 (O_1068,N_14891,N_14839);
nor UO_1069 (O_1069,N_14880,N_14826);
nand UO_1070 (O_1070,N_14985,N_14878);
and UO_1071 (O_1071,N_14937,N_14816);
and UO_1072 (O_1072,N_14816,N_14887);
xor UO_1073 (O_1073,N_14880,N_14949);
nor UO_1074 (O_1074,N_14937,N_14805);
nand UO_1075 (O_1075,N_14811,N_14871);
xnor UO_1076 (O_1076,N_14935,N_14866);
nor UO_1077 (O_1077,N_14848,N_14985);
nand UO_1078 (O_1078,N_14982,N_14998);
or UO_1079 (O_1079,N_14831,N_14914);
or UO_1080 (O_1080,N_14887,N_14867);
xor UO_1081 (O_1081,N_14892,N_14906);
nor UO_1082 (O_1082,N_14871,N_14867);
xor UO_1083 (O_1083,N_14995,N_14933);
nor UO_1084 (O_1084,N_14872,N_14961);
or UO_1085 (O_1085,N_14983,N_14996);
nand UO_1086 (O_1086,N_14863,N_14950);
nor UO_1087 (O_1087,N_14943,N_14871);
or UO_1088 (O_1088,N_14912,N_14840);
nor UO_1089 (O_1089,N_14941,N_14805);
and UO_1090 (O_1090,N_14916,N_14983);
nand UO_1091 (O_1091,N_14877,N_14868);
nor UO_1092 (O_1092,N_14901,N_14821);
nor UO_1093 (O_1093,N_14887,N_14947);
nand UO_1094 (O_1094,N_14911,N_14940);
nor UO_1095 (O_1095,N_14916,N_14865);
xnor UO_1096 (O_1096,N_14896,N_14906);
or UO_1097 (O_1097,N_14988,N_14943);
or UO_1098 (O_1098,N_14850,N_14811);
nor UO_1099 (O_1099,N_14994,N_14944);
xnor UO_1100 (O_1100,N_14957,N_14963);
nand UO_1101 (O_1101,N_14929,N_14827);
and UO_1102 (O_1102,N_14884,N_14931);
xnor UO_1103 (O_1103,N_14980,N_14949);
or UO_1104 (O_1104,N_14811,N_14866);
and UO_1105 (O_1105,N_14896,N_14925);
or UO_1106 (O_1106,N_14858,N_14892);
or UO_1107 (O_1107,N_14860,N_14994);
nand UO_1108 (O_1108,N_14900,N_14865);
xnor UO_1109 (O_1109,N_14856,N_14838);
nor UO_1110 (O_1110,N_14945,N_14925);
nand UO_1111 (O_1111,N_14837,N_14989);
or UO_1112 (O_1112,N_14927,N_14910);
nand UO_1113 (O_1113,N_14987,N_14817);
nand UO_1114 (O_1114,N_14844,N_14971);
nor UO_1115 (O_1115,N_14902,N_14848);
or UO_1116 (O_1116,N_14998,N_14969);
or UO_1117 (O_1117,N_14993,N_14875);
nand UO_1118 (O_1118,N_14892,N_14945);
and UO_1119 (O_1119,N_14825,N_14925);
or UO_1120 (O_1120,N_14876,N_14809);
xnor UO_1121 (O_1121,N_14927,N_14957);
and UO_1122 (O_1122,N_14856,N_14848);
or UO_1123 (O_1123,N_14990,N_14866);
nor UO_1124 (O_1124,N_14900,N_14831);
nor UO_1125 (O_1125,N_14838,N_14981);
nor UO_1126 (O_1126,N_14819,N_14982);
xor UO_1127 (O_1127,N_14927,N_14979);
nor UO_1128 (O_1128,N_14836,N_14842);
nand UO_1129 (O_1129,N_14926,N_14890);
xor UO_1130 (O_1130,N_14955,N_14833);
nor UO_1131 (O_1131,N_14801,N_14922);
and UO_1132 (O_1132,N_14813,N_14838);
or UO_1133 (O_1133,N_14888,N_14890);
and UO_1134 (O_1134,N_14862,N_14952);
and UO_1135 (O_1135,N_14912,N_14946);
xor UO_1136 (O_1136,N_14813,N_14814);
nor UO_1137 (O_1137,N_14984,N_14963);
xnor UO_1138 (O_1138,N_14922,N_14814);
or UO_1139 (O_1139,N_14977,N_14924);
xnor UO_1140 (O_1140,N_14865,N_14864);
nor UO_1141 (O_1141,N_14826,N_14874);
or UO_1142 (O_1142,N_14844,N_14979);
nor UO_1143 (O_1143,N_14992,N_14821);
and UO_1144 (O_1144,N_14881,N_14852);
nand UO_1145 (O_1145,N_14967,N_14882);
xnor UO_1146 (O_1146,N_14971,N_14961);
nor UO_1147 (O_1147,N_14979,N_14863);
and UO_1148 (O_1148,N_14884,N_14947);
xnor UO_1149 (O_1149,N_14983,N_14901);
and UO_1150 (O_1150,N_14948,N_14965);
or UO_1151 (O_1151,N_14811,N_14939);
nor UO_1152 (O_1152,N_14866,N_14837);
nor UO_1153 (O_1153,N_14832,N_14877);
nand UO_1154 (O_1154,N_14806,N_14960);
xnor UO_1155 (O_1155,N_14969,N_14821);
xnor UO_1156 (O_1156,N_14884,N_14812);
xor UO_1157 (O_1157,N_14848,N_14995);
nor UO_1158 (O_1158,N_14921,N_14945);
or UO_1159 (O_1159,N_14844,N_14904);
nor UO_1160 (O_1160,N_14939,N_14920);
or UO_1161 (O_1161,N_14983,N_14878);
and UO_1162 (O_1162,N_14927,N_14831);
nor UO_1163 (O_1163,N_14866,N_14885);
and UO_1164 (O_1164,N_14881,N_14872);
or UO_1165 (O_1165,N_14903,N_14824);
nand UO_1166 (O_1166,N_14970,N_14969);
nor UO_1167 (O_1167,N_14949,N_14955);
and UO_1168 (O_1168,N_14959,N_14927);
xor UO_1169 (O_1169,N_14911,N_14928);
nand UO_1170 (O_1170,N_14818,N_14826);
nor UO_1171 (O_1171,N_14951,N_14889);
nor UO_1172 (O_1172,N_14871,N_14842);
xor UO_1173 (O_1173,N_14837,N_14896);
xor UO_1174 (O_1174,N_14857,N_14965);
or UO_1175 (O_1175,N_14842,N_14906);
or UO_1176 (O_1176,N_14922,N_14962);
nand UO_1177 (O_1177,N_14918,N_14851);
nor UO_1178 (O_1178,N_14846,N_14947);
nand UO_1179 (O_1179,N_14802,N_14913);
nand UO_1180 (O_1180,N_14940,N_14879);
xnor UO_1181 (O_1181,N_14835,N_14824);
or UO_1182 (O_1182,N_14955,N_14809);
xor UO_1183 (O_1183,N_14900,N_14824);
nand UO_1184 (O_1184,N_14904,N_14973);
nor UO_1185 (O_1185,N_14860,N_14917);
xnor UO_1186 (O_1186,N_14903,N_14869);
or UO_1187 (O_1187,N_14877,N_14941);
xor UO_1188 (O_1188,N_14821,N_14857);
nand UO_1189 (O_1189,N_14943,N_14892);
nand UO_1190 (O_1190,N_14962,N_14995);
and UO_1191 (O_1191,N_14816,N_14991);
or UO_1192 (O_1192,N_14933,N_14813);
xor UO_1193 (O_1193,N_14846,N_14955);
xor UO_1194 (O_1194,N_14857,N_14860);
and UO_1195 (O_1195,N_14821,N_14825);
or UO_1196 (O_1196,N_14847,N_14856);
nor UO_1197 (O_1197,N_14853,N_14827);
or UO_1198 (O_1198,N_14982,N_14919);
nor UO_1199 (O_1199,N_14939,N_14908);
and UO_1200 (O_1200,N_14926,N_14920);
or UO_1201 (O_1201,N_14814,N_14880);
xor UO_1202 (O_1202,N_14988,N_14851);
xor UO_1203 (O_1203,N_14882,N_14949);
and UO_1204 (O_1204,N_14988,N_14927);
and UO_1205 (O_1205,N_14905,N_14993);
nor UO_1206 (O_1206,N_14975,N_14858);
or UO_1207 (O_1207,N_14992,N_14936);
nor UO_1208 (O_1208,N_14929,N_14815);
nand UO_1209 (O_1209,N_14964,N_14960);
nor UO_1210 (O_1210,N_14937,N_14864);
xor UO_1211 (O_1211,N_14809,N_14891);
nor UO_1212 (O_1212,N_14943,N_14806);
xnor UO_1213 (O_1213,N_14983,N_14841);
nand UO_1214 (O_1214,N_14807,N_14857);
nand UO_1215 (O_1215,N_14945,N_14941);
and UO_1216 (O_1216,N_14975,N_14893);
or UO_1217 (O_1217,N_14918,N_14978);
nand UO_1218 (O_1218,N_14876,N_14827);
xor UO_1219 (O_1219,N_14916,N_14947);
xor UO_1220 (O_1220,N_14931,N_14890);
and UO_1221 (O_1221,N_14917,N_14994);
xor UO_1222 (O_1222,N_14881,N_14882);
or UO_1223 (O_1223,N_14927,N_14817);
nor UO_1224 (O_1224,N_14836,N_14869);
xor UO_1225 (O_1225,N_14852,N_14974);
nor UO_1226 (O_1226,N_14942,N_14868);
xor UO_1227 (O_1227,N_14841,N_14879);
nand UO_1228 (O_1228,N_14928,N_14895);
nand UO_1229 (O_1229,N_14862,N_14933);
and UO_1230 (O_1230,N_14971,N_14990);
and UO_1231 (O_1231,N_14820,N_14963);
or UO_1232 (O_1232,N_14904,N_14879);
or UO_1233 (O_1233,N_14991,N_14902);
nand UO_1234 (O_1234,N_14936,N_14880);
xor UO_1235 (O_1235,N_14912,N_14870);
nand UO_1236 (O_1236,N_14809,N_14856);
nor UO_1237 (O_1237,N_14805,N_14801);
nor UO_1238 (O_1238,N_14900,N_14996);
nand UO_1239 (O_1239,N_14972,N_14988);
and UO_1240 (O_1240,N_14830,N_14985);
nor UO_1241 (O_1241,N_14926,N_14908);
xor UO_1242 (O_1242,N_14958,N_14857);
nor UO_1243 (O_1243,N_14922,N_14852);
nor UO_1244 (O_1244,N_14826,N_14871);
nor UO_1245 (O_1245,N_14996,N_14912);
nor UO_1246 (O_1246,N_14810,N_14903);
xnor UO_1247 (O_1247,N_14896,N_14813);
nor UO_1248 (O_1248,N_14913,N_14815);
xnor UO_1249 (O_1249,N_14963,N_14930);
nand UO_1250 (O_1250,N_14976,N_14843);
xor UO_1251 (O_1251,N_14874,N_14802);
nand UO_1252 (O_1252,N_14851,N_14923);
nand UO_1253 (O_1253,N_14969,N_14851);
and UO_1254 (O_1254,N_14928,N_14869);
or UO_1255 (O_1255,N_14863,N_14808);
nor UO_1256 (O_1256,N_14885,N_14803);
nor UO_1257 (O_1257,N_14806,N_14981);
or UO_1258 (O_1258,N_14852,N_14868);
and UO_1259 (O_1259,N_14803,N_14974);
nor UO_1260 (O_1260,N_14851,N_14806);
nor UO_1261 (O_1261,N_14952,N_14916);
nand UO_1262 (O_1262,N_14940,N_14886);
and UO_1263 (O_1263,N_14926,N_14852);
or UO_1264 (O_1264,N_14943,N_14872);
xnor UO_1265 (O_1265,N_14843,N_14866);
and UO_1266 (O_1266,N_14989,N_14906);
or UO_1267 (O_1267,N_14886,N_14851);
nand UO_1268 (O_1268,N_14946,N_14940);
or UO_1269 (O_1269,N_14993,N_14857);
or UO_1270 (O_1270,N_14983,N_14813);
and UO_1271 (O_1271,N_14856,N_14811);
nand UO_1272 (O_1272,N_14977,N_14856);
nand UO_1273 (O_1273,N_14885,N_14977);
xor UO_1274 (O_1274,N_14809,N_14951);
nand UO_1275 (O_1275,N_14890,N_14906);
nand UO_1276 (O_1276,N_14861,N_14996);
and UO_1277 (O_1277,N_14970,N_14904);
or UO_1278 (O_1278,N_14869,N_14897);
xnor UO_1279 (O_1279,N_14999,N_14938);
nor UO_1280 (O_1280,N_14958,N_14837);
xor UO_1281 (O_1281,N_14938,N_14992);
or UO_1282 (O_1282,N_14954,N_14950);
and UO_1283 (O_1283,N_14833,N_14874);
and UO_1284 (O_1284,N_14934,N_14855);
xor UO_1285 (O_1285,N_14942,N_14936);
nand UO_1286 (O_1286,N_14852,N_14981);
nand UO_1287 (O_1287,N_14822,N_14857);
and UO_1288 (O_1288,N_14928,N_14999);
and UO_1289 (O_1289,N_14836,N_14967);
nand UO_1290 (O_1290,N_14981,N_14955);
nor UO_1291 (O_1291,N_14976,N_14983);
nor UO_1292 (O_1292,N_14979,N_14894);
xor UO_1293 (O_1293,N_14841,N_14949);
or UO_1294 (O_1294,N_14966,N_14833);
or UO_1295 (O_1295,N_14871,N_14882);
or UO_1296 (O_1296,N_14983,N_14890);
xor UO_1297 (O_1297,N_14953,N_14944);
and UO_1298 (O_1298,N_14830,N_14875);
nand UO_1299 (O_1299,N_14938,N_14802);
nor UO_1300 (O_1300,N_14854,N_14994);
xnor UO_1301 (O_1301,N_14932,N_14891);
and UO_1302 (O_1302,N_14822,N_14974);
and UO_1303 (O_1303,N_14984,N_14899);
xor UO_1304 (O_1304,N_14945,N_14966);
or UO_1305 (O_1305,N_14866,N_14800);
xnor UO_1306 (O_1306,N_14949,N_14845);
and UO_1307 (O_1307,N_14923,N_14972);
xor UO_1308 (O_1308,N_14820,N_14829);
nand UO_1309 (O_1309,N_14983,N_14960);
nand UO_1310 (O_1310,N_14841,N_14945);
or UO_1311 (O_1311,N_14878,N_14893);
or UO_1312 (O_1312,N_14828,N_14836);
and UO_1313 (O_1313,N_14999,N_14909);
xnor UO_1314 (O_1314,N_14974,N_14846);
nor UO_1315 (O_1315,N_14855,N_14886);
and UO_1316 (O_1316,N_14866,N_14892);
nand UO_1317 (O_1317,N_14919,N_14855);
xor UO_1318 (O_1318,N_14865,N_14923);
and UO_1319 (O_1319,N_14886,N_14896);
nand UO_1320 (O_1320,N_14960,N_14908);
nor UO_1321 (O_1321,N_14986,N_14959);
nor UO_1322 (O_1322,N_14946,N_14932);
nor UO_1323 (O_1323,N_14966,N_14846);
or UO_1324 (O_1324,N_14952,N_14850);
and UO_1325 (O_1325,N_14894,N_14883);
nor UO_1326 (O_1326,N_14903,N_14850);
or UO_1327 (O_1327,N_14965,N_14938);
xnor UO_1328 (O_1328,N_14936,N_14982);
or UO_1329 (O_1329,N_14820,N_14952);
xnor UO_1330 (O_1330,N_14888,N_14998);
or UO_1331 (O_1331,N_14834,N_14994);
nor UO_1332 (O_1332,N_14858,N_14855);
nor UO_1333 (O_1333,N_14985,N_14933);
or UO_1334 (O_1334,N_14915,N_14800);
nand UO_1335 (O_1335,N_14899,N_14964);
nor UO_1336 (O_1336,N_14892,N_14880);
nand UO_1337 (O_1337,N_14912,N_14814);
xor UO_1338 (O_1338,N_14988,N_14949);
xnor UO_1339 (O_1339,N_14851,N_14970);
nor UO_1340 (O_1340,N_14877,N_14850);
and UO_1341 (O_1341,N_14804,N_14888);
nor UO_1342 (O_1342,N_14939,N_14848);
and UO_1343 (O_1343,N_14921,N_14979);
or UO_1344 (O_1344,N_14956,N_14975);
nand UO_1345 (O_1345,N_14989,N_14979);
xor UO_1346 (O_1346,N_14835,N_14910);
nand UO_1347 (O_1347,N_14893,N_14817);
nand UO_1348 (O_1348,N_14813,N_14976);
and UO_1349 (O_1349,N_14900,N_14884);
xor UO_1350 (O_1350,N_14872,N_14930);
xor UO_1351 (O_1351,N_14893,N_14923);
or UO_1352 (O_1352,N_14886,N_14978);
xor UO_1353 (O_1353,N_14974,N_14975);
and UO_1354 (O_1354,N_14813,N_14907);
and UO_1355 (O_1355,N_14878,N_14867);
nor UO_1356 (O_1356,N_14903,N_14808);
xor UO_1357 (O_1357,N_14991,N_14924);
nand UO_1358 (O_1358,N_14816,N_14822);
or UO_1359 (O_1359,N_14839,N_14946);
xnor UO_1360 (O_1360,N_14839,N_14920);
xor UO_1361 (O_1361,N_14981,N_14864);
and UO_1362 (O_1362,N_14997,N_14958);
xor UO_1363 (O_1363,N_14809,N_14824);
nor UO_1364 (O_1364,N_14979,N_14972);
xor UO_1365 (O_1365,N_14991,N_14860);
and UO_1366 (O_1366,N_14910,N_14945);
or UO_1367 (O_1367,N_14987,N_14865);
nand UO_1368 (O_1368,N_14944,N_14854);
xor UO_1369 (O_1369,N_14816,N_14860);
nor UO_1370 (O_1370,N_14864,N_14975);
and UO_1371 (O_1371,N_14938,N_14909);
xor UO_1372 (O_1372,N_14999,N_14844);
nand UO_1373 (O_1373,N_14828,N_14834);
nand UO_1374 (O_1374,N_14863,N_14913);
xor UO_1375 (O_1375,N_14947,N_14839);
xor UO_1376 (O_1376,N_14900,N_14853);
xor UO_1377 (O_1377,N_14970,N_14983);
or UO_1378 (O_1378,N_14997,N_14876);
or UO_1379 (O_1379,N_14800,N_14969);
nand UO_1380 (O_1380,N_14935,N_14995);
nor UO_1381 (O_1381,N_14880,N_14877);
or UO_1382 (O_1382,N_14994,N_14966);
xnor UO_1383 (O_1383,N_14877,N_14957);
and UO_1384 (O_1384,N_14998,N_14981);
nand UO_1385 (O_1385,N_14881,N_14937);
nor UO_1386 (O_1386,N_14835,N_14920);
nand UO_1387 (O_1387,N_14871,N_14878);
nand UO_1388 (O_1388,N_14936,N_14934);
xor UO_1389 (O_1389,N_14866,N_14889);
or UO_1390 (O_1390,N_14864,N_14805);
nor UO_1391 (O_1391,N_14875,N_14863);
and UO_1392 (O_1392,N_14994,N_14848);
xnor UO_1393 (O_1393,N_14803,N_14988);
nor UO_1394 (O_1394,N_14899,N_14998);
or UO_1395 (O_1395,N_14822,N_14836);
or UO_1396 (O_1396,N_14840,N_14959);
and UO_1397 (O_1397,N_14926,N_14964);
and UO_1398 (O_1398,N_14866,N_14847);
nor UO_1399 (O_1399,N_14832,N_14805);
and UO_1400 (O_1400,N_14927,N_14884);
and UO_1401 (O_1401,N_14921,N_14842);
nand UO_1402 (O_1402,N_14871,N_14887);
nor UO_1403 (O_1403,N_14840,N_14950);
nand UO_1404 (O_1404,N_14946,N_14831);
nor UO_1405 (O_1405,N_14911,N_14818);
and UO_1406 (O_1406,N_14854,N_14900);
or UO_1407 (O_1407,N_14802,N_14963);
xor UO_1408 (O_1408,N_14983,N_14837);
xor UO_1409 (O_1409,N_14843,N_14918);
and UO_1410 (O_1410,N_14982,N_14839);
and UO_1411 (O_1411,N_14868,N_14862);
xnor UO_1412 (O_1412,N_14858,N_14897);
or UO_1413 (O_1413,N_14936,N_14902);
nor UO_1414 (O_1414,N_14856,N_14955);
nand UO_1415 (O_1415,N_14981,N_14878);
nor UO_1416 (O_1416,N_14900,N_14987);
nand UO_1417 (O_1417,N_14873,N_14851);
or UO_1418 (O_1418,N_14994,N_14800);
nor UO_1419 (O_1419,N_14929,N_14868);
or UO_1420 (O_1420,N_14810,N_14895);
nand UO_1421 (O_1421,N_14845,N_14989);
nor UO_1422 (O_1422,N_14886,N_14988);
nor UO_1423 (O_1423,N_14894,N_14846);
nor UO_1424 (O_1424,N_14814,N_14849);
or UO_1425 (O_1425,N_14893,N_14805);
nor UO_1426 (O_1426,N_14954,N_14818);
or UO_1427 (O_1427,N_14905,N_14906);
nor UO_1428 (O_1428,N_14891,N_14921);
nor UO_1429 (O_1429,N_14930,N_14934);
xor UO_1430 (O_1430,N_14870,N_14841);
xnor UO_1431 (O_1431,N_14962,N_14902);
or UO_1432 (O_1432,N_14992,N_14921);
nor UO_1433 (O_1433,N_14897,N_14883);
xnor UO_1434 (O_1434,N_14986,N_14939);
or UO_1435 (O_1435,N_14929,N_14869);
or UO_1436 (O_1436,N_14858,N_14825);
and UO_1437 (O_1437,N_14908,N_14869);
nand UO_1438 (O_1438,N_14979,N_14802);
and UO_1439 (O_1439,N_14865,N_14855);
nand UO_1440 (O_1440,N_14849,N_14829);
and UO_1441 (O_1441,N_14958,N_14979);
and UO_1442 (O_1442,N_14892,N_14962);
nor UO_1443 (O_1443,N_14948,N_14971);
xnor UO_1444 (O_1444,N_14888,N_14841);
or UO_1445 (O_1445,N_14873,N_14922);
xor UO_1446 (O_1446,N_14945,N_14817);
or UO_1447 (O_1447,N_14974,N_14837);
or UO_1448 (O_1448,N_14801,N_14883);
nand UO_1449 (O_1449,N_14870,N_14941);
nor UO_1450 (O_1450,N_14869,N_14915);
xnor UO_1451 (O_1451,N_14969,N_14937);
or UO_1452 (O_1452,N_14975,N_14913);
and UO_1453 (O_1453,N_14971,N_14895);
nand UO_1454 (O_1454,N_14802,N_14919);
or UO_1455 (O_1455,N_14861,N_14842);
nor UO_1456 (O_1456,N_14924,N_14962);
xor UO_1457 (O_1457,N_14811,N_14922);
or UO_1458 (O_1458,N_14835,N_14965);
or UO_1459 (O_1459,N_14947,N_14870);
or UO_1460 (O_1460,N_14975,N_14909);
nand UO_1461 (O_1461,N_14822,N_14891);
nand UO_1462 (O_1462,N_14846,N_14870);
nor UO_1463 (O_1463,N_14994,N_14912);
nor UO_1464 (O_1464,N_14832,N_14984);
or UO_1465 (O_1465,N_14993,N_14951);
and UO_1466 (O_1466,N_14984,N_14836);
nand UO_1467 (O_1467,N_14886,N_14989);
nand UO_1468 (O_1468,N_14869,N_14973);
xnor UO_1469 (O_1469,N_14844,N_14953);
xor UO_1470 (O_1470,N_14889,N_14802);
nor UO_1471 (O_1471,N_14891,N_14853);
xnor UO_1472 (O_1472,N_14907,N_14949);
xnor UO_1473 (O_1473,N_14898,N_14994);
nor UO_1474 (O_1474,N_14999,N_14943);
and UO_1475 (O_1475,N_14812,N_14926);
and UO_1476 (O_1476,N_14901,N_14830);
nor UO_1477 (O_1477,N_14959,N_14952);
and UO_1478 (O_1478,N_14860,N_14878);
nand UO_1479 (O_1479,N_14820,N_14992);
xor UO_1480 (O_1480,N_14826,N_14945);
or UO_1481 (O_1481,N_14831,N_14814);
xor UO_1482 (O_1482,N_14937,N_14878);
nand UO_1483 (O_1483,N_14925,N_14898);
or UO_1484 (O_1484,N_14807,N_14835);
nor UO_1485 (O_1485,N_14942,N_14940);
and UO_1486 (O_1486,N_14964,N_14970);
nand UO_1487 (O_1487,N_14852,N_14867);
and UO_1488 (O_1488,N_14927,N_14836);
xnor UO_1489 (O_1489,N_14824,N_14844);
xor UO_1490 (O_1490,N_14946,N_14813);
nor UO_1491 (O_1491,N_14972,N_14805);
nor UO_1492 (O_1492,N_14851,N_14811);
or UO_1493 (O_1493,N_14979,N_14926);
xor UO_1494 (O_1494,N_14967,N_14968);
xor UO_1495 (O_1495,N_14808,N_14921);
nand UO_1496 (O_1496,N_14933,N_14805);
nand UO_1497 (O_1497,N_14967,N_14871);
xnor UO_1498 (O_1498,N_14801,N_14876);
xnor UO_1499 (O_1499,N_14877,N_14878);
xor UO_1500 (O_1500,N_14997,N_14819);
and UO_1501 (O_1501,N_14821,N_14988);
nor UO_1502 (O_1502,N_14957,N_14907);
and UO_1503 (O_1503,N_14807,N_14801);
or UO_1504 (O_1504,N_14978,N_14894);
xor UO_1505 (O_1505,N_14862,N_14951);
and UO_1506 (O_1506,N_14858,N_14962);
xnor UO_1507 (O_1507,N_14964,N_14946);
nand UO_1508 (O_1508,N_14908,N_14916);
and UO_1509 (O_1509,N_14855,N_14859);
and UO_1510 (O_1510,N_14932,N_14901);
nand UO_1511 (O_1511,N_14809,N_14986);
and UO_1512 (O_1512,N_14988,N_14876);
or UO_1513 (O_1513,N_14953,N_14912);
xnor UO_1514 (O_1514,N_14983,N_14951);
and UO_1515 (O_1515,N_14908,N_14862);
xor UO_1516 (O_1516,N_14995,N_14879);
or UO_1517 (O_1517,N_14984,N_14847);
and UO_1518 (O_1518,N_14993,N_14966);
and UO_1519 (O_1519,N_14939,N_14918);
xor UO_1520 (O_1520,N_14937,N_14854);
nand UO_1521 (O_1521,N_14994,N_14845);
and UO_1522 (O_1522,N_14832,N_14819);
xor UO_1523 (O_1523,N_14940,N_14962);
and UO_1524 (O_1524,N_14973,N_14948);
nor UO_1525 (O_1525,N_14995,N_14982);
xor UO_1526 (O_1526,N_14859,N_14910);
nor UO_1527 (O_1527,N_14990,N_14996);
or UO_1528 (O_1528,N_14860,N_14894);
or UO_1529 (O_1529,N_14922,N_14904);
and UO_1530 (O_1530,N_14832,N_14938);
xor UO_1531 (O_1531,N_14867,N_14973);
or UO_1532 (O_1532,N_14852,N_14915);
and UO_1533 (O_1533,N_14854,N_14901);
nand UO_1534 (O_1534,N_14856,N_14996);
and UO_1535 (O_1535,N_14976,N_14837);
nor UO_1536 (O_1536,N_14839,N_14807);
xor UO_1537 (O_1537,N_14996,N_14931);
and UO_1538 (O_1538,N_14844,N_14887);
and UO_1539 (O_1539,N_14835,N_14942);
or UO_1540 (O_1540,N_14866,N_14985);
or UO_1541 (O_1541,N_14970,N_14885);
nand UO_1542 (O_1542,N_14833,N_14879);
xor UO_1543 (O_1543,N_14950,N_14879);
or UO_1544 (O_1544,N_14877,N_14996);
nor UO_1545 (O_1545,N_14960,N_14993);
nand UO_1546 (O_1546,N_14912,N_14864);
nor UO_1547 (O_1547,N_14966,N_14919);
xor UO_1548 (O_1548,N_14836,N_14808);
xnor UO_1549 (O_1549,N_14914,N_14985);
and UO_1550 (O_1550,N_14971,N_14883);
and UO_1551 (O_1551,N_14949,N_14971);
nand UO_1552 (O_1552,N_14873,N_14844);
nor UO_1553 (O_1553,N_14844,N_14820);
and UO_1554 (O_1554,N_14944,N_14954);
nor UO_1555 (O_1555,N_14831,N_14830);
nor UO_1556 (O_1556,N_14930,N_14863);
nor UO_1557 (O_1557,N_14870,N_14984);
xnor UO_1558 (O_1558,N_14903,N_14998);
or UO_1559 (O_1559,N_14931,N_14964);
nor UO_1560 (O_1560,N_14897,N_14988);
nor UO_1561 (O_1561,N_14915,N_14842);
and UO_1562 (O_1562,N_14976,N_14966);
and UO_1563 (O_1563,N_14973,N_14939);
nand UO_1564 (O_1564,N_14888,N_14853);
or UO_1565 (O_1565,N_14879,N_14911);
xnor UO_1566 (O_1566,N_14873,N_14956);
and UO_1567 (O_1567,N_14911,N_14972);
nor UO_1568 (O_1568,N_14882,N_14907);
nor UO_1569 (O_1569,N_14898,N_14986);
xnor UO_1570 (O_1570,N_14922,N_14846);
or UO_1571 (O_1571,N_14970,N_14941);
and UO_1572 (O_1572,N_14883,N_14992);
or UO_1573 (O_1573,N_14991,N_14896);
nand UO_1574 (O_1574,N_14951,N_14955);
nor UO_1575 (O_1575,N_14873,N_14930);
xnor UO_1576 (O_1576,N_14942,N_14975);
and UO_1577 (O_1577,N_14888,N_14821);
or UO_1578 (O_1578,N_14863,N_14972);
nor UO_1579 (O_1579,N_14806,N_14915);
xnor UO_1580 (O_1580,N_14990,N_14948);
xnor UO_1581 (O_1581,N_14960,N_14875);
nor UO_1582 (O_1582,N_14878,N_14910);
and UO_1583 (O_1583,N_14840,N_14863);
and UO_1584 (O_1584,N_14970,N_14940);
or UO_1585 (O_1585,N_14808,N_14966);
nand UO_1586 (O_1586,N_14982,N_14996);
nand UO_1587 (O_1587,N_14927,N_14845);
nor UO_1588 (O_1588,N_14845,N_14884);
nand UO_1589 (O_1589,N_14881,N_14993);
and UO_1590 (O_1590,N_14861,N_14935);
and UO_1591 (O_1591,N_14920,N_14983);
xnor UO_1592 (O_1592,N_14863,N_14918);
nor UO_1593 (O_1593,N_14867,N_14956);
xor UO_1594 (O_1594,N_14895,N_14934);
nand UO_1595 (O_1595,N_14868,N_14943);
nand UO_1596 (O_1596,N_14999,N_14973);
xnor UO_1597 (O_1597,N_14874,N_14986);
and UO_1598 (O_1598,N_14928,N_14973);
nand UO_1599 (O_1599,N_14961,N_14941);
nand UO_1600 (O_1600,N_14855,N_14929);
xor UO_1601 (O_1601,N_14912,N_14957);
and UO_1602 (O_1602,N_14818,N_14981);
xor UO_1603 (O_1603,N_14832,N_14943);
nand UO_1604 (O_1604,N_14806,N_14884);
nand UO_1605 (O_1605,N_14856,N_14891);
xor UO_1606 (O_1606,N_14829,N_14847);
nor UO_1607 (O_1607,N_14895,N_14884);
or UO_1608 (O_1608,N_14858,N_14860);
nand UO_1609 (O_1609,N_14986,N_14895);
or UO_1610 (O_1610,N_14854,N_14825);
and UO_1611 (O_1611,N_14974,N_14906);
nor UO_1612 (O_1612,N_14816,N_14923);
or UO_1613 (O_1613,N_14965,N_14829);
nand UO_1614 (O_1614,N_14992,N_14922);
xor UO_1615 (O_1615,N_14958,N_14891);
nand UO_1616 (O_1616,N_14833,N_14937);
or UO_1617 (O_1617,N_14876,N_14855);
nand UO_1618 (O_1618,N_14838,N_14875);
or UO_1619 (O_1619,N_14851,N_14989);
nor UO_1620 (O_1620,N_14894,N_14863);
nor UO_1621 (O_1621,N_14950,N_14876);
xor UO_1622 (O_1622,N_14830,N_14969);
nor UO_1623 (O_1623,N_14896,N_14825);
xor UO_1624 (O_1624,N_14954,N_14921);
and UO_1625 (O_1625,N_14820,N_14847);
nand UO_1626 (O_1626,N_14844,N_14909);
nand UO_1627 (O_1627,N_14896,N_14936);
nor UO_1628 (O_1628,N_14942,N_14923);
xnor UO_1629 (O_1629,N_14817,N_14837);
nand UO_1630 (O_1630,N_14980,N_14924);
nor UO_1631 (O_1631,N_14899,N_14823);
nor UO_1632 (O_1632,N_14912,N_14820);
nand UO_1633 (O_1633,N_14912,N_14977);
xor UO_1634 (O_1634,N_14838,N_14836);
xnor UO_1635 (O_1635,N_14916,N_14821);
nor UO_1636 (O_1636,N_14992,N_14878);
xor UO_1637 (O_1637,N_14968,N_14932);
and UO_1638 (O_1638,N_14907,N_14875);
nor UO_1639 (O_1639,N_14840,N_14841);
or UO_1640 (O_1640,N_14917,N_14952);
and UO_1641 (O_1641,N_14960,N_14868);
xnor UO_1642 (O_1642,N_14943,N_14928);
and UO_1643 (O_1643,N_14987,N_14818);
or UO_1644 (O_1644,N_14816,N_14986);
and UO_1645 (O_1645,N_14905,N_14890);
xnor UO_1646 (O_1646,N_14946,N_14896);
nor UO_1647 (O_1647,N_14918,N_14951);
nand UO_1648 (O_1648,N_14923,N_14855);
nor UO_1649 (O_1649,N_14998,N_14882);
xnor UO_1650 (O_1650,N_14961,N_14846);
or UO_1651 (O_1651,N_14998,N_14957);
nand UO_1652 (O_1652,N_14950,N_14941);
xnor UO_1653 (O_1653,N_14844,N_14997);
nor UO_1654 (O_1654,N_14806,N_14809);
or UO_1655 (O_1655,N_14947,N_14920);
xor UO_1656 (O_1656,N_14892,N_14852);
nand UO_1657 (O_1657,N_14820,N_14838);
nor UO_1658 (O_1658,N_14856,N_14873);
nand UO_1659 (O_1659,N_14985,N_14867);
or UO_1660 (O_1660,N_14810,N_14991);
and UO_1661 (O_1661,N_14819,N_14977);
or UO_1662 (O_1662,N_14836,N_14814);
nand UO_1663 (O_1663,N_14975,N_14992);
nor UO_1664 (O_1664,N_14905,N_14855);
or UO_1665 (O_1665,N_14861,N_14883);
or UO_1666 (O_1666,N_14909,N_14885);
xor UO_1667 (O_1667,N_14919,N_14951);
and UO_1668 (O_1668,N_14855,N_14909);
nand UO_1669 (O_1669,N_14829,N_14869);
and UO_1670 (O_1670,N_14817,N_14932);
nor UO_1671 (O_1671,N_14816,N_14911);
nand UO_1672 (O_1672,N_14943,N_14981);
nor UO_1673 (O_1673,N_14882,N_14945);
nand UO_1674 (O_1674,N_14984,N_14879);
and UO_1675 (O_1675,N_14899,N_14970);
nor UO_1676 (O_1676,N_14817,N_14878);
and UO_1677 (O_1677,N_14924,N_14929);
and UO_1678 (O_1678,N_14958,N_14901);
nor UO_1679 (O_1679,N_14901,N_14914);
nand UO_1680 (O_1680,N_14941,N_14922);
or UO_1681 (O_1681,N_14871,N_14901);
nor UO_1682 (O_1682,N_14957,N_14982);
nor UO_1683 (O_1683,N_14940,N_14813);
xor UO_1684 (O_1684,N_14812,N_14962);
nor UO_1685 (O_1685,N_14820,N_14879);
nand UO_1686 (O_1686,N_14833,N_14972);
and UO_1687 (O_1687,N_14849,N_14968);
xnor UO_1688 (O_1688,N_14965,N_14937);
xor UO_1689 (O_1689,N_14884,N_14857);
or UO_1690 (O_1690,N_14843,N_14956);
and UO_1691 (O_1691,N_14823,N_14885);
or UO_1692 (O_1692,N_14914,N_14882);
nor UO_1693 (O_1693,N_14870,N_14875);
or UO_1694 (O_1694,N_14801,N_14831);
xor UO_1695 (O_1695,N_14992,N_14910);
nor UO_1696 (O_1696,N_14988,N_14891);
nand UO_1697 (O_1697,N_14940,N_14943);
xor UO_1698 (O_1698,N_14865,N_14832);
nor UO_1699 (O_1699,N_14943,N_14889);
xor UO_1700 (O_1700,N_14947,N_14987);
nand UO_1701 (O_1701,N_14845,N_14900);
nor UO_1702 (O_1702,N_14874,N_14856);
and UO_1703 (O_1703,N_14829,N_14916);
nor UO_1704 (O_1704,N_14852,N_14800);
or UO_1705 (O_1705,N_14943,N_14810);
and UO_1706 (O_1706,N_14853,N_14816);
or UO_1707 (O_1707,N_14990,N_14879);
xnor UO_1708 (O_1708,N_14903,N_14896);
nor UO_1709 (O_1709,N_14902,N_14879);
nor UO_1710 (O_1710,N_14811,N_14870);
or UO_1711 (O_1711,N_14906,N_14803);
nor UO_1712 (O_1712,N_14951,N_14988);
nor UO_1713 (O_1713,N_14897,N_14973);
nor UO_1714 (O_1714,N_14984,N_14863);
xnor UO_1715 (O_1715,N_14954,N_14826);
nand UO_1716 (O_1716,N_14970,N_14844);
nor UO_1717 (O_1717,N_14948,N_14878);
or UO_1718 (O_1718,N_14818,N_14821);
nor UO_1719 (O_1719,N_14962,N_14990);
nand UO_1720 (O_1720,N_14904,N_14983);
nor UO_1721 (O_1721,N_14990,N_14848);
nand UO_1722 (O_1722,N_14848,N_14819);
xnor UO_1723 (O_1723,N_14896,N_14994);
xor UO_1724 (O_1724,N_14949,N_14889);
and UO_1725 (O_1725,N_14871,N_14813);
and UO_1726 (O_1726,N_14996,N_14929);
and UO_1727 (O_1727,N_14950,N_14800);
and UO_1728 (O_1728,N_14992,N_14880);
xor UO_1729 (O_1729,N_14944,N_14895);
nor UO_1730 (O_1730,N_14873,N_14882);
and UO_1731 (O_1731,N_14881,N_14868);
nor UO_1732 (O_1732,N_14959,N_14827);
nand UO_1733 (O_1733,N_14964,N_14869);
and UO_1734 (O_1734,N_14936,N_14882);
and UO_1735 (O_1735,N_14906,N_14830);
xor UO_1736 (O_1736,N_14925,N_14811);
or UO_1737 (O_1737,N_14919,N_14989);
or UO_1738 (O_1738,N_14823,N_14825);
xnor UO_1739 (O_1739,N_14965,N_14922);
nand UO_1740 (O_1740,N_14832,N_14815);
nand UO_1741 (O_1741,N_14902,N_14819);
or UO_1742 (O_1742,N_14813,N_14936);
nor UO_1743 (O_1743,N_14858,N_14850);
and UO_1744 (O_1744,N_14898,N_14818);
nor UO_1745 (O_1745,N_14933,N_14835);
nand UO_1746 (O_1746,N_14823,N_14987);
and UO_1747 (O_1747,N_14881,N_14972);
nor UO_1748 (O_1748,N_14948,N_14938);
nand UO_1749 (O_1749,N_14830,N_14943);
nor UO_1750 (O_1750,N_14962,N_14802);
xor UO_1751 (O_1751,N_14988,N_14878);
or UO_1752 (O_1752,N_14835,N_14991);
xnor UO_1753 (O_1753,N_14868,N_14998);
and UO_1754 (O_1754,N_14949,N_14835);
nand UO_1755 (O_1755,N_14978,N_14802);
nor UO_1756 (O_1756,N_14887,N_14856);
nand UO_1757 (O_1757,N_14980,N_14856);
and UO_1758 (O_1758,N_14892,N_14831);
nor UO_1759 (O_1759,N_14957,N_14928);
and UO_1760 (O_1760,N_14981,N_14869);
nor UO_1761 (O_1761,N_14962,N_14972);
nand UO_1762 (O_1762,N_14954,N_14866);
or UO_1763 (O_1763,N_14916,N_14813);
xor UO_1764 (O_1764,N_14844,N_14801);
nand UO_1765 (O_1765,N_14865,N_14908);
xor UO_1766 (O_1766,N_14811,N_14877);
and UO_1767 (O_1767,N_14968,N_14808);
xor UO_1768 (O_1768,N_14920,N_14882);
or UO_1769 (O_1769,N_14867,N_14843);
and UO_1770 (O_1770,N_14934,N_14882);
xor UO_1771 (O_1771,N_14869,N_14937);
xor UO_1772 (O_1772,N_14976,N_14891);
nand UO_1773 (O_1773,N_14802,N_14866);
nor UO_1774 (O_1774,N_14841,N_14954);
and UO_1775 (O_1775,N_14826,N_14957);
xnor UO_1776 (O_1776,N_14932,N_14807);
nor UO_1777 (O_1777,N_14811,N_14863);
and UO_1778 (O_1778,N_14848,N_14989);
nand UO_1779 (O_1779,N_14936,N_14861);
and UO_1780 (O_1780,N_14824,N_14830);
or UO_1781 (O_1781,N_14934,N_14909);
or UO_1782 (O_1782,N_14828,N_14944);
and UO_1783 (O_1783,N_14858,N_14944);
and UO_1784 (O_1784,N_14927,N_14809);
xnor UO_1785 (O_1785,N_14971,N_14978);
nand UO_1786 (O_1786,N_14932,N_14825);
nand UO_1787 (O_1787,N_14941,N_14894);
or UO_1788 (O_1788,N_14949,N_14863);
or UO_1789 (O_1789,N_14958,N_14940);
and UO_1790 (O_1790,N_14982,N_14947);
nand UO_1791 (O_1791,N_14929,N_14841);
and UO_1792 (O_1792,N_14912,N_14844);
nor UO_1793 (O_1793,N_14981,N_14874);
nor UO_1794 (O_1794,N_14862,N_14854);
xnor UO_1795 (O_1795,N_14949,N_14851);
nor UO_1796 (O_1796,N_14866,N_14950);
nand UO_1797 (O_1797,N_14858,N_14921);
xnor UO_1798 (O_1798,N_14937,N_14802);
nor UO_1799 (O_1799,N_14924,N_14859);
xor UO_1800 (O_1800,N_14846,N_14953);
xor UO_1801 (O_1801,N_14979,N_14940);
and UO_1802 (O_1802,N_14866,N_14831);
and UO_1803 (O_1803,N_14829,N_14852);
xnor UO_1804 (O_1804,N_14927,N_14993);
and UO_1805 (O_1805,N_14818,N_14972);
nor UO_1806 (O_1806,N_14950,N_14945);
and UO_1807 (O_1807,N_14903,N_14973);
or UO_1808 (O_1808,N_14932,N_14811);
nand UO_1809 (O_1809,N_14947,N_14990);
nand UO_1810 (O_1810,N_14879,N_14983);
nor UO_1811 (O_1811,N_14935,N_14911);
nor UO_1812 (O_1812,N_14862,N_14912);
or UO_1813 (O_1813,N_14969,N_14861);
nor UO_1814 (O_1814,N_14908,N_14924);
nor UO_1815 (O_1815,N_14944,N_14825);
xor UO_1816 (O_1816,N_14920,N_14809);
nor UO_1817 (O_1817,N_14885,N_14818);
xor UO_1818 (O_1818,N_14992,N_14857);
xnor UO_1819 (O_1819,N_14957,N_14848);
nor UO_1820 (O_1820,N_14908,N_14843);
xor UO_1821 (O_1821,N_14969,N_14882);
and UO_1822 (O_1822,N_14939,N_14964);
nand UO_1823 (O_1823,N_14815,N_14835);
nor UO_1824 (O_1824,N_14814,N_14818);
and UO_1825 (O_1825,N_14848,N_14918);
and UO_1826 (O_1826,N_14899,N_14882);
nor UO_1827 (O_1827,N_14804,N_14902);
xor UO_1828 (O_1828,N_14963,N_14842);
nor UO_1829 (O_1829,N_14887,N_14997);
nor UO_1830 (O_1830,N_14885,N_14842);
or UO_1831 (O_1831,N_14816,N_14908);
nor UO_1832 (O_1832,N_14928,N_14994);
nand UO_1833 (O_1833,N_14835,N_14921);
and UO_1834 (O_1834,N_14989,N_14883);
nand UO_1835 (O_1835,N_14922,N_14955);
nor UO_1836 (O_1836,N_14809,N_14804);
nor UO_1837 (O_1837,N_14915,N_14956);
and UO_1838 (O_1838,N_14900,N_14818);
nand UO_1839 (O_1839,N_14976,N_14915);
or UO_1840 (O_1840,N_14807,N_14880);
nor UO_1841 (O_1841,N_14846,N_14889);
or UO_1842 (O_1842,N_14881,N_14975);
and UO_1843 (O_1843,N_14835,N_14898);
xnor UO_1844 (O_1844,N_14954,N_14925);
nand UO_1845 (O_1845,N_14864,N_14859);
or UO_1846 (O_1846,N_14906,N_14844);
and UO_1847 (O_1847,N_14907,N_14993);
or UO_1848 (O_1848,N_14960,N_14816);
nand UO_1849 (O_1849,N_14897,N_14963);
xor UO_1850 (O_1850,N_14823,N_14851);
nor UO_1851 (O_1851,N_14850,N_14801);
nand UO_1852 (O_1852,N_14835,N_14896);
nor UO_1853 (O_1853,N_14955,N_14950);
or UO_1854 (O_1854,N_14917,N_14857);
nor UO_1855 (O_1855,N_14954,N_14990);
nand UO_1856 (O_1856,N_14804,N_14947);
nand UO_1857 (O_1857,N_14959,N_14997);
or UO_1858 (O_1858,N_14815,N_14925);
nand UO_1859 (O_1859,N_14913,N_14851);
nor UO_1860 (O_1860,N_14893,N_14907);
nand UO_1861 (O_1861,N_14904,N_14915);
or UO_1862 (O_1862,N_14937,N_14950);
nor UO_1863 (O_1863,N_14945,N_14836);
and UO_1864 (O_1864,N_14920,N_14824);
xnor UO_1865 (O_1865,N_14871,N_14862);
or UO_1866 (O_1866,N_14905,N_14920);
xnor UO_1867 (O_1867,N_14870,N_14884);
xnor UO_1868 (O_1868,N_14868,N_14907);
xor UO_1869 (O_1869,N_14888,N_14936);
and UO_1870 (O_1870,N_14867,N_14862);
and UO_1871 (O_1871,N_14800,N_14883);
nor UO_1872 (O_1872,N_14940,N_14867);
and UO_1873 (O_1873,N_14892,N_14915);
xnor UO_1874 (O_1874,N_14935,N_14875);
xor UO_1875 (O_1875,N_14840,N_14886);
nand UO_1876 (O_1876,N_14843,N_14838);
nor UO_1877 (O_1877,N_14839,N_14874);
nand UO_1878 (O_1878,N_14911,N_14994);
nor UO_1879 (O_1879,N_14896,N_14841);
or UO_1880 (O_1880,N_14942,N_14857);
nor UO_1881 (O_1881,N_14943,N_14859);
nand UO_1882 (O_1882,N_14950,N_14933);
xnor UO_1883 (O_1883,N_14887,N_14878);
and UO_1884 (O_1884,N_14948,N_14968);
and UO_1885 (O_1885,N_14977,N_14979);
xor UO_1886 (O_1886,N_14895,N_14839);
xnor UO_1887 (O_1887,N_14947,N_14988);
nor UO_1888 (O_1888,N_14808,N_14894);
xnor UO_1889 (O_1889,N_14961,N_14980);
nand UO_1890 (O_1890,N_14908,N_14845);
or UO_1891 (O_1891,N_14972,N_14801);
nor UO_1892 (O_1892,N_14971,N_14888);
xor UO_1893 (O_1893,N_14803,N_14955);
nand UO_1894 (O_1894,N_14827,N_14898);
nor UO_1895 (O_1895,N_14881,N_14805);
and UO_1896 (O_1896,N_14818,N_14978);
nand UO_1897 (O_1897,N_14823,N_14973);
xor UO_1898 (O_1898,N_14911,N_14829);
xor UO_1899 (O_1899,N_14849,N_14899);
nand UO_1900 (O_1900,N_14920,N_14975);
or UO_1901 (O_1901,N_14902,N_14952);
or UO_1902 (O_1902,N_14952,N_14991);
or UO_1903 (O_1903,N_14918,N_14911);
or UO_1904 (O_1904,N_14818,N_14871);
nand UO_1905 (O_1905,N_14856,N_14903);
and UO_1906 (O_1906,N_14871,N_14824);
xor UO_1907 (O_1907,N_14964,N_14945);
nor UO_1908 (O_1908,N_14829,N_14957);
xor UO_1909 (O_1909,N_14828,N_14827);
or UO_1910 (O_1910,N_14831,N_14878);
xor UO_1911 (O_1911,N_14833,N_14822);
nand UO_1912 (O_1912,N_14849,N_14819);
or UO_1913 (O_1913,N_14832,N_14836);
xnor UO_1914 (O_1914,N_14929,N_14838);
nor UO_1915 (O_1915,N_14934,N_14947);
nand UO_1916 (O_1916,N_14920,N_14911);
and UO_1917 (O_1917,N_14906,N_14819);
nor UO_1918 (O_1918,N_14824,N_14882);
nor UO_1919 (O_1919,N_14923,N_14820);
nand UO_1920 (O_1920,N_14820,N_14817);
xor UO_1921 (O_1921,N_14842,N_14908);
xor UO_1922 (O_1922,N_14852,N_14918);
nand UO_1923 (O_1923,N_14995,N_14885);
nand UO_1924 (O_1924,N_14888,N_14822);
or UO_1925 (O_1925,N_14917,N_14937);
or UO_1926 (O_1926,N_14878,N_14998);
and UO_1927 (O_1927,N_14832,N_14927);
and UO_1928 (O_1928,N_14953,N_14840);
or UO_1929 (O_1929,N_14913,N_14954);
xnor UO_1930 (O_1930,N_14810,N_14968);
nand UO_1931 (O_1931,N_14831,N_14984);
nor UO_1932 (O_1932,N_14929,N_14802);
nand UO_1933 (O_1933,N_14800,N_14917);
and UO_1934 (O_1934,N_14987,N_14917);
xor UO_1935 (O_1935,N_14885,N_14822);
nor UO_1936 (O_1936,N_14911,N_14878);
or UO_1937 (O_1937,N_14926,N_14996);
nand UO_1938 (O_1938,N_14955,N_14816);
nor UO_1939 (O_1939,N_14846,N_14898);
and UO_1940 (O_1940,N_14979,N_14883);
nand UO_1941 (O_1941,N_14973,N_14909);
and UO_1942 (O_1942,N_14906,N_14851);
xnor UO_1943 (O_1943,N_14832,N_14994);
or UO_1944 (O_1944,N_14939,N_14943);
and UO_1945 (O_1945,N_14924,N_14838);
nand UO_1946 (O_1946,N_14988,N_14990);
xor UO_1947 (O_1947,N_14940,N_14819);
xor UO_1948 (O_1948,N_14964,N_14971);
and UO_1949 (O_1949,N_14832,N_14830);
nor UO_1950 (O_1950,N_14995,N_14992);
nand UO_1951 (O_1951,N_14941,N_14966);
nor UO_1952 (O_1952,N_14803,N_14808);
or UO_1953 (O_1953,N_14990,N_14865);
and UO_1954 (O_1954,N_14934,N_14941);
nand UO_1955 (O_1955,N_14927,N_14855);
nor UO_1956 (O_1956,N_14986,N_14812);
nand UO_1957 (O_1957,N_14961,N_14931);
or UO_1958 (O_1958,N_14831,N_14886);
nand UO_1959 (O_1959,N_14987,N_14857);
nor UO_1960 (O_1960,N_14988,N_14808);
nor UO_1961 (O_1961,N_14944,N_14887);
and UO_1962 (O_1962,N_14995,N_14968);
nand UO_1963 (O_1963,N_14972,N_14910);
or UO_1964 (O_1964,N_14890,N_14855);
nor UO_1965 (O_1965,N_14977,N_14835);
xnor UO_1966 (O_1966,N_14911,N_14955);
or UO_1967 (O_1967,N_14942,N_14947);
nor UO_1968 (O_1968,N_14971,N_14889);
or UO_1969 (O_1969,N_14951,N_14840);
nor UO_1970 (O_1970,N_14814,N_14926);
nor UO_1971 (O_1971,N_14941,N_14812);
and UO_1972 (O_1972,N_14832,N_14888);
nand UO_1973 (O_1973,N_14896,N_14957);
nor UO_1974 (O_1974,N_14934,N_14974);
xnor UO_1975 (O_1975,N_14984,N_14944);
and UO_1976 (O_1976,N_14850,N_14829);
xor UO_1977 (O_1977,N_14871,N_14817);
and UO_1978 (O_1978,N_14974,N_14987);
xnor UO_1979 (O_1979,N_14847,N_14865);
nand UO_1980 (O_1980,N_14952,N_14813);
and UO_1981 (O_1981,N_14873,N_14948);
or UO_1982 (O_1982,N_14835,N_14908);
and UO_1983 (O_1983,N_14963,N_14896);
nand UO_1984 (O_1984,N_14996,N_14995);
xnor UO_1985 (O_1985,N_14956,N_14994);
or UO_1986 (O_1986,N_14939,N_14854);
and UO_1987 (O_1987,N_14983,N_14899);
and UO_1988 (O_1988,N_14867,N_14806);
or UO_1989 (O_1989,N_14903,N_14826);
or UO_1990 (O_1990,N_14831,N_14867);
xnor UO_1991 (O_1991,N_14968,N_14840);
nor UO_1992 (O_1992,N_14932,N_14907);
xnor UO_1993 (O_1993,N_14819,N_14934);
and UO_1994 (O_1994,N_14824,N_14912);
nor UO_1995 (O_1995,N_14961,N_14963);
xnor UO_1996 (O_1996,N_14893,N_14822);
or UO_1997 (O_1997,N_14833,N_14900);
and UO_1998 (O_1998,N_14822,N_14848);
nand UO_1999 (O_1999,N_14941,N_14980);
endmodule