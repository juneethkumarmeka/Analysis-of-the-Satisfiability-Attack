module basic_500_3000_500_4_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_291,In_187);
nor U1 (N_1,In_130,In_435);
and U2 (N_2,In_135,In_229);
nor U3 (N_3,In_404,In_303);
or U4 (N_4,In_199,In_390);
or U5 (N_5,In_237,In_407);
nand U6 (N_6,In_468,In_149);
or U7 (N_7,In_112,In_129);
or U8 (N_8,In_438,In_0);
nor U9 (N_9,In_363,In_201);
and U10 (N_10,In_327,In_341);
nand U11 (N_11,In_293,In_150);
nand U12 (N_12,In_410,In_364);
nor U13 (N_13,In_85,In_428);
nand U14 (N_14,In_420,In_459);
nand U15 (N_15,In_445,In_498);
nor U16 (N_16,In_421,In_412);
and U17 (N_17,In_96,In_484);
and U18 (N_18,In_178,In_153);
nor U19 (N_19,In_324,In_145);
nand U20 (N_20,In_336,In_117);
and U21 (N_21,In_343,In_450);
nor U22 (N_22,In_13,In_335);
nor U23 (N_23,In_443,In_193);
and U24 (N_24,In_15,In_362);
nor U25 (N_25,In_417,In_176);
or U26 (N_26,In_214,In_91);
nor U27 (N_27,In_42,In_350);
nor U28 (N_28,In_62,In_133);
and U29 (N_29,In_104,In_212);
nand U30 (N_30,In_409,In_499);
and U31 (N_31,In_281,In_477);
nand U32 (N_32,In_115,In_24);
and U33 (N_33,In_126,In_299);
and U34 (N_34,In_209,In_476);
and U35 (N_35,In_306,In_330);
and U36 (N_36,In_473,In_189);
nand U37 (N_37,In_180,In_304);
nand U38 (N_38,In_332,In_31);
or U39 (N_39,In_218,In_92);
or U40 (N_40,In_56,In_136);
or U41 (N_41,In_349,In_270);
nor U42 (N_42,In_458,In_173);
and U43 (N_43,In_400,In_282);
or U44 (N_44,In_406,In_479);
nor U45 (N_45,In_455,In_4);
and U46 (N_46,In_352,In_197);
and U47 (N_47,In_396,In_278);
nor U48 (N_48,In_177,In_379);
nand U49 (N_49,In_210,In_446);
and U50 (N_50,In_383,In_80);
or U51 (N_51,In_253,In_122);
and U52 (N_52,In_174,In_82);
and U53 (N_53,In_454,In_87);
and U54 (N_54,In_219,In_340);
and U55 (N_55,In_347,In_30);
or U56 (N_56,In_485,In_273);
or U57 (N_57,In_439,In_12);
and U58 (N_58,In_156,In_329);
and U59 (N_59,In_171,In_227);
nand U60 (N_60,In_296,In_372);
or U61 (N_61,In_375,In_26);
nor U62 (N_62,In_425,In_140);
nand U63 (N_63,In_7,In_194);
nor U64 (N_64,In_211,In_295);
nor U65 (N_65,In_146,In_257);
nor U66 (N_66,In_89,In_72);
nor U67 (N_67,In_249,In_21);
or U68 (N_68,In_23,In_206);
and U69 (N_69,In_142,In_483);
and U70 (N_70,In_441,In_27);
nor U71 (N_71,In_371,In_449);
and U72 (N_72,In_243,In_461);
nor U73 (N_73,In_319,In_25);
and U74 (N_74,In_471,In_127);
and U75 (N_75,In_360,In_312);
nor U76 (N_76,In_385,In_34);
nor U77 (N_77,In_275,In_154);
nor U78 (N_78,In_318,In_298);
or U79 (N_79,In_105,In_231);
nor U80 (N_80,In_74,In_120);
and U81 (N_81,In_116,In_262);
nor U82 (N_82,In_492,In_269);
xnor U83 (N_83,In_195,In_378);
nand U84 (N_84,In_457,In_365);
or U85 (N_85,In_422,In_57);
and U86 (N_86,In_393,In_307);
nand U87 (N_87,In_285,In_71);
or U88 (N_88,In_331,In_244);
or U89 (N_89,In_49,In_490);
nor U90 (N_90,In_292,In_143);
nor U91 (N_91,In_223,In_191);
or U92 (N_92,In_467,In_192);
and U93 (N_93,In_280,In_160);
nand U94 (N_94,In_283,In_75);
nor U95 (N_95,In_381,In_286);
or U96 (N_96,In_415,In_172);
or U97 (N_97,In_297,In_203);
and U98 (N_98,In_33,In_43);
and U99 (N_99,In_22,In_83);
nand U100 (N_100,In_272,In_155);
or U101 (N_101,In_6,In_469);
and U102 (N_102,In_121,In_388);
nand U103 (N_103,In_260,In_495);
nand U104 (N_104,In_41,In_370);
and U105 (N_105,In_402,In_328);
and U106 (N_106,In_44,In_188);
nor U107 (N_107,In_345,In_208);
nor U108 (N_108,In_185,In_353);
or U109 (N_109,In_426,In_221);
nand U110 (N_110,In_40,In_58);
nand U111 (N_111,In_491,In_430);
and U112 (N_112,In_76,In_494);
nor U113 (N_113,In_239,In_124);
nand U114 (N_114,In_79,In_405);
nand U115 (N_115,In_397,In_168);
nor U116 (N_116,In_241,In_157);
or U117 (N_117,In_423,In_392);
or U118 (N_118,In_95,In_399);
nand U119 (N_119,In_261,In_207);
nand U120 (N_120,In_464,In_376);
nand U121 (N_121,In_361,In_263);
nand U122 (N_122,In_256,In_337);
and U123 (N_123,In_152,In_451);
and U124 (N_124,In_148,In_141);
nand U125 (N_125,In_63,In_240);
or U126 (N_126,In_305,In_159);
and U127 (N_127,In_138,In_414);
nor U128 (N_128,In_179,In_248);
or U129 (N_129,In_108,In_204);
and U130 (N_130,In_213,In_252);
nor U131 (N_131,In_8,In_50);
or U132 (N_132,In_10,In_308);
or U133 (N_133,In_359,In_165);
and U134 (N_134,In_496,In_250);
nand U135 (N_135,In_169,In_186);
or U136 (N_136,In_369,In_61);
and U137 (N_137,In_109,In_478);
or U138 (N_138,In_367,In_333);
nand U139 (N_139,In_114,In_131);
nor U140 (N_140,In_39,In_453);
xnor U141 (N_141,In_356,In_416);
nor U142 (N_142,In_497,In_2);
nand U143 (N_143,In_432,In_132);
or U144 (N_144,In_488,In_486);
nand U145 (N_145,In_334,In_325);
nand U146 (N_146,In_401,In_216);
nor U147 (N_147,In_475,In_366);
nor U148 (N_148,In_437,In_166);
and U149 (N_149,In_339,In_51);
nand U150 (N_150,In_35,In_20);
nor U151 (N_151,In_232,In_300);
or U152 (N_152,In_81,In_190);
or U153 (N_153,In_301,In_164);
and U154 (N_154,In_265,In_53);
nand U155 (N_155,In_128,In_230);
or U156 (N_156,In_448,In_182);
and U157 (N_157,In_103,In_36);
nor U158 (N_158,In_18,In_175);
nor U159 (N_159,In_377,In_68);
xnor U160 (N_160,In_225,In_45);
nor U161 (N_161,In_54,In_309);
or U162 (N_162,In_162,In_344);
and U163 (N_163,In_16,In_88);
nand U164 (N_164,In_384,In_493);
xnor U165 (N_165,In_137,In_274);
nand U166 (N_166,In_258,In_419);
and U167 (N_167,In_480,In_351);
nor U168 (N_168,In_245,In_37);
or U169 (N_169,In_472,In_93);
nor U170 (N_170,In_264,In_101);
xor U171 (N_171,In_102,In_357);
nand U172 (N_172,In_271,In_107);
xnor U173 (N_173,In_342,In_470);
nor U174 (N_174,In_326,In_268);
nand U175 (N_175,In_289,In_202);
or U176 (N_176,In_317,In_65);
nand U177 (N_177,In_259,In_374);
nor U178 (N_178,In_234,In_302);
and U179 (N_179,In_147,In_411);
and U180 (N_180,In_125,In_346);
nand U181 (N_181,In_77,In_163);
nor U182 (N_182,In_84,In_434);
xor U183 (N_183,In_460,In_440);
nor U184 (N_184,In_100,In_196);
nand U185 (N_185,In_474,In_14);
nand U186 (N_186,In_380,In_73);
nor U187 (N_187,In_290,In_355);
nor U188 (N_188,In_255,In_391);
and U189 (N_189,In_170,In_481);
or U190 (N_190,In_246,In_70);
nand U191 (N_191,In_442,In_46);
nor U192 (N_192,In_228,In_408);
and U193 (N_193,In_320,In_447);
and U194 (N_194,In_452,In_236);
or U195 (N_195,In_348,In_394);
and U196 (N_196,In_354,In_183);
or U197 (N_197,In_386,In_322);
and U198 (N_198,In_395,In_413);
or U199 (N_199,In_123,In_48);
or U200 (N_200,In_266,In_251);
or U201 (N_201,In_277,In_482);
nor U202 (N_202,In_99,In_418);
nand U203 (N_203,In_28,In_118);
or U204 (N_204,In_279,In_288);
nand U205 (N_205,In_1,In_487);
nor U206 (N_206,In_294,In_224);
nand U207 (N_207,In_338,In_200);
nand U208 (N_208,In_184,In_3);
nand U209 (N_209,In_161,In_463);
nor U210 (N_210,In_69,In_238);
nand U211 (N_211,In_215,In_276);
and U212 (N_212,In_19,In_60);
and U213 (N_213,In_181,In_389);
and U214 (N_214,In_134,In_316);
nor U215 (N_215,In_67,In_226);
and U216 (N_216,In_456,In_323);
nand U217 (N_217,In_489,In_151);
or U218 (N_218,In_29,In_431);
nor U219 (N_219,In_64,In_313);
and U220 (N_220,In_314,In_110);
nor U221 (N_221,In_311,In_144);
or U222 (N_222,In_94,In_167);
xnor U223 (N_223,In_32,In_17);
or U224 (N_224,In_52,In_47);
nand U225 (N_225,In_466,In_55);
and U226 (N_226,In_90,In_358);
nand U227 (N_227,In_106,In_403);
or U228 (N_228,In_38,In_382);
nand U229 (N_229,In_97,In_233);
or U230 (N_230,In_310,In_158);
nor U231 (N_231,In_222,In_235);
or U232 (N_232,In_247,In_465);
nor U233 (N_233,In_66,In_368);
nand U234 (N_234,In_424,In_217);
and U235 (N_235,In_433,In_387);
nor U236 (N_236,In_78,In_373);
nand U237 (N_237,In_119,In_98);
and U238 (N_238,In_284,In_267);
and U239 (N_239,In_198,In_9);
xnor U240 (N_240,In_220,In_321);
nand U241 (N_241,In_86,In_139);
or U242 (N_242,In_436,In_315);
nand U243 (N_243,In_462,In_242);
or U244 (N_244,In_111,In_287);
or U245 (N_245,In_205,In_59);
nor U246 (N_246,In_444,In_429);
nor U247 (N_247,In_398,In_427);
or U248 (N_248,In_254,In_5);
nand U249 (N_249,In_11,In_113);
nand U250 (N_250,In_310,In_280);
nor U251 (N_251,In_439,In_461);
or U252 (N_252,In_126,In_3);
nor U253 (N_253,In_403,In_442);
xor U254 (N_254,In_204,In_353);
or U255 (N_255,In_46,In_148);
and U256 (N_256,In_325,In_498);
or U257 (N_257,In_320,In_433);
nor U258 (N_258,In_187,In_321);
nor U259 (N_259,In_232,In_419);
or U260 (N_260,In_405,In_222);
nand U261 (N_261,In_47,In_130);
or U262 (N_262,In_209,In_107);
nor U263 (N_263,In_320,In_228);
nand U264 (N_264,In_344,In_297);
or U265 (N_265,In_60,In_421);
or U266 (N_266,In_413,In_74);
or U267 (N_267,In_154,In_314);
nand U268 (N_268,In_156,In_486);
nor U269 (N_269,In_295,In_11);
and U270 (N_270,In_210,In_257);
nor U271 (N_271,In_190,In_226);
or U272 (N_272,In_171,In_426);
nand U273 (N_273,In_214,In_442);
nor U274 (N_274,In_429,In_155);
or U275 (N_275,In_431,In_300);
nand U276 (N_276,In_379,In_26);
nand U277 (N_277,In_352,In_300);
or U278 (N_278,In_24,In_212);
nor U279 (N_279,In_168,In_408);
nor U280 (N_280,In_386,In_50);
nor U281 (N_281,In_360,In_42);
or U282 (N_282,In_322,In_425);
nor U283 (N_283,In_20,In_169);
nor U284 (N_284,In_262,In_407);
or U285 (N_285,In_430,In_178);
nor U286 (N_286,In_107,In_451);
or U287 (N_287,In_408,In_330);
and U288 (N_288,In_205,In_297);
nand U289 (N_289,In_88,In_8);
xnor U290 (N_290,In_175,In_492);
xor U291 (N_291,In_168,In_383);
nand U292 (N_292,In_99,In_462);
or U293 (N_293,In_489,In_288);
or U294 (N_294,In_349,In_430);
or U295 (N_295,In_162,In_74);
nand U296 (N_296,In_188,In_314);
and U297 (N_297,In_432,In_269);
nor U298 (N_298,In_94,In_355);
or U299 (N_299,In_303,In_376);
and U300 (N_300,In_486,In_499);
nor U301 (N_301,In_321,In_357);
or U302 (N_302,In_45,In_256);
and U303 (N_303,In_412,In_179);
and U304 (N_304,In_465,In_484);
nand U305 (N_305,In_317,In_301);
and U306 (N_306,In_391,In_137);
or U307 (N_307,In_476,In_128);
and U308 (N_308,In_63,In_307);
nand U309 (N_309,In_261,In_257);
nand U310 (N_310,In_327,In_403);
or U311 (N_311,In_261,In_264);
or U312 (N_312,In_452,In_270);
and U313 (N_313,In_201,In_339);
nor U314 (N_314,In_262,In_20);
or U315 (N_315,In_294,In_64);
xnor U316 (N_316,In_144,In_405);
or U317 (N_317,In_479,In_81);
or U318 (N_318,In_3,In_153);
nand U319 (N_319,In_370,In_49);
or U320 (N_320,In_371,In_176);
nor U321 (N_321,In_131,In_421);
or U322 (N_322,In_114,In_413);
and U323 (N_323,In_291,In_153);
and U324 (N_324,In_436,In_444);
and U325 (N_325,In_402,In_248);
nor U326 (N_326,In_467,In_34);
nor U327 (N_327,In_49,In_335);
and U328 (N_328,In_299,In_256);
or U329 (N_329,In_286,In_361);
nand U330 (N_330,In_466,In_382);
nand U331 (N_331,In_226,In_35);
nor U332 (N_332,In_257,In_32);
and U333 (N_333,In_235,In_162);
nor U334 (N_334,In_3,In_424);
or U335 (N_335,In_429,In_92);
or U336 (N_336,In_274,In_92);
nand U337 (N_337,In_268,In_57);
xnor U338 (N_338,In_166,In_352);
and U339 (N_339,In_436,In_165);
or U340 (N_340,In_79,In_201);
and U341 (N_341,In_204,In_288);
nor U342 (N_342,In_340,In_281);
and U343 (N_343,In_367,In_177);
nor U344 (N_344,In_152,In_267);
or U345 (N_345,In_58,In_322);
nor U346 (N_346,In_100,In_250);
and U347 (N_347,In_91,In_76);
or U348 (N_348,In_185,In_171);
or U349 (N_349,In_57,In_253);
nand U350 (N_350,In_329,In_20);
and U351 (N_351,In_91,In_473);
nand U352 (N_352,In_382,In_262);
nand U353 (N_353,In_115,In_329);
and U354 (N_354,In_312,In_175);
nor U355 (N_355,In_140,In_79);
nor U356 (N_356,In_120,In_223);
nand U357 (N_357,In_409,In_140);
or U358 (N_358,In_405,In_116);
nand U359 (N_359,In_171,In_461);
or U360 (N_360,In_23,In_76);
nor U361 (N_361,In_26,In_83);
nand U362 (N_362,In_265,In_248);
or U363 (N_363,In_218,In_175);
or U364 (N_364,In_22,In_79);
nand U365 (N_365,In_233,In_74);
and U366 (N_366,In_130,In_216);
nor U367 (N_367,In_14,In_310);
xnor U368 (N_368,In_155,In_296);
nand U369 (N_369,In_223,In_13);
nand U370 (N_370,In_269,In_144);
nand U371 (N_371,In_41,In_128);
or U372 (N_372,In_398,In_24);
nor U373 (N_373,In_348,In_491);
or U374 (N_374,In_387,In_326);
and U375 (N_375,In_317,In_410);
nor U376 (N_376,In_407,In_209);
and U377 (N_377,In_416,In_239);
nand U378 (N_378,In_138,In_497);
and U379 (N_379,In_492,In_302);
nor U380 (N_380,In_260,In_428);
and U381 (N_381,In_410,In_196);
nand U382 (N_382,In_461,In_334);
nand U383 (N_383,In_218,In_7);
and U384 (N_384,In_174,In_61);
nand U385 (N_385,In_330,In_264);
nor U386 (N_386,In_251,In_467);
and U387 (N_387,In_424,In_376);
nor U388 (N_388,In_286,In_300);
and U389 (N_389,In_296,In_253);
nand U390 (N_390,In_332,In_425);
or U391 (N_391,In_381,In_320);
and U392 (N_392,In_330,In_401);
and U393 (N_393,In_25,In_266);
or U394 (N_394,In_16,In_112);
nand U395 (N_395,In_10,In_263);
and U396 (N_396,In_342,In_168);
xor U397 (N_397,In_154,In_373);
nor U398 (N_398,In_239,In_289);
nand U399 (N_399,In_153,In_409);
nor U400 (N_400,In_102,In_201);
and U401 (N_401,In_49,In_296);
and U402 (N_402,In_289,In_369);
and U403 (N_403,In_362,In_346);
and U404 (N_404,In_81,In_314);
nor U405 (N_405,In_47,In_160);
nor U406 (N_406,In_305,In_134);
or U407 (N_407,In_393,In_493);
nor U408 (N_408,In_218,In_232);
nand U409 (N_409,In_80,In_461);
or U410 (N_410,In_324,In_149);
nor U411 (N_411,In_216,In_252);
and U412 (N_412,In_403,In_190);
and U413 (N_413,In_311,In_178);
or U414 (N_414,In_233,In_186);
or U415 (N_415,In_236,In_41);
nor U416 (N_416,In_120,In_206);
and U417 (N_417,In_413,In_317);
xor U418 (N_418,In_364,In_270);
nand U419 (N_419,In_263,In_161);
and U420 (N_420,In_205,In_425);
and U421 (N_421,In_418,In_35);
or U422 (N_422,In_430,In_495);
or U423 (N_423,In_108,In_301);
nand U424 (N_424,In_340,In_479);
and U425 (N_425,In_74,In_376);
nor U426 (N_426,In_432,In_453);
nor U427 (N_427,In_129,In_384);
nor U428 (N_428,In_173,In_416);
nor U429 (N_429,In_196,In_463);
nand U430 (N_430,In_15,In_181);
nand U431 (N_431,In_280,In_86);
xnor U432 (N_432,In_488,In_137);
or U433 (N_433,In_402,In_35);
nand U434 (N_434,In_171,In_430);
or U435 (N_435,In_117,In_244);
and U436 (N_436,In_5,In_348);
nand U437 (N_437,In_280,In_24);
nor U438 (N_438,In_302,In_225);
nand U439 (N_439,In_436,In_486);
nor U440 (N_440,In_332,In_311);
and U441 (N_441,In_300,In_350);
nand U442 (N_442,In_153,In_449);
nand U443 (N_443,In_179,In_40);
or U444 (N_444,In_322,In_424);
nand U445 (N_445,In_469,In_489);
nand U446 (N_446,In_435,In_493);
xor U447 (N_447,In_483,In_68);
nand U448 (N_448,In_495,In_160);
nor U449 (N_449,In_123,In_259);
nor U450 (N_450,In_72,In_491);
nor U451 (N_451,In_131,In_464);
and U452 (N_452,In_84,In_493);
and U453 (N_453,In_423,In_313);
or U454 (N_454,In_142,In_318);
and U455 (N_455,In_211,In_161);
and U456 (N_456,In_489,In_474);
nand U457 (N_457,In_10,In_315);
nand U458 (N_458,In_256,In_211);
nor U459 (N_459,In_153,In_434);
nor U460 (N_460,In_319,In_242);
and U461 (N_461,In_315,In_465);
nand U462 (N_462,In_285,In_343);
and U463 (N_463,In_62,In_192);
or U464 (N_464,In_244,In_48);
nand U465 (N_465,In_97,In_248);
or U466 (N_466,In_457,In_140);
nor U467 (N_467,In_460,In_474);
nand U468 (N_468,In_417,In_122);
or U469 (N_469,In_175,In_387);
xnor U470 (N_470,In_112,In_498);
or U471 (N_471,In_401,In_440);
nand U472 (N_472,In_356,In_376);
and U473 (N_473,In_364,In_82);
or U474 (N_474,In_219,In_155);
nor U475 (N_475,In_429,In_375);
and U476 (N_476,In_249,In_414);
or U477 (N_477,In_102,In_115);
or U478 (N_478,In_118,In_166);
nor U479 (N_479,In_393,In_376);
or U480 (N_480,In_253,In_243);
nand U481 (N_481,In_454,In_265);
nor U482 (N_482,In_429,In_349);
nor U483 (N_483,In_260,In_336);
and U484 (N_484,In_157,In_108);
and U485 (N_485,In_30,In_196);
or U486 (N_486,In_241,In_146);
or U487 (N_487,In_26,In_468);
nand U488 (N_488,In_88,In_108);
nor U489 (N_489,In_182,In_149);
nor U490 (N_490,In_100,In_156);
nor U491 (N_491,In_82,In_8);
or U492 (N_492,In_80,In_261);
nor U493 (N_493,In_58,In_16);
nand U494 (N_494,In_381,In_40);
nand U495 (N_495,In_495,In_294);
and U496 (N_496,In_261,In_203);
and U497 (N_497,In_191,In_259);
or U498 (N_498,In_250,In_48);
or U499 (N_499,In_167,In_266);
nand U500 (N_500,In_274,In_420);
xnor U501 (N_501,In_253,In_228);
or U502 (N_502,In_356,In_17);
or U503 (N_503,In_183,In_67);
xnor U504 (N_504,In_473,In_26);
nor U505 (N_505,In_471,In_356);
or U506 (N_506,In_293,In_401);
nand U507 (N_507,In_493,In_234);
nor U508 (N_508,In_295,In_389);
nor U509 (N_509,In_260,In_153);
or U510 (N_510,In_163,In_114);
nor U511 (N_511,In_255,In_306);
or U512 (N_512,In_202,In_142);
nor U513 (N_513,In_353,In_449);
nand U514 (N_514,In_15,In_445);
nand U515 (N_515,In_278,In_0);
and U516 (N_516,In_396,In_153);
nand U517 (N_517,In_373,In_68);
xnor U518 (N_518,In_304,In_8);
and U519 (N_519,In_424,In_11);
nand U520 (N_520,In_230,In_119);
or U521 (N_521,In_483,In_39);
nor U522 (N_522,In_173,In_286);
and U523 (N_523,In_136,In_440);
or U524 (N_524,In_390,In_374);
nand U525 (N_525,In_195,In_6);
or U526 (N_526,In_302,In_59);
or U527 (N_527,In_472,In_466);
nand U528 (N_528,In_374,In_441);
nand U529 (N_529,In_89,In_337);
or U530 (N_530,In_73,In_249);
nor U531 (N_531,In_277,In_330);
nor U532 (N_532,In_431,In_161);
and U533 (N_533,In_434,In_192);
nor U534 (N_534,In_399,In_124);
and U535 (N_535,In_295,In_483);
nand U536 (N_536,In_318,In_343);
nor U537 (N_537,In_257,In_218);
nor U538 (N_538,In_387,In_224);
or U539 (N_539,In_437,In_303);
nor U540 (N_540,In_165,In_156);
nand U541 (N_541,In_374,In_288);
or U542 (N_542,In_284,In_421);
nand U543 (N_543,In_377,In_229);
or U544 (N_544,In_409,In_207);
xnor U545 (N_545,In_4,In_5);
and U546 (N_546,In_89,In_123);
nand U547 (N_547,In_191,In_491);
nor U548 (N_548,In_440,In_458);
nand U549 (N_549,In_326,In_442);
and U550 (N_550,In_206,In_386);
or U551 (N_551,In_381,In_56);
and U552 (N_552,In_332,In_384);
nand U553 (N_553,In_192,In_404);
or U554 (N_554,In_259,In_499);
nor U555 (N_555,In_329,In_318);
nand U556 (N_556,In_138,In_454);
nand U557 (N_557,In_426,In_184);
nand U558 (N_558,In_80,In_235);
nand U559 (N_559,In_464,In_394);
nand U560 (N_560,In_378,In_408);
nand U561 (N_561,In_231,In_125);
nand U562 (N_562,In_230,In_304);
nand U563 (N_563,In_329,In_256);
or U564 (N_564,In_221,In_169);
nand U565 (N_565,In_205,In_421);
or U566 (N_566,In_305,In_213);
nor U567 (N_567,In_34,In_369);
nand U568 (N_568,In_236,In_333);
and U569 (N_569,In_226,In_235);
xnor U570 (N_570,In_380,In_287);
or U571 (N_571,In_112,In_258);
nand U572 (N_572,In_210,In_426);
or U573 (N_573,In_354,In_173);
nand U574 (N_574,In_369,In_391);
nor U575 (N_575,In_462,In_395);
or U576 (N_576,In_329,In_279);
nand U577 (N_577,In_171,In_422);
nor U578 (N_578,In_266,In_339);
or U579 (N_579,In_336,In_274);
or U580 (N_580,In_334,In_331);
and U581 (N_581,In_106,In_306);
nand U582 (N_582,In_479,In_234);
nand U583 (N_583,In_142,In_185);
and U584 (N_584,In_494,In_110);
nand U585 (N_585,In_109,In_279);
nand U586 (N_586,In_243,In_349);
and U587 (N_587,In_374,In_237);
or U588 (N_588,In_168,In_36);
and U589 (N_589,In_91,In_328);
nor U590 (N_590,In_410,In_342);
or U591 (N_591,In_314,In_133);
or U592 (N_592,In_59,In_9);
nor U593 (N_593,In_75,In_157);
and U594 (N_594,In_214,In_293);
and U595 (N_595,In_211,In_147);
nand U596 (N_596,In_428,In_348);
or U597 (N_597,In_434,In_420);
nand U598 (N_598,In_359,In_193);
or U599 (N_599,In_295,In_68);
and U600 (N_600,In_497,In_450);
and U601 (N_601,In_304,In_14);
nor U602 (N_602,In_356,In_12);
and U603 (N_603,In_43,In_28);
or U604 (N_604,In_423,In_407);
nor U605 (N_605,In_131,In_199);
or U606 (N_606,In_193,In_1);
and U607 (N_607,In_267,In_472);
and U608 (N_608,In_436,In_290);
nand U609 (N_609,In_206,In_24);
nand U610 (N_610,In_77,In_80);
and U611 (N_611,In_18,In_44);
and U612 (N_612,In_183,In_63);
nand U613 (N_613,In_416,In_183);
xor U614 (N_614,In_201,In_382);
nand U615 (N_615,In_252,In_404);
or U616 (N_616,In_353,In_420);
and U617 (N_617,In_460,In_472);
nor U618 (N_618,In_473,In_249);
and U619 (N_619,In_182,In_168);
nor U620 (N_620,In_149,In_224);
and U621 (N_621,In_155,In_484);
nor U622 (N_622,In_18,In_99);
nand U623 (N_623,In_174,In_233);
nor U624 (N_624,In_190,In_277);
nor U625 (N_625,In_260,In_200);
nand U626 (N_626,In_478,In_15);
nand U627 (N_627,In_353,In_355);
nor U628 (N_628,In_336,In_384);
nor U629 (N_629,In_455,In_238);
or U630 (N_630,In_492,In_210);
or U631 (N_631,In_223,In_395);
xnor U632 (N_632,In_347,In_133);
nand U633 (N_633,In_405,In_333);
nor U634 (N_634,In_330,In_479);
nor U635 (N_635,In_246,In_20);
nand U636 (N_636,In_316,In_438);
nor U637 (N_637,In_299,In_140);
nand U638 (N_638,In_465,In_86);
and U639 (N_639,In_485,In_145);
or U640 (N_640,In_201,In_139);
or U641 (N_641,In_286,In_456);
and U642 (N_642,In_93,In_113);
nor U643 (N_643,In_355,In_439);
and U644 (N_644,In_422,In_142);
nor U645 (N_645,In_370,In_301);
nand U646 (N_646,In_116,In_150);
and U647 (N_647,In_376,In_17);
nand U648 (N_648,In_197,In_212);
and U649 (N_649,In_273,In_133);
or U650 (N_650,In_380,In_60);
and U651 (N_651,In_470,In_176);
and U652 (N_652,In_250,In_162);
or U653 (N_653,In_142,In_265);
and U654 (N_654,In_42,In_283);
nand U655 (N_655,In_160,In_55);
nand U656 (N_656,In_227,In_340);
nor U657 (N_657,In_237,In_421);
xnor U658 (N_658,In_463,In_17);
nand U659 (N_659,In_349,In_85);
or U660 (N_660,In_119,In_203);
or U661 (N_661,In_250,In_119);
xnor U662 (N_662,In_485,In_408);
or U663 (N_663,In_353,In_441);
xor U664 (N_664,In_241,In_171);
nand U665 (N_665,In_75,In_94);
xnor U666 (N_666,In_390,In_333);
or U667 (N_667,In_129,In_99);
and U668 (N_668,In_41,In_184);
nand U669 (N_669,In_76,In_40);
or U670 (N_670,In_471,In_223);
nor U671 (N_671,In_146,In_366);
or U672 (N_672,In_74,In_347);
nor U673 (N_673,In_169,In_362);
nand U674 (N_674,In_306,In_50);
nand U675 (N_675,In_319,In_474);
and U676 (N_676,In_242,In_401);
nor U677 (N_677,In_21,In_174);
or U678 (N_678,In_272,In_126);
or U679 (N_679,In_387,In_84);
or U680 (N_680,In_12,In_334);
nor U681 (N_681,In_361,In_268);
nand U682 (N_682,In_172,In_290);
nor U683 (N_683,In_10,In_223);
nand U684 (N_684,In_399,In_212);
or U685 (N_685,In_328,In_138);
nand U686 (N_686,In_80,In_294);
and U687 (N_687,In_114,In_124);
nor U688 (N_688,In_392,In_477);
nor U689 (N_689,In_429,In_89);
and U690 (N_690,In_263,In_144);
and U691 (N_691,In_479,In_1);
or U692 (N_692,In_242,In_96);
nand U693 (N_693,In_38,In_97);
nand U694 (N_694,In_78,In_75);
or U695 (N_695,In_330,In_109);
nand U696 (N_696,In_432,In_158);
xnor U697 (N_697,In_341,In_258);
nor U698 (N_698,In_362,In_357);
nor U699 (N_699,In_225,In_140);
nor U700 (N_700,In_120,In_172);
and U701 (N_701,In_401,In_127);
or U702 (N_702,In_33,In_329);
or U703 (N_703,In_440,In_324);
xnor U704 (N_704,In_91,In_135);
or U705 (N_705,In_174,In_241);
or U706 (N_706,In_306,In_491);
nand U707 (N_707,In_264,In_421);
nand U708 (N_708,In_448,In_27);
nand U709 (N_709,In_276,In_383);
or U710 (N_710,In_26,In_369);
and U711 (N_711,In_180,In_444);
or U712 (N_712,In_241,In_233);
nand U713 (N_713,In_282,In_143);
nor U714 (N_714,In_327,In_337);
nand U715 (N_715,In_57,In_247);
or U716 (N_716,In_310,In_67);
and U717 (N_717,In_274,In_428);
nand U718 (N_718,In_262,In_356);
nor U719 (N_719,In_100,In_177);
nor U720 (N_720,In_427,In_485);
nor U721 (N_721,In_414,In_247);
nor U722 (N_722,In_443,In_175);
or U723 (N_723,In_429,In_221);
or U724 (N_724,In_70,In_477);
nand U725 (N_725,In_214,In_342);
nand U726 (N_726,In_214,In_173);
nor U727 (N_727,In_118,In_286);
nor U728 (N_728,In_133,In_109);
nand U729 (N_729,In_130,In_288);
nor U730 (N_730,In_379,In_336);
or U731 (N_731,In_105,In_81);
or U732 (N_732,In_16,In_470);
or U733 (N_733,In_332,In_373);
and U734 (N_734,In_326,In_409);
nand U735 (N_735,In_61,In_216);
nand U736 (N_736,In_460,In_464);
nor U737 (N_737,In_317,In_355);
and U738 (N_738,In_423,In_65);
nor U739 (N_739,In_250,In_19);
nor U740 (N_740,In_114,In_472);
nor U741 (N_741,In_183,In_328);
or U742 (N_742,In_486,In_477);
or U743 (N_743,In_214,In_373);
and U744 (N_744,In_68,In_244);
nand U745 (N_745,In_333,In_159);
nor U746 (N_746,In_105,In_116);
xnor U747 (N_747,In_439,In_292);
and U748 (N_748,In_291,In_367);
and U749 (N_749,In_421,In_341);
nand U750 (N_750,N_615,N_179);
and U751 (N_751,N_284,N_228);
nand U752 (N_752,N_117,N_486);
and U753 (N_753,N_289,N_643);
and U754 (N_754,N_20,N_349);
or U755 (N_755,N_624,N_579);
nor U756 (N_756,N_736,N_204);
nand U757 (N_757,N_544,N_336);
or U758 (N_758,N_379,N_526);
and U759 (N_759,N_97,N_594);
or U760 (N_760,N_31,N_15);
nor U761 (N_761,N_461,N_528);
and U762 (N_762,N_191,N_398);
or U763 (N_763,N_280,N_676);
nor U764 (N_764,N_21,N_671);
and U765 (N_765,N_86,N_480);
and U766 (N_766,N_57,N_704);
nor U767 (N_767,N_463,N_450);
nand U768 (N_768,N_33,N_171);
and U769 (N_769,N_50,N_68);
nand U770 (N_770,N_523,N_721);
nand U771 (N_771,N_602,N_717);
and U772 (N_772,N_128,N_361);
or U773 (N_773,N_478,N_504);
nand U774 (N_774,N_340,N_282);
and U775 (N_775,N_456,N_407);
nor U776 (N_776,N_206,N_472);
nor U777 (N_777,N_420,N_550);
nor U778 (N_778,N_642,N_513);
or U779 (N_779,N_443,N_72);
nor U780 (N_780,N_663,N_66);
or U781 (N_781,N_134,N_583);
xnor U782 (N_782,N_434,N_484);
or U783 (N_783,N_144,N_245);
nor U784 (N_784,N_559,N_259);
nor U785 (N_785,N_600,N_331);
or U786 (N_786,N_525,N_227);
nand U787 (N_787,N_652,N_328);
nor U788 (N_788,N_535,N_726);
nand U789 (N_789,N_294,N_279);
nand U790 (N_790,N_77,N_35);
or U791 (N_791,N_271,N_555);
or U792 (N_792,N_22,N_418);
and U793 (N_793,N_178,N_741);
nand U794 (N_794,N_655,N_502);
and U795 (N_795,N_692,N_410);
nor U796 (N_796,N_306,N_565);
or U797 (N_797,N_733,N_576);
nand U798 (N_798,N_503,N_684);
or U799 (N_799,N_551,N_710);
nand U800 (N_800,N_681,N_476);
nor U801 (N_801,N_452,N_441);
xnor U802 (N_802,N_272,N_714);
nand U803 (N_803,N_173,N_275);
or U804 (N_804,N_326,N_490);
nor U805 (N_805,N_651,N_69);
nand U806 (N_806,N_689,N_24);
and U807 (N_807,N_554,N_256);
nor U808 (N_808,N_333,N_578);
or U809 (N_809,N_40,N_706);
nor U810 (N_810,N_744,N_739);
nand U811 (N_811,N_589,N_101);
and U812 (N_812,N_105,N_52);
and U813 (N_813,N_103,N_353);
nand U814 (N_814,N_577,N_136);
nor U815 (N_815,N_74,N_682);
nand U816 (N_816,N_295,N_633);
nand U817 (N_817,N_121,N_713);
nor U818 (N_818,N_75,N_728);
and U819 (N_819,N_674,N_483);
and U820 (N_820,N_512,N_668);
nor U821 (N_821,N_229,N_96);
nand U822 (N_822,N_561,N_91);
nand U823 (N_823,N_266,N_670);
nor U824 (N_824,N_237,N_261);
and U825 (N_825,N_425,N_214);
nor U826 (N_826,N_386,N_380);
and U827 (N_827,N_76,N_62);
nor U828 (N_828,N_357,N_735);
nand U829 (N_829,N_310,N_320);
nand U830 (N_830,N_520,N_162);
and U831 (N_831,N_392,N_677);
nand U832 (N_832,N_240,N_672);
nand U833 (N_833,N_612,N_404);
and U834 (N_834,N_730,N_182);
nand U835 (N_835,N_219,N_164);
xnor U836 (N_836,N_177,N_318);
and U837 (N_837,N_737,N_188);
nand U838 (N_838,N_274,N_248);
xor U839 (N_839,N_309,N_46);
nor U840 (N_840,N_531,N_140);
nor U841 (N_841,N_734,N_641);
and U842 (N_842,N_451,N_429);
nand U843 (N_843,N_12,N_319);
or U844 (N_844,N_607,N_571);
and U845 (N_845,N_104,N_359);
or U846 (N_846,N_65,N_546);
nor U847 (N_847,N_193,N_92);
or U848 (N_848,N_293,N_458);
or U849 (N_849,N_627,N_87);
and U850 (N_850,N_530,N_125);
and U851 (N_851,N_343,N_497);
or U852 (N_852,N_547,N_586);
nand U853 (N_853,N_30,N_16);
or U854 (N_854,N_285,N_393);
and U855 (N_855,N_374,N_675);
nor U856 (N_856,N_347,N_464);
nor U857 (N_857,N_515,N_370);
nand U858 (N_858,N_372,N_258);
nand U859 (N_859,N_252,N_745);
and U860 (N_860,N_149,N_118);
and U861 (N_861,N_291,N_685);
nor U862 (N_862,N_378,N_473);
nor U863 (N_863,N_647,N_697);
nor U864 (N_864,N_481,N_54);
nor U865 (N_865,N_569,N_63);
and U866 (N_866,N_13,N_221);
and U867 (N_867,N_367,N_596);
nor U868 (N_868,N_678,N_189);
and U869 (N_869,N_59,N_532);
xnor U870 (N_870,N_568,N_45);
nand U871 (N_871,N_648,N_616);
and U872 (N_872,N_416,N_585);
nor U873 (N_873,N_707,N_175);
nand U874 (N_874,N_743,N_169);
or U875 (N_875,N_58,N_270);
or U876 (N_876,N_649,N_738);
or U877 (N_877,N_342,N_511);
nand U878 (N_878,N_43,N_444);
or U879 (N_879,N_541,N_29);
nor U880 (N_880,N_421,N_605);
and U881 (N_881,N_67,N_247);
nor U882 (N_882,N_222,N_746);
nor U883 (N_883,N_190,N_584);
nand U884 (N_884,N_269,N_719);
and U885 (N_885,N_351,N_199);
and U886 (N_886,N_292,N_85);
or U887 (N_887,N_354,N_564);
nand U888 (N_888,N_202,N_211);
nand U889 (N_889,N_494,N_55);
or U890 (N_890,N_61,N_308);
xor U891 (N_891,N_510,N_341);
or U892 (N_892,N_712,N_241);
nor U893 (N_893,N_110,N_283);
and U894 (N_894,N_47,N_126);
nor U895 (N_895,N_246,N_657);
nand U896 (N_896,N_462,N_453);
or U897 (N_897,N_116,N_250);
or U898 (N_898,N_427,N_466);
and U899 (N_899,N_350,N_686);
or U900 (N_900,N_84,N_618);
nor U901 (N_901,N_225,N_366);
and U902 (N_902,N_377,N_181);
and U903 (N_903,N_608,N_623);
nor U904 (N_904,N_419,N_479);
and U905 (N_905,N_303,N_720);
nor U906 (N_906,N_749,N_552);
nand U907 (N_907,N_257,N_424);
and U908 (N_908,N_150,N_196);
and U909 (N_909,N_239,N_369);
nand U910 (N_910,N_163,N_335);
xnor U911 (N_911,N_231,N_606);
and U912 (N_912,N_263,N_519);
nor U913 (N_913,N_321,N_363);
and U914 (N_914,N_558,N_298);
or U915 (N_915,N_167,N_8);
nand U916 (N_916,N_455,N_338);
or U917 (N_917,N_17,N_93);
nor U918 (N_918,N_430,N_439);
nor U919 (N_919,N_115,N_698);
xor U920 (N_920,N_708,N_412);
nor U921 (N_921,N_488,N_414);
or U922 (N_922,N_114,N_10);
and U923 (N_923,N_400,N_251);
and U924 (N_924,N_603,N_305);
and U925 (N_925,N_390,N_540);
nor U926 (N_926,N_388,N_673);
or U927 (N_927,N_312,N_42);
nor U928 (N_928,N_688,N_145);
nor U929 (N_929,N_25,N_582);
or U930 (N_930,N_711,N_539);
nor U931 (N_931,N_650,N_2);
and U932 (N_932,N_448,N_469);
nor U933 (N_933,N_37,N_1);
nor U934 (N_934,N_518,N_224);
nor U935 (N_935,N_529,N_723);
or U936 (N_936,N_203,N_127);
or U937 (N_937,N_625,N_409);
and U938 (N_938,N_73,N_687);
nand U939 (N_939,N_747,N_212);
nor U940 (N_940,N_438,N_658);
xnor U941 (N_941,N_141,N_112);
and U942 (N_942,N_56,N_669);
nor U943 (N_943,N_475,N_487);
or U944 (N_944,N_71,N_146);
nand U945 (N_945,N_152,N_591);
nand U946 (N_946,N_516,N_667);
or U947 (N_947,N_653,N_459);
nand U948 (N_948,N_27,N_135);
or U949 (N_949,N_613,N_337);
and U950 (N_950,N_521,N_384);
nor U951 (N_951,N_417,N_235);
xor U952 (N_952,N_238,N_53);
nand U953 (N_953,N_208,N_123);
nor U954 (N_954,N_183,N_527);
or U955 (N_955,N_41,N_358);
nand U956 (N_956,N_659,N_273);
nor U957 (N_957,N_299,N_281);
nor U958 (N_958,N_78,N_243);
or U959 (N_959,N_543,N_18);
xnor U960 (N_960,N_38,N_664);
and U961 (N_961,N_130,N_524);
nor U962 (N_962,N_365,N_542);
and U963 (N_963,N_597,N_680);
and U964 (N_964,N_718,N_296);
nor U965 (N_965,N_645,N_156);
and U966 (N_966,N_402,N_352);
or U967 (N_967,N_396,N_210);
nand U968 (N_968,N_588,N_142);
and U969 (N_969,N_223,N_26);
and U970 (N_970,N_133,N_288);
nand U971 (N_971,N_611,N_99);
or U972 (N_972,N_406,N_656);
xor U973 (N_973,N_415,N_151);
or U974 (N_974,N_715,N_701);
nand U975 (N_975,N_209,N_98);
or U976 (N_976,N_81,N_106);
and U977 (N_977,N_82,N_88);
and U978 (N_978,N_313,N_34);
nand U979 (N_979,N_80,N_696);
or U980 (N_980,N_348,N_428);
nor U981 (N_981,N_264,N_344);
nor U982 (N_982,N_94,N_83);
or U983 (N_983,N_195,N_267);
nand U984 (N_984,N_387,N_454);
or U985 (N_985,N_644,N_180);
or U986 (N_986,N_620,N_375);
nor U987 (N_987,N_399,N_660);
nand U988 (N_988,N_360,N_562);
nor U989 (N_989,N_381,N_637);
or U990 (N_990,N_635,N_111);
nand U991 (N_991,N_595,N_630);
or U992 (N_992,N_489,N_422);
nor U993 (N_993,N_119,N_147);
nand U994 (N_994,N_95,N_3);
nand U995 (N_995,N_411,N_640);
and U996 (N_996,N_729,N_327);
nor U997 (N_997,N_634,N_44);
nor U998 (N_998,N_170,N_482);
or U999 (N_999,N_322,N_253);
and U1000 (N_1000,N_49,N_621);
xnor U1001 (N_1001,N_548,N_356);
or U1002 (N_1002,N_722,N_90);
or U1003 (N_1003,N_614,N_185);
or U1004 (N_1004,N_506,N_500);
xor U1005 (N_1005,N_699,N_693);
nor U1006 (N_1006,N_165,N_197);
nand U1007 (N_1007,N_437,N_646);
or U1008 (N_1008,N_447,N_545);
nor U1009 (N_1009,N_495,N_100);
nor U1010 (N_1010,N_330,N_218);
nor U1011 (N_1011,N_304,N_332);
nor U1012 (N_1012,N_186,N_345);
nor U1013 (N_1013,N_124,N_700);
and U1014 (N_1014,N_485,N_23);
nor U1015 (N_1015,N_587,N_391);
nor U1016 (N_1016,N_628,N_329);
and U1017 (N_1017,N_395,N_610);
and U1018 (N_1018,N_716,N_431);
and U1019 (N_1019,N_631,N_122);
and U1020 (N_1020,N_436,N_505);
or U1021 (N_1021,N_598,N_639);
nor U1022 (N_1022,N_724,N_198);
nor U1023 (N_1023,N_514,N_200);
or U1024 (N_1024,N_5,N_638);
or U1025 (N_1025,N_573,N_262);
or U1026 (N_1026,N_236,N_373);
or U1027 (N_1027,N_695,N_70);
nor U1028 (N_1028,N_496,N_622);
and U1029 (N_1029,N_389,N_317);
nor U1030 (N_1030,N_470,N_570);
and U1031 (N_1031,N_440,N_445);
and U1032 (N_1032,N_158,N_549);
nand U1033 (N_1033,N_629,N_255);
and U1034 (N_1034,N_575,N_553);
nor U1035 (N_1035,N_538,N_148);
nand U1036 (N_1036,N_19,N_590);
nor U1037 (N_1037,N_626,N_307);
and U1038 (N_1038,N_460,N_11);
or U1039 (N_1039,N_205,N_446);
nand U1040 (N_1040,N_731,N_7);
nor U1041 (N_1041,N_435,N_268);
nor U1042 (N_1042,N_536,N_507);
and U1043 (N_1043,N_168,N_449);
nor U1044 (N_1044,N_371,N_468);
nor U1045 (N_1045,N_403,N_315);
or U1046 (N_1046,N_14,N_39);
and U1047 (N_1047,N_159,N_323);
and U1048 (N_1048,N_581,N_609);
or U1049 (N_1049,N_471,N_316);
or U1050 (N_1050,N_244,N_194);
or U1051 (N_1051,N_423,N_477);
and U1052 (N_1052,N_385,N_683);
or U1053 (N_1053,N_230,N_234);
or U1054 (N_1054,N_89,N_220);
nand U1055 (N_1055,N_28,N_566);
nand U1056 (N_1056,N_691,N_679);
and U1057 (N_1057,N_9,N_465);
and U1058 (N_1058,N_426,N_301);
nor U1059 (N_1059,N_709,N_413);
nand U1060 (N_1060,N_401,N_155);
and U1061 (N_1061,N_432,N_534);
and U1062 (N_1062,N_4,N_474);
or U1063 (N_1063,N_604,N_129);
or U1064 (N_1064,N_232,N_113);
nor U1065 (N_1065,N_742,N_302);
nand U1066 (N_1066,N_355,N_109);
nor U1067 (N_1067,N_32,N_160);
and U1068 (N_1068,N_36,N_467);
nor U1069 (N_1069,N_174,N_311);
nor U1070 (N_1070,N_740,N_533);
nand U1071 (N_1071,N_153,N_498);
nor U1072 (N_1072,N_705,N_102);
and U1073 (N_1073,N_201,N_314);
and U1074 (N_1074,N_226,N_143);
nor U1075 (N_1075,N_702,N_286);
nand U1076 (N_1076,N_216,N_166);
nand U1077 (N_1077,N_694,N_325);
or U1078 (N_1078,N_60,N_508);
nand U1079 (N_1079,N_563,N_132);
nand U1080 (N_1080,N_64,N_433);
or U1081 (N_1081,N_48,N_601);
or U1082 (N_1082,N_139,N_249);
and U1083 (N_1083,N_654,N_215);
and U1084 (N_1084,N_405,N_364);
and U1085 (N_1085,N_161,N_287);
xnor U1086 (N_1086,N_107,N_176);
nand U1087 (N_1087,N_278,N_580);
or U1088 (N_1088,N_6,N_207);
or U1089 (N_1089,N_408,N_619);
nand U1090 (N_1090,N_491,N_632);
or U1091 (N_1091,N_137,N_556);
nor U1092 (N_1092,N_690,N_703);
and U1093 (N_1093,N_265,N_233);
nand U1094 (N_1094,N_276,N_368);
and U1095 (N_1095,N_394,N_254);
or U1096 (N_1096,N_334,N_172);
or U1097 (N_1097,N_509,N_666);
and U1098 (N_1098,N_383,N_157);
or U1099 (N_1099,N_187,N_593);
nor U1100 (N_1100,N_154,N_662);
nor U1101 (N_1101,N_636,N_184);
nor U1102 (N_1102,N_108,N_324);
nor U1103 (N_1103,N_51,N_574);
nand U1104 (N_1104,N_732,N_493);
or U1105 (N_1105,N_242,N_192);
nand U1106 (N_1106,N_362,N_297);
nor U1107 (N_1107,N_260,N_492);
nor U1108 (N_1108,N_748,N_572);
nand U1109 (N_1109,N_665,N_0);
and U1110 (N_1110,N_537,N_277);
nor U1111 (N_1111,N_120,N_397);
and U1112 (N_1112,N_557,N_131);
nor U1113 (N_1113,N_457,N_560);
or U1114 (N_1114,N_617,N_727);
or U1115 (N_1115,N_567,N_599);
or U1116 (N_1116,N_501,N_522);
nor U1117 (N_1117,N_499,N_346);
nor U1118 (N_1118,N_442,N_217);
and U1119 (N_1119,N_138,N_300);
nand U1120 (N_1120,N_382,N_517);
nor U1121 (N_1121,N_79,N_213);
nor U1122 (N_1122,N_592,N_376);
nand U1123 (N_1123,N_661,N_290);
nor U1124 (N_1124,N_725,N_339);
nor U1125 (N_1125,N_397,N_749);
nor U1126 (N_1126,N_404,N_267);
nand U1127 (N_1127,N_655,N_92);
nor U1128 (N_1128,N_484,N_461);
and U1129 (N_1129,N_606,N_206);
nand U1130 (N_1130,N_609,N_165);
nor U1131 (N_1131,N_748,N_233);
or U1132 (N_1132,N_309,N_670);
nand U1133 (N_1133,N_84,N_568);
and U1134 (N_1134,N_702,N_203);
nor U1135 (N_1135,N_228,N_334);
nand U1136 (N_1136,N_12,N_613);
nand U1137 (N_1137,N_620,N_140);
nand U1138 (N_1138,N_57,N_12);
or U1139 (N_1139,N_289,N_81);
and U1140 (N_1140,N_534,N_232);
nor U1141 (N_1141,N_213,N_80);
or U1142 (N_1142,N_413,N_74);
or U1143 (N_1143,N_478,N_413);
and U1144 (N_1144,N_75,N_56);
nand U1145 (N_1145,N_469,N_545);
and U1146 (N_1146,N_378,N_397);
or U1147 (N_1147,N_121,N_729);
and U1148 (N_1148,N_428,N_659);
and U1149 (N_1149,N_331,N_54);
or U1150 (N_1150,N_215,N_692);
nand U1151 (N_1151,N_452,N_384);
or U1152 (N_1152,N_76,N_287);
nor U1153 (N_1153,N_508,N_461);
nand U1154 (N_1154,N_725,N_155);
or U1155 (N_1155,N_374,N_612);
nor U1156 (N_1156,N_114,N_388);
nor U1157 (N_1157,N_343,N_396);
nor U1158 (N_1158,N_670,N_424);
and U1159 (N_1159,N_551,N_387);
xnor U1160 (N_1160,N_198,N_728);
or U1161 (N_1161,N_618,N_441);
and U1162 (N_1162,N_58,N_417);
nand U1163 (N_1163,N_720,N_355);
nand U1164 (N_1164,N_416,N_565);
nor U1165 (N_1165,N_479,N_628);
nand U1166 (N_1166,N_399,N_382);
nand U1167 (N_1167,N_26,N_154);
or U1168 (N_1168,N_385,N_384);
or U1169 (N_1169,N_306,N_239);
nand U1170 (N_1170,N_700,N_591);
or U1171 (N_1171,N_390,N_340);
and U1172 (N_1172,N_275,N_609);
nand U1173 (N_1173,N_211,N_285);
and U1174 (N_1174,N_626,N_87);
and U1175 (N_1175,N_698,N_372);
nor U1176 (N_1176,N_392,N_657);
nor U1177 (N_1177,N_479,N_150);
nand U1178 (N_1178,N_76,N_457);
nand U1179 (N_1179,N_135,N_560);
nand U1180 (N_1180,N_544,N_47);
and U1181 (N_1181,N_428,N_566);
or U1182 (N_1182,N_92,N_149);
nor U1183 (N_1183,N_731,N_71);
nand U1184 (N_1184,N_63,N_335);
nor U1185 (N_1185,N_232,N_628);
nor U1186 (N_1186,N_5,N_711);
and U1187 (N_1187,N_571,N_214);
nand U1188 (N_1188,N_48,N_571);
and U1189 (N_1189,N_455,N_287);
or U1190 (N_1190,N_663,N_546);
xnor U1191 (N_1191,N_302,N_51);
and U1192 (N_1192,N_88,N_715);
nor U1193 (N_1193,N_735,N_576);
nor U1194 (N_1194,N_611,N_399);
and U1195 (N_1195,N_642,N_318);
and U1196 (N_1196,N_296,N_416);
nand U1197 (N_1197,N_685,N_422);
nand U1198 (N_1198,N_133,N_291);
or U1199 (N_1199,N_490,N_379);
nor U1200 (N_1200,N_360,N_702);
or U1201 (N_1201,N_741,N_198);
and U1202 (N_1202,N_209,N_327);
nand U1203 (N_1203,N_210,N_566);
nor U1204 (N_1204,N_90,N_662);
and U1205 (N_1205,N_301,N_102);
nand U1206 (N_1206,N_506,N_110);
and U1207 (N_1207,N_464,N_390);
nand U1208 (N_1208,N_427,N_381);
or U1209 (N_1209,N_136,N_632);
nor U1210 (N_1210,N_322,N_437);
and U1211 (N_1211,N_453,N_640);
nand U1212 (N_1212,N_698,N_169);
or U1213 (N_1213,N_636,N_377);
nor U1214 (N_1214,N_394,N_51);
nor U1215 (N_1215,N_620,N_500);
nand U1216 (N_1216,N_333,N_241);
nor U1217 (N_1217,N_430,N_350);
nor U1218 (N_1218,N_706,N_347);
and U1219 (N_1219,N_490,N_624);
and U1220 (N_1220,N_6,N_145);
nor U1221 (N_1221,N_148,N_7);
nor U1222 (N_1222,N_554,N_560);
xnor U1223 (N_1223,N_83,N_703);
nand U1224 (N_1224,N_157,N_626);
or U1225 (N_1225,N_240,N_351);
or U1226 (N_1226,N_473,N_220);
xor U1227 (N_1227,N_705,N_319);
nand U1228 (N_1228,N_452,N_167);
nand U1229 (N_1229,N_262,N_658);
nand U1230 (N_1230,N_330,N_275);
nor U1231 (N_1231,N_523,N_168);
nor U1232 (N_1232,N_149,N_71);
or U1233 (N_1233,N_42,N_572);
nand U1234 (N_1234,N_176,N_642);
or U1235 (N_1235,N_291,N_330);
nand U1236 (N_1236,N_41,N_549);
nand U1237 (N_1237,N_324,N_467);
and U1238 (N_1238,N_316,N_275);
or U1239 (N_1239,N_717,N_655);
nand U1240 (N_1240,N_229,N_76);
and U1241 (N_1241,N_67,N_656);
nand U1242 (N_1242,N_208,N_700);
nand U1243 (N_1243,N_312,N_335);
nor U1244 (N_1244,N_238,N_21);
nand U1245 (N_1245,N_77,N_130);
nand U1246 (N_1246,N_674,N_720);
or U1247 (N_1247,N_667,N_148);
nor U1248 (N_1248,N_425,N_193);
nor U1249 (N_1249,N_427,N_389);
and U1250 (N_1250,N_509,N_741);
or U1251 (N_1251,N_559,N_666);
or U1252 (N_1252,N_467,N_608);
nor U1253 (N_1253,N_244,N_501);
or U1254 (N_1254,N_274,N_23);
and U1255 (N_1255,N_670,N_104);
nand U1256 (N_1256,N_21,N_744);
xnor U1257 (N_1257,N_552,N_324);
and U1258 (N_1258,N_670,N_106);
nor U1259 (N_1259,N_329,N_650);
and U1260 (N_1260,N_682,N_451);
and U1261 (N_1261,N_730,N_346);
or U1262 (N_1262,N_393,N_67);
nand U1263 (N_1263,N_686,N_249);
and U1264 (N_1264,N_451,N_718);
or U1265 (N_1265,N_719,N_2);
nor U1266 (N_1266,N_679,N_391);
and U1267 (N_1267,N_441,N_235);
nand U1268 (N_1268,N_307,N_591);
nand U1269 (N_1269,N_571,N_727);
nand U1270 (N_1270,N_374,N_93);
nand U1271 (N_1271,N_149,N_413);
nor U1272 (N_1272,N_615,N_356);
and U1273 (N_1273,N_574,N_643);
nor U1274 (N_1274,N_336,N_746);
xor U1275 (N_1275,N_9,N_47);
and U1276 (N_1276,N_185,N_327);
nor U1277 (N_1277,N_343,N_368);
or U1278 (N_1278,N_501,N_5);
nor U1279 (N_1279,N_732,N_46);
nand U1280 (N_1280,N_176,N_640);
nand U1281 (N_1281,N_455,N_480);
nand U1282 (N_1282,N_543,N_315);
or U1283 (N_1283,N_307,N_463);
nand U1284 (N_1284,N_179,N_23);
nor U1285 (N_1285,N_261,N_76);
and U1286 (N_1286,N_344,N_733);
nor U1287 (N_1287,N_117,N_442);
nand U1288 (N_1288,N_141,N_74);
nand U1289 (N_1289,N_415,N_226);
or U1290 (N_1290,N_162,N_634);
nor U1291 (N_1291,N_229,N_146);
nor U1292 (N_1292,N_327,N_479);
nor U1293 (N_1293,N_77,N_94);
or U1294 (N_1294,N_749,N_523);
or U1295 (N_1295,N_74,N_182);
or U1296 (N_1296,N_129,N_593);
nand U1297 (N_1297,N_590,N_729);
nand U1298 (N_1298,N_200,N_384);
or U1299 (N_1299,N_98,N_368);
or U1300 (N_1300,N_63,N_148);
nand U1301 (N_1301,N_398,N_450);
nand U1302 (N_1302,N_183,N_39);
and U1303 (N_1303,N_272,N_538);
nor U1304 (N_1304,N_497,N_383);
or U1305 (N_1305,N_157,N_53);
and U1306 (N_1306,N_400,N_135);
nand U1307 (N_1307,N_461,N_709);
nand U1308 (N_1308,N_3,N_544);
or U1309 (N_1309,N_516,N_114);
and U1310 (N_1310,N_412,N_743);
or U1311 (N_1311,N_265,N_178);
nand U1312 (N_1312,N_93,N_491);
or U1313 (N_1313,N_675,N_146);
nand U1314 (N_1314,N_552,N_736);
or U1315 (N_1315,N_728,N_598);
and U1316 (N_1316,N_599,N_76);
or U1317 (N_1317,N_290,N_319);
and U1318 (N_1318,N_411,N_198);
xnor U1319 (N_1319,N_187,N_530);
and U1320 (N_1320,N_64,N_436);
nand U1321 (N_1321,N_61,N_289);
or U1322 (N_1322,N_316,N_521);
nor U1323 (N_1323,N_725,N_353);
nand U1324 (N_1324,N_469,N_646);
nand U1325 (N_1325,N_658,N_177);
and U1326 (N_1326,N_641,N_122);
and U1327 (N_1327,N_260,N_150);
and U1328 (N_1328,N_675,N_215);
nand U1329 (N_1329,N_450,N_221);
and U1330 (N_1330,N_77,N_144);
nor U1331 (N_1331,N_589,N_495);
nor U1332 (N_1332,N_539,N_380);
and U1333 (N_1333,N_249,N_91);
and U1334 (N_1334,N_354,N_149);
and U1335 (N_1335,N_289,N_560);
nor U1336 (N_1336,N_194,N_630);
and U1337 (N_1337,N_273,N_25);
or U1338 (N_1338,N_40,N_164);
nand U1339 (N_1339,N_498,N_64);
and U1340 (N_1340,N_277,N_60);
or U1341 (N_1341,N_440,N_182);
or U1342 (N_1342,N_281,N_508);
or U1343 (N_1343,N_123,N_546);
xnor U1344 (N_1344,N_320,N_303);
nand U1345 (N_1345,N_450,N_425);
nand U1346 (N_1346,N_595,N_394);
nor U1347 (N_1347,N_325,N_430);
nand U1348 (N_1348,N_79,N_24);
nand U1349 (N_1349,N_355,N_324);
and U1350 (N_1350,N_460,N_33);
and U1351 (N_1351,N_448,N_661);
or U1352 (N_1352,N_78,N_170);
nand U1353 (N_1353,N_567,N_126);
and U1354 (N_1354,N_102,N_430);
nand U1355 (N_1355,N_540,N_369);
nand U1356 (N_1356,N_34,N_101);
nand U1357 (N_1357,N_47,N_175);
xnor U1358 (N_1358,N_239,N_132);
nor U1359 (N_1359,N_605,N_42);
nor U1360 (N_1360,N_62,N_642);
nand U1361 (N_1361,N_594,N_365);
or U1362 (N_1362,N_119,N_394);
nor U1363 (N_1363,N_2,N_485);
or U1364 (N_1364,N_302,N_647);
or U1365 (N_1365,N_189,N_428);
nor U1366 (N_1366,N_616,N_228);
nor U1367 (N_1367,N_312,N_550);
nor U1368 (N_1368,N_312,N_452);
nand U1369 (N_1369,N_141,N_111);
nand U1370 (N_1370,N_513,N_350);
and U1371 (N_1371,N_682,N_460);
nand U1372 (N_1372,N_41,N_493);
or U1373 (N_1373,N_746,N_231);
nor U1374 (N_1374,N_720,N_579);
and U1375 (N_1375,N_86,N_511);
nand U1376 (N_1376,N_224,N_669);
and U1377 (N_1377,N_68,N_367);
nor U1378 (N_1378,N_461,N_110);
or U1379 (N_1379,N_69,N_64);
nand U1380 (N_1380,N_103,N_95);
nor U1381 (N_1381,N_9,N_491);
and U1382 (N_1382,N_73,N_34);
nor U1383 (N_1383,N_426,N_65);
or U1384 (N_1384,N_632,N_525);
and U1385 (N_1385,N_174,N_677);
and U1386 (N_1386,N_399,N_230);
or U1387 (N_1387,N_535,N_332);
and U1388 (N_1388,N_748,N_685);
nand U1389 (N_1389,N_669,N_1);
nand U1390 (N_1390,N_524,N_454);
and U1391 (N_1391,N_707,N_430);
or U1392 (N_1392,N_699,N_356);
or U1393 (N_1393,N_544,N_92);
and U1394 (N_1394,N_270,N_506);
nor U1395 (N_1395,N_114,N_47);
or U1396 (N_1396,N_51,N_511);
nor U1397 (N_1397,N_341,N_161);
nand U1398 (N_1398,N_138,N_587);
nor U1399 (N_1399,N_321,N_14);
and U1400 (N_1400,N_599,N_592);
and U1401 (N_1401,N_597,N_602);
or U1402 (N_1402,N_142,N_332);
nand U1403 (N_1403,N_354,N_410);
or U1404 (N_1404,N_483,N_157);
nand U1405 (N_1405,N_81,N_666);
nand U1406 (N_1406,N_198,N_228);
xnor U1407 (N_1407,N_694,N_342);
or U1408 (N_1408,N_633,N_357);
nor U1409 (N_1409,N_292,N_132);
and U1410 (N_1410,N_134,N_262);
or U1411 (N_1411,N_48,N_497);
or U1412 (N_1412,N_20,N_284);
and U1413 (N_1413,N_175,N_229);
or U1414 (N_1414,N_418,N_240);
nand U1415 (N_1415,N_608,N_583);
and U1416 (N_1416,N_551,N_62);
nand U1417 (N_1417,N_554,N_712);
nand U1418 (N_1418,N_279,N_411);
nand U1419 (N_1419,N_441,N_253);
and U1420 (N_1420,N_279,N_545);
nand U1421 (N_1421,N_25,N_506);
xnor U1422 (N_1422,N_48,N_657);
nor U1423 (N_1423,N_262,N_532);
nor U1424 (N_1424,N_363,N_659);
and U1425 (N_1425,N_323,N_282);
or U1426 (N_1426,N_91,N_219);
and U1427 (N_1427,N_642,N_551);
xnor U1428 (N_1428,N_133,N_261);
or U1429 (N_1429,N_108,N_381);
nor U1430 (N_1430,N_743,N_469);
nor U1431 (N_1431,N_624,N_401);
or U1432 (N_1432,N_41,N_490);
or U1433 (N_1433,N_228,N_230);
xnor U1434 (N_1434,N_506,N_673);
nand U1435 (N_1435,N_130,N_622);
nand U1436 (N_1436,N_284,N_627);
and U1437 (N_1437,N_371,N_135);
nand U1438 (N_1438,N_487,N_736);
nor U1439 (N_1439,N_121,N_608);
or U1440 (N_1440,N_125,N_74);
and U1441 (N_1441,N_154,N_659);
nand U1442 (N_1442,N_417,N_456);
nor U1443 (N_1443,N_39,N_166);
nand U1444 (N_1444,N_666,N_7);
nand U1445 (N_1445,N_349,N_174);
nand U1446 (N_1446,N_185,N_170);
or U1447 (N_1447,N_681,N_331);
or U1448 (N_1448,N_681,N_0);
and U1449 (N_1449,N_250,N_452);
nor U1450 (N_1450,N_698,N_410);
or U1451 (N_1451,N_719,N_45);
or U1452 (N_1452,N_597,N_696);
nand U1453 (N_1453,N_138,N_295);
or U1454 (N_1454,N_220,N_307);
and U1455 (N_1455,N_454,N_83);
nand U1456 (N_1456,N_75,N_484);
nand U1457 (N_1457,N_274,N_624);
or U1458 (N_1458,N_409,N_486);
and U1459 (N_1459,N_39,N_114);
nand U1460 (N_1460,N_180,N_144);
nand U1461 (N_1461,N_702,N_181);
or U1462 (N_1462,N_140,N_194);
nand U1463 (N_1463,N_73,N_211);
nand U1464 (N_1464,N_490,N_293);
or U1465 (N_1465,N_582,N_330);
nand U1466 (N_1466,N_399,N_680);
nor U1467 (N_1467,N_556,N_594);
nand U1468 (N_1468,N_689,N_262);
xnor U1469 (N_1469,N_313,N_454);
or U1470 (N_1470,N_186,N_185);
nor U1471 (N_1471,N_580,N_562);
and U1472 (N_1472,N_475,N_11);
nand U1473 (N_1473,N_293,N_242);
and U1474 (N_1474,N_67,N_333);
and U1475 (N_1475,N_402,N_692);
and U1476 (N_1476,N_611,N_520);
nand U1477 (N_1477,N_679,N_384);
nand U1478 (N_1478,N_544,N_744);
nor U1479 (N_1479,N_597,N_175);
nor U1480 (N_1480,N_741,N_641);
and U1481 (N_1481,N_682,N_334);
or U1482 (N_1482,N_639,N_163);
nand U1483 (N_1483,N_658,N_634);
nor U1484 (N_1484,N_107,N_76);
nand U1485 (N_1485,N_69,N_71);
nor U1486 (N_1486,N_700,N_620);
nand U1487 (N_1487,N_345,N_639);
nor U1488 (N_1488,N_532,N_20);
or U1489 (N_1489,N_111,N_535);
nor U1490 (N_1490,N_71,N_526);
nor U1491 (N_1491,N_528,N_589);
xnor U1492 (N_1492,N_625,N_230);
nor U1493 (N_1493,N_254,N_190);
and U1494 (N_1494,N_202,N_177);
or U1495 (N_1495,N_95,N_401);
nor U1496 (N_1496,N_426,N_274);
nor U1497 (N_1497,N_613,N_320);
and U1498 (N_1498,N_252,N_327);
or U1499 (N_1499,N_272,N_141);
nand U1500 (N_1500,N_917,N_923);
nand U1501 (N_1501,N_920,N_876);
nand U1502 (N_1502,N_1011,N_863);
or U1503 (N_1503,N_1483,N_1434);
nand U1504 (N_1504,N_1476,N_855);
or U1505 (N_1505,N_785,N_1365);
nand U1506 (N_1506,N_757,N_1376);
and U1507 (N_1507,N_853,N_985);
or U1508 (N_1508,N_1068,N_1085);
or U1509 (N_1509,N_1331,N_1119);
and U1510 (N_1510,N_1448,N_847);
and U1511 (N_1511,N_867,N_780);
xnor U1512 (N_1512,N_1008,N_758);
nand U1513 (N_1513,N_1254,N_1016);
nand U1514 (N_1514,N_882,N_1407);
nand U1515 (N_1515,N_1299,N_1169);
nor U1516 (N_1516,N_1040,N_997);
nor U1517 (N_1517,N_891,N_1189);
nor U1518 (N_1518,N_1202,N_772);
nor U1519 (N_1519,N_816,N_1444);
and U1520 (N_1520,N_1067,N_1478);
nand U1521 (N_1521,N_1081,N_1475);
nor U1522 (N_1522,N_1391,N_1193);
nor U1523 (N_1523,N_992,N_1443);
or U1524 (N_1524,N_1106,N_764);
nor U1525 (N_1525,N_1465,N_1079);
or U1526 (N_1526,N_1156,N_821);
nand U1527 (N_1527,N_1198,N_941);
or U1528 (N_1528,N_881,N_1241);
and U1529 (N_1529,N_844,N_811);
and U1530 (N_1530,N_1248,N_1394);
or U1531 (N_1531,N_1245,N_813);
nand U1532 (N_1532,N_879,N_1378);
nor U1533 (N_1533,N_902,N_1278);
nand U1534 (N_1534,N_1204,N_971);
nand U1535 (N_1535,N_1264,N_1321);
nor U1536 (N_1536,N_940,N_909);
or U1537 (N_1537,N_1025,N_1127);
and U1538 (N_1538,N_1295,N_1308);
nor U1539 (N_1539,N_954,N_931);
nand U1540 (N_1540,N_1281,N_1061);
nor U1541 (N_1541,N_1269,N_1334);
or U1542 (N_1542,N_1133,N_922);
or U1543 (N_1543,N_1201,N_825);
nand U1544 (N_1544,N_1172,N_1010);
nand U1545 (N_1545,N_1356,N_1107);
nand U1546 (N_1546,N_1153,N_1333);
or U1547 (N_1547,N_1194,N_955);
and U1548 (N_1548,N_1024,N_1195);
and U1549 (N_1549,N_1249,N_1023);
and U1550 (N_1550,N_1030,N_1028);
and U1551 (N_1551,N_1335,N_973);
nand U1552 (N_1552,N_1418,N_1151);
xor U1553 (N_1553,N_1468,N_1291);
nor U1554 (N_1554,N_1206,N_1311);
and U1555 (N_1555,N_1213,N_1284);
nand U1556 (N_1556,N_1089,N_1084);
nand U1557 (N_1557,N_823,N_1027);
nor U1558 (N_1558,N_1366,N_901);
and U1559 (N_1559,N_1446,N_1293);
and U1560 (N_1560,N_1420,N_1176);
or U1561 (N_1561,N_1439,N_1373);
and U1562 (N_1562,N_1362,N_854);
nand U1563 (N_1563,N_1041,N_766);
and U1564 (N_1564,N_978,N_1327);
xnor U1565 (N_1565,N_1124,N_1170);
or U1566 (N_1566,N_967,N_841);
nand U1567 (N_1567,N_1340,N_988);
nand U1568 (N_1568,N_1427,N_953);
and U1569 (N_1569,N_871,N_752);
or U1570 (N_1570,N_875,N_1401);
or U1571 (N_1571,N_958,N_1363);
and U1572 (N_1572,N_1111,N_1410);
nand U1573 (N_1573,N_1185,N_1228);
nor U1574 (N_1574,N_982,N_1268);
or U1575 (N_1575,N_1021,N_1073);
and U1576 (N_1576,N_1368,N_899);
nor U1577 (N_1577,N_1217,N_1005);
nand U1578 (N_1578,N_1015,N_1454);
or U1579 (N_1579,N_1052,N_1094);
and U1580 (N_1580,N_801,N_1338);
and U1581 (N_1581,N_1115,N_810);
nand U1582 (N_1582,N_1009,N_1045);
nand U1583 (N_1583,N_820,N_1088);
or U1584 (N_1584,N_1237,N_1148);
xnor U1585 (N_1585,N_1162,N_1223);
nand U1586 (N_1586,N_800,N_1285);
nor U1587 (N_1587,N_834,N_1186);
or U1588 (N_1588,N_987,N_1417);
or U1589 (N_1589,N_1398,N_1498);
nand U1590 (N_1590,N_1243,N_771);
or U1591 (N_1591,N_1354,N_1225);
nand U1592 (N_1592,N_1431,N_947);
or U1593 (N_1593,N_1236,N_1240);
or U1594 (N_1594,N_1445,N_913);
nand U1595 (N_1595,N_1014,N_832);
and U1596 (N_1596,N_884,N_1095);
nor U1597 (N_1597,N_1022,N_819);
nor U1598 (N_1598,N_932,N_1208);
and U1599 (N_1599,N_963,N_792);
nand U1600 (N_1600,N_1042,N_1182);
or U1601 (N_1601,N_945,N_1349);
nand U1602 (N_1602,N_1116,N_979);
and U1603 (N_1603,N_1215,N_984);
and U1604 (N_1604,N_1013,N_960);
or U1605 (N_1605,N_928,N_1210);
nor U1606 (N_1606,N_1357,N_860);
and U1607 (N_1607,N_1121,N_1406);
or U1608 (N_1608,N_1132,N_1090);
nor U1609 (N_1609,N_1075,N_1481);
nand U1610 (N_1610,N_1017,N_1004);
and U1611 (N_1611,N_1322,N_1031);
nand U1612 (N_1612,N_848,N_1246);
nand U1613 (N_1613,N_1272,N_1294);
or U1614 (N_1614,N_1110,N_1386);
nand U1615 (N_1615,N_750,N_1310);
nor U1616 (N_1616,N_843,N_1424);
and U1617 (N_1617,N_1377,N_944);
or U1618 (N_1618,N_1054,N_1163);
and U1619 (N_1619,N_1043,N_1422);
and U1620 (N_1620,N_1065,N_999);
and U1621 (N_1621,N_808,N_1477);
and U1622 (N_1622,N_1051,N_1305);
and U1623 (N_1623,N_898,N_1205);
or U1624 (N_1624,N_989,N_1425);
nand U1625 (N_1625,N_1487,N_894);
and U1626 (N_1626,N_1267,N_1072);
or U1627 (N_1627,N_1192,N_1097);
or U1628 (N_1628,N_956,N_938);
nor U1629 (N_1629,N_1399,N_1428);
or U1630 (N_1630,N_1037,N_1282);
nand U1631 (N_1631,N_1480,N_769);
nor U1632 (N_1632,N_1411,N_974);
nor U1633 (N_1633,N_1370,N_935);
nand U1634 (N_1634,N_939,N_1066);
and U1635 (N_1635,N_1346,N_1449);
nor U1636 (N_1636,N_1474,N_1280);
nor U1637 (N_1637,N_1277,N_1160);
nand U1638 (N_1638,N_1062,N_1227);
or U1639 (N_1639,N_1047,N_1258);
and U1640 (N_1640,N_906,N_1155);
nor U1641 (N_1641,N_1146,N_1108);
nor U1642 (N_1642,N_934,N_930);
xnor U1643 (N_1643,N_1224,N_768);
nor U1644 (N_1644,N_948,N_1292);
or U1645 (N_1645,N_1057,N_790);
nor U1646 (N_1646,N_957,N_1207);
nand U1647 (N_1647,N_1053,N_802);
and U1648 (N_1648,N_857,N_1056);
and U1649 (N_1649,N_1120,N_1390);
nand U1650 (N_1650,N_1479,N_1029);
nor U1651 (N_1651,N_1492,N_924);
nand U1652 (N_1652,N_755,N_1143);
or U1653 (N_1653,N_788,N_1113);
nand U1654 (N_1654,N_1279,N_842);
and U1655 (N_1655,N_1329,N_885);
nor U1656 (N_1656,N_1125,N_976);
or U1657 (N_1657,N_1490,N_1301);
nand U1658 (N_1658,N_870,N_903);
nor U1659 (N_1659,N_831,N_1191);
nor U1660 (N_1660,N_1188,N_1382);
nand U1661 (N_1661,N_1307,N_993);
or U1662 (N_1662,N_1467,N_777);
and U1663 (N_1663,N_1247,N_775);
nor U1664 (N_1664,N_1459,N_1485);
nor U1665 (N_1665,N_910,N_996);
or U1666 (N_1666,N_1309,N_1164);
and U1667 (N_1667,N_798,N_856);
nand U1668 (N_1668,N_1218,N_1463);
and U1669 (N_1669,N_828,N_1287);
and U1670 (N_1670,N_1069,N_1130);
and U1671 (N_1671,N_1315,N_1470);
and U1672 (N_1672,N_1405,N_1252);
nand U1673 (N_1673,N_833,N_1298);
and U1674 (N_1674,N_795,N_1137);
nor U1675 (N_1675,N_818,N_760);
nand U1676 (N_1676,N_878,N_1226);
and U1677 (N_1677,N_1128,N_975);
nor U1678 (N_1678,N_1001,N_1134);
and U1679 (N_1679,N_951,N_1472);
and U1680 (N_1680,N_918,N_933);
and U1681 (N_1681,N_1300,N_1136);
nand U1682 (N_1682,N_1060,N_1184);
or U1683 (N_1683,N_1239,N_861);
nor U1684 (N_1684,N_805,N_1101);
nand U1685 (N_1685,N_1020,N_846);
and U1686 (N_1686,N_1288,N_897);
and U1687 (N_1687,N_959,N_994);
xor U1688 (N_1688,N_1093,N_972);
nor U1689 (N_1689,N_794,N_990);
and U1690 (N_1690,N_1395,N_907);
and U1691 (N_1691,N_1426,N_1087);
nor U1692 (N_1692,N_925,N_830);
xor U1693 (N_1693,N_1423,N_892);
nand U1694 (N_1694,N_1083,N_1145);
nand U1695 (N_1695,N_1438,N_1319);
and U1696 (N_1696,N_926,N_1166);
nand U1697 (N_1697,N_986,N_782);
or U1698 (N_1698,N_1318,N_895);
nand U1699 (N_1699,N_797,N_1266);
nand U1700 (N_1700,N_1235,N_1242);
and U1701 (N_1701,N_968,N_1413);
and U1702 (N_1702,N_1038,N_1385);
nand U1703 (N_1703,N_1450,N_1152);
or U1704 (N_1704,N_849,N_1456);
and U1705 (N_1705,N_1351,N_822);
xnor U1706 (N_1706,N_1233,N_1187);
nor U1707 (N_1707,N_1400,N_1437);
and U1708 (N_1708,N_1343,N_1402);
or U1709 (N_1709,N_1044,N_904);
nor U1710 (N_1710,N_950,N_852);
nor U1711 (N_1711,N_781,N_806);
nand U1712 (N_1712,N_905,N_763);
or U1713 (N_1713,N_1149,N_845);
nor U1714 (N_1714,N_762,N_1289);
or U1715 (N_1715,N_1353,N_1175);
or U1716 (N_1716,N_796,N_1165);
and U1717 (N_1717,N_1499,N_1064);
nand U1718 (N_1718,N_962,N_1050);
and U1719 (N_1719,N_1099,N_1000);
and U1720 (N_1720,N_1436,N_817);
and U1721 (N_1721,N_1036,N_859);
or U1722 (N_1722,N_1058,N_1473);
nor U1723 (N_1723,N_1347,N_1379);
and U1724 (N_1724,N_1341,N_1493);
and U1725 (N_1725,N_1002,N_1105);
nand U1726 (N_1726,N_1232,N_1147);
and U1727 (N_1727,N_1117,N_983);
xnor U1728 (N_1728,N_961,N_1404);
or U1729 (N_1729,N_1220,N_838);
nand U1730 (N_1730,N_1471,N_1460);
nand U1731 (N_1731,N_1323,N_936);
nor U1732 (N_1732,N_1348,N_1482);
nand U1733 (N_1733,N_1297,N_1034);
nand U1734 (N_1734,N_1414,N_872);
nand U1735 (N_1735,N_1180,N_1109);
nor U1736 (N_1736,N_1344,N_1167);
nand U1737 (N_1737,N_1096,N_1486);
nand U1738 (N_1738,N_1039,N_942);
nor U1739 (N_1739,N_1129,N_1352);
nor U1740 (N_1740,N_908,N_900);
xor U1741 (N_1741,N_753,N_1082);
or U1742 (N_1742,N_1229,N_1496);
and U1743 (N_1743,N_864,N_1290);
and U1744 (N_1744,N_804,N_1003);
nor U1745 (N_1745,N_1491,N_778);
nand U1746 (N_1746,N_1432,N_1257);
nand U1747 (N_1747,N_1212,N_840);
or U1748 (N_1748,N_1330,N_927);
nand U1749 (N_1749,N_1469,N_791);
and U1750 (N_1750,N_1055,N_1171);
and U1751 (N_1751,N_783,N_767);
or U1752 (N_1752,N_865,N_1118);
and U1753 (N_1753,N_1397,N_826);
and U1754 (N_1754,N_1387,N_1371);
nor U1755 (N_1755,N_1158,N_1336);
nand U1756 (N_1756,N_1126,N_1203);
nand U1757 (N_1757,N_866,N_1380);
or U1758 (N_1758,N_1306,N_770);
nand U1759 (N_1759,N_793,N_1157);
or U1760 (N_1760,N_765,N_1265);
and U1761 (N_1761,N_1433,N_787);
nor U1762 (N_1762,N_1412,N_1230);
nor U1763 (N_1763,N_807,N_886);
nor U1764 (N_1764,N_1074,N_889);
nor U1765 (N_1765,N_980,N_1360);
or U1766 (N_1766,N_756,N_915);
or U1767 (N_1767,N_929,N_851);
or U1768 (N_1768,N_1135,N_1332);
and U1769 (N_1769,N_998,N_1372);
nor U1770 (N_1770,N_1100,N_836);
and U1771 (N_1771,N_1048,N_995);
or U1772 (N_1772,N_1286,N_1447);
or U1773 (N_1773,N_1141,N_1421);
nor U1774 (N_1774,N_946,N_1388);
and U1775 (N_1775,N_1345,N_1367);
and U1776 (N_1776,N_779,N_1092);
and U1777 (N_1777,N_1019,N_1409);
nor U1778 (N_1778,N_1102,N_1262);
nor U1779 (N_1779,N_1026,N_981);
nor U1780 (N_1780,N_803,N_1464);
nand U1781 (N_1781,N_877,N_1320);
nor U1782 (N_1782,N_1324,N_1154);
nand U1783 (N_1783,N_786,N_1263);
xor U1784 (N_1784,N_1159,N_1144);
nand U1785 (N_1785,N_896,N_1080);
nor U1786 (N_1786,N_1112,N_893);
or U1787 (N_1787,N_809,N_1392);
and U1788 (N_1788,N_1441,N_1453);
and U1789 (N_1789,N_1389,N_964);
or U1790 (N_1790,N_1484,N_1374);
and U1791 (N_1791,N_1442,N_873);
xor U1792 (N_1792,N_965,N_1276);
nor U1793 (N_1793,N_1046,N_815);
and U1794 (N_1794,N_916,N_1098);
nor U1795 (N_1795,N_1337,N_888);
nand U1796 (N_1796,N_1359,N_1489);
or U1797 (N_1797,N_1006,N_1161);
nor U1798 (N_1798,N_1190,N_1222);
or U1799 (N_1799,N_1261,N_1316);
or U1800 (N_1800,N_1140,N_970);
nor U1801 (N_1801,N_1403,N_1179);
or U1802 (N_1802,N_1440,N_1494);
or U1803 (N_1803,N_1457,N_1488);
and U1804 (N_1804,N_1435,N_789);
xnor U1805 (N_1805,N_1071,N_883);
and U1806 (N_1806,N_1381,N_837);
nand U1807 (N_1807,N_1078,N_1430);
nor U1808 (N_1808,N_1077,N_774);
nor U1809 (N_1809,N_952,N_921);
and U1810 (N_1810,N_890,N_1314);
and U1811 (N_1811,N_1012,N_977);
nor U1812 (N_1812,N_814,N_1032);
nand U1813 (N_1813,N_1275,N_919);
nand U1814 (N_1814,N_1178,N_1452);
nand U1815 (N_1815,N_1304,N_1033);
xor U1816 (N_1816,N_1114,N_1018);
nand U1817 (N_1817,N_1408,N_874);
and U1818 (N_1818,N_1173,N_1350);
or U1819 (N_1819,N_812,N_991);
and U1820 (N_1820,N_1244,N_835);
or U1821 (N_1821,N_1260,N_751);
or U1822 (N_1822,N_1059,N_1384);
and U1823 (N_1823,N_1251,N_1209);
or U1824 (N_1824,N_1123,N_1063);
nor U1825 (N_1825,N_1273,N_1296);
nand U1826 (N_1826,N_880,N_1255);
or U1827 (N_1827,N_1429,N_937);
and U1828 (N_1828,N_1091,N_1076);
nor U1829 (N_1829,N_850,N_1461);
or U1830 (N_1830,N_773,N_1364);
nor U1831 (N_1831,N_1256,N_1302);
nor U1832 (N_1832,N_1326,N_1216);
nand U1833 (N_1833,N_1086,N_911);
nor U1834 (N_1834,N_1419,N_869);
or U1835 (N_1835,N_1131,N_1462);
nand U1836 (N_1836,N_1312,N_1451);
or U1837 (N_1837,N_1196,N_1495);
or U1838 (N_1838,N_1369,N_827);
or U1839 (N_1839,N_1183,N_1122);
and U1840 (N_1840,N_1250,N_1219);
and U1841 (N_1841,N_1138,N_1325);
nand U1842 (N_1842,N_1355,N_1234);
and U1843 (N_1843,N_862,N_1375);
or U1844 (N_1844,N_1253,N_912);
and U1845 (N_1845,N_1383,N_1313);
nor U1846 (N_1846,N_1317,N_887);
and U1847 (N_1847,N_761,N_1070);
nor U1848 (N_1848,N_1497,N_1271);
nand U1849 (N_1849,N_1221,N_1104);
nor U1850 (N_1850,N_969,N_1142);
nor U1851 (N_1851,N_1035,N_759);
xnor U1852 (N_1852,N_1393,N_1049);
or U1853 (N_1853,N_1466,N_1455);
nand U1854 (N_1854,N_839,N_1339);
or U1855 (N_1855,N_1231,N_754);
nand U1856 (N_1856,N_824,N_1181);
or U1857 (N_1857,N_1197,N_1270);
nand U1858 (N_1858,N_1139,N_1007);
and U1859 (N_1859,N_1259,N_799);
and U1860 (N_1860,N_1200,N_914);
or U1861 (N_1861,N_829,N_1274);
and U1862 (N_1862,N_1342,N_1358);
or U1863 (N_1863,N_949,N_1177);
or U1864 (N_1864,N_1174,N_858);
nand U1865 (N_1865,N_868,N_1361);
or U1866 (N_1866,N_1303,N_943);
and U1867 (N_1867,N_1238,N_966);
nand U1868 (N_1868,N_1150,N_1283);
nand U1869 (N_1869,N_776,N_1328);
and U1870 (N_1870,N_1396,N_1168);
or U1871 (N_1871,N_1458,N_1211);
nand U1872 (N_1872,N_1199,N_1415);
nor U1873 (N_1873,N_1103,N_1214);
and U1874 (N_1874,N_1416,N_784);
and U1875 (N_1875,N_1020,N_1425);
nor U1876 (N_1876,N_1045,N_1352);
nor U1877 (N_1877,N_812,N_1150);
or U1878 (N_1878,N_838,N_970);
nor U1879 (N_1879,N_1055,N_1297);
nor U1880 (N_1880,N_988,N_856);
and U1881 (N_1881,N_1134,N_757);
or U1882 (N_1882,N_1158,N_1126);
nor U1883 (N_1883,N_1303,N_1176);
nand U1884 (N_1884,N_1013,N_1349);
and U1885 (N_1885,N_900,N_1213);
nor U1886 (N_1886,N_1394,N_1281);
nor U1887 (N_1887,N_948,N_781);
nand U1888 (N_1888,N_873,N_1491);
or U1889 (N_1889,N_1003,N_1026);
and U1890 (N_1890,N_784,N_983);
and U1891 (N_1891,N_1360,N_984);
and U1892 (N_1892,N_1242,N_1088);
and U1893 (N_1893,N_1333,N_1289);
xnor U1894 (N_1894,N_1157,N_840);
or U1895 (N_1895,N_1368,N_804);
or U1896 (N_1896,N_784,N_1489);
nor U1897 (N_1897,N_855,N_1220);
or U1898 (N_1898,N_1259,N_1014);
or U1899 (N_1899,N_829,N_806);
or U1900 (N_1900,N_783,N_807);
and U1901 (N_1901,N_854,N_1146);
or U1902 (N_1902,N_1111,N_855);
xnor U1903 (N_1903,N_986,N_1176);
nand U1904 (N_1904,N_940,N_1364);
and U1905 (N_1905,N_925,N_1134);
or U1906 (N_1906,N_1225,N_846);
and U1907 (N_1907,N_982,N_1014);
nand U1908 (N_1908,N_1035,N_1000);
nand U1909 (N_1909,N_1491,N_1036);
nor U1910 (N_1910,N_1011,N_1158);
nor U1911 (N_1911,N_1012,N_876);
nor U1912 (N_1912,N_1101,N_1375);
nand U1913 (N_1913,N_1024,N_1375);
or U1914 (N_1914,N_926,N_1460);
nor U1915 (N_1915,N_1449,N_1407);
or U1916 (N_1916,N_795,N_879);
or U1917 (N_1917,N_1238,N_924);
nor U1918 (N_1918,N_1454,N_761);
or U1919 (N_1919,N_1285,N_1083);
and U1920 (N_1920,N_861,N_1151);
or U1921 (N_1921,N_787,N_978);
nor U1922 (N_1922,N_1426,N_1061);
nor U1923 (N_1923,N_1243,N_943);
and U1924 (N_1924,N_1453,N_1397);
and U1925 (N_1925,N_1081,N_1458);
nor U1926 (N_1926,N_1498,N_805);
nand U1927 (N_1927,N_1078,N_1377);
nand U1928 (N_1928,N_1052,N_1348);
nor U1929 (N_1929,N_1201,N_936);
nand U1930 (N_1930,N_1471,N_1031);
and U1931 (N_1931,N_1281,N_1284);
or U1932 (N_1932,N_1272,N_1113);
nand U1933 (N_1933,N_1338,N_1094);
and U1934 (N_1934,N_1455,N_1109);
and U1935 (N_1935,N_1365,N_1325);
and U1936 (N_1936,N_1374,N_1252);
nor U1937 (N_1937,N_1251,N_870);
nor U1938 (N_1938,N_1271,N_1214);
or U1939 (N_1939,N_1013,N_1205);
or U1940 (N_1940,N_767,N_1180);
nand U1941 (N_1941,N_1408,N_1336);
and U1942 (N_1942,N_1345,N_1300);
nor U1943 (N_1943,N_1165,N_968);
and U1944 (N_1944,N_1447,N_891);
or U1945 (N_1945,N_1340,N_1137);
xnor U1946 (N_1946,N_766,N_1026);
and U1947 (N_1947,N_1255,N_1401);
nor U1948 (N_1948,N_1381,N_1328);
nor U1949 (N_1949,N_831,N_1473);
nor U1950 (N_1950,N_1316,N_1240);
and U1951 (N_1951,N_876,N_919);
or U1952 (N_1952,N_1165,N_1153);
nor U1953 (N_1953,N_754,N_805);
and U1954 (N_1954,N_1336,N_1135);
nor U1955 (N_1955,N_1010,N_1245);
or U1956 (N_1956,N_984,N_1279);
or U1957 (N_1957,N_982,N_1465);
nor U1958 (N_1958,N_1496,N_1198);
or U1959 (N_1959,N_1280,N_1084);
or U1960 (N_1960,N_924,N_1241);
or U1961 (N_1961,N_910,N_1160);
nor U1962 (N_1962,N_1167,N_967);
nand U1963 (N_1963,N_1172,N_1245);
nand U1964 (N_1964,N_1005,N_1487);
nor U1965 (N_1965,N_1198,N_1294);
or U1966 (N_1966,N_762,N_1414);
nand U1967 (N_1967,N_817,N_1367);
nand U1968 (N_1968,N_1375,N_1436);
nand U1969 (N_1969,N_1078,N_1191);
or U1970 (N_1970,N_1141,N_1462);
nor U1971 (N_1971,N_1414,N_1392);
nor U1972 (N_1972,N_938,N_950);
or U1973 (N_1973,N_917,N_803);
or U1974 (N_1974,N_895,N_840);
and U1975 (N_1975,N_816,N_1234);
or U1976 (N_1976,N_913,N_799);
nand U1977 (N_1977,N_755,N_1334);
nor U1978 (N_1978,N_1093,N_768);
nand U1979 (N_1979,N_827,N_977);
and U1980 (N_1980,N_895,N_757);
or U1981 (N_1981,N_1419,N_856);
nor U1982 (N_1982,N_1001,N_1198);
nor U1983 (N_1983,N_1023,N_969);
nand U1984 (N_1984,N_967,N_1212);
nand U1985 (N_1985,N_970,N_1114);
nor U1986 (N_1986,N_1074,N_791);
nand U1987 (N_1987,N_1073,N_766);
nand U1988 (N_1988,N_944,N_1154);
or U1989 (N_1989,N_853,N_928);
and U1990 (N_1990,N_772,N_1070);
and U1991 (N_1991,N_1136,N_1050);
nor U1992 (N_1992,N_872,N_1103);
nor U1993 (N_1993,N_1050,N_772);
or U1994 (N_1994,N_874,N_1362);
nand U1995 (N_1995,N_884,N_1362);
nand U1996 (N_1996,N_925,N_953);
and U1997 (N_1997,N_1223,N_1132);
nand U1998 (N_1998,N_987,N_1146);
or U1999 (N_1999,N_1047,N_1421);
and U2000 (N_2000,N_1313,N_1421);
and U2001 (N_2001,N_1049,N_1374);
nand U2002 (N_2002,N_1434,N_1364);
nor U2003 (N_2003,N_1358,N_812);
and U2004 (N_2004,N_778,N_991);
nand U2005 (N_2005,N_924,N_1408);
nor U2006 (N_2006,N_1393,N_759);
xor U2007 (N_2007,N_961,N_1196);
nand U2008 (N_2008,N_840,N_792);
or U2009 (N_2009,N_759,N_893);
nor U2010 (N_2010,N_813,N_810);
and U2011 (N_2011,N_1148,N_1182);
nand U2012 (N_2012,N_1322,N_1081);
nand U2013 (N_2013,N_1015,N_1117);
or U2014 (N_2014,N_961,N_1043);
nand U2015 (N_2015,N_1105,N_1336);
nor U2016 (N_2016,N_1239,N_1085);
nor U2017 (N_2017,N_947,N_1238);
and U2018 (N_2018,N_860,N_1473);
or U2019 (N_2019,N_797,N_875);
or U2020 (N_2020,N_1149,N_1457);
nand U2021 (N_2021,N_1466,N_1378);
or U2022 (N_2022,N_820,N_1341);
nand U2023 (N_2023,N_1457,N_853);
or U2024 (N_2024,N_1168,N_1277);
nand U2025 (N_2025,N_972,N_1102);
and U2026 (N_2026,N_788,N_1274);
nand U2027 (N_2027,N_787,N_1401);
nor U2028 (N_2028,N_1354,N_1307);
and U2029 (N_2029,N_1404,N_1031);
or U2030 (N_2030,N_1119,N_851);
and U2031 (N_2031,N_1451,N_1230);
xnor U2032 (N_2032,N_825,N_1302);
nand U2033 (N_2033,N_1065,N_1279);
and U2034 (N_2034,N_919,N_877);
nor U2035 (N_2035,N_751,N_1154);
nand U2036 (N_2036,N_1028,N_1437);
nand U2037 (N_2037,N_755,N_1234);
nor U2038 (N_2038,N_1411,N_807);
and U2039 (N_2039,N_1111,N_1309);
nand U2040 (N_2040,N_1132,N_1157);
and U2041 (N_2041,N_960,N_1281);
or U2042 (N_2042,N_767,N_1404);
nor U2043 (N_2043,N_957,N_1470);
nor U2044 (N_2044,N_871,N_792);
and U2045 (N_2045,N_1446,N_1387);
nor U2046 (N_2046,N_1211,N_1104);
and U2047 (N_2047,N_1046,N_1065);
and U2048 (N_2048,N_1380,N_1393);
nand U2049 (N_2049,N_797,N_808);
and U2050 (N_2050,N_1156,N_1279);
and U2051 (N_2051,N_834,N_960);
and U2052 (N_2052,N_949,N_785);
nand U2053 (N_2053,N_1396,N_1006);
or U2054 (N_2054,N_820,N_1186);
nand U2055 (N_2055,N_1310,N_1491);
nand U2056 (N_2056,N_1032,N_1142);
or U2057 (N_2057,N_815,N_1320);
nand U2058 (N_2058,N_1030,N_927);
nor U2059 (N_2059,N_1182,N_1184);
and U2060 (N_2060,N_1125,N_778);
nor U2061 (N_2061,N_1231,N_955);
nand U2062 (N_2062,N_783,N_1022);
or U2063 (N_2063,N_1211,N_779);
nor U2064 (N_2064,N_1052,N_1112);
and U2065 (N_2065,N_789,N_1062);
and U2066 (N_2066,N_1071,N_1362);
nand U2067 (N_2067,N_1002,N_1201);
and U2068 (N_2068,N_846,N_1143);
nor U2069 (N_2069,N_1202,N_998);
xnor U2070 (N_2070,N_1397,N_1266);
and U2071 (N_2071,N_1203,N_781);
and U2072 (N_2072,N_1094,N_1329);
or U2073 (N_2073,N_1254,N_827);
and U2074 (N_2074,N_1149,N_775);
or U2075 (N_2075,N_1422,N_1007);
and U2076 (N_2076,N_1149,N_1121);
or U2077 (N_2077,N_810,N_801);
nor U2078 (N_2078,N_914,N_918);
nand U2079 (N_2079,N_1307,N_1398);
nand U2080 (N_2080,N_1495,N_985);
nand U2081 (N_2081,N_929,N_1299);
nand U2082 (N_2082,N_1129,N_1255);
and U2083 (N_2083,N_1087,N_977);
and U2084 (N_2084,N_940,N_1466);
and U2085 (N_2085,N_1223,N_799);
and U2086 (N_2086,N_1397,N_1383);
nor U2087 (N_2087,N_1091,N_1206);
nand U2088 (N_2088,N_885,N_1430);
nor U2089 (N_2089,N_783,N_1097);
nand U2090 (N_2090,N_1418,N_854);
xor U2091 (N_2091,N_1498,N_1009);
or U2092 (N_2092,N_1187,N_1238);
nor U2093 (N_2093,N_913,N_1078);
nor U2094 (N_2094,N_1256,N_895);
or U2095 (N_2095,N_837,N_764);
and U2096 (N_2096,N_1451,N_1044);
and U2097 (N_2097,N_1427,N_1008);
or U2098 (N_2098,N_1342,N_1165);
nand U2099 (N_2099,N_761,N_1118);
or U2100 (N_2100,N_1364,N_1201);
and U2101 (N_2101,N_1177,N_959);
or U2102 (N_2102,N_1236,N_1467);
nand U2103 (N_2103,N_1195,N_1406);
xor U2104 (N_2104,N_1498,N_1458);
nand U2105 (N_2105,N_889,N_1235);
nand U2106 (N_2106,N_1416,N_1338);
and U2107 (N_2107,N_1169,N_1156);
nor U2108 (N_2108,N_1225,N_811);
nand U2109 (N_2109,N_913,N_1326);
nor U2110 (N_2110,N_831,N_1238);
and U2111 (N_2111,N_765,N_1318);
xnor U2112 (N_2112,N_1063,N_1194);
and U2113 (N_2113,N_762,N_1026);
or U2114 (N_2114,N_1156,N_1163);
xnor U2115 (N_2115,N_1073,N_1034);
nor U2116 (N_2116,N_875,N_898);
nand U2117 (N_2117,N_1042,N_803);
nor U2118 (N_2118,N_926,N_1396);
nand U2119 (N_2119,N_1035,N_929);
nor U2120 (N_2120,N_979,N_1248);
or U2121 (N_2121,N_1113,N_1038);
or U2122 (N_2122,N_1176,N_1448);
xor U2123 (N_2123,N_764,N_758);
and U2124 (N_2124,N_842,N_1229);
nand U2125 (N_2125,N_1173,N_1170);
and U2126 (N_2126,N_1337,N_1413);
and U2127 (N_2127,N_1171,N_1411);
and U2128 (N_2128,N_1163,N_1157);
nand U2129 (N_2129,N_905,N_1258);
nor U2130 (N_2130,N_1051,N_982);
nor U2131 (N_2131,N_1327,N_1392);
or U2132 (N_2132,N_1358,N_1062);
xor U2133 (N_2133,N_1064,N_1246);
nand U2134 (N_2134,N_815,N_1345);
nor U2135 (N_2135,N_1465,N_836);
xor U2136 (N_2136,N_947,N_882);
nand U2137 (N_2137,N_880,N_1241);
nor U2138 (N_2138,N_841,N_927);
and U2139 (N_2139,N_1495,N_907);
nor U2140 (N_2140,N_1325,N_1157);
nand U2141 (N_2141,N_794,N_1067);
or U2142 (N_2142,N_1488,N_1176);
nand U2143 (N_2143,N_1104,N_1102);
and U2144 (N_2144,N_830,N_1140);
nor U2145 (N_2145,N_1495,N_1005);
and U2146 (N_2146,N_1270,N_1116);
or U2147 (N_2147,N_766,N_810);
nand U2148 (N_2148,N_1040,N_1164);
and U2149 (N_2149,N_850,N_1083);
nor U2150 (N_2150,N_1328,N_1005);
nand U2151 (N_2151,N_1069,N_877);
and U2152 (N_2152,N_814,N_787);
nor U2153 (N_2153,N_957,N_905);
nand U2154 (N_2154,N_1456,N_1054);
nor U2155 (N_2155,N_1358,N_1340);
or U2156 (N_2156,N_893,N_1370);
nand U2157 (N_2157,N_962,N_1070);
nor U2158 (N_2158,N_1439,N_1222);
nand U2159 (N_2159,N_1016,N_908);
nand U2160 (N_2160,N_1367,N_1152);
nand U2161 (N_2161,N_1089,N_1182);
nand U2162 (N_2162,N_1164,N_987);
nand U2163 (N_2163,N_785,N_935);
or U2164 (N_2164,N_1085,N_1016);
nor U2165 (N_2165,N_1108,N_1310);
or U2166 (N_2166,N_1474,N_1098);
and U2167 (N_2167,N_1380,N_1377);
or U2168 (N_2168,N_997,N_1151);
nand U2169 (N_2169,N_1270,N_1461);
nor U2170 (N_2170,N_1253,N_1011);
and U2171 (N_2171,N_981,N_1497);
nand U2172 (N_2172,N_885,N_1224);
nor U2173 (N_2173,N_1337,N_1102);
nor U2174 (N_2174,N_1042,N_828);
nor U2175 (N_2175,N_1154,N_991);
nor U2176 (N_2176,N_1164,N_896);
nand U2177 (N_2177,N_757,N_1192);
nor U2178 (N_2178,N_841,N_906);
or U2179 (N_2179,N_796,N_958);
and U2180 (N_2180,N_1081,N_1216);
nand U2181 (N_2181,N_1349,N_834);
or U2182 (N_2182,N_917,N_1320);
and U2183 (N_2183,N_1477,N_799);
nor U2184 (N_2184,N_1129,N_757);
nor U2185 (N_2185,N_1237,N_772);
nor U2186 (N_2186,N_764,N_1126);
or U2187 (N_2187,N_1228,N_976);
nand U2188 (N_2188,N_976,N_1062);
and U2189 (N_2189,N_1350,N_774);
and U2190 (N_2190,N_1242,N_1110);
and U2191 (N_2191,N_963,N_1459);
or U2192 (N_2192,N_903,N_1093);
nand U2193 (N_2193,N_931,N_1323);
nand U2194 (N_2194,N_1133,N_1249);
and U2195 (N_2195,N_1169,N_1086);
and U2196 (N_2196,N_1257,N_1397);
nand U2197 (N_2197,N_1171,N_970);
and U2198 (N_2198,N_1179,N_1017);
and U2199 (N_2199,N_1406,N_1099);
nand U2200 (N_2200,N_866,N_947);
or U2201 (N_2201,N_895,N_850);
xnor U2202 (N_2202,N_1448,N_1064);
and U2203 (N_2203,N_1406,N_1101);
or U2204 (N_2204,N_1447,N_1135);
or U2205 (N_2205,N_1331,N_1296);
and U2206 (N_2206,N_1033,N_853);
nor U2207 (N_2207,N_1242,N_945);
nor U2208 (N_2208,N_1229,N_926);
nand U2209 (N_2209,N_987,N_1292);
or U2210 (N_2210,N_1301,N_784);
or U2211 (N_2211,N_1089,N_1497);
and U2212 (N_2212,N_1047,N_1392);
nor U2213 (N_2213,N_987,N_781);
nor U2214 (N_2214,N_1199,N_1098);
and U2215 (N_2215,N_1025,N_1353);
and U2216 (N_2216,N_1061,N_1045);
xnor U2217 (N_2217,N_1325,N_1014);
or U2218 (N_2218,N_1224,N_1423);
and U2219 (N_2219,N_1124,N_820);
and U2220 (N_2220,N_979,N_863);
nand U2221 (N_2221,N_1143,N_1024);
and U2222 (N_2222,N_980,N_1392);
and U2223 (N_2223,N_1106,N_1172);
or U2224 (N_2224,N_916,N_755);
and U2225 (N_2225,N_951,N_1150);
and U2226 (N_2226,N_805,N_865);
nor U2227 (N_2227,N_989,N_1403);
or U2228 (N_2228,N_781,N_849);
nor U2229 (N_2229,N_895,N_1163);
nand U2230 (N_2230,N_1435,N_778);
nor U2231 (N_2231,N_1322,N_1484);
nand U2232 (N_2232,N_874,N_955);
or U2233 (N_2233,N_1332,N_815);
nand U2234 (N_2234,N_1269,N_1104);
or U2235 (N_2235,N_833,N_1338);
and U2236 (N_2236,N_1300,N_1483);
nand U2237 (N_2237,N_920,N_1133);
nor U2238 (N_2238,N_864,N_890);
and U2239 (N_2239,N_1291,N_786);
or U2240 (N_2240,N_1127,N_1344);
nor U2241 (N_2241,N_1041,N_1336);
or U2242 (N_2242,N_1118,N_1249);
or U2243 (N_2243,N_804,N_1047);
nor U2244 (N_2244,N_914,N_1390);
nand U2245 (N_2245,N_1323,N_1184);
nor U2246 (N_2246,N_958,N_1300);
nand U2247 (N_2247,N_894,N_801);
xor U2248 (N_2248,N_998,N_802);
xnor U2249 (N_2249,N_937,N_765);
and U2250 (N_2250,N_1790,N_2230);
xnor U2251 (N_2251,N_1521,N_1843);
or U2252 (N_2252,N_2199,N_2012);
nor U2253 (N_2253,N_1886,N_1771);
nor U2254 (N_2254,N_1587,N_2138);
or U2255 (N_2255,N_2167,N_2223);
xnor U2256 (N_2256,N_2202,N_2131);
or U2257 (N_2257,N_1541,N_1702);
nor U2258 (N_2258,N_2150,N_1750);
nor U2259 (N_2259,N_1980,N_2044);
nand U2260 (N_2260,N_1954,N_1532);
and U2261 (N_2261,N_1503,N_2217);
nand U2262 (N_2262,N_2075,N_1996);
xnor U2263 (N_2263,N_1549,N_2218);
or U2264 (N_2264,N_1709,N_1870);
and U2265 (N_2265,N_2105,N_2060);
or U2266 (N_2266,N_2221,N_1792);
nand U2267 (N_2267,N_2233,N_1795);
nand U2268 (N_2268,N_2173,N_1791);
and U2269 (N_2269,N_2224,N_1612);
nand U2270 (N_2270,N_1669,N_2078);
or U2271 (N_2271,N_1995,N_2137);
xor U2272 (N_2272,N_2245,N_1821);
nor U2273 (N_2273,N_1674,N_1559);
and U2274 (N_2274,N_1933,N_1845);
nand U2275 (N_2275,N_2070,N_1751);
nor U2276 (N_2276,N_2094,N_2184);
and U2277 (N_2277,N_1544,N_1606);
xnor U2278 (N_2278,N_2031,N_1682);
nand U2279 (N_2279,N_1923,N_1912);
xnor U2280 (N_2280,N_1951,N_1648);
or U2281 (N_2281,N_1830,N_1784);
nor U2282 (N_2282,N_1740,N_1525);
nor U2283 (N_2283,N_2166,N_2144);
and U2284 (N_2284,N_1691,N_1676);
or U2285 (N_2285,N_2129,N_1734);
nor U2286 (N_2286,N_2093,N_1937);
or U2287 (N_2287,N_1839,N_1572);
or U2288 (N_2288,N_1566,N_2182);
or U2289 (N_2289,N_2063,N_2164);
nand U2290 (N_2290,N_1965,N_1852);
and U2291 (N_2291,N_1949,N_2151);
or U2292 (N_2292,N_1584,N_2141);
nor U2293 (N_2293,N_1514,N_1862);
and U2294 (N_2294,N_1553,N_1938);
nand U2295 (N_2295,N_1913,N_1901);
and U2296 (N_2296,N_1652,N_1992);
nand U2297 (N_2297,N_1573,N_1962);
and U2298 (N_2298,N_1890,N_1947);
nor U2299 (N_2299,N_1959,N_2046);
xor U2300 (N_2300,N_1783,N_1785);
or U2301 (N_2301,N_2118,N_2187);
nor U2302 (N_2302,N_1766,N_1920);
nand U2303 (N_2303,N_1824,N_1581);
nand U2304 (N_2304,N_1643,N_2237);
nand U2305 (N_2305,N_1671,N_2239);
or U2306 (N_2306,N_2027,N_1561);
or U2307 (N_2307,N_2020,N_1769);
nand U2308 (N_2308,N_1952,N_1958);
and U2309 (N_2309,N_2231,N_2103);
xor U2310 (N_2310,N_1859,N_1687);
and U2311 (N_2311,N_1898,N_2128);
nor U2312 (N_2312,N_1893,N_1582);
and U2313 (N_2313,N_1679,N_1774);
nor U2314 (N_2314,N_1689,N_2039);
nand U2315 (N_2315,N_1626,N_2073);
or U2316 (N_2316,N_1803,N_1723);
and U2317 (N_2317,N_2148,N_1835);
nand U2318 (N_2318,N_1999,N_1720);
and U2319 (N_2319,N_2069,N_1555);
nor U2320 (N_2320,N_1888,N_1595);
xor U2321 (N_2321,N_1925,N_1737);
nor U2322 (N_2322,N_2168,N_1801);
and U2323 (N_2323,N_2076,N_1660);
nor U2324 (N_2324,N_1551,N_1724);
and U2325 (N_2325,N_1617,N_1787);
and U2326 (N_2326,N_1873,N_1825);
nor U2327 (N_2327,N_1861,N_1904);
nand U2328 (N_2328,N_1994,N_1692);
or U2329 (N_2329,N_1611,N_1736);
or U2330 (N_2330,N_1700,N_2127);
nand U2331 (N_2331,N_1817,N_1694);
and U2332 (N_2332,N_2211,N_1563);
nand U2333 (N_2333,N_1810,N_2000);
and U2334 (N_2334,N_1748,N_1654);
nand U2335 (N_2335,N_1819,N_1984);
or U2336 (N_2336,N_1823,N_2049);
nor U2337 (N_2337,N_1688,N_1761);
or U2338 (N_2338,N_2159,N_1616);
and U2339 (N_2339,N_2102,N_2149);
nor U2340 (N_2340,N_1829,N_2024);
and U2341 (N_2341,N_2050,N_1746);
and U2342 (N_2342,N_1697,N_2232);
nor U2343 (N_2343,N_1666,N_2117);
or U2344 (N_2344,N_2064,N_1762);
and U2345 (N_2345,N_1653,N_1630);
and U2346 (N_2346,N_1779,N_2214);
or U2347 (N_2347,N_1754,N_1850);
or U2348 (N_2348,N_1647,N_1625);
nand U2349 (N_2349,N_2037,N_1699);
nor U2350 (N_2350,N_1812,N_1698);
nor U2351 (N_2351,N_2162,N_1714);
nor U2352 (N_2352,N_2215,N_1828);
nor U2353 (N_2353,N_1855,N_1877);
or U2354 (N_2354,N_1781,N_1858);
and U2355 (N_2355,N_2013,N_1554);
and U2356 (N_2356,N_1849,N_2241);
nor U2357 (N_2357,N_2190,N_2018);
or U2358 (N_2358,N_1908,N_1928);
nand U2359 (N_2359,N_1944,N_2043);
nor U2360 (N_2360,N_2176,N_1827);
nor U2361 (N_2361,N_1657,N_2210);
nor U2362 (N_2362,N_1583,N_1664);
nand U2363 (N_2363,N_1523,N_1507);
nand U2364 (N_2364,N_1622,N_2236);
or U2365 (N_2365,N_1650,N_1872);
nand U2366 (N_2366,N_1651,N_2116);
nand U2367 (N_2367,N_2066,N_1887);
xor U2368 (N_2368,N_2101,N_1518);
nor U2369 (N_2369,N_1897,N_1929);
nor U2370 (N_2370,N_1602,N_2071);
nand U2371 (N_2371,N_1537,N_2008);
or U2372 (N_2372,N_2216,N_1655);
nand U2373 (N_2373,N_1701,N_2225);
and U2374 (N_2374,N_1706,N_1725);
and U2375 (N_2375,N_1517,N_1597);
nand U2376 (N_2376,N_2189,N_1976);
or U2377 (N_2377,N_1605,N_1543);
or U2378 (N_2378,N_1987,N_1970);
nor U2379 (N_2379,N_2068,N_1867);
nand U2380 (N_2380,N_2041,N_1799);
or U2381 (N_2381,N_1631,N_1600);
nor U2382 (N_2382,N_2026,N_2004);
and U2383 (N_2383,N_1826,N_2002);
and U2384 (N_2384,N_2157,N_1816);
and U2385 (N_2385,N_1534,N_2047);
nor U2386 (N_2386,N_1550,N_1708);
nand U2387 (N_2387,N_2015,N_1627);
xor U2388 (N_2388,N_2086,N_1950);
and U2389 (N_2389,N_1747,N_1842);
and U2390 (N_2390,N_1636,N_1865);
or U2391 (N_2391,N_2001,N_1895);
nand U2392 (N_2392,N_1713,N_2130);
nor U2393 (N_2393,N_1501,N_1834);
or U2394 (N_2394,N_1820,N_2053);
nor U2395 (N_2395,N_1509,N_1807);
nor U2396 (N_2396,N_1538,N_1763);
or U2397 (N_2397,N_1866,N_2121);
and U2398 (N_2398,N_1990,N_2247);
nor U2399 (N_2399,N_2192,N_2052);
or U2400 (N_2400,N_2055,N_2096);
and U2401 (N_2401,N_2212,N_2005);
and U2402 (N_2402,N_1545,N_1571);
nand U2403 (N_2403,N_1782,N_1863);
and U2404 (N_2404,N_1608,N_1633);
and U2405 (N_2405,N_1985,N_1506);
xnor U2406 (N_2406,N_2206,N_1847);
and U2407 (N_2407,N_1967,N_1978);
nor U2408 (N_2408,N_2054,N_1732);
and U2409 (N_2409,N_1936,N_1715);
or U2410 (N_2410,N_1607,N_1742);
nand U2411 (N_2411,N_2126,N_2133);
nor U2412 (N_2412,N_2109,N_1739);
nand U2413 (N_2413,N_1589,N_1993);
or U2414 (N_2414,N_1749,N_2185);
and U2415 (N_2415,N_1946,N_1562);
nor U2416 (N_2416,N_1530,N_2034);
nand U2417 (N_2417,N_1510,N_2081);
nor U2418 (N_2418,N_1695,N_1768);
nor U2419 (N_2419,N_1909,N_2095);
xnor U2420 (N_2420,N_1644,N_1975);
nand U2421 (N_2421,N_1727,N_2139);
nor U2422 (N_2422,N_1811,N_2025);
xnor U2423 (N_2423,N_2106,N_1690);
nor U2424 (N_2424,N_1634,N_1776);
and U2425 (N_2425,N_1599,N_1667);
nand U2426 (N_2426,N_1942,N_1729);
or U2427 (N_2427,N_2120,N_1880);
or U2428 (N_2428,N_2065,N_2119);
nand U2429 (N_2429,N_1922,N_2135);
nand U2430 (N_2430,N_2198,N_1693);
and U2431 (N_2431,N_2023,N_1528);
or U2432 (N_2432,N_1678,N_1618);
or U2433 (N_2433,N_2188,N_2136);
and U2434 (N_2434,N_2028,N_2006);
and U2435 (N_2435,N_1963,N_2074);
and U2436 (N_2436,N_1719,N_1902);
or U2437 (N_2437,N_1857,N_1527);
or U2438 (N_2438,N_2179,N_2194);
nand U2439 (N_2439,N_2249,N_1560);
nand U2440 (N_2440,N_1884,N_2227);
and U2441 (N_2441,N_1814,N_1759);
nor U2442 (N_2442,N_1540,N_1593);
nor U2443 (N_2443,N_2088,N_1542);
nand U2444 (N_2444,N_1973,N_1894);
or U2445 (N_2445,N_1773,N_2032);
nand U2446 (N_2446,N_1511,N_2110);
nand U2447 (N_2447,N_1539,N_2204);
nand U2448 (N_2448,N_2177,N_1683);
nand U2449 (N_2449,N_1670,N_1557);
nor U2450 (N_2450,N_2158,N_1753);
nand U2451 (N_2451,N_1752,N_2056);
nand U2452 (N_2452,N_1570,N_2042);
or U2453 (N_2453,N_1869,N_1743);
nor U2454 (N_2454,N_1956,N_1711);
or U2455 (N_2455,N_1638,N_2195);
and U2456 (N_2456,N_2080,N_1982);
or U2457 (N_2457,N_1778,N_1726);
and U2458 (N_2458,N_2170,N_2220);
and U2459 (N_2459,N_1519,N_1868);
nor U2460 (N_2460,N_2033,N_1645);
and U2461 (N_2461,N_1991,N_1649);
and U2462 (N_2462,N_1860,N_1900);
xor U2463 (N_2463,N_1755,N_2057);
nor U2464 (N_2464,N_1881,N_1558);
or U2465 (N_2465,N_1926,N_2238);
and U2466 (N_2466,N_1547,N_1885);
or U2467 (N_2467,N_1848,N_1939);
and U2468 (N_2468,N_2089,N_1822);
or U2469 (N_2469,N_1818,N_1610);
nor U2470 (N_2470,N_1960,N_2174);
and U2471 (N_2471,N_1705,N_2246);
and U2472 (N_2472,N_1662,N_1940);
and U2473 (N_2473,N_2040,N_1966);
and U2474 (N_2474,N_1896,N_1815);
or U2475 (N_2475,N_1601,N_2219);
nand U2476 (N_2476,N_1567,N_2207);
and U2477 (N_2477,N_1505,N_2067);
nor U2478 (N_2478,N_2156,N_1983);
or U2479 (N_2479,N_2208,N_1577);
nand U2480 (N_2480,N_2205,N_1906);
or U2481 (N_2481,N_2155,N_1831);
and U2482 (N_2482,N_2222,N_2123);
and U2483 (N_2483,N_1738,N_1998);
or U2484 (N_2484,N_1672,N_1640);
and U2485 (N_2485,N_1686,N_1961);
or U2486 (N_2486,N_2235,N_1813);
nand U2487 (N_2487,N_2193,N_1680);
and U2488 (N_2488,N_1879,N_1916);
and U2489 (N_2489,N_2108,N_2242);
nand U2490 (N_2490,N_1770,N_1878);
and U2491 (N_2491,N_2014,N_1721);
or U2492 (N_2492,N_2180,N_1837);
and U2493 (N_2493,N_1800,N_2243);
nor U2494 (N_2494,N_1722,N_2181);
nor U2495 (N_2495,N_1945,N_1556);
and U2496 (N_2496,N_2152,N_1793);
nand U2497 (N_2497,N_1535,N_2048);
and U2498 (N_2498,N_2240,N_1758);
nand U2499 (N_2499,N_2196,N_1892);
nor U2500 (N_2500,N_2175,N_1635);
nor U2501 (N_2501,N_1977,N_2009);
or U2502 (N_2502,N_2058,N_2079);
nor U2503 (N_2503,N_1846,N_2017);
nand U2504 (N_2504,N_1522,N_2111);
xnor U2505 (N_2505,N_2045,N_1716);
and U2506 (N_2506,N_2160,N_1665);
nor U2507 (N_2507,N_1911,N_2097);
nand U2508 (N_2508,N_1798,N_2124);
and U2509 (N_2509,N_1986,N_1564);
or U2510 (N_2510,N_1953,N_2010);
nand U2511 (N_2511,N_1574,N_1910);
or U2512 (N_2512,N_1552,N_1656);
and U2513 (N_2513,N_2143,N_1907);
nand U2514 (N_2514,N_1696,N_1931);
and U2515 (N_2515,N_1760,N_1780);
nand U2516 (N_2516,N_1915,N_1673);
or U2517 (N_2517,N_1590,N_1808);
or U2518 (N_2518,N_1579,N_1710);
nand U2519 (N_2519,N_1588,N_2113);
nor U2520 (N_2520,N_1943,N_1735);
nor U2521 (N_2521,N_2036,N_1851);
or U2522 (N_2522,N_2122,N_1621);
and U2523 (N_2523,N_1974,N_1924);
or U2524 (N_2524,N_1972,N_1917);
xnor U2525 (N_2525,N_2077,N_1874);
or U2526 (N_2526,N_1598,N_2016);
nor U2527 (N_2527,N_2092,N_1513);
nand U2528 (N_2528,N_1788,N_1596);
nand U2529 (N_2529,N_1903,N_1932);
nor U2530 (N_2530,N_2090,N_1809);
nand U2531 (N_2531,N_1764,N_1526);
nand U2532 (N_2532,N_1789,N_2087);
nor U2533 (N_2533,N_1615,N_2035);
and U2534 (N_2534,N_2145,N_2147);
nand U2535 (N_2535,N_1592,N_1632);
nor U2536 (N_2536,N_2234,N_1832);
nand U2537 (N_2537,N_1744,N_1875);
and U2538 (N_2538,N_1536,N_1745);
nor U2539 (N_2539,N_1524,N_1919);
nand U2540 (N_2540,N_2022,N_1585);
and U2541 (N_2541,N_1646,N_2115);
nand U2542 (N_2542,N_1969,N_2226);
and U2543 (N_2543,N_1717,N_1728);
nor U2544 (N_2544,N_2178,N_1568);
and U2545 (N_2545,N_2200,N_1957);
or U2546 (N_2546,N_1997,N_1914);
and U2547 (N_2547,N_2107,N_1731);
nor U2548 (N_2548,N_2134,N_1604);
nor U2549 (N_2549,N_1899,N_1575);
nand U2550 (N_2550,N_1704,N_1668);
and U2551 (N_2551,N_1854,N_1883);
nor U2552 (N_2552,N_1934,N_1979);
and U2553 (N_2553,N_1504,N_1756);
and U2554 (N_2554,N_2186,N_2244);
nand U2555 (N_2555,N_2209,N_1775);
and U2556 (N_2556,N_1594,N_2029);
and U2557 (N_2557,N_1772,N_1889);
nand U2558 (N_2558,N_1876,N_1637);
or U2559 (N_2559,N_1730,N_2172);
or U2560 (N_2560,N_2154,N_1629);
nor U2561 (N_2561,N_1712,N_2171);
and U2562 (N_2562,N_1804,N_1882);
and U2563 (N_2563,N_1981,N_2125);
nand U2564 (N_2564,N_1613,N_1703);
and U2565 (N_2565,N_1639,N_1641);
or U2566 (N_2566,N_1786,N_2161);
and U2567 (N_2567,N_1603,N_2112);
and U2568 (N_2568,N_2229,N_2007);
xnor U2569 (N_2569,N_1619,N_1891);
nor U2570 (N_2570,N_1733,N_2051);
and U2571 (N_2571,N_2132,N_1580);
or U2572 (N_2572,N_1757,N_2100);
and U2573 (N_2573,N_2061,N_1578);
and U2574 (N_2574,N_1586,N_1508);
and U2575 (N_2575,N_1591,N_1853);
or U2576 (N_2576,N_2062,N_2104);
or U2577 (N_2577,N_1905,N_1569);
and U2578 (N_2578,N_1623,N_2197);
or U2579 (N_2579,N_1948,N_2085);
nor U2580 (N_2580,N_2163,N_1659);
nor U2581 (N_2581,N_1658,N_2248);
or U2582 (N_2582,N_1841,N_2114);
nand U2583 (N_2583,N_1516,N_1806);
nor U2584 (N_2584,N_2003,N_2030);
or U2585 (N_2585,N_1515,N_2011);
or U2586 (N_2586,N_1968,N_2153);
nor U2587 (N_2587,N_1864,N_1805);
nor U2588 (N_2588,N_1765,N_2165);
or U2589 (N_2589,N_1988,N_1971);
and U2590 (N_2590,N_1844,N_1533);
or U2591 (N_2591,N_1796,N_1927);
nand U2592 (N_2592,N_2059,N_1833);
or U2593 (N_2593,N_2084,N_1794);
or U2594 (N_2594,N_1685,N_2201);
nand U2595 (N_2595,N_1767,N_1935);
nand U2596 (N_2596,N_1500,N_1856);
nand U2597 (N_2597,N_2142,N_2203);
nor U2598 (N_2598,N_2191,N_1548);
or U2599 (N_2599,N_1707,N_1512);
and U2600 (N_2600,N_2098,N_2083);
nand U2601 (N_2601,N_1871,N_1941);
xor U2602 (N_2602,N_2146,N_1502);
nor U2603 (N_2603,N_1642,N_1565);
nand U2604 (N_2604,N_1802,N_1663);
nor U2605 (N_2605,N_1930,N_1921);
and U2606 (N_2606,N_2038,N_1741);
nand U2607 (N_2607,N_2082,N_1609);
nor U2608 (N_2608,N_1684,N_1797);
or U2609 (N_2609,N_2228,N_1840);
or U2610 (N_2610,N_1628,N_1531);
nand U2611 (N_2611,N_2213,N_1677);
and U2612 (N_2612,N_1520,N_1777);
nand U2613 (N_2613,N_2019,N_2140);
nor U2614 (N_2614,N_1614,N_2021);
nand U2615 (N_2615,N_1838,N_1989);
nand U2616 (N_2616,N_1675,N_1546);
nand U2617 (N_2617,N_1718,N_2099);
and U2618 (N_2618,N_2183,N_1576);
nor U2619 (N_2619,N_2091,N_1836);
nor U2620 (N_2620,N_1964,N_1529);
or U2621 (N_2621,N_1624,N_2072);
nor U2622 (N_2622,N_1661,N_1955);
and U2623 (N_2623,N_2169,N_1918);
nand U2624 (N_2624,N_1681,N_1620);
nor U2625 (N_2625,N_2071,N_1850);
and U2626 (N_2626,N_1614,N_1766);
nand U2627 (N_2627,N_1562,N_2173);
and U2628 (N_2628,N_1616,N_2087);
nand U2629 (N_2629,N_1516,N_1584);
nor U2630 (N_2630,N_2135,N_1986);
or U2631 (N_2631,N_1639,N_1812);
or U2632 (N_2632,N_2165,N_1972);
and U2633 (N_2633,N_2140,N_1567);
and U2634 (N_2634,N_2110,N_1903);
nor U2635 (N_2635,N_1576,N_2139);
or U2636 (N_2636,N_1767,N_1574);
nor U2637 (N_2637,N_1878,N_1680);
or U2638 (N_2638,N_2249,N_1754);
nor U2639 (N_2639,N_2195,N_2043);
nor U2640 (N_2640,N_1579,N_1959);
or U2641 (N_2641,N_1506,N_1721);
or U2642 (N_2642,N_1767,N_2003);
or U2643 (N_2643,N_1557,N_2155);
or U2644 (N_2644,N_2247,N_2043);
and U2645 (N_2645,N_2122,N_2091);
nor U2646 (N_2646,N_2137,N_1953);
and U2647 (N_2647,N_1576,N_2115);
or U2648 (N_2648,N_1642,N_1911);
nor U2649 (N_2649,N_1788,N_1928);
nand U2650 (N_2650,N_2186,N_1563);
or U2651 (N_2651,N_1712,N_1652);
nor U2652 (N_2652,N_1751,N_1600);
or U2653 (N_2653,N_2241,N_1683);
nor U2654 (N_2654,N_1847,N_1795);
nand U2655 (N_2655,N_2191,N_1661);
nand U2656 (N_2656,N_1760,N_2139);
nand U2657 (N_2657,N_1862,N_1746);
and U2658 (N_2658,N_1736,N_1741);
nand U2659 (N_2659,N_1864,N_1957);
nor U2660 (N_2660,N_1757,N_2106);
nand U2661 (N_2661,N_2168,N_2217);
or U2662 (N_2662,N_2139,N_1735);
and U2663 (N_2663,N_1767,N_1813);
nor U2664 (N_2664,N_1911,N_1638);
or U2665 (N_2665,N_1579,N_1968);
and U2666 (N_2666,N_2020,N_1579);
nor U2667 (N_2667,N_2063,N_1568);
nand U2668 (N_2668,N_1944,N_1829);
nand U2669 (N_2669,N_2013,N_2004);
nand U2670 (N_2670,N_2208,N_1972);
and U2671 (N_2671,N_1579,N_1812);
nor U2672 (N_2672,N_1838,N_1589);
nor U2673 (N_2673,N_1978,N_1531);
nor U2674 (N_2674,N_1952,N_1641);
or U2675 (N_2675,N_2102,N_2231);
nor U2676 (N_2676,N_1517,N_1842);
and U2677 (N_2677,N_1535,N_1812);
and U2678 (N_2678,N_1595,N_1910);
nand U2679 (N_2679,N_2151,N_2198);
nand U2680 (N_2680,N_2228,N_1597);
nand U2681 (N_2681,N_2166,N_1810);
nor U2682 (N_2682,N_1997,N_1888);
or U2683 (N_2683,N_1853,N_1545);
or U2684 (N_2684,N_1877,N_2124);
nor U2685 (N_2685,N_1928,N_2218);
and U2686 (N_2686,N_2018,N_1928);
nor U2687 (N_2687,N_1943,N_1818);
nand U2688 (N_2688,N_1611,N_2195);
nand U2689 (N_2689,N_1558,N_1676);
nand U2690 (N_2690,N_1979,N_1778);
and U2691 (N_2691,N_2139,N_1975);
and U2692 (N_2692,N_1586,N_1971);
or U2693 (N_2693,N_1801,N_1945);
and U2694 (N_2694,N_1530,N_1776);
and U2695 (N_2695,N_2090,N_1583);
nand U2696 (N_2696,N_1852,N_1799);
nand U2697 (N_2697,N_2186,N_1900);
nand U2698 (N_2698,N_2053,N_2107);
and U2699 (N_2699,N_1510,N_1624);
and U2700 (N_2700,N_1901,N_2245);
nor U2701 (N_2701,N_1521,N_1694);
or U2702 (N_2702,N_1742,N_2077);
nor U2703 (N_2703,N_2100,N_1586);
nor U2704 (N_2704,N_1984,N_1780);
xnor U2705 (N_2705,N_1695,N_2178);
and U2706 (N_2706,N_1899,N_2001);
xor U2707 (N_2707,N_1869,N_1558);
or U2708 (N_2708,N_1984,N_2180);
and U2709 (N_2709,N_2216,N_2243);
or U2710 (N_2710,N_2001,N_1663);
or U2711 (N_2711,N_1784,N_1519);
nor U2712 (N_2712,N_1501,N_1944);
and U2713 (N_2713,N_1989,N_2097);
nor U2714 (N_2714,N_2203,N_1950);
or U2715 (N_2715,N_1518,N_1923);
nor U2716 (N_2716,N_2039,N_1538);
and U2717 (N_2717,N_1579,N_1619);
and U2718 (N_2718,N_2093,N_1974);
or U2719 (N_2719,N_2161,N_2065);
nand U2720 (N_2720,N_1662,N_2154);
nand U2721 (N_2721,N_1677,N_1780);
or U2722 (N_2722,N_1805,N_1842);
and U2723 (N_2723,N_1815,N_1542);
and U2724 (N_2724,N_1527,N_1993);
and U2725 (N_2725,N_1829,N_2122);
or U2726 (N_2726,N_1610,N_1701);
or U2727 (N_2727,N_1591,N_1639);
xor U2728 (N_2728,N_2119,N_1961);
or U2729 (N_2729,N_2121,N_2119);
nor U2730 (N_2730,N_1606,N_1983);
nor U2731 (N_2731,N_1502,N_1558);
and U2732 (N_2732,N_1676,N_1624);
and U2733 (N_2733,N_2124,N_1905);
and U2734 (N_2734,N_2105,N_1712);
or U2735 (N_2735,N_1693,N_1813);
and U2736 (N_2736,N_1620,N_2079);
or U2737 (N_2737,N_1780,N_2112);
nand U2738 (N_2738,N_1513,N_2052);
nor U2739 (N_2739,N_1837,N_2209);
nor U2740 (N_2740,N_1991,N_1887);
nand U2741 (N_2741,N_2111,N_1598);
and U2742 (N_2742,N_2005,N_2146);
nor U2743 (N_2743,N_1579,N_1814);
or U2744 (N_2744,N_2138,N_1607);
or U2745 (N_2745,N_1665,N_2164);
nand U2746 (N_2746,N_1563,N_2219);
nand U2747 (N_2747,N_2053,N_2088);
xnor U2748 (N_2748,N_1638,N_2245);
and U2749 (N_2749,N_1723,N_1728);
or U2750 (N_2750,N_2119,N_1655);
nor U2751 (N_2751,N_2188,N_2072);
and U2752 (N_2752,N_1824,N_1716);
and U2753 (N_2753,N_2015,N_2113);
or U2754 (N_2754,N_1952,N_1552);
nor U2755 (N_2755,N_1916,N_1774);
nand U2756 (N_2756,N_2158,N_1667);
nand U2757 (N_2757,N_1771,N_2112);
nand U2758 (N_2758,N_1641,N_1942);
nor U2759 (N_2759,N_1735,N_2101);
nand U2760 (N_2760,N_1556,N_2028);
or U2761 (N_2761,N_1901,N_2173);
nand U2762 (N_2762,N_1979,N_2052);
or U2763 (N_2763,N_2157,N_1787);
or U2764 (N_2764,N_2241,N_1890);
nand U2765 (N_2765,N_1702,N_1731);
nor U2766 (N_2766,N_1805,N_1861);
nor U2767 (N_2767,N_1859,N_1655);
nand U2768 (N_2768,N_1661,N_1755);
nand U2769 (N_2769,N_1536,N_1982);
or U2770 (N_2770,N_2156,N_2031);
nor U2771 (N_2771,N_1510,N_2056);
nand U2772 (N_2772,N_2087,N_1529);
nor U2773 (N_2773,N_1640,N_2197);
nor U2774 (N_2774,N_2109,N_2034);
or U2775 (N_2775,N_1760,N_1883);
nand U2776 (N_2776,N_2063,N_2142);
or U2777 (N_2777,N_1669,N_1954);
nor U2778 (N_2778,N_1664,N_1826);
nand U2779 (N_2779,N_1948,N_2008);
or U2780 (N_2780,N_2236,N_1644);
or U2781 (N_2781,N_1800,N_1868);
nor U2782 (N_2782,N_1785,N_2169);
or U2783 (N_2783,N_1905,N_1772);
and U2784 (N_2784,N_2206,N_1770);
nor U2785 (N_2785,N_2224,N_1520);
nand U2786 (N_2786,N_1960,N_1931);
nor U2787 (N_2787,N_2236,N_1938);
and U2788 (N_2788,N_1723,N_1664);
and U2789 (N_2789,N_1614,N_1589);
nand U2790 (N_2790,N_2181,N_1906);
or U2791 (N_2791,N_1972,N_1911);
nand U2792 (N_2792,N_1698,N_2188);
or U2793 (N_2793,N_2086,N_2189);
nor U2794 (N_2794,N_1524,N_2091);
nand U2795 (N_2795,N_1883,N_2066);
nand U2796 (N_2796,N_1703,N_1538);
nand U2797 (N_2797,N_1897,N_1883);
and U2798 (N_2798,N_2126,N_1559);
and U2799 (N_2799,N_1770,N_1538);
xnor U2800 (N_2800,N_1836,N_1649);
xnor U2801 (N_2801,N_1766,N_1845);
nand U2802 (N_2802,N_2151,N_1638);
nand U2803 (N_2803,N_1928,N_2054);
and U2804 (N_2804,N_2151,N_1935);
and U2805 (N_2805,N_1825,N_1662);
nand U2806 (N_2806,N_1881,N_2038);
and U2807 (N_2807,N_1822,N_1637);
or U2808 (N_2808,N_1842,N_2106);
xor U2809 (N_2809,N_1673,N_1735);
or U2810 (N_2810,N_2126,N_1744);
or U2811 (N_2811,N_1830,N_1797);
and U2812 (N_2812,N_1950,N_2042);
or U2813 (N_2813,N_1670,N_2110);
or U2814 (N_2814,N_1859,N_1999);
xor U2815 (N_2815,N_2039,N_2239);
nor U2816 (N_2816,N_1568,N_2105);
or U2817 (N_2817,N_2248,N_2163);
and U2818 (N_2818,N_2123,N_1627);
or U2819 (N_2819,N_1812,N_1713);
or U2820 (N_2820,N_2011,N_1712);
and U2821 (N_2821,N_1741,N_2031);
nand U2822 (N_2822,N_1530,N_1582);
and U2823 (N_2823,N_1924,N_1878);
nor U2824 (N_2824,N_2040,N_1993);
and U2825 (N_2825,N_2221,N_1624);
and U2826 (N_2826,N_1586,N_1534);
nand U2827 (N_2827,N_2154,N_1906);
nor U2828 (N_2828,N_1737,N_1663);
nand U2829 (N_2829,N_2015,N_1589);
or U2830 (N_2830,N_1947,N_1835);
or U2831 (N_2831,N_2038,N_1506);
or U2832 (N_2832,N_1682,N_1781);
xnor U2833 (N_2833,N_2229,N_1785);
and U2834 (N_2834,N_2167,N_2183);
or U2835 (N_2835,N_1758,N_2034);
nand U2836 (N_2836,N_1541,N_1696);
and U2837 (N_2837,N_2056,N_2176);
or U2838 (N_2838,N_2194,N_2051);
nand U2839 (N_2839,N_2181,N_2035);
and U2840 (N_2840,N_1829,N_1567);
nor U2841 (N_2841,N_2025,N_1735);
nand U2842 (N_2842,N_1947,N_1526);
and U2843 (N_2843,N_1834,N_1695);
nand U2844 (N_2844,N_1963,N_1703);
nor U2845 (N_2845,N_2149,N_1803);
or U2846 (N_2846,N_1528,N_2145);
and U2847 (N_2847,N_2194,N_1931);
nand U2848 (N_2848,N_1540,N_2017);
nor U2849 (N_2849,N_2066,N_1840);
or U2850 (N_2850,N_2173,N_2162);
nand U2851 (N_2851,N_2150,N_2005);
nor U2852 (N_2852,N_1617,N_1531);
nor U2853 (N_2853,N_1916,N_1557);
and U2854 (N_2854,N_1558,N_2041);
nand U2855 (N_2855,N_1595,N_1841);
nor U2856 (N_2856,N_2238,N_1994);
and U2857 (N_2857,N_2001,N_1543);
or U2858 (N_2858,N_2117,N_2095);
or U2859 (N_2859,N_1748,N_2060);
nand U2860 (N_2860,N_2210,N_1929);
or U2861 (N_2861,N_2225,N_2151);
or U2862 (N_2862,N_2148,N_1896);
nand U2863 (N_2863,N_2092,N_2201);
nand U2864 (N_2864,N_1949,N_1646);
or U2865 (N_2865,N_1860,N_1661);
and U2866 (N_2866,N_1986,N_2120);
nor U2867 (N_2867,N_1571,N_1517);
nand U2868 (N_2868,N_1720,N_2043);
nand U2869 (N_2869,N_1757,N_2009);
and U2870 (N_2870,N_2175,N_2177);
or U2871 (N_2871,N_2094,N_1952);
nor U2872 (N_2872,N_1615,N_1543);
or U2873 (N_2873,N_2154,N_2103);
nor U2874 (N_2874,N_2203,N_1668);
or U2875 (N_2875,N_1518,N_1501);
nor U2876 (N_2876,N_1804,N_2168);
or U2877 (N_2877,N_1818,N_1698);
or U2878 (N_2878,N_2085,N_2102);
or U2879 (N_2879,N_1553,N_1878);
nor U2880 (N_2880,N_2166,N_2196);
and U2881 (N_2881,N_1799,N_1914);
or U2882 (N_2882,N_1548,N_1664);
and U2883 (N_2883,N_2176,N_1760);
and U2884 (N_2884,N_1990,N_2044);
or U2885 (N_2885,N_1856,N_2159);
nand U2886 (N_2886,N_1847,N_2043);
and U2887 (N_2887,N_1649,N_1603);
nor U2888 (N_2888,N_2039,N_1527);
nor U2889 (N_2889,N_1564,N_1524);
nor U2890 (N_2890,N_2026,N_1937);
or U2891 (N_2891,N_1986,N_2044);
nor U2892 (N_2892,N_2001,N_1813);
or U2893 (N_2893,N_1874,N_1771);
nand U2894 (N_2894,N_1671,N_1645);
nor U2895 (N_2895,N_1871,N_1511);
and U2896 (N_2896,N_1556,N_2048);
or U2897 (N_2897,N_1575,N_1943);
or U2898 (N_2898,N_1870,N_1688);
and U2899 (N_2899,N_1620,N_2144);
and U2900 (N_2900,N_2198,N_1767);
and U2901 (N_2901,N_1696,N_2172);
and U2902 (N_2902,N_1888,N_1752);
or U2903 (N_2903,N_2036,N_2069);
and U2904 (N_2904,N_2155,N_2169);
nand U2905 (N_2905,N_1623,N_1770);
or U2906 (N_2906,N_1680,N_2207);
or U2907 (N_2907,N_1609,N_1743);
and U2908 (N_2908,N_1979,N_1924);
nor U2909 (N_2909,N_1815,N_1651);
or U2910 (N_2910,N_2246,N_2124);
xnor U2911 (N_2911,N_1740,N_1511);
and U2912 (N_2912,N_2200,N_1672);
nand U2913 (N_2913,N_1595,N_2106);
nand U2914 (N_2914,N_1711,N_1974);
nand U2915 (N_2915,N_1897,N_1500);
and U2916 (N_2916,N_1643,N_1669);
and U2917 (N_2917,N_2160,N_2156);
nand U2918 (N_2918,N_1997,N_1656);
nand U2919 (N_2919,N_1604,N_2038);
and U2920 (N_2920,N_2225,N_2196);
nand U2921 (N_2921,N_1839,N_1925);
nor U2922 (N_2922,N_2058,N_2162);
nand U2923 (N_2923,N_1953,N_2211);
or U2924 (N_2924,N_2086,N_1623);
or U2925 (N_2925,N_1524,N_1874);
or U2926 (N_2926,N_2078,N_1723);
nor U2927 (N_2927,N_2060,N_1971);
nor U2928 (N_2928,N_1661,N_1866);
nand U2929 (N_2929,N_1734,N_1561);
nand U2930 (N_2930,N_1722,N_1810);
nand U2931 (N_2931,N_2213,N_1534);
and U2932 (N_2932,N_2187,N_1773);
and U2933 (N_2933,N_1775,N_1997);
nor U2934 (N_2934,N_1655,N_1718);
nand U2935 (N_2935,N_1525,N_1937);
xor U2936 (N_2936,N_1964,N_1582);
nor U2937 (N_2937,N_1883,N_1797);
nand U2938 (N_2938,N_1817,N_1607);
and U2939 (N_2939,N_1917,N_1571);
or U2940 (N_2940,N_1523,N_2075);
nor U2941 (N_2941,N_2003,N_1705);
and U2942 (N_2942,N_2085,N_2143);
nor U2943 (N_2943,N_1839,N_1714);
or U2944 (N_2944,N_1870,N_1756);
nand U2945 (N_2945,N_1968,N_1790);
or U2946 (N_2946,N_1683,N_2094);
and U2947 (N_2947,N_1630,N_1658);
nand U2948 (N_2948,N_2140,N_1623);
and U2949 (N_2949,N_1650,N_1987);
nor U2950 (N_2950,N_1576,N_2007);
nand U2951 (N_2951,N_1983,N_1570);
or U2952 (N_2952,N_1887,N_1734);
nand U2953 (N_2953,N_1724,N_1854);
or U2954 (N_2954,N_2187,N_2244);
or U2955 (N_2955,N_1573,N_1850);
nor U2956 (N_2956,N_1808,N_1900);
nand U2957 (N_2957,N_2078,N_1556);
nor U2958 (N_2958,N_1971,N_2174);
nor U2959 (N_2959,N_2130,N_1654);
nand U2960 (N_2960,N_1587,N_2034);
nor U2961 (N_2961,N_2133,N_1924);
nor U2962 (N_2962,N_1895,N_1753);
and U2963 (N_2963,N_1770,N_2208);
nand U2964 (N_2964,N_1777,N_2238);
and U2965 (N_2965,N_1760,N_1514);
and U2966 (N_2966,N_2198,N_2221);
nor U2967 (N_2967,N_1844,N_1700);
and U2968 (N_2968,N_2026,N_1561);
nand U2969 (N_2969,N_2120,N_2145);
nor U2970 (N_2970,N_1771,N_2128);
and U2971 (N_2971,N_1586,N_1723);
nor U2972 (N_2972,N_2187,N_2221);
nand U2973 (N_2973,N_1886,N_1703);
xnor U2974 (N_2974,N_2148,N_1807);
or U2975 (N_2975,N_1699,N_2131);
or U2976 (N_2976,N_1805,N_1605);
and U2977 (N_2977,N_1558,N_1525);
or U2978 (N_2978,N_2000,N_1980);
or U2979 (N_2979,N_1697,N_2074);
nor U2980 (N_2980,N_1715,N_2176);
nand U2981 (N_2981,N_2236,N_1865);
and U2982 (N_2982,N_1707,N_2093);
nand U2983 (N_2983,N_2089,N_1509);
or U2984 (N_2984,N_1924,N_2197);
xnor U2985 (N_2985,N_1599,N_1592);
or U2986 (N_2986,N_1809,N_2147);
nor U2987 (N_2987,N_1769,N_2248);
or U2988 (N_2988,N_1861,N_2190);
nand U2989 (N_2989,N_1752,N_1521);
nand U2990 (N_2990,N_2003,N_1617);
nand U2991 (N_2991,N_2243,N_1734);
nand U2992 (N_2992,N_2111,N_2020);
or U2993 (N_2993,N_2158,N_1922);
or U2994 (N_2994,N_1749,N_1689);
or U2995 (N_2995,N_1634,N_1500);
or U2996 (N_2996,N_1827,N_1713);
or U2997 (N_2997,N_1882,N_1793);
or U2998 (N_2998,N_2001,N_2156);
nor U2999 (N_2999,N_2063,N_2141);
and UO_0 (O_0,N_2405,N_2493);
nor UO_1 (O_1,N_2372,N_2956);
and UO_2 (O_2,N_2615,N_2285);
nand UO_3 (O_3,N_2789,N_2921);
nor UO_4 (O_4,N_2588,N_2552);
nand UO_5 (O_5,N_2254,N_2577);
nand UO_6 (O_6,N_2265,N_2337);
and UO_7 (O_7,N_2797,N_2748);
or UO_8 (O_8,N_2884,N_2987);
or UO_9 (O_9,N_2466,N_2482);
nand UO_10 (O_10,N_2486,N_2593);
nor UO_11 (O_11,N_2270,N_2346);
nand UO_12 (O_12,N_2375,N_2643);
and UO_13 (O_13,N_2299,N_2656);
and UO_14 (O_14,N_2424,N_2566);
and UO_15 (O_15,N_2312,N_2431);
or UO_16 (O_16,N_2929,N_2521);
or UO_17 (O_17,N_2835,N_2351);
or UO_18 (O_18,N_2589,N_2983);
or UO_19 (O_19,N_2638,N_2878);
nand UO_20 (O_20,N_2870,N_2449);
and UO_21 (O_21,N_2894,N_2652);
or UO_22 (O_22,N_2840,N_2551);
nand UO_23 (O_23,N_2947,N_2649);
nand UO_24 (O_24,N_2707,N_2496);
and UO_25 (O_25,N_2562,N_2487);
and UO_26 (O_26,N_2497,N_2730);
nor UO_27 (O_27,N_2595,N_2683);
nor UO_28 (O_28,N_2934,N_2988);
nor UO_29 (O_29,N_2474,N_2542);
and UO_30 (O_30,N_2286,N_2480);
xor UO_31 (O_31,N_2525,N_2903);
nor UO_32 (O_32,N_2569,N_2338);
nor UO_33 (O_33,N_2289,N_2268);
nand UO_34 (O_34,N_2256,N_2791);
and UO_35 (O_35,N_2607,N_2612);
or UO_36 (O_36,N_2689,N_2845);
nor UO_37 (O_37,N_2253,N_2839);
or UO_38 (O_38,N_2933,N_2874);
nand UO_39 (O_39,N_2796,N_2288);
xnor UO_40 (O_40,N_2995,N_2526);
nand UO_41 (O_41,N_2782,N_2483);
nand UO_42 (O_42,N_2655,N_2781);
and UO_43 (O_43,N_2668,N_2650);
nor UO_44 (O_44,N_2583,N_2883);
nor UO_45 (O_45,N_2777,N_2920);
and UO_46 (O_46,N_2358,N_2645);
or UO_47 (O_47,N_2898,N_2659);
or UO_48 (O_48,N_2842,N_2618);
nand UO_49 (O_49,N_2634,N_2460);
or UO_50 (O_50,N_2602,N_2553);
and UO_51 (O_51,N_2477,N_2769);
and UO_52 (O_52,N_2413,N_2274);
nor UO_53 (O_53,N_2913,N_2524);
and UO_54 (O_54,N_2365,N_2805);
nor UO_55 (O_55,N_2567,N_2317);
or UO_56 (O_56,N_2957,N_2331);
and UO_57 (O_57,N_2505,N_2808);
and UO_58 (O_58,N_2742,N_2681);
nor UO_59 (O_59,N_2627,N_2812);
nor UO_60 (O_60,N_2339,N_2290);
or UO_61 (O_61,N_2579,N_2963);
nand UO_62 (O_62,N_2775,N_2440);
nor UO_63 (O_63,N_2648,N_2904);
nor UO_64 (O_64,N_2386,N_2815);
and UO_65 (O_65,N_2370,N_2547);
and UO_66 (O_66,N_2905,N_2900);
nor UO_67 (O_67,N_2379,N_2434);
nor UO_68 (O_68,N_2374,N_2837);
xnor UO_69 (O_69,N_2733,N_2258);
and UO_70 (O_70,N_2565,N_2600);
nand UO_71 (O_71,N_2294,N_2457);
or UO_72 (O_72,N_2251,N_2546);
nor UO_73 (O_73,N_2908,N_2488);
or UO_74 (O_74,N_2669,N_2470);
or UO_75 (O_75,N_2529,N_2662);
nor UO_76 (O_76,N_2794,N_2978);
or UO_77 (O_77,N_2427,N_2303);
nand UO_78 (O_78,N_2522,N_2676);
or UO_79 (O_79,N_2262,N_2320);
nor UO_80 (O_80,N_2397,N_2484);
nand UO_81 (O_81,N_2369,N_2793);
and UO_82 (O_82,N_2550,N_2385);
or UO_83 (O_83,N_2611,N_2384);
nor UO_84 (O_84,N_2932,N_2519);
and UO_85 (O_85,N_2902,N_2768);
nand UO_86 (O_86,N_2887,N_2863);
and UO_87 (O_87,N_2364,N_2786);
and UO_88 (O_88,N_2964,N_2972);
and UO_89 (O_89,N_2624,N_2401);
or UO_90 (O_90,N_2330,N_2347);
nor UO_91 (O_91,N_2927,N_2468);
and UO_92 (O_92,N_2727,N_2500);
and UO_93 (O_93,N_2412,N_2642);
or UO_94 (O_94,N_2272,N_2387);
nor UO_95 (O_95,N_2784,N_2680);
nor UO_96 (O_96,N_2471,N_2378);
nor UO_97 (O_97,N_2628,N_2545);
nor UO_98 (O_98,N_2451,N_2930);
nand UO_99 (O_99,N_2419,N_2335);
nor UO_100 (O_100,N_2925,N_2275);
nand UO_101 (O_101,N_2381,N_2937);
nor UO_102 (O_102,N_2296,N_2968);
nor UO_103 (O_103,N_2392,N_2435);
and UO_104 (O_104,N_2907,N_2635);
and UO_105 (O_105,N_2584,N_2914);
or UO_106 (O_106,N_2721,N_2459);
nand UO_107 (O_107,N_2561,N_2574);
nand UO_108 (O_108,N_2509,N_2536);
xnor UO_109 (O_109,N_2432,N_2657);
and UO_110 (O_110,N_2663,N_2818);
or UO_111 (O_111,N_2672,N_2445);
nor UO_112 (O_112,N_2757,N_2700);
nand UO_113 (O_113,N_2362,N_2311);
nand UO_114 (O_114,N_2520,N_2325);
nor UO_115 (O_115,N_2350,N_2341);
and UO_116 (O_116,N_2984,N_2792);
or UO_117 (O_117,N_2531,N_2877);
and UO_118 (O_118,N_2605,N_2323);
or UO_119 (O_119,N_2620,N_2368);
nand UO_120 (O_120,N_2758,N_2410);
and UO_121 (O_121,N_2264,N_2834);
nor UO_122 (O_122,N_2388,N_2910);
nor UO_123 (O_123,N_2633,N_2918);
and UO_124 (O_124,N_2982,N_2617);
nor UO_125 (O_125,N_2585,N_2454);
xnor UO_126 (O_126,N_2951,N_2478);
or UO_127 (O_127,N_2587,N_2590);
or UO_128 (O_128,N_2363,N_2436);
nand UO_129 (O_129,N_2508,N_2755);
nor UO_130 (O_130,N_2785,N_2608);
nand UO_131 (O_131,N_2847,N_2686);
or UO_132 (O_132,N_2527,N_2799);
and UO_133 (O_133,N_2996,N_2879);
or UO_134 (O_134,N_2489,N_2557);
nor UO_135 (O_135,N_2804,N_2670);
and UO_136 (O_136,N_2621,N_2261);
nor UO_137 (O_137,N_2813,N_2543);
and UO_138 (O_138,N_2352,N_2534);
or UO_139 (O_139,N_2967,N_2698);
and UO_140 (O_140,N_2301,N_2899);
and UO_141 (O_141,N_2773,N_2776);
nand UO_142 (O_142,N_2414,N_2267);
nor UO_143 (O_143,N_2532,N_2257);
and UO_144 (O_144,N_2896,N_2462);
nand UO_145 (O_145,N_2959,N_2958);
and UO_146 (O_146,N_2671,N_2919);
and UO_147 (O_147,N_2622,N_2269);
and UO_148 (O_148,N_2667,N_2753);
and UO_149 (O_149,N_2640,N_2823);
nor UO_150 (O_150,N_2740,N_2438);
nor UO_151 (O_151,N_2283,N_2833);
and UO_152 (O_152,N_2568,N_2549);
and UO_153 (O_153,N_2336,N_2518);
xnor UO_154 (O_154,N_2399,N_2407);
nor UO_155 (O_155,N_2409,N_2450);
nor UO_156 (O_156,N_2690,N_2810);
nor UO_157 (O_157,N_2788,N_2997);
or UO_158 (O_158,N_2644,N_2357);
or UO_159 (O_159,N_2580,N_2880);
and UO_160 (O_160,N_2291,N_2430);
and UO_161 (O_161,N_2806,N_2637);
nor UO_162 (O_162,N_2315,N_2609);
nand UO_163 (O_163,N_2917,N_2660);
and UO_164 (O_164,N_2770,N_2586);
and UO_165 (O_165,N_2429,N_2390);
nor UO_166 (O_166,N_2575,N_2827);
and UO_167 (O_167,N_2674,N_2772);
nand UO_168 (O_168,N_2979,N_2598);
nor UO_169 (O_169,N_2393,N_2928);
nor UO_170 (O_170,N_2467,N_2974);
or UO_171 (O_171,N_2687,N_2795);
or UO_172 (O_172,N_2949,N_2857);
nand UO_173 (O_173,N_2380,N_2761);
or UO_174 (O_174,N_2666,N_2528);
nor UO_175 (O_175,N_2359,N_2860);
nand UO_176 (O_176,N_2825,N_2821);
and UO_177 (O_177,N_2464,N_2475);
and UO_178 (O_178,N_2647,N_2779);
nor UO_179 (O_179,N_2415,N_2625);
and UO_180 (O_180,N_2843,N_2911);
and UO_181 (O_181,N_2737,N_2537);
nor UO_182 (O_182,N_2292,N_2564);
and UO_183 (O_183,N_2836,N_2992);
or UO_184 (O_184,N_2811,N_2456);
or UO_185 (O_185,N_2846,N_2377);
nor UO_186 (O_186,N_2719,N_2861);
or UO_187 (O_187,N_2893,N_2945);
nor UO_188 (O_188,N_2807,N_2309);
nor UO_189 (O_189,N_2306,N_2280);
nor UO_190 (O_190,N_2916,N_2771);
and UO_191 (O_191,N_2616,N_2329);
or UO_192 (O_192,N_2559,N_2334);
or UO_193 (O_193,N_2631,N_2876);
nor UO_194 (O_194,N_2849,N_2867);
and UO_195 (O_195,N_2851,N_2485);
nand UO_196 (O_196,N_2856,N_2639);
nand UO_197 (O_197,N_2349,N_2504);
nand UO_198 (O_198,N_2926,N_2855);
nand UO_199 (O_199,N_2872,N_2400);
xnor UO_200 (O_200,N_2408,N_2512);
nor UO_201 (O_201,N_2455,N_2971);
nor UO_202 (O_202,N_2591,N_2989);
nor UO_203 (O_203,N_2703,N_2844);
nor UO_204 (O_204,N_2554,N_2780);
and UO_205 (O_205,N_2540,N_2367);
nor UO_206 (O_206,N_2322,N_2739);
or UO_207 (O_207,N_2922,N_2441);
and UO_208 (O_208,N_2476,N_2382);
nand UO_209 (O_209,N_2985,N_2886);
or UO_210 (O_210,N_2327,N_2859);
xnor UO_211 (O_211,N_2962,N_2479);
xnor UO_212 (O_212,N_2749,N_2724);
nand UO_213 (O_213,N_2308,N_2720);
and UO_214 (O_214,N_2935,N_2340);
or UO_215 (O_215,N_2344,N_2688);
and UO_216 (O_216,N_2754,N_2305);
or UO_217 (O_217,N_2538,N_2428);
or UO_218 (O_218,N_2866,N_2875);
xor UO_219 (O_219,N_2658,N_2389);
nand UO_220 (O_220,N_2417,N_2723);
and UO_221 (O_221,N_2970,N_2915);
nand UO_222 (O_222,N_2864,N_2743);
nor UO_223 (O_223,N_2396,N_2882);
nor UO_224 (O_224,N_2831,N_2885);
nor UO_225 (O_225,N_2912,N_2324);
nor UO_226 (O_226,N_2333,N_2582);
or UO_227 (O_227,N_2715,N_2848);
nand UO_228 (O_228,N_2318,N_2741);
nand UO_229 (O_229,N_2502,N_2778);
nor UO_230 (O_230,N_2544,N_2800);
and UO_231 (O_231,N_2398,N_2422);
nand UO_232 (O_232,N_2871,N_2986);
nor UO_233 (O_233,N_2641,N_2766);
or UO_234 (O_234,N_2418,N_2490);
nor UO_235 (O_235,N_2439,N_2714);
nor UO_236 (O_236,N_2708,N_2960);
nand UO_237 (O_237,N_2767,N_2701);
xnor UO_238 (O_238,N_2302,N_2682);
or UO_239 (O_239,N_2383,N_2250);
nand UO_240 (O_240,N_2498,N_2371);
or UO_241 (O_241,N_2973,N_2924);
nand UO_242 (O_242,N_2646,N_2798);
nand UO_243 (O_243,N_2709,N_2993);
nor UO_244 (O_244,N_2950,N_2759);
or UO_245 (O_245,N_2745,N_2853);
nand UO_246 (O_246,N_2822,N_2437);
or UO_247 (O_247,N_2613,N_2953);
nand UO_248 (O_248,N_2726,N_2817);
nand UO_249 (O_249,N_2510,N_2906);
and UO_250 (O_250,N_2404,N_2492);
nand UO_251 (O_251,N_2969,N_2623);
or UO_252 (O_252,N_2814,N_2300);
xnor UO_253 (O_253,N_2548,N_2517);
or UO_254 (O_254,N_2573,N_2391);
nand UO_255 (O_255,N_2354,N_2936);
nor UO_256 (O_256,N_2763,N_2691);
or UO_257 (O_257,N_2696,N_2751);
nor UO_258 (O_258,N_2541,N_2684);
nor UO_259 (O_259,N_2980,N_2416);
nor UO_260 (O_260,N_2361,N_2923);
and UO_261 (O_261,N_2728,N_2994);
xnor UO_262 (O_262,N_2854,N_2348);
nor UO_263 (O_263,N_2446,N_2629);
nand UO_264 (O_264,N_2735,N_2803);
and UO_265 (O_265,N_2494,N_2802);
and UO_266 (O_266,N_2736,N_2705);
xnor UO_267 (O_267,N_2816,N_2991);
or UO_268 (O_268,N_2604,N_2411);
or UO_269 (O_269,N_2717,N_2673);
nor UO_270 (O_270,N_2287,N_2444);
and UO_271 (O_271,N_2343,N_2353);
or UO_272 (O_272,N_2626,N_2284);
and UO_273 (O_273,N_2661,N_2693);
nand UO_274 (O_274,N_2865,N_2838);
nor UO_275 (O_275,N_2603,N_2718);
or UO_276 (O_276,N_2495,N_2328);
nor UO_277 (O_277,N_2281,N_2423);
or UO_278 (O_278,N_2694,N_2961);
nor UO_279 (O_279,N_2571,N_2998);
nand UO_280 (O_280,N_2578,N_2402);
and UO_281 (O_281,N_2809,N_2515);
nand UO_282 (O_282,N_2293,N_2895);
nand UO_283 (O_283,N_2679,N_2889);
xnor UO_284 (O_284,N_2255,N_2345);
or UO_285 (O_285,N_2897,N_2712);
nor UO_286 (O_286,N_2403,N_2862);
or UO_287 (O_287,N_2976,N_2463);
nor UO_288 (O_288,N_2734,N_2732);
or UO_289 (O_289,N_2319,N_2630);
nor UO_290 (O_290,N_2533,N_2356);
xnor UO_291 (O_291,N_2263,N_2828);
nand UO_292 (O_292,N_2832,N_2752);
or UO_293 (O_293,N_2266,N_2881);
nor UO_294 (O_294,N_2276,N_2954);
nand UO_295 (O_295,N_2426,N_2252);
nand UO_296 (O_296,N_2738,N_2975);
nor UO_297 (O_297,N_2503,N_2981);
and UO_298 (O_298,N_2523,N_2764);
nor UO_299 (O_299,N_2499,N_2888);
nor UO_300 (O_300,N_2819,N_2943);
and UO_301 (O_301,N_2314,N_2511);
nor UO_302 (O_302,N_2558,N_2572);
xor UO_303 (O_303,N_2297,N_2820);
nor UO_304 (O_304,N_2941,N_2260);
or UO_305 (O_305,N_2539,N_2373);
or UO_306 (O_306,N_2692,N_2614);
nand UO_307 (O_307,N_2420,N_2830);
and UO_308 (O_308,N_2452,N_2952);
nor UO_309 (O_309,N_2729,N_2581);
nor UO_310 (O_310,N_2801,N_2762);
nand UO_311 (O_311,N_2722,N_2790);
xor UO_312 (O_312,N_2619,N_2942);
nand UO_313 (O_313,N_2355,N_2279);
and UO_314 (O_314,N_2841,N_2295);
and UO_315 (O_315,N_2599,N_2891);
or UO_316 (O_316,N_2664,N_2946);
and UO_317 (O_317,N_2697,N_2756);
or UO_318 (O_318,N_2892,N_2597);
and UO_319 (O_319,N_2774,N_2535);
nor UO_320 (O_320,N_2596,N_2706);
nand UO_321 (O_321,N_2321,N_2725);
and UO_322 (O_322,N_2901,N_2273);
or UO_323 (O_323,N_2869,N_2278);
or UO_324 (O_324,N_2472,N_2282);
nor UO_325 (O_325,N_2744,N_2442);
and UO_326 (O_326,N_2516,N_2665);
or UO_327 (O_327,N_2277,N_2826);
nor UO_328 (O_328,N_2699,N_2829);
nand UO_329 (O_329,N_2506,N_2453);
nor UO_330 (O_330,N_2395,N_2491);
or UO_331 (O_331,N_2873,N_2465);
and UO_332 (O_332,N_2342,N_2563);
and UO_333 (O_333,N_2704,N_2458);
nand UO_334 (O_334,N_2360,N_2965);
nand UO_335 (O_335,N_2858,N_2990);
nor UO_336 (O_336,N_2850,N_2473);
and UO_337 (O_337,N_2461,N_2447);
nor UO_338 (O_338,N_2695,N_2713);
nor UO_339 (O_339,N_2570,N_2601);
xnor UO_340 (O_340,N_2594,N_2555);
and UO_341 (O_341,N_2868,N_2999);
nand UO_342 (O_342,N_2654,N_2443);
and UO_343 (O_343,N_2955,N_2421);
or UO_344 (O_344,N_2747,N_2939);
nor UO_345 (O_345,N_2501,N_2530);
and UO_346 (O_346,N_2406,N_2944);
nand UO_347 (O_347,N_2576,N_2787);
or UO_348 (O_348,N_2448,N_2710);
nand UO_349 (O_349,N_2514,N_2271);
or UO_350 (O_350,N_2556,N_2746);
and UO_351 (O_351,N_2481,N_2702);
nand UO_352 (O_352,N_2469,N_2966);
xor UO_353 (O_353,N_2948,N_2313);
nand UO_354 (O_354,N_2716,N_2677);
nor UO_355 (O_355,N_2310,N_2783);
nand UO_356 (O_356,N_2307,N_2394);
nor UO_357 (O_357,N_2376,N_2366);
and UO_358 (O_358,N_2750,N_2592);
nor UO_359 (O_359,N_2606,N_2675);
or UO_360 (O_360,N_2940,N_2636);
and UO_361 (O_361,N_2610,N_2433);
and UO_362 (O_362,N_2560,N_2938);
and UO_363 (O_363,N_2765,N_2977);
nand UO_364 (O_364,N_2685,N_2632);
nand UO_365 (O_365,N_2259,N_2304);
nand UO_366 (O_366,N_2711,N_2909);
and UO_367 (O_367,N_2651,N_2513);
nand UO_368 (O_368,N_2678,N_2731);
xnor UO_369 (O_369,N_2931,N_2425);
or UO_370 (O_370,N_2824,N_2852);
nand UO_371 (O_371,N_2298,N_2316);
nor UO_372 (O_372,N_2760,N_2653);
or UO_373 (O_373,N_2332,N_2326);
nand UO_374 (O_374,N_2890,N_2507);
nor UO_375 (O_375,N_2291,N_2774);
nand UO_376 (O_376,N_2413,N_2630);
nand UO_377 (O_377,N_2433,N_2775);
or UO_378 (O_378,N_2396,N_2418);
nand UO_379 (O_379,N_2655,N_2362);
or UO_380 (O_380,N_2429,N_2898);
nor UO_381 (O_381,N_2589,N_2624);
xnor UO_382 (O_382,N_2445,N_2737);
or UO_383 (O_383,N_2876,N_2727);
nand UO_384 (O_384,N_2790,N_2804);
nand UO_385 (O_385,N_2417,N_2534);
or UO_386 (O_386,N_2865,N_2840);
nor UO_387 (O_387,N_2928,N_2957);
nand UO_388 (O_388,N_2619,N_2789);
nand UO_389 (O_389,N_2615,N_2512);
nor UO_390 (O_390,N_2924,N_2387);
and UO_391 (O_391,N_2630,N_2683);
nand UO_392 (O_392,N_2513,N_2278);
and UO_393 (O_393,N_2302,N_2550);
nor UO_394 (O_394,N_2547,N_2925);
nor UO_395 (O_395,N_2861,N_2603);
and UO_396 (O_396,N_2897,N_2902);
nand UO_397 (O_397,N_2626,N_2681);
or UO_398 (O_398,N_2769,N_2299);
and UO_399 (O_399,N_2328,N_2468);
or UO_400 (O_400,N_2890,N_2292);
and UO_401 (O_401,N_2922,N_2583);
nor UO_402 (O_402,N_2406,N_2443);
nor UO_403 (O_403,N_2638,N_2812);
or UO_404 (O_404,N_2749,N_2346);
or UO_405 (O_405,N_2701,N_2888);
and UO_406 (O_406,N_2389,N_2320);
or UO_407 (O_407,N_2791,N_2711);
nor UO_408 (O_408,N_2812,N_2930);
nand UO_409 (O_409,N_2254,N_2903);
and UO_410 (O_410,N_2571,N_2801);
or UO_411 (O_411,N_2375,N_2696);
or UO_412 (O_412,N_2787,N_2606);
nand UO_413 (O_413,N_2927,N_2274);
or UO_414 (O_414,N_2983,N_2470);
nor UO_415 (O_415,N_2349,N_2957);
and UO_416 (O_416,N_2398,N_2763);
and UO_417 (O_417,N_2530,N_2993);
or UO_418 (O_418,N_2960,N_2771);
nor UO_419 (O_419,N_2874,N_2605);
nand UO_420 (O_420,N_2276,N_2576);
nor UO_421 (O_421,N_2564,N_2313);
nor UO_422 (O_422,N_2263,N_2583);
and UO_423 (O_423,N_2489,N_2403);
nand UO_424 (O_424,N_2366,N_2701);
nand UO_425 (O_425,N_2948,N_2483);
nor UO_426 (O_426,N_2618,N_2443);
and UO_427 (O_427,N_2992,N_2620);
and UO_428 (O_428,N_2399,N_2472);
nand UO_429 (O_429,N_2681,N_2717);
or UO_430 (O_430,N_2579,N_2802);
nor UO_431 (O_431,N_2576,N_2867);
or UO_432 (O_432,N_2348,N_2658);
nor UO_433 (O_433,N_2799,N_2939);
nor UO_434 (O_434,N_2897,N_2888);
nor UO_435 (O_435,N_2896,N_2507);
and UO_436 (O_436,N_2971,N_2511);
and UO_437 (O_437,N_2999,N_2836);
nand UO_438 (O_438,N_2985,N_2714);
nor UO_439 (O_439,N_2396,N_2853);
nor UO_440 (O_440,N_2291,N_2370);
nor UO_441 (O_441,N_2741,N_2722);
nand UO_442 (O_442,N_2398,N_2278);
nand UO_443 (O_443,N_2364,N_2796);
and UO_444 (O_444,N_2347,N_2931);
and UO_445 (O_445,N_2319,N_2920);
nor UO_446 (O_446,N_2552,N_2482);
nor UO_447 (O_447,N_2984,N_2318);
or UO_448 (O_448,N_2932,N_2455);
xor UO_449 (O_449,N_2830,N_2736);
or UO_450 (O_450,N_2852,N_2417);
nand UO_451 (O_451,N_2402,N_2422);
and UO_452 (O_452,N_2591,N_2861);
nand UO_453 (O_453,N_2643,N_2371);
and UO_454 (O_454,N_2574,N_2384);
nand UO_455 (O_455,N_2794,N_2624);
and UO_456 (O_456,N_2736,N_2323);
nand UO_457 (O_457,N_2306,N_2676);
and UO_458 (O_458,N_2730,N_2802);
nand UO_459 (O_459,N_2759,N_2427);
nand UO_460 (O_460,N_2647,N_2942);
or UO_461 (O_461,N_2941,N_2904);
nand UO_462 (O_462,N_2685,N_2711);
nand UO_463 (O_463,N_2665,N_2715);
and UO_464 (O_464,N_2900,N_2352);
or UO_465 (O_465,N_2252,N_2735);
nor UO_466 (O_466,N_2662,N_2697);
nor UO_467 (O_467,N_2255,N_2738);
nor UO_468 (O_468,N_2940,N_2935);
nand UO_469 (O_469,N_2643,N_2420);
nand UO_470 (O_470,N_2656,N_2488);
xor UO_471 (O_471,N_2543,N_2957);
nor UO_472 (O_472,N_2279,N_2650);
nand UO_473 (O_473,N_2504,N_2539);
and UO_474 (O_474,N_2514,N_2598);
nand UO_475 (O_475,N_2505,N_2644);
or UO_476 (O_476,N_2692,N_2635);
nor UO_477 (O_477,N_2662,N_2915);
and UO_478 (O_478,N_2355,N_2913);
or UO_479 (O_479,N_2424,N_2471);
and UO_480 (O_480,N_2965,N_2466);
and UO_481 (O_481,N_2792,N_2325);
nor UO_482 (O_482,N_2555,N_2394);
or UO_483 (O_483,N_2402,N_2834);
nor UO_484 (O_484,N_2379,N_2600);
xnor UO_485 (O_485,N_2628,N_2313);
and UO_486 (O_486,N_2426,N_2987);
nand UO_487 (O_487,N_2304,N_2512);
and UO_488 (O_488,N_2339,N_2647);
nor UO_489 (O_489,N_2590,N_2847);
and UO_490 (O_490,N_2869,N_2864);
and UO_491 (O_491,N_2998,N_2635);
nor UO_492 (O_492,N_2700,N_2413);
or UO_493 (O_493,N_2803,N_2967);
nand UO_494 (O_494,N_2329,N_2448);
and UO_495 (O_495,N_2618,N_2885);
or UO_496 (O_496,N_2725,N_2483);
nor UO_497 (O_497,N_2744,N_2921);
and UO_498 (O_498,N_2909,N_2877);
nor UO_499 (O_499,N_2544,N_2584);
endmodule