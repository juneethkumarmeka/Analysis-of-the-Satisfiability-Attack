module basic_750_5000_1000_25_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_576,In_3);
and U1 (N_1,In_716,In_316);
nor U2 (N_2,In_382,In_232);
nor U3 (N_3,In_643,In_214);
nand U4 (N_4,In_538,In_283);
or U5 (N_5,In_34,In_439);
or U6 (N_6,In_460,In_174);
or U7 (N_7,In_677,In_471);
or U8 (N_8,In_70,In_104);
or U9 (N_9,In_199,In_203);
or U10 (N_10,In_710,In_707);
or U11 (N_11,In_17,In_600);
or U12 (N_12,In_709,In_519);
nor U13 (N_13,In_90,In_544);
nor U14 (N_14,In_46,In_428);
or U15 (N_15,In_671,In_490);
nand U16 (N_16,In_44,In_638);
nor U17 (N_17,In_75,In_429);
nand U18 (N_18,In_72,In_637);
and U19 (N_19,In_73,In_607);
nand U20 (N_20,In_84,In_28);
or U21 (N_21,In_590,In_178);
xor U22 (N_22,In_634,In_474);
nand U23 (N_23,In_156,In_237);
or U24 (N_24,In_14,In_489);
and U25 (N_25,In_185,In_680);
nor U26 (N_26,In_242,In_191);
and U27 (N_27,In_651,In_582);
and U28 (N_28,In_15,In_7);
and U29 (N_29,In_365,In_226);
or U30 (N_30,In_197,In_278);
nor U31 (N_31,In_211,In_273);
nand U32 (N_32,In_624,In_697);
or U33 (N_33,In_155,In_683);
and U34 (N_34,In_476,In_290);
or U35 (N_35,In_531,In_121);
and U36 (N_36,In_373,In_287);
or U37 (N_37,In_526,In_13);
nand U38 (N_38,In_142,In_605);
nand U39 (N_39,In_417,In_173);
nor U40 (N_40,In_451,In_599);
nand U41 (N_41,In_681,In_189);
and U42 (N_42,In_371,In_678);
and U43 (N_43,In_604,In_375);
nand U44 (N_44,In_55,In_105);
nand U45 (N_45,In_655,In_508);
or U46 (N_46,In_459,In_669);
or U47 (N_47,In_292,In_12);
nor U48 (N_48,In_695,In_684);
and U49 (N_49,In_357,In_466);
nor U50 (N_50,In_547,In_546);
nor U51 (N_51,In_285,In_386);
nand U52 (N_52,In_517,In_201);
nand U53 (N_53,In_253,In_220);
nand U54 (N_54,In_183,In_502);
and U55 (N_55,In_618,In_210);
or U56 (N_56,In_659,In_503);
and U57 (N_57,In_380,In_136);
nand U58 (N_58,In_470,In_550);
and U59 (N_59,In_463,In_652);
xnor U60 (N_60,In_704,In_113);
and U61 (N_61,In_510,In_564);
nor U62 (N_62,In_625,In_88);
and U63 (N_63,In_415,In_109);
nor U64 (N_64,In_92,In_454);
nand U65 (N_65,In_478,In_532);
and U66 (N_66,In_480,In_228);
nor U67 (N_67,In_93,In_140);
or U68 (N_68,In_2,In_686);
nor U69 (N_69,In_555,In_412);
and U70 (N_70,In_218,In_672);
or U71 (N_71,In_694,In_107);
and U72 (N_72,In_658,In_315);
or U73 (N_73,In_536,In_613);
nor U74 (N_74,In_233,In_616);
nand U75 (N_75,In_215,In_376);
nand U76 (N_76,In_79,In_359);
nand U77 (N_77,In_487,In_225);
nand U78 (N_78,In_263,In_56);
nand U79 (N_79,In_453,In_615);
nor U80 (N_80,In_339,In_317);
nor U81 (N_81,In_575,In_356);
and U82 (N_82,In_128,In_736);
or U83 (N_83,In_112,In_322);
and U84 (N_84,In_126,In_268);
nor U85 (N_85,In_527,In_379);
or U86 (N_86,In_494,In_612);
nor U87 (N_87,In_441,In_628);
nand U88 (N_88,In_256,In_633);
and U89 (N_89,In_22,In_350);
nor U90 (N_90,In_170,In_192);
and U91 (N_91,In_654,In_43);
xnor U92 (N_92,In_80,In_469);
xor U93 (N_93,In_588,In_35);
xor U94 (N_94,In_449,In_20);
nor U95 (N_95,In_496,In_366);
or U96 (N_96,In_57,In_110);
and U97 (N_97,In_120,In_563);
nand U98 (N_98,In_161,In_687);
nor U99 (N_99,In_394,In_137);
or U100 (N_100,In_516,In_257);
or U101 (N_101,In_81,In_676);
and U102 (N_102,In_746,In_403);
nor U103 (N_103,In_498,In_741);
and U104 (N_104,In_690,In_343);
and U105 (N_105,In_135,In_304);
and U106 (N_106,In_335,In_323);
nand U107 (N_107,In_21,In_611);
nor U108 (N_108,In_217,In_326);
or U109 (N_109,In_723,In_579);
and U110 (N_110,In_99,In_358);
and U111 (N_111,In_689,In_724);
and U112 (N_112,In_577,In_648);
nand U113 (N_113,In_325,In_311);
and U114 (N_114,In_640,In_32);
and U115 (N_115,In_314,In_103);
or U116 (N_116,In_586,In_398);
or U117 (N_117,In_370,In_61);
and U118 (N_118,In_312,In_83);
xor U119 (N_119,In_167,In_175);
and U120 (N_120,In_608,In_574);
or U121 (N_121,In_172,In_601);
and U122 (N_122,In_702,In_448);
or U123 (N_123,In_435,In_372);
nor U124 (N_124,In_506,In_444);
nor U125 (N_125,In_727,In_713);
nand U126 (N_126,In_195,In_499);
or U127 (N_127,In_205,In_9);
nor U128 (N_128,In_390,In_302);
nand U129 (N_129,In_541,In_632);
nor U130 (N_130,In_742,In_138);
or U131 (N_131,In_533,In_297);
and U132 (N_132,In_129,In_513);
nand U133 (N_133,In_406,In_206);
nand U134 (N_134,In_10,In_250);
and U135 (N_135,In_363,In_53);
or U136 (N_136,In_539,In_700);
nand U137 (N_137,In_647,In_213);
or U138 (N_138,In_60,In_200);
nand U139 (N_139,In_102,In_610);
nand U140 (N_140,In_277,In_246);
nand U141 (N_141,In_298,In_45);
and U142 (N_142,In_324,In_168);
or U143 (N_143,In_229,In_33);
and U144 (N_144,In_447,In_352);
and U145 (N_145,In_348,In_86);
nand U146 (N_146,In_149,In_332);
nor U147 (N_147,In_388,In_492);
nor U148 (N_148,In_653,In_391);
nand U149 (N_149,In_275,In_560);
nand U150 (N_150,In_475,In_421);
and U151 (N_151,In_130,In_342);
nor U152 (N_152,In_208,In_525);
or U153 (N_153,In_708,In_118);
or U154 (N_154,In_67,In_23);
xor U155 (N_155,In_204,In_74);
or U156 (N_156,In_662,In_318);
or U157 (N_157,In_743,In_181);
nor U158 (N_158,In_272,In_196);
or U159 (N_159,In_24,In_207);
nor U160 (N_160,In_212,In_749);
or U161 (N_161,In_606,In_281);
and U162 (N_162,In_5,In_407);
nor U163 (N_163,In_571,In_688);
nor U164 (N_164,In_578,In_271);
and U165 (N_165,In_549,In_642);
nor U166 (N_166,In_561,In_505);
nand U167 (N_167,In_572,In_562);
nand U168 (N_168,In_221,In_300);
or U169 (N_169,In_346,In_8);
nand U170 (N_170,In_733,In_667);
nand U171 (N_171,In_673,In_334);
or U172 (N_172,In_160,In_554);
or U173 (N_173,In_255,In_231);
or U174 (N_174,In_106,In_280);
nand U175 (N_175,In_82,In_286);
nor U176 (N_176,In_402,In_715);
or U177 (N_177,In_739,In_158);
or U178 (N_178,In_523,In_269);
or U179 (N_179,In_666,In_165);
or U180 (N_180,In_157,In_223);
nor U181 (N_181,In_306,In_265);
or U182 (N_182,In_98,In_30);
or U183 (N_183,In_116,In_224);
nor U184 (N_184,In_87,In_392);
and U185 (N_185,In_665,In_726);
or U186 (N_186,In_166,In_276);
nor U187 (N_187,In_552,In_535);
and U188 (N_188,In_133,In_147);
nor U189 (N_189,In_59,In_411);
nand U190 (N_190,In_521,In_674);
nand U191 (N_191,In_62,In_568);
nand U192 (N_192,In_718,In_473);
nand U193 (N_193,In_19,In_94);
and U194 (N_194,In_252,In_626);
nor U195 (N_195,In_31,In_479);
or U196 (N_196,In_11,In_328);
nor U197 (N_197,In_127,In_180);
nand U198 (N_198,In_458,In_202);
nand U199 (N_199,In_51,In_450);
nor U200 (N_200,N_77,N_64);
or U201 (N_201,In_566,In_401);
nor U202 (N_202,In_512,In_509);
nor U203 (N_203,In_714,In_719);
nand U204 (N_204,In_438,N_155);
or U205 (N_205,In_656,In_279);
nor U206 (N_206,In_260,In_425);
or U207 (N_207,N_184,N_80);
xor U208 (N_208,In_150,N_68);
and U209 (N_209,In_301,In_1);
xor U210 (N_210,N_23,N_75);
or U211 (N_211,In_289,N_185);
nand U212 (N_212,N_31,N_122);
and U213 (N_213,In_725,In_493);
and U214 (N_214,In_239,In_663);
or U215 (N_215,N_90,In_420);
nor U216 (N_216,In_36,In_703);
nand U217 (N_217,N_22,In_48);
or U218 (N_218,N_3,In_511);
nand U219 (N_219,In_293,In_691);
and U220 (N_220,In_468,In_364);
nor U221 (N_221,N_25,In_426);
nor U222 (N_222,N_91,In_179);
and U223 (N_223,In_596,In_591);
nand U224 (N_224,N_52,In_182);
or U225 (N_225,N_7,N_87);
or U226 (N_226,In_261,In_330);
or U227 (N_227,In_491,In_153);
or U228 (N_228,In_485,In_565);
nor U229 (N_229,In_345,In_661);
or U230 (N_230,In_528,In_69);
nor U231 (N_231,N_97,In_501);
nor U232 (N_232,In_436,N_195);
nand U233 (N_233,N_189,In_396);
nor U234 (N_234,In_437,In_518);
nor U235 (N_235,N_71,In_631);
or U236 (N_236,In_177,In_668);
and U237 (N_237,N_120,N_73);
and U238 (N_238,In_488,N_99);
and U239 (N_239,N_1,In_484);
and U240 (N_240,In_132,In_620);
nor U241 (N_241,In_405,In_679);
nor U242 (N_242,In_481,In_594);
and U243 (N_243,N_86,N_163);
nand U244 (N_244,In_47,In_685);
nand U245 (N_245,N_58,In_592);
or U246 (N_246,In_699,N_104);
nand U247 (N_247,In_557,In_465);
nand U248 (N_248,In_698,In_583);
nor U249 (N_249,In_321,In_299);
and U250 (N_250,In_198,In_537);
nand U251 (N_251,In_97,In_559);
xnor U252 (N_252,In_416,In_483);
and U253 (N_253,In_40,In_467);
nor U254 (N_254,N_59,N_61);
or U255 (N_255,In_209,In_529);
and U256 (N_256,N_191,N_112);
or U257 (N_257,N_67,N_100);
nand U258 (N_258,In_65,N_56);
and U259 (N_259,In_455,N_124);
nand U260 (N_260,In_646,In_216);
nand U261 (N_261,In_734,In_593);
or U262 (N_262,In_163,N_116);
nor U263 (N_263,In_545,In_515);
nand U264 (N_264,N_160,In_117);
and U265 (N_265,In_383,N_103);
xor U266 (N_266,In_721,N_130);
xor U267 (N_267,N_156,In_248);
or U268 (N_268,N_158,N_186);
nor U269 (N_269,In_139,In_96);
nor U270 (N_270,In_717,N_39);
nand U271 (N_271,In_433,N_149);
and U272 (N_272,In_29,In_657);
or U273 (N_273,N_151,In_602);
nand U274 (N_274,In_187,In_63);
nand U275 (N_275,In_682,N_55);
or U276 (N_276,N_2,In_354);
or U277 (N_277,In_692,N_96);
nand U278 (N_278,In_235,In_122);
or U279 (N_279,N_43,N_132);
nand U280 (N_280,N_178,In_567);
or U281 (N_281,N_107,N_102);
nand U282 (N_282,In_598,N_117);
nor U283 (N_283,In_570,In_452);
or U284 (N_284,N_44,In_381);
and U285 (N_285,N_41,In_744);
nand U286 (N_286,In_341,N_4);
and U287 (N_287,In_675,In_431);
nand U288 (N_288,N_111,In_639);
nand U289 (N_289,In_184,N_114);
and U290 (N_290,In_446,In_308);
nor U291 (N_291,N_27,N_175);
or U292 (N_292,In_630,In_188);
or U293 (N_293,N_144,In_551);
nand U294 (N_294,N_50,In_664);
or U295 (N_295,N_159,In_422);
or U296 (N_296,N_162,N_48);
or U297 (N_297,N_167,N_92);
and U298 (N_298,In_442,N_115);
nand U299 (N_299,In_635,In_123);
nor U300 (N_300,N_119,N_69);
or U301 (N_301,In_58,N_150);
and U302 (N_302,In_349,In_729);
or U303 (N_303,N_142,N_154);
and U304 (N_304,In_274,In_738);
nor U305 (N_305,N_135,In_387);
and U306 (N_306,In_711,N_165);
and U307 (N_307,In_410,N_110);
nand U308 (N_308,In_264,In_696);
and U309 (N_309,In_146,In_38);
or U310 (N_310,In_740,N_76);
or U311 (N_311,In_85,N_190);
nand U312 (N_312,In_440,N_16);
and U313 (N_313,N_109,In_303);
nor U314 (N_314,N_5,N_169);
or U315 (N_315,N_113,N_14);
or U316 (N_316,In_145,N_177);
or U317 (N_317,N_53,In_482);
and U318 (N_318,In_369,N_172);
nand U319 (N_319,In_39,In_558);
and U320 (N_320,In_385,In_748);
nor U321 (N_321,In_423,In_234);
nor U322 (N_322,In_336,In_514);
and U323 (N_323,N_29,N_133);
nand U324 (N_324,In_553,In_645);
nand U325 (N_325,In_222,In_238);
nor U326 (N_326,In_413,In_50);
nand U327 (N_327,In_266,In_362);
and U328 (N_328,N_136,N_131);
or U329 (N_329,In_712,In_331);
xnor U330 (N_330,In_504,N_152);
nand U331 (N_331,In_745,In_240);
nor U332 (N_332,In_171,In_462);
xor U333 (N_333,N_40,In_310);
nand U334 (N_334,In_18,In_267);
nor U335 (N_335,In_259,In_159);
and U336 (N_336,In_64,In_585);
nand U337 (N_337,In_115,N_63);
or U338 (N_338,N_143,In_542);
or U339 (N_339,N_79,In_219);
nand U340 (N_340,In_445,N_11);
or U341 (N_341,In_186,In_730);
nand U342 (N_342,N_128,In_374);
xor U343 (N_343,In_456,In_520);
nor U344 (N_344,N_65,In_486);
nand U345 (N_345,In_95,In_0);
nor U346 (N_346,N_145,In_495);
and U347 (N_347,In_731,N_192);
nor U348 (N_348,N_60,In_101);
and U349 (N_349,In_430,In_377);
nor U350 (N_350,In_91,In_534);
and U351 (N_351,In_581,N_30);
or U352 (N_352,In_621,In_154);
and U353 (N_353,In_728,In_337);
or U354 (N_354,In_309,In_644);
nor U355 (N_355,N_147,In_706);
or U356 (N_356,In_609,In_355);
or U357 (N_357,In_477,In_507);
nor U358 (N_358,In_125,In_397);
nand U359 (N_359,N_161,In_162);
nand U360 (N_360,In_236,In_409);
and U361 (N_361,In_66,In_243);
nand U362 (N_362,N_8,N_45);
or U363 (N_363,N_197,In_89);
and U364 (N_364,In_254,N_196);
nor U365 (N_365,N_28,In_307);
and U366 (N_366,In_548,In_4);
or U367 (N_367,N_170,In_148);
nand U368 (N_368,In_25,N_194);
nand U369 (N_369,In_408,N_179);
or U370 (N_370,N_164,In_124);
and U371 (N_371,In_580,N_93);
nor U372 (N_372,In_327,In_595);
nor U373 (N_373,N_126,In_427);
and U374 (N_374,In_569,In_747);
or U375 (N_375,In_284,In_587);
nor U376 (N_376,In_660,In_540);
or U377 (N_377,In_617,In_641);
nand U378 (N_378,In_340,N_95);
nor U379 (N_379,In_584,In_313);
xor U380 (N_380,In_368,N_33);
or U381 (N_381,N_168,N_66);
or U382 (N_382,N_139,N_141);
nand U383 (N_383,N_146,In_176);
nand U384 (N_384,N_88,In_461);
and U385 (N_385,N_101,In_320);
or U386 (N_386,N_15,N_54);
nor U387 (N_387,N_62,N_85);
or U388 (N_388,N_24,N_17);
nor U389 (N_389,In_6,N_121);
nand U390 (N_390,N_78,In_52);
or U391 (N_391,In_597,In_119);
or U392 (N_392,N_123,In_190);
nand U393 (N_393,N_6,In_247);
nand U394 (N_394,N_129,In_732);
and U395 (N_395,In_424,In_693);
nand U396 (N_396,In_378,N_19);
nand U397 (N_397,In_353,N_34);
or U398 (N_398,In_251,In_230);
and U399 (N_399,In_522,In_144);
nor U400 (N_400,N_344,N_399);
and U401 (N_401,N_338,In_164);
nand U402 (N_402,N_232,N_258);
and U403 (N_403,N_216,N_313);
or U404 (N_404,In_344,N_286);
nand U405 (N_405,In_556,In_434);
nand U406 (N_406,N_312,N_397);
nor U407 (N_407,N_74,In_443);
or U408 (N_408,N_84,N_108);
and U409 (N_409,N_381,N_94);
nand U410 (N_410,In_457,In_41);
nor U411 (N_411,N_297,In_131);
and U412 (N_412,N_275,N_317);
nor U413 (N_413,N_208,In_227);
or U414 (N_414,In_393,In_270);
nand U415 (N_415,N_244,N_398);
nor U416 (N_416,N_82,N_362);
and U417 (N_417,N_310,N_336);
nor U418 (N_418,In_432,N_276);
and U419 (N_419,N_322,N_292);
nand U420 (N_420,In_319,N_347);
and U421 (N_421,N_212,N_203);
nor U422 (N_422,N_254,In_614);
or U423 (N_423,In_530,N_273);
and U424 (N_424,N_188,N_346);
or U425 (N_425,In_54,N_393);
or U426 (N_426,N_385,N_199);
and U427 (N_427,N_183,N_251);
or U428 (N_428,N_9,N_301);
or U429 (N_429,N_35,N_390);
nor U430 (N_430,In_395,N_348);
or U431 (N_431,N_173,N_304);
nor U432 (N_432,N_321,N_382);
nor U433 (N_433,N_298,N_118);
and U434 (N_434,N_315,N_361);
and U435 (N_435,N_372,N_370);
and U436 (N_436,N_307,N_371);
or U437 (N_437,N_256,N_243);
or U438 (N_438,N_269,N_51);
nor U439 (N_439,N_289,N_350);
nand U440 (N_440,N_246,N_140);
or U441 (N_441,N_284,N_200);
or U442 (N_442,N_280,N_396);
nand U443 (N_443,N_323,In_288);
nor U444 (N_444,N_89,N_288);
nand U445 (N_445,N_320,N_13);
nand U446 (N_446,N_153,N_283);
xnor U447 (N_447,N_180,N_277);
nor U448 (N_448,N_330,In_701);
and U449 (N_449,N_314,N_296);
nor U450 (N_450,In_367,In_26);
nor U451 (N_451,In_705,N_0);
nand U452 (N_452,N_358,In_464);
or U453 (N_453,In_589,N_220);
nor U454 (N_454,In_245,N_237);
and U455 (N_455,N_227,N_238);
and U456 (N_456,N_72,N_334);
or U457 (N_457,N_264,N_166);
nand U458 (N_458,N_386,N_255);
or U459 (N_459,N_324,N_377);
nand U460 (N_460,N_222,In_389);
nor U461 (N_461,N_217,In_351);
and U462 (N_462,N_105,N_305);
and U463 (N_463,In_497,In_143);
nor U464 (N_464,N_295,In_244);
or U465 (N_465,N_294,N_46);
nor U466 (N_466,N_378,N_300);
or U467 (N_467,In_151,N_209);
nor U468 (N_468,In_735,In_623);
nand U469 (N_469,N_225,In_76);
and U470 (N_470,N_271,N_319);
xnor U471 (N_471,N_327,N_234);
or U472 (N_472,N_228,N_70);
nor U473 (N_473,N_260,N_37);
and U474 (N_474,In_573,In_329);
nand U475 (N_475,N_356,N_215);
nand U476 (N_476,N_268,In_418);
nor U477 (N_477,N_302,N_389);
nand U478 (N_478,N_206,N_270);
nor U479 (N_479,In_295,In_78);
nor U480 (N_480,N_354,In_333);
nor U481 (N_481,N_32,In_111);
or U482 (N_482,N_279,N_221);
or U483 (N_483,In_399,N_281);
xor U484 (N_484,N_360,N_214);
or U485 (N_485,In_543,N_303);
and U486 (N_486,In_603,N_211);
nor U487 (N_487,N_308,N_125);
nand U488 (N_488,N_242,N_249);
nor U489 (N_489,N_337,N_329);
or U490 (N_490,N_207,N_98);
nor U491 (N_491,In_338,N_252);
nand U492 (N_492,In_193,N_335);
nor U493 (N_493,N_49,N_369);
and U494 (N_494,N_21,In_37);
and U495 (N_495,In_720,In_249);
and U496 (N_496,N_325,N_198);
and U497 (N_497,N_379,N_331);
nand U498 (N_498,N_213,N_230);
nand U499 (N_499,In_360,N_374);
and U500 (N_500,In_108,In_114);
nor U501 (N_501,N_223,N_394);
nand U502 (N_502,N_253,In_400);
or U503 (N_503,N_218,N_343);
nor U504 (N_504,N_387,N_359);
nor U505 (N_505,In_68,N_193);
nor U506 (N_506,N_257,N_247);
nand U507 (N_507,N_388,N_328);
nor U508 (N_508,In_619,N_26);
and U509 (N_509,N_42,In_472);
nand U510 (N_510,N_375,N_299);
or U511 (N_511,N_182,In_42);
and U512 (N_512,N_205,N_81);
nor U513 (N_513,N_248,In_152);
xor U514 (N_514,N_345,N_47);
nand U515 (N_515,In_71,In_347);
nand U516 (N_516,N_20,In_305);
or U517 (N_517,N_181,In_258);
and U518 (N_518,N_363,N_266);
nor U519 (N_519,N_290,N_148);
and U520 (N_520,N_341,In_737);
or U521 (N_521,N_287,N_137);
and U522 (N_522,N_395,N_57);
nor U523 (N_523,In_670,N_368);
nand U524 (N_524,In_500,N_236);
or U525 (N_525,N_127,N_274);
nand U526 (N_526,N_339,N_171);
and U527 (N_527,In_100,N_351);
and U528 (N_528,In_627,N_259);
and U529 (N_529,N_380,In_27);
nor U530 (N_530,N_278,In_649);
nand U531 (N_531,N_383,In_282);
or U532 (N_532,N_333,In_722);
and U533 (N_533,N_176,N_134);
nor U534 (N_534,In_291,In_77);
nand U535 (N_535,N_201,In_169);
and U536 (N_536,N_326,N_226);
or U537 (N_537,In_241,N_272);
and U538 (N_538,N_187,N_250);
nand U539 (N_539,N_293,N_355);
and U540 (N_540,N_263,N_83);
nor U541 (N_541,N_229,In_134);
nor U542 (N_542,N_204,N_384);
and U543 (N_543,N_240,N_18);
or U544 (N_544,In_141,N_342);
or U545 (N_545,N_235,N_291);
nand U546 (N_546,In_16,In_419);
nand U547 (N_547,N_241,N_202);
xnor U548 (N_548,N_239,N_340);
nor U549 (N_549,N_353,N_357);
and U550 (N_550,N_366,N_233);
or U551 (N_551,In_361,In_49);
nor U552 (N_552,N_245,N_306);
or U553 (N_553,N_364,N_10);
nor U554 (N_554,In_194,N_265);
nand U555 (N_555,In_384,In_262);
or U556 (N_556,N_174,N_219);
nand U557 (N_557,N_138,N_231);
or U558 (N_558,N_392,N_267);
nand U559 (N_559,In_636,N_282);
nand U560 (N_560,N_262,N_332);
nand U561 (N_561,In_524,In_296);
nor U562 (N_562,N_210,N_352);
or U563 (N_563,N_318,N_373);
and U564 (N_564,In_404,N_157);
nand U565 (N_565,N_391,N_309);
or U566 (N_566,N_12,N_367);
and U567 (N_567,N_224,N_38);
or U568 (N_568,In_294,In_414);
and U569 (N_569,N_316,N_311);
nor U570 (N_570,N_106,N_285);
and U571 (N_571,N_36,In_629);
nor U572 (N_572,N_349,N_365);
or U573 (N_573,N_261,N_376);
xor U574 (N_574,In_650,In_622);
nor U575 (N_575,N_290,N_344);
nand U576 (N_576,N_298,N_391);
nor U577 (N_577,In_720,N_249);
nand U578 (N_578,N_323,N_297);
or U579 (N_579,N_211,N_157);
and U580 (N_580,N_237,N_241);
or U581 (N_581,N_72,In_245);
nor U582 (N_582,N_307,In_650);
xnor U583 (N_583,N_314,N_216);
or U584 (N_584,N_335,N_222);
or U585 (N_585,N_0,N_342);
nand U586 (N_586,N_384,N_205);
nand U587 (N_587,N_345,N_206);
or U588 (N_588,N_279,N_287);
nand U589 (N_589,In_722,N_348);
or U590 (N_590,N_392,N_379);
or U591 (N_591,N_285,N_390);
and U592 (N_592,N_245,N_89);
nor U593 (N_593,N_272,N_327);
and U594 (N_594,In_169,In_291);
or U595 (N_595,N_212,N_395);
nand U596 (N_596,N_202,N_385);
and U597 (N_597,N_383,In_169);
and U598 (N_598,In_111,In_288);
nor U599 (N_599,N_296,N_229);
nand U600 (N_600,N_430,N_562);
nand U601 (N_601,N_574,N_442);
or U602 (N_602,N_417,N_493);
and U603 (N_603,N_412,N_481);
and U604 (N_604,N_587,N_454);
and U605 (N_605,N_411,N_579);
nand U606 (N_606,N_443,N_451);
nand U607 (N_607,N_536,N_463);
or U608 (N_608,N_457,N_419);
and U609 (N_609,N_471,N_427);
or U610 (N_610,N_588,N_473);
or U611 (N_611,N_445,N_597);
or U612 (N_612,N_566,N_549);
and U613 (N_613,N_494,N_534);
nand U614 (N_614,N_528,N_472);
and U615 (N_615,N_516,N_543);
nand U616 (N_616,N_533,N_462);
nand U617 (N_617,N_489,N_487);
nor U618 (N_618,N_467,N_475);
nor U619 (N_619,N_551,N_586);
or U620 (N_620,N_582,N_482);
or U621 (N_621,N_416,N_595);
and U622 (N_622,N_418,N_581);
nand U623 (N_623,N_450,N_490);
and U624 (N_624,N_422,N_440);
nand U625 (N_625,N_437,N_537);
nand U626 (N_626,N_514,N_453);
or U627 (N_627,N_441,N_452);
and U628 (N_628,N_464,N_403);
nor U629 (N_629,N_518,N_477);
nor U630 (N_630,N_401,N_438);
and U631 (N_631,N_448,N_492);
and U632 (N_632,N_527,N_599);
nor U633 (N_633,N_592,N_577);
or U634 (N_634,N_569,N_436);
nor U635 (N_635,N_415,N_555);
or U636 (N_636,N_540,N_486);
and U637 (N_637,N_515,N_575);
nor U638 (N_638,N_425,N_439);
nand U639 (N_639,N_589,N_408);
nand U640 (N_640,N_433,N_404);
or U641 (N_641,N_512,N_447);
nand U642 (N_642,N_402,N_495);
or U643 (N_643,N_478,N_524);
nand U644 (N_644,N_497,N_421);
nor U645 (N_645,N_572,N_550);
or U646 (N_646,N_585,N_470);
and U647 (N_647,N_558,N_517);
nor U648 (N_648,N_520,N_499);
and U649 (N_649,N_508,N_510);
nor U650 (N_650,N_500,N_590);
or U651 (N_651,N_519,N_544);
and U652 (N_652,N_431,N_598);
xnor U653 (N_653,N_584,N_563);
and U654 (N_654,N_541,N_531);
nor U655 (N_655,N_560,N_444);
nand U656 (N_656,N_458,N_409);
or U657 (N_657,N_591,N_428);
or U658 (N_658,N_465,N_542);
or U659 (N_659,N_511,N_567);
and U660 (N_660,N_571,N_460);
nand U661 (N_661,N_545,N_506);
or U662 (N_662,N_580,N_459);
or U663 (N_663,N_406,N_523);
and U664 (N_664,N_434,N_414);
nand U665 (N_665,N_535,N_413);
or U666 (N_666,N_480,N_556);
or U667 (N_667,N_570,N_539);
nor U668 (N_668,N_559,N_484);
xor U669 (N_669,N_505,N_507);
and U670 (N_670,N_468,N_446);
or U671 (N_671,N_496,N_522);
or U672 (N_672,N_538,N_564);
nand U673 (N_673,N_491,N_532);
or U674 (N_674,N_498,N_521);
and U675 (N_675,N_449,N_420);
or U676 (N_676,N_525,N_483);
nand U677 (N_677,N_568,N_432);
nand U678 (N_678,N_546,N_565);
and U679 (N_679,N_469,N_547);
and U680 (N_680,N_461,N_400);
nand U681 (N_681,N_502,N_593);
and U682 (N_682,N_530,N_426);
xnor U683 (N_683,N_424,N_410);
nand U684 (N_684,N_573,N_576);
nand U685 (N_685,N_429,N_455);
and U686 (N_686,N_435,N_485);
and U687 (N_687,N_594,N_548);
or U688 (N_688,N_583,N_504);
xor U689 (N_689,N_578,N_513);
or U690 (N_690,N_456,N_423);
nor U691 (N_691,N_474,N_479);
or U692 (N_692,N_407,N_501);
nor U693 (N_693,N_596,N_509);
or U694 (N_694,N_554,N_476);
or U695 (N_695,N_405,N_488);
nand U696 (N_696,N_526,N_557);
or U697 (N_697,N_561,N_466);
nor U698 (N_698,N_503,N_552);
nand U699 (N_699,N_529,N_553);
and U700 (N_700,N_410,N_576);
or U701 (N_701,N_448,N_592);
or U702 (N_702,N_539,N_577);
and U703 (N_703,N_439,N_411);
nand U704 (N_704,N_459,N_506);
and U705 (N_705,N_597,N_411);
or U706 (N_706,N_565,N_494);
xor U707 (N_707,N_503,N_414);
and U708 (N_708,N_543,N_527);
or U709 (N_709,N_537,N_524);
nand U710 (N_710,N_503,N_567);
nor U711 (N_711,N_565,N_457);
and U712 (N_712,N_588,N_557);
and U713 (N_713,N_574,N_483);
nor U714 (N_714,N_414,N_579);
nand U715 (N_715,N_491,N_456);
or U716 (N_716,N_591,N_561);
nand U717 (N_717,N_421,N_564);
and U718 (N_718,N_530,N_492);
or U719 (N_719,N_506,N_535);
or U720 (N_720,N_495,N_508);
or U721 (N_721,N_562,N_415);
or U722 (N_722,N_501,N_465);
nand U723 (N_723,N_496,N_543);
nor U724 (N_724,N_429,N_408);
xnor U725 (N_725,N_506,N_596);
and U726 (N_726,N_470,N_409);
or U727 (N_727,N_537,N_470);
and U728 (N_728,N_425,N_400);
and U729 (N_729,N_552,N_548);
nand U730 (N_730,N_453,N_590);
and U731 (N_731,N_405,N_521);
nand U732 (N_732,N_431,N_563);
and U733 (N_733,N_479,N_583);
nand U734 (N_734,N_552,N_546);
or U735 (N_735,N_404,N_571);
or U736 (N_736,N_562,N_490);
xor U737 (N_737,N_550,N_423);
xnor U738 (N_738,N_568,N_450);
or U739 (N_739,N_452,N_516);
and U740 (N_740,N_407,N_558);
nand U741 (N_741,N_442,N_509);
nor U742 (N_742,N_454,N_552);
or U743 (N_743,N_481,N_559);
or U744 (N_744,N_480,N_444);
and U745 (N_745,N_492,N_486);
and U746 (N_746,N_445,N_555);
nand U747 (N_747,N_417,N_499);
xnor U748 (N_748,N_410,N_440);
xnor U749 (N_749,N_500,N_408);
nor U750 (N_750,N_502,N_410);
nand U751 (N_751,N_482,N_441);
nor U752 (N_752,N_421,N_538);
or U753 (N_753,N_466,N_578);
and U754 (N_754,N_486,N_496);
or U755 (N_755,N_409,N_449);
and U756 (N_756,N_455,N_438);
nand U757 (N_757,N_511,N_432);
nand U758 (N_758,N_502,N_437);
nor U759 (N_759,N_405,N_595);
nor U760 (N_760,N_455,N_451);
nand U761 (N_761,N_522,N_555);
and U762 (N_762,N_518,N_454);
nand U763 (N_763,N_497,N_564);
nor U764 (N_764,N_547,N_559);
or U765 (N_765,N_583,N_574);
and U766 (N_766,N_576,N_591);
nor U767 (N_767,N_543,N_541);
nand U768 (N_768,N_421,N_560);
or U769 (N_769,N_420,N_467);
and U770 (N_770,N_419,N_485);
or U771 (N_771,N_573,N_408);
nor U772 (N_772,N_495,N_541);
nor U773 (N_773,N_493,N_432);
or U774 (N_774,N_452,N_424);
or U775 (N_775,N_461,N_579);
or U776 (N_776,N_536,N_532);
or U777 (N_777,N_483,N_590);
nor U778 (N_778,N_574,N_410);
and U779 (N_779,N_488,N_471);
nand U780 (N_780,N_408,N_413);
or U781 (N_781,N_583,N_461);
nor U782 (N_782,N_488,N_511);
nand U783 (N_783,N_401,N_537);
xnor U784 (N_784,N_485,N_563);
nor U785 (N_785,N_537,N_448);
nand U786 (N_786,N_465,N_477);
or U787 (N_787,N_502,N_455);
and U788 (N_788,N_508,N_497);
nor U789 (N_789,N_540,N_555);
and U790 (N_790,N_520,N_506);
or U791 (N_791,N_459,N_500);
nand U792 (N_792,N_519,N_438);
nor U793 (N_793,N_577,N_452);
or U794 (N_794,N_455,N_581);
nand U795 (N_795,N_451,N_465);
nand U796 (N_796,N_509,N_439);
nand U797 (N_797,N_581,N_520);
nand U798 (N_798,N_582,N_512);
or U799 (N_799,N_524,N_597);
and U800 (N_800,N_736,N_607);
nand U801 (N_801,N_724,N_770);
and U802 (N_802,N_777,N_663);
nor U803 (N_803,N_690,N_750);
nor U804 (N_804,N_665,N_629);
and U805 (N_805,N_788,N_696);
or U806 (N_806,N_605,N_766);
nor U807 (N_807,N_742,N_717);
nand U808 (N_808,N_687,N_704);
nand U809 (N_809,N_713,N_721);
nand U810 (N_810,N_727,N_772);
or U811 (N_811,N_719,N_796);
nand U812 (N_812,N_695,N_739);
and U813 (N_813,N_723,N_706);
or U814 (N_814,N_753,N_653);
nand U815 (N_815,N_678,N_793);
and U816 (N_816,N_748,N_685);
nor U817 (N_817,N_784,N_708);
nor U818 (N_818,N_670,N_794);
nor U819 (N_819,N_632,N_751);
nor U820 (N_820,N_780,N_700);
nand U821 (N_821,N_641,N_759);
nor U822 (N_822,N_684,N_631);
and U823 (N_823,N_611,N_646);
and U824 (N_824,N_762,N_640);
and U825 (N_825,N_621,N_636);
xnor U826 (N_826,N_712,N_740);
nor U827 (N_827,N_707,N_789);
and U828 (N_828,N_741,N_764);
nor U829 (N_829,N_783,N_656);
nand U830 (N_830,N_697,N_725);
nor U831 (N_831,N_676,N_643);
or U832 (N_832,N_603,N_668);
nor U833 (N_833,N_658,N_767);
nand U834 (N_834,N_768,N_699);
and U835 (N_835,N_617,N_672);
or U836 (N_836,N_771,N_642);
nor U837 (N_837,N_667,N_775);
nor U838 (N_838,N_756,N_635);
or U839 (N_839,N_730,N_701);
nor U840 (N_840,N_720,N_675);
nor U841 (N_841,N_614,N_798);
nor U842 (N_842,N_630,N_639);
nor U843 (N_843,N_735,N_660);
nor U844 (N_844,N_662,N_615);
and U845 (N_845,N_619,N_681);
xor U846 (N_846,N_627,N_623);
nand U847 (N_847,N_715,N_743);
and U848 (N_848,N_792,N_761);
or U849 (N_849,N_638,N_781);
nor U850 (N_850,N_738,N_674);
and U851 (N_851,N_757,N_763);
nand U852 (N_852,N_673,N_671);
nor U853 (N_853,N_749,N_722);
nand U854 (N_854,N_683,N_732);
or U855 (N_855,N_791,N_774);
nor U856 (N_856,N_659,N_785);
and U857 (N_857,N_729,N_797);
nand U858 (N_858,N_604,N_733);
nand U859 (N_859,N_679,N_714);
nor U860 (N_860,N_666,N_645);
or U861 (N_861,N_693,N_705);
nand U862 (N_862,N_652,N_716);
nor U863 (N_863,N_664,N_694);
or U864 (N_864,N_692,N_612);
nand U865 (N_865,N_769,N_610);
nor U866 (N_866,N_609,N_649);
nor U867 (N_867,N_747,N_710);
and U868 (N_868,N_731,N_795);
or U869 (N_869,N_600,N_778);
and U870 (N_870,N_786,N_625);
or U871 (N_871,N_702,N_765);
nand U872 (N_872,N_752,N_628);
nand U873 (N_873,N_728,N_620);
or U874 (N_874,N_626,N_650);
nor U875 (N_875,N_624,N_654);
and U876 (N_876,N_644,N_754);
nand U877 (N_877,N_776,N_703);
or U878 (N_878,N_709,N_682);
and U879 (N_879,N_634,N_613);
or U880 (N_880,N_618,N_608);
or U881 (N_881,N_773,N_746);
nor U882 (N_882,N_755,N_686);
and U883 (N_883,N_657,N_760);
or U884 (N_884,N_637,N_787);
nand U885 (N_885,N_799,N_779);
nor U886 (N_886,N_745,N_655);
or U887 (N_887,N_698,N_790);
and U888 (N_888,N_689,N_734);
nor U889 (N_889,N_782,N_758);
and U890 (N_890,N_633,N_718);
and U891 (N_891,N_688,N_648);
or U892 (N_892,N_744,N_677);
nor U893 (N_893,N_651,N_711);
or U894 (N_894,N_737,N_602);
and U895 (N_895,N_661,N_616);
or U896 (N_896,N_606,N_601);
xor U897 (N_897,N_726,N_622);
nand U898 (N_898,N_691,N_680);
nor U899 (N_899,N_669,N_647);
or U900 (N_900,N_701,N_746);
nor U901 (N_901,N_634,N_633);
and U902 (N_902,N_653,N_752);
nand U903 (N_903,N_611,N_647);
nor U904 (N_904,N_768,N_721);
xor U905 (N_905,N_651,N_637);
and U906 (N_906,N_736,N_671);
or U907 (N_907,N_618,N_698);
nand U908 (N_908,N_779,N_733);
nor U909 (N_909,N_729,N_637);
and U910 (N_910,N_708,N_757);
nor U911 (N_911,N_766,N_756);
nor U912 (N_912,N_662,N_790);
or U913 (N_913,N_785,N_769);
nand U914 (N_914,N_736,N_724);
and U915 (N_915,N_708,N_731);
nand U916 (N_916,N_735,N_788);
nor U917 (N_917,N_796,N_639);
nand U918 (N_918,N_670,N_775);
nand U919 (N_919,N_674,N_616);
or U920 (N_920,N_686,N_761);
or U921 (N_921,N_674,N_610);
or U922 (N_922,N_798,N_690);
or U923 (N_923,N_728,N_744);
or U924 (N_924,N_621,N_773);
or U925 (N_925,N_708,N_680);
and U926 (N_926,N_752,N_686);
nand U927 (N_927,N_723,N_661);
and U928 (N_928,N_789,N_764);
nor U929 (N_929,N_725,N_683);
and U930 (N_930,N_780,N_692);
and U931 (N_931,N_608,N_668);
nor U932 (N_932,N_781,N_676);
nor U933 (N_933,N_739,N_742);
nand U934 (N_934,N_770,N_700);
nand U935 (N_935,N_671,N_640);
or U936 (N_936,N_636,N_653);
nand U937 (N_937,N_719,N_652);
nand U938 (N_938,N_686,N_749);
nand U939 (N_939,N_645,N_604);
and U940 (N_940,N_668,N_625);
or U941 (N_941,N_721,N_691);
or U942 (N_942,N_771,N_755);
nand U943 (N_943,N_743,N_789);
and U944 (N_944,N_636,N_788);
or U945 (N_945,N_767,N_652);
or U946 (N_946,N_626,N_604);
xor U947 (N_947,N_680,N_747);
or U948 (N_948,N_725,N_616);
nor U949 (N_949,N_737,N_606);
or U950 (N_950,N_736,N_617);
and U951 (N_951,N_621,N_614);
and U952 (N_952,N_767,N_736);
and U953 (N_953,N_635,N_608);
nand U954 (N_954,N_759,N_651);
and U955 (N_955,N_668,N_712);
nor U956 (N_956,N_774,N_601);
nor U957 (N_957,N_601,N_760);
nand U958 (N_958,N_646,N_600);
nand U959 (N_959,N_763,N_663);
or U960 (N_960,N_628,N_770);
nand U961 (N_961,N_785,N_691);
and U962 (N_962,N_739,N_774);
xnor U963 (N_963,N_730,N_685);
nand U964 (N_964,N_689,N_779);
and U965 (N_965,N_703,N_775);
nor U966 (N_966,N_614,N_694);
and U967 (N_967,N_640,N_668);
nor U968 (N_968,N_636,N_684);
and U969 (N_969,N_676,N_746);
nor U970 (N_970,N_732,N_673);
nor U971 (N_971,N_774,N_737);
nand U972 (N_972,N_766,N_714);
or U973 (N_973,N_606,N_642);
xnor U974 (N_974,N_749,N_693);
and U975 (N_975,N_710,N_705);
nand U976 (N_976,N_643,N_645);
and U977 (N_977,N_681,N_651);
nor U978 (N_978,N_734,N_635);
nor U979 (N_979,N_624,N_621);
or U980 (N_980,N_675,N_739);
nand U981 (N_981,N_716,N_784);
or U982 (N_982,N_775,N_613);
and U983 (N_983,N_680,N_693);
nand U984 (N_984,N_710,N_693);
and U985 (N_985,N_783,N_637);
xor U986 (N_986,N_776,N_791);
and U987 (N_987,N_648,N_684);
and U988 (N_988,N_655,N_674);
and U989 (N_989,N_694,N_612);
nor U990 (N_990,N_664,N_725);
or U991 (N_991,N_670,N_624);
and U992 (N_992,N_704,N_640);
nor U993 (N_993,N_676,N_791);
and U994 (N_994,N_789,N_767);
and U995 (N_995,N_660,N_773);
nor U996 (N_996,N_780,N_719);
nor U997 (N_997,N_724,N_729);
nor U998 (N_998,N_775,N_655);
or U999 (N_999,N_703,N_684);
nand U1000 (N_1000,N_974,N_874);
nor U1001 (N_1001,N_800,N_868);
nand U1002 (N_1002,N_946,N_987);
nor U1003 (N_1003,N_847,N_842);
or U1004 (N_1004,N_919,N_840);
and U1005 (N_1005,N_837,N_979);
or U1006 (N_1006,N_869,N_852);
xnor U1007 (N_1007,N_918,N_948);
nand U1008 (N_1008,N_932,N_975);
and U1009 (N_1009,N_968,N_831);
and U1010 (N_1010,N_835,N_970);
nor U1011 (N_1011,N_870,N_891);
and U1012 (N_1012,N_862,N_923);
or U1013 (N_1013,N_810,N_957);
nand U1014 (N_1014,N_882,N_899);
or U1015 (N_1015,N_898,N_966);
nor U1016 (N_1016,N_942,N_982);
xnor U1017 (N_1017,N_836,N_865);
or U1018 (N_1018,N_990,N_993);
and U1019 (N_1019,N_821,N_921);
nand U1020 (N_1020,N_926,N_927);
or U1021 (N_1021,N_901,N_943);
nand U1022 (N_1022,N_910,N_886);
and U1023 (N_1023,N_823,N_839);
or U1024 (N_1024,N_965,N_929);
and U1025 (N_1025,N_834,N_995);
nor U1026 (N_1026,N_955,N_854);
or U1027 (N_1027,N_937,N_888);
or U1028 (N_1028,N_963,N_801);
and U1029 (N_1029,N_947,N_833);
or U1030 (N_1030,N_879,N_817);
nand U1031 (N_1031,N_900,N_972);
or U1032 (N_1032,N_892,N_904);
nor U1033 (N_1033,N_895,N_941);
nor U1034 (N_1034,N_939,N_832);
xor U1035 (N_1035,N_804,N_952);
nor U1036 (N_1036,N_997,N_911);
nor U1037 (N_1037,N_885,N_916);
and U1038 (N_1038,N_820,N_934);
nand U1039 (N_1039,N_983,N_838);
nor U1040 (N_1040,N_962,N_944);
nor U1041 (N_1041,N_878,N_897);
or U1042 (N_1042,N_826,N_864);
nand U1043 (N_1043,N_913,N_851);
or U1044 (N_1044,N_920,N_863);
or U1045 (N_1045,N_848,N_805);
nand U1046 (N_1046,N_860,N_813);
and U1047 (N_1047,N_917,N_845);
or U1048 (N_1048,N_871,N_950);
and U1049 (N_1049,N_827,N_954);
or U1050 (N_1050,N_930,N_802);
or U1051 (N_1051,N_998,N_841);
or U1052 (N_1052,N_956,N_857);
nand U1053 (N_1053,N_894,N_844);
nand U1054 (N_1054,N_830,N_825);
nor U1055 (N_1055,N_806,N_843);
nand U1056 (N_1056,N_877,N_872);
nand U1057 (N_1057,N_978,N_907);
nand U1058 (N_1058,N_822,N_992);
nor U1059 (N_1059,N_807,N_873);
or U1060 (N_1060,N_986,N_960);
xnor U1061 (N_1061,N_818,N_816);
and U1062 (N_1062,N_914,N_936);
and U1063 (N_1063,N_915,N_858);
nand U1064 (N_1064,N_967,N_912);
nor U1065 (N_1065,N_876,N_933);
and U1066 (N_1066,N_803,N_828);
nor U1067 (N_1067,N_884,N_856);
or U1068 (N_1068,N_976,N_971);
nor U1069 (N_1069,N_940,N_853);
and U1070 (N_1070,N_938,N_969);
nor U1071 (N_1071,N_893,N_924);
and U1072 (N_1072,N_849,N_931);
and U1073 (N_1073,N_973,N_906);
nor U1074 (N_1074,N_994,N_908);
nor U1075 (N_1075,N_903,N_988);
xor U1076 (N_1076,N_953,N_855);
or U1077 (N_1077,N_935,N_815);
nand U1078 (N_1078,N_964,N_925);
and U1079 (N_1079,N_859,N_846);
or U1080 (N_1080,N_824,N_961);
and U1081 (N_1081,N_881,N_819);
nor U1082 (N_1082,N_812,N_850);
nor U1083 (N_1083,N_808,N_980);
and U1084 (N_1084,N_958,N_875);
nor U1085 (N_1085,N_829,N_991);
and U1086 (N_1086,N_880,N_890);
nand U1087 (N_1087,N_909,N_981);
or U1088 (N_1088,N_959,N_984);
or U1089 (N_1089,N_811,N_985);
and U1090 (N_1090,N_989,N_928);
nor U1091 (N_1091,N_866,N_999);
xnor U1092 (N_1092,N_951,N_996);
nand U1093 (N_1093,N_809,N_887);
and U1094 (N_1094,N_922,N_889);
nand U1095 (N_1095,N_861,N_867);
and U1096 (N_1096,N_949,N_945);
nor U1097 (N_1097,N_902,N_896);
nor U1098 (N_1098,N_814,N_905);
and U1099 (N_1099,N_883,N_977);
nand U1100 (N_1100,N_996,N_862);
nand U1101 (N_1101,N_806,N_833);
nand U1102 (N_1102,N_909,N_921);
nand U1103 (N_1103,N_834,N_830);
nor U1104 (N_1104,N_899,N_874);
and U1105 (N_1105,N_914,N_851);
or U1106 (N_1106,N_816,N_939);
nand U1107 (N_1107,N_985,N_897);
nand U1108 (N_1108,N_861,N_975);
or U1109 (N_1109,N_959,N_944);
and U1110 (N_1110,N_902,N_805);
nand U1111 (N_1111,N_995,N_843);
and U1112 (N_1112,N_877,N_911);
or U1113 (N_1113,N_895,N_954);
or U1114 (N_1114,N_907,N_948);
and U1115 (N_1115,N_991,N_896);
or U1116 (N_1116,N_881,N_957);
nor U1117 (N_1117,N_828,N_862);
nand U1118 (N_1118,N_910,N_853);
nand U1119 (N_1119,N_850,N_967);
and U1120 (N_1120,N_839,N_843);
or U1121 (N_1121,N_875,N_897);
nor U1122 (N_1122,N_940,N_875);
or U1123 (N_1123,N_835,N_802);
or U1124 (N_1124,N_880,N_963);
xor U1125 (N_1125,N_856,N_876);
nand U1126 (N_1126,N_999,N_933);
or U1127 (N_1127,N_896,N_931);
nand U1128 (N_1128,N_951,N_962);
nand U1129 (N_1129,N_991,N_927);
nand U1130 (N_1130,N_948,N_802);
and U1131 (N_1131,N_924,N_844);
nor U1132 (N_1132,N_884,N_971);
and U1133 (N_1133,N_868,N_949);
or U1134 (N_1134,N_970,N_883);
and U1135 (N_1135,N_939,N_884);
nand U1136 (N_1136,N_827,N_936);
nand U1137 (N_1137,N_865,N_833);
nand U1138 (N_1138,N_959,N_840);
or U1139 (N_1139,N_973,N_916);
and U1140 (N_1140,N_807,N_932);
nand U1141 (N_1141,N_837,N_898);
xor U1142 (N_1142,N_869,N_807);
nor U1143 (N_1143,N_991,N_992);
nor U1144 (N_1144,N_872,N_948);
and U1145 (N_1145,N_956,N_873);
or U1146 (N_1146,N_826,N_808);
and U1147 (N_1147,N_948,N_951);
and U1148 (N_1148,N_932,N_853);
or U1149 (N_1149,N_981,N_846);
nand U1150 (N_1150,N_865,N_979);
and U1151 (N_1151,N_978,N_976);
and U1152 (N_1152,N_957,N_853);
or U1153 (N_1153,N_882,N_948);
and U1154 (N_1154,N_855,N_963);
nand U1155 (N_1155,N_993,N_874);
xnor U1156 (N_1156,N_939,N_921);
and U1157 (N_1157,N_971,N_982);
and U1158 (N_1158,N_911,N_845);
and U1159 (N_1159,N_998,N_904);
or U1160 (N_1160,N_937,N_865);
nand U1161 (N_1161,N_829,N_913);
and U1162 (N_1162,N_900,N_817);
xnor U1163 (N_1163,N_948,N_878);
or U1164 (N_1164,N_823,N_926);
and U1165 (N_1165,N_865,N_919);
nor U1166 (N_1166,N_983,N_803);
and U1167 (N_1167,N_973,N_850);
or U1168 (N_1168,N_872,N_964);
or U1169 (N_1169,N_820,N_951);
and U1170 (N_1170,N_870,N_939);
nor U1171 (N_1171,N_806,N_860);
or U1172 (N_1172,N_821,N_954);
nand U1173 (N_1173,N_907,N_818);
nand U1174 (N_1174,N_973,N_921);
or U1175 (N_1175,N_937,N_877);
nand U1176 (N_1176,N_980,N_959);
nor U1177 (N_1177,N_932,N_934);
xor U1178 (N_1178,N_855,N_964);
and U1179 (N_1179,N_994,N_921);
and U1180 (N_1180,N_801,N_909);
nand U1181 (N_1181,N_902,N_837);
nor U1182 (N_1182,N_872,N_972);
nor U1183 (N_1183,N_921,N_854);
nand U1184 (N_1184,N_818,N_951);
and U1185 (N_1185,N_939,N_989);
nor U1186 (N_1186,N_866,N_987);
nor U1187 (N_1187,N_897,N_986);
nand U1188 (N_1188,N_912,N_936);
and U1189 (N_1189,N_951,N_805);
nor U1190 (N_1190,N_819,N_824);
or U1191 (N_1191,N_975,N_912);
or U1192 (N_1192,N_844,N_987);
nor U1193 (N_1193,N_832,N_844);
and U1194 (N_1194,N_874,N_836);
or U1195 (N_1195,N_855,N_933);
and U1196 (N_1196,N_968,N_834);
nor U1197 (N_1197,N_850,N_854);
nand U1198 (N_1198,N_932,N_889);
or U1199 (N_1199,N_973,N_901);
nand U1200 (N_1200,N_1168,N_1042);
and U1201 (N_1201,N_1022,N_1175);
or U1202 (N_1202,N_1186,N_1161);
and U1203 (N_1203,N_1153,N_1148);
nand U1204 (N_1204,N_1061,N_1034);
or U1205 (N_1205,N_1129,N_1033);
nor U1206 (N_1206,N_1071,N_1036);
and U1207 (N_1207,N_1182,N_1086);
nand U1208 (N_1208,N_1039,N_1140);
and U1209 (N_1209,N_1013,N_1045);
nor U1210 (N_1210,N_1193,N_1081);
and U1211 (N_1211,N_1038,N_1110);
nor U1212 (N_1212,N_1128,N_1195);
nor U1213 (N_1213,N_1112,N_1184);
xor U1214 (N_1214,N_1047,N_1088);
xnor U1215 (N_1215,N_1080,N_1040);
nand U1216 (N_1216,N_1165,N_1017);
nand U1217 (N_1217,N_1111,N_1123);
nand U1218 (N_1218,N_1062,N_1104);
nand U1219 (N_1219,N_1027,N_1023);
or U1220 (N_1220,N_1196,N_1149);
and U1221 (N_1221,N_1041,N_1199);
or U1222 (N_1222,N_1142,N_1152);
nand U1223 (N_1223,N_1019,N_1162);
and U1224 (N_1224,N_1091,N_1114);
or U1225 (N_1225,N_1026,N_1069);
and U1226 (N_1226,N_1093,N_1085);
or U1227 (N_1227,N_1126,N_1057);
nor U1228 (N_1228,N_1049,N_1108);
nor U1229 (N_1229,N_1191,N_1054);
nor U1230 (N_1230,N_1089,N_1079);
xor U1231 (N_1231,N_1192,N_1117);
nand U1232 (N_1232,N_1084,N_1058);
nor U1233 (N_1233,N_1167,N_1095);
nor U1234 (N_1234,N_1075,N_1147);
or U1235 (N_1235,N_1030,N_1092);
or U1236 (N_1236,N_1124,N_1083);
and U1237 (N_1237,N_1109,N_1094);
and U1238 (N_1238,N_1107,N_1014);
nand U1239 (N_1239,N_1125,N_1174);
or U1240 (N_1240,N_1187,N_1063);
and U1241 (N_1241,N_1068,N_1133);
nor U1242 (N_1242,N_1181,N_1105);
nor U1243 (N_1243,N_1053,N_1159);
nand U1244 (N_1244,N_1066,N_1177);
nor U1245 (N_1245,N_1031,N_1003);
nor U1246 (N_1246,N_1012,N_1180);
or U1247 (N_1247,N_1096,N_1144);
or U1248 (N_1248,N_1119,N_1158);
or U1249 (N_1249,N_1064,N_1029);
or U1250 (N_1250,N_1115,N_1001);
or U1251 (N_1251,N_1130,N_1150);
and U1252 (N_1252,N_1028,N_1009);
nor U1253 (N_1253,N_1032,N_1122);
xor U1254 (N_1254,N_1078,N_1157);
or U1255 (N_1255,N_1137,N_1116);
and U1256 (N_1256,N_1076,N_1050);
nand U1257 (N_1257,N_1018,N_1008);
and U1258 (N_1258,N_1006,N_1141);
and U1259 (N_1259,N_1102,N_1067);
xnor U1260 (N_1260,N_1021,N_1059);
nor U1261 (N_1261,N_1048,N_1188);
or U1262 (N_1262,N_1198,N_1143);
nor U1263 (N_1263,N_1035,N_1185);
nand U1264 (N_1264,N_1051,N_1146);
and U1265 (N_1265,N_1024,N_1160);
and U1266 (N_1266,N_1015,N_1169);
or U1267 (N_1267,N_1100,N_1052);
nor U1268 (N_1268,N_1055,N_1189);
or U1269 (N_1269,N_1010,N_1135);
and U1270 (N_1270,N_1127,N_1139);
nor U1271 (N_1271,N_1000,N_1002);
nor U1272 (N_1272,N_1007,N_1164);
nand U1273 (N_1273,N_1090,N_1172);
and U1274 (N_1274,N_1082,N_1178);
nor U1275 (N_1275,N_1087,N_1155);
and U1276 (N_1276,N_1005,N_1043);
nand U1277 (N_1277,N_1136,N_1132);
and U1278 (N_1278,N_1197,N_1138);
or U1279 (N_1279,N_1037,N_1170);
or U1280 (N_1280,N_1103,N_1163);
nand U1281 (N_1281,N_1118,N_1176);
and U1282 (N_1282,N_1156,N_1065);
nor U1283 (N_1283,N_1131,N_1070);
nor U1284 (N_1284,N_1044,N_1166);
nor U1285 (N_1285,N_1074,N_1120);
nand U1286 (N_1286,N_1020,N_1025);
or U1287 (N_1287,N_1179,N_1099);
or U1288 (N_1288,N_1171,N_1154);
or U1289 (N_1289,N_1097,N_1113);
or U1290 (N_1290,N_1183,N_1151);
and U1291 (N_1291,N_1190,N_1073);
and U1292 (N_1292,N_1173,N_1121);
or U1293 (N_1293,N_1060,N_1098);
or U1294 (N_1294,N_1101,N_1011);
nor U1295 (N_1295,N_1016,N_1046);
or U1296 (N_1296,N_1056,N_1145);
nand U1297 (N_1297,N_1194,N_1106);
nor U1298 (N_1298,N_1072,N_1077);
and U1299 (N_1299,N_1134,N_1004);
nor U1300 (N_1300,N_1018,N_1056);
nand U1301 (N_1301,N_1156,N_1141);
nand U1302 (N_1302,N_1054,N_1031);
nand U1303 (N_1303,N_1116,N_1028);
nand U1304 (N_1304,N_1090,N_1007);
nand U1305 (N_1305,N_1192,N_1163);
xnor U1306 (N_1306,N_1097,N_1178);
or U1307 (N_1307,N_1031,N_1189);
and U1308 (N_1308,N_1068,N_1153);
and U1309 (N_1309,N_1162,N_1058);
nor U1310 (N_1310,N_1044,N_1058);
nand U1311 (N_1311,N_1116,N_1063);
nand U1312 (N_1312,N_1145,N_1140);
nor U1313 (N_1313,N_1023,N_1126);
nand U1314 (N_1314,N_1063,N_1120);
and U1315 (N_1315,N_1191,N_1126);
nand U1316 (N_1316,N_1085,N_1167);
and U1317 (N_1317,N_1006,N_1115);
or U1318 (N_1318,N_1151,N_1191);
and U1319 (N_1319,N_1034,N_1148);
and U1320 (N_1320,N_1007,N_1072);
nor U1321 (N_1321,N_1080,N_1134);
nor U1322 (N_1322,N_1052,N_1132);
nor U1323 (N_1323,N_1049,N_1064);
or U1324 (N_1324,N_1010,N_1190);
or U1325 (N_1325,N_1185,N_1123);
nand U1326 (N_1326,N_1112,N_1072);
nor U1327 (N_1327,N_1142,N_1053);
or U1328 (N_1328,N_1024,N_1138);
or U1329 (N_1329,N_1080,N_1181);
or U1330 (N_1330,N_1143,N_1032);
or U1331 (N_1331,N_1090,N_1196);
and U1332 (N_1332,N_1131,N_1097);
nor U1333 (N_1333,N_1191,N_1063);
and U1334 (N_1334,N_1023,N_1145);
nor U1335 (N_1335,N_1128,N_1098);
or U1336 (N_1336,N_1177,N_1046);
nand U1337 (N_1337,N_1120,N_1183);
nand U1338 (N_1338,N_1035,N_1080);
and U1339 (N_1339,N_1015,N_1179);
nand U1340 (N_1340,N_1060,N_1150);
xnor U1341 (N_1341,N_1082,N_1021);
or U1342 (N_1342,N_1106,N_1111);
nand U1343 (N_1343,N_1093,N_1169);
or U1344 (N_1344,N_1101,N_1111);
nand U1345 (N_1345,N_1076,N_1031);
nor U1346 (N_1346,N_1060,N_1114);
or U1347 (N_1347,N_1033,N_1041);
nand U1348 (N_1348,N_1031,N_1049);
or U1349 (N_1349,N_1002,N_1117);
and U1350 (N_1350,N_1066,N_1055);
nor U1351 (N_1351,N_1088,N_1160);
or U1352 (N_1352,N_1102,N_1029);
nor U1353 (N_1353,N_1114,N_1038);
and U1354 (N_1354,N_1133,N_1120);
nand U1355 (N_1355,N_1032,N_1006);
nand U1356 (N_1356,N_1054,N_1123);
nand U1357 (N_1357,N_1068,N_1061);
and U1358 (N_1358,N_1058,N_1086);
or U1359 (N_1359,N_1115,N_1039);
or U1360 (N_1360,N_1184,N_1175);
and U1361 (N_1361,N_1143,N_1145);
nor U1362 (N_1362,N_1194,N_1186);
or U1363 (N_1363,N_1139,N_1016);
nand U1364 (N_1364,N_1026,N_1194);
and U1365 (N_1365,N_1040,N_1162);
and U1366 (N_1366,N_1021,N_1176);
nand U1367 (N_1367,N_1120,N_1118);
nor U1368 (N_1368,N_1124,N_1161);
nor U1369 (N_1369,N_1005,N_1087);
and U1370 (N_1370,N_1001,N_1103);
and U1371 (N_1371,N_1092,N_1017);
nand U1372 (N_1372,N_1014,N_1096);
and U1373 (N_1373,N_1056,N_1092);
and U1374 (N_1374,N_1064,N_1066);
and U1375 (N_1375,N_1017,N_1005);
nor U1376 (N_1376,N_1171,N_1186);
and U1377 (N_1377,N_1119,N_1099);
or U1378 (N_1378,N_1129,N_1031);
and U1379 (N_1379,N_1020,N_1002);
nor U1380 (N_1380,N_1067,N_1179);
nand U1381 (N_1381,N_1046,N_1182);
nand U1382 (N_1382,N_1086,N_1018);
nor U1383 (N_1383,N_1064,N_1095);
nor U1384 (N_1384,N_1104,N_1167);
or U1385 (N_1385,N_1094,N_1026);
or U1386 (N_1386,N_1008,N_1118);
nand U1387 (N_1387,N_1068,N_1108);
or U1388 (N_1388,N_1021,N_1143);
and U1389 (N_1389,N_1081,N_1031);
or U1390 (N_1390,N_1188,N_1028);
nand U1391 (N_1391,N_1075,N_1196);
and U1392 (N_1392,N_1114,N_1155);
nor U1393 (N_1393,N_1010,N_1179);
nor U1394 (N_1394,N_1001,N_1105);
and U1395 (N_1395,N_1043,N_1074);
or U1396 (N_1396,N_1105,N_1008);
nand U1397 (N_1397,N_1154,N_1079);
nor U1398 (N_1398,N_1106,N_1066);
nor U1399 (N_1399,N_1154,N_1175);
nand U1400 (N_1400,N_1291,N_1357);
or U1401 (N_1401,N_1277,N_1319);
nand U1402 (N_1402,N_1379,N_1265);
or U1403 (N_1403,N_1311,N_1245);
nand U1404 (N_1404,N_1275,N_1316);
and U1405 (N_1405,N_1307,N_1303);
or U1406 (N_1406,N_1358,N_1312);
nor U1407 (N_1407,N_1289,N_1306);
or U1408 (N_1408,N_1239,N_1323);
or U1409 (N_1409,N_1349,N_1278);
and U1410 (N_1410,N_1346,N_1288);
or U1411 (N_1411,N_1330,N_1264);
or U1412 (N_1412,N_1372,N_1226);
nand U1413 (N_1413,N_1284,N_1356);
nand U1414 (N_1414,N_1370,N_1282);
nor U1415 (N_1415,N_1293,N_1329);
and U1416 (N_1416,N_1242,N_1213);
nor U1417 (N_1417,N_1220,N_1224);
xnor U1418 (N_1418,N_1261,N_1201);
and U1419 (N_1419,N_1233,N_1260);
nand U1420 (N_1420,N_1371,N_1396);
or U1421 (N_1421,N_1361,N_1309);
or U1422 (N_1422,N_1366,N_1318);
or U1423 (N_1423,N_1281,N_1297);
nor U1424 (N_1424,N_1292,N_1302);
and U1425 (N_1425,N_1285,N_1287);
nor U1426 (N_1426,N_1283,N_1328);
and U1427 (N_1427,N_1204,N_1249);
and U1428 (N_1428,N_1397,N_1270);
or U1429 (N_1429,N_1359,N_1387);
or U1430 (N_1430,N_1335,N_1229);
nor U1431 (N_1431,N_1376,N_1207);
nor U1432 (N_1432,N_1389,N_1324);
or U1433 (N_1433,N_1232,N_1365);
nor U1434 (N_1434,N_1255,N_1295);
nand U1435 (N_1435,N_1258,N_1344);
and U1436 (N_1436,N_1217,N_1345);
or U1437 (N_1437,N_1222,N_1206);
or U1438 (N_1438,N_1325,N_1313);
nand U1439 (N_1439,N_1314,N_1263);
and U1440 (N_1440,N_1210,N_1266);
xnor U1441 (N_1441,N_1205,N_1342);
and U1442 (N_1442,N_1360,N_1398);
nor U1443 (N_1443,N_1305,N_1355);
and U1444 (N_1444,N_1271,N_1351);
nand U1445 (N_1445,N_1272,N_1280);
and U1446 (N_1446,N_1269,N_1251);
and U1447 (N_1447,N_1394,N_1273);
or U1448 (N_1448,N_1214,N_1254);
or U1449 (N_1449,N_1378,N_1338);
or U1450 (N_1450,N_1363,N_1294);
nand U1451 (N_1451,N_1375,N_1352);
nand U1452 (N_1452,N_1274,N_1267);
and U1453 (N_1453,N_1384,N_1334);
nand U1454 (N_1454,N_1348,N_1276);
xnor U1455 (N_1455,N_1399,N_1320);
nand U1456 (N_1456,N_1364,N_1225);
nand U1457 (N_1457,N_1317,N_1230);
or U1458 (N_1458,N_1347,N_1354);
nand U1459 (N_1459,N_1315,N_1202);
nand U1460 (N_1460,N_1308,N_1337);
nor U1461 (N_1461,N_1259,N_1333);
nor U1462 (N_1462,N_1322,N_1250);
or U1463 (N_1463,N_1368,N_1331);
xnor U1464 (N_1464,N_1253,N_1310);
nand U1465 (N_1465,N_1301,N_1290);
nor U1466 (N_1466,N_1248,N_1246);
or U1467 (N_1467,N_1223,N_1390);
nor U1468 (N_1468,N_1383,N_1208);
nor U1469 (N_1469,N_1388,N_1238);
nand U1470 (N_1470,N_1200,N_1286);
nand U1471 (N_1471,N_1227,N_1377);
or U1472 (N_1472,N_1367,N_1216);
nor U1473 (N_1473,N_1326,N_1211);
nor U1474 (N_1474,N_1252,N_1257);
nor U1475 (N_1475,N_1296,N_1298);
and U1476 (N_1476,N_1236,N_1393);
nor U1477 (N_1477,N_1374,N_1234);
or U1478 (N_1478,N_1237,N_1300);
and U1479 (N_1479,N_1268,N_1304);
nand U1480 (N_1480,N_1262,N_1341);
and U1481 (N_1481,N_1299,N_1340);
or U1482 (N_1482,N_1256,N_1332);
nor U1483 (N_1483,N_1391,N_1279);
and U1484 (N_1484,N_1221,N_1395);
nand U1485 (N_1485,N_1362,N_1219);
nand U1486 (N_1486,N_1209,N_1392);
and U1487 (N_1487,N_1369,N_1240);
nand U1488 (N_1488,N_1235,N_1382);
and U1489 (N_1489,N_1386,N_1231);
or U1490 (N_1490,N_1228,N_1212);
nor U1491 (N_1491,N_1385,N_1343);
nand U1492 (N_1492,N_1241,N_1203);
and U1493 (N_1493,N_1373,N_1243);
nor U1494 (N_1494,N_1336,N_1244);
and U1495 (N_1495,N_1327,N_1247);
or U1496 (N_1496,N_1380,N_1321);
and U1497 (N_1497,N_1218,N_1215);
nor U1498 (N_1498,N_1381,N_1339);
nand U1499 (N_1499,N_1350,N_1353);
and U1500 (N_1500,N_1299,N_1232);
nand U1501 (N_1501,N_1278,N_1335);
and U1502 (N_1502,N_1269,N_1209);
or U1503 (N_1503,N_1339,N_1357);
nor U1504 (N_1504,N_1230,N_1365);
or U1505 (N_1505,N_1230,N_1369);
nor U1506 (N_1506,N_1348,N_1375);
or U1507 (N_1507,N_1232,N_1352);
and U1508 (N_1508,N_1289,N_1347);
nor U1509 (N_1509,N_1380,N_1290);
and U1510 (N_1510,N_1283,N_1373);
nor U1511 (N_1511,N_1287,N_1388);
nor U1512 (N_1512,N_1265,N_1388);
or U1513 (N_1513,N_1231,N_1311);
nor U1514 (N_1514,N_1331,N_1261);
or U1515 (N_1515,N_1340,N_1266);
nand U1516 (N_1516,N_1255,N_1329);
nand U1517 (N_1517,N_1307,N_1262);
nor U1518 (N_1518,N_1269,N_1211);
or U1519 (N_1519,N_1353,N_1392);
nor U1520 (N_1520,N_1227,N_1273);
nor U1521 (N_1521,N_1264,N_1328);
nand U1522 (N_1522,N_1355,N_1363);
xnor U1523 (N_1523,N_1213,N_1234);
nand U1524 (N_1524,N_1326,N_1320);
nor U1525 (N_1525,N_1327,N_1365);
nor U1526 (N_1526,N_1397,N_1277);
nand U1527 (N_1527,N_1369,N_1394);
or U1528 (N_1528,N_1274,N_1227);
nor U1529 (N_1529,N_1266,N_1215);
xor U1530 (N_1530,N_1360,N_1283);
nand U1531 (N_1531,N_1386,N_1294);
and U1532 (N_1532,N_1335,N_1208);
nand U1533 (N_1533,N_1221,N_1255);
nand U1534 (N_1534,N_1220,N_1375);
or U1535 (N_1535,N_1214,N_1289);
nand U1536 (N_1536,N_1272,N_1278);
nor U1537 (N_1537,N_1262,N_1223);
or U1538 (N_1538,N_1368,N_1395);
and U1539 (N_1539,N_1295,N_1357);
nor U1540 (N_1540,N_1261,N_1369);
or U1541 (N_1541,N_1225,N_1283);
nand U1542 (N_1542,N_1303,N_1372);
or U1543 (N_1543,N_1305,N_1384);
and U1544 (N_1544,N_1259,N_1350);
nor U1545 (N_1545,N_1248,N_1231);
nor U1546 (N_1546,N_1353,N_1279);
or U1547 (N_1547,N_1364,N_1294);
nor U1548 (N_1548,N_1210,N_1213);
nand U1549 (N_1549,N_1353,N_1352);
or U1550 (N_1550,N_1391,N_1300);
nand U1551 (N_1551,N_1320,N_1219);
and U1552 (N_1552,N_1265,N_1397);
and U1553 (N_1553,N_1354,N_1350);
nand U1554 (N_1554,N_1207,N_1315);
nand U1555 (N_1555,N_1298,N_1293);
or U1556 (N_1556,N_1365,N_1253);
and U1557 (N_1557,N_1391,N_1267);
nand U1558 (N_1558,N_1290,N_1345);
nor U1559 (N_1559,N_1227,N_1277);
nand U1560 (N_1560,N_1399,N_1270);
nor U1561 (N_1561,N_1382,N_1219);
nand U1562 (N_1562,N_1319,N_1326);
or U1563 (N_1563,N_1397,N_1286);
nand U1564 (N_1564,N_1205,N_1349);
or U1565 (N_1565,N_1233,N_1267);
nor U1566 (N_1566,N_1284,N_1285);
and U1567 (N_1567,N_1322,N_1309);
nand U1568 (N_1568,N_1369,N_1347);
and U1569 (N_1569,N_1235,N_1393);
nand U1570 (N_1570,N_1347,N_1330);
or U1571 (N_1571,N_1366,N_1305);
and U1572 (N_1572,N_1358,N_1224);
xor U1573 (N_1573,N_1301,N_1355);
and U1574 (N_1574,N_1254,N_1244);
nor U1575 (N_1575,N_1364,N_1388);
nor U1576 (N_1576,N_1289,N_1354);
nor U1577 (N_1577,N_1388,N_1322);
nand U1578 (N_1578,N_1352,N_1237);
and U1579 (N_1579,N_1323,N_1217);
or U1580 (N_1580,N_1209,N_1247);
nand U1581 (N_1581,N_1376,N_1380);
nand U1582 (N_1582,N_1259,N_1263);
or U1583 (N_1583,N_1348,N_1236);
and U1584 (N_1584,N_1320,N_1247);
or U1585 (N_1585,N_1237,N_1319);
or U1586 (N_1586,N_1292,N_1284);
nor U1587 (N_1587,N_1388,N_1230);
nor U1588 (N_1588,N_1294,N_1322);
nand U1589 (N_1589,N_1357,N_1276);
nand U1590 (N_1590,N_1391,N_1381);
or U1591 (N_1591,N_1384,N_1306);
or U1592 (N_1592,N_1371,N_1389);
and U1593 (N_1593,N_1302,N_1255);
nor U1594 (N_1594,N_1336,N_1353);
and U1595 (N_1595,N_1313,N_1314);
nor U1596 (N_1596,N_1324,N_1260);
and U1597 (N_1597,N_1216,N_1206);
or U1598 (N_1598,N_1360,N_1368);
nand U1599 (N_1599,N_1296,N_1284);
nor U1600 (N_1600,N_1592,N_1436);
or U1601 (N_1601,N_1596,N_1482);
nor U1602 (N_1602,N_1548,N_1559);
nand U1603 (N_1603,N_1506,N_1431);
nand U1604 (N_1604,N_1529,N_1423);
nand U1605 (N_1605,N_1453,N_1552);
nor U1606 (N_1606,N_1459,N_1472);
or U1607 (N_1607,N_1427,N_1512);
and U1608 (N_1608,N_1510,N_1590);
or U1609 (N_1609,N_1542,N_1434);
nor U1610 (N_1610,N_1464,N_1477);
nor U1611 (N_1611,N_1583,N_1538);
nor U1612 (N_1612,N_1569,N_1415);
or U1613 (N_1613,N_1425,N_1483);
and U1614 (N_1614,N_1413,N_1401);
nand U1615 (N_1615,N_1406,N_1561);
or U1616 (N_1616,N_1437,N_1543);
nor U1617 (N_1617,N_1519,N_1547);
nand U1618 (N_1618,N_1443,N_1549);
nor U1619 (N_1619,N_1585,N_1424);
nand U1620 (N_1620,N_1422,N_1435);
xnor U1621 (N_1621,N_1518,N_1479);
nand U1622 (N_1622,N_1446,N_1591);
nor U1623 (N_1623,N_1462,N_1491);
nand U1624 (N_1624,N_1553,N_1454);
and U1625 (N_1625,N_1579,N_1540);
nand U1626 (N_1626,N_1456,N_1545);
nor U1627 (N_1627,N_1408,N_1452);
or U1628 (N_1628,N_1485,N_1532);
nor U1629 (N_1629,N_1572,N_1449);
nor U1630 (N_1630,N_1516,N_1567);
and U1631 (N_1631,N_1587,N_1495);
and U1632 (N_1632,N_1418,N_1576);
nand U1633 (N_1633,N_1439,N_1457);
or U1634 (N_1634,N_1588,N_1577);
and U1635 (N_1635,N_1544,N_1410);
or U1636 (N_1636,N_1531,N_1499);
and U1637 (N_1637,N_1503,N_1556);
or U1638 (N_1638,N_1411,N_1507);
and U1639 (N_1639,N_1550,N_1526);
nand U1640 (N_1640,N_1575,N_1470);
nand U1641 (N_1641,N_1511,N_1541);
and U1642 (N_1642,N_1484,N_1451);
nand U1643 (N_1643,N_1461,N_1586);
nor U1644 (N_1644,N_1487,N_1473);
nor U1645 (N_1645,N_1494,N_1574);
nor U1646 (N_1646,N_1403,N_1471);
nor U1647 (N_1647,N_1476,N_1426);
or U1648 (N_1648,N_1525,N_1417);
and U1649 (N_1649,N_1475,N_1407);
or U1650 (N_1650,N_1489,N_1536);
or U1651 (N_1651,N_1441,N_1509);
nand U1652 (N_1652,N_1496,N_1515);
and U1653 (N_1653,N_1508,N_1402);
nand U1654 (N_1654,N_1492,N_1432);
and U1655 (N_1655,N_1527,N_1584);
nor U1656 (N_1656,N_1563,N_1595);
or U1657 (N_1657,N_1478,N_1420);
nand U1658 (N_1658,N_1551,N_1480);
or U1659 (N_1659,N_1474,N_1593);
nor U1660 (N_1660,N_1488,N_1568);
nor U1661 (N_1661,N_1502,N_1400);
nand U1662 (N_1662,N_1493,N_1497);
and U1663 (N_1663,N_1571,N_1481);
nor U1664 (N_1664,N_1486,N_1524);
and U1665 (N_1665,N_1537,N_1513);
or U1666 (N_1666,N_1465,N_1555);
nor U1667 (N_1667,N_1594,N_1460);
nor U1668 (N_1668,N_1533,N_1501);
and U1669 (N_1669,N_1438,N_1500);
nor U1670 (N_1670,N_1463,N_1554);
or U1671 (N_1671,N_1578,N_1564);
nor U1672 (N_1672,N_1444,N_1409);
nand U1673 (N_1673,N_1430,N_1570);
or U1674 (N_1674,N_1522,N_1404);
and U1675 (N_1675,N_1448,N_1469);
xnor U1676 (N_1676,N_1514,N_1517);
xor U1677 (N_1677,N_1546,N_1530);
nand U1678 (N_1678,N_1428,N_1589);
nand U1679 (N_1679,N_1557,N_1405);
and U1680 (N_1680,N_1520,N_1505);
nor U1681 (N_1681,N_1458,N_1429);
or U1682 (N_1682,N_1534,N_1581);
and U1683 (N_1683,N_1599,N_1504);
and U1684 (N_1684,N_1573,N_1562);
or U1685 (N_1685,N_1566,N_1558);
nor U1686 (N_1686,N_1445,N_1421);
nand U1687 (N_1687,N_1414,N_1467);
nor U1688 (N_1688,N_1433,N_1442);
and U1689 (N_1689,N_1560,N_1597);
nand U1690 (N_1690,N_1582,N_1447);
or U1691 (N_1691,N_1539,N_1468);
nor U1692 (N_1692,N_1565,N_1440);
nor U1693 (N_1693,N_1521,N_1580);
and U1694 (N_1694,N_1523,N_1455);
and U1695 (N_1695,N_1450,N_1412);
nor U1696 (N_1696,N_1498,N_1535);
nor U1697 (N_1697,N_1466,N_1528);
nand U1698 (N_1698,N_1598,N_1419);
and U1699 (N_1699,N_1416,N_1490);
nor U1700 (N_1700,N_1513,N_1526);
or U1701 (N_1701,N_1504,N_1595);
nand U1702 (N_1702,N_1593,N_1540);
nand U1703 (N_1703,N_1428,N_1579);
nor U1704 (N_1704,N_1599,N_1545);
nor U1705 (N_1705,N_1492,N_1449);
nor U1706 (N_1706,N_1456,N_1491);
or U1707 (N_1707,N_1440,N_1519);
and U1708 (N_1708,N_1500,N_1577);
or U1709 (N_1709,N_1540,N_1556);
and U1710 (N_1710,N_1599,N_1429);
and U1711 (N_1711,N_1451,N_1550);
nand U1712 (N_1712,N_1500,N_1564);
or U1713 (N_1713,N_1423,N_1594);
or U1714 (N_1714,N_1591,N_1417);
nand U1715 (N_1715,N_1508,N_1510);
nand U1716 (N_1716,N_1580,N_1599);
or U1717 (N_1717,N_1540,N_1468);
or U1718 (N_1718,N_1565,N_1538);
and U1719 (N_1719,N_1410,N_1576);
and U1720 (N_1720,N_1564,N_1475);
nand U1721 (N_1721,N_1424,N_1474);
nor U1722 (N_1722,N_1554,N_1426);
xor U1723 (N_1723,N_1470,N_1558);
xor U1724 (N_1724,N_1480,N_1594);
nor U1725 (N_1725,N_1539,N_1442);
xnor U1726 (N_1726,N_1512,N_1565);
nor U1727 (N_1727,N_1528,N_1546);
and U1728 (N_1728,N_1412,N_1495);
nand U1729 (N_1729,N_1548,N_1462);
nand U1730 (N_1730,N_1440,N_1485);
nor U1731 (N_1731,N_1538,N_1539);
or U1732 (N_1732,N_1599,N_1400);
and U1733 (N_1733,N_1514,N_1478);
nor U1734 (N_1734,N_1542,N_1598);
nand U1735 (N_1735,N_1403,N_1470);
or U1736 (N_1736,N_1481,N_1519);
nand U1737 (N_1737,N_1567,N_1433);
nand U1738 (N_1738,N_1486,N_1538);
nor U1739 (N_1739,N_1443,N_1417);
and U1740 (N_1740,N_1434,N_1510);
and U1741 (N_1741,N_1540,N_1542);
and U1742 (N_1742,N_1581,N_1491);
and U1743 (N_1743,N_1508,N_1509);
or U1744 (N_1744,N_1525,N_1534);
and U1745 (N_1745,N_1492,N_1575);
nor U1746 (N_1746,N_1583,N_1422);
nor U1747 (N_1747,N_1550,N_1529);
nor U1748 (N_1748,N_1458,N_1455);
nand U1749 (N_1749,N_1416,N_1468);
nand U1750 (N_1750,N_1542,N_1413);
nand U1751 (N_1751,N_1483,N_1410);
nand U1752 (N_1752,N_1532,N_1455);
nand U1753 (N_1753,N_1546,N_1591);
or U1754 (N_1754,N_1548,N_1524);
nand U1755 (N_1755,N_1431,N_1532);
nand U1756 (N_1756,N_1552,N_1579);
nand U1757 (N_1757,N_1503,N_1427);
and U1758 (N_1758,N_1416,N_1567);
nor U1759 (N_1759,N_1404,N_1519);
or U1760 (N_1760,N_1478,N_1565);
nor U1761 (N_1761,N_1409,N_1501);
or U1762 (N_1762,N_1427,N_1527);
and U1763 (N_1763,N_1596,N_1587);
nand U1764 (N_1764,N_1467,N_1552);
nor U1765 (N_1765,N_1488,N_1422);
xor U1766 (N_1766,N_1551,N_1514);
nor U1767 (N_1767,N_1582,N_1477);
or U1768 (N_1768,N_1574,N_1436);
or U1769 (N_1769,N_1555,N_1545);
nand U1770 (N_1770,N_1515,N_1427);
and U1771 (N_1771,N_1516,N_1596);
nand U1772 (N_1772,N_1413,N_1501);
nor U1773 (N_1773,N_1574,N_1463);
and U1774 (N_1774,N_1508,N_1594);
nor U1775 (N_1775,N_1581,N_1560);
nand U1776 (N_1776,N_1533,N_1410);
and U1777 (N_1777,N_1475,N_1483);
nor U1778 (N_1778,N_1510,N_1571);
nor U1779 (N_1779,N_1539,N_1490);
nor U1780 (N_1780,N_1479,N_1429);
or U1781 (N_1781,N_1597,N_1450);
nor U1782 (N_1782,N_1462,N_1549);
nor U1783 (N_1783,N_1556,N_1537);
or U1784 (N_1784,N_1551,N_1506);
nand U1785 (N_1785,N_1535,N_1423);
nor U1786 (N_1786,N_1537,N_1421);
or U1787 (N_1787,N_1481,N_1496);
or U1788 (N_1788,N_1452,N_1592);
or U1789 (N_1789,N_1477,N_1442);
nand U1790 (N_1790,N_1498,N_1540);
or U1791 (N_1791,N_1433,N_1580);
nor U1792 (N_1792,N_1585,N_1572);
nand U1793 (N_1793,N_1489,N_1530);
and U1794 (N_1794,N_1559,N_1589);
or U1795 (N_1795,N_1545,N_1457);
xor U1796 (N_1796,N_1562,N_1548);
or U1797 (N_1797,N_1534,N_1408);
or U1798 (N_1798,N_1434,N_1426);
or U1799 (N_1799,N_1486,N_1418);
nor U1800 (N_1800,N_1761,N_1793);
nand U1801 (N_1801,N_1647,N_1622);
or U1802 (N_1802,N_1774,N_1737);
nor U1803 (N_1803,N_1659,N_1694);
nor U1804 (N_1804,N_1658,N_1777);
or U1805 (N_1805,N_1670,N_1617);
nor U1806 (N_1806,N_1764,N_1619);
nand U1807 (N_1807,N_1615,N_1701);
nor U1808 (N_1808,N_1707,N_1719);
nand U1809 (N_1809,N_1790,N_1778);
nand U1810 (N_1810,N_1709,N_1648);
and U1811 (N_1811,N_1607,N_1728);
nand U1812 (N_1812,N_1725,N_1779);
and U1813 (N_1813,N_1632,N_1634);
or U1814 (N_1814,N_1652,N_1679);
nand U1815 (N_1815,N_1721,N_1757);
nor U1816 (N_1816,N_1646,N_1748);
nor U1817 (N_1817,N_1600,N_1673);
and U1818 (N_1818,N_1769,N_1667);
xor U1819 (N_1819,N_1651,N_1765);
and U1820 (N_1820,N_1669,N_1781);
or U1821 (N_1821,N_1754,N_1794);
nor U1822 (N_1822,N_1636,N_1742);
nor U1823 (N_1823,N_1708,N_1727);
and U1824 (N_1824,N_1678,N_1773);
nand U1825 (N_1825,N_1653,N_1677);
nor U1826 (N_1826,N_1705,N_1642);
nand U1827 (N_1827,N_1620,N_1702);
nand U1828 (N_1828,N_1723,N_1660);
and U1829 (N_1829,N_1602,N_1641);
or U1830 (N_1830,N_1676,N_1629);
or U1831 (N_1831,N_1771,N_1716);
nor U1832 (N_1832,N_1724,N_1776);
nor U1833 (N_1833,N_1656,N_1782);
nor U1834 (N_1834,N_1689,N_1655);
and U1835 (N_1835,N_1681,N_1668);
nor U1836 (N_1836,N_1743,N_1780);
nand U1837 (N_1837,N_1644,N_1758);
or U1838 (N_1838,N_1797,N_1718);
nor U1839 (N_1839,N_1783,N_1795);
and U1840 (N_1840,N_1796,N_1746);
nor U1841 (N_1841,N_1744,N_1755);
or U1842 (N_1842,N_1735,N_1663);
or U1843 (N_1843,N_1700,N_1710);
nor U1844 (N_1844,N_1692,N_1618);
nor U1845 (N_1845,N_1784,N_1661);
nor U1846 (N_1846,N_1760,N_1601);
and U1847 (N_1847,N_1616,N_1604);
and U1848 (N_1848,N_1666,N_1713);
nor U1849 (N_1849,N_1751,N_1635);
or U1850 (N_1850,N_1714,N_1682);
or U1851 (N_1851,N_1739,N_1736);
nand U1852 (N_1852,N_1674,N_1785);
or U1853 (N_1853,N_1726,N_1772);
nor U1854 (N_1854,N_1691,N_1608);
or U1855 (N_1855,N_1638,N_1690);
or U1856 (N_1856,N_1639,N_1624);
nand U1857 (N_1857,N_1697,N_1770);
nor U1858 (N_1858,N_1704,N_1625);
nand U1859 (N_1859,N_1703,N_1627);
or U1860 (N_1860,N_1664,N_1745);
or U1861 (N_1861,N_1603,N_1753);
nor U1862 (N_1862,N_1637,N_1611);
or U1863 (N_1863,N_1741,N_1775);
nand U1864 (N_1864,N_1729,N_1752);
and U1865 (N_1865,N_1633,N_1763);
nand U1866 (N_1866,N_1657,N_1749);
nor U1867 (N_1867,N_1738,N_1799);
nor U1868 (N_1868,N_1649,N_1706);
and U1869 (N_1869,N_1722,N_1747);
or U1870 (N_1870,N_1605,N_1762);
nand U1871 (N_1871,N_1614,N_1683);
or U1872 (N_1872,N_1789,N_1675);
nor U1873 (N_1873,N_1698,N_1766);
nor U1874 (N_1874,N_1643,N_1680);
or U1875 (N_1875,N_1628,N_1613);
and U1876 (N_1876,N_1720,N_1672);
nor U1877 (N_1877,N_1630,N_1750);
or U1878 (N_1878,N_1609,N_1712);
nand U1879 (N_1879,N_1767,N_1786);
and U1880 (N_1880,N_1798,N_1711);
or U1881 (N_1881,N_1693,N_1792);
or U1882 (N_1882,N_1623,N_1671);
or U1883 (N_1883,N_1731,N_1734);
nor U1884 (N_1884,N_1732,N_1759);
nor U1885 (N_1885,N_1631,N_1791);
and U1886 (N_1886,N_1654,N_1699);
nor U1887 (N_1887,N_1650,N_1610);
or U1888 (N_1888,N_1787,N_1740);
nand U1889 (N_1889,N_1626,N_1696);
and U1890 (N_1890,N_1662,N_1715);
nand U1891 (N_1891,N_1768,N_1788);
and U1892 (N_1892,N_1756,N_1717);
and U1893 (N_1893,N_1684,N_1733);
or U1894 (N_1894,N_1730,N_1640);
or U1895 (N_1895,N_1606,N_1687);
or U1896 (N_1896,N_1685,N_1645);
nor U1897 (N_1897,N_1686,N_1665);
xnor U1898 (N_1898,N_1612,N_1695);
and U1899 (N_1899,N_1688,N_1621);
and U1900 (N_1900,N_1782,N_1678);
nand U1901 (N_1901,N_1767,N_1777);
nand U1902 (N_1902,N_1724,N_1773);
or U1903 (N_1903,N_1700,N_1711);
nor U1904 (N_1904,N_1633,N_1645);
and U1905 (N_1905,N_1747,N_1758);
nand U1906 (N_1906,N_1750,N_1682);
nor U1907 (N_1907,N_1784,N_1777);
and U1908 (N_1908,N_1712,N_1690);
nor U1909 (N_1909,N_1622,N_1681);
and U1910 (N_1910,N_1728,N_1799);
nor U1911 (N_1911,N_1780,N_1665);
and U1912 (N_1912,N_1657,N_1778);
nor U1913 (N_1913,N_1748,N_1694);
and U1914 (N_1914,N_1715,N_1655);
nand U1915 (N_1915,N_1641,N_1753);
nor U1916 (N_1916,N_1744,N_1637);
nand U1917 (N_1917,N_1731,N_1709);
nand U1918 (N_1918,N_1793,N_1618);
nor U1919 (N_1919,N_1611,N_1692);
nand U1920 (N_1920,N_1719,N_1657);
nor U1921 (N_1921,N_1634,N_1689);
and U1922 (N_1922,N_1722,N_1751);
and U1923 (N_1923,N_1615,N_1780);
nor U1924 (N_1924,N_1664,N_1640);
nand U1925 (N_1925,N_1773,N_1741);
nand U1926 (N_1926,N_1629,N_1728);
or U1927 (N_1927,N_1776,N_1756);
or U1928 (N_1928,N_1674,N_1726);
and U1929 (N_1929,N_1680,N_1723);
and U1930 (N_1930,N_1740,N_1680);
or U1931 (N_1931,N_1768,N_1795);
nor U1932 (N_1932,N_1616,N_1636);
nand U1933 (N_1933,N_1697,N_1620);
nand U1934 (N_1934,N_1768,N_1652);
and U1935 (N_1935,N_1712,N_1634);
and U1936 (N_1936,N_1652,N_1754);
and U1937 (N_1937,N_1656,N_1617);
or U1938 (N_1938,N_1603,N_1604);
xnor U1939 (N_1939,N_1643,N_1767);
nor U1940 (N_1940,N_1706,N_1790);
nor U1941 (N_1941,N_1621,N_1690);
nand U1942 (N_1942,N_1767,N_1710);
or U1943 (N_1943,N_1741,N_1712);
nor U1944 (N_1944,N_1776,N_1632);
and U1945 (N_1945,N_1691,N_1659);
nor U1946 (N_1946,N_1648,N_1795);
nand U1947 (N_1947,N_1622,N_1760);
nor U1948 (N_1948,N_1656,N_1752);
or U1949 (N_1949,N_1748,N_1675);
nand U1950 (N_1950,N_1612,N_1737);
nand U1951 (N_1951,N_1694,N_1634);
nand U1952 (N_1952,N_1787,N_1736);
nor U1953 (N_1953,N_1797,N_1753);
and U1954 (N_1954,N_1787,N_1673);
nand U1955 (N_1955,N_1796,N_1771);
or U1956 (N_1956,N_1617,N_1611);
nand U1957 (N_1957,N_1742,N_1760);
and U1958 (N_1958,N_1734,N_1770);
and U1959 (N_1959,N_1651,N_1779);
xor U1960 (N_1960,N_1703,N_1717);
or U1961 (N_1961,N_1616,N_1697);
nand U1962 (N_1962,N_1787,N_1705);
or U1963 (N_1963,N_1635,N_1661);
nand U1964 (N_1964,N_1756,N_1758);
or U1965 (N_1965,N_1600,N_1692);
or U1966 (N_1966,N_1791,N_1710);
nand U1967 (N_1967,N_1782,N_1683);
xor U1968 (N_1968,N_1644,N_1664);
and U1969 (N_1969,N_1678,N_1735);
and U1970 (N_1970,N_1606,N_1723);
nand U1971 (N_1971,N_1781,N_1627);
or U1972 (N_1972,N_1793,N_1747);
or U1973 (N_1973,N_1742,N_1715);
nand U1974 (N_1974,N_1684,N_1721);
nor U1975 (N_1975,N_1611,N_1671);
nand U1976 (N_1976,N_1689,N_1760);
nand U1977 (N_1977,N_1659,N_1675);
or U1978 (N_1978,N_1604,N_1618);
nor U1979 (N_1979,N_1777,N_1664);
and U1980 (N_1980,N_1677,N_1615);
and U1981 (N_1981,N_1744,N_1612);
or U1982 (N_1982,N_1786,N_1750);
nand U1983 (N_1983,N_1648,N_1760);
nand U1984 (N_1984,N_1721,N_1620);
nor U1985 (N_1985,N_1744,N_1710);
nor U1986 (N_1986,N_1747,N_1632);
nand U1987 (N_1987,N_1608,N_1674);
or U1988 (N_1988,N_1766,N_1756);
nand U1989 (N_1989,N_1645,N_1763);
or U1990 (N_1990,N_1796,N_1635);
or U1991 (N_1991,N_1772,N_1615);
nand U1992 (N_1992,N_1676,N_1775);
nand U1993 (N_1993,N_1668,N_1648);
nand U1994 (N_1994,N_1651,N_1722);
nor U1995 (N_1995,N_1765,N_1688);
nand U1996 (N_1996,N_1685,N_1600);
or U1997 (N_1997,N_1600,N_1606);
nand U1998 (N_1998,N_1716,N_1601);
nor U1999 (N_1999,N_1652,N_1796);
and U2000 (N_2000,N_1962,N_1940);
nand U2001 (N_2001,N_1934,N_1812);
and U2002 (N_2002,N_1802,N_1897);
nand U2003 (N_2003,N_1807,N_1917);
nor U2004 (N_2004,N_1989,N_1896);
nand U2005 (N_2005,N_1955,N_1904);
nand U2006 (N_2006,N_1863,N_1979);
and U2007 (N_2007,N_1980,N_1957);
nor U2008 (N_2008,N_1935,N_1860);
or U2009 (N_2009,N_1998,N_1872);
nor U2010 (N_2010,N_1987,N_1942);
or U2011 (N_2011,N_1894,N_1887);
nor U2012 (N_2012,N_1965,N_1824);
nor U2013 (N_2013,N_1866,N_1994);
and U2014 (N_2014,N_1950,N_1912);
and U2015 (N_2015,N_1918,N_1846);
nor U2016 (N_2016,N_1902,N_1815);
nor U2017 (N_2017,N_1855,N_1971);
nor U2018 (N_2018,N_1944,N_1837);
nand U2019 (N_2019,N_1926,N_1985);
nor U2020 (N_2020,N_1862,N_1829);
or U2021 (N_2021,N_1927,N_1975);
or U2022 (N_2022,N_1840,N_1868);
nand U2023 (N_2023,N_1891,N_1990);
nor U2024 (N_2024,N_1805,N_1974);
and U2025 (N_2025,N_1895,N_1931);
and U2026 (N_2026,N_1825,N_1937);
nand U2027 (N_2027,N_1910,N_1925);
nand U2028 (N_2028,N_1864,N_1819);
nor U2029 (N_2029,N_1869,N_1905);
nand U2030 (N_2030,N_1839,N_1859);
nand U2031 (N_2031,N_1976,N_1997);
nand U2032 (N_2032,N_1883,N_1876);
or U2033 (N_2033,N_1977,N_1803);
and U2034 (N_2034,N_1958,N_1884);
or U2035 (N_2035,N_1890,N_1875);
nand U2036 (N_2036,N_1936,N_1908);
nor U2037 (N_2037,N_1889,N_1967);
and U2038 (N_2038,N_1809,N_1827);
and U2039 (N_2039,N_1988,N_1814);
and U2040 (N_2040,N_1813,N_1849);
nand U2041 (N_2041,N_1993,N_1892);
nor U2042 (N_2042,N_1885,N_1938);
nor U2043 (N_2043,N_1949,N_1948);
nand U2044 (N_2044,N_1995,N_1960);
nand U2045 (N_2045,N_1870,N_1899);
or U2046 (N_2046,N_1953,N_1847);
nand U2047 (N_2047,N_1867,N_1821);
or U2048 (N_2048,N_1834,N_1920);
nand U2049 (N_2049,N_1991,N_1841);
and U2050 (N_2050,N_1861,N_1945);
nor U2051 (N_2051,N_1930,N_1911);
nor U2052 (N_2052,N_1969,N_1820);
or U2053 (N_2053,N_1959,N_1838);
and U2054 (N_2054,N_1843,N_1941);
and U2055 (N_2055,N_1877,N_1933);
nor U2056 (N_2056,N_1810,N_1832);
nand U2057 (N_2057,N_1924,N_1893);
and U2058 (N_2058,N_1836,N_1857);
nand U2059 (N_2059,N_1811,N_1888);
nor U2060 (N_2060,N_1921,N_1984);
nand U2061 (N_2061,N_1804,N_1986);
nor U2062 (N_2062,N_1886,N_1966);
nand U2063 (N_2063,N_1801,N_1946);
or U2064 (N_2064,N_1844,N_1858);
and U2065 (N_2065,N_1845,N_1800);
nor U2066 (N_2066,N_1928,N_1828);
nand U2067 (N_2067,N_1947,N_1964);
nor U2068 (N_2068,N_1853,N_1956);
nand U2069 (N_2069,N_1831,N_1865);
and U2070 (N_2070,N_1873,N_1981);
xnor U2071 (N_2071,N_1806,N_1880);
and U2072 (N_2072,N_1922,N_1848);
nand U2073 (N_2073,N_1901,N_1919);
or U2074 (N_2074,N_1833,N_1907);
and U2075 (N_2075,N_1854,N_1850);
nor U2076 (N_2076,N_1808,N_1879);
nor U2077 (N_2077,N_1903,N_1932);
nor U2078 (N_2078,N_1943,N_1818);
or U2079 (N_2079,N_1968,N_1999);
and U2080 (N_2080,N_1961,N_1978);
and U2081 (N_2081,N_1826,N_1816);
nor U2082 (N_2082,N_1916,N_1952);
and U2083 (N_2083,N_1856,N_1973);
and U2084 (N_2084,N_1881,N_1996);
and U2085 (N_2085,N_1983,N_1914);
nor U2086 (N_2086,N_1817,N_1822);
and U2087 (N_2087,N_1830,N_1900);
nand U2088 (N_2088,N_1823,N_1913);
and U2089 (N_2089,N_1851,N_1898);
and U2090 (N_2090,N_1842,N_1954);
nand U2091 (N_2091,N_1852,N_1951);
nand U2092 (N_2092,N_1992,N_1871);
nor U2093 (N_2093,N_1970,N_1915);
or U2094 (N_2094,N_1972,N_1982);
nor U2095 (N_2095,N_1906,N_1939);
or U2096 (N_2096,N_1923,N_1963);
and U2097 (N_2097,N_1874,N_1835);
and U2098 (N_2098,N_1929,N_1878);
nand U2099 (N_2099,N_1882,N_1909);
nor U2100 (N_2100,N_1808,N_1849);
and U2101 (N_2101,N_1818,N_1949);
or U2102 (N_2102,N_1844,N_1884);
nor U2103 (N_2103,N_1819,N_1849);
or U2104 (N_2104,N_1937,N_1963);
and U2105 (N_2105,N_1884,N_1998);
nand U2106 (N_2106,N_1968,N_1875);
or U2107 (N_2107,N_1969,N_1959);
and U2108 (N_2108,N_1804,N_1805);
and U2109 (N_2109,N_1856,N_1847);
nand U2110 (N_2110,N_1805,N_1910);
nor U2111 (N_2111,N_1969,N_1972);
nand U2112 (N_2112,N_1925,N_1970);
nor U2113 (N_2113,N_1852,N_1837);
nor U2114 (N_2114,N_1957,N_1908);
and U2115 (N_2115,N_1806,N_1888);
and U2116 (N_2116,N_1947,N_1840);
and U2117 (N_2117,N_1993,N_1809);
nor U2118 (N_2118,N_1983,N_1864);
nand U2119 (N_2119,N_1825,N_1963);
and U2120 (N_2120,N_1962,N_1924);
or U2121 (N_2121,N_1880,N_1836);
and U2122 (N_2122,N_1963,N_1837);
or U2123 (N_2123,N_1861,N_1910);
and U2124 (N_2124,N_1978,N_1911);
nand U2125 (N_2125,N_1966,N_1937);
nand U2126 (N_2126,N_1876,N_1829);
or U2127 (N_2127,N_1898,N_1896);
nand U2128 (N_2128,N_1989,N_1978);
and U2129 (N_2129,N_1801,N_1931);
nor U2130 (N_2130,N_1884,N_1883);
nand U2131 (N_2131,N_1902,N_1908);
or U2132 (N_2132,N_1929,N_1962);
nand U2133 (N_2133,N_1803,N_1844);
and U2134 (N_2134,N_1871,N_1971);
or U2135 (N_2135,N_1874,N_1974);
nor U2136 (N_2136,N_1885,N_1831);
and U2137 (N_2137,N_1835,N_1897);
nor U2138 (N_2138,N_1961,N_1908);
nor U2139 (N_2139,N_1997,N_1800);
and U2140 (N_2140,N_1825,N_1814);
nand U2141 (N_2141,N_1869,N_1916);
nand U2142 (N_2142,N_1983,N_1850);
or U2143 (N_2143,N_1993,N_1808);
nand U2144 (N_2144,N_1824,N_1929);
nor U2145 (N_2145,N_1908,N_1804);
nand U2146 (N_2146,N_1991,N_1921);
nand U2147 (N_2147,N_1860,N_1925);
nand U2148 (N_2148,N_1865,N_1917);
nand U2149 (N_2149,N_1837,N_1814);
nor U2150 (N_2150,N_1947,N_1960);
and U2151 (N_2151,N_1968,N_1834);
nand U2152 (N_2152,N_1956,N_1811);
and U2153 (N_2153,N_1855,N_1951);
or U2154 (N_2154,N_1949,N_1959);
and U2155 (N_2155,N_1861,N_1929);
and U2156 (N_2156,N_1863,N_1889);
nor U2157 (N_2157,N_1859,N_1904);
nand U2158 (N_2158,N_1847,N_1815);
and U2159 (N_2159,N_1995,N_1870);
nand U2160 (N_2160,N_1803,N_1842);
xor U2161 (N_2161,N_1948,N_1811);
or U2162 (N_2162,N_1872,N_1889);
or U2163 (N_2163,N_1961,N_1855);
nand U2164 (N_2164,N_1909,N_1936);
nand U2165 (N_2165,N_1847,N_1930);
and U2166 (N_2166,N_1911,N_1899);
and U2167 (N_2167,N_1977,N_1824);
nand U2168 (N_2168,N_1947,N_1995);
and U2169 (N_2169,N_1888,N_1875);
and U2170 (N_2170,N_1842,N_1911);
or U2171 (N_2171,N_1815,N_1877);
nand U2172 (N_2172,N_1900,N_1996);
nor U2173 (N_2173,N_1867,N_1853);
or U2174 (N_2174,N_1935,N_1939);
xnor U2175 (N_2175,N_1813,N_1966);
or U2176 (N_2176,N_1931,N_1889);
nor U2177 (N_2177,N_1997,N_1973);
nor U2178 (N_2178,N_1968,N_1976);
nand U2179 (N_2179,N_1973,N_1949);
and U2180 (N_2180,N_1908,N_1929);
nor U2181 (N_2181,N_1899,N_1916);
nor U2182 (N_2182,N_1873,N_1980);
and U2183 (N_2183,N_1984,N_1899);
and U2184 (N_2184,N_1820,N_1854);
and U2185 (N_2185,N_1862,N_1894);
or U2186 (N_2186,N_1875,N_1911);
xor U2187 (N_2187,N_1989,N_1813);
or U2188 (N_2188,N_1829,N_1855);
and U2189 (N_2189,N_1912,N_1881);
or U2190 (N_2190,N_1906,N_1901);
nand U2191 (N_2191,N_1954,N_1925);
nand U2192 (N_2192,N_1926,N_1922);
and U2193 (N_2193,N_1980,N_1882);
nor U2194 (N_2194,N_1867,N_1912);
and U2195 (N_2195,N_1805,N_1988);
or U2196 (N_2196,N_1988,N_1957);
and U2197 (N_2197,N_1920,N_1888);
nand U2198 (N_2198,N_1826,N_1987);
nor U2199 (N_2199,N_1931,N_1868);
or U2200 (N_2200,N_2031,N_2158);
nor U2201 (N_2201,N_2192,N_2037);
and U2202 (N_2202,N_2047,N_2036);
or U2203 (N_2203,N_2069,N_2067);
or U2204 (N_2204,N_2176,N_2062);
nand U2205 (N_2205,N_2020,N_2074);
nand U2206 (N_2206,N_2081,N_2018);
nor U2207 (N_2207,N_2131,N_2169);
or U2208 (N_2208,N_2053,N_2121);
and U2209 (N_2209,N_2086,N_2068);
or U2210 (N_2210,N_2174,N_2085);
and U2211 (N_2211,N_2024,N_2122);
nor U2212 (N_2212,N_2083,N_2161);
and U2213 (N_2213,N_2138,N_2061);
and U2214 (N_2214,N_2105,N_2159);
nand U2215 (N_2215,N_2017,N_2019);
and U2216 (N_2216,N_2154,N_2147);
nor U2217 (N_2217,N_2092,N_2189);
and U2218 (N_2218,N_2143,N_2029);
nor U2219 (N_2219,N_2119,N_2065);
nand U2220 (N_2220,N_2127,N_2120);
and U2221 (N_2221,N_2001,N_2040);
nor U2222 (N_2222,N_2155,N_2148);
or U2223 (N_2223,N_2152,N_2052);
and U2224 (N_2224,N_2051,N_2100);
and U2225 (N_2225,N_2116,N_2103);
and U2226 (N_2226,N_2087,N_2175);
or U2227 (N_2227,N_2165,N_2114);
nor U2228 (N_2228,N_2023,N_2091);
and U2229 (N_2229,N_2072,N_2125);
or U2230 (N_2230,N_2195,N_2022);
or U2231 (N_2231,N_2184,N_2049);
nand U2232 (N_2232,N_2115,N_2188);
nand U2233 (N_2233,N_2130,N_2044);
nor U2234 (N_2234,N_2177,N_2102);
nor U2235 (N_2235,N_2071,N_2133);
or U2236 (N_2236,N_2144,N_2060);
nand U2237 (N_2237,N_2027,N_2117);
nand U2238 (N_2238,N_2076,N_2066);
or U2239 (N_2239,N_2096,N_2182);
nand U2240 (N_2240,N_2097,N_2098);
nand U2241 (N_2241,N_2190,N_2151);
nor U2242 (N_2242,N_2039,N_2135);
nand U2243 (N_2243,N_2166,N_2185);
and U2244 (N_2244,N_2129,N_2181);
or U2245 (N_2245,N_2187,N_2070);
nor U2246 (N_2246,N_2183,N_2137);
or U2247 (N_2247,N_2043,N_2055);
or U2248 (N_2248,N_2179,N_2149);
nand U2249 (N_2249,N_2004,N_2101);
nor U2250 (N_2250,N_2141,N_2168);
or U2251 (N_2251,N_2045,N_2012);
nor U2252 (N_2252,N_2164,N_2107);
nor U2253 (N_2253,N_2082,N_2048);
and U2254 (N_2254,N_2173,N_2197);
nand U2255 (N_2255,N_2078,N_2199);
or U2256 (N_2256,N_2075,N_2058);
nor U2257 (N_2257,N_2106,N_2104);
and U2258 (N_2258,N_2057,N_2178);
nor U2259 (N_2259,N_2134,N_2080);
or U2260 (N_2260,N_2021,N_2128);
nor U2261 (N_2261,N_2109,N_2180);
nor U2262 (N_2262,N_2145,N_2006);
xnor U2263 (N_2263,N_2099,N_2026);
or U2264 (N_2264,N_2196,N_2198);
or U2265 (N_2265,N_2136,N_2132);
nor U2266 (N_2266,N_2016,N_2010);
nor U2267 (N_2267,N_2033,N_2124);
and U2268 (N_2268,N_2008,N_2156);
nand U2269 (N_2269,N_2153,N_2110);
or U2270 (N_2270,N_2163,N_2015);
nor U2271 (N_2271,N_2157,N_2108);
or U2272 (N_2272,N_2041,N_2095);
and U2273 (N_2273,N_2186,N_2193);
and U2274 (N_2274,N_2194,N_2003);
nand U2275 (N_2275,N_2084,N_2077);
and U2276 (N_2276,N_2088,N_2063);
nand U2277 (N_2277,N_2140,N_2035);
or U2278 (N_2278,N_2126,N_2112);
and U2279 (N_2279,N_2094,N_2011);
nand U2280 (N_2280,N_2007,N_2160);
nor U2281 (N_2281,N_2089,N_2032);
and U2282 (N_2282,N_2030,N_2014);
nor U2283 (N_2283,N_2056,N_2038);
nand U2284 (N_2284,N_2172,N_2118);
nor U2285 (N_2285,N_2162,N_2054);
and U2286 (N_2286,N_2113,N_2073);
and U2287 (N_2287,N_2171,N_2139);
and U2288 (N_2288,N_2064,N_2050);
or U2289 (N_2289,N_2090,N_2025);
nor U2290 (N_2290,N_2079,N_2000);
and U2291 (N_2291,N_2111,N_2142);
or U2292 (N_2292,N_2009,N_2002);
nor U2293 (N_2293,N_2167,N_2042);
nand U2294 (N_2294,N_2034,N_2028);
and U2295 (N_2295,N_2150,N_2093);
and U2296 (N_2296,N_2123,N_2046);
or U2297 (N_2297,N_2170,N_2146);
or U2298 (N_2298,N_2013,N_2191);
and U2299 (N_2299,N_2059,N_2005);
and U2300 (N_2300,N_2092,N_2191);
nor U2301 (N_2301,N_2131,N_2126);
nand U2302 (N_2302,N_2071,N_2024);
nor U2303 (N_2303,N_2179,N_2092);
and U2304 (N_2304,N_2026,N_2087);
or U2305 (N_2305,N_2143,N_2010);
nand U2306 (N_2306,N_2029,N_2194);
nand U2307 (N_2307,N_2088,N_2074);
or U2308 (N_2308,N_2005,N_2189);
nand U2309 (N_2309,N_2062,N_2191);
xor U2310 (N_2310,N_2129,N_2114);
and U2311 (N_2311,N_2163,N_2000);
or U2312 (N_2312,N_2009,N_2032);
nor U2313 (N_2313,N_2058,N_2014);
nand U2314 (N_2314,N_2040,N_2012);
nand U2315 (N_2315,N_2108,N_2042);
and U2316 (N_2316,N_2025,N_2128);
and U2317 (N_2317,N_2171,N_2143);
and U2318 (N_2318,N_2018,N_2155);
and U2319 (N_2319,N_2018,N_2139);
or U2320 (N_2320,N_2136,N_2138);
or U2321 (N_2321,N_2021,N_2062);
and U2322 (N_2322,N_2012,N_2078);
nand U2323 (N_2323,N_2191,N_2163);
and U2324 (N_2324,N_2160,N_2060);
or U2325 (N_2325,N_2035,N_2061);
or U2326 (N_2326,N_2017,N_2095);
and U2327 (N_2327,N_2149,N_2068);
nor U2328 (N_2328,N_2169,N_2186);
nand U2329 (N_2329,N_2027,N_2134);
and U2330 (N_2330,N_2089,N_2128);
nand U2331 (N_2331,N_2016,N_2186);
nor U2332 (N_2332,N_2148,N_2015);
and U2333 (N_2333,N_2141,N_2156);
nand U2334 (N_2334,N_2007,N_2094);
and U2335 (N_2335,N_2147,N_2132);
nor U2336 (N_2336,N_2027,N_2129);
and U2337 (N_2337,N_2066,N_2059);
or U2338 (N_2338,N_2177,N_2109);
nor U2339 (N_2339,N_2044,N_2189);
or U2340 (N_2340,N_2071,N_2063);
or U2341 (N_2341,N_2109,N_2153);
nand U2342 (N_2342,N_2148,N_2059);
and U2343 (N_2343,N_2112,N_2034);
and U2344 (N_2344,N_2104,N_2190);
and U2345 (N_2345,N_2160,N_2194);
nand U2346 (N_2346,N_2126,N_2088);
nand U2347 (N_2347,N_2047,N_2098);
nor U2348 (N_2348,N_2119,N_2031);
or U2349 (N_2349,N_2097,N_2111);
or U2350 (N_2350,N_2065,N_2042);
or U2351 (N_2351,N_2125,N_2017);
nor U2352 (N_2352,N_2018,N_2189);
or U2353 (N_2353,N_2010,N_2150);
nand U2354 (N_2354,N_2010,N_2079);
nand U2355 (N_2355,N_2146,N_2016);
nor U2356 (N_2356,N_2096,N_2119);
and U2357 (N_2357,N_2056,N_2115);
nand U2358 (N_2358,N_2058,N_2118);
and U2359 (N_2359,N_2088,N_2085);
or U2360 (N_2360,N_2087,N_2080);
and U2361 (N_2361,N_2146,N_2194);
and U2362 (N_2362,N_2086,N_2117);
nor U2363 (N_2363,N_2026,N_2197);
nor U2364 (N_2364,N_2044,N_2101);
and U2365 (N_2365,N_2061,N_2118);
nand U2366 (N_2366,N_2029,N_2017);
nor U2367 (N_2367,N_2170,N_2006);
or U2368 (N_2368,N_2079,N_2162);
and U2369 (N_2369,N_2049,N_2160);
or U2370 (N_2370,N_2066,N_2087);
nor U2371 (N_2371,N_2085,N_2046);
or U2372 (N_2372,N_2128,N_2002);
or U2373 (N_2373,N_2127,N_2180);
nand U2374 (N_2374,N_2161,N_2073);
or U2375 (N_2375,N_2129,N_2162);
nand U2376 (N_2376,N_2177,N_2080);
or U2377 (N_2377,N_2076,N_2171);
nand U2378 (N_2378,N_2161,N_2003);
nor U2379 (N_2379,N_2022,N_2082);
or U2380 (N_2380,N_2149,N_2119);
nand U2381 (N_2381,N_2108,N_2191);
nand U2382 (N_2382,N_2030,N_2040);
and U2383 (N_2383,N_2026,N_2169);
nand U2384 (N_2384,N_2075,N_2142);
nor U2385 (N_2385,N_2195,N_2000);
nand U2386 (N_2386,N_2095,N_2091);
or U2387 (N_2387,N_2105,N_2094);
nand U2388 (N_2388,N_2089,N_2018);
and U2389 (N_2389,N_2177,N_2064);
or U2390 (N_2390,N_2016,N_2054);
and U2391 (N_2391,N_2001,N_2050);
nand U2392 (N_2392,N_2097,N_2042);
and U2393 (N_2393,N_2109,N_2151);
or U2394 (N_2394,N_2050,N_2000);
or U2395 (N_2395,N_2197,N_2067);
and U2396 (N_2396,N_2099,N_2198);
nand U2397 (N_2397,N_2191,N_2078);
or U2398 (N_2398,N_2026,N_2091);
nor U2399 (N_2399,N_2101,N_2182);
nor U2400 (N_2400,N_2257,N_2386);
nand U2401 (N_2401,N_2384,N_2247);
nor U2402 (N_2402,N_2211,N_2399);
nand U2403 (N_2403,N_2239,N_2360);
nor U2404 (N_2404,N_2346,N_2303);
nand U2405 (N_2405,N_2341,N_2311);
or U2406 (N_2406,N_2245,N_2297);
or U2407 (N_2407,N_2389,N_2294);
nor U2408 (N_2408,N_2235,N_2228);
and U2409 (N_2409,N_2323,N_2373);
nor U2410 (N_2410,N_2327,N_2213);
xnor U2411 (N_2411,N_2387,N_2291);
nor U2412 (N_2412,N_2209,N_2280);
xnor U2413 (N_2413,N_2278,N_2325);
xor U2414 (N_2414,N_2250,N_2249);
nor U2415 (N_2415,N_2261,N_2275);
nand U2416 (N_2416,N_2216,N_2292);
and U2417 (N_2417,N_2259,N_2331);
or U2418 (N_2418,N_2299,N_2304);
and U2419 (N_2419,N_2312,N_2279);
and U2420 (N_2420,N_2368,N_2340);
nand U2421 (N_2421,N_2370,N_2301);
and U2422 (N_2422,N_2240,N_2324);
nor U2423 (N_2423,N_2365,N_2263);
and U2424 (N_2424,N_2273,N_2210);
and U2425 (N_2425,N_2295,N_2395);
and U2426 (N_2426,N_2351,N_2356);
nor U2427 (N_2427,N_2318,N_2313);
nand U2428 (N_2428,N_2272,N_2253);
nor U2429 (N_2429,N_2322,N_2366);
or U2430 (N_2430,N_2338,N_2353);
nand U2431 (N_2431,N_2363,N_2337);
nand U2432 (N_2432,N_2252,N_2359);
nand U2433 (N_2433,N_2394,N_2305);
nand U2434 (N_2434,N_2317,N_2264);
xor U2435 (N_2435,N_2201,N_2220);
or U2436 (N_2436,N_2336,N_2343);
nand U2437 (N_2437,N_2329,N_2350);
and U2438 (N_2438,N_2270,N_2241);
nor U2439 (N_2439,N_2284,N_2229);
nand U2440 (N_2440,N_2334,N_2277);
or U2441 (N_2441,N_2372,N_2208);
and U2442 (N_2442,N_2357,N_2379);
or U2443 (N_2443,N_2282,N_2224);
and U2444 (N_2444,N_2255,N_2276);
nor U2445 (N_2445,N_2328,N_2339);
or U2446 (N_2446,N_2237,N_2333);
or U2447 (N_2447,N_2367,N_2238);
nand U2448 (N_2448,N_2369,N_2335);
nand U2449 (N_2449,N_2381,N_2265);
and U2450 (N_2450,N_2262,N_2388);
nor U2451 (N_2451,N_2308,N_2218);
nor U2452 (N_2452,N_2254,N_2246);
and U2453 (N_2453,N_2309,N_2214);
xor U2454 (N_2454,N_2364,N_2378);
nand U2455 (N_2455,N_2215,N_2287);
nor U2456 (N_2456,N_2227,N_2345);
and U2457 (N_2457,N_2260,N_2298);
and U2458 (N_2458,N_2231,N_2354);
nor U2459 (N_2459,N_2319,N_2377);
nor U2460 (N_2460,N_2385,N_2269);
nand U2461 (N_2461,N_2206,N_2281);
and U2462 (N_2462,N_2212,N_2347);
and U2463 (N_2463,N_2285,N_2217);
nand U2464 (N_2464,N_2314,N_2274);
and U2465 (N_2465,N_2243,N_2266);
nor U2466 (N_2466,N_2236,N_2290);
or U2467 (N_2467,N_2310,N_2267);
and U2468 (N_2468,N_2205,N_2221);
or U2469 (N_2469,N_2283,N_2202);
nor U2470 (N_2470,N_2390,N_2232);
nand U2471 (N_2471,N_2326,N_2315);
and U2472 (N_2472,N_2256,N_2248);
and U2473 (N_2473,N_2306,N_2219);
or U2474 (N_2474,N_2391,N_2271);
and U2475 (N_2475,N_2375,N_2383);
and U2476 (N_2476,N_2234,N_2293);
or U2477 (N_2477,N_2332,N_2223);
and U2478 (N_2478,N_2316,N_2398);
and U2479 (N_2479,N_2230,N_2371);
and U2480 (N_2480,N_2251,N_2362);
nand U2481 (N_2481,N_2396,N_2244);
nor U2482 (N_2482,N_2204,N_2288);
or U2483 (N_2483,N_2330,N_2352);
or U2484 (N_2484,N_2200,N_2374);
nor U2485 (N_2485,N_2307,N_2289);
and U2486 (N_2486,N_2380,N_2397);
and U2487 (N_2487,N_2302,N_2355);
or U2488 (N_2488,N_2376,N_2226);
and U2489 (N_2489,N_2225,N_2348);
or U2490 (N_2490,N_2258,N_2296);
nor U2491 (N_2491,N_2233,N_2358);
or U2492 (N_2492,N_2349,N_2342);
and U2493 (N_2493,N_2382,N_2242);
nor U2494 (N_2494,N_2320,N_2203);
and U2495 (N_2495,N_2393,N_2392);
nor U2496 (N_2496,N_2286,N_2321);
nor U2497 (N_2497,N_2268,N_2207);
nor U2498 (N_2498,N_2222,N_2344);
nor U2499 (N_2499,N_2300,N_2361);
and U2500 (N_2500,N_2322,N_2257);
or U2501 (N_2501,N_2227,N_2349);
nand U2502 (N_2502,N_2312,N_2340);
or U2503 (N_2503,N_2267,N_2326);
or U2504 (N_2504,N_2393,N_2304);
and U2505 (N_2505,N_2373,N_2268);
nand U2506 (N_2506,N_2208,N_2387);
and U2507 (N_2507,N_2223,N_2327);
or U2508 (N_2508,N_2300,N_2265);
or U2509 (N_2509,N_2236,N_2213);
and U2510 (N_2510,N_2307,N_2372);
nor U2511 (N_2511,N_2351,N_2205);
and U2512 (N_2512,N_2352,N_2370);
xor U2513 (N_2513,N_2377,N_2276);
and U2514 (N_2514,N_2271,N_2238);
and U2515 (N_2515,N_2383,N_2261);
nand U2516 (N_2516,N_2281,N_2256);
and U2517 (N_2517,N_2257,N_2312);
and U2518 (N_2518,N_2277,N_2209);
nor U2519 (N_2519,N_2351,N_2311);
or U2520 (N_2520,N_2278,N_2249);
or U2521 (N_2521,N_2322,N_2270);
or U2522 (N_2522,N_2364,N_2356);
or U2523 (N_2523,N_2371,N_2258);
and U2524 (N_2524,N_2337,N_2211);
or U2525 (N_2525,N_2223,N_2305);
xor U2526 (N_2526,N_2372,N_2210);
nand U2527 (N_2527,N_2354,N_2394);
and U2528 (N_2528,N_2330,N_2397);
or U2529 (N_2529,N_2371,N_2305);
nand U2530 (N_2530,N_2220,N_2313);
nand U2531 (N_2531,N_2235,N_2229);
or U2532 (N_2532,N_2324,N_2283);
and U2533 (N_2533,N_2308,N_2314);
or U2534 (N_2534,N_2384,N_2279);
and U2535 (N_2535,N_2319,N_2328);
nand U2536 (N_2536,N_2362,N_2366);
and U2537 (N_2537,N_2298,N_2258);
nor U2538 (N_2538,N_2296,N_2384);
and U2539 (N_2539,N_2232,N_2391);
or U2540 (N_2540,N_2392,N_2321);
or U2541 (N_2541,N_2256,N_2314);
and U2542 (N_2542,N_2324,N_2348);
nor U2543 (N_2543,N_2279,N_2217);
and U2544 (N_2544,N_2289,N_2353);
nand U2545 (N_2545,N_2211,N_2323);
xor U2546 (N_2546,N_2238,N_2311);
nor U2547 (N_2547,N_2322,N_2355);
nand U2548 (N_2548,N_2342,N_2366);
nor U2549 (N_2549,N_2398,N_2273);
and U2550 (N_2550,N_2226,N_2342);
and U2551 (N_2551,N_2357,N_2359);
nand U2552 (N_2552,N_2382,N_2280);
or U2553 (N_2553,N_2274,N_2285);
xnor U2554 (N_2554,N_2226,N_2228);
nand U2555 (N_2555,N_2322,N_2341);
nor U2556 (N_2556,N_2357,N_2203);
or U2557 (N_2557,N_2260,N_2215);
nand U2558 (N_2558,N_2200,N_2357);
or U2559 (N_2559,N_2304,N_2286);
nor U2560 (N_2560,N_2326,N_2260);
nor U2561 (N_2561,N_2292,N_2261);
nor U2562 (N_2562,N_2266,N_2382);
nor U2563 (N_2563,N_2319,N_2330);
or U2564 (N_2564,N_2316,N_2350);
and U2565 (N_2565,N_2334,N_2396);
nor U2566 (N_2566,N_2291,N_2228);
or U2567 (N_2567,N_2286,N_2324);
nor U2568 (N_2568,N_2287,N_2390);
or U2569 (N_2569,N_2210,N_2256);
or U2570 (N_2570,N_2231,N_2287);
and U2571 (N_2571,N_2378,N_2230);
nand U2572 (N_2572,N_2399,N_2296);
and U2573 (N_2573,N_2249,N_2367);
and U2574 (N_2574,N_2366,N_2348);
xnor U2575 (N_2575,N_2320,N_2384);
or U2576 (N_2576,N_2274,N_2230);
nand U2577 (N_2577,N_2208,N_2399);
nand U2578 (N_2578,N_2372,N_2201);
and U2579 (N_2579,N_2269,N_2367);
nand U2580 (N_2580,N_2205,N_2226);
nand U2581 (N_2581,N_2292,N_2257);
nand U2582 (N_2582,N_2304,N_2292);
and U2583 (N_2583,N_2281,N_2243);
or U2584 (N_2584,N_2224,N_2309);
nor U2585 (N_2585,N_2384,N_2235);
nor U2586 (N_2586,N_2287,N_2255);
nor U2587 (N_2587,N_2295,N_2217);
nor U2588 (N_2588,N_2272,N_2387);
nand U2589 (N_2589,N_2250,N_2206);
nand U2590 (N_2590,N_2327,N_2235);
and U2591 (N_2591,N_2294,N_2396);
or U2592 (N_2592,N_2340,N_2392);
nand U2593 (N_2593,N_2343,N_2328);
xnor U2594 (N_2594,N_2211,N_2313);
xor U2595 (N_2595,N_2262,N_2285);
nor U2596 (N_2596,N_2368,N_2298);
or U2597 (N_2597,N_2241,N_2394);
or U2598 (N_2598,N_2233,N_2258);
nor U2599 (N_2599,N_2249,N_2228);
and U2600 (N_2600,N_2544,N_2581);
nand U2601 (N_2601,N_2573,N_2506);
and U2602 (N_2602,N_2424,N_2489);
nand U2603 (N_2603,N_2413,N_2599);
nand U2604 (N_2604,N_2476,N_2449);
and U2605 (N_2605,N_2456,N_2467);
or U2606 (N_2606,N_2479,N_2543);
and U2607 (N_2607,N_2488,N_2561);
nor U2608 (N_2608,N_2509,N_2576);
nand U2609 (N_2609,N_2407,N_2433);
nor U2610 (N_2610,N_2463,N_2500);
nor U2611 (N_2611,N_2527,N_2510);
xor U2612 (N_2612,N_2414,N_2498);
nor U2613 (N_2613,N_2590,N_2437);
or U2614 (N_2614,N_2550,N_2443);
nand U2615 (N_2615,N_2555,N_2459);
nand U2616 (N_2616,N_2520,N_2432);
nor U2617 (N_2617,N_2587,N_2487);
or U2618 (N_2618,N_2406,N_2533);
and U2619 (N_2619,N_2585,N_2570);
nand U2620 (N_2620,N_2503,N_2538);
nand U2621 (N_2621,N_2480,N_2451);
and U2622 (N_2622,N_2472,N_2470);
nor U2623 (N_2623,N_2507,N_2551);
nor U2624 (N_2624,N_2572,N_2468);
nand U2625 (N_2625,N_2534,N_2542);
and U2626 (N_2626,N_2589,N_2401);
nand U2627 (N_2627,N_2427,N_2532);
nor U2628 (N_2628,N_2558,N_2531);
nor U2629 (N_2629,N_2436,N_2548);
nand U2630 (N_2630,N_2522,N_2416);
nand U2631 (N_2631,N_2492,N_2528);
nor U2632 (N_2632,N_2598,N_2518);
nand U2633 (N_2633,N_2428,N_2505);
nand U2634 (N_2634,N_2417,N_2588);
and U2635 (N_2635,N_2577,N_2517);
and U2636 (N_2636,N_2557,N_2495);
or U2637 (N_2637,N_2422,N_2466);
or U2638 (N_2638,N_2482,N_2584);
or U2639 (N_2639,N_2493,N_2594);
nor U2640 (N_2640,N_2567,N_2419);
and U2641 (N_2641,N_2515,N_2425);
nor U2642 (N_2642,N_2485,N_2420);
or U2643 (N_2643,N_2516,N_2444);
or U2644 (N_2644,N_2582,N_2439);
nor U2645 (N_2645,N_2502,N_2474);
and U2646 (N_2646,N_2546,N_2521);
and U2647 (N_2647,N_2409,N_2595);
nand U2648 (N_2648,N_2559,N_2536);
nand U2649 (N_2649,N_2481,N_2494);
or U2650 (N_2650,N_2440,N_2565);
nor U2651 (N_2651,N_2450,N_2513);
nand U2652 (N_2652,N_2402,N_2471);
nand U2653 (N_2653,N_2434,N_2415);
or U2654 (N_2654,N_2569,N_2501);
or U2655 (N_2655,N_2554,N_2537);
or U2656 (N_2656,N_2529,N_2458);
and U2657 (N_2657,N_2597,N_2575);
nand U2658 (N_2658,N_2473,N_2483);
and U2659 (N_2659,N_2423,N_2447);
and U2660 (N_2660,N_2418,N_2579);
and U2661 (N_2661,N_2591,N_2486);
nor U2662 (N_2662,N_2421,N_2519);
or U2663 (N_2663,N_2574,N_2566);
nand U2664 (N_2664,N_2496,N_2469);
nand U2665 (N_2665,N_2553,N_2545);
nor U2666 (N_2666,N_2524,N_2523);
nor U2667 (N_2667,N_2540,N_2526);
and U2668 (N_2668,N_2478,N_2491);
nand U2669 (N_2669,N_2484,N_2441);
nand U2670 (N_2670,N_2455,N_2465);
nor U2671 (N_2671,N_2462,N_2563);
nor U2672 (N_2672,N_2549,N_2556);
nor U2673 (N_2673,N_2435,N_2504);
nor U2674 (N_2674,N_2535,N_2431);
nor U2675 (N_2675,N_2448,N_2512);
nor U2676 (N_2676,N_2541,N_2514);
nor U2677 (N_2677,N_2564,N_2453);
or U2678 (N_2678,N_2580,N_2426);
and U2679 (N_2679,N_2445,N_2410);
nand U2680 (N_2680,N_2454,N_2429);
or U2681 (N_2681,N_2457,N_2530);
nor U2682 (N_2682,N_2430,N_2403);
and U2683 (N_2683,N_2568,N_2405);
or U2684 (N_2684,N_2525,N_2586);
and U2685 (N_2685,N_2552,N_2461);
nor U2686 (N_2686,N_2477,N_2442);
or U2687 (N_2687,N_2475,N_2560);
or U2688 (N_2688,N_2592,N_2547);
or U2689 (N_2689,N_2571,N_2593);
or U2690 (N_2690,N_2508,N_2497);
nor U2691 (N_2691,N_2411,N_2400);
and U2692 (N_2692,N_2490,N_2578);
and U2693 (N_2693,N_2460,N_2446);
nand U2694 (N_2694,N_2562,N_2404);
or U2695 (N_2695,N_2464,N_2408);
nand U2696 (N_2696,N_2499,N_2511);
or U2697 (N_2697,N_2412,N_2583);
or U2698 (N_2698,N_2452,N_2438);
nor U2699 (N_2699,N_2539,N_2596);
nor U2700 (N_2700,N_2409,N_2512);
xor U2701 (N_2701,N_2468,N_2526);
and U2702 (N_2702,N_2576,N_2598);
nor U2703 (N_2703,N_2403,N_2537);
nand U2704 (N_2704,N_2480,N_2563);
nor U2705 (N_2705,N_2533,N_2434);
and U2706 (N_2706,N_2412,N_2509);
and U2707 (N_2707,N_2492,N_2566);
xor U2708 (N_2708,N_2567,N_2444);
or U2709 (N_2709,N_2438,N_2539);
nor U2710 (N_2710,N_2446,N_2573);
xor U2711 (N_2711,N_2412,N_2476);
or U2712 (N_2712,N_2584,N_2513);
nand U2713 (N_2713,N_2469,N_2454);
and U2714 (N_2714,N_2597,N_2588);
nand U2715 (N_2715,N_2519,N_2463);
nor U2716 (N_2716,N_2598,N_2563);
nand U2717 (N_2717,N_2561,N_2464);
and U2718 (N_2718,N_2473,N_2429);
nand U2719 (N_2719,N_2559,N_2512);
or U2720 (N_2720,N_2590,N_2477);
nand U2721 (N_2721,N_2538,N_2489);
nand U2722 (N_2722,N_2576,N_2529);
or U2723 (N_2723,N_2444,N_2574);
and U2724 (N_2724,N_2456,N_2518);
nor U2725 (N_2725,N_2573,N_2483);
nor U2726 (N_2726,N_2525,N_2428);
nand U2727 (N_2727,N_2544,N_2503);
nor U2728 (N_2728,N_2418,N_2456);
nor U2729 (N_2729,N_2498,N_2449);
nand U2730 (N_2730,N_2474,N_2485);
nand U2731 (N_2731,N_2510,N_2519);
nor U2732 (N_2732,N_2574,N_2505);
nand U2733 (N_2733,N_2568,N_2483);
or U2734 (N_2734,N_2491,N_2420);
nor U2735 (N_2735,N_2441,N_2558);
or U2736 (N_2736,N_2554,N_2574);
nand U2737 (N_2737,N_2527,N_2598);
nand U2738 (N_2738,N_2595,N_2411);
or U2739 (N_2739,N_2546,N_2414);
nand U2740 (N_2740,N_2590,N_2424);
and U2741 (N_2741,N_2509,N_2444);
and U2742 (N_2742,N_2534,N_2402);
and U2743 (N_2743,N_2513,N_2511);
or U2744 (N_2744,N_2493,N_2413);
and U2745 (N_2745,N_2442,N_2523);
nor U2746 (N_2746,N_2457,N_2527);
xnor U2747 (N_2747,N_2479,N_2485);
nand U2748 (N_2748,N_2536,N_2579);
nor U2749 (N_2749,N_2553,N_2593);
or U2750 (N_2750,N_2565,N_2529);
nand U2751 (N_2751,N_2583,N_2507);
and U2752 (N_2752,N_2517,N_2560);
nand U2753 (N_2753,N_2479,N_2524);
and U2754 (N_2754,N_2440,N_2525);
and U2755 (N_2755,N_2471,N_2588);
or U2756 (N_2756,N_2506,N_2548);
nand U2757 (N_2757,N_2451,N_2404);
and U2758 (N_2758,N_2487,N_2582);
nand U2759 (N_2759,N_2567,N_2529);
or U2760 (N_2760,N_2413,N_2516);
nor U2761 (N_2761,N_2519,N_2415);
and U2762 (N_2762,N_2577,N_2493);
nor U2763 (N_2763,N_2520,N_2583);
nand U2764 (N_2764,N_2489,N_2401);
or U2765 (N_2765,N_2423,N_2476);
and U2766 (N_2766,N_2468,N_2532);
and U2767 (N_2767,N_2553,N_2469);
and U2768 (N_2768,N_2561,N_2421);
nand U2769 (N_2769,N_2506,N_2558);
nand U2770 (N_2770,N_2444,N_2507);
nand U2771 (N_2771,N_2592,N_2447);
nand U2772 (N_2772,N_2426,N_2522);
and U2773 (N_2773,N_2419,N_2458);
nor U2774 (N_2774,N_2409,N_2496);
and U2775 (N_2775,N_2593,N_2435);
or U2776 (N_2776,N_2407,N_2525);
or U2777 (N_2777,N_2592,N_2549);
or U2778 (N_2778,N_2419,N_2432);
nor U2779 (N_2779,N_2428,N_2443);
nand U2780 (N_2780,N_2408,N_2466);
xnor U2781 (N_2781,N_2536,N_2465);
nor U2782 (N_2782,N_2457,N_2496);
or U2783 (N_2783,N_2484,N_2488);
nand U2784 (N_2784,N_2509,N_2474);
or U2785 (N_2785,N_2590,N_2498);
nor U2786 (N_2786,N_2568,N_2502);
nor U2787 (N_2787,N_2567,N_2554);
nand U2788 (N_2788,N_2432,N_2445);
or U2789 (N_2789,N_2415,N_2496);
and U2790 (N_2790,N_2590,N_2406);
nand U2791 (N_2791,N_2408,N_2475);
and U2792 (N_2792,N_2404,N_2590);
nand U2793 (N_2793,N_2542,N_2570);
nand U2794 (N_2794,N_2476,N_2521);
and U2795 (N_2795,N_2545,N_2579);
nor U2796 (N_2796,N_2572,N_2523);
nor U2797 (N_2797,N_2480,N_2562);
nor U2798 (N_2798,N_2468,N_2576);
nand U2799 (N_2799,N_2444,N_2480);
or U2800 (N_2800,N_2731,N_2743);
nor U2801 (N_2801,N_2721,N_2610);
nand U2802 (N_2802,N_2631,N_2628);
nor U2803 (N_2803,N_2671,N_2755);
nor U2804 (N_2804,N_2772,N_2738);
nor U2805 (N_2805,N_2616,N_2652);
nand U2806 (N_2806,N_2670,N_2717);
nor U2807 (N_2807,N_2748,N_2793);
and U2808 (N_2808,N_2645,N_2678);
nand U2809 (N_2809,N_2653,N_2725);
nor U2810 (N_2810,N_2632,N_2712);
nand U2811 (N_2811,N_2716,N_2714);
and U2812 (N_2812,N_2781,N_2629);
or U2813 (N_2813,N_2609,N_2744);
and U2814 (N_2814,N_2760,N_2777);
and U2815 (N_2815,N_2704,N_2683);
nand U2816 (N_2816,N_2786,N_2727);
nor U2817 (N_2817,N_2797,N_2762);
or U2818 (N_2818,N_2764,N_2633);
nand U2819 (N_2819,N_2680,N_2602);
or U2820 (N_2820,N_2788,N_2695);
and U2821 (N_2821,N_2690,N_2757);
or U2822 (N_2822,N_2728,N_2729);
nand U2823 (N_2823,N_2742,N_2737);
nand U2824 (N_2824,N_2622,N_2649);
nor U2825 (N_2825,N_2705,N_2644);
nand U2826 (N_2826,N_2775,N_2681);
nor U2827 (N_2827,N_2771,N_2794);
nor U2828 (N_2828,N_2657,N_2706);
nand U2829 (N_2829,N_2668,N_2615);
nor U2830 (N_2830,N_2639,N_2654);
nand U2831 (N_2831,N_2650,N_2600);
nand U2832 (N_2832,N_2713,N_2621);
and U2833 (N_2833,N_2720,N_2673);
nand U2834 (N_2834,N_2761,N_2641);
or U2835 (N_2835,N_2611,N_2791);
nor U2836 (N_2836,N_2637,N_2656);
nand U2837 (N_2837,N_2626,N_2672);
nand U2838 (N_2838,N_2686,N_2752);
or U2839 (N_2839,N_2736,N_2784);
or U2840 (N_2840,N_2724,N_2607);
and U2841 (N_2841,N_2711,N_2674);
nor U2842 (N_2842,N_2798,N_2642);
and U2843 (N_2843,N_2799,N_2691);
or U2844 (N_2844,N_2643,N_2785);
and U2845 (N_2845,N_2702,N_2790);
nor U2846 (N_2846,N_2679,N_2718);
or U2847 (N_2847,N_2710,N_2770);
nor U2848 (N_2848,N_2774,N_2665);
nand U2849 (N_2849,N_2659,N_2792);
nand U2850 (N_2850,N_2620,N_2694);
and U2851 (N_2851,N_2676,N_2606);
or U2852 (N_2852,N_2779,N_2789);
or U2853 (N_2853,N_2617,N_2740);
or U2854 (N_2854,N_2783,N_2739);
nand U2855 (N_2855,N_2778,N_2648);
and U2856 (N_2856,N_2701,N_2624);
nand U2857 (N_2857,N_2754,N_2707);
or U2858 (N_2858,N_2758,N_2635);
nor U2859 (N_2859,N_2663,N_2759);
and U2860 (N_2860,N_2708,N_2723);
or U2861 (N_2861,N_2699,N_2769);
nand U2862 (N_2862,N_2741,N_2776);
nor U2863 (N_2863,N_2604,N_2664);
or U2864 (N_2864,N_2638,N_2655);
and U2865 (N_2865,N_2618,N_2608);
and U2866 (N_2866,N_2647,N_2719);
nor U2867 (N_2867,N_2746,N_2756);
and U2868 (N_2868,N_2627,N_2693);
and U2869 (N_2869,N_2750,N_2662);
nand U2870 (N_2870,N_2601,N_2733);
nand U2871 (N_2871,N_2603,N_2796);
nor U2872 (N_2872,N_2749,N_2661);
nor U2873 (N_2873,N_2734,N_2651);
nor U2874 (N_2874,N_2795,N_2605);
nand U2875 (N_2875,N_2625,N_2700);
or U2876 (N_2876,N_2747,N_2667);
and U2877 (N_2877,N_2715,N_2787);
or U2878 (N_2878,N_2636,N_2773);
and U2879 (N_2879,N_2677,N_2732);
and U2880 (N_2880,N_2696,N_2767);
xor U2881 (N_2881,N_2768,N_2692);
nand U2882 (N_2882,N_2730,N_2640);
or U2883 (N_2883,N_2709,N_2684);
or U2884 (N_2884,N_2619,N_2763);
nand U2885 (N_2885,N_2703,N_2623);
or U2886 (N_2886,N_2613,N_2687);
and U2887 (N_2887,N_2630,N_2675);
and U2888 (N_2888,N_2766,N_2780);
or U2889 (N_2889,N_2669,N_2682);
nor U2890 (N_2890,N_2634,N_2745);
xnor U2891 (N_2891,N_2765,N_2697);
and U2892 (N_2892,N_2614,N_2722);
nor U2893 (N_2893,N_2689,N_2726);
or U2894 (N_2894,N_2751,N_2646);
xor U2895 (N_2895,N_2735,N_2698);
nand U2896 (N_2896,N_2658,N_2782);
and U2897 (N_2897,N_2612,N_2685);
nor U2898 (N_2898,N_2660,N_2688);
and U2899 (N_2899,N_2666,N_2753);
or U2900 (N_2900,N_2677,N_2643);
and U2901 (N_2901,N_2650,N_2676);
or U2902 (N_2902,N_2630,N_2741);
nand U2903 (N_2903,N_2767,N_2676);
or U2904 (N_2904,N_2743,N_2786);
or U2905 (N_2905,N_2697,N_2653);
or U2906 (N_2906,N_2694,N_2761);
nor U2907 (N_2907,N_2732,N_2728);
and U2908 (N_2908,N_2688,N_2603);
nand U2909 (N_2909,N_2671,N_2705);
nand U2910 (N_2910,N_2688,N_2780);
or U2911 (N_2911,N_2655,N_2616);
or U2912 (N_2912,N_2779,N_2724);
nor U2913 (N_2913,N_2643,N_2697);
and U2914 (N_2914,N_2600,N_2772);
nor U2915 (N_2915,N_2780,N_2755);
nor U2916 (N_2916,N_2702,N_2646);
and U2917 (N_2917,N_2602,N_2791);
nand U2918 (N_2918,N_2744,N_2700);
nand U2919 (N_2919,N_2668,N_2631);
or U2920 (N_2920,N_2732,N_2617);
and U2921 (N_2921,N_2621,N_2726);
and U2922 (N_2922,N_2761,N_2781);
and U2923 (N_2923,N_2602,N_2705);
or U2924 (N_2924,N_2744,N_2678);
nor U2925 (N_2925,N_2768,N_2769);
nor U2926 (N_2926,N_2732,N_2766);
and U2927 (N_2927,N_2798,N_2613);
and U2928 (N_2928,N_2779,N_2677);
and U2929 (N_2929,N_2729,N_2787);
nand U2930 (N_2930,N_2654,N_2742);
nor U2931 (N_2931,N_2619,N_2738);
xor U2932 (N_2932,N_2610,N_2763);
and U2933 (N_2933,N_2709,N_2668);
nor U2934 (N_2934,N_2623,N_2676);
and U2935 (N_2935,N_2683,N_2710);
nand U2936 (N_2936,N_2791,N_2644);
nor U2937 (N_2937,N_2759,N_2656);
and U2938 (N_2938,N_2783,N_2781);
nand U2939 (N_2939,N_2728,N_2691);
and U2940 (N_2940,N_2751,N_2665);
nor U2941 (N_2941,N_2684,N_2772);
nand U2942 (N_2942,N_2715,N_2618);
nor U2943 (N_2943,N_2623,N_2627);
or U2944 (N_2944,N_2739,N_2629);
or U2945 (N_2945,N_2603,N_2659);
or U2946 (N_2946,N_2600,N_2613);
nor U2947 (N_2947,N_2617,N_2627);
and U2948 (N_2948,N_2675,N_2665);
and U2949 (N_2949,N_2686,N_2714);
nor U2950 (N_2950,N_2648,N_2750);
and U2951 (N_2951,N_2733,N_2698);
and U2952 (N_2952,N_2681,N_2720);
and U2953 (N_2953,N_2772,N_2693);
and U2954 (N_2954,N_2691,N_2623);
and U2955 (N_2955,N_2727,N_2701);
nor U2956 (N_2956,N_2679,N_2794);
nor U2957 (N_2957,N_2703,N_2682);
or U2958 (N_2958,N_2799,N_2656);
or U2959 (N_2959,N_2759,N_2778);
or U2960 (N_2960,N_2654,N_2609);
nand U2961 (N_2961,N_2742,N_2659);
nand U2962 (N_2962,N_2603,N_2673);
nor U2963 (N_2963,N_2716,N_2635);
nor U2964 (N_2964,N_2770,N_2609);
and U2965 (N_2965,N_2747,N_2716);
or U2966 (N_2966,N_2614,N_2727);
and U2967 (N_2967,N_2617,N_2770);
and U2968 (N_2968,N_2716,N_2601);
and U2969 (N_2969,N_2662,N_2789);
nor U2970 (N_2970,N_2609,N_2712);
nand U2971 (N_2971,N_2720,N_2758);
nor U2972 (N_2972,N_2718,N_2659);
nor U2973 (N_2973,N_2781,N_2625);
nand U2974 (N_2974,N_2649,N_2742);
or U2975 (N_2975,N_2733,N_2751);
nand U2976 (N_2976,N_2684,N_2673);
and U2977 (N_2977,N_2700,N_2663);
and U2978 (N_2978,N_2700,N_2604);
and U2979 (N_2979,N_2741,N_2685);
nand U2980 (N_2980,N_2600,N_2666);
nand U2981 (N_2981,N_2739,N_2662);
or U2982 (N_2982,N_2687,N_2756);
nor U2983 (N_2983,N_2788,N_2707);
nor U2984 (N_2984,N_2795,N_2665);
or U2985 (N_2985,N_2724,N_2780);
nor U2986 (N_2986,N_2791,N_2652);
nand U2987 (N_2987,N_2749,N_2630);
nor U2988 (N_2988,N_2610,N_2744);
nor U2989 (N_2989,N_2783,N_2680);
or U2990 (N_2990,N_2785,N_2698);
or U2991 (N_2991,N_2768,N_2792);
and U2992 (N_2992,N_2739,N_2799);
nor U2993 (N_2993,N_2642,N_2693);
and U2994 (N_2994,N_2743,N_2697);
or U2995 (N_2995,N_2755,N_2797);
nand U2996 (N_2996,N_2666,N_2618);
nor U2997 (N_2997,N_2691,N_2746);
or U2998 (N_2998,N_2603,N_2710);
xor U2999 (N_2999,N_2676,N_2741);
or U3000 (N_3000,N_2935,N_2955);
nand U3001 (N_3001,N_2843,N_2862);
or U3002 (N_3002,N_2907,N_2884);
or U3003 (N_3003,N_2880,N_2952);
or U3004 (N_3004,N_2906,N_2897);
nor U3005 (N_3005,N_2981,N_2826);
or U3006 (N_3006,N_2943,N_2921);
or U3007 (N_3007,N_2805,N_2970);
or U3008 (N_3008,N_2854,N_2829);
and U3009 (N_3009,N_2992,N_2817);
nand U3010 (N_3010,N_2890,N_2808);
nand U3011 (N_3011,N_2813,N_2998);
nand U3012 (N_3012,N_2911,N_2987);
or U3013 (N_3013,N_2836,N_2940);
nor U3014 (N_3014,N_2942,N_2807);
nor U3015 (N_3015,N_2840,N_2929);
and U3016 (N_3016,N_2923,N_2954);
and U3017 (N_3017,N_2971,N_2913);
nor U3018 (N_3018,N_2920,N_2861);
nor U3019 (N_3019,N_2977,N_2865);
and U3020 (N_3020,N_2956,N_2803);
nor U3021 (N_3021,N_2902,N_2887);
nor U3022 (N_3022,N_2868,N_2881);
nor U3023 (N_3023,N_2975,N_2823);
and U3024 (N_3024,N_2866,N_2922);
nor U3025 (N_3025,N_2997,N_2983);
nor U3026 (N_3026,N_2818,N_2848);
nand U3027 (N_3027,N_2816,N_2908);
or U3028 (N_3028,N_2969,N_2859);
nand U3029 (N_3029,N_2910,N_2972);
or U3030 (N_3030,N_2994,N_2978);
or U3031 (N_3031,N_2871,N_2979);
or U3032 (N_3032,N_2869,N_2968);
or U3033 (N_3033,N_2842,N_2939);
nand U3034 (N_3034,N_2945,N_2837);
or U3035 (N_3035,N_2849,N_2901);
nand U3036 (N_3036,N_2927,N_2928);
nor U3037 (N_3037,N_2894,N_2967);
and U3038 (N_3038,N_2980,N_2905);
or U3039 (N_3039,N_2919,N_2814);
and U3040 (N_3040,N_2909,N_2985);
xor U3041 (N_3041,N_2915,N_2825);
or U3042 (N_3042,N_2851,N_2999);
nand U3043 (N_3043,N_2889,N_2879);
nor U3044 (N_3044,N_2873,N_2930);
nand U3045 (N_3045,N_2802,N_2858);
nor U3046 (N_3046,N_2827,N_2917);
nand U3047 (N_3047,N_2860,N_2811);
nor U3048 (N_3048,N_2990,N_2820);
or U3049 (N_3049,N_2918,N_2872);
or U3050 (N_3050,N_2850,N_2900);
nor U3051 (N_3051,N_2875,N_2870);
nand U3052 (N_3052,N_2941,N_2988);
nand U3053 (N_3053,N_2847,N_2853);
and U3054 (N_3054,N_2833,N_2839);
nand U3055 (N_3055,N_2916,N_2828);
and U3056 (N_3056,N_2931,N_2976);
nor U3057 (N_3057,N_2856,N_2964);
nor U3058 (N_3058,N_2953,N_2819);
and U3059 (N_3059,N_2821,N_2996);
and U3060 (N_3060,N_2835,N_2896);
or U3061 (N_3061,N_2891,N_2801);
and U3062 (N_3062,N_2885,N_2882);
and U3063 (N_3063,N_2950,N_2863);
and U3064 (N_3064,N_2946,N_2838);
nand U3065 (N_3065,N_2960,N_2937);
nand U3066 (N_3066,N_2834,N_2841);
nor U3067 (N_3067,N_2831,N_2852);
nand U3068 (N_3068,N_2957,N_2895);
nor U3069 (N_3069,N_2804,N_2948);
and U3070 (N_3070,N_2993,N_2810);
and U3071 (N_3071,N_2925,N_2857);
and U3072 (N_3072,N_2892,N_2878);
nor U3073 (N_3073,N_2926,N_2989);
or U3074 (N_3074,N_2883,N_2966);
nand U3075 (N_3075,N_2800,N_2973);
nand U3076 (N_3076,N_2904,N_2991);
or U3077 (N_3077,N_2877,N_2903);
or U3078 (N_3078,N_2876,N_2951);
nor U3079 (N_3079,N_2944,N_2888);
nor U3080 (N_3080,N_2914,N_2893);
and U3081 (N_3081,N_2898,N_2959);
nand U3082 (N_3082,N_2958,N_2899);
and U3083 (N_3083,N_2965,N_2832);
nand U3084 (N_3084,N_2995,N_2886);
nor U3085 (N_3085,N_2963,N_2844);
or U3086 (N_3086,N_2830,N_2806);
and U3087 (N_3087,N_2962,N_2932);
nor U3088 (N_3088,N_2845,N_2822);
and U3089 (N_3089,N_2934,N_2933);
nand U3090 (N_3090,N_2974,N_2984);
nor U3091 (N_3091,N_2874,N_2986);
nand U3092 (N_3092,N_2947,N_2936);
and U3093 (N_3093,N_2961,N_2949);
nand U3094 (N_3094,N_2812,N_2982);
and U3095 (N_3095,N_2867,N_2938);
or U3096 (N_3096,N_2855,N_2912);
nand U3097 (N_3097,N_2864,N_2924);
nor U3098 (N_3098,N_2815,N_2824);
nand U3099 (N_3099,N_2809,N_2846);
or U3100 (N_3100,N_2954,N_2827);
or U3101 (N_3101,N_2936,N_2873);
xnor U3102 (N_3102,N_2973,N_2963);
nor U3103 (N_3103,N_2945,N_2991);
or U3104 (N_3104,N_2959,N_2887);
nor U3105 (N_3105,N_2879,N_2806);
or U3106 (N_3106,N_2879,N_2995);
nor U3107 (N_3107,N_2974,N_2989);
or U3108 (N_3108,N_2885,N_2913);
nor U3109 (N_3109,N_2993,N_2897);
nand U3110 (N_3110,N_2869,N_2925);
nor U3111 (N_3111,N_2948,N_2836);
nor U3112 (N_3112,N_2801,N_2924);
nor U3113 (N_3113,N_2914,N_2865);
nor U3114 (N_3114,N_2825,N_2829);
nor U3115 (N_3115,N_2883,N_2841);
nor U3116 (N_3116,N_2953,N_2970);
nand U3117 (N_3117,N_2941,N_2879);
nor U3118 (N_3118,N_2847,N_2998);
nand U3119 (N_3119,N_2915,N_2927);
nor U3120 (N_3120,N_2856,N_2867);
and U3121 (N_3121,N_2914,N_2835);
or U3122 (N_3122,N_2978,N_2893);
nor U3123 (N_3123,N_2926,N_2978);
and U3124 (N_3124,N_2973,N_2997);
xnor U3125 (N_3125,N_2931,N_2860);
and U3126 (N_3126,N_2870,N_2928);
or U3127 (N_3127,N_2977,N_2911);
nand U3128 (N_3128,N_2998,N_2953);
nand U3129 (N_3129,N_2955,N_2849);
nand U3130 (N_3130,N_2807,N_2818);
or U3131 (N_3131,N_2876,N_2873);
or U3132 (N_3132,N_2960,N_2866);
or U3133 (N_3133,N_2952,N_2872);
nand U3134 (N_3134,N_2873,N_2932);
nor U3135 (N_3135,N_2853,N_2902);
nand U3136 (N_3136,N_2862,N_2893);
or U3137 (N_3137,N_2867,N_2909);
and U3138 (N_3138,N_2881,N_2802);
or U3139 (N_3139,N_2837,N_2927);
nand U3140 (N_3140,N_2898,N_2904);
and U3141 (N_3141,N_2930,N_2998);
or U3142 (N_3142,N_2820,N_2926);
nand U3143 (N_3143,N_2955,N_2963);
nand U3144 (N_3144,N_2916,N_2889);
or U3145 (N_3145,N_2815,N_2808);
or U3146 (N_3146,N_2829,N_2981);
or U3147 (N_3147,N_2951,N_2866);
or U3148 (N_3148,N_2885,N_2952);
or U3149 (N_3149,N_2817,N_2833);
nor U3150 (N_3150,N_2899,N_2866);
nor U3151 (N_3151,N_2850,N_2963);
and U3152 (N_3152,N_2916,N_2854);
nor U3153 (N_3153,N_2906,N_2991);
xnor U3154 (N_3154,N_2977,N_2899);
or U3155 (N_3155,N_2929,N_2995);
and U3156 (N_3156,N_2843,N_2916);
and U3157 (N_3157,N_2803,N_2976);
nor U3158 (N_3158,N_2926,N_2807);
or U3159 (N_3159,N_2902,N_2952);
nor U3160 (N_3160,N_2988,N_2893);
and U3161 (N_3161,N_2961,N_2883);
nand U3162 (N_3162,N_2866,N_2875);
nor U3163 (N_3163,N_2997,N_2851);
nor U3164 (N_3164,N_2895,N_2894);
nor U3165 (N_3165,N_2913,N_2908);
or U3166 (N_3166,N_2930,N_2986);
and U3167 (N_3167,N_2833,N_2807);
or U3168 (N_3168,N_2924,N_2998);
and U3169 (N_3169,N_2905,N_2812);
or U3170 (N_3170,N_2854,N_2889);
nor U3171 (N_3171,N_2959,N_2990);
and U3172 (N_3172,N_2825,N_2875);
nand U3173 (N_3173,N_2918,N_2853);
or U3174 (N_3174,N_2878,N_2936);
and U3175 (N_3175,N_2833,N_2842);
or U3176 (N_3176,N_2890,N_2935);
or U3177 (N_3177,N_2966,N_2952);
or U3178 (N_3178,N_2904,N_2936);
nand U3179 (N_3179,N_2910,N_2854);
or U3180 (N_3180,N_2863,N_2908);
nor U3181 (N_3181,N_2961,N_2890);
nor U3182 (N_3182,N_2903,N_2935);
nand U3183 (N_3183,N_2916,N_2894);
xnor U3184 (N_3184,N_2853,N_2928);
or U3185 (N_3185,N_2941,N_2947);
nand U3186 (N_3186,N_2963,N_2950);
or U3187 (N_3187,N_2939,N_2817);
nand U3188 (N_3188,N_2951,N_2810);
or U3189 (N_3189,N_2924,N_2867);
nor U3190 (N_3190,N_2999,N_2915);
and U3191 (N_3191,N_2833,N_2902);
nand U3192 (N_3192,N_2945,N_2912);
and U3193 (N_3193,N_2826,N_2866);
and U3194 (N_3194,N_2980,N_2951);
xor U3195 (N_3195,N_2907,N_2845);
nand U3196 (N_3196,N_2999,N_2907);
and U3197 (N_3197,N_2817,N_2912);
and U3198 (N_3198,N_2963,N_2992);
and U3199 (N_3199,N_2832,N_2990);
nor U3200 (N_3200,N_3115,N_3029);
nand U3201 (N_3201,N_3132,N_3060);
or U3202 (N_3202,N_3116,N_3030);
or U3203 (N_3203,N_3001,N_3148);
or U3204 (N_3204,N_3051,N_3179);
or U3205 (N_3205,N_3174,N_3171);
or U3206 (N_3206,N_3099,N_3150);
nor U3207 (N_3207,N_3141,N_3111);
and U3208 (N_3208,N_3002,N_3126);
nand U3209 (N_3209,N_3197,N_3076);
xor U3210 (N_3210,N_3033,N_3080);
or U3211 (N_3211,N_3130,N_3008);
or U3212 (N_3212,N_3067,N_3157);
or U3213 (N_3213,N_3125,N_3146);
or U3214 (N_3214,N_3101,N_3084);
nor U3215 (N_3215,N_3155,N_3050);
nand U3216 (N_3216,N_3059,N_3164);
nor U3217 (N_3217,N_3031,N_3068);
and U3218 (N_3218,N_3052,N_3118);
nand U3219 (N_3219,N_3172,N_3124);
nor U3220 (N_3220,N_3131,N_3191);
nor U3221 (N_3221,N_3088,N_3158);
nor U3222 (N_3222,N_3165,N_3036);
or U3223 (N_3223,N_3134,N_3138);
or U3224 (N_3224,N_3018,N_3014);
nor U3225 (N_3225,N_3144,N_3110);
nand U3226 (N_3226,N_3169,N_3047);
and U3227 (N_3227,N_3085,N_3093);
nand U3228 (N_3228,N_3135,N_3090);
nand U3229 (N_3229,N_3069,N_3079);
or U3230 (N_3230,N_3034,N_3046);
or U3231 (N_3231,N_3178,N_3058);
nor U3232 (N_3232,N_3007,N_3025);
nor U3233 (N_3233,N_3021,N_3037);
nor U3234 (N_3234,N_3063,N_3077);
or U3235 (N_3235,N_3082,N_3071);
and U3236 (N_3236,N_3012,N_3166);
or U3237 (N_3237,N_3055,N_3020);
nor U3238 (N_3238,N_3149,N_3054);
nor U3239 (N_3239,N_3039,N_3106);
and U3240 (N_3240,N_3086,N_3173);
or U3241 (N_3241,N_3154,N_3091);
nor U3242 (N_3242,N_3167,N_3035);
or U3243 (N_3243,N_3064,N_3040);
nand U3244 (N_3244,N_3177,N_3081);
nand U3245 (N_3245,N_3100,N_3128);
or U3246 (N_3246,N_3153,N_3075);
and U3247 (N_3247,N_3123,N_3083);
nand U3248 (N_3248,N_3094,N_3187);
or U3249 (N_3249,N_3041,N_3193);
nand U3250 (N_3250,N_3192,N_3194);
nor U3251 (N_3251,N_3000,N_3022);
nor U3252 (N_3252,N_3010,N_3015);
or U3253 (N_3253,N_3142,N_3161);
nand U3254 (N_3254,N_3023,N_3038);
and U3255 (N_3255,N_3114,N_3070);
or U3256 (N_3256,N_3105,N_3016);
and U3257 (N_3257,N_3113,N_3073);
and U3258 (N_3258,N_3107,N_3143);
nor U3259 (N_3259,N_3098,N_3043);
and U3260 (N_3260,N_3185,N_3056);
or U3261 (N_3261,N_3074,N_3104);
and U3262 (N_3262,N_3163,N_3019);
nor U3263 (N_3263,N_3089,N_3097);
and U3264 (N_3264,N_3117,N_3199);
and U3265 (N_3265,N_3180,N_3109);
nand U3266 (N_3266,N_3186,N_3184);
nor U3267 (N_3267,N_3182,N_3065);
nor U3268 (N_3268,N_3151,N_3017);
or U3269 (N_3269,N_3120,N_3170);
and U3270 (N_3270,N_3156,N_3072);
and U3271 (N_3271,N_3032,N_3042);
and U3272 (N_3272,N_3139,N_3009);
nor U3273 (N_3273,N_3121,N_3048);
nand U3274 (N_3274,N_3159,N_3112);
nor U3275 (N_3275,N_3137,N_3103);
nor U3276 (N_3276,N_3175,N_3006);
nand U3277 (N_3277,N_3176,N_3005);
nand U3278 (N_3278,N_3162,N_3053);
nor U3279 (N_3279,N_3061,N_3108);
nor U3280 (N_3280,N_3027,N_3057);
nand U3281 (N_3281,N_3140,N_3196);
or U3282 (N_3282,N_3102,N_3013);
xor U3283 (N_3283,N_3092,N_3127);
and U3284 (N_3284,N_3049,N_3122);
nor U3285 (N_3285,N_3062,N_3096);
or U3286 (N_3286,N_3147,N_3066);
nor U3287 (N_3287,N_3045,N_3044);
nor U3288 (N_3288,N_3095,N_3133);
nand U3289 (N_3289,N_3004,N_3003);
nand U3290 (N_3290,N_3190,N_3188);
or U3291 (N_3291,N_3087,N_3181);
nand U3292 (N_3292,N_3011,N_3160);
or U3293 (N_3293,N_3024,N_3026);
or U3294 (N_3294,N_3145,N_3198);
and U3295 (N_3295,N_3078,N_3119);
and U3296 (N_3296,N_3028,N_3152);
nor U3297 (N_3297,N_3183,N_3168);
nand U3298 (N_3298,N_3189,N_3136);
nand U3299 (N_3299,N_3195,N_3129);
nor U3300 (N_3300,N_3055,N_3009);
nand U3301 (N_3301,N_3051,N_3184);
nor U3302 (N_3302,N_3064,N_3173);
nand U3303 (N_3303,N_3168,N_3158);
nor U3304 (N_3304,N_3013,N_3059);
nor U3305 (N_3305,N_3130,N_3159);
nand U3306 (N_3306,N_3010,N_3077);
or U3307 (N_3307,N_3016,N_3122);
nand U3308 (N_3308,N_3054,N_3138);
nor U3309 (N_3309,N_3093,N_3105);
and U3310 (N_3310,N_3032,N_3084);
nor U3311 (N_3311,N_3060,N_3103);
nand U3312 (N_3312,N_3042,N_3157);
and U3313 (N_3313,N_3065,N_3184);
and U3314 (N_3314,N_3003,N_3134);
nand U3315 (N_3315,N_3049,N_3066);
nand U3316 (N_3316,N_3189,N_3054);
nor U3317 (N_3317,N_3080,N_3027);
nand U3318 (N_3318,N_3007,N_3090);
or U3319 (N_3319,N_3019,N_3167);
nand U3320 (N_3320,N_3162,N_3197);
or U3321 (N_3321,N_3192,N_3199);
and U3322 (N_3322,N_3057,N_3124);
nand U3323 (N_3323,N_3087,N_3138);
nor U3324 (N_3324,N_3099,N_3098);
nand U3325 (N_3325,N_3185,N_3093);
nand U3326 (N_3326,N_3045,N_3049);
nor U3327 (N_3327,N_3193,N_3095);
or U3328 (N_3328,N_3067,N_3011);
and U3329 (N_3329,N_3184,N_3149);
nand U3330 (N_3330,N_3176,N_3024);
nor U3331 (N_3331,N_3152,N_3106);
and U3332 (N_3332,N_3174,N_3054);
nand U3333 (N_3333,N_3058,N_3082);
nor U3334 (N_3334,N_3086,N_3183);
nand U3335 (N_3335,N_3149,N_3099);
nor U3336 (N_3336,N_3072,N_3031);
nand U3337 (N_3337,N_3096,N_3053);
and U3338 (N_3338,N_3009,N_3015);
nor U3339 (N_3339,N_3084,N_3135);
or U3340 (N_3340,N_3006,N_3157);
or U3341 (N_3341,N_3153,N_3134);
and U3342 (N_3342,N_3164,N_3023);
or U3343 (N_3343,N_3166,N_3154);
or U3344 (N_3344,N_3148,N_3008);
nor U3345 (N_3345,N_3061,N_3188);
nor U3346 (N_3346,N_3093,N_3086);
and U3347 (N_3347,N_3090,N_3122);
or U3348 (N_3348,N_3030,N_3160);
nor U3349 (N_3349,N_3113,N_3165);
and U3350 (N_3350,N_3156,N_3022);
and U3351 (N_3351,N_3190,N_3009);
nand U3352 (N_3352,N_3125,N_3133);
or U3353 (N_3353,N_3127,N_3186);
nand U3354 (N_3354,N_3133,N_3035);
and U3355 (N_3355,N_3045,N_3167);
nand U3356 (N_3356,N_3020,N_3007);
and U3357 (N_3357,N_3052,N_3117);
and U3358 (N_3358,N_3147,N_3122);
nor U3359 (N_3359,N_3091,N_3070);
and U3360 (N_3360,N_3138,N_3012);
nand U3361 (N_3361,N_3125,N_3030);
nor U3362 (N_3362,N_3007,N_3141);
or U3363 (N_3363,N_3093,N_3177);
nor U3364 (N_3364,N_3081,N_3162);
nand U3365 (N_3365,N_3075,N_3099);
nor U3366 (N_3366,N_3014,N_3070);
or U3367 (N_3367,N_3155,N_3187);
nor U3368 (N_3368,N_3104,N_3060);
and U3369 (N_3369,N_3012,N_3074);
and U3370 (N_3370,N_3125,N_3005);
or U3371 (N_3371,N_3041,N_3002);
nand U3372 (N_3372,N_3198,N_3110);
and U3373 (N_3373,N_3039,N_3154);
nor U3374 (N_3374,N_3076,N_3041);
nand U3375 (N_3375,N_3053,N_3150);
and U3376 (N_3376,N_3198,N_3190);
nor U3377 (N_3377,N_3098,N_3093);
and U3378 (N_3378,N_3089,N_3026);
or U3379 (N_3379,N_3128,N_3145);
or U3380 (N_3380,N_3143,N_3164);
nor U3381 (N_3381,N_3064,N_3013);
nor U3382 (N_3382,N_3024,N_3061);
or U3383 (N_3383,N_3066,N_3118);
nand U3384 (N_3384,N_3079,N_3112);
nor U3385 (N_3385,N_3005,N_3114);
nand U3386 (N_3386,N_3016,N_3037);
nand U3387 (N_3387,N_3160,N_3190);
nor U3388 (N_3388,N_3099,N_3118);
nor U3389 (N_3389,N_3195,N_3067);
and U3390 (N_3390,N_3166,N_3165);
nand U3391 (N_3391,N_3123,N_3036);
nor U3392 (N_3392,N_3036,N_3038);
nand U3393 (N_3393,N_3117,N_3136);
and U3394 (N_3394,N_3196,N_3056);
nand U3395 (N_3395,N_3090,N_3148);
nand U3396 (N_3396,N_3153,N_3149);
and U3397 (N_3397,N_3042,N_3183);
nor U3398 (N_3398,N_3199,N_3091);
or U3399 (N_3399,N_3026,N_3169);
nand U3400 (N_3400,N_3226,N_3372);
nor U3401 (N_3401,N_3223,N_3275);
nand U3402 (N_3402,N_3325,N_3356);
and U3403 (N_3403,N_3228,N_3334);
nand U3404 (N_3404,N_3368,N_3268);
or U3405 (N_3405,N_3305,N_3218);
nor U3406 (N_3406,N_3363,N_3350);
and U3407 (N_3407,N_3213,N_3291);
or U3408 (N_3408,N_3256,N_3339);
and U3409 (N_3409,N_3319,N_3234);
nand U3410 (N_3410,N_3253,N_3353);
and U3411 (N_3411,N_3239,N_3297);
nand U3412 (N_3412,N_3248,N_3358);
or U3413 (N_3413,N_3202,N_3338);
or U3414 (N_3414,N_3337,N_3381);
nand U3415 (N_3415,N_3365,N_3307);
and U3416 (N_3416,N_3242,N_3207);
xor U3417 (N_3417,N_3205,N_3317);
nand U3418 (N_3418,N_3298,N_3238);
xor U3419 (N_3419,N_3294,N_3236);
or U3420 (N_3420,N_3329,N_3378);
and U3421 (N_3421,N_3391,N_3231);
nor U3422 (N_3422,N_3394,N_3349);
xor U3423 (N_3423,N_3357,N_3251);
and U3424 (N_3424,N_3336,N_3264);
nor U3425 (N_3425,N_3392,N_3227);
and U3426 (N_3426,N_3295,N_3375);
and U3427 (N_3427,N_3217,N_3209);
nand U3428 (N_3428,N_3398,N_3343);
and U3429 (N_3429,N_3206,N_3221);
and U3430 (N_3430,N_3265,N_3254);
or U3431 (N_3431,N_3322,N_3214);
nor U3432 (N_3432,N_3237,N_3282);
xor U3433 (N_3433,N_3321,N_3200);
nand U3434 (N_3434,N_3335,N_3276);
xnor U3435 (N_3435,N_3257,N_3341);
nor U3436 (N_3436,N_3272,N_3299);
nand U3437 (N_3437,N_3230,N_3311);
and U3438 (N_3438,N_3313,N_3367);
or U3439 (N_3439,N_3283,N_3285);
nor U3440 (N_3440,N_3352,N_3287);
nor U3441 (N_3441,N_3323,N_3346);
nor U3442 (N_3442,N_3373,N_3312);
and U3443 (N_3443,N_3211,N_3278);
nand U3444 (N_3444,N_3360,N_3284);
and U3445 (N_3445,N_3304,N_3219);
nor U3446 (N_3446,N_3377,N_3288);
or U3447 (N_3447,N_3252,N_3271);
nand U3448 (N_3448,N_3387,N_3233);
nand U3449 (N_3449,N_3386,N_3263);
nand U3450 (N_3450,N_3382,N_3309);
nor U3451 (N_3451,N_3222,N_3332);
or U3452 (N_3452,N_3361,N_3260);
and U3453 (N_3453,N_3303,N_3240);
nand U3454 (N_3454,N_3399,N_3302);
and U3455 (N_3455,N_3362,N_3310);
nand U3456 (N_3456,N_3280,N_3220);
and U3457 (N_3457,N_3397,N_3286);
nand U3458 (N_3458,N_3374,N_3210);
and U3459 (N_3459,N_3243,N_3347);
nor U3460 (N_3460,N_3201,N_3203);
and U3461 (N_3461,N_3333,N_3208);
or U3462 (N_3462,N_3270,N_3384);
nand U3463 (N_3463,N_3340,N_3245);
nor U3464 (N_3464,N_3315,N_3212);
or U3465 (N_3465,N_3232,N_3216);
nor U3466 (N_3466,N_3290,N_3229);
xor U3467 (N_3467,N_3296,N_3348);
and U3468 (N_3468,N_3390,N_3277);
nor U3469 (N_3469,N_3261,N_3327);
nand U3470 (N_3470,N_3306,N_3293);
nor U3471 (N_3471,N_3273,N_3393);
and U3472 (N_3472,N_3345,N_3318);
xnor U3473 (N_3473,N_3289,N_3262);
nand U3474 (N_3474,N_3344,N_3316);
and U3475 (N_3475,N_3331,N_3269);
xor U3476 (N_3476,N_3235,N_3292);
nand U3477 (N_3477,N_3314,N_3355);
nor U3478 (N_3478,N_3351,N_3225);
nor U3479 (N_3479,N_3249,N_3267);
or U3480 (N_3480,N_3215,N_3300);
nor U3481 (N_3481,N_3244,N_3383);
or U3482 (N_3482,N_3204,N_3342);
nor U3483 (N_3483,N_3369,N_3395);
nand U3484 (N_3484,N_3255,N_3241);
or U3485 (N_3485,N_3281,N_3224);
and U3486 (N_3486,N_3246,N_3379);
and U3487 (N_3487,N_3301,N_3266);
and U3488 (N_3488,N_3376,N_3308);
and U3489 (N_3489,N_3326,N_3371);
and U3490 (N_3490,N_3250,N_3328);
nor U3491 (N_3491,N_3354,N_3320);
nor U3492 (N_3492,N_3324,N_3396);
or U3493 (N_3493,N_3259,N_3258);
nand U3494 (N_3494,N_3366,N_3364);
nand U3495 (N_3495,N_3380,N_3330);
or U3496 (N_3496,N_3389,N_3385);
and U3497 (N_3497,N_3274,N_3388);
nand U3498 (N_3498,N_3370,N_3279);
and U3499 (N_3499,N_3247,N_3359);
nor U3500 (N_3500,N_3296,N_3280);
and U3501 (N_3501,N_3337,N_3249);
or U3502 (N_3502,N_3340,N_3258);
nor U3503 (N_3503,N_3380,N_3350);
nand U3504 (N_3504,N_3333,N_3367);
xnor U3505 (N_3505,N_3374,N_3310);
or U3506 (N_3506,N_3326,N_3203);
nor U3507 (N_3507,N_3267,N_3285);
nor U3508 (N_3508,N_3207,N_3399);
nor U3509 (N_3509,N_3313,N_3239);
or U3510 (N_3510,N_3305,N_3223);
nor U3511 (N_3511,N_3258,N_3384);
and U3512 (N_3512,N_3386,N_3348);
xnor U3513 (N_3513,N_3332,N_3233);
and U3514 (N_3514,N_3347,N_3293);
nor U3515 (N_3515,N_3254,N_3306);
nand U3516 (N_3516,N_3350,N_3265);
or U3517 (N_3517,N_3270,N_3389);
or U3518 (N_3518,N_3200,N_3204);
xor U3519 (N_3519,N_3224,N_3249);
nor U3520 (N_3520,N_3203,N_3290);
nand U3521 (N_3521,N_3364,N_3383);
nor U3522 (N_3522,N_3307,N_3204);
and U3523 (N_3523,N_3269,N_3236);
xnor U3524 (N_3524,N_3376,N_3278);
nand U3525 (N_3525,N_3284,N_3202);
or U3526 (N_3526,N_3371,N_3236);
nor U3527 (N_3527,N_3283,N_3274);
nor U3528 (N_3528,N_3262,N_3318);
nand U3529 (N_3529,N_3352,N_3373);
nand U3530 (N_3530,N_3234,N_3260);
nand U3531 (N_3531,N_3212,N_3235);
and U3532 (N_3532,N_3222,N_3246);
nor U3533 (N_3533,N_3328,N_3244);
nand U3534 (N_3534,N_3236,N_3226);
nor U3535 (N_3535,N_3348,N_3325);
or U3536 (N_3536,N_3306,N_3246);
or U3537 (N_3537,N_3239,N_3272);
nor U3538 (N_3538,N_3228,N_3234);
nor U3539 (N_3539,N_3267,N_3261);
nand U3540 (N_3540,N_3321,N_3399);
xnor U3541 (N_3541,N_3321,N_3347);
nand U3542 (N_3542,N_3280,N_3382);
nand U3543 (N_3543,N_3332,N_3265);
and U3544 (N_3544,N_3283,N_3213);
or U3545 (N_3545,N_3373,N_3258);
and U3546 (N_3546,N_3314,N_3329);
or U3547 (N_3547,N_3281,N_3385);
nand U3548 (N_3548,N_3271,N_3234);
nand U3549 (N_3549,N_3328,N_3205);
or U3550 (N_3550,N_3366,N_3334);
nor U3551 (N_3551,N_3258,N_3398);
and U3552 (N_3552,N_3344,N_3318);
nor U3553 (N_3553,N_3310,N_3277);
nand U3554 (N_3554,N_3263,N_3235);
xnor U3555 (N_3555,N_3230,N_3215);
and U3556 (N_3556,N_3343,N_3272);
or U3557 (N_3557,N_3207,N_3276);
and U3558 (N_3558,N_3392,N_3375);
or U3559 (N_3559,N_3357,N_3328);
nand U3560 (N_3560,N_3252,N_3295);
xor U3561 (N_3561,N_3256,N_3319);
and U3562 (N_3562,N_3292,N_3391);
nor U3563 (N_3563,N_3230,N_3251);
nor U3564 (N_3564,N_3235,N_3358);
nand U3565 (N_3565,N_3396,N_3237);
nor U3566 (N_3566,N_3218,N_3204);
nor U3567 (N_3567,N_3383,N_3396);
or U3568 (N_3568,N_3375,N_3274);
nor U3569 (N_3569,N_3226,N_3290);
and U3570 (N_3570,N_3253,N_3336);
nand U3571 (N_3571,N_3205,N_3365);
and U3572 (N_3572,N_3371,N_3374);
nand U3573 (N_3573,N_3213,N_3382);
and U3574 (N_3574,N_3326,N_3254);
nor U3575 (N_3575,N_3327,N_3366);
and U3576 (N_3576,N_3279,N_3379);
and U3577 (N_3577,N_3203,N_3395);
or U3578 (N_3578,N_3310,N_3201);
nor U3579 (N_3579,N_3205,N_3222);
and U3580 (N_3580,N_3218,N_3262);
and U3581 (N_3581,N_3323,N_3381);
nor U3582 (N_3582,N_3385,N_3206);
nand U3583 (N_3583,N_3275,N_3312);
nand U3584 (N_3584,N_3288,N_3389);
and U3585 (N_3585,N_3355,N_3337);
and U3586 (N_3586,N_3219,N_3380);
and U3587 (N_3587,N_3325,N_3247);
nand U3588 (N_3588,N_3387,N_3269);
xor U3589 (N_3589,N_3245,N_3366);
and U3590 (N_3590,N_3241,N_3275);
and U3591 (N_3591,N_3329,N_3256);
and U3592 (N_3592,N_3266,N_3310);
or U3593 (N_3593,N_3237,N_3325);
and U3594 (N_3594,N_3375,N_3298);
and U3595 (N_3595,N_3262,N_3263);
nand U3596 (N_3596,N_3235,N_3253);
nor U3597 (N_3597,N_3392,N_3341);
nor U3598 (N_3598,N_3202,N_3331);
nand U3599 (N_3599,N_3223,N_3287);
nor U3600 (N_3600,N_3542,N_3493);
and U3601 (N_3601,N_3440,N_3581);
or U3602 (N_3602,N_3519,N_3481);
and U3603 (N_3603,N_3462,N_3489);
nand U3604 (N_3604,N_3591,N_3575);
nor U3605 (N_3605,N_3419,N_3594);
or U3606 (N_3606,N_3566,N_3514);
nor U3607 (N_3607,N_3459,N_3523);
nor U3608 (N_3608,N_3404,N_3592);
nor U3609 (N_3609,N_3507,N_3454);
nor U3610 (N_3610,N_3551,N_3495);
or U3611 (N_3611,N_3573,N_3416);
and U3612 (N_3612,N_3490,N_3472);
and U3613 (N_3613,N_3401,N_3593);
or U3614 (N_3614,N_3429,N_3587);
and U3615 (N_3615,N_3569,N_3570);
nand U3616 (N_3616,N_3485,N_3470);
or U3617 (N_3617,N_3518,N_3576);
or U3618 (N_3618,N_3497,N_3565);
or U3619 (N_3619,N_3492,N_3448);
xnor U3620 (N_3620,N_3502,N_3484);
nor U3621 (N_3621,N_3597,N_3482);
nor U3622 (N_3622,N_3579,N_3550);
nand U3623 (N_3623,N_3410,N_3577);
and U3624 (N_3624,N_3450,N_3438);
and U3625 (N_3625,N_3421,N_3457);
nand U3626 (N_3626,N_3595,N_3557);
xor U3627 (N_3627,N_3411,N_3553);
and U3628 (N_3628,N_3415,N_3406);
and U3629 (N_3629,N_3451,N_3418);
and U3630 (N_3630,N_3494,N_3455);
and U3631 (N_3631,N_3473,N_3412);
or U3632 (N_3632,N_3467,N_3478);
and U3633 (N_3633,N_3430,N_3505);
nand U3634 (N_3634,N_3476,N_3506);
nand U3635 (N_3635,N_3503,N_3483);
or U3636 (N_3636,N_3538,N_3558);
nand U3637 (N_3637,N_3555,N_3517);
or U3638 (N_3638,N_3487,N_3532);
nor U3639 (N_3639,N_3586,N_3515);
nand U3640 (N_3640,N_3414,N_3516);
nor U3641 (N_3641,N_3449,N_3425);
xnor U3642 (N_3642,N_3402,N_3545);
nor U3643 (N_3643,N_3442,N_3567);
nand U3644 (N_3644,N_3536,N_3599);
or U3645 (N_3645,N_3413,N_3544);
or U3646 (N_3646,N_3578,N_3443);
or U3647 (N_3647,N_3403,N_3469);
nor U3648 (N_3648,N_3496,N_3466);
and U3649 (N_3649,N_3564,N_3480);
nand U3650 (N_3650,N_3491,N_3585);
nor U3651 (N_3651,N_3409,N_3488);
or U3652 (N_3652,N_3486,N_3471);
or U3653 (N_3653,N_3468,N_3511);
and U3654 (N_3654,N_3537,N_3441);
or U3655 (N_3655,N_3400,N_3498);
nor U3656 (N_3656,N_3431,N_3549);
or U3657 (N_3657,N_3420,N_3408);
or U3658 (N_3658,N_3439,N_3583);
nand U3659 (N_3659,N_3479,N_3590);
or U3660 (N_3660,N_3547,N_3526);
or U3661 (N_3661,N_3562,N_3530);
nand U3662 (N_3662,N_3465,N_3509);
and U3663 (N_3663,N_3463,N_3433);
or U3664 (N_3664,N_3571,N_3444);
nor U3665 (N_3665,N_3531,N_3461);
nor U3666 (N_3666,N_3572,N_3426);
nor U3667 (N_3667,N_3422,N_3525);
nor U3668 (N_3668,N_3554,N_3546);
and U3669 (N_3669,N_3520,N_3522);
nor U3670 (N_3670,N_3453,N_3574);
nor U3671 (N_3671,N_3500,N_3452);
or U3672 (N_3672,N_3533,N_3582);
nand U3673 (N_3673,N_3475,N_3513);
and U3674 (N_3674,N_3543,N_3499);
and U3675 (N_3675,N_3435,N_3501);
and U3676 (N_3676,N_3437,N_3596);
nor U3677 (N_3677,N_3539,N_3588);
nand U3678 (N_3678,N_3512,N_3504);
and U3679 (N_3679,N_3589,N_3434);
or U3680 (N_3680,N_3598,N_3527);
or U3681 (N_3681,N_3427,N_3432);
nand U3682 (N_3682,N_3584,N_3529);
and U3683 (N_3683,N_3464,N_3460);
and U3684 (N_3684,N_3560,N_3477);
and U3685 (N_3685,N_3456,N_3508);
nand U3686 (N_3686,N_3417,N_3563);
nand U3687 (N_3687,N_3446,N_3568);
nand U3688 (N_3688,N_3474,N_3559);
and U3689 (N_3689,N_3540,N_3407);
and U3690 (N_3690,N_3445,N_3534);
nor U3691 (N_3691,N_3580,N_3428);
nand U3692 (N_3692,N_3510,N_3524);
or U3693 (N_3693,N_3541,N_3535);
nand U3694 (N_3694,N_3521,N_3423);
nor U3695 (N_3695,N_3556,N_3447);
nand U3696 (N_3696,N_3548,N_3561);
or U3697 (N_3697,N_3424,N_3528);
nor U3698 (N_3698,N_3552,N_3458);
and U3699 (N_3699,N_3436,N_3405);
nor U3700 (N_3700,N_3502,N_3400);
or U3701 (N_3701,N_3576,N_3594);
and U3702 (N_3702,N_3441,N_3582);
and U3703 (N_3703,N_3419,N_3513);
nand U3704 (N_3704,N_3491,N_3521);
and U3705 (N_3705,N_3448,N_3409);
or U3706 (N_3706,N_3500,N_3592);
nor U3707 (N_3707,N_3487,N_3461);
nor U3708 (N_3708,N_3584,N_3425);
and U3709 (N_3709,N_3512,N_3425);
or U3710 (N_3710,N_3407,N_3505);
and U3711 (N_3711,N_3418,N_3485);
nor U3712 (N_3712,N_3412,N_3510);
nand U3713 (N_3713,N_3475,N_3528);
and U3714 (N_3714,N_3533,N_3484);
and U3715 (N_3715,N_3519,N_3598);
or U3716 (N_3716,N_3510,N_3476);
xnor U3717 (N_3717,N_3582,N_3574);
or U3718 (N_3718,N_3407,N_3583);
or U3719 (N_3719,N_3443,N_3521);
nor U3720 (N_3720,N_3528,N_3577);
nor U3721 (N_3721,N_3482,N_3592);
nor U3722 (N_3722,N_3520,N_3400);
nand U3723 (N_3723,N_3529,N_3485);
nand U3724 (N_3724,N_3404,N_3561);
or U3725 (N_3725,N_3543,N_3512);
and U3726 (N_3726,N_3414,N_3496);
nand U3727 (N_3727,N_3562,N_3535);
and U3728 (N_3728,N_3554,N_3523);
or U3729 (N_3729,N_3554,N_3417);
nand U3730 (N_3730,N_3431,N_3578);
and U3731 (N_3731,N_3462,N_3448);
or U3732 (N_3732,N_3493,N_3517);
or U3733 (N_3733,N_3425,N_3578);
nand U3734 (N_3734,N_3593,N_3574);
nor U3735 (N_3735,N_3524,N_3499);
or U3736 (N_3736,N_3581,N_3562);
nor U3737 (N_3737,N_3535,N_3546);
nor U3738 (N_3738,N_3541,N_3457);
or U3739 (N_3739,N_3491,N_3457);
nand U3740 (N_3740,N_3417,N_3444);
or U3741 (N_3741,N_3473,N_3493);
nand U3742 (N_3742,N_3469,N_3507);
or U3743 (N_3743,N_3535,N_3504);
nand U3744 (N_3744,N_3403,N_3576);
and U3745 (N_3745,N_3440,N_3403);
and U3746 (N_3746,N_3557,N_3462);
nand U3747 (N_3747,N_3422,N_3508);
xnor U3748 (N_3748,N_3456,N_3478);
nor U3749 (N_3749,N_3529,N_3474);
or U3750 (N_3750,N_3595,N_3548);
and U3751 (N_3751,N_3478,N_3463);
nor U3752 (N_3752,N_3432,N_3466);
and U3753 (N_3753,N_3572,N_3467);
or U3754 (N_3754,N_3530,N_3575);
xnor U3755 (N_3755,N_3437,N_3421);
xnor U3756 (N_3756,N_3540,N_3403);
or U3757 (N_3757,N_3545,N_3531);
nand U3758 (N_3758,N_3562,N_3409);
or U3759 (N_3759,N_3549,N_3512);
nand U3760 (N_3760,N_3405,N_3540);
and U3761 (N_3761,N_3572,N_3401);
nor U3762 (N_3762,N_3455,N_3498);
nor U3763 (N_3763,N_3499,N_3451);
nand U3764 (N_3764,N_3550,N_3485);
nor U3765 (N_3765,N_3563,N_3578);
nor U3766 (N_3766,N_3458,N_3402);
or U3767 (N_3767,N_3513,N_3545);
nand U3768 (N_3768,N_3498,N_3487);
nor U3769 (N_3769,N_3528,N_3597);
nand U3770 (N_3770,N_3511,N_3502);
nor U3771 (N_3771,N_3421,N_3577);
or U3772 (N_3772,N_3585,N_3424);
or U3773 (N_3773,N_3452,N_3583);
nor U3774 (N_3774,N_3541,N_3440);
or U3775 (N_3775,N_3559,N_3435);
nor U3776 (N_3776,N_3460,N_3438);
nor U3777 (N_3777,N_3559,N_3411);
or U3778 (N_3778,N_3427,N_3442);
nand U3779 (N_3779,N_3524,N_3432);
and U3780 (N_3780,N_3447,N_3504);
nor U3781 (N_3781,N_3505,N_3516);
and U3782 (N_3782,N_3590,N_3550);
and U3783 (N_3783,N_3439,N_3429);
nand U3784 (N_3784,N_3463,N_3436);
nand U3785 (N_3785,N_3524,N_3558);
and U3786 (N_3786,N_3487,N_3442);
or U3787 (N_3787,N_3452,N_3536);
or U3788 (N_3788,N_3461,N_3585);
nand U3789 (N_3789,N_3529,N_3502);
and U3790 (N_3790,N_3492,N_3428);
or U3791 (N_3791,N_3524,N_3435);
nor U3792 (N_3792,N_3535,N_3433);
and U3793 (N_3793,N_3550,N_3596);
nor U3794 (N_3794,N_3414,N_3590);
or U3795 (N_3795,N_3535,N_3522);
nand U3796 (N_3796,N_3588,N_3597);
and U3797 (N_3797,N_3510,N_3436);
nand U3798 (N_3798,N_3425,N_3494);
xor U3799 (N_3799,N_3521,N_3546);
or U3800 (N_3800,N_3770,N_3634);
and U3801 (N_3801,N_3755,N_3718);
nor U3802 (N_3802,N_3762,N_3607);
or U3803 (N_3803,N_3749,N_3776);
or U3804 (N_3804,N_3766,N_3631);
and U3805 (N_3805,N_3761,N_3681);
xnor U3806 (N_3806,N_3656,N_3626);
nor U3807 (N_3807,N_3719,N_3696);
or U3808 (N_3808,N_3715,N_3621);
or U3809 (N_3809,N_3791,N_3627);
and U3810 (N_3810,N_3654,N_3773);
nor U3811 (N_3811,N_3793,N_3643);
and U3812 (N_3812,N_3614,N_3774);
and U3813 (N_3813,N_3660,N_3727);
nand U3814 (N_3814,N_3694,N_3688);
and U3815 (N_3815,N_3737,N_3658);
nor U3816 (N_3816,N_3690,N_3796);
and U3817 (N_3817,N_3680,N_3742);
nor U3818 (N_3818,N_3610,N_3780);
nor U3819 (N_3819,N_3635,N_3782);
nor U3820 (N_3820,N_3600,N_3752);
and U3821 (N_3821,N_3760,N_3717);
and U3822 (N_3822,N_3666,N_3733);
or U3823 (N_3823,N_3701,N_3726);
or U3824 (N_3824,N_3678,N_3601);
nand U3825 (N_3825,N_3675,N_3662);
nand U3826 (N_3826,N_3655,N_3778);
and U3827 (N_3827,N_3728,N_3744);
and U3828 (N_3828,N_3753,N_3630);
and U3829 (N_3829,N_3628,N_3757);
or U3830 (N_3830,N_3732,N_3608);
or U3831 (N_3831,N_3671,N_3673);
and U3832 (N_3832,N_3798,N_3619);
and U3833 (N_3833,N_3731,N_3786);
nor U3834 (N_3834,N_3777,N_3613);
nor U3835 (N_3835,N_3652,N_3764);
nand U3836 (N_3836,N_3784,N_3771);
or U3837 (N_3837,N_3637,N_3738);
or U3838 (N_3838,N_3699,N_3772);
nand U3839 (N_3839,N_3788,N_3661);
nor U3840 (N_3840,N_3783,N_3676);
nand U3841 (N_3841,N_3704,N_3792);
nor U3842 (N_3842,N_3725,N_3768);
and U3843 (N_3843,N_3674,N_3657);
nand U3844 (N_3844,N_3743,N_3650);
and U3845 (N_3845,N_3629,N_3741);
nor U3846 (N_3846,N_3713,N_3767);
nor U3847 (N_3847,N_3708,N_3616);
and U3848 (N_3848,N_3735,N_3703);
or U3849 (N_3849,N_3721,N_3724);
xor U3850 (N_3850,N_3602,N_3633);
nand U3851 (N_3851,N_3611,N_3645);
and U3852 (N_3852,N_3695,N_3759);
and U3853 (N_3853,N_3697,N_3706);
or U3854 (N_3854,N_3711,N_3740);
and U3855 (N_3855,N_3730,N_3640);
nor U3856 (N_3856,N_3624,N_3687);
nor U3857 (N_3857,N_3682,N_3797);
or U3858 (N_3858,N_3606,N_3604);
and U3859 (N_3859,N_3736,N_3605);
nand U3860 (N_3860,N_3765,N_3641);
and U3861 (N_3861,N_3679,N_3622);
and U3862 (N_3862,N_3653,N_3729);
and U3863 (N_3863,N_3663,N_3720);
nand U3864 (N_3864,N_3665,N_3707);
nor U3865 (N_3865,N_3638,N_3689);
nor U3866 (N_3866,N_3644,N_3672);
or U3867 (N_3867,N_3615,N_3603);
or U3868 (N_3868,N_3789,N_3705);
or U3869 (N_3869,N_3714,N_3642);
nand U3870 (N_3870,N_3648,N_3787);
or U3871 (N_3871,N_3751,N_3794);
or U3872 (N_3872,N_3739,N_3659);
and U3873 (N_3873,N_3785,N_3667);
nand U3874 (N_3874,N_3691,N_3748);
and U3875 (N_3875,N_3779,N_3781);
and U3876 (N_3876,N_3790,N_3612);
nor U3877 (N_3877,N_3693,N_3683);
nor U3878 (N_3878,N_3763,N_3775);
nor U3879 (N_3879,N_3636,N_3686);
nand U3880 (N_3880,N_3722,N_3684);
nor U3881 (N_3881,N_3692,N_3632);
nand U3882 (N_3882,N_3620,N_3754);
and U3883 (N_3883,N_3723,N_3639);
or U3884 (N_3884,N_3685,N_3664);
nor U3885 (N_3885,N_3747,N_3617);
and U3886 (N_3886,N_3702,N_3649);
nor U3887 (N_3887,N_3799,N_3625);
nor U3888 (N_3888,N_3618,N_3758);
or U3889 (N_3889,N_3609,N_3677);
nor U3890 (N_3890,N_3669,N_3746);
xnor U3891 (N_3891,N_3712,N_3670);
nand U3892 (N_3892,N_3710,N_3647);
and U3893 (N_3893,N_3750,N_3716);
or U3894 (N_3894,N_3709,N_3668);
nor U3895 (N_3895,N_3795,N_3651);
nor U3896 (N_3896,N_3623,N_3646);
nand U3897 (N_3897,N_3700,N_3756);
or U3898 (N_3898,N_3769,N_3745);
nor U3899 (N_3899,N_3734,N_3698);
and U3900 (N_3900,N_3633,N_3776);
and U3901 (N_3901,N_3727,N_3634);
nor U3902 (N_3902,N_3797,N_3740);
xor U3903 (N_3903,N_3656,N_3760);
and U3904 (N_3904,N_3733,N_3781);
nor U3905 (N_3905,N_3651,N_3686);
and U3906 (N_3906,N_3787,N_3783);
xor U3907 (N_3907,N_3618,N_3784);
nor U3908 (N_3908,N_3616,N_3680);
nor U3909 (N_3909,N_3726,N_3723);
or U3910 (N_3910,N_3633,N_3706);
nand U3911 (N_3911,N_3772,N_3634);
or U3912 (N_3912,N_3654,N_3777);
nand U3913 (N_3913,N_3658,N_3799);
or U3914 (N_3914,N_3727,N_3756);
and U3915 (N_3915,N_3717,N_3666);
and U3916 (N_3916,N_3655,N_3618);
nand U3917 (N_3917,N_3611,N_3720);
nor U3918 (N_3918,N_3653,N_3642);
nor U3919 (N_3919,N_3601,N_3788);
and U3920 (N_3920,N_3665,N_3658);
xnor U3921 (N_3921,N_3678,N_3615);
nor U3922 (N_3922,N_3630,N_3791);
nor U3923 (N_3923,N_3790,N_3652);
xnor U3924 (N_3924,N_3781,N_3710);
and U3925 (N_3925,N_3790,N_3684);
nor U3926 (N_3926,N_3782,N_3715);
nand U3927 (N_3927,N_3606,N_3677);
or U3928 (N_3928,N_3749,N_3618);
or U3929 (N_3929,N_3749,N_3682);
nor U3930 (N_3930,N_3695,N_3725);
and U3931 (N_3931,N_3732,N_3696);
and U3932 (N_3932,N_3695,N_3743);
or U3933 (N_3933,N_3690,N_3671);
nor U3934 (N_3934,N_3659,N_3729);
nand U3935 (N_3935,N_3631,N_3731);
and U3936 (N_3936,N_3695,N_3717);
nor U3937 (N_3937,N_3779,N_3620);
nand U3938 (N_3938,N_3717,N_3715);
nand U3939 (N_3939,N_3638,N_3602);
and U3940 (N_3940,N_3770,N_3648);
nand U3941 (N_3941,N_3777,N_3667);
nand U3942 (N_3942,N_3631,N_3724);
nor U3943 (N_3943,N_3793,N_3632);
or U3944 (N_3944,N_3682,N_3720);
nand U3945 (N_3945,N_3636,N_3757);
or U3946 (N_3946,N_3668,N_3756);
or U3947 (N_3947,N_3776,N_3613);
and U3948 (N_3948,N_3673,N_3634);
nand U3949 (N_3949,N_3782,N_3647);
or U3950 (N_3950,N_3733,N_3752);
nor U3951 (N_3951,N_3615,N_3662);
or U3952 (N_3952,N_3668,N_3670);
or U3953 (N_3953,N_3746,N_3605);
nor U3954 (N_3954,N_3747,N_3623);
and U3955 (N_3955,N_3761,N_3643);
nor U3956 (N_3956,N_3758,N_3722);
or U3957 (N_3957,N_3730,N_3787);
xnor U3958 (N_3958,N_3614,N_3624);
xor U3959 (N_3959,N_3761,N_3655);
and U3960 (N_3960,N_3741,N_3720);
nor U3961 (N_3961,N_3693,N_3624);
nor U3962 (N_3962,N_3700,N_3694);
or U3963 (N_3963,N_3770,N_3799);
or U3964 (N_3964,N_3635,N_3682);
nand U3965 (N_3965,N_3692,N_3773);
nand U3966 (N_3966,N_3784,N_3651);
nor U3967 (N_3967,N_3670,N_3635);
nor U3968 (N_3968,N_3691,N_3614);
nand U3969 (N_3969,N_3663,N_3677);
and U3970 (N_3970,N_3638,N_3722);
and U3971 (N_3971,N_3670,N_3751);
and U3972 (N_3972,N_3713,N_3678);
nor U3973 (N_3973,N_3708,N_3670);
and U3974 (N_3974,N_3704,N_3744);
nand U3975 (N_3975,N_3780,N_3663);
or U3976 (N_3976,N_3785,N_3728);
nor U3977 (N_3977,N_3673,N_3715);
and U3978 (N_3978,N_3677,N_3630);
nand U3979 (N_3979,N_3673,N_3663);
and U3980 (N_3980,N_3657,N_3652);
nand U3981 (N_3981,N_3719,N_3714);
nand U3982 (N_3982,N_3612,N_3686);
or U3983 (N_3983,N_3681,N_3613);
or U3984 (N_3984,N_3697,N_3625);
and U3985 (N_3985,N_3763,N_3671);
nor U3986 (N_3986,N_3730,N_3624);
nand U3987 (N_3987,N_3659,N_3755);
nand U3988 (N_3988,N_3779,N_3629);
and U3989 (N_3989,N_3667,N_3703);
nand U3990 (N_3990,N_3684,N_3732);
nand U3991 (N_3991,N_3768,N_3778);
nor U3992 (N_3992,N_3661,N_3601);
nor U3993 (N_3993,N_3696,N_3665);
or U3994 (N_3994,N_3714,N_3706);
or U3995 (N_3995,N_3778,N_3697);
nor U3996 (N_3996,N_3611,N_3723);
nor U3997 (N_3997,N_3646,N_3666);
or U3998 (N_3998,N_3756,N_3725);
nor U3999 (N_3999,N_3637,N_3662);
and U4000 (N_4000,N_3922,N_3959);
nor U4001 (N_4001,N_3894,N_3900);
or U4002 (N_4002,N_3826,N_3984);
or U4003 (N_4003,N_3853,N_3884);
or U4004 (N_4004,N_3839,N_3941);
nand U4005 (N_4005,N_3964,N_3869);
and U4006 (N_4006,N_3997,N_3801);
or U4007 (N_4007,N_3851,N_3908);
or U4008 (N_4008,N_3842,N_3887);
and U4009 (N_4009,N_3892,N_3995);
and U4010 (N_4010,N_3871,N_3863);
and U4011 (N_4011,N_3850,N_3870);
or U4012 (N_4012,N_3819,N_3923);
or U4013 (N_4013,N_3823,N_3909);
nor U4014 (N_4014,N_3800,N_3919);
xor U4015 (N_4015,N_3879,N_3804);
or U4016 (N_4016,N_3898,N_3963);
nor U4017 (N_4017,N_3938,N_3873);
and U4018 (N_4018,N_3927,N_3837);
or U4019 (N_4019,N_3974,N_3802);
nand U4020 (N_4020,N_3981,N_3817);
and U4021 (N_4021,N_3972,N_3916);
nor U4022 (N_4022,N_3921,N_3950);
nor U4023 (N_4023,N_3913,N_3814);
xor U4024 (N_4024,N_3838,N_3936);
nor U4025 (N_4025,N_3910,N_3957);
nand U4026 (N_4026,N_3889,N_3880);
and U4027 (N_4027,N_3890,N_3882);
nand U4028 (N_4028,N_3973,N_3815);
or U4029 (N_4029,N_3874,N_3975);
or U4030 (N_4030,N_3846,N_3834);
and U4031 (N_4031,N_3821,N_3867);
nor U4032 (N_4032,N_3847,N_3946);
and U4033 (N_4033,N_3856,N_3977);
nor U4034 (N_4034,N_3808,N_3830);
nor U4035 (N_4035,N_3831,N_3809);
or U4036 (N_4036,N_3862,N_3849);
or U4037 (N_4037,N_3960,N_3929);
nor U4038 (N_4038,N_3967,N_3952);
nand U4039 (N_4039,N_3996,N_3833);
nor U4040 (N_4040,N_3987,N_3843);
nor U4041 (N_4041,N_3990,N_3978);
and U4042 (N_4042,N_3955,N_3881);
nand U4043 (N_4043,N_3812,N_3822);
nor U4044 (N_4044,N_3998,N_3926);
or U4045 (N_4045,N_3876,N_3925);
nor U4046 (N_4046,N_3939,N_3947);
xor U4047 (N_4047,N_3915,N_3983);
xnor U4048 (N_4048,N_3845,N_3994);
nand U4049 (N_4049,N_3848,N_3832);
or U4050 (N_4050,N_3989,N_3827);
nor U4051 (N_4051,N_3979,N_3860);
xor U4052 (N_4052,N_3864,N_3944);
nor U4053 (N_4053,N_3866,N_3852);
or U4054 (N_4054,N_3875,N_3965);
nand U4055 (N_4055,N_3855,N_3859);
and U4056 (N_4056,N_3897,N_3982);
and U4057 (N_4057,N_3906,N_3918);
and U4058 (N_4058,N_3899,N_3858);
nand U4059 (N_4059,N_3888,N_3883);
nor U4060 (N_4060,N_3828,N_3935);
nand U4061 (N_4061,N_3954,N_3953);
or U4062 (N_4062,N_3811,N_3907);
or U4063 (N_4063,N_3904,N_3968);
and U4064 (N_4064,N_3956,N_3886);
nand U4065 (N_4065,N_3825,N_3942);
xor U4066 (N_4066,N_3920,N_3912);
or U4067 (N_4067,N_3854,N_3992);
or U4068 (N_4068,N_3999,N_3969);
and U4069 (N_4069,N_3932,N_3928);
xor U4070 (N_4070,N_3868,N_3807);
and U4071 (N_4071,N_3948,N_3933);
nand U4072 (N_4072,N_3917,N_3962);
nand U4073 (N_4073,N_3940,N_3857);
nor U4074 (N_4074,N_3902,N_3970);
and U4075 (N_4075,N_3958,N_3980);
nand U4076 (N_4076,N_3878,N_3971);
nand U4077 (N_4077,N_3914,N_3885);
nand U4078 (N_4078,N_3816,N_3861);
or U4079 (N_4079,N_3951,N_3810);
or U4080 (N_4080,N_3891,N_3865);
nand U4081 (N_4081,N_3905,N_3986);
and U4082 (N_4082,N_3877,N_3805);
and U4083 (N_4083,N_3901,N_3976);
nor U4084 (N_4084,N_3836,N_3988);
nor U4085 (N_4085,N_3961,N_3945);
nor U4086 (N_4086,N_3985,N_3803);
xor U4087 (N_4087,N_3820,N_3806);
or U4088 (N_4088,N_3991,N_3930);
or U4089 (N_4089,N_3813,N_3829);
nor U4090 (N_4090,N_3896,N_3943);
and U4091 (N_4091,N_3993,N_3903);
or U4092 (N_4092,N_3934,N_3835);
nor U4093 (N_4093,N_3949,N_3893);
or U4094 (N_4094,N_3895,N_3818);
nor U4095 (N_4095,N_3937,N_3824);
nand U4096 (N_4096,N_3872,N_3844);
and U4097 (N_4097,N_3911,N_3924);
nand U4098 (N_4098,N_3966,N_3841);
nand U4099 (N_4099,N_3840,N_3931);
nand U4100 (N_4100,N_3862,N_3842);
nor U4101 (N_4101,N_3960,N_3956);
and U4102 (N_4102,N_3833,N_3851);
and U4103 (N_4103,N_3927,N_3841);
and U4104 (N_4104,N_3913,N_3851);
and U4105 (N_4105,N_3969,N_3892);
and U4106 (N_4106,N_3970,N_3912);
nand U4107 (N_4107,N_3856,N_3958);
nand U4108 (N_4108,N_3949,N_3843);
nor U4109 (N_4109,N_3901,N_3952);
or U4110 (N_4110,N_3955,N_3825);
nand U4111 (N_4111,N_3994,N_3834);
nand U4112 (N_4112,N_3907,N_3905);
nor U4113 (N_4113,N_3984,N_3909);
xnor U4114 (N_4114,N_3998,N_3809);
or U4115 (N_4115,N_3929,N_3931);
nand U4116 (N_4116,N_3848,N_3817);
and U4117 (N_4117,N_3861,N_3987);
or U4118 (N_4118,N_3929,N_3940);
nand U4119 (N_4119,N_3989,N_3996);
nand U4120 (N_4120,N_3817,N_3900);
and U4121 (N_4121,N_3961,N_3834);
or U4122 (N_4122,N_3969,N_3804);
or U4123 (N_4123,N_3828,N_3977);
or U4124 (N_4124,N_3974,N_3800);
nor U4125 (N_4125,N_3944,N_3851);
or U4126 (N_4126,N_3983,N_3911);
nor U4127 (N_4127,N_3842,N_3953);
xor U4128 (N_4128,N_3959,N_3807);
or U4129 (N_4129,N_3815,N_3952);
or U4130 (N_4130,N_3813,N_3980);
or U4131 (N_4131,N_3907,N_3960);
or U4132 (N_4132,N_3888,N_3811);
nand U4133 (N_4133,N_3891,N_3820);
and U4134 (N_4134,N_3974,N_3836);
and U4135 (N_4135,N_3978,N_3928);
or U4136 (N_4136,N_3903,N_3925);
or U4137 (N_4137,N_3814,N_3838);
or U4138 (N_4138,N_3840,N_3898);
nand U4139 (N_4139,N_3864,N_3874);
or U4140 (N_4140,N_3813,N_3808);
nor U4141 (N_4141,N_3886,N_3962);
nand U4142 (N_4142,N_3807,N_3826);
and U4143 (N_4143,N_3862,N_3911);
nor U4144 (N_4144,N_3860,N_3899);
and U4145 (N_4145,N_3883,N_3809);
or U4146 (N_4146,N_3925,N_3947);
and U4147 (N_4147,N_3958,N_3802);
nor U4148 (N_4148,N_3898,N_3985);
nand U4149 (N_4149,N_3912,N_3888);
and U4150 (N_4150,N_3946,N_3863);
and U4151 (N_4151,N_3936,N_3890);
nor U4152 (N_4152,N_3988,N_3998);
or U4153 (N_4153,N_3821,N_3928);
or U4154 (N_4154,N_3961,N_3812);
xnor U4155 (N_4155,N_3884,N_3980);
nor U4156 (N_4156,N_3842,N_3850);
and U4157 (N_4157,N_3864,N_3986);
nor U4158 (N_4158,N_3857,N_3934);
nand U4159 (N_4159,N_3956,N_3875);
nand U4160 (N_4160,N_3833,N_3875);
nand U4161 (N_4161,N_3888,N_3872);
or U4162 (N_4162,N_3928,N_3878);
or U4163 (N_4163,N_3869,N_3848);
nand U4164 (N_4164,N_3820,N_3983);
nor U4165 (N_4165,N_3952,N_3848);
or U4166 (N_4166,N_3976,N_3815);
nand U4167 (N_4167,N_3923,N_3802);
nor U4168 (N_4168,N_3942,N_3824);
and U4169 (N_4169,N_3859,N_3849);
and U4170 (N_4170,N_3831,N_3913);
nand U4171 (N_4171,N_3902,N_3985);
or U4172 (N_4172,N_3900,N_3961);
nand U4173 (N_4173,N_3898,N_3934);
nand U4174 (N_4174,N_3980,N_3867);
nand U4175 (N_4175,N_3920,N_3939);
and U4176 (N_4176,N_3883,N_3873);
nand U4177 (N_4177,N_3820,N_3878);
and U4178 (N_4178,N_3996,N_3901);
and U4179 (N_4179,N_3845,N_3960);
nand U4180 (N_4180,N_3912,N_3856);
and U4181 (N_4181,N_3818,N_3975);
xor U4182 (N_4182,N_3801,N_3834);
nor U4183 (N_4183,N_3954,N_3833);
or U4184 (N_4184,N_3824,N_3941);
or U4185 (N_4185,N_3993,N_3966);
nand U4186 (N_4186,N_3807,N_3811);
and U4187 (N_4187,N_3806,N_3944);
or U4188 (N_4188,N_3868,N_3890);
nand U4189 (N_4189,N_3988,N_3933);
and U4190 (N_4190,N_3841,N_3837);
or U4191 (N_4191,N_3875,N_3892);
nor U4192 (N_4192,N_3989,N_3976);
nor U4193 (N_4193,N_3890,N_3834);
and U4194 (N_4194,N_3911,N_3806);
nor U4195 (N_4195,N_3943,N_3908);
and U4196 (N_4196,N_3937,N_3886);
nor U4197 (N_4197,N_3883,N_3820);
and U4198 (N_4198,N_3982,N_3981);
or U4199 (N_4199,N_3818,N_3972);
nor U4200 (N_4200,N_4194,N_4085);
or U4201 (N_4201,N_4136,N_4193);
or U4202 (N_4202,N_4140,N_4087);
and U4203 (N_4203,N_4090,N_4078);
and U4204 (N_4204,N_4051,N_4190);
nand U4205 (N_4205,N_4132,N_4118);
and U4206 (N_4206,N_4061,N_4153);
and U4207 (N_4207,N_4144,N_4106);
nor U4208 (N_4208,N_4148,N_4006);
or U4209 (N_4209,N_4170,N_4126);
or U4210 (N_4210,N_4198,N_4063);
nand U4211 (N_4211,N_4151,N_4199);
and U4212 (N_4212,N_4089,N_4159);
and U4213 (N_4213,N_4056,N_4023);
and U4214 (N_4214,N_4071,N_4157);
nor U4215 (N_4215,N_4142,N_4017);
nand U4216 (N_4216,N_4066,N_4003);
nand U4217 (N_4217,N_4113,N_4083);
and U4218 (N_4218,N_4031,N_4008);
xnor U4219 (N_4219,N_4044,N_4169);
nor U4220 (N_4220,N_4001,N_4027);
nor U4221 (N_4221,N_4020,N_4036);
nor U4222 (N_4222,N_4077,N_4129);
nor U4223 (N_4223,N_4068,N_4101);
and U4224 (N_4224,N_4168,N_4117);
nand U4225 (N_4225,N_4111,N_4131);
or U4226 (N_4226,N_4011,N_4120);
or U4227 (N_4227,N_4091,N_4004);
or U4228 (N_4228,N_4156,N_4135);
nor U4229 (N_4229,N_4145,N_4139);
nand U4230 (N_4230,N_4035,N_4041);
nor U4231 (N_4231,N_4098,N_4074);
and U4232 (N_4232,N_4103,N_4015);
nor U4233 (N_4233,N_4143,N_4097);
or U4234 (N_4234,N_4161,N_4045);
nand U4235 (N_4235,N_4110,N_4012);
nand U4236 (N_4236,N_4180,N_4123);
and U4237 (N_4237,N_4178,N_4073);
or U4238 (N_4238,N_4029,N_4160);
nor U4239 (N_4239,N_4185,N_4171);
or U4240 (N_4240,N_4146,N_4076);
or U4241 (N_4241,N_4149,N_4105);
or U4242 (N_4242,N_4081,N_4086);
or U4243 (N_4243,N_4095,N_4165);
and U4244 (N_4244,N_4039,N_4112);
nand U4245 (N_4245,N_4043,N_4107);
and U4246 (N_4246,N_4124,N_4080);
nand U4247 (N_4247,N_4115,N_4021);
nor U4248 (N_4248,N_4025,N_4184);
nand U4249 (N_4249,N_4166,N_4192);
and U4250 (N_4250,N_4067,N_4072);
and U4251 (N_4251,N_4028,N_4055);
nand U4252 (N_4252,N_4128,N_4047);
or U4253 (N_4253,N_4053,N_4064);
or U4254 (N_4254,N_4177,N_4150);
nor U4255 (N_4255,N_4121,N_4164);
nor U4256 (N_4256,N_4094,N_4033);
or U4257 (N_4257,N_4130,N_4092);
nand U4258 (N_4258,N_4138,N_4099);
or U4259 (N_4259,N_4009,N_4050);
nor U4260 (N_4260,N_4127,N_4102);
nand U4261 (N_4261,N_4175,N_4010);
or U4262 (N_4262,N_4007,N_4026);
or U4263 (N_4263,N_4155,N_4186);
nand U4264 (N_4264,N_4059,N_4125);
nand U4265 (N_4265,N_4162,N_4042);
nor U4266 (N_4266,N_4013,N_4084);
or U4267 (N_4267,N_4119,N_4134);
nor U4268 (N_4268,N_4030,N_4163);
nor U4269 (N_4269,N_4195,N_4114);
and U4270 (N_4270,N_4188,N_4196);
or U4271 (N_4271,N_4189,N_4093);
and U4272 (N_4272,N_4082,N_4022);
nor U4273 (N_4273,N_4070,N_4191);
nor U4274 (N_4274,N_4000,N_4016);
or U4275 (N_4275,N_4057,N_4062);
nand U4276 (N_4276,N_4049,N_4079);
and U4277 (N_4277,N_4032,N_4034);
nor U4278 (N_4278,N_4147,N_4154);
nand U4279 (N_4279,N_4133,N_4075);
and U4280 (N_4280,N_4046,N_4152);
or U4281 (N_4281,N_4141,N_4048);
and U4282 (N_4282,N_4108,N_4018);
nor U4283 (N_4283,N_4052,N_4182);
nand U4284 (N_4284,N_4024,N_4109);
or U4285 (N_4285,N_4116,N_4060);
or U4286 (N_4286,N_4065,N_4174);
nor U4287 (N_4287,N_4197,N_4137);
or U4288 (N_4288,N_4100,N_4069);
nand U4289 (N_4289,N_4179,N_4104);
and U4290 (N_4290,N_4172,N_4088);
and U4291 (N_4291,N_4040,N_4096);
nor U4292 (N_4292,N_4167,N_4176);
xor U4293 (N_4293,N_4019,N_4122);
nand U4294 (N_4294,N_4038,N_4002);
nor U4295 (N_4295,N_4181,N_4158);
nand U4296 (N_4296,N_4054,N_4187);
nand U4297 (N_4297,N_4173,N_4005);
and U4298 (N_4298,N_4058,N_4037);
nand U4299 (N_4299,N_4183,N_4014);
or U4300 (N_4300,N_4153,N_4131);
nor U4301 (N_4301,N_4009,N_4102);
nand U4302 (N_4302,N_4137,N_4013);
or U4303 (N_4303,N_4104,N_4007);
and U4304 (N_4304,N_4038,N_4022);
xnor U4305 (N_4305,N_4113,N_4035);
and U4306 (N_4306,N_4158,N_4118);
nor U4307 (N_4307,N_4035,N_4064);
xor U4308 (N_4308,N_4091,N_4022);
or U4309 (N_4309,N_4063,N_4047);
xor U4310 (N_4310,N_4019,N_4173);
nor U4311 (N_4311,N_4173,N_4110);
nand U4312 (N_4312,N_4016,N_4023);
nand U4313 (N_4313,N_4018,N_4045);
nand U4314 (N_4314,N_4111,N_4184);
or U4315 (N_4315,N_4115,N_4071);
or U4316 (N_4316,N_4041,N_4115);
nor U4317 (N_4317,N_4145,N_4182);
and U4318 (N_4318,N_4003,N_4156);
nand U4319 (N_4319,N_4037,N_4014);
nor U4320 (N_4320,N_4125,N_4137);
or U4321 (N_4321,N_4122,N_4027);
nand U4322 (N_4322,N_4110,N_4062);
nand U4323 (N_4323,N_4023,N_4093);
or U4324 (N_4324,N_4035,N_4045);
or U4325 (N_4325,N_4114,N_4012);
nand U4326 (N_4326,N_4088,N_4170);
nand U4327 (N_4327,N_4163,N_4197);
nor U4328 (N_4328,N_4089,N_4194);
nand U4329 (N_4329,N_4066,N_4148);
or U4330 (N_4330,N_4124,N_4119);
and U4331 (N_4331,N_4197,N_4080);
or U4332 (N_4332,N_4023,N_4078);
nand U4333 (N_4333,N_4198,N_4115);
nand U4334 (N_4334,N_4175,N_4143);
nand U4335 (N_4335,N_4048,N_4062);
nor U4336 (N_4336,N_4122,N_4099);
xnor U4337 (N_4337,N_4082,N_4061);
or U4338 (N_4338,N_4028,N_4125);
nand U4339 (N_4339,N_4043,N_4127);
nor U4340 (N_4340,N_4029,N_4161);
nand U4341 (N_4341,N_4102,N_4027);
and U4342 (N_4342,N_4037,N_4125);
nor U4343 (N_4343,N_4071,N_4179);
nand U4344 (N_4344,N_4165,N_4198);
nor U4345 (N_4345,N_4041,N_4158);
and U4346 (N_4346,N_4054,N_4016);
xor U4347 (N_4347,N_4051,N_4028);
nand U4348 (N_4348,N_4075,N_4033);
nor U4349 (N_4349,N_4008,N_4116);
or U4350 (N_4350,N_4166,N_4011);
and U4351 (N_4351,N_4191,N_4153);
or U4352 (N_4352,N_4157,N_4086);
nand U4353 (N_4353,N_4197,N_4068);
and U4354 (N_4354,N_4049,N_4074);
or U4355 (N_4355,N_4066,N_4045);
nand U4356 (N_4356,N_4155,N_4027);
or U4357 (N_4357,N_4101,N_4026);
nor U4358 (N_4358,N_4132,N_4111);
nor U4359 (N_4359,N_4167,N_4026);
and U4360 (N_4360,N_4099,N_4013);
and U4361 (N_4361,N_4151,N_4197);
nand U4362 (N_4362,N_4165,N_4195);
nor U4363 (N_4363,N_4133,N_4080);
and U4364 (N_4364,N_4027,N_4012);
and U4365 (N_4365,N_4049,N_4141);
nand U4366 (N_4366,N_4198,N_4061);
nand U4367 (N_4367,N_4181,N_4045);
or U4368 (N_4368,N_4080,N_4081);
nor U4369 (N_4369,N_4024,N_4019);
nand U4370 (N_4370,N_4092,N_4180);
nor U4371 (N_4371,N_4102,N_4018);
nand U4372 (N_4372,N_4079,N_4095);
nor U4373 (N_4373,N_4175,N_4098);
nand U4374 (N_4374,N_4054,N_4156);
or U4375 (N_4375,N_4033,N_4001);
nor U4376 (N_4376,N_4191,N_4170);
or U4377 (N_4377,N_4110,N_4052);
and U4378 (N_4378,N_4073,N_4188);
and U4379 (N_4379,N_4158,N_4156);
or U4380 (N_4380,N_4026,N_4131);
and U4381 (N_4381,N_4189,N_4039);
or U4382 (N_4382,N_4158,N_4128);
nand U4383 (N_4383,N_4109,N_4116);
or U4384 (N_4384,N_4167,N_4178);
and U4385 (N_4385,N_4187,N_4140);
nor U4386 (N_4386,N_4151,N_4044);
and U4387 (N_4387,N_4166,N_4125);
or U4388 (N_4388,N_4009,N_4144);
or U4389 (N_4389,N_4036,N_4038);
nor U4390 (N_4390,N_4033,N_4092);
or U4391 (N_4391,N_4167,N_4195);
and U4392 (N_4392,N_4038,N_4047);
xor U4393 (N_4393,N_4011,N_4104);
or U4394 (N_4394,N_4096,N_4184);
and U4395 (N_4395,N_4139,N_4147);
nand U4396 (N_4396,N_4148,N_4020);
xor U4397 (N_4397,N_4103,N_4034);
or U4398 (N_4398,N_4013,N_4086);
nor U4399 (N_4399,N_4182,N_4016);
nand U4400 (N_4400,N_4242,N_4358);
nor U4401 (N_4401,N_4300,N_4389);
and U4402 (N_4402,N_4210,N_4265);
nand U4403 (N_4403,N_4287,N_4267);
nor U4404 (N_4404,N_4316,N_4248);
and U4405 (N_4405,N_4335,N_4288);
nor U4406 (N_4406,N_4253,N_4392);
nor U4407 (N_4407,N_4268,N_4315);
and U4408 (N_4408,N_4246,N_4299);
and U4409 (N_4409,N_4282,N_4213);
nand U4410 (N_4410,N_4396,N_4276);
and U4411 (N_4411,N_4226,N_4269);
nor U4412 (N_4412,N_4245,N_4214);
or U4413 (N_4413,N_4314,N_4381);
and U4414 (N_4414,N_4223,N_4355);
or U4415 (N_4415,N_4377,N_4260);
or U4416 (N_4416,N_4391,N_4339);
and U4417 (N_4417,N_4313,N_4376);
or U4418 (N_4418,N_4394,N_4329);
or U4419 (N_4419,N_4207,N_4380);
nand U4420 (N_4420,N_4322,N_4304);
and U4421 (N_4421,N_4349,N_4218);
or U4422 (N_4422,N_4326,N_4307);
or U4423 (N_4423,N_4310,N_4221);
nor U4424 (N_4424,N_4270,N_4222);
nor U4425 (N_4425,N_4318,N_4227);
and U4426 (N_4426,N_4364,N_4371);
and U4427 (N_4427,N_4366,N_4343);
nor U4428 (N_4428,N_4271,N_4284);
or U4429 (N_4429,N_4258,N_4395);
or U4430 (N_4430,N_4306,N_4361);
nor U4431 (N_4431,N_4212,N_4348);
nand U4432 (N_4432,N_4219,N_4387);
or U4433 (N_4433,N_4390,N_4312);
nor U4434 (N_4434,N_4235,N_4263);
nor U4435 (N_4435,N_4200,N_4372);
nor U4436 (N_4436,N_4294,N_4256);
and U4437 (N_4437,N_4374,N_4243);
nand U4438 (N_4438,N_4388,N_4290);
and U4439 (N_4439,N_4386,N_4296);
and U4440 (N_4440,N_4398,N_4217);
nand U4441 (N_4441,N_4231,N_4337);
nor U4442 (N_4442,N_4251,N_4280);
and U4443 (N_4443,N_4375,N_4297);
or U4444 (N_4444,N_4399,N_4345);
and U4445 (N_4445,N_4356,N_4239);
nand U4446 (N_4446,N_4341,N_4277);
or U4447 (N_4447,N_4274,N_4334);
and U4448 (N_4448,N_4309,N_4354);
nor U4449 (N_4449,N_4308,N_4359);
nand U4450 (N_4450,N_4321,N_4261);
nor U4451 (N_4451,N_4220,N_4273);
nand U4452 (N_4452,N_4292,N_4232);
nor U4453 (N_4453,N_4230,N_4379);
and U4454 (N_4454,N_4238,N_4209);
or U4455 (N_4455,N_4216,N_4266);
xor U4456 (N_4456,N_4254,N_4360);
or U4457 (N_4457,N_4211,N_4249);
nand U4458 (N_4458,N_4302,N_4208);
nand U4459 (N_4459,N_4281,N_4373);
or U4460 (N_4460,N_4205,N_4275);
or U4461 (N_4461,N_4336,N_4224);
and U4462 (N_4462,N_4206,N_4264);
or U4463 (N_4463,N_4252,N_4332);
nand U4464 (N_4464,N_4384,N_4283);
nor U4465 (N_4465,N_4262,N_4383);
nor U4466 (N_4466,N_4225,N_4240);
and U4467 (N_4467,N_4328,N_4363);
nor U4468 (N_4468,N_4317,N_4344);
nand U4469 (N_4469,N_4385,N_4293);
or U4470 (N_4470,N_4201,N_4234);
and U4471 (N_4471,N_4320,N_4286);
and U4472 (N_4472,N_4357,N_4368);
nand U4473 (N_4473,N_4353,N_4204);
nand U4474 (N_4474,N_4325,N_4303);
nor U4475 (N_4475,N_4393,N_4241);
nor U4476 (N_4476,N_4330,N_4250);
or U4477 (N_4477,N_4347,N_4247);
and U4478 (N_4478,N_4291,N_4203);
nor U4479 (N_4479,N_4331,N_4285);
or U4480 (N_4480,N_4362,N_4229);
and U4481 (N_4481,N_4301,N_4397);
and U4482 (N_4482,N_4279,N_4237);
nand U4483 (N_4483,N_4323,N_4295);
nor U4484 (N_4484,N_4233,N_4327);
and U4485 (N_4485,N_4319,N_4272);
and U4486 (N_4486,N_4338,N_4352);
nor U4487 (N_4487,N_4346,N_4367);
or U4488 (N_4488,N_4350,N_4370);
or U4489 (N_4489,N_4259,N_4382);
nor U4490 (N_4490,N_4228,N_4257);
or U4491 (N_4491,N_4255,N_4340);
or U4492 (N_4492,N_4236,N_4378);
or U4493 (N_4493,N_4365,N_4369);
nand U4494 (N_4494,N_4289,N_4333);
nor U4495 (N_4495,N_4342,N_4351);
and U4496 (N_4496,N_4305,N_4311);
or U4497 (N_4497,N_4324,N_4202);
and U4498 (N_4498,N_4298,N_4215);
and U4499 (N_4499,N_4278,N_4244);
or U4500 (N_4500,N_4387,N_4310);
nand U4501 (N_4501,N_4304,N_4305);
and U4502 (N_4502,N_4237,N_4366);
or U4503 (N_4503,N_4356,N_4338);
nand U4504 (N_4504,N_4345,N_4295);
nand U4505 (N_4505,N_4210,N_4391);
and U4506 (N_4506,N_4213,N_4378);
and U4507 (N_4507,N_4321,N_4332);
nand U4508 (N_4508,N_4389,N_4255);
and U4509 (N_4509,N_4309,N_4380);
nand U4510 (N_4510,N_4380,N_4382);
nor U4511 (N_4511,N_4277,N_4260);
and U4512 (N_4512,N_4220,N_4305);
or U4513 (N_4513,N_4361,N_4255);
nor U4514 (N_4514,N_4353,N_4286);
nor U4515 (N_4515,N_4248,N_4276);
or U4516 (N_4516,N_4321,N_4349);
nor U4517 (N_4517,N_4392,N_4272);
nor U4518 (N_4518,N_4236,N_4362);
or U4519 (N_4519,N_4293,N_4399);
or U4520 (N_4520,N_4375,N_4235);
and U4521 (N_4521,N_4392,N_4274);
or U4522 (N_4522,N_4353,N_4328);
nand U4523 (N_4523,N_4215,N_4284);
nand U4524 (N_4524,N_4372,N_4219);
or U4525 (N_4525,N_4371,N_4266);
nor U4526 (N_4526,N_4244,N_4379);
and U4527 (N_4527,N_4318,N_4379);
nor U4528 (N_4528,N_4394,N_4323);
and U4529 (N_4529,N_4370,N_4295);
and U4530 (N_4530,N_4252,N_4335);
nand U4531 (N_4531,N_4361,N_4246);
nand U4532 (N_4532,N_4336,N_4243);
and U4533 (N_4533,N_4229,N_4297);
nand U4534 (N_4534,N_4375,N_4261);
and U4535 (N_4535,N_4240,N_4235);
nand U4536 (N_4536,N_4369,N_4307);
nand U4537 (N_4537,N_4279,N_4271);
nor U4538 (N_4538,N_4372,N_4327);
and U4539 (N_4539,N_4393,N_4228);
nor U4540 (N_4540,N_4247,N_4358);
nor U4541 (N_4541,N_4355,N_4351);
and U4542 (N_4542,N_4391,N_4324);
and U4543 (N_4543,N_4288,N_4227);
nand U4544 (N_4544,N_4228,N_4213);
or U4545 (N_4545,N_4332,N_4257);
and U4546 (N_4546,N_4316,N_4219);
or U4547 (N_4547,N_4273,N_4354);
and U4548 (N_4548,N_4397,N_4313);
nor U4549 (N_4549,N_4247,N_4319);
and U4550 (N_4550,N_4316,N_4229);
or U4551 (N_4551,N_4336,N_4335);
nand U4552 (N_4552,N_4205,N_4357);
nor U4553 (N_4553,N_4339,N_4301);
nand U4554 (N_4554,N_4328,N_4281);
nand U4555 (N_4555,N_4348,N_4320);
nor U4556 (N_4556,N_4229,N_4334);
and U4557 (N_4557,N_4304,N_4388);
or U4558 (N_4558,N_4329,N_4265);
nand U4559 (N_4559,N_4296,N_4300);
or U4560 (N_4560,N_4347,N_4390);
nor U4561 (N_4561,N_4385,N_4230);
nand U4562 (N_4562,N_4223,N_4370);
nand U4563 (N_4563,N_4379,N_4287);
nand U4564 (N_4564,N_4215,N_4256);
nand U4565 (N_4565,N_4240,N_4304);
nand U4566 (N_4566,N_4365,N_4217);
nor U4567 (N_4567,N_4272,N_4245);
nand U4568 (N_4568,N_4277,N_4374);
nor U4569 (N_4569,N_4349,N_4318);
nor U4570 (N_4570,N_4317,N_4322);
nand U4571 (N_4571,N_4376,N_4348);
nor U4572 (N_4572,N_4393,N_4339);
nor U4573 (N_4573,N_4340,N_4209);
or U4574 (N_4574,N_4222,N_4373);
nor U4575 (N_4575,N_4309,N_4353);
or U4576 (N_4576,N_4204,N_4356);
and U4577 (N_4577,N_4379,N_4259);
or U4578 (N_4578,N_4225,N_4367);
or U4579 (N_4579,N_4284,N_4318);
nor U4580 (N_4580,N_4328,N_4386);
or U4581 (N_4581,N_4250,N_4347);
xnor U4582 (N_4582,N_4334,N_4363);
xnor U4583 (N_4583,N_4345,N_4262);
or U4584 (N_4584,N_4374,N_4337);
and U4585 (N_4585,N_4300,N_4254);
or U4586 (N_4586,N_4270,N_4291);
nor U4587 (N_4587,N_4305,N_4210);
nand U4588 (N_4588,N_4257,N_4325);
and U4589 (N_4589,N_4360,N_4367);
and U4590 (N_4590,N_4304,N_4279);
and U4591 (N_4591,N_4209,N_4293);
and U4592 (N_4592,N_4254,N_4317);
nor U4593 (N_4593,N_4264,N_4335);
nand U4594 (N_4594,N_4326,N_4398);
and U4595 (N_4595,N_4229,N_4318);
and U4596 (N_4596,N_4316,N_4295);
or U4597 (N_4597,N_4369,N_4330);
nand U4598 (N_4598,N_4296,N_4269);
or U4599 (N_4599,N_4245,N_4313);
or U4600 (N_4600,N_4590,N_4511);
or U4601 (N_4601,N_4404,N_4463);
or U4602 (N_4602,N_4556,N_4525);
nor U4603 (N_4603,N_4548,N_4427);
nor U4604 (N_4604,N_4417,N_4588);
and U4605 (N_4605,N_4473,N_4448);
and U4606 (N_4606,N_4421,N_4596);
or U4607 (N_4607,N_4503,N_4526);
nand U4608 (N_4608,N_4595,N_4405);
nor U4609 (N_4609,N_4411,N_4562);
and U4610 (N_4610,N_4521,N_4578);
and U4611 (N_4611,N_4458,N_4514);
or U4612 (N_4612,N_4439,N_4489);
or U4613 (N_4613,N_4500,N_4557);
or U4614 (N_4614,N_4586,N_4579);
nor U4615 (N_4615,N_4583,N_4599);
nand U4616 (N_4616,N_4508,N_4451);
or U4617 (N_4617,N_4453,N_4549);
nand U4618 (N_4618,N_4495,N_4460);
or U4619 (N_4619,N_4573,N_4512);
and U4620 (N_4620,N_4499,N_4510);
nand U4621 (N_4621,N_4485,N_4457);
and U4622 (N_4622,N_4479,N_4401);
nor U4623 (N_4623,N_4542,N_4465);
nor U4624 (N_4624,N_4440,N_4509);
nand U4625 (N_4625,N_4516,N_4428);
xor U4626 (N_4626,N_4493,N_4478);
nand U4627 (N_4627,N_4409,N_4433);
and U4628 (N_4628,N_4425,N_4498);
nor U4629 (N_4629,N_4436,N_4561);
and U4630 (N_4630,N_4407,N_4502);
nand U4631 (N_4631,N_4501,N_4536);
and U4632 (N_4632,N_4545,N_4575);
or U4633 (N_4633,N_4587,N_4515);
and U4634 (N_4634,N_4437,N_4554);
or U4635 (N_4635,N_4480,N_4544);
nand U4636 (N_4636,N_4444,N_4532);
nand U4637 (N_4637,N_4490,N_4581);
and U4638 (N_4638,N_4567,N_4414);
and U4639 (N_4639,N_4402,N_4564);
nand U4640 (N_4640,N_4455,N_4423);
or U4641 (N_4641,N_4543,N_4540);
and U4642 (N_4642,N_4408,N_4442);
nand U4643 (N_4643,N_4412,N_4560);
nand U4644 (N_4644,N_4547,N_4531);
nor U4645 (N_4645,N_4580,N_4566);
nand U4646 (N_4646,N_4406,N_4420);
nand U4647 (N_4647,N_4565,N_4558);
nor U4648 (N_4648,N_4418,N_4534);
nor U4649 (N_4649,N_4528,N_4577);
nand U4650 (N_4650,N_4505,N_4416);
nor U4651 (N_4651,N_4435,N_4584);
xnor U4652 (N_4652,N_4400,N_4593);
or U4653 (N_4653,N_4429,N_4487);
nor U4654 (N_4654,N_4415,N_4486);
nor U4655 (N_4655,N_4546,N_4585);
and U4656 (N_4656,N_4449,N_4483);
or U4657 (N_4657,N_4452,N_4431);
nand U4658 (N_4658,N_4441,N_4563);
or U4659 (N_4659,N_4506,N_4422);
or U4660 (N_4660,N_4475,N_4494);
or U4661 (N_4661,N_4555,N_4527);
and U4662 (N_4662,N_4469,N_4426);
or U4663 (N_4663,N_4459,N_4598);
nor U4664 (N_4664,N_4434,N_4445);
or U4665 (N_4665,N_4492,N_4535);
nand U4666 (N_4666,N_4552,N_4504);
nor U4667 (N_4667,N_4488,N_4438);
nor U4668 (N_4668,N_4550,N_4574);
nor U4669 (N_4669,N_4530,N_4582);
nor U4670 (N_4670,N_4589,N_4523);
and U4671 (N_4671,N_4553,N_4529);
nor U4672 (N_4672,N_4474,N_4413);
nor U4673 (N_4673,N_4446,N_4592);
and U4674 (N_4674,N_4519,N_4410);
and U4675 (N_4675,N_4539,N_4522);
or U4676 (N_4676,N_4484,N_4569);
or U4677 (N_4677,N_4456,N_4571);
nand U4678 (N_4678,N_4430,N_4559);
or U4679 (N_4679,N_4432,N_4513);
and U4680 (N_4680,N_4461,N_4424);
nor U4681 (N_4681,N_4517,N_4594);
nor U4682 (N_4682,N_4472,N_4470);
or U4683 (N_4683,N_4462,N_4568);
and U4684 (N_4684,N_4597,N_4518);
and U4685 (N_4685,N_4520,N_4467);
nand U4686 (N_4686,N_4454,N_4570);
nor U4687 (N_4687,N_4476,N_4538);
nand U4688 (N_4688,N_4447,N_4551);
nor U4689 (N_4689,N_4591,N_4533);
and U4690 (N_4690,N_4471,N_4464);
xor U4691 (N_4691,N_4524,N_4541);
nor U4692 (N_4692,N_4466,N_4497);
nor U4693 (N_4693,N_4572,N_4576);
and U4694 (N_4694,N_4482,N_4403);
nor U4695 (N_4695,N_4491,N_4496);
nand U4696 (N_4696,N_4468,N_4443);
nor U4697 (N_4697,N_4419,N_4477);
and U4698 (N_4698,N_4481,N_4537);
or U4699 (N_4699,N_4507,N_4450);
nand U4700 (N_4700,N_4462,N_4585);
nor U4701 (N_4701,N_4473,N_4460);
or U4702 (N_4702,N_4476,N_4502);
nor U4703 (N_4703,N_4400,N_4417);
or U4704 (N_4704,N_4557,N_4489);
and U4705 (N_4705,N_4403,N_4483);
or U4706 (N_4706,N_4446,N_4412);
and U4707 (N_4707,N_4434,N_4496);
xor U4708 (N_4708,N_4528,N_4421);
nand U4709 (N_4709,N_4481,N_4496);
or U4710 (N_4710,N_4589,N_4483);
or U4711 (N_4711,N_4521,N_4518);
nor U4712 (N_4712,N_4480,N_4407);
or U4713 (N_4713,N_4571,N_4599);
or U4714 (N_4714,N_4436,N_4415);
and U4715 (N_4715,N_4501,N_4477);
nand U4716 (N_4716,N_4574,N_4543);
or U4717 (N_4717,N_4598,N_4551);
nand U4718 (N_4718,N_4493,N_4590);
and U4719 (N_4719,N_4438,N_4447);
nand U4720 (N_4720,N_4497,N_4495);
nor U4721 (N_4721,N_4576,N_4548);
and U4722 (N_4722,N_4576,N_4411);
or U4723 (N_4723,N_4450,N_4562);
nand U4724 (N_4724,N_4555,N_4494);
and U4725 (N_4725,N_4502,N_4411);
xor U4726 (N_4726,N_4428,N_4574);
or U4727 (N_4727,N_4522,N_4524);
or U4728 (N_4728,N_4454,N_4509);
or U4729 (N_4729,N_4416,N_4419);
or U4730 (N_4730,N_4553,N_4537);
nand U4731 (N_4731,N_4433,N_4526);
nor U4732 (N_4732,N_4448,N_4475);
or U4733 (N_4733,N_4401,N_4483);
nand U4734 (N_4734,N_4586,N_4501);
and U4735 (N_4735,N_4468,N_4598);
nor U4736 (N_4736,N_4536,N_4517);
and U4737 (N_4737,N_4576,N_4527);
nand U4738 (N_4738,N_4423,N_4446);
nor U4739 (N_4739,N_4522,N_4480);
or U4740 (N_4740,N_4432,N_4487);
nor U4741 (N_4741,N_4421,N_4590);
and U4742 (N_4742,N_4423,N_4565);
and U4743 (N_4743,N_4425,N_4512);
and U4744 (N_4744,N_4435,N_4595);
and U4745 (N_4745,N_4580,N_4530);
nor U4746 (N_4746,N_4543,N_4456);
nor U4747 (N_4747,N_4584,N_4547);
and U4748 (N_4748,N_4593,N_4557);
and U4749 (N_4749,N_4559,N_4549);
nand U4750 (N_4750,N_4542,N_4406);
nand U4751 (N_4751,N_4450,N_4463);
xor U4752 (N_4752,N_4541,N_4530);
or U4753 (N_4753,N_4440,N_4521);
and U4754 (N_4754,N_4444,N_4415);
nand U4755 (N_4755,N_4521,N_4432);
and U4756 (N_4756,N_4553,N_4570);
nand U4757 (N_4757,N_4508,N_4403);
and U4758 (N_4758,N_4468,N_4461);
nor U4759 (N_4759,N_4455,N_4596);
nor U4760 (N_4760,N_4401,N_4579);
and U4761 (N_4761,N_4506,N_4442);
xnor U4762 (N_4762,N_4479,N_4516);
or U4763 (N_4763,N_4547,N_4554);
nand U4764 (N_4764,N_4500,N_4445);
nor U4765 (N_4765,N_4494,N_4426);
nand U4766 (N_4766,N_4583,N_4448);
or U4767 (N_4767,N_4553,N_4500);
nand U4768 (N_4768,N_4586,N_4521);
nor U4769 (N_4769,N_4591,N_4458);
or U4770 (N_4770,N_4560,N_4534);
and U4771 (N_4771,N_4458,N_4568);
or U4772 (N_4772,N_4428,N_4532);
and U4773 (N_4773,N_4508,N_4562);
nor U4774 (N_4774,N_4542,N_4565);
nor U4775 (N_4775,N_4487,N_4439);
nand U4776 (N_4776,N_4526,N_4427);
nand U4777 (N_4777,N_4459,N_4435);
nand U4778 (N_4778,N_4544,N_4448);
nand U4779 (N_4779,N_4409,N_4460);
or U4780 (N_4780,N_4514,N_4534);
xor U4781 (N_4781,N_4550,N_4524);
nand U4782 (N_4782,N_4452,N_4522);
or U4783 (N_4783,N_4533,N_4569);
or U4784 (N_4784,N_4546,N_4540);
nand U4785 (N_4785,N_4518,N_4472);
nor U4786 (N_4786,N_4471,N_4493);
and U4787 (N_4787,N_4578,N_4454);
and U4788 (N_4788,N_4588,N_4589);
nor U4789 (N_4789,N_4429,N_4518);
nand U4790 (N_4790,N_4401,N_4415);
or U4791 (N_4791,N_4412,N_4468);
or U4792 (N_4792,N_4553,N_4556);
nand U4793 (N_4793,N_4462,N_4407);
and U4794 (N_4794,N_4538,N_4553);
nand U4795 (N_4795,N_4414,N_4416);
and U4796 (N_4796,N_4486,N_4406);
nand U4797 (N_4797,N_4584,N_4482);
nand U4798 (N_4798,N_4464,N_4477);
and U4799 (N_4799,N_4410,N_4545);
or U4800 (N_4800,N_4669,N_4787);
nor U4801 (N_4801,N_4663,N_4629);
or U4802 (N_4802,N_4735,N_4795);
or U4803 (N_4803,N_4677,N_4727);
nor U4804 (N_4804,N_4765,N_4699);
or U4805 (N_4805,N_4732,N_4611);
nand U4806 (N_4806,N_4722,N_4682);
nor U4807 (N_4807,N_4644,N_4734);
and U4808 (N_4808,N_4675,N_4607);
and U4809 (N_4809,N_4604,N_4637);
nor U4810 (N_4810,N_4763,N_4646);
nor U4811 (N_4811,N_4660,N_4662);
and U4812 (N_4812,N_4724,N_4634);
nand U4813 (N_4813,N_4761,N_4719);
nand U4814 (N_4814,N_4605,N_4784);
nand U4815 (N_4815,N_4626,N_4661);
nand U4816 (N_4816,N_4650,N_4757);
nor U4817 (N_4817,N_4658,N_4756);
nand U4818 (N_4818,N_4630,N_4683);
or U4819 (N_4819,N_4603,N_4745);
nand U4820 (N_4820,N_4743,N_4668);
nor U4821 (N_4821,N_4744,N_4705);
and U4822 (N_4822,N_4747,N_4779);
or U4823 (N_4823,N_4600,N_4681);
nor U4824 (N_4824,N_4615,N_4733);
xnor U4825 (N_4825,N_4748,N_4692);
and U4826 (N_4826,N_4655,N_4642);
or U4827 (N_4827,N_4647,N_4654);
and U4828 (N_4828,N_4753,N_4760);
nor U4829 (N_4829,N_4782,N_4726);
and U4830 (N_4830,N_4664,N_4645);
or U4831 (N_4831,N_4672,N_4752);
and U4832 (N_4832,N_4693,N_4674);
nor U4833 (N_4833,N_4691,N_4689);
nor U4834 (N_4834,N_4742,N_4776);
and U4835 (N_4835,N_4627,N_4746);
or U4836 (N_4836,N_4749,N_4715);
nand U4837 (N_4837,N_4686,N_4631);
nand U4838 (N_4838,N_4792,N_4780);
nor U4839 (N_4839,N_4643,N_4670);
or U4840 (N_4840,N_4641,N_4609);
and U4841 (N_4841,N_4736,N_4778);
or U4842 (N_4842,N_4614,N_4718);
and U4843 (N_4843,N_4720,N_4676);
nand U4844 (N_4844,N_4790,N_4767);
or U4845 (N_4845,N_4771,N_4602);
nor U4846 (N_4846,N_4659,N_4740);
nand U4847 (N_4847,N_4636,N_4608);
nor U4848 (N_4848,N_4758,N_4678);
nand U4849 (N_4849,N_4695,N_4694);
nor U4850 (N_4850,N_4775,N_4680);
nand U4851 (N_4851,N_4794,N_4710);
nand U4852 (N_4852,N_4711,N_4781);
nand U4853 (N_4853,N_4762,N_4737);
nand U4854 (N_4854,N_4638,N_4786);
nor U4855 (N_4855,N_4704,N_4652);
or U4856 (N_4856,N_4738,N_4616);
nor U4857 (N_4857,N_4751,N_4716);
nand U4858 (N_4858,N_4766,N_4684);
or U4859 (N_4859,N_4701,N_4639);
nor U4860 (N_4860,N_4796,N_4725);
nand U4861 (N_4861,N_4700,N_4723);
nand U4862 (N_4862,N_4685,N_4709);
or U4863 (N_4863,N_4708,N_4619);
nor U4864 (N_4864,N_4754,N_4713);
nand U4865 (N_4865,N_4657,N_4785);
or U4866 (N_4866,N_4791,N_4799);
or U4867 (N_4867,N_4730,N_4640);
nor U4868 (N_4868,N_4741,N_4798);
nor U4869 (N_4869,N_4728,N_4688);
nor U4870 (N_4870,N_4653,N_4618);
nor U4871 (N_4871,N_4632,N_4617);
nor U4872 (N_4872,N_4690,N_4625);
nor U4873 (N_4873,N_4750,N_4755);
nand U4874 (N_4874,N_4773,N_4696);
and U4875 (N_4875,N_4777,N_4712);
nor U4876 (N_4876,N_4612,N_4628);
nor U4877 (N_4877,N_4721,N_4624);
nor U4878 (N_4878,N_4703,N_4622);
or U4879 (N_4879,N_4679,N_4601);
and U4880 (N_4880,N_4739,N_4613);
nand U4881 (N_4881,N_4633,N_4729);
and U4882 (N_4882,N_4623,N_4687);
nand U4883 (N_4883,N_4648,N_4772);
nor U4884 (N_4884,N_4768,N_4635);
and U4885 (N_4885,N_4774,N_4665);
and U4886 (N_4886,N_4783,N_4789);
nand U4887 (N_4887,N_4671,N_4606);
nor U4888 (N_4888,N_4731,N_4649);
nor U4889 (N_4889,N_4797,N_4656);
or U4890 (N_4890,N_4793,N_4717);
nand U4891 (N_4891,N_4620,N_4764);
xor U4892 (N_4892,N_4702,N_4667);
and U4893 (N_4893,N_4770,N_4673);
or U4894 (N_4894,N_4759,N_4714);
and U4895 (N_4895,N_4788,N_4666);
nand U4896 (N_4896,N_4621,N_4697);
or U4897 (N_4897,N_4769,N_4707);
and U4898 (N_4898,N_4698,N_4706);
and U4899 (N_4899,N_4651,N_4610);
and U4900 (N_4900,N_4647,N_4643);
or U4901 (N_4901,N_4607,N_4773);
and U4902 (N_4902,N_4747,N_4660);
nor U4903 (N_4903,N_4604,N_4718);
nand U4904 (N_4904,N_4627,N_4721);
and U4905 (N_4905,N_4630,N_4757);
xnor U4906 (N_4906,N_4740,N_4728);
or U4907 (N_4907,N_4675,N_4657);
nand U4908 (N_4908,N_4790,N_4660);
nand U4909 (N_4909,N_4694,N_4790);
nor U4910 (N_4910,N_4611,N_4749);
nand U4911 (N_4911,N_4614,N_4603);
or U4912 (N_4912,N_4616,N_4667);
or U4913 (N_4913,N_4703,N_4705);
nand U4914 (N_4914,N_4639,N_4685);
and U4915 (N_4915,N_4605,N_4715);
nand U4916 (N_4916,N_4775,N_4700);
nand U4917 (N_4917,N_4725,N_4615);
or U4918 (N_4918,N_4653,N_4670);
and U4919 (N_4919,N_4691,N_4708);
nand U4920 (N_4920,N_4689,N_4734);
or U4921 (N_4921,N_4673,N_4736);
and U4922 (N_4922,N_4765,N_4774);
nand U4923 (N_4923,N_4649,N_4656);
nand U4924 (N_4924,N_4648,N_4627);
xnor U4925 (N_4925,N_4767,N_4740);
xor U4926 (N_4926,N_4791,N_4610);
or U4927 (N_4927,N_4723,N_4603);
and U4928 (N_4928,N_4766,N_4709);
or U4929 (N_4929,N_4611,N_4793);
and U4930 (N_4930,N_4605,N_4799);
nand U4931 (N_4931,N_4651,N_4767);
nor U4932 (N_4932,N_4778,N_4644);
nor U4933 (N_4933,N_4628,N_4672);
nand U4934 (N_4934,N_4794,N_4729);
nor U4935 (N_4935,N_4746,N_4762);
or U4936 (N_4936,N_4760,N_4610);
nor U4937 (N_4937,N_4652,N_4622);
nor U4938 (N_4938,N_4637,N_4628);
or U4939 (N_4939,N_4720,N_4729);
nand U4940 (N_4940,N_4691,N_4633);
nand U4941 (N_4941,N_4656,N_4720);
nand U4942 (N_4942,N_4716,N_4761);
or U4943 (N_4943,N_4640,N_4665);
nor U4944 (N_4944,N_4683,N_4603);
or U4945 (N_4945,N_4730,N_4764);
or U4946 (N_4946,N_4644,N_4614);
and U4947 (N_4947,N_4694,N_4604);
nor U4948 (N_4948,N_4642,N_4613);
nand U4949 (N_4949,N_4731,N_4624);
and U4950 (N_4950,N_4780,N_4634);
nor U4951 (N_4951,N_4772,N_4669);
nor U4952 (N_4952,N_4779,N_4611);
nand U4953 (N_4953,N_4692,N_4721);
nor U4954 (N_4954,N_4678,N_4748);
or U4955 (N_4955,N_4617,N_4724);
nand U4956 (N_4956,N_4681,N_4724);
or U4957 (N_4957,N_4792,N_4672);
nor U4958 (N_4958,N_4671,N_4786);
nor U4959 (N_4959,N_4680,N_4748);
or U4960 (N_4960,N_4755,N_4668);
nor U4961 (N_4961,N_4793,N_4678);
nor U4962 (N_4962,N_4716,N_4798);
nor U4963 (N_4963,N_4756,N_4729);
or U4964 (N_4964,N_4651,N_4604);
and U4965 (N_4965,N_4610,N_4775);
and U4966 (N_4966,N_4695,N_4735);
and U4967 (N_4967,N_4630,N_4734);
or U4968 (N_4968,N_4681,N_4750);
nor U4969 (N_4969,N_4706,N_4797);
or U4970 (N_4970,N_4622,N_4662);
and U4971 (N_4971,N_4796,N_4607);
nand U4972 (N_4972,N_4777,N_4747);
nand U4973 (N_4973,N_4639,N_4715);
nor U4974 (N_4974,N_4618,N_4718);
nand U4975 (N_4975,N_4774,N_4729);
and U4976 (N_4976,N_4711,N_4670);
or U4977 (N_4977,N_4705,N_4719);
and U4978 (N_4978,N_4773,N_4608);
nand U4979 (N_4979,N_4746,N_4660);
nand U4980 (N_4980,N_4743,N_4628);
and U4981 (N_4981,N_4738,N_4799);
nand U4982 (N_4982,N_4643,N_4794);
and U4983 (N_4983,N_4702,N_4766);
nor U4984 (N_4984,N_4754,N_4735);
and U4985 (N_4985,N_4739,N_4687);
and U4986 (N_4986,N_4785,N_4755);
or U4987 (N_4987,N_4681,N_4735);
nand U4988 (N_4988,N_4752,N_4739);
nor U4989 (N_4989,N_4777,N_4682);
or U4990 (N_4990,N_4631,N_4627);
and U4991 (N_4991,N_4659,N_4750);
xnor U4992 (N_4992,N_4745,N_4733);
nand U4993 (N_4993,N_4676,N_4723);
and U4994 (N_4994,N_4677,N_4651);
and U4995 (N_4995,N_4746,N_4681);
nor U4996 (N_4996,N_4700,N_4688);
or U4997 (N_4997,N_4764,N_4777);
and U4998 (N_4998,N_4783,N_4674);
and U4999 (N_4999,N_4694,N_4672);
and UO_0 (O_0,N_4979,N_4921);
and UO_1 (O_1,N_4966,N_4851);
nand UO_2 (O_2,N_4812,N_4822);
nor UO_3 (O_3,N_4916,N_4882);
and UO_4 (O_4,N_4900,N_4955);
nor UO_5 (O_5,N_4805,N_4821);
nor UO_6 (O_6,N_4904,N_4907);
xor UO_7 (O_7,N_4923,N_4930);
nand UO_8 (O_8,N_4967,N_4952);
and UO_9 (O_9,N_4880,N_4884);
nand UO_10 (O_10,N_4852,N_4867);
and UO_11 (O_11,N_4908,N_4943);
and UO_12 (O_12,N_4847,N_4849);
or UO_13 (O_13,N_4948,N_4811);
nand UO_14 (O_14,N_4878,N_4906);
or UO_15 (O_15,N_4868,N_4942);
nor UO_16 (O_16,N_4848,N_4935);
nor UO_17 (O_17,N_4996,N_4910);
and UO_18 (O_18,N_4919,N_4912);
nor UO_19 (O_19,N_4991,N_4890);
and UO_20 (O_20,N_4939,N_4972);
nand UO_21 (O_21,N_4808,N_4889);
nand UO_22 (O_22,N_4950,N_4938);
or UO_23 (O_23,N_4850,N_4839);
xnor UO_24 (O_24,N_4976,N_4920);
and UO_25 (O_25,N_4817,N_4940);
or UO_26 (O_26,N_4818,N_4947);
nand UO_27 (O_27,N_4989,N_4885);
nor UO_28 (O_28,N_4854,N_4892);
or UO_29 (O_29,N_4974,N_4862);
nor UO_30 (O_30,N_4816,N_4977);
or UO_31 (O_31,N_4896,N_4980);
or UO_32 (O_32,N_4872,N_4963);
and UO_33 (O_33,N_4925,N_4936);
nand UO_34 (O_34,N_4829,N_4926);
or UO_35 (O_35,N_4866,N_4843);
or UO_36 (O_36,N_4951,N_4834);
or UO_37 (O_37,N_4835,N_4914);
nor UO_38 (O_38,N_4993,N_4901);
nor UO_39 (O_39,N_4982,N_4917);
or UO_40 (O_40,N_4937,N_4870);
or UO_41 (O_41,N_4842,N_4804);
or UO_42 (O_42,N_4858,N_4807);
nor UO_43 (O_43,N_4864,N_4911);
and UO_44 (O_44,N_4819,N_4975);
nand UO_45 (O_45,N_4954,N_4863);
nor UO_46 (O_46,N_4823,N_4944);
or UO_47 (O_47,N_4814,N_4869);
and UO_48 (O_48,N_4856,N_4928);
nor UO_49 (O_49,N_4957,N_4845);
nand UO_50 (O_50,N_4932,N_4992);
and UO_51 (O_51,N_4853,N_4860);
and UO_52 (O_52,N_4883,N_4994);
and UO_53 (O_53,N_4987,N_4960);
and UO_54 (O_54,N_4855,N_4833);
and UO_55 (O_55,N_4832,N_4809);
nor UO_56 (O_56,N_4813,N_4873);
and UO_57 (O_57,N_4981,N_4897);
nor UO_58 (O_58,N_4985,N_4838);
or UO_59 (O_59,N_4801,N_4941);
nor UO_60 (O_60,N_4828,N_4934);
nand UO_61 (O_61,N_4995,N_4964);
or UO_62 (O_62,N_4998,N_4978);
or UO_63 (O_63,N_4879,N_4830);
or UO_64 (O_64,N_4893,N_4961);
or UO_65 (O_65,N_4837,N_4962);
or UO_66 (O_66,N_4810,N_4969);
nor UO_67 (O_67,N_4931,N_4905);
and UO_68 (O_68,N_4970,N_4999);
or UO_69 (O_69,N_4800,N_4899);
nand UO_70 (O_70,N_4913,N_4841);
and UO_71 (O_71,N_4806,N_4857);
nand UO_72 (O_72,N_4895,N_4988);
or UO_73 (O_73,N_4874,N_4953);
and UO_74 (O_74,N_4903,N_4918);
and UO_75 (O_75,N_4997,N_4902);
xor UO_76 (O_76,N_4949,N_4881);
nand UO_77 (O_77,N_4803,N_4827);
or UO_78 (O_78,N_4887,N_4861);
nor UO_79 (O_79,N_4965,N_4836);
and UO_80 (O_80,N_4859,N_4891);
nand UO_81 (O_81,N_4933,N_4915);
xnor UO_82 (O_82,N_4871,N_4824);
or UO_83 (O_83,N_4973,N_4894);
or UO_84 (O_84,N_4984,N_4826);
and UO_85 (O_85,N_4958,N_4986);
nand UO_86 (O_86,N_4815,N_4971);
and UO_87 (O_87,N_4831,N_4922);
nand UO_88 (O_88,N_4945,N_4825);
nor UO_89 (O_89,N_4877,N_4865);
and UO_90 (O_90,N_4886,N_4820);
and UO_91 (O_91,N_4875,N_4844);
and UO_92 (O_92,N_4898,N_4802);
and UO_93 (O_93,N_4990,N_4909);
nand UO_94 (O_94,N_4983,N_4888);
nor UO_95 (O_95,N_4929,N_4959);
and UO_96 (O_96,N_4968,N_4927);
and UO_97 (O_97,N_4840,N_4876);
or UO_98 (O_98,N_4956,N_4846);
or UO_99 (O_99,N_4924,N_4946);
and UO_100 (O_100,N_4949,N_4942);
nor UO_101 (O_101,N_4866,N_4886);
nor UO_102 (O_102,N_4971,N_4827);
or UO_103 (O_103,N_4823,N_4982);
nor UO_104 (O_104,N_4878,N_4945);
or UO_105 (O_105,N_4918,N_4901);
nor UO_106 (O_106,N_4929,N_4817);
nand UO_107 (O_107,N_4957,N_4932);
nor UO_108 (O_108,N_4960,N_4876);
and UO_109 (O_109,N_4977,N_4827);
and UO_110 (O_110,N_4841,N_4977);
nand UO_111 (O_111,N_4953,N_4912);
or UO_112 (O_112,N_4961,N_4910);
xnor UO_113 (O_113,N_4973,N_4833);
and UO_114 (O_114,N_4888,N_4942);
and UO_115 (O_115,N_4893,N_4850);
nor UO_116 (O_116,N_4939,N_4877);
or UO_117 (O_117,N_4870,N_4888);
nand UO_118 (O_118,N_4973,N_4852);
or UO_119 (O_119,N_4917,N_4814);
nand UO_120 (O_120,N_4858,N_4854);
nand UO_121 (O_121,N_4897,N_4820);
nor UO_122 (O_122,N_4989,N_4987);
or UO_123 (O_123,N_4939,N_4840);
xnor UO_124 (O_124,N_4916,N_4949);
nor UO_125 (O_125,N_4866,N_4925);
nor UO_126 (O_126,N_4806,N_4931);
nor UO_127 (O_127,N_4819,N_4853);
or UO_128 (O_128,N_4843,N_4954);
and UO_129 (O_129,N_4917,N_4975);
nor UO_130 (O_130,N_4864,N_4810);
and UO_131 (O_131,N_4884,N_4830);
nand UO_132 (O_132,N_4938,N_4876);
or UO_133 (O_133,N_4824,N_4825);
or UO_134 (O_134,N_4976,N_4955);
or UO_135 (O_135,N_4827,N_4979);
and UO_136 (O_136,N_4836,N_4980);
nor UO_137 (O_137,N_4833,N_4853);
nor UO_138 (O_138,N_4866,N_4819);
and UO_139 (O_139,N_4803,N_4937);
nor UO_140 (O_140,N_4905,N_4985);
nand UO_141 (O_141,N_4960,N_4975);
or UO_142 (O_142,N_4976,N_4882);
or UO_143 (O_143,N_4886,N_4883);
nor UO_144 (O_144,N_4974,N_4806);
nand UO_145 (O_145,N_4865,N_4998);
and UO_146 (O_146,N_4984,N_4893);
or UO_147 (O_147,N_4954,N_4887);
and UO_148 (O_148,N_4992,N_4951);
nand UO_149 (O_149,N_4835,N_4862);
nor UO_150 (O_150,N_4914,N_4886);
nor UO_151 (O_151,N_4921,N_4934);
and UO_152 (O_152,N_4915,N_4922);
nor UO_153 (O_153,N_4897,N_4994);
nor UO_154 (O_154,N_4816,N_4953);
and UO_155 (O_155,N_4961,N_4952);
nor UO_156 (O_156,N_4898,N_4974);
nor UO_157 (O_157,N_4938,N_4942);
nand UO_158 (O_158,N_4820,N_4828);
nand UO_159 (O_159,N_4918,N_4822);
nand UO_160 (O_160,N_4845,N_4854);
and UO_161 (O_161,N_4823,N_4812);
and UO_162 (O_162,N_4854,N_4976);
nand UO_163 (O_163,N_4837,N_4899);
nand UO_164 (O_164,N_4901,N_4804);
and UO_165 (O_165,N_4962,N_4933);
or UO_166 (O_166,N_4947,N_4867);
nand UO_167 (O_167,N_4908,N_4964);
nand UO_168 (O_168,N_4972,N_4969);
nand UO_169 (O_169,N_4939,N_4893);
nand UO_170 (O_170,N_4819,N_4901);
or UO_171 (O_171,N_4832,N_4908);
and UO_172 (O_172,N_4810,N_4954);
nor UO_173 (O_173,N_4810,N_4846);
nand UO_174 (O_174,N_4885,N_4873);
and UO_175 (O_175,N_4992,N_4853);
and UO_176 (O_176,N_4961,N_4860);
or UO_177 (O_177,N_4936,N_4898);
nand UO_178 (O_178,N_4974,N_4988);
nor UO_179 (O_179,N_4998,N_4899);
nor UO_180 (O_180,N_4965,N_4951);
nor UO_181 (O_181,N_4928,N_4895);
or UO_182 (O_182,N_4960,N_4820);
and UO_183 (O_183,N_4817,N_4862);
or UO_184 (O_184,N_4812,N_4887);
or UO_185 (O_185,N_4969,N_4970);
or UO_186 (O_186,N_4896,N_4974);
nor UO_187 (O_187,N_4976,N_4980);
nor UO_188 (O_188,N_4991,N_4962);
nand UO_189 (O_189,N_4900,N_4922);
nor UO_190 (O_190,N_4903,N_4834);
nand UO_191 (O_191,N_4961,N_4821);
nor UO_192 (O_192,N_4873,N_4970);
nor UO_193 (O_193,N_4822,N_4834);
or UO_194 (O_194,N_4923,N_4959);
or UO_195 (O_195,N_4842,N_4926);
and UO_196 (O_196,N_4914,N_4849);
or UO_197 (O_197,N_4874,N_4986);
and UO_198 (O_198,N_4955,N_4865);
or UO_199 (O_199,N_4922,N_4849);
or UO_200 (O_200,N_4969,N_4832);
xnor UO_201 (O_201,N_4903,N_4958);
xor UO_202 (O_202,N_4844,N_4983);
or UO_203 (O_203,N_4978,N_4808);
nand UO_204 (O_204,N_4865,N_4838);
and UO_205 (O_205,N_4854,N_4890);
and UO_206 (O_206,N_4804,N_4853);
and UO_207 (O_207,N_4837,N_4845);
or UO_208 (O_208,N_4938,N_4852);
and UO_209 (O_209,N_4819,N_4856);
nor UO_210 (O_210,N_4888,N_4926);
nor UO_211 (O_211,N_4960,N_4962);
nand UO_212 (O_212,N_4886,N_4958);
or UO_213 (O_213,N_4931,N_4800);
nor UO_214 (O_214,N_4887,N_4808);
and UO_215 (O_215,N_4944,N_4879);
nor UO_216 (O_216,N_4810,N_4901);
and UO_217 (O_217,N_4924,N_4992);
nand UO_218 (O_218,N_4928,N_4964);
nand UO_219 (O_219,N_4930,N_4836);
and UO_220 (O_220,N_4865,N_4947);
nand UO_221 (O_221,N_4971,N_4805);
or UO_222 (O_222,N_4974,N_4866);
or UO_223 (O_223,N_4985,N_4981);
nand UO_224 (O_224,N_4808,N_4882);
nand UO_225 (O_225,N_4988,N_4933);
nand UO_226 (O_226,N_4826,N_4860);
xnor UO_227 (O_227,N_4994,N_4970);
nand UO_228 (O_228,N_4832,N_4883);
nand UO_229 (O_229,N_4994,N_4995);
nand UO_230 (O_230,N_4966,N_4809);
nor UO_231 (O_231,N_4991,N_4995);
nor UO_232 (O_232,N_4927,N_4812);
and UO_233 (O_233,N_4915,N_4902);
nor UO_234 (O_234,N_4854,N_4894);
nor UO_235 (O_235,N_4857,N_4990);
or UO_236 (O_236,N_4828,N_4801);
nor UO_237 (O_237,N_4802,N_4984);
and UO_238 (O_238,N_4851,N_4859);
and UO_239 (O_239,N_4903,N_4971);
nor UO_240 (O_240,N_4819,N_4849);
and UO_241 (O_241,N_4940,N_4937);
nand UO_242 (O_242,N_4941,N_4999);
nand UO_243 (O_243,N_4888,N_4880);
nand UO_244 (O_244,N_4988,N_4812);
nand UO_245 (O_245,N_4959,N_4960);
and UO_246 (O_246,N_4923,N_4855);
nor UO_247 (O_247,N_4874,N_4966);
nor UO_248 (O_248,N_4897,N_4993);
nand UO_249 (O_249,N_4869,N_4885);
or UO_250 (O_250,N_4977,N_4808);
nand UO_251 (O_251,N_4850,N_4988);
nor UO_252 (O_252,N_4861,N_4985);
and UO_253 (O_253,N_4840,N_4801);
or UO_254 (O_254,N_4930,N_4907);
xor UO_255 (O_255,N_4994,N_4968);
and UO_256 (O_256,N_4909,N_4904);
nor UO_257 (O_257,N_4890,N_4905);
nor UO_258 (O_258,N_4993,N_4898);
nor UO_259 (O_259,N_4953,N_4966);
xor UO_260 (O_260,N_4842,N_4800);
nand UO_261 (O_261,N_4875,N_4988);
nand UO_262 (O_262,N_4938,N_4895);
or UO_263 (O_263,N_4832,N_4853);
xnor UO_264 (O_264,N_4810,N_4833);
and UO_265 (O_265,N_4993,N_4980);
or UO_266 (O_266,N_4950,N_4986);
nor UO_267 (O_267,N_4990,N_4902);
or UO_268 (O_268,N_4853,N_4908);
xor UO_269 (O_269,N_4897,N_4900);
and UO_270 (O_270,N_4880,N_4917);
and UO_271 (O_271,N_4989,N_4809);
or UO_272 (O_272,N_4839,N_4801);
nand UO_273 (O_273,N_4821,N_4982);
nand UO_274 (O_274,N_4988,N_4989);
and UO_275 (O_275,N_4810,N_4855);
and UO_276 (O_276,N_4918,N_4965);
or UO_277 (O_277,N_4917,N_4862);
nand UO_278 (O_278,N_4942,N_4987);
and UO_279 (O_279,N_4862,N_4884);
or UO_280 (O_280,N_4831,N_4880);
or UO_281 (O_281,N_4954,N_4809);
nor UO_282 (O_282,N_4836,N_4931);
nor UO_283 (O_283,N_4819,N_4871);
nand UO_284 (O_284,N_4893,N_4922);
and UO_285 (O_285,N_4803,N_4928);
and UO_286 (O_286,N_4941,N_4868);
or UO_287 (O_287,N_4918,N_4885);
or UO_288 (O_288,N_4857,N_4870);
and UO_289 (O_289,N_4800,N_4986);
nor UO_290 (O_290,N_4903,N_4975);
and UO_291 (O_291,N_4941,N_4919);
or UO_292 (O_292,N_4863,N_4884);
and UO_293 (O_293,N_4869,N_4870);
nand UO_294 (O_294,N_4988,N_4805);
nand UO_295 (O_295,N_4871,N_4970);
nor UO_296 (O_296,N_4876,N_4804);
nand UO_297 (O_297,N_4988,N_4900);
and UO_298 (O_298,N_4862,N_4935);
or UO_299 (O_299,N_4873,N_4878);
and UO_300 (O_300,N_4962,N_4834);
or UO_301 (O_301,N_4926,N_4937);
and UO_302 (O_302,N_4983,N_4929);
xnor UO_303 (O_303,N_4971,N_4895);
nand UO_304 (O_304,N_4965,N_4938);
nor UO_305 (O_305,N_4945,N_4974);
nand UO_306 (O_306,N_4887,N_4952);
and UO_307 (O_307,N_4863,N_4966);
nor UO_308 (O_308,N_4893,N_4904);
and UO_309 (O_309,N_4908,N_4884);
nor UO_310 (O_310,N_4944,N_4912);
nand UO_311 (O_311,N_4912,N_4921);
nand UO_312 (O_312,N_4909,N_4846);
and UO_313 (O_313,N_4978,N_4873);
nand UO_314 (O_314,N_4986,N_4862);
nor UO_315 (O_315,N_4835,N_4913);
xnor UO_316 (O_316,N_4965,N_4900);
nor UO_317 (O_317,N_4854,N_4810);
nor UO_318 (O_318,N_4979,N_4887);
and UO_319 (O_319,N_4984,N_4830);
or UO_320 (O_320,N_4816,N_4911);
and UO_321 (O_321,N_4937,N_4850);
nor UO_322 (O_322,N_4974,N_4983);
nand UO_323 (O_323,N_4911,N_4994);
or UO_324 (O_324,N_4879,N_4934);
nor UO_325 (O_325,N_4808,N_4822);
and UO_326 (O_326,N_4880,N_4809);
nor UO_327 (O_327,N_4868,N_4881);
and UO_328 (O_328,N_4904,N_4863);
and UO_329 (O_329,N_4980,N_4995);
nor UO_330 (O_330,N_4954,N_4845);
nor UO_331 (O_331,N_4895,N_4825);
and UO_332 (O_332,N_4848,N_4880);
nor UO_333 (O_333,N_4830,N_4988);
and UO_334 (O_334,N_4932,N_4916);
nor UO_335 (O_335,N_4961,N_4964);
nor UO_336 (O_336,N_4949,N_4911);
nor UO_337 (O_337,N_4870,N_4896);
xnor UO_338 (O_338,N_4905,N_4891);
nand UO_339 (O_339,N_4948,N_4883);
and UO_340 (O_340,N_4963,N_4991);
or UO_341 (O_341,N_4887,N_4888);
and UO_342 (O_342,N_4909,N_4928);
or UO_343 (O_343,N_4999,N_4887);
or UO_344 (O_344,N_4899,N_4881);
and UO_345 (O_345,N_4819,N_4872);
and UO_346 (O_346,N_4867,N_4935);
nand UO_347 (O_347,N_4993,N_4877);
nor UO_348 (O_348,N_4928,N_4910);
nand UO_349 (O_349,N_4868,N_4865);
or UO_350 (O_350,N_4977,N_4843);
nand UO_351 (O_351,N_4876,N_4902);
nor UO_352 (O_352,N_4922,N_4975);
and UO_353 (O_353,N_4907,N_4846);
and UO_354 (O_354,N_4853,N_4813);
nand UO_355 (O_355,N_4828,N_4916);
and UO_356 (O_356,N_4800,N_4948);
nand UO_357 (O_357,N_4826,N_4805);
nand UO_358 (O_358,N_4814,N_4952);
or UO_359 (O_359,N_4884,N_4886);
nand UO_360 (O_360,N_4937,N_4953);
and UO_361 (O_361,N_4811,N_4895);
nand UO_362 (O_362,N_4981,N_4900);
nand UO_363 (O_363,N_4977,N_4833);
nand UO_364 (O_364,N_4908,N_4841);
and UO_365 (O_365,N_4938,N_4906);
and UO_366 (O_366,N_4884,N_4945);
xnor UO_367 (O_367,N_4895,N_4902);
nand UO_368 (O_368,N_4825,N_4817);
and UO_369 (O_369,N_4991,N_4977);
nand UO_370 (O_370,N_4929,N_4979);
nor UO_371 (O_371,N_4954,N_4867);
nand UO_372 (O_372,N_4970,N_4818);
nand UO_373 (O_373,N_4827,N_4853);
nand UO_374 (O_374,N_4873,N_4899);
or UO_375 (O_375,N_4896,N_4963);
or UO_376 (O_376,N_4933,N_4836);
nand UO_377 (O_377,N_4859,N_4955);
nor UO_378 (O_378,N_4874,N_4844);
nand UO_379 (O_379,N_4950,N_4955);
nor UO_380 (O_380,N_4800,N_4984);
nor UO_381 (O_381,N_4832,N_4847);
nor UO_382 (O_382,N_4813,N_4884);
nor UO_383 (O_383,N_4881,N_4810);
nand UO_384 (O_384,N_4990,N_4989);
and UO_385 (O_385,N_4876,N_4945);
nor UO_386 (O_386,N_4916,N_4840);
nand UO_387 (O_387,N_4962,N_4953);
nor UO_388 (O_388,N_4854,N_4939);
nand UO_389 (O_389,N_4874,N_4976);
and UO_390 (O_390,N_4926,N_4802);
or UO_391 (O_391,N_4905,N_4886);
nand UO_392 (O_392,N_4908,N_4879);
and UO_393 (O_393,N_4988,N_4982);
nand UO_394 (O_394,N_4902,N_4894);
and UO_395 (O_395,N_4818,N_4990);
and UO_396 (O_396,N_4822,N_4852);
nand UO_397 (O_397,N_4944,N_4926);
xor UO_398 (O_398,N_4979,N_4811);
and UO_399 (O_399,N_4843,N_4856);
and UO_400 (O_400,N_4910,N_4858);
nor UO_401 (O_401,N_4922,N_4832);
nand UO_402 (O_402,N_4842,N_4878);
and UO_403 (O_403,N_4921,N_4893);
or UO_404 (O_404,N_4954,N_4908);
or UO_405 (O_405,N_4905,N_4910);
and UO_406 (O_406,N_4837,N_4968);
nor UO_407 (O_407,N_4855,N_4841);
or UO_408 (O_408,N_4941,N_4879);
nor UO_409 (O_409,N_4883,N_4810);
or UO_410 (O_410,N_4865,N_4837);
or UO_411 (O_411,N_4894,N_4976);
or UO_412 (O_412,N_4892,N_4999);
nor UO_413 (O_413,N_4839,N_4988);
nor UO_414 (O_414,N_4800,N_4993);
or UO_415 (O_415,N_4967,N_4942);
nor UO_416 (O_416,N_4858,N_4947);
nor UO_417 (O_417,N_4830,N_4820);
and UO_418 (O_418,N_4838,N_4873);
nor UO_419 (O_419,N_4856,N_4858);
nand UO_420 (O_420,N_4866,N_4921);
nor UO_421 (O_421,N_4913,N_4979);
nand UO_422 (O_422,N_4802,N_4983);
nand UO_423 (O_423,N_4962,N_4886);
nor UO_424 (O_424,N_4832,N_4813);
nor UO_425 (O_425,N_4829,N_4910);
or UO_426 (O_426,N_4927,N_4964);
nor UO_427 (O_427,N_4929,N_4890);
or UO_428 (O_428,N_4841,N_4974);
and UO_429 (O_429,N_4824,N_4961);
and UO_430 (O_430,N_4873,N_4938);
nor UO_431 (O_431,N_4960,N_4842);
nand UO_432 (O_432,N_4929,N_4942);
nand UO_433 (O_433,N_4892,N_4960);
nand UO_434 (O_434,N_4907,N_4815);
nor UO_435 (O_435,N_4947,N_4975);
or UO_436 (O_436,N_4803,N_4942);
nand UO_437 (O_437,N_4842,N_4820);
xor UO_438 (O_438,N_4959,N_4926);
nand UO_439 (O_439,N_4934,N_4813);
nand UO_440 (O_440,N_4910,N_4993);
nor UO_441 (O_441,N_4812,N_4984);
and UO_442 (O_442,N_4814,N_4864);
and UO_443 (O_443,N_4837,N_4891);
nand UO_444 (O_444,N_4955,N_4909);
or UO_445 (O_445,N_4900,N_4848);
nor UO_446 (O_446,N_4940,N_4899);
and UO_447 (O_447,N_4905,N_4837);
and UO_448 (O_448,N_4834,N_4976);
nor UO_449 (O_449,N_4835,N_4901);
nor UO_450 (O_450,N_4906,N_4855);
nand UO_451 (O_451,N_4824,N_4968);
or UO_452 (O_452,N_4979,N_4985);
nand UO_453 (O_453,N_4824,N_4866);
and UO_454 (O_454,N_4966,N_4929);
and UO_455 (O_455,N_4951,N_4840);
nor UO_456 (O_456,N_4987,N_4864);
nand UO_457 (O_457,N_4914,N_4945);
nor UO_458 (O_458,N_4921,N_4831);
or UO_459 (O_459,N_4813,N_4886);
and UO_460 (O_460,N_4987,N_4847);
nand UO_461 (O_461,N_4936,N_4917);
or UO_462 (O_462,N_4850,N_4921);
nand UO_463 (O_463,N_4958,N_4997);
nor UO_464 (O_464,N_4949,N_4808);
nand UO_465 (O_465,N_4895,N_4889);
or UO_466 (O_466,N_4966,N_4800);
nor UO_467 (O_467,N_4940,N_4933);
nor UO_468 (O_468,N_4859,N_4882);
nand UO_469 (O_469,N_4824,N_4925);
nor UO_470 (O_470,N_4925,N_4995);
nand UO_471 (O_471,N_4865,N_4885);
nand UO_472 (O_472,N_4893,N_4872);
and UO_473 (O_473,N_4914,N_4959);
or UO_474 (O_474,N_4832,N_4934);
nand UO_475 (O_475,N_4964,N_4832);
nand UO_476 (O_476,N_4980,N_4848);
or UO_477 (O_477,N_4931,N_4855);
nor UO_478 (O_478,N_4873,N_4939);
or UO_479 (O_479,N_4828,N_4927);
or UO_480 (O_480,N_4916,N_4879);
or UO_481 (O_481,N_4909,N_4937);
xor UO_482 (O_482,N_4822,N_4969);
nand UO_483 (O_483,N_4923,N_4921);
nand UO_484 (O_484,N_4977,N_4984);
nor UO_485 (O_485,N_4965,N_4864);
and UO_486 (O_486,N_4995,N_4936);
nor UO_487 (O_487,N_4897,N_4920);
and UO_488 (O_488,N_4838,N_4937);
or UO_489 (O_489,N_4854,N_4885);
or UO_490 (O_490,N_4864,N_4986);
and UO_491 (O_491,N_4853,N_4855);
nor UO_492 (O_492,N_4863,N_4902);
nor UO_493 (O_493,N_4955,N_4957);
nor UO_494 (O_494,N_4817,N_4868);
and UO_495 (O_495,N_4825,N_4813);
nor UO_496 (O_496,N_4974,N_4814);
nand UO_497 (O_497,N_4832,N_4956);
nand UO_498 (O_498,N_4821,N_4994);
or UO_499 (O_499,N_4829,N_4820);
nor UO_500 (O_500,N_4964,N_4920);
nand UO_501 (O_501,N_4866,N_4935);
nand UO_502 (O_502,N_4946,N_4995);
nand UO_503 (O_503,N_4845,N_4849);
nand UO_504 (O_504,N_4952,N_4835);
and UO_505 (O_505,N_4974,N_4836);
nor UO_506 (O_506,N_4993,N_4803);
or UO_507 (O_507,N_4919,N_4840);
or UO_508 (O_508,N_4948,N_4810);
nor UO_509 (O_509,N_4923,N_4883);
nand UO_510 (O_510,N_4826,N_4890);
nor UO_511 (O_511,N_4971,N_4845);
or UO_512 (O_512,N_4989,N_4870);
nor UO_513 (O_513,N_4969,N_4895);
or UO_514 (O_514,N_4961,N_4906);
and UO_515 (O_515,N_4881,N_4848);
or UO_516 (O_516,N_4842,N_4970);
nor UO_517 (O_517,N_4909,N_4878);
nand UO_518 (O_518,N_4924,N_4908);
nor UO_519 (O_519,N_4976,N_4977);
and UO_520 (O_520,N_4884,N_4850);
or UO_521 (O_521,N_4968,N_4967);
nand UO_522 (O_522,N_4997,N_4979);
nand UO_523 (O_523,N_4901,N_4826);
and UO_524 (O_524,N_4824,N_4999);
and UO_525 (O_525,N_4949,N_4876);
nand UO_526 (O_526,N_4803,N_4941);
nand UO_527 (O_527,N_4832,N_4914);
and UO_528 (O_528,N_4913,N_4929);
nand UO_529 (O_529,N_4912,N_4896);
and UO_530 (O_530,N_4808,N_4898);
and UO_531 (O_531,N_4882,N_4969);
or UO_532 (O_532,N_4932,N_4946);
and UO_533 (O_533,N_4901,N_4896);
nor UO_534 (O_534,N_4885,N_4859);
nand UO_535 (O_535,N_4815,N_4809);
or UO_536 (O_536,N_4961,N_4985);
nand UO_537 (O_537,N_4931,N_4960);
nand UO_538 (O_538,N_4958,N_4862);
nor UO_539 (O_539,N_4980,N_4912);
or UO_540 (O_540,N_4828,N_4898);
or UO_541 (O_541,N_4932,N_4833);
and UO_542 (O_542,N_4913,N_4941);
and UO_543 (O_543,N_4940,N_4870);
or UO_544 (O_544,N_4974,N_4959);
nor UO_545 (O_545,N_4942,N_4885);
and UO_546 (O_546,N_4920,N_4992);
and UO_547 (O_547,N_4880,N_4815);
or UO_548 (O_548,N_4925,N_4879);
and UO_549 (O_549,N_4841,N_4920);
nor UO_550 (O_550,N_4928,N_4862);
or UO_551 (O_551,N_4912,N_4887);
or UO_552 (O_552,N_4892,N_4866);
nor UO_553 (O_553,N_4908,N_4968);
nor UO_554 (O_554,N_4910,N_4919);
nand UO_555 (O_555,N_4998,N_4884);
nor UO_556 (O_556,N_4949,N_4910);
nand UO_557 (O_557,N_4834,N_4901);
nor UO_558 (O_558,N_4872,N_4838);
and UO_559 (O_559,N_4918,N_4989);
nand UO_560 (O_560,N_4887,N_4950);
and UO_561 (O_561,N_4972,N_4871);
nand UO_562 (O_562,N_4861,N_4941);
nor UO_563 (O_563,N_4818,N_4957);
nand UO_564 (O_564,N_4940,N_4909);
nor UO_565 (O_565,N_4860,N_4948);
and UO_566 (O_566,N_4920,N_4991);
or UO_567 (O_567,N_4925,N_4867);
nand UO_568 (O_568,N_4938,N_4949);
and UO_569 (O_569,N_4924,N_4942);
and UO_570 (O_570,N_4854,N_4809);
and UO_571 (O_571,N_4986,N_4913);
and UO_572 (O_572,N_4897,N_4810);
and UO_573 (O_573,N_4816,N_4899);
nor UO_574 (O_574,N_4958,N_4831);
or UO_575 (O_575,N_4980,N_4890);
nor UO_576 (O_576,N_4803,N_4904);
nand UO_577 (O_577,N_4911,N_4956);
nand UO_578 (O_578,N_4996,N_4836);
and UO_579 (O_579,N_4985,N_4875);
nand UO_580 (O_580,N_4865,N_4978);
nor UO_581 (O_581,N_4943,N_4910);
or UO_582 (O_582,N_4928,N_4946);
or UO_583 (O_583,N_4845,N_4961);
or UO_584 (O_584,N_4837,N_4939);
or UO_585 (O_585,N_4840,N_4827);
or UO_586 (O_586,N_4890,N_4947);
nand UO_587 (O_587,N_4809,N_4950);
nand UO_588 (O_588,N_4944,N_4960);
and UO_589 (O_589,N_4926,N_4859);
xor UO_590 (O_590,N_4967,N_4851);
and UO_591 (O_591,N_4994,N_4988);
and UO_592 (O_592,N_4825,N_4893);
and UO_593 (O_593,N_4903,N_4934);
or UO_594 (O_594,N_4918,N_4964);
or UO_595 (O_595,N_4880,N_4858);
nor UO_596 (O_596,N_4849,N_4876);
nand UO_597 (O_597,N_4919,N_4870);
nor UO_598 (O_598,N_4918,N_4934);
nand UO_599 (O_599,N_4856,N_4869);
nor UO_600 (O_600,N_4970,N_4952);
nand UO_601 (O_601,N_4987,N_4924);
nand UO_602 (O_602,N_4972,N_4944);
nand UO_603 (O_603,N_4958,N_4906);
nor UO_604 (O_604,N_4882,N_4807);
nor UO_605 (O_605,N_4840,N_4830);
nor UO_606 (O_606,N_4874,N_4867);
and UO_607 (O_607,N_4821,N_4962);
nor UO_608 (O_608,N_4972,N_4994);
and UO_609 (O_609,N_4907,N_4922);
and UO_610 (O_610,N_4919,N_4994);
nor UO_611 (O_611,N_4947,N_4907);
and UO_612 (O_612,N_4840,N_4832);
or UO_613 (O_613,N_4937,N_4871);
nor UO_614 (O_614,N_4873,N_4918);
or UO_615 (O_615,N_4813,N_4992);
and UO_616 (O_616,N_4834,N_4968);
and UO_617 (O_617,N_4841,N_4859);
nand UO_618 (O_618,N_4877,N_4874);
and UO_619 (O_619,N_4872,N_4895);
nor UO_620 (O_620,N_4913,N_4854);
or UO_621 (O_621,N_4872,N_4874);
nor UO_622 (O_622,N_4852,N_4995);
nor UO_623 (O_623,N_4976,N_4832);
or UO_624 (O_624,N_4896,N_4855);
nand UO_625 (O_625,N_4981,N_4852);
or UO_626 (O_626,N_4995,N_4960);
nor UO_627 (O_627,N_4952,N_4902);
or UO_628 (O_628,N_4860,N_4973);
or UO_629 (O_629,N_4988,N_4866);
nand UO_630 (O_630,N_4848,N_4812);
nor UO_631 (O_631,N_4982,N_4878);
nand UO_632 (O_632,N_4971,N_4964);
nand UO_633 (O_633,N_4905,N_4821);
nand UO_634 (O_634,N_4802,N_4988);
nor UO_635 (O_635,N_4847,N_4853);
or UO_636 (O_636,N_4802,N_4839);
or UO_637 (O_637,N_4937,N_4828);
nand UO_638 (O_638,N_4877,N_4806);
and UO_639 (O_639,N_4879,N_4948);
and UO_640 (O_640,N_4812,N_4862);
or UO_641 (O_641,N_4934,N_4806);
nand UO_642 (O_642,N_4931,N_4924);
nor UO_643 (O_643,N_4946,N_4884);
or UO_644 (O_644,N_4955,N_4864);
and UO_645 (O_645,N_4997,N_4815);
or UO_646 (O_646,N_4857,N_4888);
and UO_647 (O_647,N_4866,N_4882);
nand UO_648 (O_648,N_4911,N_4811);
or UO_649 (O_649,N_4859,N_4877);
or UO_650 (O_650,N_4824,N_4918);
or UO_651 (O_651,N_4998,N_4903);
xor UO_652 (O_652,N_4948,N_4996);
nand UO_653 (O_653,N_4880,N_4902);
or UO_654 (O_654,N_4958,N_4968);
nor UO_655 (O_655,N_4930,N_4941);
nand UO_656 (O_656,N_4829,N_4984);
nor UO_657 (O_657,N_4862,N_4984);
or UO_658 (O_658,N_4954,N_4969);
and UO_659 (O_659,N_4957,N_4998);
and UO_660 (O_660,N_4949,N_4860);
nand UO_661 (O_661,N_4953,N_4822);
and UO_662 (O_662,N_4947,N_4849);
nor UO_663 (O_663,N_4974,N_4891);
nor UO_664 (O_664,N_4878,N_4985);
nor UO_665 (O_665,N_4887,N_4822);
or UO_666 (O_666,N_4834,N_4825);
and UO_667 (O_667,N_4825,N_4931);
nor UO_668 (O_668,N_4810,N_4807);
and UO_669 (O_669,N_4996,N_4981);
nor UO_670 (O_670,N_4924,N_4991);
or UO_671 (O_671,N_4921,N_4878);
nand UO_672 (O_672,N_4932,N_4919);
nand UO_673 (O_673,N_4877,N_4966);
nand UO_674 (O_674,N_4839,N_4918);
and UO_675 (O_675,N_4897,N_4808);
xnor UO_676 (O_676,N_4960,N_4806);
and UO_677 (O_677,N_4855,N_4993);
nand UO_678 (O_678,N_4821,N_4988);
nor UO_679 (O_679,N_4966,N_4965);
nand UO_680 (O_680,N_4894,N_4968);
or UO_681 (O_681,N_4879,N_4851);
xnor UO_682 (O_682,N_4914,N_4808);
or UO_683 (O_683,N_4871,N_4850);
nor UO_684 (O_684,N_4847,N_4882);
nor UO_685 (O_685,N_4924,N_4962);
and UO_686 (O_686,N_4980,N_4899);
and UO_687 (O_687,N_4946,N_4867);
and UO_688 (O_688,N_4805,N_4945);
or UO_689 (O_689,N_4923,N_4952);
or UO_690 (O_690,N_4869,N_4876);
nand UO_691 (O_691,N_4905,N_4992);
and UO_692 (O_692,N_4952,N_4943);
nor UO_693 (O_693,N_4818,N_4828);
nor UO_694 (O_694,N_4948,N_4918);
nor UO_695 (O_695,N_4839,N_4813);
or UO_696 (O_696,N_4971,N_4965);
or UO_697 (O_697,N_4809,N_4830);
nand UO_698 (O_698,N_4927,N_4979);
nand UO_699 (O_699,N_4994,N_4892);
and UO_700 (O_700,N_4809,N_4995);
and UO_701 (O_701,N_4908,N_4828);
or UO_702 (O_702,N_4934,N_4850);
nor UO_703 (O_703,N_4839,N_4955);
nand UO_704 (O_704,N_4821,N_4957);
and UO_705 (O_705,N_4950,N_4903);
nand UO_706 (O_706,N_4894,N_4800);
nor UO_707 (O_707,N_4821,N_4864);
or UO_708 (O_708,N_4958,N_4813);
nand UO_709 (O_709,N_4941,N_4841);
nand UO_710 (O_710,N_4867,N_4969);
nor UO_711 (O_711,N_4865,N_4874);
nor UO_712 (O_712,N_4892,N_4801);
nand UO_713 (O_713,N_4899,N_4844);
xor UO_714 (O_714,N_4903,N_4895);
or UO_715 (O_715,N_4805,N_4998);
nor UO_716 (O_716,N_4905,N_4802);
nand UO_717 (O_717,N_4986,N_4974);
or UO_718 (O_718,N_4840,N_4988);
and UO_719 (O_719,N_4862,N_4993);
nand UO_720 (O_720,N_4836,N_4942);
and UO_721 (O_721,N_4966,N_4980);
or UO_722 (O_722,N_4879,N_4920);
nor UO_723 (O_723,N_4988,N_4856);
nor UO_724 (O_724,N_4893,N_4830);
nor UO_725 (O_725,N_4925,N_4998);
and UO_726 (O_726,N_4918,N_4931);
and UO_727 (O_727,N_4838,N_4911);
nand UO_728 (O_728,N_4805,N_4891);
nand UO_729 (O_729,N_4928,N_4918);
nand UO_730 (O_730,N_4879,N_4893);
nand UO_731 (O_731,N_4850,N_4851);
and UO_732 (O_732,N_4805,N_4933);
or UO_733 (O_733,N_4971,N_4861);
or UO_734 (O_734,N_4880,N_4890);
or UO_735 (O_735,N_4898,N_4931);
nor UO_736 (O_736,N_4819,N_4962);
nand UO_737 (O_737,N_4970,N_4813);
and UO_738 (O_738,N_4895,N_4835);
nand UO_739 (O_739,N_4816,N_4908);
nor UO_740 (O_740,N_4809,N_4909);
nor UO_741 (O_741,N_4867,N_4979);
nand UO_742 (O_742,N_4837,N_4946);
or UO_743 (O_743,N_4886,N_4845);
and UO_744 (O_744,N_4883,N_4918);
or UO_745 (O_745,N_4854,N_4911);
or UO_746 (O_746,N_4874,N_4907);
or UO_747 (O_747,N_4896,N_4959);
nand UO_748 (O_748,N_4971,N_4867);
and UO_749 (O_749,N_4849,N_4978);
or UO_750 (O_750,N_4879,N_4995);
nor UO_751 (O_751,N_4973,N_4989);
and UO_752 (O_752,N_4970,N_4827);
nand UO_753 (O_753,N_4823,N_4846);
xor UO_754 (O_754,N_4831,N_4935);
and UO_755 (O_755,N_4850,N_4857);
and UO_756 (O_756,N_4975,N_4964);
or UO_757 (O_757,N_4959,N_4941);
nand UO_758 (O_758,N_4944,N_4983);
and UO_759 (O_759,N_4853,N_4898);
nor UO_760 (O_760,N_4961,N_4982);
or UO_761 (O_761,N_4923,N_4859);
and UO_762 (O_762,N_4831,N_4815);
nand UO_763 (O_763,N_4979,N_4871);
and UO_764 (O_764,N_4867,N_4910);
and UO_765 (O_765,N_4818,N_4921);
nand UO_766 (O_766,N_4995,N_4801);
or UO_767 (O_767,N_4898,N_4852);
nor UO_768 (O_768,N_4935,N_4991);
or UO_769 (O_769,N_4900,N_4966);
nand UO_770 (O_770,N_4985,N_4888);
nand UO_771 (O_771,N_4949,N_4832);
nand UO_772 (O_772,N_4891,N_4851);
nor UO_773 (O_773,N_4974,N_4927);
or UO_774 (O_774,N_4822,N_4886);
nand UO_775 (O_775,N_4945,N_4928);
nor UO_776 (O_776,N_4811,N_4844);
and UO_777 (O_777,N_4873,N_4995);
and UO_778 (O_778,N_4804,N_4833);
nor UO_779 (O_779,N_4858,N_4818);
or UO_780 (O_780,N_4982,N_4983);
or UO_781 (O_781,N_4912,N_4891);
nand UO_782 (O_782,N_4991,N_4941);
nor UO_783 (O_783,N_4869,N_4992);
or UO_784 (O_784,N_4998,N_4993);
and UO_785 (O_785,N_4814,N_4993);
nand UO_786 (O_786,N_4962,N_4811);
nor UO_787 (O_787,N_4808,N_4968);
nand UO_788 (O_788,N_4857,N_4960);
nor UO_789 (O_789,N_4941,N_4975);
or UO_790 (O_790,N_4976,N_4921);
and UO_791 (O_791,N_4959,N_4887);
or UO_792 (O_792,N_4905,N_4924);
nand UO_793 (O_793,N_4954,N_4818);
or UO_794 (O_794,N_4866,N_4993);
and UO_795 (O_795,N_4939,N_4849);
nor UO_796 (O_796,N_4852,N_4943);
xnor UO_797 (O_797,N_4950,N_4995);
nor UO_798 (O_798,N_4848,N_4845);
and UO_799 (O_799,N_4960,N_4888);
or UO_800 (O_800,N_4948,N_4901);
or UO_801 (O_801,N_4838,N_4906);
or UO_802 (O_802,N_4985,N_4900);
nand UO_803 (O_803,N_4913,N_4827);
nand UO_804 (O_804,N_4991,N_4815);
or UO_805 (O_805,N_4962,N_4992);
or UO_806 (O_806,N_4852,N_4829);
or UO_807 (O_807,N_4996,N_4879);
or UO_808 (O_808,N_4849,N_4881);
nor UO_809 (O_809,N_4896,N_4885);
or UO_810 (O_810,N_4912,N_4994);
nor UO_811 (O_811,N_4941,N_4830);
nor UO_812 (O_812,N_4980,N_4958);
nand UO_813 (O_813,N_4890,N_4804);
nor UO_814 (O_814,N_4938,N_4855);
nand UO_815 (O_815,N_4821,N_4929);
nor UO_816 (O_816,N_4958,N_4979);
nand UO_817 (O_817,N_4851,N_4800);
nand UO_818 (O_818,N_4816,N_4886);
and UO_819 (O_819,N_4976,N_4926);
nor UO_820 (O_820,N_4826,N_4932);
nor UO_821 (O_821,N_4936,N_4812);
and UO_822 (O_822,N_4898,N_4965);
nand UO_823 (O_823,N_4908,N_4957);
nor UO_824 (O_824,N_4840,N_4949);
or UO_825 (O_825,N_4838,N_4929);
nor UO_826 (O_826,N_4919,N_4992);
xnor UO_827 (O_827,N_4895,N_4966);
xor UO_828 (O_828,N_4854,N_4872);
nand UO_829 (O_829,N_4991,N_4904);
or UO_830 (O_830,N_4942,N_4954);
nand UO_831 (O_831,N_4876,N_4844);
nor UO_832 (O_832,N_4936,N_4938);
nand UO_833 (O_833,N_4903,N_4893);
nand UO_834 (O_834,N_4845,N_4868);
nor UO_835 (O_835,N_4969,N_4933);
and UO_836 (O_836,N_4972,N_4983);
nand UO_837 (O_837,N_4913,N_4921);
nand UO_838 (O_838,N_4818,N_4978);
or UO_839 (O_839,N_4826,N_4849);
or UO_840 (O_840,N_4934,N_4861);
and UO_841 (O_841,N_4827,N_4928);
nor UO_842 (O_842,N_4999,N_4878);
and UO_843 (O_843,N_4974,N_4870);
or UO_844 (O_844,N_4818,N_4950);
xnor UO_845 (O_845,N_4933,N_4847);
nand UO_846 (O_846,N_4990,N_4872);
nor UO_847 (O_847,N_4949,N_4892);
nand UO_848 (O_848,N_4906,N_4967);
nand UO_849 (O_849,N_4885,N_4976);
nand UO_850 (O_850,N_4801,N_4953);
and UO_851 (O_851,N_4866,N_4840);
and UO_852 (O_852,N_4815,N_4919);
nor UO_853 (O_853,N_4990,N_4972);
xnor UO_854 (O_854,N_4800,N_4914);
nand UO_855 (O_855,N_4849,N_4977);
nor UO_856 (O_856,N_4904,N_4908);
nor UO_857 (O_857,N_4825,N_4845);
or UO_858 (O_858,N_4973,N_4831);
or UO_859 (O_859,N_4943,N_4989);
and UO_860 (O_860,N_4964,N_4912);
nand UO_861 (O_861,N_4896,N_4940);
nand UO_862 (O_862,N_4822,N_4839);
or UO_863 (O_863,N_4809,N_4825);
nor UO_864 (O_864,N_4814,N_4951);
or UO_865 (O_865,N_4886,N_4810);
nor UO_866 (O_866,N_4818,N_4946);
nand UO_867 (O_867,N_4839,N_4898);
or UO_868 (O_868,N_4960,N_4824);
nand UO_869 (O_869,N_4999,N_4800);
and UO_870 (O_870,N_4819,N_4923);
nand UO_871 (O_871,N_4909,N_4862);
or UO_872 (O_872,N_4918,N_4974);
nor UO_873 (O_873,N_4833,N_4955);
or UO_874 (O_874,N_4973,N_4996);
xnor UO_875 (O_875,N_4903,N_4896);
nor UO_876 (O_876,N_4922,N_4987);
and UO_877 (O_877,N_4808,N_4870);
or UO_878 (O_878,N_4911,N_4860);
nor UO_879 (O_879,N_4896,N_4931);
or UO_880 (O_880,N_4992,N_4885);
nand UO_881 (O_881,N_4902,N_4817);
nor UO_882 (O_882,N_4950,N_4819);
and UO_883 (O_883,N_4927,N_4845);
nor UO_884 (O_884,N_4884,N_4970);
nor UO_885 (O_885,N_4846,N_4828);
or UO_886 (O_886,N_4897,N_4889);
or UO_887 (O_887,N_4931,N_4865);
nand UO_888 (O_888,N_4997,N_4931);
nand UO_889 (O_889,N_4902,N_4845);
nand UO_890 (O_890,N_4864,N_4920);
or UO_891 (O_891,N_4801,N_4852);
nor UO_892 (O_892,N_4900,N_4957);
nor UO_893 (O_893,N_4984,N_4805);
nand UO_894 (O_894,N_4929,N_4946);
and UO_895 (O_895,N_4820,N_4899);
and UO_896 (O_896,N_4908,N_4851);
nor UO_897 (O_897,N_4907,N_4813);
or UO_898 (O_898,N_4983,N_4836);
and UO_899 (O_899,N_4856,N_4803);
nor UO_900 (O_900,N_4815,N_4884);
nand UO_901 (O_901,N_4808,N_4907);
nand UO_902 (O_902,N_4887,N_4937);
and UO_903 (O_903,N_4808,N_4893);
nor UO_904 (O_904,N_4917,N_4829);
nor UO_905 (O_905,N_4801,N_4999);
nor UO_906 (O_906,N_4978,N_4979);
nand UO_907 (O_907,N_4823,N_4949);
nand UO_908 (O_908,N_4973,N_4892);
nor UO_909 (O_909,N_4976,N_4860);
nor UO_910 (O_910,N_4919,N_4900);
or UO_911 (O_911,N_4855,N_4974);
nand UO_912 (O_912,N_4869,N_4895);
or UO_913 (O_913,N_4975,N_4845);
and UO_914 (O_914,N_4952,N_4947);
nor UO_915 (O_915,N_4957,N_4963);
and UO_916 (O_916,N_4953,N_4965);
xor UO_917 (O_917,N_4823,N_4904);
nor UO_918 (O_918,N_4851,N_4952);
and UO_919 (O_919,N_4864,N_4848);
nand UO_920 (O_920,N_4882,N_4945);
nand UO_921 (O_921,N_4940,N_4815);
or UO_922 (O_922,N_4995,N_4969);
nand UO_923 (O_923,N_4970,N_4957);
and UO_924 (O_924,N_4833,N_4813);
and UO_925 (O_925,N_4990,N_4913);
nand UO_926 (O_926,N_4974,N_4931);
nand UO_927 (O_927,N_4893,N_4946);
and UO_928 (O_928,N_4935,N_4930);
or UO_929 (O_929,N_4995,N_4985);
xnor UO_930 (O_930,N_4969,N_4918);
or UO_931 (O_931,N_4858,N_4857);
or UO_932 (O_932,N_4979,N_4986);
or UO_933 (O_933,N_4937,N_4927);
nand UO_934 (O_934,N_4850,N_4816);
nor UO_935 (O_935,N_4906,N_4808);
and UO_936 (O_936,N_4983,N_4977);
and UO_937 (O_937,N_4963,N_4900);
and UO_938 (O_938,N_4931,N_4917);
nor UO_939 (O_939,N_4999,N_4850);
nand UO_940 (O_940,N_4901,N_4862);
nand UO_941 (O_941,N_4820,N_4922);
and UO_942 (O_942,N_4880,N_4979);
and UO_943 (O_943,N_4802,N_4927);
and UO_944 (O_944,N_4992,N_4880);
and UO_945 (O_945,N_4986,N_4843);
and UO_946 (O_946,N_4919,N_4955);
nand UO_947 (O_947,N_4809,N_4988);
and UO_948 (O_948,N_4897,N_4966);
nor UO_949 (O_949,N_4948,N_4886);
nor UO_950 (O_950,N_4948,N_4855);
nand UO_951 (O_951,N_4847,N_4952);
nor UO_952 (O_952,N_4806,N_4936);
nand UO_953 (O_953,N_4922,N_4811);
xnor UO_954 (O_954,N_4831,N_4993);
and UO_955 (O_955,N_4968,N_4953);
and UO_956 (O_956,N_4991,N_4931);
xnor UO_957 (O_957,N_4815,N_4900);
nand UO_958 (O_958,N_4918,N_4999);
nand UO_959 (O_959,N_4946,N_4940);
nor UO_960 (O_960,N_4833,N_4919);
nand UO_961 (O_961,N_4883,N_4895);
or UO_962 (O_962,N_4872,N_4800);
nor UO_963 (O_963,N_4836,N_4869);
and UO_964 (O_964,N_4959,N_4831);
xnor UO_965 (O_965,N_4905,N_4887);
nand UO_966 (O_966,N_4827,N_4825);
and UO_967 (O_967,N_4952,N_4818);
nor UO_968 (O_968,N_4814,N_4950);
or UO_969 (O_969,N_4943,N_4832);
or UO_970 (O_970,N_4895,N_4907);
or UO_971 (O_971,N_4918,N_4955);
nor UO_972 (O_972,N_4898,N_4837);
and UO_973 (O_973,N_4947,N_4870);
nor UO_974 (O_974,N_4925,N_4903);
or UO_975 (O_975,N_4892,N_4842);
and UO_976 (O_976,N_4923,N_4944);
nor UO_977 (O_977,N_4934,N_4935);
or UO_978 (O_978,N_4935,N_4815);
nand UO_979 (O_979,N_4910,N_4921);
or UO_980 (O_980,N_4846,N_4940);
and UO_981 (O_981,N_4962,N_4892);
or UO_982 (O_982,N_4999,N_4975);
nand UO_983 (O_983,N_4889,N_4999);
and UO_984 (O_984,N_4807,N_4809);
nor UO_985 (O_985,N_4997,N_4959);
nor UO_986 (O_986,N_4989,N_4935);
or UO_987 (O_987,N_4926,N_4940);
and UO_988 (O_988,N_4942,N_4873);
nor UO_989 (O_989,N_4952,N_4973);
and UO_990 (O_990,N_4884,N_4940);
nand UO_991 (O_991,N_4814,N_4883);
nor UO_992 (O_992,N_4901,N_4990);
nor UO_993 (O_993,N_4869,N_4851);
nand UO_994 (O_994,N_4953,N_4961);
nand UO_995 (O_995,N_4872,N_4806);
and UO_996 (O_996,N_4984,N_4825);
nand UO_997 (O_997,N_4934,N_4920);
or UO_998 (O_998,N_4997,N_4804);
nand UO_999 (O_999,N_4833,N_4956);
endmodule