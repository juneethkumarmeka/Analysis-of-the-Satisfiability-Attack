module basic_750_5000_1000_10_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xnor U0 (N_0,In_731,In_163);
nand U1 (N_1,In_481,In_143);
xor U2 (N_2,In_589,In_431);
and U3 (N_3,In_345,In_661);
or U4 (N_4,In_720,In_99);
or U5 (N_5,In_166,In_16);
nor U6 (N_6,In_286,In_502);
xor U7 (N_7,In_477,In_562);
and U8 (N_8,In_214,In_637);
and U9 (N_9,In_56,In_256);
or U10 (N_10,In_83,In_740);
or U11 (N_11,In_538,In_625);
nor U12 (N_12,In_660,In_691);
and U13 (N_13,In_483,In_692);
nand U14 (N_14,In_631,In_612);
nand U15 (N_15,In_215,In_123);
or U16 (N_16,In_383,In_485);
nand U17 (N_17,In_197,In_87);
nand U18 (N_18,In_743,In_742);
or U19 (N_19,In_261,In_162);
nor U20 (N_20,In_192,In_218);
nand U21 (N_21,In_198,In_330);
or U22 (N_22,In_668,In_333);
and U23 (N_23,In_216,In_405);
nor U24 (N_24,In_86,In_316);
xnor U25 (N_25,In_125,In_274);
and U26 (N_26,In_103,In_540);
nor U27 (N_27,In_548,In_91);
or U28 (N_28,In_194,In_2);
nand U29 (N_29,In_124,In_68);
nand U30 (N_30,In_242,In_257);
xnor U31 (N_31,In_558,In_642);
nand U32 (N_32,In_12,In_524);
or U33 (N_33,In_335,In_526);
or U34 (N_34,In_394,In_587);
and U35 (N_35,In_13,In_357);
nand U36 (N_36,In_325,In_133);
xor U37 (N_37,In_728,In_453);
nor U38 (N_38,In_654,In_493);
or U39 (N_39,In_259,In_672);
nor U40 (N_40,In_377,In_293);
nand U41 (N_41,In_469,In_295);
nor U42 (N_42,In_456,In_559);
nand U43 (N_43,In_421,In_26);
xnor U44 (N_44,In_449,In_73);
xor U45 (N_45,In_423,In_420);
or U46 (N_46,In_544,In_213);
and U47 (N_47,In_307,In_250);
and U48 (N_48,In_641,In_247);
nor U49 (N_49,In_80,In_306);
nor U50 (N_50,In_535,In_248);
and U51 (N_51,In_600,In_181);
or U52 (N_52,In_28,In_165);
or U53 (N_53,In_288,In_365);
or U54 (N_54,In_406,In_14);
and U55 (N_55,In_713,In_348);
nand U56 (N_56,In_161,In_496);
and U57 (N_57,In_200,In_463);
or U58 (N_58,In_37,In_734);
xor U59 (N_59,In_499,In_520);
and U60 (N_60,In_188,In_311);
or U61 (N_61,In_53,In_573);
nor U62 (N_62,In_690,In_171);
or U63 (N_63,In_82,In_252);
nand U64 (N_64,In_627,In_22);
xnor U65 (N_65,In_390,In_706);
nor U66 (N_66,In_225,In_310);
and U67 (N_67,In_336,In_9);
xnor U68 (N_68,In_506,In_131);
or U69 (N_69,In_135,In_364);
and U70 (N_70,In_164,In_623);
or U71 (N_71,In_684,In_458);
and U72 (N_72,In_615,In_253);
xor U73 (N_73,In_422,In_55);
or U74 (N_74,In_238,In_111);
or U75 (N_75,In_211,In_566);
and U76 (N_76,In_403,In_292);
or U77 (N_77,In_237,In_598);
nor U78 (N_78,In_104,In_552);
and U79 (N_79,In_533,In_318);
nand U80 (N_80,In_355,In_117);
or U81 (N_81,In_592,In_351);
nand U82 (N_82,In_694,In_514);
and U83 (N_83,In_11,In_110);
nand U84 (N_84,In_650,In_255);
or U85 (N_85,In_475,In_50);
or U86 (N_86,In_314,In_379);
or U87 (N_87,In_128,In_399);
nand U88 (N_88,In_374,In_685);
nand U89 (N_89,In_705,In_205);
and U90 (N_90,In_85,In_435);
and U91 (N_91,In_378,In_150);
and U92 (N_92,In_262,In_354);
or U93 (N_93,In_636,In_346);
nor U94 (N_94,In_33,In_301);
and U95 (N_95,In_386,In_490);
nand U96 (N_96,In_294,In_8);
nand U97 (N_97,In_34,In_375);
or U98 (N_98,In_582,In_302);
nand U99 (N_99,In_560,In_368);
and U100 (N_100,In_509,In_279);
or U101 (N_101,In_140,In_66);
nor U102 (N_102,In_107,In_681);
nor U103 (N_103,In_465,In_596);
and U104 (N_104,In_507,In_670);
nor U105 (N_105,In_411,In_460);
nand U106 (N_106,In_519,In_608);
xnor U107 (N_107,In_682,In_510);
nand U108 (N_108,In_737,In_64);
xor U109 (N_109,In_84,In_652);
and U110 (N_110,In_438,In_715);
or U111 (N_111,In_576,In_480);
and U112 (N_112,In_504,In_696);
nor U113 (N_113,In_381,In_602);
xor U114 (N_114,In_572,In_425);
nor U115 (N_115,In_699,In_462);
and U116 (N_116,In_227,In_605);
or U117 (N_117,In_450,In_349);
nor U118 (N_118,In_268,In_467);
and U119 (N_119,In_707,In_141);
and U120 (N_120,In_347,In_733);
xor U121 (N_121,In_601,In_69);
xor U122 (N_122,In_554,In_233);
or U123 (N_123,In_142,In_254);
or U124 (N_124,In_749,In_353);
nand U125 (N_125,In_428,In_443);
and U126 (N_126,In_183,In_235);
nand U127 (N_127,In_223,In_474);
nand U128 (N_128,In_424,In_640);
nand U129 (N_129,In_49,In_338);
or U130 (N_130,In_380,In_284);
or U131 (N_131,In_398,In_167);
or U132 (N_132,In_352,In_470);
nand U133 (N_133,In_624,In_436);
or U134 (N_134,In_178,In_437);
nor U135 (N_135,In_714,In_639);
nor U136 (N_136,In_291,In_290);
and U137 (N_137,In_39,In_471);
nor U138 (N_138,In_100,In_645);
or U139 (N_139,In_617,In_173);
xnor U140 (N_140,In_169,In_657);
nand U141 (N_141,In_275,In_102);
xnor U142 (N_142,In_426,In_182);
and U143 (N_143,In_669,In_630);
nand U144 (N_144,In_258,In_444);
nor U145 (N_145,In_18,In_210);
xor U146 (N_146,In_663,In_92);
nand U147 (N_147,In_747,In_3);
and U148 (N_148,In_675,In_67);
nand U149 (N_149,In_716,In_446);
nor U150 (N_150,In_129,In_146);
xor U151 (N_151,In_666,In_413);
and U152 (N_152,In_704,In_145);
or U153 (N_153,In_323,In_479);
and U154 (N_154,In_410,In_79);
or U155 (N_155,In_695,In_303);
nor U156 (N_156,In_531,In_246);
or U157 (N_157,In_196,In_6);
nand U158 (N_158,In_584,In_571);
and U159 (N_159,In_676,In_62);
or U160 (N_160,In_47,In_580);
and U161 (N_161,In_54,In_546);
and U162 (N_162,In_702,In_270);
and U163 (N_163,In_241,In_429);
or U164 (N_164,In_468,In_189);
or U165 (N_165,In_698,In_452);
and U166 (N_166,In_498,In_484);
nand U167 (N_167,In_667,In_144);
nand U168 (N_168,In_209,In_719);
and U169 (N_169,In_384,In_25);
nor U170 (N_170,In_473,In_220);
nand U171 (N_171,In_539,In_563);
nand U172 (N_172,In_57,In_319);
nand U173 (N_173,In_635,In_711);
xnor U174 (N_174,In_680,In_387);
or U175 (N_175,In_15,In_500);
nand U176 (N_176,In_611,In_120);
and U177 (N_177,In_505,In_95);
xnor U178 (N_178,In_81,In_606);
nor U179 (N_179,In_23,In_172);
and U180 (N_180,In_727,In_595);
or U181 (N_181,In_697,In_432);
nand U182 (N_182,In_170,In_597);
or U183 (N_183,In_689,In_151);
and U184 (N_184,In_108,In_289);
or U185 (N_185,In_362,In_708);
nor U186 (N_186,In_190,In_542);
nor U187 (N_187,In_187,In_551);
and U188 (N_188,In_412,In_679);
xnor U189 (N_189,In_441,In_52);
nor U190 (N_190,In_646,In_735);
and U191 (N_191,In_360,In_59);
xor U192 (N_192,In_430,In_653);
or U193 (N_193,In_723,In_409);
or U194 (N_194,In_334,In_76);
and U195 (N_195,In_260,In_287);
or U196 (N_196,In_71,In_358);
and U197 (N_197,In_89,In_647);
nand U198 (N_198,In_494,In_119);
or U199 (N_199,In_344,In_547);
nand U200 (N_200,In_243,In_603);
nand U201 (N_201,In_72,In_495);
nor U202 (N_202,In_4,In_557);
xnor U203 (N_203,In_701,In_46);
nor U204 (N_204,In_326,In_664);
or U205 (N_205,In_251,In_382);
xnor U206 (N_206,In_553,In_320);
or U207 (N_207,In_315,In_370);
xnor U208 (N_208,In_414,In_512);
nor U209 (N_209,In_492,In_231);
or U210 (N_210,In_298,In_296);
nand U211 (N_211,In_417,In_401);
nand U212 (N_212,In_363,In_583);
nand U213 (N_213,In_322,In_543);
xor U214 (N_214,In_276,In_127);
and U215 (N_215,In_175,In_523);
xnor U216 (N_216,In_249,In_193);
and U217 (N_217,In_497,In_244);
and U218 (N_218,In_10,In_581);
nor U219 (N_219,In_264,In_725);
nand U220 (N_220,In_40,In_281);
nand U221 (N_221,In_204,In_439);
or U222 (N_222,In_313,In_299);
xnor U223 (N_223,In_155,In_78);
and U224 (N_224,In_65,In_208);
nor U225 (N_225,In_651,In_221);
nand U226 (N_226,In_232,In_112);
nor U227 (N_227,In_516,In_638);
and U228 (N_228,In_36,In_622);
and U229 (N_229,In_659,In_245);
nand U230 (N_230,In_472,In_137);
or U231 (N_231,In_152,In_674);
or U232 (N_232,In_525,In_199);
or U233 (N_233,In_17,In_101);
xnor U234 (N_234,In_388,In_722);
and U235 (N_235,In_457,In_570);
nor U236 (N_236,In_732,In_447);
or U237 (N_237,In_487,In_272);
nand U238 (N_238,In_226,In_356);
and U239 (N_239,In_105,In_139);
xor U240 (N_240,In_561,In_219);
nand U241 (N_241,In_738,In_515);
nor U242 (N_242,In_109,In_545);
and U243 (N_243,In_748,In_649);
or U244 (N_244,In_74,In_361);
nor U245 (N_245,In_565,In_343);
nor U246 (N_246,In_230,In_1);
nor U247 (N_247,In_454,In_568);
and U248 (N_248,In_138,In_369);
nand U249 (N_249,In_38,In_41);
or U250 (N_250,In_709,In_700);
or U251 (N_251,In_459,In_195);
and U252 (N_252,In_376,In_550);
and U253 (N_253,In_207,In_304);
xor U254 (N_254,In_522,In_671);
nor U255 (N_255,In_407,In_445);
nor U256 (N_256,In_574,In_32);
or U257 (N_257,In_564,In_317);
nor U258 (N_258,In_419,In_621);
or U259 (N_259,In_312,In_180);
xnor U260 (N_260,In_229,In_404);
nor U261 (N_261,In_359,In_517);
nand U262 (N_262,In_27,In_393);
and U263 (N_263,In_35,In_130);
nand U264 (N_264,In_511,In_741);
or U265 (N_265,In_367,In_433);
or U266 (N_266,In_5,In_385);
nand U267 (N_267,In_427,In_159);
and U268 (N_268,In_285,In_686);
xnor U269 (N_269,In_341,In_331);
and U270 (N_270,In_478,In_416);
nand U271 (N_271,In_594,In_30);
nor U272 (N_272,In_739,In_97);
xnor U273 (N_273,In_488,In_618);
nand U274 (N_274,In_116,In_578);
nand U275 (N_275,In_521,In_461);
nor U276 (N_276,In_541,In_44);
nand U277 (N_277,In_342,In_308);
and U278 (N_278,In_154,In_19);
or U279 (N_279,In_212,In_201);
nand U280 (N_280,In_729,In_632);
xor U281 (N_281,In_392,In_29);
or U282 (N_282,In_577,In_489);
or U283 (N_283,In_389,In_662);
or U284 (N_284,In_98,In_93);
and U285 (N_285,In_328,In_324);
xnor U286 (N_286,In_549,In_185);
and U287 (N_287,In_282,In_567);
and U288 (N_288,In_263,In_327);
nor U289 (N_289,In_45,In_58);
nor U290 (N_290,In_147,In_300);
nand U291 (N_291,In_217,In_156);
nand U292 (N_292,In_96,In_528);
xnor U293 (N_293,In_332,In_202);
nand U294 (N_294,In_277,In_466);
or U295 (N_295,In_575,In_616);
xnor U296 (N_296,In_136,In_114);
and U297 (N_297,In_234,In_77);
and U298 (N_298,In_486,In_665);
and U299 (N_299,In_132,In_31);
or U300 (N_300,In_75,In_527);
or U301 (N_301,In_337,In_113);
or U302 (N_302,In_633,In_297);
and U303 (N_303,In_0,In_745);
or U304 (N_304,In_513,In_121);
or U305 (N_305,In_203,In_501);
nor U306 (N_306,In_21,In_518);
and U307 (N_307,In_350,In_191);
nand U308 (N_308,In_7,In_148);
and U309 (N_309,In_391,In_585);
and U310 (N_310,In_532,In_122);
or U311 (N_311,In_48,In_569);
or U312 (N_312,In_442,In_280);
and U313 (N_313,In_643,In_366);
and U314 (N_314,In_599,In_464);
or U315 (N_315,In_717,In_157);
nand U316 (N_316,In_556,In_373);
or U317 (N_317,In_94,In_683);
and U318 (N_318,In_688,In_586);
xnor U319 (N_319,In_371,In_476);
nand U320 (N_320,In_530,In_395);
xor U321 (N_321,In_179,In_160);
or U322 (N_322,In_176,In_309);
nor U323 (N_323,In_656,In_60);
nor U324 (N_324,In_730,In_712);
nor U325 (N_325,In_613,In_174);
or U326 (N_326,In_408,In_222);
or U327 (N_327,In_628,In_61);
or U328 (N_328,In_415,In_455);
or U329 (N_329,In_434,In_534);
or U330 (N_330,In_149,In_491);
nand U331 (N_331,In_158,In_88);
nor U332 (N_332,In_448,In_440);
nand U333 (N_333,In_206,In_655);
nand U334 (N_334,In_609,In_746);
nand U335 (N_335,In_51,In_724);
or U336 (N_336,In_24,In_153);
nand U337 (N_337,In_590,In_591);
and U338 (N_338,In_20,In_115);
xor U339 (N_339,In_677,In_619);
xnor U340 (N_340,In_673,In_168);
xor U341 (N_341,In_239,In_106);
and U342 (N_342,In_482,In_503);
and U343 (N_343,In_634,In_693);
nand U344 (N_344,In_42,In_43);
nand U345 (N_345,In_579,In_271);
and U346 (N_346,In_658,In_536);
nand U347 (N_347,In_118,In_278);
or U348 (N_348,In_372,In_228);
xnor U349 (N_349,In_744,In_269);
and U350 (N_350,In_236,In_678);
and U351 (N_351,In_687,In_451);
nand U352 (N_352,In_90,In_321);
nand U353 (N_353,In_397,In_644);
nand U354 (N_354,In_710,In_126);
or U355 (N_355,In_593,In_555);
and U356 (N_356,In_529,In_726);
or U357 (N_357,In_186,In_177);
and U358 (N_358,In_224,In_607);
or U359 (N_359,In_63,In_273);
nand U360 (N_360,In_134,In_604);
or U361 (N_361,In_703,In_240);
and U362 (N_362,In_340,In_184);
and U363 (N_363,In_400,In_648);
xnor U364 (N_364,In_537,In_736);
nand U365 (N_365,In_588,In_329);
nor U366 (N_366,In_396,In_614);
nand U367 (N_367,In_70,In_620);
and U368 (N_368,In_265,In_305);
or U369 (N_369,In_339,In_402);
nor U370 (N_370,In_718,In_266);
nand U371 (N_371,In_629,In_267);
or U372 (N_372,In_508,In_626);
nor U373 (N_373,In_418,In_721);
or U374 (N_374,In_283,In_610);
and U375 (N_375,In_281,In_58);
nor U376 (N_376,In_244,In_442);
nand U377 (N_377,In_179,In_76);
xor U378 (N_378,In_154,In_705);
nand U379 (N_379,In_320,In_188);
nor U380 (N_380,In_514,In_597);
or U381 (N_381,In_140,In_40);
nor U382 (N_382,In_741,In_596);
nand U383 (N_383,In_728,In_711);
nand U384 (N_384,In_125,In_702);
nand U385 (N_385,In_448,In_347);
xor U386 (N_386,In_465,In_441);
and U387 (N_387,In_587,In_172);
and U388 (N_388,In_154,In_612);
or U389 (N_389,In_665,In_188);
or U390 (N_390,In_538,In_394);
and U391 (N_391,In_689,In_353);
nor U392 (N_392,In_632,In_593);
nor U393 (N_393,In_99,In_532);
and U394 (N_394,In_723,In_636);
nor U395 (N_395,In_247,In_736);
and U396 (N_396,In_460,In_383);
nand U397 (N_397,In_142,In_471);
nor U398 (N_398,In_598,In_145);
or U399 (N_399,In_21,In_586);
nand U400 (N_400,In_712,In_105);
xnor U401 (N_401,In_366,In_530);
nand U402 (N_402,In_257,In_379);
and U403 (N_403,In_302,In_216);
and U404 (N_404,In_104,In_208);
and U405 (N_405,In_496,In_603);
nor U406 (N_406,In_662,In_359);
or U407 (N_407,In_386,In_338);
nor U408 (N_408,In_412,In_703);
and U409 (N_409,In_35,In_499);
and U410 (N_410,In_644,In_575);
or U411 (N_411,In_722,In_740);
or U412 (N_412,In_166,In_448);
nand U413 (N_413,In_363,In_184);
nor U414 (N_414,In_91,In_628);
and U415 (N_415,In_31,In_84);
nor U416 (N_416,In_21,In_330);
nor U417 (N_417,In_412,In_211);
nor U418 (N_418,In_666,In_389);
nand U419 (N_419,In_645,In_202);
or U420 (N_420,In_321,In_507);
or U421 (N_421,In_386,In_372);
nor U422 (N_422,In_721,In_455);
nand U423 (N_423,In_363,In_687);
nor U424 (N_424,In_393,In_682);
or U425 (N_425,In_384,In_249);
nor U426 (N_426,In_19,In_417);
and U427 (N_427,In_331,In_227);
nand U428 (N_428,In_291,In_533);
xnor U429 (N_429,In_197,In_600);
and U430 (N_430,In_685,In_509);
and U431 (N_431,In_553,In_747);
and U432 (N_432,In_680,In_185);
nand U433 (N_433,In_277,In_665);
and U434 (N_434,In_551,In_429);
nor U435 (N_435,In_323,In_141);
or U436 (N_436,In_548,In_71);
nand U437 (N_437,In_48,In_121);
nand U438 (N_438,In_328,In_393);
or U439 (N_439,In_451,In_167);
nand U440 (N_440,In_285,In_185);
nand U441 (N_441,In_746,In_515);
and U442 (N_442,In_626,In_578);
xor U443 (N_443,In_391,In_621);
nor U444 (N_444,In_156,In_381);
nand U445 (N_445,In_254,In_582);
and U446 (N_446,In_455,In_394);
or U447 (N_447,In_280,In_286);
nand U448 (N_448,In_42,In_430);
and U449 (N_449,In_381,In_426);
nor U450 (N_450,In_92,In_711);
nand U451 (N_451,In_98,In_470);
nand U452 (N_452,In_448,In_212);
and U453 (N_453,In_184,In_695);
xor U454 (N_454,In_418,In_588);
and U455 (N_455,In_402,In_476);
xor U456 (N_456,In_708,In_19);
nor U457 (N_457,In_607,In_11);
nand U458 (N_458,In_328,In_363);
nand U459 (N_459,In_194,In_58);
and U460 (N_460,In_516,In_459);
xor U461 (N_461,In_423,In_614);
xor U462 (N_462,In_562,In_312);
and U463 (N_463,In_275,In_671);
and U464 (N_464,In_261,In_482);
or U465 (N_465,In_323,In_348);
nor U466 (N_466,In_487,In_351);
nand U467 (N_467,In_657,In_472);
nand U468 (N_468,In_309,In_167);
or U469 (N_469,In_469,In_587);
or U470 (N_470,In_735,In_60);
or U471 (N_471,In_186,In_184);
or U472 (N_472,In_399,In_8);
nor U473 (N_473,In_680,In_602);
nor U474 (N_474,In_601,In_660);
and U475 (N_475,In_647,In_154);
or U476 (N_476,In_115,In_302);
or U477 (N_477,In_661,In_421);
and U478 (N_478,In_740,In_316);
nand U479 (N_479,In_448,In_491);
nor U480 (N_480,In_281,In_742);
xnor U481 (N_481,In_311,In_366);
and U482 (N_482,In_613,In_621);
nor U483 (N_483,In_77,In_303);
nand U484 (N_484,In_429,In_332);
and U485 (N_485,In_207,In_332);
nand U486 (N_486,In_395,In_67);
xor U487 (N_487,In_36,In_83);
and U488 (N_488,In_662,In_0);
nor U489 (N_489,In_129,In_567);
nor U490 (N_490,In_39,In_134);
nor U491 (N_491,In_655,In_93);
nor U492 (N_492,In_100,In_193);
nor U493 (N_493,In_513,In_501);
or U494 (N_494,In_285,In_375);
nor U495 (N_495,In_223,In_183);
nand U496 (N_496,In_349,In_161);
or U497 (N_497,In_684,In_530);
nand U498 (N_498,In_197,In_713);
or U499 (N_499,In_723,In_118);
nand U500 (N_500,N_376,N_208);
nor U501 (N_501,N_192,N_462);
xor U502 (N_502,N_85,N_33);
and U503 (N_503,N_206,N_443);
nor U504 (N_504,N_482,N_8);
and U505 (N_505,N_143,N_497);
or U506 (N_506,N_254,N_100);
and U507 (N_507,N_223,N_12);
nand U508 (N_508,N_127,N_160);
nor U509 (N_509,N_40,N_377);
and U510 (N_510,N_179,N_409);
and U511 (N_511,N_251,N_315);
or U512 (N_512,N_398,N_450);
nor U513 (N_513,N_296,N_330);
nor U514 (N_514,N_467,N_322);
nand U515 (N_515,N_129,N_280);
nand U516 (N_516,N_426,N_123);
nand U517 (N_517,N_386,N_42);
nand U518 (N_518,N_29,N_381);
nand U519 (N_519,N_117,N_360);
and U520 (N_520,N_263,N_422);
nand U521 (N_521,N_397,N_256);
nand U522 (N_522,N_162,N_358);
nor U523 (N_523,N_199,N_444);
nor U524 (N_524,N_483,N_420);
or U525 (N_525,N_135,N_364);
nand U526 (N_526,N_425,N_156);
and U527 (N_527,N_18,N_242);
and U528 (N_528,N_101,N_212);
and U529 (N_529,N_11,N_114);
and U530 (N_530,N_459,N_173);
or U531 (N_531,N_16,N_436);
and U532 (N_532,N_357,N_204);
and U533 (N_533,N_168,N_41);
nor U534 (N_534,N_267,N_488);
or U535 (N_535,N_468,N_83);
xor U536 (N_536,N_189,N_217);
nor U537 (N_537,N_105,N_463);
and U538 (N_538,N_164,N_258);
and U539 (N_539,N_132,N_421);
nand U540 (N_540,N_55,N_466);
nor U541 (N_541,N_495,N_356);
or U542 (N_542,N_210,N_261);
nor U543 (N_543,N_23,N_485);
xnor U544 (N_544,N_22,N_266);
nor U545 (N_545,N_219,N_452);
nand U546 (N_546,N_379,N_26);
nor U547 (N_547,N_6,N_259);
or U548 (N_548,N_367,N_170);
or U549 (N_549,N_408,N_298);
xnor U550 (N_550,N_318,N_64);
or U551 (N_551,N_139,N_257);
nand U552 (N_552,N_154,N_137);
or U553 (N_553,N_404,N_337);
or U554 (N_554,N_227,N_278);
nor U555 (N_555,N_411,N_60);
nand U556 (N_556,N_405,N_182);
or U557 (N_557,N_230,N_56);
xnor U558 (N_558,N_191,N_43);
and U559 (N_559,N_39,N_423);
nand U560 (N_560,N_287,N_141);
and U561 (N_561,N_240,N_150);
nand U562 (N_562,N_70,N_118);
and U563 (N_563,N_447,N_17);
nand U564 (N_564,N_338,N_48);
nand U565 (N_565,N_348,N_82);
or U566 (N_566,N_172,N_46);
xor U567 (N_567,N_312,N_218);
or U568 (N_568,N_209,N_310);
nor U569 (N_569,N_63,N_387);
nand U570 (N_570,N_95,N_451);
or U571 (N_571,N_14,N_92);
and U572 (N_572,N_311,N_388);
and U573 (N_573,N_461,N_439);
or U574 (N_574,N_27,N_198);
or U575 (N_575,N_49,N_188);
or U576 (N_576,N_285,N_126);
and U577 (N_577,N_20,N_197);
nand U578 (N_578,N_228,N_75);
or U579 (N_579,N_301,N_32);
xor U580 (N_580,N_15,N_472);
nor U581 (N_581,N_97,N_442);
xnor U582 (N_582,N_340,N_317);
nand U583 (N_583,N_342,N_76);
nand U584 (N_584,N_238,N_104);
nand U585 (N_585,N_96,N_246);
and U586 (N_586,N_406,N_415);
xnor U587 (N_587,N_323,N_99);
and U588 (N_588,N_313,N_414);
nand U589 (N_589,N_326,N_292);
nor U590 (N_590,N_243,N_341);
or U591 (N_591,N_166,N_302);
nor U592 (N_592,N_125,N_430);
or U593 (N_593,N_87,N_382);
or U594 (N_594,N_62,N_111);
and U595 (N_595,N_116,N_320);
nor U596 (N_596,N_345,N_57);
or U597 (N_597,N_366,N_34);
and U598 (N_598,N_30,N_25);
xnor U599 (N_599,N_474,N_353);
or U600 (N_600,N_184,N_331);
nor U601 (N_601,N_339,N_215);
and U602 (N_602,N_252,N_53);
nand U603 (N_603,N_475,N_44);
nor U604 (N_604,N_145,N_390);
or U605 (N_605,N_122,N_113);
or U606 (N_606,N_303,N_289);
and U607 (N_607,N_253,N_418);
nor U608 (N_608,N_50,N_363);
and U609 (N_609,N_457,N_383);
and U610 (N_610,N_155,N_226);
or U611 (N_611,N_213,N_328);
xor U612 (N_612,N_394,N_274);
or U613 (N_613,N_66,N_81);
or U614 (N_614,N_362,N_171);
or U615 (N_615,N_350,N_417);
and U616 (N_616,N_214,N_454);
nor U617 (N_617,N_45,N_498);
and U618 (N_618,N_181,N_458);
and U619 (N_619,N_440,N_275);
or U620 (N_620,N_282,N_58);
and U621 (N_621,N_371,N_389);
or U622 (N_622,N_236,N_499);
nor U623 (N_623,N_144,N_107);
nor U624 (N_624,N_260,N_365);
nor U625 (N_625,N_224,N_24);
and U626 (N_626,N_361,N_429);
xnor U627 (N_627,N_147,N_158);
and U628 (N_628,N_419,N_65);
nand U629 (N_629,N_351,N_36);
and U630 (N_630,N_391,N_232);
or U631 (N_631,N_121,N_324);
nor U632 (N_632,N_159,N_470);
and U633 (N_633,N_157,N_464);
nand U634 (N_634,N_67,N_247);
nand U635 (N_635,N_61,N_165);
nand U636 (N_636,N_180,N_200);
xor U637 (N_637,N_346,N_378);
and U638 (N_638,N_374,N_91);
or U639 (N_639,N_349,N_321);
xnor U640 (N_640,N_175,N_399);
xor U641 (N_641,N_21,N_202);
nand U642 (N_642,N_148,N_2);
nand U643 (N_643,N_441,N_161);
or U644 (N_644,N_307,N_167);
nand U645 (N_645,N_433,N_124);
nor U646 (N_646,N_255,N_407);
and U647 (N_647,N_262,N_69);
nand U648 (N_648,N_86,N_245);
or U649 (N_649,N_201,N_384);
nand U650 (N_650,N_190,N_38);
and U651 (N_651,N_432,N_130);
and U652 (N_652,N_77,N_103);
nand U653 (N_653,N_434,N_131);
nor U654 (N_654,N_110,N_220);
nand U655 (N_655,N_413,N_133);
nand U656 (N_656,N_370,N_244);
and U657 (N_657,N_277,N_146);
nor U658 (N_658,N_73,N_268);
nand U659 (N_659,N_297,N_327);
or U660 (N_660,N_465,N_187);
xnor U661 (N_661,N_51,N_336);
xnor U662 (N_662,N_460,N_355);
and U663 (N_663,N_211,N_305);
nand U664 (N_664,N_487,N_481);
nand U665 (N_665,N_271,N_424);
nand U666 (N_666,N_235,N_489);
and U667 (N_667,N_140,N_193);
and U668 (N_668,N_88,N_286);
or U669 (N_669,N_335,N_207);
nor U670 (N_670,N_334,N_134);
and U671 (N_671,N_269,N_446);
nand U672 (N_672,N_479,N_250);
nand U673 (N_673,N_290,N_106);
or U674 (N_674,N_329,N_343);
nor U675 (N_675,N_0,N_9);
nand U676 (N_676,N_486,N_372);
and U677 (N_677,N_300,N_480);
nor U678 (N_678,N_233,N_54);
nor U679 (N_679,N_295,N_112);
nand U680 (N_680,N_35,N_283);
nor U681 (N_681,N_281,N_437);
or U682 (N_682,N_368,N_153);
nand U683 (N_683,N_19,N_473);
xnor U684 (N_684,N_272,N_108);
nor U685 (N_685,N_186,N_142);
or U686 (N_686,N_152,N_72);
nor U687 (N_687,N_299,N_352);
or U688 (N_688,N_293,N_71);
or U689 (N_689,N_239,N_291);
nor U690 (N_690,N_237,N_494);
nand U691 (N_691,N_354,N_332);
nand U692 (N_692,N_80,N_375);
nor U693 (N_693,N_306,N_431);
or U694 (N_694,N_169,N_373);
xnor U695 (N_695,N_493,N_120);
nor U696 (N_696,N_435,N_216);
and U697 (N_697,N_484,N_448);
and U698 (N_698,N_279,N_119);
and U699 (N_699,N_284,N_229);
nor U700 (N_700,N_151,N_94);
nor U701 (N_701,N_456,N_102);
nor U702 (N_702,N_234,N_196);
nand U703 (N_703,N_449,N_98);
and U704 (N_704,N_347,N_89);
nor U705 (N_705,N_385,N_496);
and U706 (N_706,N_225,N_231);
and U707 (N_707,N_138,N_10);
and U708 (N_708,N_4,N_1);
nor U709 (N_709,N_3,N_7);
or U710 (N_710,N_205,N_194);
nor U711 (N_711,N_222,N_393);
and U712 (N_712,N_314,N_248);
nand U713 (N_713,N_478,N_396);
xor U714 (N_714,N_490,N_445);
and U715 (N_715,N_308,N_90);
xnor U716 (N_716,N_78,N_270);
and U717 (N_717,N_403,N_203);
nand U718 (N_718,N_344,N_333);
nor U719 (N_719,N_400,N_392);
or U720 (N_720,N_288,N_476);
nor U721 (N_721,N_427,N_115);
nor U722 (N_722,N_109,N_273);
nor U723 (N_723,N_369,N_380);
nand U724 (N_724,N_174,N_195);
and U725 (N_725,N_402,N_241);
or U726 (N_726,N_428,N_469);
nand U727 (N_727,N_178,N_176);
nor U728 (N_728,N_177,N_47);
nor U729 (N_729,N_304,N_316);
nand U730 (N_730,N_453,N_249);
or U731 (N_731,N_13,N_416);
nor U732 (N_732,N_79,N_37);
and U733 (N_733,N_163,N_438);
or U734 (N_734,N_319,N_276);
nor U735 (N_735,N_294,N_136);
or U736 (N_736,N_5,N_52);
or U737 (N_737,N_93,N_221);
or U738 (N_738,N_471,N_74);
or U739 (N_739,N_325,N_410);
nor U740 (N_740,N_395,N_84);
nand U741 (N_741,N_128,N_491);
and U742 (N_742,N_265,N_401);
and U743 (N_743,N_185,N_477);
nand U744 (N_744,N_309,N_412);
or U745 (N_745,N_492,N_149);
nor U746 (N_746,N_68,N_183);
nor U747 (N_747,N_359,N_59);
and U748 (N_748,N_28,N_455);
and U749 (N_749,N_31,N_264);
nor U750 (N_750,N_107,N_280);
xnor U751 (N_751,N_218,N_202);
or U752 (N_752,N_37,N_315);
nand U753 (N_753,N_89,N_207);
xor U754 (N_754,N_20,N_30);
nor U755 (N_755,N_342,N_350);
nor U756 (N_756,N_8,N_397);
or U757 (N_757,N_38,N_54);
or U758 (N_758,N_275,N_226);
and U759 (N_759,N_163,N_462);
nor U760 (N_760,N_300,N_109);
or U761 (N_761,N_339,N_30);
and U762 (N_762,N_133,N_365);
and U763 (N_763,N_138,N_279);
nand U764 (N_764,N_65,N_102);
nand U765 (N_765,N_292,N_236);
or U766 (N_766,N_200,N_405);
nand U767 (N_767,N_75,N_242);
nand U768 (N_768,N_174,N_496);
or U769 (N_769,N_258,N_88);
nor U770 (N_770,N_421,N_301);
nor U771 (N_771,N_401,N_390);
nor U772 (N_772,N_77,N_1);
and U773 (N_773,N_43,N_399);
nor U774 (N_774,N_369,N_445);
nor U775 (N_775,N_201,N_446);
and U776 (N_776,N_432,N_400);
and U777 (N_777,N_102,N_471);
nor U778 (N_778,N_414,N_312);
nor U779 (N_779,N_342,N_290);
and U780 (N_780,N_419,N_68);
and U781 (N_781,N_307,N_214);
nand U782 (N_782,N_387,N_104);
and U783 (N_783,N_168,N_469);
nand U784 (N_784,N_382,N_315);
nand U785 (N_785,N_36,N_74);
nand U786 (N_786,N_54,N_390);
nand U787 (N_787,N_311,N_364);
nor U788 (N_788,N_42,N_280);
and U789 (N_789,N_401,N_376);
nand U790 (N_790,N_467,N_88);
nor U791 (N_791,N_2,N_183);
nor U792 (N_792,N_222,N_209);
nand U793 (N_793,N_323,N_0);
or U794 (N_794,N_274,N_195);
nor U795 (N_795,N_442,N_457);
and U796 (N_796,N_356,N_446);
nand U797 (N_797,N_62,N_488);
or U798 (N_798,N_421,N_440);
and U799 (N_799,N_225,N_112);
or U800 (N_800,N_136,N_191);
nor U801 (N_801,N_24,N_345);
or U802 (N_802,N_251,N_268);
and U803 (N_803,N_11,N_98);
or U804 (N_804,N_99,N_172);
or U805 (N_805,N_131,N_412);
or U806 (N_806,N_457,N_210);
nor U807 (N_807,N_182,N_175);
nand U808 (N_808,N_336,N_278);
xnor U809 (N_809,N_340,N_228);
nor U810 (N_810,N_222,N_25);
nand U811 (N_811,N_312,N_83);
nor U812 (N_812,N_109,N_217);
nor U813 (N_813,N_10,N_460);
nor U814 (N_814,N_185,N_66);
xor U815 (N_815,N_69,N_369);
xor U816 (N_816,N_233,N_362);
nand U817 (N_817,N_443,N_281);
and U818 (N_818,N_259,N_343);
nand U819 (N_819,N_366,N_356);
or U820 (N_820,N_431,N_264);
and U821 (N_821,N_380,N_61);
nor U822 (N_822,N_312,N_55);
and U823 (N_823,N_470,N_20);
xor U824 (N_824,N_452,N_344);
xor U825 (N_825,N_60,N_87);
or U826 (N_826,N_466,N_33);
nand U827 (N_827,N_144,N_6);
nor U828 (N_828,N_68,N_105);
and U829 (N_829,N_2,N_134);
nand U830 (N_830,N_156,N_63);
nand U831 (N_831,N_348,N_120);
nor U832 (N_832,N_466,N_65);
nor U833 (N_833,N_63,N_137);
or U834 (N_834,N_133,N_366);
xnor U835 (N_835,N_14,N_86);
or U836 (N_836,N_457,N_159);
and U837 (N_837,N_416,N_434);
or U838 (N_838,N_331,N_245);
nor U839 (N_839,N_457,N_236);
and U840 (N_840,N_66,N_77);
or U841 (N_841,N_190,N_232);
nor U842 (N_842,N_90,N_141);
nand U843 (N_843,N_485,N_462);
nand U844 (N_844,N_299,N_418);
or U845 (N_845,N_476,N_214);
or U846 (N_846,N_301,N_182);
nor U847 (N_847,N_137,N_177);
and U848 (N_848,N_269,N_175);
and U849 (N_849,N_181,N_163);
nand U850 (N_850,N_12,N_217);
nand U851 (N_851,N_234,N_430);
nand U852 (N_852,N_296,N_44);
and U853 (N_853,N_45,N_318);
nor U854 (N_854,N_395,N_120);
nand U855 (N_855,N_168,N_452);
nand U856 (N_856,N_198,N_115);
nor U857 (N_857,N_173,N_345);
and U858 (N_858,N_484,N_39);
nor U859 (N_859,N_184,N_333);
and U860 (N_860,N_109,N_222);
nor U861 (N_861,N_11,N_465);
nand U862 (N_862,N_450,N_482);
nor U863 (N_863,N_149,N_37);
or U864 (N_864,N_330,N_481);
nor U865 (N_865,N_411,N_378);
and U866 (N_866,N_492,N_285);
and U867 (N_867,N_316,N_105);
nor U868 (N_868,N_210,N_69);
nand U869 (N_869,N_202,N_155);
or U870 (N_870,N_241,N_401);
xnor U871 (N_871,N_171,N_436);
and U872 (N_872,N_162,N_144);
xnor U873 (N_873,N_67,N_465);
nor U874 (N_874,N_121,N_23);
nor U875 (N_875,N_371,N_498);
nand U876 (N_876,N_339,N_320);
nand U877 (N_877,N_236,N_184);
xnor U878 (N_878,N_428,N_434);
or U879 (N_879,N_403,N_373);
nand U880 (N_880,N_84,N_277);
or U881 (N_881,N_105,N_214);
nand U882 (N_882,N_290,N_125);
nand U883 (N_883,N_383,N_460);
and U884 (N_884,N_217,N_242);
xor U885 (N_885,N_390,N_335);
nand U886 (N_886,N_188,N_150);
nor U887 (N_887,N_215,N_450);
nor U888 (N_888,N_223,N_402);
and U889 (N_889,N_221,N_493);
or U890 (N_890,N_126,N_392);
nor U891 (N_891,N_3,N_283);
or U892 (N_892,N_423,N_42);
and U893 (N_893,N_236,N_125);
xor U894 (N_894,N_113,N_372);
xor U895 (N_895,N_484,N_173);
and U896 (N_896,N_112,N_303);
nor U897 (N_897,N_403,N_89);
and U898 (N_898,N_91,N_313);
or U899 (N_899,N_96,N_339);
or U900 (N_900,N_216,N_151);
xor U901 (N_901,N_66,N_140);
or U902 (N_902,N_67,N_188);
or U903 (N_903,N_165,N_3);
nand U904 (N_904,N_290,N_251);
or U905 (N_905,N_186,N_35);
or U906 (N_906,N_449,N_381);
nand U907 (N_907,N_10,N_349);
and U908 (N_908,N_409,N_379);
or U909 (N_909,N_132,N_325);
or U910 (N_910,N_474,N_286);
nand U911 (N_911,N_23,N_257);
nor U912 (N_912,N_267,N_312);
nor U913 (N_913,N_298,N_363);
or U914 (N_914,N_213,N_66);
and U915 (N_915,N_26,N_471);
or U916 (N_916,N_442,N_26);
xor U917 (N_917,N_210,N_431);
and U918 (N_918,N_397,N_330);
nor U919 (N_919,N_301,N_142);
or U920 (N_920,N_491,N_243);
and U921 (N_921,N_318,N_462);
nor U922 (N_922,N_261,N_268);
and U923 (N_923,N_190,N_130);
and U924 (N_924,N_337,N_12);
or U925 (N_925,N_34,N_344);
and U926 (N_926,N_498,N_125);
nand U927 (N_927,N_151,N_469);
xnor U928 (N_928,N_345,N_59);
or U929 (N_929,N_165,N_50);
and U930 (N_930,N_223,N_384);
nand U931 (N_931,N_420,N_435);
nand U932 (N_932,N_251,N_276);
nor U933 (N_933,N_419,N_478);
and U934 (N_934,N_440,N_298);
nand U935 (N_935,N_340,N_356);
nand U936 (N_936,N_493,N_301);
or U937 (N_937,N_432,N_46);
and U938 (N_938,N_103,N_147);
or U939 (N_939,N_165,N_140);
xnor U940 (N_940,N_107,N_478);
xnor U941 (N_941,N_446,N_380);
nand U942 (N_942,N_21,N_449);
nand U943 (N_943,N_280,N_418);
nand U944 (N_944,N_264,N_415);
or U945 (N_945,N_303,N_64);
and U946 (N_946,N_460,N_375);
nor U947 (N_947,N_77,N_460);
and U948 (N_948,N_407,N_122);
and U949 (N_949,N_447,N_74);
xor U950 (N_950,N_44,N_382);
and U951 (N_951,N_280,N_34);
nand U952 (N_952,N_483,N_346);
xnor U953 (N_953,N_350,N_303);
and U954 (N_954,N_294,N_207);
nor U955 (N_955,N_454,N_293);
and U956 (N_956,N_192,N_215);
nor U957 (N_957,N_463,N_443);
nand U958 (N_958,N_118,N_313);
nor U959 (N_959,N_119,N_272);
or U960 (N_960,N_399,N_480);
and U961 (N_961,N_449,N_9);
or U962 (N_962,N_424,N_45);
and U963 (N_963,N_339,N_440);
and U964 (N_964,N_45,N_9);
or U965 (N_965,N_49,N_106);
nand U966 (N_966,N_295,N_408);
or U967 (N_967,N_164,N_202);
nand U968 (N_968,N_282,N_183);
and U969 (N_969,N_463,N_385);
nor U970 (N_970,N_75,N_455);
and U971 (N_971,N_374,N_350);
nand U972 (N_972,N_376,N_461);
nand U973 (N_973,N_116,N_494);
nand U974 (N_974,N_382,N_158);
and U975 (N_975,N_341,N_496);
nand U976 (N_976,N_281,N_440);
or U977 (N_977,N_60,N_133);
and U978 (N_978,N_307,N_439);
or U979 (N_979,N_383,N_49);
nor U980 (N_980,N_356,N_307);
xor U981 (N_981,N_392,N_475);
or U982 (N_982,N_131,N_351);
or U983 (N_983,N_458,N_152);
or U984 (N_984,N_435,N_64);
and U985 (N_985,N_306,N_445);
nor U986 (N_986,N_482,N_352);
or U987 (N_987,N_148,N_349);
nor U988 (N_988,N_93,N_210);
xor U989 (N_989,N_298,N_259);
xnor U990 (N_990,N_43,N_159);
and U991 (N_991,N_498,N_408);
or U992 (N_992,N_392,N_422);
nand U993 (N_993,N_463,N_205);
and U994 (N_994,N_410,N_103);
and U995 (N_995,N_478,N_180);
or U996 (N_996,N_133,N_410);
nand U997 (N_997,N_101,N_358);
xnor U998 (N_998,N_287,N_221);
or U999 (N_999,N_465,N_229);
nor U1000 (N_1000,N_690,N_989);
or U1001 (N_1001,N_915,N_651);
and U1002 (N_1002,N_772,N_947);
or U1003 (N_1003,N_673,N_624);
xnor U1004 (N_1004,N_940,N_896);
or U1005 (N_1005,N_903,N_842);
or U1006 (N_1006,N_794,N_710);
nand U1007 (N_1007,N_613,N_824);
or U1008 (N_1008,N_725,N_751);
xnor U1009 (N_1009,N_600,N_758);
nor U1010 (N_1010,N_978,N_693);
and U1011 (N_1011,N_942,N_788);
or U1012 (N_1012,N_713,N_771);
nand U1013 (N_1013,N_700,N_535);
nor U1014 (N_1014,N_546,N_987);
and U1015 (N_1015,N_962,N_626);
and U1016 (N_1016,N_573,N_707);
nor U1017 (N_1017,N_506,N_729);
and U1018 (N_1018,N_877,N_657);
xor U1019 (N_1019,N_930,N_647);
or U1020 (N_1020,N_604,N_872);
nor U1021 (N_1021,N_599,N_721);
nand U1022 (N_1022,N_649,N_765);
and U1023 (N_1023,N_584,N_924);
nor U1024 (N_1024,N_534,N_752);
or U1025 (N_1025,N_681,N_910);
nor U1026 (N_1026,N_526,N_868);
nand U1027 (N_1027,N_997,N_652);
nand U1028 (N_1028,N_735,N_509);
xnor U1029 (N_1029,N_577,N_938);
xor U1030 (N_1030,N_741,N_922);
nor U1031 (N_1031,N_750,N_780);
and U1032 (N_1032,N_553,N_988);
nand U1033 (N_1033,N_799,N_656);
nand U1034 (N_1034,N_547,N_542);
and U1035 (N_1035,N_668,N_928);
and U1036 (N_1036,N_691,N_897);
or U1037 (N_1037,N_504,N_986);
nand U1038 (N_1038,N_871,N_723);
or U1039 (N_1039,N_636,N_782);
and U1040 (N_1040,N_863,N_538);
or U1041 (N_1041,N_798,N_909);
and U1042 (N_1042,N_831,N_703);
xor U1043 (N_1043,N_557,N_807);
and U1044 (N_1044,N_620,N_802);
nand U1045 (N_1045,N_929,N_778);
nor U1046 (N_1046,N_718,N_839);
or U1047 (N_1047,N_753,N_914);
or U1048 (N_1048,N_679,N_687);
nand U1049 (N_1049,N_843,N_611);
xor U1050 (N_1050,N_976,N_932);
and U1051 (N_1051,N_822,N_738);
or U1052 (N_1052,N_663,N_812);
or U1053 (N_1053,N_856,N_826);
xnor U1054 (N_1054,N_916,N_682);
or U1055 (N_1055,N_724,N_887);
and U1056 (N_1056,N_874,N_904);
and U1057 (N_1057,N_792,N_888);
nand U1058 (N_1058,N_803,N_737);
and U1059 (N_1059,N_736,N_530);
or U1060 (N_1060,N_879,N_745);
or U1061 (N_1061,N_865,N_572);
or U1062 (N_1062,N_776,N_519);
xor U1063 (N_1063,N_576,N_770);
nand U1064 (N_1064,N_800,N_943);
nor U1065 (N_1065,N_715,N_632);
nor U1066 (N_1066,N_590,N_789);
nor U1067 (N_1067,N_864,N_653);
nor U1068 (N_1068,N_979,N_827);
and U1069 (N_1069,N_983,N_834);
nor U1070 (N_1070,N_701,N_844);
or U1071 (N_1071,N_621,N_622);
nor U1072 (N_1072,N_804,N_764);
xor U1073 (N_1073,N_775,N_501);
nand U1074 (N_1074,N_810,N_511);
xor U1075 (N_1075,N_541,N_708);
nand U1076 (N_1076,N_667,N_610);
nor U1077 (N_1077,N_912,N_680);
xnor U1078 (N_1078,N_855,N_763);
nor U1079 (N_1079,N_591,N_515);
and U1080 (N_1080,N_769,N_974);
or U1081 (N_1081,N_537,N_985);
xor U1082 (N_1082,N_523,N_975);
and U1083 (N_1083,N_766,N_900);
or U1084 (N_1084,N_968,N_637);
or U1085 (N_1085,N_934,N_823);
nor U1086 (N_1086,N_650,N_671);
nand U1087 (N_1087,N_586,N_953);
or U1088 (N_1088,N_734,N_966);
nor U1089 (N_1089,N_993,N_786);
and U1090 (N_1090,N_588,N_555);
and U1091 (N_1091,N_919,N_532);
and U1092 (N_1092,N_956,N_744);
and U1093 (N_1093,N_779,N_732);
or U1094 (N_1094,N_528,N_890);
and U1095 (N_1095,N_911,N_818);
nor U1096 (N_1096,N_731,N_961);
or U1097 (N_1097,N_992,N_609);
nand U1098 (N_1098,N_683,N_500);
nor U1099 (N_1099,N_664,N_574);
nand U1100 (N_1100,N_615,N_793);
nor U1101 (N_1101,N_935,N_702);
nand U1102 (N_1102,N_579,N_633);
and U1103 (N_1103,N_561,N_832);
or U1104 (N_1104,N_524,N_845);
and U1105 (N_1105,N_920,N_655);
or U1106 (N_1106,N_630,N_562);
xnor U1107 (N_1107,N_836,N_891);
nand U1108 (N_1108,N_939,N_892);
or U1109 (N_1109,N_767,N_881);
nand U1110 (N_1110,N_949,N_886);
xor U1111 (N_1111,N_642,N_885);
and U1112 (N_1112,N_560,N_848);
nor U1113 (N_1113,N_805,N_720);
xor U1114 (N_1114,N_659,N_631);
and U1115 (N_1115,N_840,N_616);
or U1116 (N_1116,N_774,N_952);
nor U1117 (N_1117,N_869,N_847);
nor U1118 (N_1118,N_944,N_955);
nor U1119 (N_1119,N_899,N_518);
or U1120 (N_1120,N_617,N_905);
nor U1121 (N_1121,N_882,N_685);
nor U1122 (N_1122,N_739,N_578);
or U1123 (N_1123,N_996,N_684);
nand U1124 (N_1124,N_627,N_699);
nand U1125 (N_1125,N_984,N_596);
and U1126 (N_1126,N_913,N_921);
nand U1127 (N_1127,N_565,N_605);
and U1128 (N_1128,N_754,N_704);
nand U1129 (N_1129,N_566,N_665);
or U1130 (N_1130,N_925,N_846);
nand U1131 (N_1131,N_876,N_815);
or U1132 (N_1132,N_821,N_759);
or U1133 (N_1133,N_806,N_757);
or U1134 (N_1134,N_606,N_790);
or U1135 (N_1135,N_743,N_851);
nor U1136 (N_1136,N_918,N_850);
nor U1137 (N_1137,N_728,N_860);
and U1138 (N_1138,N_862,N_858);
and U1139 (N_1139,N_536,N_884);
nor U1140 (N_1140,N_677,N_873);
nand U1141 (N_1141,N_933,N_648);
and U1142 (N_1142,N_706,N_958);
and U1143 (N_1143,N_705,N_973);
or U1144 (N_1144,N_517,N_676);
and U1145 (N_1145,N_575,N_817);
and U1146 (N_1146,N_960,N_880);
or U1147 (N_1147,N_959,N_623);
and U1148 (N_1148,N_520,N_835);
xnor U1149 (N_1149,N_522,N_963);
nand U1150 (N_1150,N_867,N_601);
nor U1151 (N_1151,N_946,N_964);
nand U1152 (N_1152,N_990,N_908);
and U1153 (N_1153,N_999,N_889);
nand U1154 (N_1154,N_580,N_977);
nand U1155 (N_1155,N_998,N_625);
nand U1156 (N_1156,N_917,N_503);
xor U1157 (N_1157,N_556,N_995);
xor U1158 (N_1158,N_854,N_628);
nor U1159 (N_1159,N_597,N_670);
and U1160 (N_1160,N_666,N_982);
or U1161 (N_1161,N_678,N_957);
and U1162 (N_1162,N_830,N_781);
or U1163 (N_1163,N_857,N_711);
and U1164 (N_1164,N_994,N_635);
and U1165 (N_1165,N_797,N_505);
nor U1166 (N_1166,N_583,N_969);
nor U1167 (N_1167,N_548,N_747);
xnor U1168 (N_1168,N_714,N_618);
or U1169 (N_1169,N_608,N_849);
or U1170 (N_1170,N_569,N_967);
nand U1171 (N_1171,N_722,N_571);
nand U1172 (N_1172,N_951,N_748);
or U1173 (N_1173,N_712,N_733);
nand U1174 (N_1174,N_950,N_593);
nand U1175 (N_1175,N_695,N_820);
and U1176 (N_1176,N_638,N_893);
nor U1177 (N_1177,N_598,N_948);
or U1178 (N_1178,N_906,N_746);
nand U1179 (N_1179,N_540,N_761);
or U1180 (N_1180,N_602,N_740);
nor U1181 (N_1181,N_841,N_833);
and U1182 (N_1182,N_658,N_531);
and U1183 (N_1183,N_672,N_589);
and U1184 (N_1184,N_612,N_936);
nor U1185 (N_1185,N_660,N_965);
and U1186 (N_1186,N_727,N_694);
nand U1187 (N_1187,N_716,N_785);
xor U1188 (N_1188,N_895,N_927);
nand U1189 (N_1189,N_829,N_883);
nand U1190 (N_1190,N_742,N_641);
and U1191 (N_1191,N_756,N_603);
or U1192 (N_1192,N_796,N_816);
and U1193 (N_1193,N_545,N_634);
or U1194 (N_1194,N_582,N_931);
or U1195 (N_1195,N_549,N_502);
nand U1196 (N_1196,N_675,N_558);
nor U1197 (N_1197,N_859,N_595);
nor U1198 (N_1198,N_811,N_688);
nand U1199 (N_1199,N_592,N_514);
nand U1200 (N_1200,N_581,N_870);
and U1201 (N_1201,N_825,N_525);
nor U1202 (N_1202,N_991,N_550);
nand U1203 (N_1203,N_941,N_760);
or U1204 (N_1204,N_878,N_837);
and U1205 (N_1205,N_539,N_686);
xor U1206 (N_1206,N_972,N_801);
and U1207 (N_1207,N_762,N_644);
nand U1208 (N_1208,N_901,N_814);
or U1209 (N_1209,N_981,N_563);
nand U1210 (N_1210,N_689,N_838);
nor U1211 (N_1211,N_567,N_508);
nand U1212 (N_1212,N_866,N_937);
and U1213 (N_1213,N_510,N_852);
and U1214 (N_1214,N_777,N_551);
nand U1215 (N_1215,N_980,N_730);
xor U1216 (N_1216,N_614,N_512);
nor U1217 (N_1217,N_692,N_587);
nand U1218 (N_1218,N_619,N_813);
and U1219 (N_1219,N_945,N_926);
nand U1220 (N_1220,N_654,N_507);
or U1221 (N_1221,N_521,N_585);
and U1222 (N_1222,N_828,N_568);
nand U1223 (N_1223,N_923,N_697);
or U1224 (N_1224,N_554,N_787);
nand U1225 (N_1225,N_552,N_898);
nor U1226 (N_1226,N_564,N_533);
nand U1227 (N_1227,N_809,N_795);
nand U1228 (N_1228,N_768,N_894);
nor U1229 (N_1229,N_559,N_674);
nor U1230 (N_1230,N_662,N_819);
and U1231 (N_1231,N_544,N_516);
xor U1232 (N_1232,N_629,N_594);
nand U1233 (N_1233,N_902,N_709);
nor U1234 (N_1234,N_749,N_719);
nor U1235 (N_1235,N_543,N_527);
nor U1236 (N_1236,N_784,N_773);
or U1237 (N_1237,N_970,N_717);
nand U1238 (N_1238,N_971,N_639);
nand U1239 (N_1239,N_513,N_726);
nor U1240 (N_1240,N_783,N_755);
or U1241 (N_1241,N_954,N_808);
nor U1242 (N_1242,N_861,N_698);
nand U1243 (N_1243,N_669,N_607);
nor U1244 (N_1244,N_646,N_645);
nand U1245 (N_1245,N_853,N_661);
nand U1246 (N_1246,N_529,N_791);
nand U1247 (N_1247,N_696,N_643);
and U1248 (N_1248,N_907,N_640);
nor U1249 (N_1249,N_875,N_570);
and U1250 (N_1250,N_521,N_898);
or U1251 (N_1251,N_997,N_639);
nor U1252 (N_1252,N_717,N_732);
and U1253 (N_1253,N_867,N_905);
and U1254 (N_1254,N_942,N_995);
nor U1255 (N_1255,N_809,N_734);
and U1256 (N_1256,N_743,N_986);
nor U1257 (N_1257,N_632,N_519);
or U1258 (N_1258,N_730,N_981);
nand U1259 (N_1259,N_648,N_749);
and U1260 (N_1260,N_730,N_673);
xnor U1261 (N_1261,N_763,N_843);
and U1262 (N_1262,N_517,N_736);
nand U1263 (N_1263,N_708,N_996);
nor U1264 (N_1264,N_918,N_697);
and U1265 (N_1265,N_585,N_779);
nand U1266 (N_1266,N_645,N_859);
nand U1267 (N_1267,N_657,N_892);
and U1268 (N_1268,N_974,N_829);
xnor U1269 (N_1269,N_674,N_856);
nor U1270 (N_1270,N_824,N_614);
or U1271 (N_1271,N_902,N_868);
nor U1272 (N_1272,N_913,N_911);
xor U1273 (N_1273,N_770,N_505);
or U1274 (N_1274,N_662,N_899);
nand U1275 (N_1275,N_879,N_840);
and U1276 (N_1276,N_656,N_528);
nand U1277 (N_1277,N_683,N_754);
and U1278 (N_1278,N_621,N_741);
and U1279 (N_1279,N_616,N_584);
nand U1280 (N_1280,N_572,N_757);
and U1281 (N_1281,N_665,N_745);
nand U1282 (N_1282,N_940,N_904);
xnor U1283 (N_1283,N_739,N_692);
or U1284 (N_1284,N_968,N_744);
or U1285 (N_1285,N_582,N_886);
nand U1286 (N_1286,N_977,N_508);
or U1287 (N_1287,N_675,N_597);
nor U1288 (N_1288,N_999,N_690);
or U1289 (N_1289,N_549,N_774);
xor U1290 (N_1290,N_937,N_998);
and U1291 (N_1291,N_618,N_734);
and U1292 (N_1292,N_636,N_926);
or U1293 (N_1293,N_777,N_891);
nor U1294 (N_1294,N_833,N_760);
nand U1295 (N_1295,N_985,N_865);
nor U1296 (N_1296,N_613,N_623);
and U1297 (N_1297,N_607,N_573);
or U1298 (N_1298,N_817,N_932);
nand U1299 (N_1299,N_862,N_952);
nand U1300 (N_1300,N_617,N_553);
or U1301 (N_1301,N_508,N_823);
or U1302 (N_1302,N_586,N_823);
and U1303 (N_1303,N_581,N_975);
and U1304 (N_1304,N_516,N_583);
and U1305 (N_1305,N_913,N_519);
or U1306 (N_1306,N_765,N_950);
or U1307 (N_1307,N_601,N_577);
nand U1308 (N_1308,N_592,N_934);
nand U1309 (N_1309,N_881,N_841);
nand U1310 (N_1310,N_788,N_902);
nand U1311 (N_1311,N_531,N_953);
or U1312 (N_1312,N_510,N_694);
nor U1313 (N_1313,N_714,N_914);
nor U1314 (N_1314,N_866,N_806);
and U1315 (N_1315,N_712,N_519);
xnor U1316 (N_1316,N_725,N_577);
and U1317 (N_1317,N_659,N_630);
or U1318 (N_1318,N_926,N_674);
nor U1319 (N_1319,N_794,N_861);
nor U1320 (N_1320,N_670,N_844);
nor U1321 (N_1321,N_549,N_850);
nor U1322 (N_1322,N_528,N_786);
nand U1323 (N_1323,N_809,N_804);
or U1324 (N_1324,N_673,N_685);
and U1325 (N_1325,N_682,N_608);
nor U1326 (N_1326,N_938,N_610);
or U1327 (N_1327,N_754,N_648);
nand U1328 (N_1328,N_923,N_573);
and U1329 (N_1329,N_770,N_926);
or U1330 (N_1330,N_698,N_643);
and U1331 (N_1331,N_791,N_572);
nor U1332 (N_1332,N_678,N_966);
or U1333 (N_1333,N_631,N_833);
and U1334 (N_1334,N_596,N_826);
and U1335 (N_1335,N_983,N_667);
or U1336 (N_1336,N_842,N_990);
nand U1337 (N_1337,N_523,N_710);
or U1338 (N_1338,N_644,N_549);
and U1339 (N_1339,N_631,N_673);
and U1340 (N_1340,N_551,N_690);
or U1341 (N_1341,N_940,N_586);
or U1342 (N_1342,N_984,N_619);
nor U1343 (N_1343,N_919,N_560);
or U1344 (N_1344,N_667,N_566);
nor U1345 (N_1345,N_817,N_893);
nand U1346 (N_1346,N_690,N_762);
nand U1347 (N_1347,N_850,N_962);
or U1348 (N_1348,N_654,N_906);
nand U1349 (N_1349,N_540,N_976);
and U1350 (N_1350,N_654,N_736);
or U1351 (N_1351,N_758,N_902);
xnor U1352 (N_1352,N_637,N_681);
or U1353 (N_1353,N_766,N_720);
and U1354 (N_1354,N_727,N_767);
and U1355 (N_1355,N_555,N_568);
and U1356 (N_1356,N_653,N_724);
nor U1357 (N_1357,N_545,N_978);
or U1358 (N_1358,N_749,N_766);
nand U1359 (N_1359,N_943,N_737);
nand U1360 (N_1360,N_967,N_697);
nand U1361 (N_1361,N_885,N_826);
and U1362 (N_1362,N_986,N_683);
nand U1363 (N_1363,N_633,N_612);
nor U1364 (N_1364,N_527,N_630);
and U1365 (N_1365,N_949,N_531);
or U1366 (N_1366,N_931,N_861);
xnor U1367 (N_1367,N_736,N_641);
nor U1368 (N_1368,N_679,N_937);
nor U1369 (N_1369,N_621,N_974);
or U1370 (N_1370,N_567,N_745);
nand U1371 (N_1371,N_729,N_605);
nand U1372 (N_1372,N_710,N_657);
or U1373 (N_1373,N_828,N_617);
and U1374 (N_1374,N_738,N_955);
and U1375 (N_1375,N_931,N_712);
or U1376 (N_1376,N_828,N_879);
and U1377 (N_1377,N_541,N_638);
and U1378 (N_1378,N_577,N_929);
nor U1379 (N_1379,N_782,N_634);
or U1380 (N_1380,N_872,N_770);
and U1381 (N_1381,N_902,N_523);
or U1382 (N_1382,N_568,N_563);
nand U1383 (N_1383,N_858,N_760);
or U1384 (N_1384,N_796,N_942);
nand U1385 (N_1385,N_808,N_605);
xor U1386 (N_1386,N_708,N_864);
or U1387 (N_1387,N_753,N_822);
nor U1388 (N_1388,N_624,N_905);
or U1389 (N_1389,N_583,N_671);
nor U1390 (N_1390,N_585,N_869);
and U1391 (N_1391,N_600,N_510);
nor U1392 (N_1392,N_667,N_999);
nand U1393 (N_1393,N_765,N_988);
nor U1394 (N_1394,N_592,N_972);
or U1395 (N_1395,N_711,N_921);
or U1396 (N_1396,N_797,N_960);
xnor U1397 (N_1397,N_840,N_567);
or U1398 (N_1398,N_611,N_844);
or U1399 (N_1399,N_958,N_957);
or U1400 (N_1400,N_593,N_955);
or U1401 (N_1401,N_798,N_889);
nor U1402 (N_1402,N_522,N_819);
and U1403 (N_1403,N_830,N_661);
xor U1404 (N_1404,N_568,N_594);
nand U1405 (N_1405,N_697,N_830);
nand U1406 (N_1406,N_735,N_879);
nand U1407 (N_1407,N_761,N_644);
or U1408 (N_1408,N_972,N_674);
nand U1409 (N_1409,N_567,N_852);
xnor U1410 (N_1410,N_733,N_568);
nand U1411 (N_1411,N_872,N_549);
and U1412 (N_1412,N_550,N_920);
and U1413 (N_1413,N_686,N_622);
nand U1414 (N_1414,N_942,N_734);
xnor U1415 (N_1415,N_971,N_993);
or U1416 (N_1416,N_869,N_992);
nand U1417 (N_1417,N_626,N_875);
or U1418 (N_1418,N_735,N_682);
and U1419 (N_1419,N_559,N_650);
and U1420 (N_1420,N_977,N_627);
nand U1421 (N_1421,N_666,N_842);
or U1422 (N_1422,N_648,N_929);
and U1423 (N_1423,N_768,N_856);
nand U1424 (N_1424,N_914,N_631);
or U1425 (N_1425,N_940,N_918);
nor U1426 (N_1426,N_601,N_694);
nor U1427 (N_1427,N_513,N_607);
or U1428 (N_1428,N_677,N_688);
and U1429 (N_1429,N_824,N_547);
nor U1430 (N_1430,N_813,N_984);
nor U1431 (N_1431,N_660,N_753);
nand U1432 (N_1432,N_946,N_716);
and U1433 (N_1433,N_524,N_683);
and U1434 (N_1434,N_960,N_652);
xor U1435 (N_1435,N_857,N_909);
nor U1436 (N_1436,N_828,N_822);
nor U1437 (N_1437,N_561,N_536);
and U1438 (N_1438,N_955,N_830);
nor U1439 (N_1439,N_918,N_644);
xor U1440 (N_1440,N_667,N_699);
nand U1441 (N_1441,N_980,N_558);
or U1442 (N_1442,N_954,N_793);
or U1443 (N_1443,N_938,N_652);
and U1444 (N_1444,N_858,N_814);
and U1445 (N_1445,N_898,N_571);
or U1446 (N_1446,N_525,N_959);
or U1447 (N_1447,N_604,N_923);
nand U1448 (N_1448,N_547,N_647);
nand U1449 (N_1449,N_621,N_876);
xnor U1450 (N_1450,N_675,N_575);
or U1451 (N_1451,N_703,N_661);
and U1452 (N_1452,N_717,N_878);
nand U1453 (N_1453,N_530,N_563);
xnor U1454 (N_1454,N_750,N_834);
or U1455 (N_1455,N_511,N_827);
or U1456 (N_1456,N_845,N_659);
or U1457 (N_1457,N_564,N_629);
or U1458 (N_1458,N_725,N_808);
xnor U1459 (N_1459,N_962,N_693);
nand U1460 (N_1460,N_706,N_897);
and U1461 (N_1461,N_697,N_964);
and U1462 (N_1462,N_780,N_596);
nor U1463 (N_1463,N_528,N_955);
and U1464 (N_1464,N_885,N_512);
xnor U1465 (N_1465,N_694,N_551);
nand U1466 (N_1466,N_601,N_542);
or U1467 (N_1467,N_557,N_951);
nor U1468 (N_1468,N_541,N_821);
nand U1469 (N_1469,N_883,N_919);
xor U1470 (N_1470,N_897,N_657);
and U1471 (N_1471,N_719,N_961);
nand U1472 (N_1472,N_676,N_600);
xor U1473 (N_1473,N_596,N_777);
nor U1474 (N_1474,N_887,N_622);
and U1475 (N_1475,N_750,N_807);
nand U1476 (N_1476,N_736,N_843);
nor U1477 (N_1477,N_953,N_517);
or U1478 (N_1478,N_926,N_850);
nor U1479 (N_1479,N_728,N_751);
and U1480 (N_1480,N_739,N_976);
or U1481 (N_1481,N_768,N_726);
nand U1482 (N_1482,N_917,N_918);
nand U1483 (N_1483,N_831,N_721);
nand U1484 (N_1484,N_581,N_938);
or U1485 (N_1485,N_744,N_947);
and U1486 (N_1486,N_617,N_928);
nand U1487 (N_1487,N_848,N_792);
or U1488 (N_1488,N_703,N_750);
nand U1489 (N_1489,N_665,N_971);
nor U1490 (N_1490,N_515,N_848);
or U1491 (N_1491,N_879,N_744);
xor U1492 (N_1492,N_550,N_681);
xnor U1493 (N_1493,N_932,N_873);
xnor U1494 (N_1494,N_553,N_872);
nor U1495 (N_1495,N_807,N_543);
xor U1496 (N_1496,N_762,N_993);
nor U1497 (N_1497,N_589,N_514);
nor U1498 (N_1498,N_761,N_643);
and U1499 (N_1499,N_529,N_543);
or U1500 (N_1500,N_1374,N_1159);
or U1501 (N_1501,N_1312,N_1129);
and U1502 (N_1502,N_1424,N_1400);
nand U1503 (N_1503,N_1082,N_1363);
nor U1504 (N_1504,N_1409,N_1151);
xnor U1505 (N_1505,N_1176,N_1279);
or U1506 (N_1506,N_1496,N_1283);
nand U1507 (N_1507,N_1354,N_1055);
or U1508 (N_1508,N_1124,N_1138);
nand U1509 (N_1509,N_1019,N_1073);
xnor U1510 (N_1510,N_1321,N_1278);
and U1511 (N_1511,N_1222,N_1047);
nor U1512 (N_1512,N_1095,N_1116);
xor U1513 (N_1513,N_1032,N_1280);
xnor U1514 (N_1514,N_1296,N_1271);
and U1515 (N_1515,N_1075,N_1240);
or U1516 (N_1516,N_1391,N_1269);
nand U1517 (N_1517,N_1200,N_1437);
nor U1518 (N_1518,N_1265,N_1253);
nor U1519 (N_1519,N_1356,N_1315);
nor U1520 (N_1520,N_1066,N_1079);
nor U1521 (N_1521,N_1475,N_1173);
nor U1522 (N_1522,N_1347,N_1218);
or U1523 (N_1523,N_1247,N_1262);
nand U1524 (N_1524,N_1168,N_1130);
nor U1525 (N_1525,N_1489,N_1167);
xor U1526 (N_1526,N_1304,N_1494);
nor U1527 (N_1527,N_1087,N_1461);
and U1528 (N_1528,N_1418,N_1195);
nor U1529 (N_1529,N_1171,N_1415);
or U1530 (N_1530,N_1027,N_1157);
nor U1531 (N_1531,N_1086,N_1408);
and U1532 (N_1532,N_1015,N_1012);
and U1533 (N_1533,N_1219,N_1038);
and U1534 (N_1534,N_1479,N_1263);
or U1535 (N_1535,N_1028,N_1045);
and U1536 (N_1536,N_1360,N_1237);
and U1537 (N_1537,N_1314,N_1266);
nor U1538 (N_1538,N_1110,N_1106);
nor U1539 (N_1539,N_1215,N_1049);
and U1540 (N_1540,N_1302,N_1146);
nor U1541 (N_1541,N_1319,N_1348);
nand U1542 (N_1542,N_1270,N_1371);
or U1543 (N_1543,N_1036,N_1022);
nand U1544 (N_1544,N_1472,N_1212);
and U1545 (N_1545,N_1272,N_1490);
and U1546 (N_1546,N_1076,N_1465);
and U1547 (N_1547,N_1469,N_1425);
or U1548 (N_1548,N_1459,N_1034);
nand U1549 (N_1549,N_1037,N_1099);
nand U1550 (N_1550,N_1333,N_1048);
or U1551 (N_1551,N_1261,N_1370);
and U1552 (N_1552,N_1142,N_1120);
xor U1553 (N_1553,N_1414,N_1096);
xor U1554 (N_1554,N_1382,N_1202);
xnor U1555 (N_1555,N_1063,N_1236);
nor U1556 (N_1556,N_1350,N_1405);
nand U1557 (N_1557,N_1131,N_1104);
and U1558 (N_1558,N_1463,N_1401);
and U1559 (N_1559,N_1089,N_1144);
xnor U1560 (N_1560,N_1125,N_1232);
and U1561 (N_1561,N_1477,N_1207);
nor U1562 (N_1562,N_1325,N_1123);
xor U1563 (N_1563,N_1478,N_1121);
or U1564 (N_1564,N_1362,N_1018);
xnor U1565 (N_1565,N_1072,N_1188);
nand U1566 (N_1566,N_1085,N_1389);
nand U1567 (N_1567,N_1118,N_1198);
nand U1568 (N_1568,N_1134,N_1115);
or U1569 (N_1569,N_1326,N_1238);
nor U1570 (N_1570,N_1090,N_1139);
and U1571 (N_1571,N_1070,N_1416);
or U1572 (N_1572,N_1064,N_1242);
nand U1573 (N_1573,N_1373,N_1054);
xor U1574 (N_1574,N_1381,N_1339);
nand U1575 (N_1575,N_1349,N_1396);
or U1576 (N_1576,N_1052,N_1248);
nand U1577 (N_1577,N_1482,N_1030);
and U1578 (N_1578,N_1281,N_1344);
and U1579 (N_1579,N_1456,N_1295);
nor U1580 (N_1580,N_1084,N_1119);
nor U1581 (N_1581,N_1403,N_1254);
nand U1582 (N_1582,N_1336,N_1031);
or U1583 (N_1583,N_1448,N_1444);
nand U1584 (N_1584,N_1107,N_1343);
and U1585 (N_1585,N_1203,N_1141);
nor U1586 (N_1586,N_1259,N_1290);
nor U1587 (N_1587,N_1431,N_1361);
or U1588 (N_1588,N_1040,N_1402);
nor U1589 (N_1589,N_1136,N_1029);
nand U1590 (N_1590,N_1397,N_1108);
and U1591 (N_1591,N_1065,N_1282);
xnor U1592 (N_1592,N_1446,N_1256);
or U1593 (N_1593,N_1398,N_1100);
or U1594 (N_1594,N_1308,N_1005);
or U1595 (N_1595,N_1340,N_1033);
and U1596 (N_1596,N_1094,N_1150);
nand U1597 (N_1597,N_1183,N_1193);
or U1598 (N_1598,N_1413,N_1365);
or U1599 (N_1599,N_1467,N_1154);
and U1600 (N_1600,N_1187,N_1208);
and U1601 (N_1601,N_1433,N_1322);
and U1602 (N_1602,N_1145,N_1069);
nor U1603 (N_1603,N_1196,N_1334);
nand U1604 (N_1604,N_1423,N_1216);
nand U1605 (N_1605,N_1491,N_1149);
and U1606 (N_1606,N_1239,N_1303);
and U1607 (N_1607,N_1367,N_1024);
nor U1608 (N_1608,N_1293,N_1455);
and U1609 (N_1609,N_1417,N_1184);
nand U1610 (N_1610,N_1481,N_1345);
nor U1611 (N_1611,N_1013,N_1376);
and U1612 (N_1612,N_1229,N_1352);
nand U1613 (N_1613,N_1080,N_1231);
or U1614 (N_1614,N_1411,N_1039);
xor U1615 (N_1615,N_1499,N_1143);
or U1616 (N_1616,N_1379,N_1386);
nor U1617 (N_1617,N_1014,N_1109);
or U1618 (N_1618,N_1436,N_1017);
and U1619 (N_1619,N_1488,N_1434);
and U1620 (N_1620,N_1117,N_1058);
or U1621 (N_1621,N_1174,N_1466);
nand U1622 (N_1622,N_1162,N_1179);
nand U1623 (N_1623,N_1378,N_1355);
xnor U1624 (N_1624,N_1211,N_1357);
or U1625 (N_1625,N_1163,N_1480);
or U1626 (N_1626,N_1227,N_1166);
nor U1627 (N_1627,N_1074,N_1369);
xnor U1628 (N_1628,N_1288,N_1061);
or U1629 (N_1629,N_1358,N_1335);
nand U1630 (N_1630,N_1009,N_1368);
or U1631 (N_1631,N_1301,N_1449);
nand U1632 (N_1632,N_1294,N_1128);
or U1633 (N_1633,N_1126,N_1485);
or U1634 (N_1634,N_1419,N_1153);
nor U1635 (N_1635,N_1346,N_1375);
xor U1636 (N_1636,N_1050,N_1046);
nor U1637 (N_1637,N_1366,N_1394);
nand U1638 (N_1638,N_1292,N_1316);
or U1639 (N_1639,N_1457,N_1062);
nor U1640 (N_1640,N_1377,N_1317);
nor U1641 (N_1641,N_1338,N_1180);
or U1642 (N_1642,N_1372,N_1044);
nor U1643 (N_1643,N_1468,N_1426);
or U1644 (N_1644,N_1251,N_1291);
xor U1645 (N_1645,N_1297,N_1148);
xnor U1646 (N_1646,N_1042,N_1008);
and U1647 (N_1647,N_1205,N_1410);
and U1648 (N_1648,N_1201,N_1313);
nor U1649 (N_1649,N_1245,N_1083);
nand U1650 (N_1650,N_1430,N_1233);
nand U1651 (N_1651,N_1388,N_1092);
nand U1652 (N_1652,N_1450,N_1194);
and U1653 (N_1653,N_1289,N_1497);
or U1654 (N_1654,N_1023,N_1067);
and U1655 (N_1655,N_1137,N_1439);
nand U1656 (N_1656,N_1421,N_1445);
xnor U1657 (N_1657,N_1487,N_1309);
and U1658 (N_1658,N_1182,N_1432);
nor U1659 (N_1659,N_1181,N_1053);
and U1660 (N_1660,N_1330,N_1328);
or U1661 (N_1661,N_1241,N_1001);
xnor U1662 (N_1662,N_1209,N_1310);
or U1663 (N_1663,N_1003,N_1223);
nand U1664 (N_1664,N_1225,N_1091);
nor U1665 (N_1665,N_1006,N_1453);
nor U1666 (N_1666,N_1429,N_1011);
and U1667 (N_1667,N_1021,N_1447);
and U1668 (N_1668,N_1442,N_1165);
nand U1669 (N_1669,N_1364,N_1311);
nor U1670 (N_1670,N_1443,N_1041);
or U1671 (N_1671,N_1327,N_1160);
and U1672 (N_1672,N_1390,N_1060);
or U1673 (N_1673,N_1329,N_1454);
and U1674 (N_1674,N_1035,N_1077);
nor U1675 (N_1675,N_1406,N_1016);
and U1676 (N_1676,N_1111,N_1007);
and U1677 (N_1677,N_1493,N_1155);
or U1678 (N_1678,N_1392,N_1217);
nand U1679 (N_1679,N_1192,N_1088);
nand U1680 (N_1680,N_1399,N_1081);
nor U1681 (N_1681,N_1206,N_1221);
or U1682 (N_1682,N_1286,N_1275);
nor U1683 (N_1683,N_1422,N_1393);
nor U1684 (N_1684,N_1189,N_1113);
and U1685 (N_1685,N_1428,N_1498);
and U1686 (N_1686,N_1486,N_1010);
or U1687 (N_1687,N_1268,N_1078);
and U1688 (N_1688,N_1051,N_1056);
nor U1689 (N_1689,N_1464,N_1299);
nand U1690 (N_1690,N_1249,N_1257);
and U1691 (N_1691,N_1127,N_1451);
nand U1692 (N_1692,N_1452,N_1170);
nand U1693 (N_1693,N_1385,N_1341);
or U1694 (N_1694,N_1101,N_1152);
and U1695 (N_1695,N_1191,N_1220);
nor U1696 (N_1696,N_1004,N_1135);
and U1697 (N_1697,N_1473,N_1285);
and U1698 (N_1698,N_1140,N_1230);
and U1699 (N_1699,N_1175,N_1440);
nand U1700 (N_1700,N_1412,N_1103);
nand U1701 (N_1701,N_1204,N_1228);
xnor U1702 (N_1702,N_1133,N_1097);
nand U1703 (N_1703,N_1342,N_1258);
or U1704 (N_1704,N_1224,N_1300);
nor U1705 (N_1705,N_1147,N_1071);
or U1706 (N_1706,N_1380,N_1458);
nor U1707 (N_1707,N_1156,N_1057);
nand U1708 (N_1708,N_1059,N_1332);
nor U1709 (N_1709,N_1000,N_1020);
nor U1710 (N_1710,N_1492,N_1210);
nand U1711 (N_1711,N_1114,N_1161);
and U1712 (N_1712,N_1384,N_1484);
nor U1713 (N_1713,N_1420,N_1305);
nand U1714 (N_1714,N_1172,N_1264);
nand U1715 (N_1715,N_1323,N_1252);
xnor U1716 (N_1716,N_1260,N_1197);
nand U1717 (N_1717,N_1359,N_1383);
or U1718 (N_1718,N_1387,N_1471);
and U1719 (N_1719,N_1025,N_1284);
or U1720 (N_1720,N_1250,N_1351);
nor U1721 (N_1721,N_1395,N_1320);
nor U1722 (N_1722,N_1132,N_1255);
or U1723 (N_1723,N_1435,N_1177);
nand U1724 (N_1724,N_1105,N_1273);
nand U1725 (N_1725,N_1331,N_1407);
nand U1726 (N_1726,N_1353,N_1318);
nor U1727 (N_1727,N_1274,N_1178);
nand U1728 (N_1728,N_1438,N_1306);
or U1729 (N_1729,N_1476,N_1474);
and U1730 (N_1730,N_1068,N_1226);
or U1731 (N_1731,N_1298,N_1234);
nor U1732 (N_1732,N_1337,N_1214);
xnor U1733 (N_1733,N_1093,N_1307);
and U1734 (N_1734,N_1462,N_1460);
xor U1735 (N_1735,N_1246,N_1043);
nand U1736 (N_1736,N_1267,N_1190);
or U1737 (N_1737,N_1158,N_1427);
and U1738 (N_1738,N_1244,N_1324);
and U1739 (N_1739,N_1243,N_1169);
nand U1740 (N_1740,N_1287,N_1213);
nand U1741 (N_1741,N_1002,N_1164);
nand U1742 (N_1742,N_1441,N_1235);
nand U1743 (N_1743,N_1185,N_1483);
or U1744 (N_1744,N_1122,N_1199);
and U1745 (N_1745,N_1277,N_1112);
and U1746 (N_1746,N_1026,N_1102);
nor U1747 (N_1747,N_1098,N_1495);
nor U1748 (N_1748,N_1276,N_1186);
and U1749 (N_1749,N_1470,N_1404);
nand U1750 (N_1750,N_1110,N_1274);
nand U1751 (N_1751,N_1193,N_1041);
and U1752 (N_1752,N_1169,N_1361);
and U1753 (N_1753,N_1268,N_1269);
or U1754 (N_1754,N_1408,N_1493);
xnor U1755 (N_1755,N_1200,N_1090);
nand U1756 (N_1756,N_1278,N_1368);
or U1757 (N_1757,N_1166,N_1245);
nor U1758 (N_1758,N_1445,N_1338);
nand U1759 (N_1759,N_1215,N_1253);
and U1760 (N_1760,N_1314,N_1471);
nor U1761 (N_1761,N_1365,N_1370);
xor U1762 (N_1762,N_1078,N_1087);
xnor U1763 (N_1763,N_1163,N_1304);
or U1764 (N_1764,N_1003,N_1443);
nand U1765 (N_1765,N_1273,N_1372);
or U1766 (N_1766,N_1003,N_1099);
nand U1767 (N_1767,N_1072,N_1151);
xor U1768 (N_1768,N_1213,N_1123);
or U1769 (N_1769,N_1467,N_1021);
and U1770 (N_1770,N_1497,N_1489);
or U1771 (N_1771,N_1371,N_1271);
and U1772 (N_1772,N_1002,N_1245);
nor U1773 (N_1773,N_1378,N_1046);
or U1774 (N_1774,N_1225,N_1393);
and U1775 (N_1775,N_1144,N_1284);
nand U1776 (N_1776,N_1161,N_1277);
xnor U1777 (N_1777,N_1009,N_1171);
and U1778 (N_1778,N_1333,N_1035);
and U1779 (N_1779,N_1039,N_1403);
nand U1780 (N_1780,N_1472,N_1293);
or U1781 (N_1781,N_1414,N_1495);
nor U1782 (N_1782,N_1354,N_1001);
nor U1783 (N_1783,N_1316,N_1222);
and U1784 (N_1784,N_1295,N_1106);
xnor U1785 (N_1785,N_1266,N_1489);
nor U1786 (N_1786,N_1123,N_1234);
or U1787 (N_1787,N_1424,N_1489);
nor U1788 (N_1788,N_1179,N_1203);
nor U1789 (N_1789,N_1374,N_1060);
nor U1790 (N_1790,N_1267,N_1248);
or U1791 (N_1791,N_1113,N_1194);
and U1792 (N_1792,N_1220,N_1015);
or U1793 (N_1793,N_1090,N_1483);
and U1794 (N_1794,N_1391,N_1358);
nor U1795 (N_1795,N_1205,N_1326);
or U1796 (N_1796,N_1132,N_1096);
nand U1797 (N_1797,N_1243,N_1183);
or U1798 (N_1798,N_1454,N_1146);
nand U1799 (N_1799,N_1481,N_1439);
or U1800 (N_1800,N_1409,N_1086);
nand U1801 (N_1801,N_1268,N_1175);
or U1802 (N_1802,N_1401,N_1306);
and U1803 (N_1803,N_1344,N_1417);
or U1804 (N_1804,N_1335,N_1305);
nor U1805 (N_1805,N_1043,N_1008);
nor U1806 (N_1806,N_1447,N_1277);
or U1807 (N_1807,N_1446,N_1238);
or U1808 (N_1808,N_1195,N_1298);
nor U1809 (N_1809,N_1311,N_1160);
xor U1810 (N_1810,N_1232,N_1126);
nand U1811 (N_1811,N_1151,N_1425);
nand U1812 (N_1812,N_1361,N_1265);
and U1813 (N_1813,N_1335,N_1199);
xor U1814 (N_1814,N_1249,N_1425);
nor U1815 (N_1815,N_1087,N_1307);
nand U1816 (N_1816,N_1222,N_1124);
nor U1817 (N_1817,N_1369,N_1021);
or U1818 (N_1818,N_1436,N_1131);
and U1819 (N_1819,N_1260,N_1160);
nand U1820 (N_1820,N_1085,N_1135);
and U1821 (N_1821,N_1465,N_1423);
nand U1822 (N_1822,N_1182,N_1154);
nor U1823 (N_1823,N_1374,N_1429);
or U1824 (N_1824,N_1133,N_1437);
nand U1825 (N_1825,N_1294,N_1038);
nand U1826 (N_1826,N_1439,N_1126);
nand U1827 (N_1827,N_1499,N_1070);
and U1828 (N_1828,N_1450,N_1178);
nand U1829 (N_1829,N_1013,N_1299);
nor U1830 (N_1830,N_1208,N_1055);
nand U1831 (N_1831,N_1154,N_1489);
or U1832 (N_1832,N_1398,N_1419);
xor U1833 (N_1833,N_1276,N_1374);
nand U1834 (N_1834,N_1337,N_1265);
xor U1835 (N_1835,N_1446,N_1010);
nand U1836 (N_1836,N_1186,N_1385);
or U1837 (N_1837,N_1047,N_1268);
xor U1838 (N_1838,N_1320,N_1333);
nand U1839 (N_1839,N_1108,N_1193);
nand U1840 (N_1840,N_1179,N_1219);
nor U1841 (N_1841,N_1140,N_1294);
and U1842 (N_1842,N_1125,N_1310);
and U1843 (N_1843,N_1080,N_1458);
nand U1844 (N_1844,N_1213,N_1413);
and U1845 (N_1845,N_1408,N_1465);
nand U1846 (N_1846,N_1398,N_1148);
or U1847 (N_1847,N_1155,N_1189);
nor U1848 (N_1848,N_1183,N_1439);
and U1849 (N_1849,N_1145,N_1297);
or U1850 (N_1850,N_1422,N_1147);
or U1851 (N_1851,N_1233,N_1428);
nand U1852 (N_1852,N_1133,N_1228);
and U1853 (N_1853,N_1196,N_1215);
or U1854 (N_1854,N_1346,N_1105);
nand U1855 (N_1855,N_1043,N_1101);
and U1856 (N_1856,N_1067,N_1159);
or U1857 (N_1857,N_1218,N_1457);
or U1858 (N_1858,N_1461,N_1247);
or U1859 (N_1859,N_1082,N_1248);
nor U1860 (N_1860,N_1191,N_1493);
nor U1861 (N_1861,N_1025,N_1129);
and U1862 (N_1862,N_1091,N_1414);
xnor U1863 (N_1863,N_1323,N_1301);
and U1864 (N_1864,N_1052,N_1259);
xor U1865 (N_1865,N_1484,N_1368);
nand U1866 (N_1866,N_1017,N_1472);
nand U1867 (N_1867,N_1150,N_1009);
nand U1868 (N_1868,N_1188,N_1331);
and U1869 (N_1869,N_1017,N_1205);
xor U1870 (N_1870,N_1223,N_1080);
nand U1871 (N_1871,N_1056,N_1044);
nor U1872 (N_1872,N_1413,N_1294);
nand U1873 (N_1873,N_1367,N_1171);
nor U1874 (N_1874,N_1409,N_1449);
nand U1875 (N_1875,N_1319,N_1160);
and U1876 (N_1876,N_1161,N_1126);
nor U1877 (N_1877,N_1381,N_1063);
nand U1878 (N_1878,N_1067,N_1011);
and U1879 (N_1879,N_1486,N_1134);
or U1880 (N_1880,N_1397,N_1228);
nand U1881 (N_1881,N_1363,N_1243);
or U1882 (N_1882,N_1429,N_1114);
nand U1883 (N_1883,N_1209,N_1229);
nand U1884 (N_1884,N_1101,N_1212);
xnor U1885 (N_1885,N_1077,N_1482);
or U1886 (N_1886,N_1270,N_1109);
nor U1887 (N_1887,N_1187,N_1412);
nand U1888 (N_1888,N_1355,N_1010);
or U1889 (N_1889,N_1445,N_1187);
nand U1890 (N_1890,N_1308,N_1441);
nor U1891 (N_1891,N_1495,N_1072);
xnor U1892 (N_1892,N_1335,N_1459);
or U1893 (N_1893,N_1149,N_1461);
nor U1894 (N_1894,N_1457,N_1095);
nand U1895 (N_1895,N_1260,N_1158);
nor U1896 (N_1896,N_1248,N_1395);
nor U1897 (N_1897,N_1113,N_1469);
or U1898 (N_1898,N_1216,N_1418);
or U1899 (N_1899,N_1238,N_1415);
nor U1900 (N_1900,N_1072,N_1158);
nor U1901 (N_1901,N_1405,N_1089);
or U1902 (N_1902,N_1084,N_1237);
or U1903 (N_1903,N_1231,N_1458);
or U1904 (N_1904,N_1360,N_1470);
nor U1905 (N_1905,N_1497,N_1017);
nand U1906 (N_1906,N_1076,N_1468);
nor U1907 (N_1907,N_1429,N_1006);
nand U1908 (N_1908,N_1154,N_1062);
nor U1909 (N_1909,N_1005,N_1282);
and U1910 (N_1910,N_1100,N_1051);
nand U1911 (N_1911,N_1136,N_1350);
or U1912 (N_1912,N_1384,N_1143);
nor U1913 (N_1913,N_1359,N_1095);
nand U1914 (N_1914,N_1026,N_1270);
and U1915 (N_1915,N_1002,N_1103);
and U1916 (N_1916,N_1360,N_1358);
nand U1917 (N_1917,N_1392,N_1483);
nor U1918 (N_1918,N_1038,N_1493);
nor U1919 (N_1919,N_1451,N_1485);
or U1920 (N_1920,N_1323,N_1415);
nor U1921 (N_1921,N_1096,N_1369);
xnor U1922 (N_1922,N_1062,N_1481);
nor U1923 (N_1923,N_1106,N_1301);
nor U1924 (N_1924,N_1036,N_1264);
and U1925 (N_1925,N_1315,N_1209);
or U1926 (N_1926,N_1400,N_1413);
nand U1927 (N_1927,N_1395,N_1490);
or U1928 (N_1928,N_1433,N_1225);
xor U1929 (N_1929,N_1404,N_1043);
nand U1930 (N_1930,N_1006,N_1065);
nand U1931 (N_1931,N_1413,N_1307);
nor U1932 (N_1932,N_1358,N_1218);
and U1933 (N_1933,N_1220,N_1492);
or U1934 (N_1934,N_1488,N_1092);
and U1935 (N_1935,N_1378,N_1398);
and U1936 (N_1936,N_1029,N_1292);
or U1937 (N_1937,N_1073,N_1115);
nand U1938 (N_1938,N_1469,N_1203);
nand U1939 (N_1939,N_1383,N_1316);
nor U1940 (N_1940,N_1349,N_1150);
or U1941 (N_1941,N_1066,N_1470);
nor U1942 (N_1942,N_1281,N_1228);
xnor U1943 (N_1943,N_1355,N_1324);
xnor U1944 (N_1944,N_1077,N_1259);
and U1945 (N_1945,N_1001,N_1191);
and U1946 (N_1946,N_1088,N_1263);
nand U1947 (N_1947,N_1119,N_1257);
nand U1948 (N_1948,N_1181,N_1397);
nand U1949 (N_1949,N_1014,N_1358);
nor U1950 (N_1950,N_1030,N_1361);
nor U1951 (N_1951,N_1301,N_1177);
nor U1952 (N_1952,N_1108,N_1166);
nor U1953 (N_1953,N_1440,N_1125);
or U1954 (N_1954,N_1311,N_1454);
and U1955 (N_1955,N_1167,N_1373);
nor U1956 (N_1956,N_1020,N_1195);
nor U1957 (N_1957,N_1430,N_1177);
xnor U1958 (N_1958,N_1335,N_1230);
or U1959 (N_1959,N_1407,N_1462);
or U1960 (N_1960,N_1454,N_1465);
nor U1961 (N_1961,N_1131,N_1245);
nor U1962 (N_1962,N_1330,N_1095);
xnor U1963 (N_1963,N_1449,N_1311);
nand U1964 (N_1964,N_1408,N_1101);
nor U1965 (N_1965,N_1301,N_1179);
or U1966 (N_1966,N_1141,N_1419);
or U1967 (N_1967,N_1361,N_1353);
nor U1968 (N_1968,N_1109,N_1311);
and U1969 (N_1969,N_1172,N_1377);
or U1970 (N_1970,N_1389,N_1232);
nor U1971 (N_1971,N_1156,N_1472);
or U1972 (N_1972,N_1435,N_1483);
or U1973 (N_1973,N_1286,N_1044);
or U1974 (N_1974,N_1365,N_1352);
and U1975 (N_1975,N_1241,N_1219);
and U1976 (N_1976,N_1088,N_1152);
nand U1977 (N_1977,N_1377,N_1487);
and U1978 (N_1978,N_1487,N_1466);
or U1979 (N_1979,N_1483,N_1258);
or U1980 (N_1980,N_1258,N_1241);
or U1981 (N_1981,N_1263,N_1481);
xnor U1982 (N_1982,N_1178,N_1427);
or U1983 (N_1983,N_1013,N_1288);
nor U1984 (N_1984,N_1404,N_1172);
nor U1985 (N_1985,N_1012,N_1344);
nand U1986 (N_1986,N_1153,N_1379);
or U1987 (N_1987,N_1040,N_1395);
or U1988 (N_1988,N_1187,N_1437);
or U1989 (N_1989,N_1216,N_1241);
and U1990 (N_1990,N_1370,N_1247);
nand U1991 (N_1991,N_1172,N_1118);
nand U1992 (N_1992,N_1405,N_1117);
nor U1993 (N_1993,N_1322,N_1038);
and U1994 (N_1994,N_1104,N_1491);
nand U1995 (N_1995,N_1314,N_1132);
nor U1996 (N_1996,N_1280,N_1234);
xnor U1997 (N_1997,N_1037,N_1236);
nor U1998 (N_1998,N_1407,N_1119);
nor U1999 (N_1999,N_1434,N_1253);
or U2000 (N_2000,N_1602,N_1508);
and U2001 (N_2001,N_1789,N_1858);
nand U2002 (N_2002,N_1964,N_1919);
and U2003 (N_2003,N_1968,N_1900);
or U2004 (N_2004,N_1957,N_1679);
nand U2005 (N_2005,N_1888,N_1887);
and U2006 (N_2006,N_1871,N_1688);
nand U2007 (N_2007,N_1661,N_1956);
and U2008 (N_2008,N_1958,N_1922);
and U2009 (N_2009,N_1593,N_1934);
nor U2010 (N_2010,N_1659,N_1836);
nor U2011 (N_2011,N_1945,N_1827);
and U2012 (N_2012,N_1708,N_1924);
and U2013 (N_2013,N_1723,N_1705);
or U2014 (N_2014,N_1638,N_1833);
or U2015 (N_2015,N_1687,N_1624);
xor U2016 (N_2016,N_1883,N_1840);
nand U2017 (N_2017,N_1648,N_1930);
or U2018 (N_2018,N_1910,N_1588);
and U2019 (N_2019,N_1763,N_1890);
and U2020 (N_2020,N_1989,N_1579);
or U2021 (N_2021,N_1605,N_1757);
and U2022 (N_2022,N_1783,N_1851);
or U2023 (N_2023,N_1891,N_1750);
nor U2024 (N_2024,N_1854,N_1967);
and U2025 (N_2025,N_1960,N_1549);
nand U2026 (N_2026,N_1632,N_1722);
or U2027 (N_2027,N_1849,N_1741);
or U2028 (N_2028,N_1601,N_1935);
or U2029 (N_2029,N_1907,N_1905);
nor U2030 (N_2030,N_1850,N_1716);
and U2031 (N_2031,N_1999,N_1842);
or U2032 (N_2032,N_1585,N_1525);
and U2033 (N_2033,N_1509,N_1726);
and U2034 (N_2034,N_1787,N_1813);
and U2035 (N_2035,N_1595,N_1812);
nor U2036 (N_2036,N_1558,N_1564);
and U2037 (N_2037,N_1954,N_1870);
and U2038 (N_2038,N_1927,N_1516);
xor U2039 (N_2039,N_1942,N_1537);
nand U2040 (N_2040,N_1686,N_1590);
nor U2041 (N_2041,N_1879,N_1559);
and U2042 (N_2042,N_1589,N_1550);
nand U2043 (N_2043,N_1546,N_1796);
nor U2044 (N_2044,N_1758,N_1583);
or U2045 (N_2045,N_1665,N_1754);
or U2046 (N_2046,N_1540,N_1520);
nor U2047 (N_2047,N_1738,N_1551);
and U2048 (N_2048,N_1785,N_1568);
and U2049 (N_2049,N_1501,N_1683);
nand U2050 (N_2050,N_1697,N_1777);
xor U2051 (N_2051,N_1894,N_1734);
nand U2052 (N_2052,N_1664,N_1896);
or U2053 (N_2053,N_1507,N_1528);
xor U2054 (N_2054,N_1510,N_1543);
nand U2055 (N_2055,N_1644,N_1994);
and U2056 (N_2056,N_1557,N_1881);
xor U2057 (N_2057,N_1929,N_1662);
or U2058 (N_2058,N_1569,N_1859);
nand U2059 (N_2059,N_1502,N_1959);
and U2060 (N_2060,N_1869,N_1656);
or U2061 (N_2061,N_1966,N_1639);
nor U2062 (N_2062,N_1682,N_1594);
nor U2063 (N_2063,N_1591,N_1715);
or U2064 (N_2064,N_1992,N_1725);
nor U2065 (N_2065,N_1824,N_1802);
and U2066 (N_2066,N_1643,N_1645);
or U2067 (N_2067,N_1611,N_1831);
and U2068 (N_2068,N_1848,N_1646);
or U2069 (N_2069,N_1839,N_1993);
nor U2070 (N_2070,N_1852,N_1673);
or U2071 (N_2071,N_1599,N_1577);
and U2072 (N_2072,N_1744,N_1616);
or U2073 (N_2073,N_1529,N_1668);
nor U2074 (N_2074,N_1675,N_1765);
nor U2075 (N_2075,N_1556,N_1823);
nand U2076 (N_2076,N_1768,N_1774);
and U2077 (N_2077,N_1914,N_1707);
and U2078 (N_2078,N_1838,N_1511);
or U2079 (N_2079,N_1915,N_1971);
nor U2080 (N_2080,N_1953,N_1933);
and U2081 (N_2081,N_1925,N_1533);
or U2082 (N_2082,N_1737,N_1753);
nand U2083 (N_2083,N_1685,N_1514);
or U2084 (N_2084,N_1955,N_1906);
or U2085 (N_2085,N_1633,N_1926);
nor U2086 (N_2086,N_1710,N_1610);
and U2087 (N_2087,N_1988,N_1658);
and U2088 (N_2088,N_1819,N_1619);
or U2089 (N_2089,N_1554,N_1666);
nor U2090 (N_2090,N_1652,N_1820);
nand U2091 (N_2091,N_1776,N_1635);
and U2092 (N_2092,N_1853,N_1884);
and U2093 (N_2093,N_1649,N_1563);
nand U2094 (N_2094,N_1573,N_1739);
or U2095 (N_2095,N_1604,N_1628);
nor U2096 (N_2096,N_1713,N_1779);
and U2097 (N_2097,N_1825,N_1822);
nand U2098 (N_2098,N_1855,N_1637);
nand U2099 (N_2099,N_1598,N_1752);
or U2100 (N_2100,N_1747,N_1578);
nor U2101 (N_2101,N_1703,N_1863);
nor U2102 (N_2102,N_1614,N_1818);
nor U2103 (N_2103,N_1788,N_1641);
nor U2104 (N_2104,N_1948,N_1584);
nor U2105 (N_2105,N_1817,N_1834);
xnor U2106 (N_2106,N_1609,N_1830);
nand U2107 (N_2107,N_1745,N_1718);
or U2108 (N_2108,N_1545,N_1524);
nor U2109 (N_2109,N_1672,N_1983);
and U2110 (N_2110,N_1943,N_1553);
or U2111 (N_2111,N_1721,N_1762);
nor U2112 (N_2112,N_1913,N_1560);
and U2113 (N_2113,N_1576,N_1872);
nor U2114 (N_2114,N_1607,N_1691);
or U2115 (N_2115,N_1519,N_1760);
xor U2116 (N_2116,N_1908,N_1606);
nor U2117 (N_2117,N_1808,N_1677);
nand U2118 (N_2118,N_1909,N_1775);
and U2119 (N_2119,N_1944,N_1868);
and U2120 (N_2120,N_1847,N_1902);
nand U2121 (N_2121,N_1972,N_1596);
nand U2122 (N_2122,N_1640,N_1692);
or U2123 (N_2123,N_1978,N_1899);
nor U2124 (N_2124,N_1660,N_1617);
nand U2125 (N_2125,N_1742,N_1521);
nand U2126 (N_2126,N_1998,N_1527);
nand U2127 (N_2127,N_1866,N_1636);
and U2128 (N_2128,N_1903,N_1620);
and U2129 (N_2129,N_1570,N_1571);
or U2130 (N_2130,N_1809,N_1980);
nor U2131 (N_2131,N_1976,N_1729);
xnor U2132 (N_2132,N_1965,N_1506);
or U2133 (N_2133,N_1987,N_1795);
nor U2134 (N_2134,N_1642,N_1699);
nand U2135 (N_2135,N_1766,N_1719);
or U2136 (N_2136,N_1650,N_1975);
or U2137 (N_2137,N_1990,N_1751);
or U2138 (N_2138,N_1886,N_1949);
nor U2139 (N_2139,N_1518,N_1829);
and U2140 (N_2140,N_1936,N_1709);
nand U2141 (N_2141,N_1689,N_1904);
and U2142 (N_2142,N_1653,N_1567);
nand U2143 (N_2143,N_1912,N_1864);
nand U2144 (N_2144,N_1951,N_1669);
xor U2145 (N_2145,N_1878,N_1512);
nor U2146 (N_2146,N_1676,N_1698);
and U2147 (N_2147,N_1627,N_1773);
or U2148 (N_2148,N_1678,N_1655);
or U2149 (N_2149,N_1844,N_1803);
nand U2150 (N_2150,N_1748,N_1963);
nand U2151 (N_2151,N_1608,N_1982);
or U2152 (N_2152,N_1928,N_1671);
nor U2153 (N_2153,N_1874,N_1523);
or U2154 (N_2154,N_1732,N_1625);
nand U2155 (N_2155,N_1937,N_1892);
and U2156 (N_2156,N_1592,N_1946);
or U2157 (N_2157,N_1740,N_1674);
or U2158 (N_2158,N_1701,N_1897);
or U2159 (N_2159,N_1974,N_1950);
nand U2160 (N_2160,N_1746,N_1889);
nand U2161 (N_2161,N_1513,N_1805);
nor U2162 (N_2162,N_1535,N_1735);
nor U2163 (N_2163,N_1837,N_1806);
nand U2164 (N_2164,N_1505,N_1544);
and U2165 (N_2165,N_1811,N_1939);
nor U2166 (N_2166,N_1728,N_1986);
nand U2167 (N_2167,N_1970,N_1804);
or U2168 (N_2168,N_1696,N_1843);
nand U2169 (N_2169,N_1684,N_1981);
nand U2170 (N_2170,N_1730,N_1828);
and U2171 (N_2171,N_1700,N_1756);
and U2172 (N_2172,N_1603,N_1565);
nand U2173 (N_2173,N_1657,N_1706);
nand U2174 (N_2174,N_1630,N_1997);
and U2175 (N_2175,N_1938,N_1799);
nand U2176 (N_2176,N_1694,N_1736);
nand U2177 (N_2177,N_1821,N_1500);
nand U2178 (N_2178,N_1724,N_1597);
nor U2179 (N_2179,N_1634,N_1873);
nor U2180 (N_2180,N_1712,N_1784);
and U2181 (N_2181,N_1704,N_1932);
or U2182 (N_2182,N_1711,N_1552);
or U2183 (N_2183,N_1893,N_1876);
nor U2184 (N_2184,N_1875,N_1612);
or U2185 (N_2185,N_1917,N_1586);
and U2186 (N_2186,N_1901,N_1670);
nand U2187 (N_2187,N_1767,N_1654);
nand U2188 (N_2188,N_1931,N_1856);
and U2189 (N_2189,N_1566,N_1526);
xnor U2190 (N_2190,N_1798,N_1845);
and U2191 (N_2191,N_1581,N_1538);
nand U2192 (N_2192,N_1952,N_1769);
or U2193 (N_2193,N_1727,N_1522);
nand U2194 (N_2194,N_1921,N_1898);
xnor U2195 (N_2195,N_1790,N_1786);
nand U2196 (N_2196,N_1920,N_1962);
nand U2197 (N_2197,N_1717,N_1996);
or U2198 (N_2198,N_1814,N_1749);
xnor U2199 (N_2199,N_1810,N_1923);
nor U2200 (N_2200,N_1984,N_1861);
or U2201 (N_2201,N_1780,N_1714);
and U2202 (N_2202,N_1582,N_1503);
nand U2203 (N_2203,N_1695,N_1680);
nand U2204 (N_2204,N_1792,N_1663);
or U2205 (N_2205,N_1860,N_1977);
nor U2206 (N_2206,N_1807,N_1969);
or U2207 (N_2207,N_1548,N_1743);
and U2208 (N_2208,N_1877,N_1794);
xnor U2209 (N_2209,N_1562,N_1622);
or U2210 (N_2210,N_1764,N_1561);
nor U2211 (N_2211,N_1755,N_1613);
xor U2212 (N_2212,N_1895,N_1555);
and U2213 (N_2213,N_1991,N_1761);
or U2214 (N_2214,N_1882,N_1885);
nand U2215 (N_2215,N_1846,N_1542);
or U2216 (N_2216,N_1916,N_1572);
and U2217 (N_2217,N_1575,N_1880);
or U2218 (N_2218,N_1541,N_1574);
nand U2219 (N_2219,N_1759,N_1800);
nand U2220 (N_2220,N_1731,N_1770);
or U2221 (N_2221,N_1615,N_1778);
nor U2222 (N_2222,N_1539,N_1947);
and U2223 (N_2223,N_1797,N_1720);
nand U2224 (N_2224,N_1702,N_1651);
or U2225 (N_2225,N_1826,N_1531);
nor U2226 (N_2226,N_1681,N_1623);
nand U2227 (N_2227,N_1536,N_1793);
or U2228 (N_2228,N_1772,N_1782);
and U2229 (N_2229,N_1580,N_1530);
or U2230 (N_2230,N_1600,N_1862);
nor U2231 (N_2231,N_1816,N_1865);
nand U2232 (N_2232,N_1781,N_1835);
and U2233 (N_2233,N_1626,N_1504);
nand U2234 (N_2234,N_1647,N_1547);
or U2235 (N_2235,N_1621,N_1918);
nor U2236 (N_2236,N_1867,N_1841);
xnor U2237 (N_2237,N_1979,N_1941);
or U2238 (N_2238,N_1629,N_1515);
or U2239 (N_2239,N_1995,N_1973);
nand U2240 (N_2240,N_1517,N_1690);
nand U2241 (N_2241,N_1940,N_1832);
nor U2242 (N_2242,N_1667,N_1791);
nor U2243 (N_2243,N_1911,N_1631);
or U2244 (N_2244,N_1733,N_1771);
nor U2245 (N_2245,N_1985,N_1961);
and U2246 (N_2246,N_1532,N_1587);
or U2247 (N_2247,N_1618,N_1534);
nor U2248 (N_2248,N_1693,N_1857);
or U2249 (N_2249,N_1815,N_1801);
and U2250 (N_2250,N_1878,N_1664);
xnor U2251 (N_2251,N_1510,N_1503);
nor U2252 (N_2252,N_1827,N_1799);
nand U2253 (N_2253,N_1649,N_1776);
and U2254 (N_2254,N_1873,N_1705);
or U2255 (N_2255,N_1897,N_1950);
nand U2256 (N_2256,N_1986,N_1602);
or U2257 (N_2257,N_1999,N_1958);
xnor U2258 (N_2258,N_1593,N_1532);
or U2259 (N_2259,N_1507,N_1692);
or U2260 (N_2260,N_1896,N_1532);
nor U2261 (N_2261,N_1507,N_1909);
nor U2262 (N_2262,N_1735,N_1667);
nor U2263 (N_2263,N_1999,N_1818);
nor U2264 (N_2264,N_1669,N_1760);
xor U2265 (N_2265,N_1741,N_1507);
and U2266 (N_2266,N_1714,N_1637);
nand U2267 (N_2267,N_1764,N_1588);
and U2268 (N_2268,N_1768,N_1751);
xor U2269 (N_2269,N_1522,N_1926);
or U2270 (N_2270,N_1672,N_1806);
and U2271 (N_2271,N_1764,N_1720);
nand U2272 (N_2272,N_1536,N_1551);
nor U2273 (N_2273,N_1760,N_1928);
nand U2274 (N_2274,N_1836,N_1567);
or U2275 (N_2275,N_1516,N_1814);
nand U2276 (N_2276,N_1623,N_1625);
nor U2277 (N_2277,N_1557,N_1622);
or U2278 (N_2278,N_1531,N_1692);
and U2279 (N_2279,N_1811,N_1848);
or U2280 (N_2280,N_1941,N_1592);
or U2281 (N_2281,N_1841,N_1686);
and U2282 (N_2282,N_1668,N_1727);
nor U2283 (N_2283,N_1871,N_1888);
nor U2284 (N_2284,N_1810,N_1500);
and U2285 (N_2285,N_1626,N_1664);
or U2286 (N_2286,N_1805,N_1585);
nand U2287 (N_2287,N_1851,N_1714);
nand U2288 (N_2288,N_1625,N_1519);
and U2289 (N_2289,N_1885,N_1820);
or U2290 (N_2290,N_1944,N_1817);
or U2291 (N_2291,N_1544,N_1989);
nand U2292 (N_2292,N_1981,N_1783);
and U2293 (N_2293,N_1897,N_1903);
nor U2294 (N_2294,N_1766,N_1938);
and U2295 (N_2295,N_1801,N_1602);
or U2296 (N_2296,N_1581,N_1893);
and U2297 (N_2297,N_1927,N_1634);
and U2298 (N_2298,N_1985,N_1561);
or U2299 (N_2299,N_1541,N_1778);
or U2300 (N_2300,N_1774,N_1650);
xnor U2301 (N_2301,N_1668,N_1737);
or U2302 (N_2302,N_1578,N_1753);
nand U2303 (N_2303,N_1637,N_1630);
nand U2304 (N_2304,N_1885,N_1863);
or U2305 (N_2305,N_1564,N_1689);
nand U2306 (N_2306,N_1903,N_1695);
nand U2307 (N_2307,N_1934,N_1884);
nand U2308 (N_2308,N_1984,N_1917);
nor U2309 (N_2309,N_1768,N_1857);
and U2310 (N_2310,N_1589,N_1531);
nand U2311 (N_2311,N_1784,N_1732);
xor U2312 (N_2312,N_1779,N_1932);
or U2313 (N_2313,N_1792,N_1807);
nand U2314 (N_2314,N_1958,N_1786);
nor U2315 (N_2315,N_1645,N_1767);
or U2316 (N_2316,N_1756,N_1752);
nor U2317 (N_2317,N_1963,N_1823);
and U2318 (N_2318,N_1773,N_1555);
nor U2319 (N_2319,N_1847,N_1844);
xnor U2320 (N_2320,N_1604,N_1691);
or U2321 (N_2321,N_1862,N_1863);
or U2322 (N_2322,N_1533,N_1966);
nor U2323 (N_2323,N_1682,N_1759);
nand U2324 (N_2324,N_1905,N_1545);
nor U2325 (N_2325,N_1770,N_1521);
or U2326 (N_2326,N_1648,N_1543);
or U2327 (N_2327,N_1652,N_1918);
or U2328 (N_2328,N_1682,N_1677);
nand U2329 (N_2329,N_1807,N_1531);
and U2330 (N_2330,N_1535,N_1744);
or U2331 (N_2331,N_1673,N_1904);
xnor U2332 (N_2332,N_1908,N_1797);
or U2333 (N_2333,N_1798,N_1994);
and U2334 (N_2334,N_1888,N_1566);
nor U2335 (N_2335,N_1650,N_1848);
xor U2336 (N_2336,N_1586,N_1703);
nand U2337 (N_2337,N_1834,N_1995);
and U2338 (N_2338,N_1727,N_1928);
or U2339 (N_2339,N_1555,N_1614);
nor U2340 (N_2340,N_1816,N_1747);
and U2341 (N_2341,N_1559,N_1957);
nand U2342 (N_2342,N_1671,N_1870);
nand U2343 (N_2343,N_1753,N_1532);
and U2344 (N_2344,N_1991,N_1822);
and U2345 (N_2345,N_1665,N_1988);
nand U2346 (N_2346,N_1950,N_1642);
and U2347 (N_2347,N_1854,N_1766);
and U2348 (N_2348,N_1911,N_1558);
and U2349 (N_2349,N_1773,N_1758);
nor U2350 (N_2350,N_1760,N_1537);
nor U2351 (N_2351,N_1681,N_1970);
nand U2352 (N_2352,N_1618,N_1908);
nand U2353 (N_2353,N_1984,N_1688);
and U2354 (N_2354,N_1528,N_1601);
and U2355 (N_2355,N_1509,N_1974);
xnor U2356 (N_2356,N_1588,N_1500);
and U2357 (N_2357,N_1845,N_1987);
nand U2358 (N_2358,N_1907,N_1932);
nor U2359 (N_2359,N_1504,N_1806);
nor U2360 (N_2360,N_1871,N_1719);
nand U2361 (N_2361,N_1594,N_1832);
nor U2362 (N_2362,N_1861,N_1767);
xor U2363 (N_2363,N_1618,N_1902);
xnor U2364 (N_2364,N_1507,N_1676);
or U2365 (N_2365,N_1660,N_1752);
nor U2366 (N_2366,N_1860,N_1868);
nor U2367 (N_2367,N_1971,N_1974);
nor U2368 (N_2368,N_1597,N_1879);
nand U2369 (N_2369,N_1559,N_1587);
or U2370 (N_2370,N_1793,N_1705);
and U2371 (N_2371,N_1699,N_1525);
and U2372 (N_2372,N_1681,N_1723);
and U2373 (N_2373,N_1509,N_1990);
nor U2374 (N_2374,N_1572,N_1718);
or U2375 (N_2375,N_1512,N_1920);
and U2376 (N_2376,N_1855,N_1733);
nor U2377 (N_2377,N_1840,N_1971);
xnor U2378 (N_2378,N_1996,N_1707);
nand U2379 (N_2379,N_1696,N_1977);
nand U2380 (N_2380,N_1654,N_1814);
nor U2381 (N_2381,N_1598,N_1681);
and U2382 (N_2382,N_1765,N_1857);
nor U2383 (N_2383,N_1755,N_1950);
or U2384 (N_2384,N_1801,N_1925);
xnor U2385 (N_2385,N_1660,N_1943);
or U2386 (N_2386,N_1913,N_1515);
and U2387 (N_2387,N_1821,N_1515);
nor U2388 (N_2388,N_1762,N_1680);
or U2389 (N_2389,N_1562,N_1852);
or U2390 (N_2390,N_1651,N_1792);
xnor U2391 (N_2391,N_1526,N_1630);
nand U2392 (N_2392,N_1851,N_1904);
xor U2393 (N_2393,N_1526,N_1531);
and U2394 (N_2394,N_1552,N_1748);
xnor U2395 (N_2395,N_1704,N_1504);
nand U2396 (N_2396,N_1814,N_1817);
nor U2397 (N_2397,N_1598,N_1595);
and U2398 (N_2398,N_1644,N_1683);
or U2399 (N_2399,N_1859,N_1605);
or U2400 (N_2400,N_1672,N_1859);
nor U2401 (N_2401,N_1793,N_1595);
or U2402 (N_2402,N_1591,N_1653);
nand U2403 (N_2403,N_1853,N_1800);
nor U2404 (N_2404,N_1689,N_1817);
and U2405 (N_2405,N_1550,N_1826);
xor U2406 (N_2406,N_1513,N_1928);
nand U2407 (N_2407,N_1983,N_1894);
nand U2408 (N_2408,N_1969,N_1875);
and U2409 (N_2409,N_1959,N_1932);
nor U2410 (N_2410,N_1650,N_1768);
and U2411 (N_2411,N_1996,N_1660);
or U2412 (N_2412,N_1890,N_1526);
or U2413 (N_2413,N_1764,N_1944);
xnor U2414 (N_2414,N_1527,N_1802);
and U2415 (N_2415,N_1511,N_1571);
and U2416 (N_2416,N_1713,N_1806);
nor U2417 (N_2417,N_1759,N_1597);
xor U2418 (N_2418,N_1961,N_1892);
nor U2419 (N_2419,N_1528,N_1503);
and U2420 (N_2420,N_1571,N_1857);
nand U2421 (N_2421,N_1807,N_1732);
and U2422 (N_2422,N_1868,N_1688);
nor U2423 (N_2423,N_1636,N_1810);
or U2424 (N_2424,N_1802,N_1921);
nand U2425 (N_2425,N_1916,N_1886);
and U2426 (N_2426,N_1546,N_1569);
xnor U2427 (N_2427,N_1654,N_1882);
xor U2428 (N_2428,N_1654,N_1929);
xnor U2429 (N_2429,N_1889,N_1764);
nor U2430 (N_2430,N_1718,N_1917);
nand U2431 (N_2431,N_1706,N_1569);
nor U2432 (N_2432,N_1860,N_1614);
xor U2433 (N_2433,N_1694,N_1764);
nand U2434 (N_2434,N_1954,N_1518);
or U2435 (N_2435,N_1956,N_1517);
or U2436 (N_2436,N_1618,N_1788);
xnor U2437 (N_2437,N_1840,N_1675);
or U2438 (N_2438,N_1846,N_1693);
nand U2439 (N_2439,N_1931,N_1847);
or U2440 (N_2440,N_1572,N_1887);
nor U2441 (N_2441,N_1908,N_1822);
and U2442 (N_2442,N_1671,N_1971);
nand U2443 (N_2443,N_1520,N_1551);
nor U2444 (N_2444,N_1536,N_1994);
nor U2445 (N_2445,N_1881,N_1566);
nor U2446 (N_2446,N_1905,N_1799);
and U2447 (N_2447,N_1746,N_1796);
and U2448 (N_2448,N_1893,N_1775);
or U2449 (N_2449,N_1666,N_1713);
nor U2450 (N_2450,N_1905,N_1862);
nor U2451 (N_2451,N_1678,N_1812);
nor U2452 (N_2452,N_1682,N_1583);
nand U2453 (N_2453,N_1642,N_1864);
nand U2454 (N_2454,N_1829,N_1781);
or U2455 (N_2455,N_1722,N_1763);
xor U2456 (N_2456,N_1562,N_1992);
nand U2457 (N_2457,N_1832,N_1888);
or U2458 (N_2458,N_1814,N_1925);
nor U2459 (N_2459,N_1904,N_1508);
nand U2460 (N_2460,N_1816,N_1881);
or U2461 (N_2461,N_1953,N_1719);
and U2462 (N_2462,N_1712,N_1621);
nand U2463 (N_2463,N_1840,N_1657);
and U2464 (N_2464,N_1974,N_1586);
xnor U2465 (N_2465,N_1824,N_1847);
nor U2466 (N_2466,N_1620,N_1655);
nor U2467 (N_2467,N_1771,N_1992);
nand U2468 (N_2468,N_1993,N_1604);
nor U2469 (N_2469,N_1596,N_1837);
nand U2470 (N_2470,N_1581,N_1559);
and U2471 (N_2471,N_1730,N_1928);
nor U2472 (N_2472,N_1582,N_1903);
or U2473 (N_2473,N_1734,N_1981);
nor U2474 (N_2474,N_1637,N_1713);
or U2475 (N_2475,N_1796,N_1801);
nand U2476 (N_2476,N_1585,N_1859);
and U2477 (N_2477,N_1977,N_1890);
nand U2478 (N_2478,N_1881,N_1915);
or U2479 (N_2479,N_1836,N_1871);
nor U2480 (N_2480,N_1958,N_1784);
and U2481 (N_2481,N_1678,N_1741);
nand U2482 (N_2482,N_1725,N_1831);
and U2483 (N_2483,N_1727,N_1989);
nand U2484 (N_2484,N_1738,N_1520);
or U2485 (N_2485,N_1947,N_1736);
or U2486 (N_2486,N_1759,N_1985);
xnor U2487 (N_2487,N_1552,N_1731);
or U2488 (N_2488,N_1636,N_1998);
and U2489 (N_2489,N_1530,N_1963);
or U2490 (N_2490,N_1642,N_1577);
xnor U2491 (N_2491,N_1797,N_1669);
and U2492 (N_2492,N_1684,N_1823);
and U2493 (N_2493,N_1927,N_1796);
and U2494 (N_2494,N_1879,N_1880);
or U2495 (N_2495,N_1636,N_1534);
and U2496 (N_2496,N_1700,N_1558);
and U2497 (N_2497,N_1552,N_1907);
nor U2498 (N_2498,N_1847,N_1948);
or U2499 (N_2499,N_1588,N_1609);
or U2500 (N_2500,N_2472,N_2376);
or U2501 (N_2501,N_2145,N_2367);
or U2502 (N_2502,N_2392,N_2110);
nor U2503 (N_2503,N_2259,N_2002);
nand U2504 (N_2504,N_2418,N_2091);
nand U2505 (N_2505,N_2374,N_2056);
xor U2506 (N_2506,N_2288,N_2203);
and U2507 (N_2507,N_2005,N_2213);
and U2508 (N_2508,N_2297,N_2190);
nand U2509 (N_2509,N_2432,N_2391);
nand U2510 (N_2510,N_2184,N_2017);
nor U2511 (N_2511,N_2076,N_2386);
nand U2512 (N_2512,N_2188,N_2434);
xnor U2513 (N_2513,N_2283,N_2322);
or U2514 (N_2514,N_2113,N_2117);
nand U2515 (N_2515,N_2115,N_2032);
nand U2516 (N_2516,N_2426,N_2130);
nor U2517 (N_2517,N_2157,N_2300);
or U2518 (N_2518,N_2205,N_2294);
and U2519 (N_2519,N_2422,N_2202);
nand U2520 (N_2520,N_2015,N_2372);
and U2521 (N_2521,N_2178,N_2354);
nor U2522 (N_2522,N_2067,N_2256);
nor U2523 (N_2523,N_2233,N_2482);
nand U2524 (N_2524,N_2065,N_2116);
or U2525 (N_2525,N_2247,N_2468);
nor U2526 (N_2526,N_2445,N_2104);
xor U2527 (N_2527,N_2201,N_2086);
nand U2528 (N_2528,N_2061,N_2244);
nor U2529 (N_2529,N_2438,N_2403);
and U2530 (N_2530,N_2339,N_2395);
or U2531 (N_2531,N_2143,N_2041);
or U2532 (N_2532,N_2142,N_2436);
or U2533 (N_2533,N_2320,N_2364);
nor U2534 (N_2534,N_2087,N_2016);
or U2535 (N_2535,N_2165,N_2211);
xnor U2536 (N_2536,N_2088,N_2228);
or U2537 (N_2537,N_2410,N_2057);
or U2538 (N_2538,N_2359,N_2132);
xor U2539 (N_2539,N_2160,N_2030);
nand U2540 (N_2540,N_2136,N_2199);
nand U2541 (N_2541,N_2207,N_2192);
and U2542 (N_2542,N_2266,N_2350);
or U2543 (N_2543,N_2133,N_2053);
nand U2544 (N_2544,N_2457,N_2357);
nand U2545 (N_2545,N_2384,N_2271);
nand U2546 (N_2546,N_2295,N_2062);
and U2547 (N_2547,N_2109,N_2236);
nor U2548 (N_2548,N_2147,N_2382);
and U2549 (N_2549,N_2006,N_2170);
nor U2550 (N_2550,N_2011,N_2269);
or U2551 (N_2551,N_2282,N_2416);
and U2552 (N_2552,N_2361,N_2388);
nor U2553 (N_2553,N_2024,N_2358);
and U2554 (N_2554,N_2253,N_2325);
xor U2555 (N_2555,N_2135,N_2013);
nor U2556 (N_2556,N_2314,N_2012);
nor U2557 (N_2557,N_2027,N_2083);
or U2558 (N_2558,N_2007,N_2186);
and U2559 (N_2559,N_2345,N_2366);
and U2560 (N_2560,N_2383,N_2260);
nor U2561 (N_2561,N_2490,N_2450);
and U2562 (N_2562,N_2368,N_2210);
xor U2563 (N_2563,N_2235,N_2324);
or U2564 (N_2564,N_2491,N_2352);
nor U2565 (N_2565,N_2270,N_2347);
nand U2566 (N_2566,N_2209,N_2315);
xnor U2567 (N_2567,N_2101,N_2274);
or U2568 (N_2568,N_2499,N_2097);
or U2569 (N_2569,N_2159,N_2498);
or U2570 (N_2570,N_2050,N_2318);
or U2571 (N_2571,N_2477,N_2289);
nand U2572 (N_2572,N_2028,N_2483);
nor U2573 (N_2573,N_2363,N_2250);
nor U2574 (N_2574,N_2390,N_2066);
and U2575 (N_2575,N_2185,N_2268);
and U2576 (N_2576,N_2375,N_2279);
nand U2577 (N_2577,N_2068,N_2313);
or U2578 (N_2578,N_2037,N_2112);
nand U2579 (N_2579,N_2331,N_2461);
nand U2580 (N_2580,N_2038,N_2129);
xor U2581 (N_2581,N_2049,N_2411);
or U2582 (N_2582,N_2355,N_2340);
nand U2583 (N_2583,N_2231,N_2310);
nor U2584 (N_2584,N_2082,N_2342);
nor U2585 (N_2585,N_2304,N_2029);
or U2586 (N_2586,N_2400,N_2127);
nor U2587 (N_2587,N_2423,N_2153);
nor U2588 (N_2588,N_2173,N_2177);
xnor U2589 (N_2589,N_2328,N_2452);
or U2590 (N_2590,N_2240,N_2196);
nand U2591 (N_2591,N_2385,N_2470);
or U2592 (N_2592,N_2077,N_2369);
or U2593 (N_2593,N_2371,N_2446);
xnor U2594 (N_2594,N_2154,N_2149);
nor U2595 (N_2595,N_2220,N_2281);
or U2596 (N_2596,N_2481,N_2084);
nor U2597 (N_2597,N_2280,N_2316);
or U2598 (N_2598,N_2290,N_2025);
xor U2599 (N_2599,N_2152,N_2332);
or U2600 (N_2600,N_2431,N_2487);
or U2601 (N_2601,N_2493,N_2413);
and U2602 (N_2602,N_2380,N_2081);
and U2603 (N_2603,N_2485,N_2248);
nor U2604 (N_2604,N_2180,N_2484);
or U2605 (N_2605,N_2344,N_2150);
nand U2606 (N_2606,N_2258,N_2118);
nor U2607 (N_2607,N_2095,N_2141);
or U2608 (N_2608,N_2427,N_2000);
nand U2609 (N_2609,N_2401,N_2107);
and U2610 (N_2610,N_2351,N_2305);
nand U2611 (N_2611,N_2409,N_2198);
and U2612 (N_2612,N_2218,N_2040);
and U2613 (N_2613,N_2285,N_2467);
or U2614 (N_2614,N_2430,N_2321);
or U2615 (N_2615,N_2478,N_2343);
nor U2616 (N_2616,N_2175,N_2138);
and U2617 (N_2617,N_2408,N_2215);
and U2618 (N_2618,N_2064,N_2080);
xor U2619 (N_2619,N_2469,N_2058);
or U2620 (N_2620,N_2105,N_2302);
nor U2621 (N_2621,N_2089,N_2497);
and U2622 (N_2622,N_2022,N_2034);
or U2623 (N_2623,N_2075,N_2122);
nor U2624 (N_2624,N_2172,N_2412);
or U2625 (N_2625,N_2193,N_2241);
xor U2626 (N_2626,N_2214,N_2448);
and U2627 (N_2627,N_2148,N_2106);
nor U2628 (N_2628,N_2362,N_2301);
or U2629 (N_2629,N_2308,N_2287);
xor U2630 (N_2630,N_2039,N_2051);
or U2631 (N_2631,N_2216,N_2272);
nand U2632 (N_2632,N_2292,N_2415);
and U2633 (N_2633,N_2488,N_2405);
and U2634 (N_2634,N_2229,N_2257);
and U2635 (N_2635,N_2496,N_2338);
nand U2636 (N_2636,N_2492,N_2458);
nor U2637 (N_2637,N_2335,N_2164);
or U2638 (N_2638,N_2168,N_2307);
xor U2639 (N_2639,N_2454,N_2181);
or U2640 (N_2640,N_2336,N_2046);
nor U2641 (N_2641,N_2045,N_2286);
nor U2642 (N_2642,N_2167,N_2219);
nor U2643 (N_2643,N_2365,N_2009);
xnor U2644 (N_2644,N_2451,N_2019);
nor U2645 (N_2645,N_2001,N_2134);
and U2646 (N_2646,N_2278,N_2381);
xnor U2647 (N_2647,N_2212,N_2123);
xnor U2648 (N_2648,N_2234,N_2495);
or U2649 (N_2649,N_2125,N_2230);
or U2650 (N_2650,N_2071,N_2402);
or U2651 (N_2651,N_2407,N_2245);
or U2652 (N_2652,N_2090,N_2174);
and U2653 (N_2653,N_2020,N_2428);
nor U2654 (N_2654,N_2182,N_2298);
nand U2655 (N_2655,N_2189,N_2333);
nand U2656 (N_2656,N_2254,N_2284);
or U2657 (N_2657,N_2311,N_2424);
or U2658 (N_2658,N_2474,N_2008);
nand U2659 (N_2659,N_2242,N_2486);
nand U2660 (N_2660,N_2440,N_2063);
xor U2661 (N_2661,N_2466,N_2393);
nand U2662 (N_2662,N_2479,N_2471);
and U2663 (N_2663,N_2070,N_2102);
and U2664 (N_2664,N_2158,N_2346);
nor U2665 (N_2665,N_2093,N_2033);
nor U2666 (N_2666,N_2111,N_2464);
nor U2667 (N_2667,N_2026,N_2429);
nor U2668 (N_2668,N_2309,N_2303);
nand U2669 (N_2669,N_2096,N_2420);
nand U2670 (N_2670,N_2059,N_2387);
and U2671 (N_2671,N_2421,N_2223);
and U2672 (N_2672,N_2163,N_2267);
or U2673 (N_2673,N_2121,N_2246);
and U2674 (N_2674,N_2317,N_2124);
nand U2675 (N_2675,N_2264,N_2191);
nor U2676 (N_2676,N_2047,N_2463);
and U2677 (N_2677,N_2263,N_2378);
nor U2678 (N_2678,N_2265,N_2226);
and U2679 (N_2679,N_2225,N_2291);
xnor U2680 (N_2680,N_2156,N_2319);
nor U2681 (N_2681,N_2139,N_2161);
nand U2682 (N_2682,N_2444,N_2480);
or U2683 (N_2683,N_2389,N_2100);
nor U2684 (N_2684,N_2055,N_2334);
nor U2685 (N_2685,N_2373,N_2459);
and U2686 (N_2686,N_2072,N_2473);
xnor U2687 (N_2687,N_2277,N_2074);
or U2688 (N_2688,N_2098,N_2255);
nand U2689 (N_2689,N_2262,N_2069);
and U2690 (N_2690,N_2453,N_2085);
nand U2691 (N_2691,N_2146,N_2078);
and U2692 (N_2692,N_2128,N_2460);
or U2693 (N_2693,N_2010,N_2273);
nor U2694 (N_2694,N_2323,N_2194);
xor U2695 (N_2695,N_2406,N_2447);
and U2696 (N_2696,N_2054,N_2224);
or U2697 (N_2697,N_2103,N_2433);
or U2698 (N_2698,N_2494,N_2036);
nor U2699 (N_2699,N_2261,N_2394);
and U2700 (N_2700,N_2462,N_2023);
xor U2701 (N_2701,N_2419,N_2243);
nand U2702 (N_2702,N_2370,N_2425);
nor U2703 (N_2703,N_2204,N_2014);
and U2704 (N_2704,N_2079,N_2035);
or U2705 (N_2705,N_2360,N_2353);
or U2706 (N_2706,N_2042,N_2099);
or U2707 (N_2707,N_2221,N_2465);
nor U2708 (N_2708,N_2404,N_2208);
nor U2709 (N_2709,N_2217,N_2004);
or U2710 (N_2710,N_2238,N_2326);
nand U2711 (N_2711,N_2414,N_2144);
nor U2712 (N_2712,N_2043,N_2151);
and U2713 (N_2713,N_2443,N_2252);
or U2714 (N_2714,N_2417,N_2439);
nand U2715 (N_2715,N_2183,N_2187);
nor U2716 (N_2716,N_2299,N_2155);
xnor U2717 (N_2717,N_2048,N_2327);
or U2718 (N_2718,N_2031,N_2162);
and U2719 (N_2719,N_2349,N_2251);
or U2720 (N_2720,N_2021,N_2435);
and U2721 (N_2721,N_2094,N_2293);
and U2722 (N_2722,N_2126,N_2222);
or U2723 (N_2723,N_2108,N_2449);
nand U2724 (N_2724,N_2169,N_2476);
nand U2725 (N_2725,N_2249,N_2206);
nand U2726 (N_2726,N_2455,N_2239);
nor U2727 (N_2727,N_2137,N_2171);
nand U2728 (N_2728,N_2166,N_2356);
nor U2729 (N_2729,N_2197,N_2312);
nand U2730 (N_2730,N_2306,N_2398);
nor U2731 (N_2731,N_2018,N_2119);
nor U2732 (N_2732,N_2092,N_2227);
and U2733 (N_2733,N_2237,N_2060);
nand U2734 (N_2734,N_2329,N_2489);
and U2735 (N_2735,N_2437,N_2379);
or U2736 (N_2736,N_2348,N_2179);
nand U2737 (N_2737,N_2140,N_2232);
nor U2738 (N_2738,N_2052,N_2114);
and U2739 (N_2739,N_2456,N_2275);
nand U2740 (N_2740,N_2399,N_2330);
xor U2741 (N_2741,N_2296,N_2337);
or U2742 (N_2742,N_2396,N_2441);
or U2743 (N_2743,N_2176,N_2131);
nor U2744 (N_2744,N_2073,N_2200);
nor U2745 (N_2745,N_2195,N_2120);
nor U2746 (N_2746,N_2044,N_2442);
xnor U2747 (N_2747,N_2276,N_2475);
or U2748 (N_2748,N_2341,N_2397);
nor U2749 (N_2749,N_2003,N_2377);
nor U2750 (N_2750,N_2036,N_2484);
xor U2751 (N_2751,N_2448,N_2105);
nor U2752 (N_2752,N_2052,N_2204);
nand U2753 (N_2753,N_2372,N_2383);
xor U2754 (N_2754,N_2020,N_2396);
nor U2755 (N_2755,N_2464,N_2197);
or U2756 (N_2756,N_2008,N_2454);
or U2757 (N_2757,N_2068,N_2181);
nand U2758 (N_2758,N_2161,N_2280);
xor U2759 (N_2759,N_2263,N_2072);
and U2760 (N_2760,N_2124,N_2228);
xnor U2761 (N_2761,N_2078,N_2153);
and U2762 (N_2762,N_2393,N_2264);
nor U2763 (N_2763,N_2041,N_2244);
and U2764 (N_2764,N_2286,N_2459);
nor U2765 (N_2765,N_2233,N_2278);
or U2766 (N_2766,N_2261,N_2129);
nor U2767 (N_2767,N_2459,N_2357);
nor U2768 (N_2768,N_2453,N_2278);
nor U2769 (N_2769,N_2496,N_2347);
nand U2770 (N_2770,N_2420,N_2147);
and U2771 (N_2771,N_2115,N_2024);
or U2772 (N_2772,N_2375,N_2466);
xnor U2773 (N_2773,N_2163,N_2264);
nor U2774 (N_2774,N_2461,N_2338);
nor U2775 (N_2775,N_2003,N_2075);
nand U2776 (N_2776,N_2304,N_2162);
nor U2777 (N_2777,N_2214,N_2000);
xor U2778 (N_2778,N_2392,N_2065);
nand U2779 (N_2779,N_2483,N_2187);
nand U2780 (N_2780,N_2312,N_2042);
xor U2781 (N_2781,N_2223,N_2080);
nor U2782 (N_2782,N_2443,N_2356);
xor U2783 (N_2783,N_2103,N_2203);
and U2784 (N_2784,N_2305,N_2496);
nor U2785 (N_2785,N_2225,N_2379);
or U2786 (N_2786,N_2474,N_2187);
and U2787 (N_2787,N_2252,N_2422);
nor U2788 (N_2788,N_2137,N_2190);
nand U2789 (N_2789,N_2156,N_2475);
xnor U2790 (N_2790,N_2412,N_2408);
xor U2791 (N_2791,N_2016,N_2208);
xnor U2792 (N_2792,N_2412,N_2332);
or U2793 (N_2793,N_2430,N_2119);
xnor U2794 (N_2794,N_2043,N_2009);
nor U2795 (N_2795,N_2111,N_2154);
or U2796 (N_2796,N_2109,N_2427);
or U2797 (N_2797,N_2274,N_2163);
nor U2798 (N_2798,N_2164,N_2352);
nor U2799 (N_2799,N_2206,N_2496);
and U2800 (N_2800,N_2330,N_2436);
nor U2801 (N_2801,N_2201,N_2025);
and U2802 (N_2802,N_2180,N_2120);
or U2803 (N_2803,N_2344,N_2440);
xor U2804 (N_2804,N_2319,N_2228);
or U2805 (N_2805,N_2007,N_2371);
nor U2806 (N_2806,N_2006,N_2411);
and U2807 (N_2807,N_2262,N_2426);
or U2808 (N_2808,N_2183,N_2017);
nand U2809 (N_2809,N_2194,N_2248);
and U2810 (N_2810,N_2369,N_2243);
or U2811 (N_2811,N_2471,N_2200);
and U2812 (N_2812,N_2315,N_2262);
nor U2813 (N_2813,N_2387,N_2318);
nand U2814 (N_2814,N_2487,N_2002);
nor U2815 (N_2815,N_2479,N_2161);
or U2816 (N_2816,N_2026,N_2218);
nand U2817 (N_2817,N_2031,N_2024);
nand U2818 (N_2818,N_2338,N_2392);
nor U2819 (N_2819,N_2263,N_2133);
or U2820 (N_2820,N_2047,N_2205);
nor U2821 (N_2821,N_2471,N_2010);
nand U2822 (N_2822,N_2346,N_2197);
or U2823 (N_2823,N_2018,N_2159);
xor U2824 (N_2824,N_2009,N_2013);
or U2825 (N_2825,N_2137,N_2478);
nand U2826 (N_2826,N_2186,N_2032);
and U2827 (N_2827,N_2003,N_2336);
or U2828 (N_2828,N_2218,N_2058);
and U2829 (N_2829,N_2264,N_2489);
nor U2830 (N_2830,N_2427,N_2426);
nor U2831 (N_2831,N_2102,N_2455);
and U2832 (N_2832,N_2320,N_2409);
nor U2833 (N_2833,N_2182,N_2187);
xnor U2834 (N_2834,N_2208,N_2212);
and U2835 (N_2835,N_2034,N_2044);
nor U2836 (N_2836,N_2258,N_2482);
nand U2837 (N_2837,N_2397,N_2335);
and U2838 (N_2838,N_2046,N_2237);
or U2839 (N_2839,N_2477,N_2220);
nor U2840 (N_2840,N_2058,N_2333);
nand U2841 (N_2841,N_2164,N_2478);
nor U2842 (N_2842,N_2336,N_2467);
and U2843 (N_2843,N_2222,N_2382);
nand U2844 (N_2844,N_2241,N_2447);
nand U2845 (N_2845,N_2044,N_2426);
nor U2846 (N_2846,N_2178,N_2452);
and U2847 (N_2847,N_2368,N_2273);
or U2848 (N_2848,N_2171,N_2069);
and U2849 (N_2849,N_2183,N_2382);
and U2850 (N_2850,N_2394,N_2040);
nor U2851 (N_2851,N_2252,N_2292);
xor U2852 (N_2852,N_2358,N_2202);
nor U2853 (N_2853,N_2225,N_2088);
xor U2854 (N_2854,N_2285,N_2187);
or U2855 (N_2855,N_2362,N_2380);
or U2856 (N_2856,N_2045,N_2104);
and U2857 (N_2857,N_2438,N_2180);
nor U2858 (N_2858,N_2242,N_2285);
nor U2859 (N_2859,N_2296,N_2273);
and U2860 (N_2860,N_2320,N_2352);
nor U2861 (N_2861,N_2180,N_2347);
nand U2862 (N_2862,N_2477,N_2488);
nor U2863 (N_2863,N_2102,N_2319);
xnor U2864 (N_2864,N_2298,N_2170);
nand U2865 (N_2865,N_2266,N_2404);
and U2866 (N_2866,N_2262,N_2445);
nor U2867 (N_2867,N_2277,N_2046);
nand U2868 (N_2868,N_2140,N_2396);
nor U2869 (N_2869,N_2373,N_2104);
nor U2870 (N_2870,N_2189,N_2198);
or U2871 (N_2871,N_2401,N_2007);
nand U2872 (N_2872,N_2327,N_2140);
nor U2873 (N_2873,N_2173,N_2171);
and U2874 (N_2874,N_2152,N_2100);
xor U2875 (N_2875,N_2133,N_2271);
nand U2876 (N_2876,N_2117,N_2118);
nand U2877 (N_2877,N_2163,N_2273);
nand U2878 (N_2878,N_2423,N_2048);
or U2879 (N_2879,N_2071,N_2049);
or U2880 (N_2880,N_2367,N_2095);
nor U2881 (N_2881,N_2464,N_2127);
or U2882 (N_2882,N_2421,N_2462);
and U2883 (N_2883,N_2082,N_2189);
or U2884 (N_2884,N_2325,N_2260);
nor U2885 (N_2885,N_2380,N_2321);
or U2886 (N_2886,N_2241,N_2439);
nand U2887 (N_2887,N_2314,N_2299);
nand U2888 (N_2888,N_2449,N_2164);
or U2889 (N_2889,N_2155,N_2340);
nor U2890 (N_2890,N_2195,N_2402);
or U2891 (N_2891,N_2002,N_2177);
nand U2892 (N_2892,N_2257,N_2389);
or U2893 (N_2893,N_2075,N_2135);
nor U2894 (N_2894,N_2303,N_2287);
and U2895 (N_2895,N_2226,N_2464);
or U2896 (N_2896,N_2372,N_2361);
and U2897 (N_2897,N_2277,N_2077);
nor U2898 (N_2898,N_2313,N_2292);
and U2899 (N_2899,N_2208,N_2479);
and U2900 (N_2900,N_2115,N_2392);
and U2901 (N_2901,N_2299,N_2364);
nand U2902 (N_2902,N_2449,N_2488);
nor U2903 (N_2903,N_2272,N_2328);
nand U2904 (N_2904,N_2290,N_2268);
nor U2905 (N_2905,N_2353,N_2277);
nand U2906 (N_2906,N_2324,N_2297);
nand U2907 (N_2907,N_2153,N_2489);
nor U2908 (N_2908,N_2163,N_2106);
nor U2909 (N_2909,N_2244,N_2418);
xor U2910 (N_2910,N_2176,N_2367);
xnor U2911 (N_2911,N_2226,N_2470);
or U2912 (N_2912,N_2353,N_2257);
nand U2913 (N_2913,N_2409,N_2348);
xnor U2914 (N_2914,N_2428,N_2445);
and U2915 (N_2915,N_2059,N_2051);
or U2916 (N_2916,N_2052,N_2110);
xnor U2917 (N_2917,N_2397,N_2300);
and U2918 (N_2918,N_2201,N_2042);
nor U2919 (N_2919,N_2085,N_2385);
or U2920 (N_2920,N_2132,N_2212);
nand U2921 (N_2921,N_2106,N_2409);
nand U2922 (N_2922,N_2109,N_2371);
nor U2923 (N_2923,N_2410,N_2212);
or U2924 (N_2924,N_2128,N_2175);
or U2925 (N_2925,N_2327,N_2306);
and U2926 (N_2926,N_2130,N_2242);
or U2927 (N_2927,N_2304,N_2099);
xor U2928 (N_2928,N_2454,N_2164);
nor U2929 (N_2929,N_2167,N_2339);
nor U2930 (N_2930,N_2401,N_2475);
or U2931 (N_2931,N_2001,N_2295);
nand U2932 (N_2932,N_2339,N_2075);
nand U2933 (N_2933,N_2438,N_2241);
nand U2934 (N_2934,N_2207,N_2457);
nor U2935 (N_2935,N_2329,N_2052);
nor U2936 (N_2936,N_2495,N_2156);
and U2937 (N_2937,N_2267,N_2183);
nand U2938 (N_2938,N_2396,N_2378);
and U2939 (N_2939,N_2144,N_2486);
nor U2940 (N_2940,N_2388,N_2349);
nor U2941 (N_2941,N_2285,N_2331);
nand U2942 (N_2942,N_2269,N_2475);
xor U2943 (N_2943,N_2398,N_2290);
and U2944 (N_2944,N_2048,N_2148);
xnor U2945 (N_2945,N_2063,N_2191);
nor U2946 (N_2946,N_2219,N_2240);
nor U2947 (N_2947,N_2467,N_2083);
nor U2948 (N_2948,N_2002,N_2173);
and U2949 (N_2949,N_2064,N_2288);
xnor U2950 (N_2950,N_2359,N_2007);
and U2951 (N_2951,N_2128,N_2368);
or U2952 (N_2952,N_2437,N_2407);
nand U2953 (N_2953,N_2135,N_2100);
nor U2954 (N_2954,N_2204,N_2189);
nor U2955 (N_2955,N_2199,N_2053);
nand U2956 (N_2956,N_2176,N_2450);
and U2957 (N_2957,N_2030,N_2185);
xnor U2958 (N_2958,N_2378,N_2274);
and U2959 (N_2959,N_2245,N_2250);
or U2960 (N_2960,N_2001,N_2393);
xor U2961 (N_2961,N_2147,N_2497);
nand U2962 (N_2962,N_2300,N_2286);
nand U2963 (N_2963,N_2443,N_2362);
and U2964 (N_2964,N_2340,N_2297);
and U2965 (N_2965,N_2386,N_2411);
and U2966 (N_2966,N_2472,N_2117);
or U2967 (N_2967,N_2350,N_2299);
and U2968 (N_2968,N_2075,N_2140);
and U2969 (N_2969,N_2278,N_2254);
xnor U2970 (N_2970,N_2344,N_2118);
or U2971 (N_2971,N_2284,N_2128);
nand U2972 (N_2972,N_2337,N_2387);
and U2973 (N_2973,N_2445,N_2140);
nand U2974 (N_2974,N_2303,N_2377);
or U2975 (N_2975,N_2072,N_2153);
nand U2976 (N_2976,N_2148,N_2041);
nand U2977 (N_2977,N_2223,N_2009);
and U2978 (N_2978,N_2495,N_2466);
and U2979 (N_2979,N_2148,N_2056);
nand U2980 (N_2980,N_2107,N_2270);
nor U2981 (N_2981,N_2143,N_2230);
xnor U2982 (N_2982,N_2139,N_2043);
nand U2983 (N_2983,N_2213,N_2080);
or U2984 (N_2984,N_2180,N_2190);
or U2985 (N_2985,N_2163,N_2418);
nand U2986 (N_2986,N_2352,N_2259);
and U2987 (N_2987,N_2019,N_2307);
nand U2988 (N_2988,N_2274,N_2341);
nor U2989 (N_2989,N_2130,N_2340);
nor U2990 (N_2990,N_2201,N_2333);
nand U2991 (N_2991,N_2461,N_2254);
and U2992 (N_2992,N_2466,N_2088);
or U2993 (N_2993,N_2227,N_2246);
xor U2994 (N_2994,N_2240,N_2143);
nor U2995 (N_2995,N_2029,N_2257);
nor U2996 (N_2996,N_2475,N_2480);
nand U2997 (N_2997,N_2266,N_2487);
nand U2998 (N_2998,N_2447,N_2231);
nor U2999 (N_2999,N_2314,N_2009);
nand U3000 (N_3000,N_2681,N_2641);
nor U3001 (N_3001,N_2543,N_2520);
and U3002 (N_3002,N_2845,N_2966);
or U3003 (N_3003,N_2531,N_2889);
or U3004 (N_3004,N_2776,N_2713);
and U3005 (N_3005,N_2784,N_2545);
xor U3006 (N_3006,N_2977,N_2636);
nor U3007 (N_3007,N_2563,N_2710);
nor U3008 (N_3008,N_2518,N_2555);
or U3009 (N_3009,N_2558,N_2647);
nor U3010 (N_3010,N_2975,N_2799);
nor U3011 (N_3011,N_2901,N_2706);
nor U3012 (N_3012,N_2753,N_2965);
or U3013 (N_3013,N_2870,N_2691);
nor U3014 (N_3014,N_2742,N_2831);
or U3015 (N_3015,N_2622,N_2868);
and U3016 (N_3016,N_2628,N_2662);
and U3017 (N_3017,N_2639,N_2572);
and U3018 (N_3018,N_2697,N_2803);
and U3019 (N_3019,N_2653,N_2967);
or U3020 (N_3020,N_2733,N_2943);
or U3021 (N_3021,N_2738,N_2542);
nor U3022 (N_3022,N_2729,N_2552);
nor U3023 (N_3023,N_2727,N_2813);
and U3024 (N_3024,N_2817,N_2587);
or U3025 (N_3025,N_2728,N_2880);
nand U3026 (N_3026,N_2856,N_2719);
xnor U3027 (N_3027,N_2948,N_2834);
nor U3028 (N_3028,N_2841,N_2758);
or U3029 (N_3029,N_2933,N_2707);
xor U3030 (N_3030,N_2862,N_2582);
and U3031 (N_3031,N_2819,N_2785);
nand U3032 (N_3032,N_2617,N_2839);
or U3033 (N_3033,N_2867,N_2940);
or U3034 (N_3034,N_2743,N_2594);
and U3035 (N_3035,N_2593,N_2954);
nand U3036 (N_3036,N_2741,N_2995);
nand U3037 (N_3037,N_2693,N_2579);
nand U3038 (N_3038,N_2575,N_2698);
nand U3039 (N_3039,N_2771,N_2649);
or U3040 (N_3040,N_2704,N_2844);
or U3041 (N_3041,N_2765,N_2999);
nor U3042 (N_3042,N_2757,N_2983);
and U3043 (N_3043,N_2692,N_2723);
and U3044 (N_3044,N_2936,N_2953);
or U3045 (N_3045,N_2956,N_2915);
nor U3046 (N_3046,N_2985,N_2567);
xnor U3047 (N_3047,N_2506,N_2778);
or U3048 (N_3048,N_2529,N_2926);
and U3049 (N_3049,N_2873,N_2525);
or U3050 (N_3050,N_2871,N_2686);
xnor U3051 (N_3051,N_2960,N_2809);
nor U3052 (N_3052,N_2625,N_2610);
xnor U3053 (N_3053,N_2554,N_2774);
or U3054 (N_3054,N_2508,N_2749);
nand U3055 (N_3055,N_2672,N_2634);
xnor U3056 (N_3056,N_2800,N_2802);
xnor U3057 (N_3057,N_2604,N_2703);
nor U3058 (N_3058,N_2951,N_2937);
nor U3059 (N_3059,N_2860,N_2551);
nand U3060 (N_3060,N_2827,N_2928);
and U3061 (N_3061,N_2602,N_2516);
and U3062 (N_3062,N_2919,N_2761);
nand U3063 (N_3063,N_2524,N_2509);
nand U3064 (N_3064,N_2671,N_2872);
and U3065 (N_3065,N_2734,N_2925);
xor U3066 (N_3066,N_2996,N_2833);
and U3067 (N_3067,N_2846,N_2557);
nor U3068 (N_3068,N_2592,N_2623);
nand U3069 (N_3069,N_2890,N_2961);
nor U3070 (N_3070,N_2984,N_2882);
and U3071 (N_3071,N_2934,N_2796);
and U3072 (N_3072,N_2705,N_2869);
nand U3073 (N_3073,N_2964,N_2777);
and U3074 (N_3074,N_2603,N_2565);
nand U3075 (N_3075,N_2535,N_2665);
nor U3076 (N_3076,N_2682,N_2709);
and U3077 (N_3077,N_2849,N_2945);
nor U3078 (N_3078,N_2721,N_2621);
or U3079 (N_3079,N_2807,N_2614);
nor U3080 (N_3080,N_2998,N_2988);
and U3081 (N_3081,N_2585,N_2790);
and U3082 (N_3082,N_2752,N_2675);
xnor U3083 (N_3083,N_2981,N_2549);
nand U3084 (N_3084,N_2982,N_2989);
nand U3085 (N_3085,N_2566,N_2787);
or U3086 (N_3086,N_2969,N_2657);
or U3087 (N_3087,N_2938,N_2895);
or U3088 (N_3088,N_2608,N_2972);
or U3089 (N_3089,N_2583,N_2611);
nand U3090 (N_3090,N_2883,N_2644);
nand U3091 (N_3091,N_2576,N_2892);
and U3092 (N_3092,N_2921,N_2843);
or U3093 (N_3093,N_2795,N_2929);
and U3094 (N_3094,N_2842,N_2650);
or U3095 (N_3095,N_2789,N_2801);
xor U3096 (N_3096,N_2864,N_2505);
or U3097 (N_3097,N_2651,N_2976);
xnor U3098 (N_3098,N_2922,N_2768);
and U3099 (N_3099,N_2523,N_2854);
nor U3100 (N_3100,N_2927,N_2772);
nand U3101 (N_3101,N_2595,N_2917);
nand U3102 (N_3102,N_2627,N_2923);
nand U3103 (N_3103,N_2910,N_2640);
xor U3104 (N_3104,N_2823,N_2720);
nor U3105 (N_3105,N_2687,N_2852);
nor U3106 (N_3106,N_2820,N_2855);
xor U3107 (N_3107,N_2577,N_2537);
xor U3108 (N_3108,N_2737,N_2599);
nor U3109 (N_3109,N_2712,N_2539);
and U3110 (N_3110,N_2600,N_2673);
and U3111 (N_3111,N_2755,N_2994);
nand U3112 (N_3112,N_2835,N_2955);
and U3113 (N_3113,N_2732,N_2909);
and U3114 (N_3114,N_2638,N_2830);
or U3115 (N_3115,N_2971,N_2946);
and U3116 (N_3116,N_2797,N_2679);
nor U3117 (N_3117,N_2747,N_2837);
and U3118 (N_3118,N_2760,N_2824);
nor U3119 (N_3119,N_2782,N_2898);
nand U3120 (N_3120,N_2918,N_2502);
and U3121 (N_3121,N_2788,N_2533);
or U3122 (N_3122,N_2962,N_2891);
xor U3123 (N_3123,N_2958,N_2896);
or U3124 (N_3124,N_2979,N_2596);
and U3125 (N_3125,N_2810,N_2974);
nand U3126 (N_3126,N_2884,N_2805);
and U3127 (N_3127,N_2521,N_2877);
nand U3128 (N_3128,N_2798,N_2536);
nor U3129 (N_3129,N_2916,N_2781);
nor U3130 (N_3130,N_2526,N_2993);
xor U3131 (N_3131,N_2735,N_2661);
nand U3132 (N_3132,N_2847,N_2806);
nor U3133 (N_3133,N_2875,N_2851);
or U3134 (N_3134,N_2818,N_2822);
nor U3135 (N_3135,N_2540,N_2598);
or U3136 (N_3136,N_2793,N_2894);
xor U3137 (N_3137,N_2762,N_2730);
nand U3138 (N_3138,N_2514,N_2689);
or U3139 (N_3139,N_2553,N_2808);
nor U3140 (N_3140,N_2786,N_2652);
nand U3141 (N_3141,N_2659,N_2930);
and U3142 (N_3142,N_2511,N_2838);
and U3143 (N_3143,N_2694,N_2544);
nor U3144 (N_3144,N_2571,N_2668);
and U3145 (N_3145,N_2522,N_2631);
xnor U3146 (N_3146,N_2804,N_2538);
nor U3147 (N_3147,N_2914,N_2912);
or U3148 (N_3148,N_2547,N_2669);
xnor U3149 (N_3149,N_2612,N_2950);
nor U3150 (N_3150,N_2885,N_2708);
nor U3151 (N_3151,N_2897,N_2646);
nand U3152 (N_3152,N_2766,N_2811);
or U3153 (N_3153,N_2767,N_2968);
nand U3154 (N_3154,N_2980,N_2913);
or U3155 (N_3155,N_2939,N_2501);
nand U3156 (N_3156,N_2590,N_2601);
xor U3157 (N_3157,N_2959,N_2941);
nor U3158 (N_3158,N_2648,N_2597);
nor U3159 (N_3159,N_2534,N_2635);
and U3160 (N_3160,N_2680,N_2722);
nor U3161 (N_3161,N_2826,N_2836);
or U3162 (N_3162,N_2740,N_2548);
and U3163 (N_3163,N_2857,N_2556);
nand U3164 (N_3164,N_2792,N_2908);
and U3165 (N_3165,N_2863,N_2986);
nor U3166 (N_3166,N_2683,N_2911);
or U3167 (N_3167,N_2580,N_2699);
and U3168 (N_3168,N_2739,N_2530);
nor U3169 (N_3169,N_2702,N_2899);
and U3170 (N_3170,N_2773,N_2578);
and U3171 (N_3171,N_2828,N_2783);
nand U3172 (N_3172,N_2903,N_2658);
or U3173 (N_3173,N_2952,N_2568);
nand U3174 (N_3174,N_2620,N_2716);
nor U3175 (N_3175,N_2715,N_2920);
and U3176 (N_3176,N_2666,N_2717);
nor U3177 (N_3177,N_2931,N_2814);
xnor U3178 (N_3178,N_2527,N_2550);
nand U3179 (N_3179,N_2677,N_2748);
nor U3180 (N_3180,N_2678,N_2512);
nor U3181 (N_3181,N_2858,N_2987);
nor U3182 (N_3182,N_2656,N_2606);
or U3183 (N_3183,N_2581,N_2670);
and U3184 (N_3184,N_2637,N_2750);
or U3185 (N_3185,N_2812,N_2779);
or U3186 (N_3186,N_2688,N_2645);
nand U3187 (N_3187,N_2724,N_2907);
and U3188 (N_3188,N_2624,N_2667);
nor U3189 (N_3189,N_2564,N_2924);
or U3190 (N_3190,N_2725,N_2500);
nor U3191 (N_3191,N_2881,N_2629);
nand U3192 (N_3192,N_2850,N_2609);
nand U3193 (N_3193,N_2840,N_2906);
nand U3194 (N_3194,N_2584,N_2643);
and U3195 (N_3195,N_2570,N_2978);
nand U3196 (N_3196,N_2507,N_2949);
or U3197 (N_3197,N_2775,N_2701);
nor U3198 (N_3198,N_2973,N_2888);
and U3199 (N_3199,N_2944,N_2886);
and U3200 (N_3200,N_2794,N_2700);
and U3201 (N_3201,N_2562,N_2791);
or U3202 (N_3202,N_2992,N_2588);
or U3203 (N_3203,N_2780,N_2696);
nand U3204 (N_3204,N_2726,N_2654);
nand U3205 (N_3205,N_2660,N_2902);
nor U3206 (N_3206,N_2821,N_2893);
nor U3207 (N_3207,N_2859,N_2997);
and U3208 (N_3208,N_2685,N_2561);
or U3209 (N_3209,N_2630,N_2695);
or U3210 (N_3210,N_2589,N_2905);
or U3211 (N_3211,N_2816,N_2746);
xnor U3212 (N_3212,N_2528,N_2663);
and U3213 (N_3213,N_2744,N_2769);
xnor U3214 (N_3214,N_2866,N_2560);
nor U3215 (N_3215,N_2642,N_2756);
xnor U3216 (N_3216,N_2616,N_2947);
and U3217 (N_3217,N_2990,N_2676);
nand U3218 (N_3218,N_2879,N_2853);
or U3219 (N_3219,N_2613,N_2632);
nor U3220 (N_3220,N_2825,N_2605);
nand U3221 (N_3221,N_2626,N_2513);
and U3222 (N_3222,N_2754,N_2618);
nor U3223 (N_3223,N_2815,N_2559);
nand U3224 (N_3224,N_2770,N_2510);
nor U3225 (N_3225,N_2591,N_2569);
nor U3226 (N_3226,N_2684,N_2957);
nand U3227 (N_3227,N_2664,N_2764);
nand U3228 (N_3228,N_2848,N_2861);
nand U3229 (N_3229,N_2874,N_2546);
and U3230 (N_3230,N_2878,N_2718);
nand U3231 (N_3231,N_2731,N_2963);
and U3232 (N_3232,N_2745,N_2504);
or U3233 (N_3233,N_2532,N_2991);
and U3234 (N_3234,N_2900,N_2970);
and U3235 (N_3235,N_2876,N_2615);
nor U3236 (N_3236,N_2887,N_2714);
and U3237 (N_3237,N_2832,N_2541);
and U3238 (N_3238,N_2586,N_2904);
or U3239 (N_3239,N_2829,N_2515);
nand U3240 (N_3240,N_2759,N_2655);
or U3241 (N_3241,N_2633,N_2763);
and U3242 (N_3242,N_2517,N_2751);
xor U3243 (N_3243,N_2942,N_2865);
nand U3244 (N_3244,N_2932,N_2574);
or U3245 (N_3245,N_2736,N_2519);
nand U3246 (N_3246,N_2619,N_2607);
and U3247 (N_3247,N_2674,N_2711);
nand U3248 (N_3248,N_2573,N_2690);
nand U3249 (N_3249,N_2503,N_2935);
and U3250 (N_3250,N_2723,N_2668);
and U3251 (N_3251,N_2802,N_2805);
or U3252 (N_3252,N_2726,N_2722);
or U3253 (N_3253,N_2584,N_2508);
xnor U3254 (N_3254,N_2918,N_2629);
nor U3255 (N_3255,N_2888,N_2900);
nor U3256 (N_3256,N_2758,N_2540);
or U3257 (N_3257,N_2949,N_2503);
and U3258 (N_3258,N_2846,N_2941);
and U3259 (N_3259,N_2998,N_2575);
or U3260 (N_3260,N_2930,N_2731);
or U3261 (N_3261,N_2552,N_2659);
and U3262 (N_3262,N_2798,N_2972);
and U3263 (N_3263,N_2658,N_2828);
nand U3264 (N_3264,N_2784,N_2821);
or U3265 (N_3265,N_2861,N_2805);
nand U3266 (N_3266,N_2989,N_2904);
or U3267 (N_3267,N_2532,N_2701);
nor U3268 (N_3268,N_2802,N_2788);
xnor U3269 (N_3269,N_2879,N_2770);
or U3270 (N_3270,N_2749,N_2984);
and U3271 (N_3271,N_2582,N_2930);
or U3272 (N_3272,N_2998,N_2749);
or U3273 (N_3273,N_2710,N_2777);
nor U3274 (N_3274,N_2773,N_2736);
nand U3275 (N_3275,N_2792,N_2960);
nor U3276 (N_3276,N_2624,N_2567);
or U3277 (N_3277,N_2831,N_2829);
nand U3278 (N_3278,N_2572,N_2948);
or U3279 (N_3279,N_2628,N_2766);
and U3280 (N_3280,N_2747,N_2947);
and U3281 (N_3281,N_2818,N_2713);
nand U3282 (N_3282,N_2869,N_2936);
nor U3283 (N_3283,N_2956,N_2887);
xor U3284 (N_3284,N_2665,N_2619);
nor U3285 (N_3285,N_2569,N_2911);
or U3286 (N_3286,N_2877,N_2692);
nor U3287 (N_3287,N_2983,N_2799);
or U3288 (N_3288,N_2989,N_2959);
and U3289 (N_3289,N_2812,N_2600);
nand U3290 (N_3290,N_2890,N_2713);
and U3291 (N_3291,N_2597,N_2779);
nand U3292 (N_3292,N_2858,N_2738);
nand U3293 (N_3293,N_2861,N_2647);
xor U3294 (N_3294,N_2748,N_2982);
nand U3295 (N_3295,N_2887,N_2998);
or U3296 (N_3296,N_2958,N_2664);
nand U3297 (N_3297,N_2717,N_2841);
nor U3298 (N_3298,N_2830,N_2736);
and U3299 (N_3299,N_2905,N_2940);
and U3300 (N_3300,N_2696,N_2880);
nor U3301 (N_3301,N_2522,N_2934);
xor U3302 (N_3302,N_2713,N_2706);
and U3303 (N_3303,N_2763,N_2595);
and U3304 (N_3304,N_2630,N_2579);
and U3305 (N_3305,N_2672,N_2500);
nor U3306 (N_3306,N_2738,N_2811);
or U3307 (N_3307,N_2944,N_2760);
nand U3308 (N_3308,N_2795,N_2780);
nor U3309 (N_3309,N_2571,N_2903);
xnor U3310 (N_3310,N_2978,N_2787);
and U3311 (N_3311,N_2589,N_2563);
or U3312 (N_3312,N_2766,N_2617);
or U3313 (N_3313,N_2635,N_2606);
or U3314 (N_3314,N_2531,N_2945);
xnor U3315 (N_3315,N_2512,N_2936);
or U3316 (N_3316,N_2645,N_2976);
nor U3317 (N_3317,N_2531,N_2802);
or U3318 (N_3318,N_2741,N_2512);
and U3319 (N_3319,N_2541,N_2723);
or U3320 (N_3320,N_2734,N_2893);
or U3321 (N_3321,N_2611,N_2607);
or U3322 (N_3322,N_2733,N_2887);
or U3323 (N_3323,N_2677,N_2688);
nand U3324 (N_3324,N_2512,N_2676);
or U3325 (N_3325,N_2736,N_2965);
or U3326 (N_3326,N_2664,N_2945);
nor U3327 (N_3327,N_2710,N_2873);
nor U3328 (N_3328,N_2688,N_2906);
xnor U3329 (N_3329,N_2686,N_2506);
nand U3330 (N_3330,N_2769,N_2631);
nor U3331 (N_3331,N_2634,N_2669);
nor U3332 (N_3332,N_2519,N_2558);
or U3333 (N_3333,N_2612,N_2616);
or U3334 (N_3334,N_2747,N_2565);
or U3335 (N_3335,N_2529,N_2506);
or U3336 (N_3336,N_2994,N_2892);
nor U3337 (N_3337,N_2591,N_2664);
nand U3338 (N_3338,N_2968,N_2543);
and U3339 (N_3339,N_2558,N_2835);
and U3340 (N_3340,N_2710,N_2854);
nand U3341 (N_3341,N_2668,N_2946);
nor U3342 (N_3342,N_2524,N_2585);
nor U3343 (N_3343,N_2875,N_2962);
or U3344 (N_3344,N_2950,N_2626);
or U3345 (N_3345,N_2765,N_2506);
and U3346 (N_3346,N_2764,N_2603);
and U3347 (N_3347,N_2971,N_2605);
or U3348 (N_3348,N_2901,N_2829);
nor U3349 (N_3349,N_2550,N_2623);
nand U3350 (N_3350,N_2519,N_2588);
or U3351 (N_3351,N_2916,N_2676);
or U3352 (N_3352,N_2742,N_2655);
and U3353 (N_3353,N_2727,N_2520);
and U3354 (N_3354,N_2795,N_2735);
and U3355 (N_3355,N_2740,N_2665);
nand U3356 (N_3356,N_2816,N_2515);
nor U3357 (N_3357,N_2779,N_2571);
and U3358 (N_3358,N_2547,N_2770);
xnor U3359 (N_3359,N_2826,N_2914);
and U3360 (N_3360,N_2901,N_2659);
or U3361 (N_3361,N_2872,N_2682);
nor U3362 (N_3362,N_2758,N_2864);
nor U3363 (N_3363,N_2862,N_2628);
or U3364 (N_3364,N_2761,N_2883);
nand U3365 (N_3365,N_2989,N_2587);
nand U3366 (N_3366,N_2970,N_2770);
and U3367 (N_3367,N_2832,N_2746);
nor U3368 (N_3368,N_2772,N_2839);
and U3369 (N_3369,N_2953,N_2791);
nand U3370 (N_3370,N_2873,N_2741);
nor U3371 (N_3371,N_2929,N_2570);
nor U3372 (N_3372,N_2774,N_2729);
nand U3373 (N_3373,N_2599,N_2527);
and U3374 (N_3374,N_2633,N_2569);
nand U3375 (N_3375,N_2751,N_2838);
and U3376 (N_3376,N_2694,N_2992);
nor U3377 (N_3377,N_2657,N_2955);
and U3378 (N_3378,N_2748,N_2912);
and U3379 (N_3379,N_2852,N_2627);
nor U3380 (N_3380,N_2820,N_2758);
or U3381 (N_3381,N_2615,N_2959);
nand U3382 (N_3382,N_2734,N_2710);
xnor U3383 (N_3383,N_2544,N_2661);
nand U3384 (N_3384,N_2884,N_2591);
nor U3385 (N_3385,N_2826,N_2630);
nand U3386 (N_3386,N_2890,N_2949);
nor U3387 (N_3387,N_2865,N_2967);
nand U3388 (N_3388,N_2942,N_2813);
or U3389 (N_3389,N_2951,N_2688);
nor U3390 (N_3390,N_2581,N_2675);
nand U3391 (N_3391,N_2552,N_2685);
and U3392 (N_3392,N_2927,N_2729);
or U3393 (N_3393,N_2587,N_2857);
nand U3394 (N_3394,N_2547,N_2611);
or U3395 (N_3395,N_2883,N_2821);
nand U3396 (N_3396,N_2572,N_2710);
and U3397 (N_3397,N_2775,N_2754);
or U3398 (N_3398,N_2560,N_2892);
nor U3399 (N_3399,N_2817,N_2594);
nand U3400 (N_3400,N_2555,N_2927);
xor U3401 (N_3401,N_2582,N_2810);
nand U3402 (N_3402,N_2979,N_2804);
and U3403 (N_3403,N_2539,N_2630);
nand U3404 (N_3404,N_2827,N_2645);
and U3405 (N_3405,N_2960,N_2705);
or U3406 (N_3406,N_2775,N_2568);
nor U3407 (N_3407,N_2804,N_2545);
nor U3408 (N_3408,N_2888,N_2591);
nand U3409 (N_3409,N_2978,N_2578);
xnor U3410 (N_3410,N_2937,N_2822);
nor U3411 (N_3411,N_2734,N_2694);
nand U3412 (N_3412,N_2876,N_2865);
nor U3413 (N_3413,N_2580,N_2944);
xor U3414 (N_3414,N_2654,N_2501);
nand U3415 (N_3415,N_2943,N_2697);
and U3416 (N_3416,N_2827,N_2694);
or U3417 (N_3417,N_2808,N_2899);
xor U3418 (N_3418,N_2998,N_2928);
and U3419 (N_3419,N_2789,N_2838);
or U3420 (N_3420,N_2760,N_2560);
nand U3421 (N_3421,N_2572,N_2977);
or U3422 (N_3422,N_2903,N_2871);
and U3423 (N_3423,N_2853,N_2826);
nor U3424 (N_3424,N_2923,N_2977);
nor U3425 (N_3425,N_2518,N_2876);
nor U3426 (N_3426,N_2808,N_2858);
nand U3427 (N_3427,N_2883,N_2979);
or U3428 (N_3428,N_2590,N_2775);
xnor U3429 (N_3429,N_2742,N_2837);
and U3430 (N_3430,N_2520,N_2971);
nor U3431 (N_3431,N_2898,N_2518);
nand U3432 (N_3432,N_2695,N_2852);
nor U3433 (N_3433,N_2820,N_2609);
nand U3434 (N_3434,N_2896,N_2723);
nor U3435 (N_3435,N_2894,N_2849);
and U3436 (N_3436,N_2755,N_2626);
nor U3437 (N_3437,N_2909,N_2779);
nand U3438 (N_3438,N_2894,N_2586);
and U3439 (N_3439,N_2668,N_2616);
and U3440 (N_3440,N_2844,N_2880);
nor U3441 (N_3441,N_2892,N_2930);
nand U3442 (N_3442,N_2592,N_2868);
nand U3443 (N_3443,N_2844,N_2684);
and U3444 (N_3444,N_2695,N_2975);
or U3445 (N_3445,N_2571,N_2834);
or U3446 (N_3446,N_2916,N_2522);
nor U3447 (N_3447,N_2935,N_2773);
or U3448 (N_3448,N_2973,N_2537);
nor U3449 (N_3449,N_2729,N_2804);
nor U3450 (N_3450,N_2772,N_2999);
nand U3451 (N_3451,N_2693,N_2518);
nor U3452 (N_3452,N_2513,N_2699);
or U3453 (N_3453,N_2816,N_2640);
nand U3454 (N_3454,N_2942,N_2601);
nor U3455 (N_3455,N_2701,N_2769);
and U3456 (N_3456,N_2912,N_2649);
nor U3457 (N_3457,N_2639,N_2801);
nor U3458 (N_3458,N_2991,N_2911);
nor U3459 (N_3459,N_2903,N_2641);
or U3460 (N_3460,N_2685,N_2895);
or U3461 (N_3461,N_2750,N_2961);
nand U3462 (N_3462,N_2503,N_2739);
nor U3463 (N_3463,N_2829,N_2524);
nand U3464 (N_3464,N_2984,N_2761);
or U3465 (N_3465,N_2525,N_2632);
nor U3466 (N_3466,N_2647,N_2752);
or U3467 (N_3467,N_2883,N_2687);
and U3468 (N_3468,N_2772,N_2556);
or U3469 (N_3469,N_2674,N_2897);
or U3470 (N_3470,N_2617,N_2790);
and U3471 (N_3471,N_2585,N_2964);
nand U3472 (N_3472,N_2835,N_2627);
or U3473 (N_3473,N_2739,N_2994);
nor U3474 (N_3474,N_2896,N_2750);
nor U3475 (N_3475,N_2520,N_2909);
nor U3476 (N_3476,N_2767,N_2647);
nand U3477 (N_3477,N_2559,N_2925);
nor U3478 (N_3478,N_2990,N_2587);
nor U3479 (N_3479,N_2854,N_2814);
nor U3480 (N_3480,N_2850,N_2508);
nand U3481 (N_3481,N_2708,N_2997);
or U3482 (N_3482,N_2803,N_2658);
and U3483 (N_3483,N_2550,N_2581);
nor U3484 (N_3484,N_2722,N_2511);
nor U3485 (N_3485,N_2854,N_2567);
or U3486 (N_3486,N_2549,N_2816);
nor U3487 (N_3487,N_2653,N_2835);
nand U3488 (N_3488,N_2825,N_2980);
and U3489 (N_3489,N_2641,N_2700);
or U3490 (N_3490,N_2725,N_2869);
or U3491 (N_3491,N_2931,N_2993);
and U3492 (N_3492,N_2753,N_2943);
and U3493 (N_3493,N_2888,N_2717);
xnor U3494 (N_3494,N_2546,N_2526);
nand U3495 (N_3495,N_2742,N_2650);
and U3496 (N_3496,N_2769,N_2544);
and U3497 (N_3497,N_2967,N_2670);
or U3498 (N_3498,N_2843,N_2938);
and U3499 (N_3499,N_2573,N_2552);
xor U3500 (N_3500,N_3168,N_3219);
or U3501 (N_3501,N_3485,N_3013);
and U3502 (N_3502,N_3154,N_3398);
nor U3503 (N_3503,N_3489,N_3084);
and U3504 (N_3504,N_3425,N_3011);
xnor U3505 (N_3505,N_3263,N_3478);
nand U3506 (N_3506,N_3041,N_3271);
or U3507 (N_3507,N_3109,N_3407);
nand U3508 (N_3508,N_3225,N_3418);
or U3509 (N_3509,N_3309,N_3320);
nor U3510 (N_3510,N_3055,N_3172);
nor U3511 (N_3511,N_3188,N_3187);
and U3512 (N_3512,N_3260,N_3195);
nand U3513 (N_3513,N_3155,N_3242);
nand U3514 (N_3514,N_3295,N_3118);
xor U3515 (N_3515,N_3021,N_3427);
and U3516 (N_3516,N_3259,N_3361);
xor U3517 (N_3517,N_3341,N_3088);
xor U3518 (N_3518,N_3421,N_3467);
and U3519 (N_3519,N_3324,N_3032);
nand U3520 (N_3520,N_3076,N_3022);
nand U3521 (N_3521,N_3157,N_3357);
nand U3522 (N_3522,N_3001,N_3176);
nor U3523 (N_3523,N_3085,N_3229);
or U3524 (N_3524,N_3371,N_3005);
and U3525 (N_3525,N_3405,N_3132);
nor U3526 (N_3526,N_3122,N_3441);
nor U3527 (N_3527,N_3406,N_3101);
nor U3528 (N_3528,N_3420,N_3382);
xor U3529 (N_3529,N_3311,N_3075);
and U3530 (N_3530,N_3432,N_3003);
and U3531 (N_3531,N_3125,N_3040);
and U3532 (N_3532,N_3196,N_3020);
and U3533 (N_3533,N_3480,N_3447);
and U3534 (N_3534,N_3174,N_3061);
xor U3535 (N_3535,N_3419,N_3378);
and U3536 (N_3536,N_3198,N_3129);
nand U3537 (N_3537,N_3140,N_3221);
or U3538 (N_3538,N_3004,N_3135);
nor U3539 (N_3539,N_3352,N_3182);
xor U3540 (N_3540,N_3440,N_3156);
or U3541 (N_3541,N_3346,N_3326);
nor U3542 (N_3542,N_3026,N_3164);
and U3543 (N_3543,N_3218,N_3099);
and U3544 (N_3544,N_3019,N_3178);
nand U3545 (N_3545,N_3289,N_3018);
and U3546 (N_3546,N_3124,N_3037);
nor U3547 (N_3547,N_3095,N_3208);
and U3548 (N_3548,N_3136,N_3308);
and U3549 (N_3549,N_3171,N_3054);
nor U3550 (N_3550,N_3365,N_3192);
nor U3551 (N_3551,N_3284,N_3241);
nor U3552 (N_3552,N_3413,N_3399);
nand U3553 (N_3553,N_3264,N_3223);
nor U3554 (N_3554,N_3276,N_3321);
nor U3555 (N_3555,N_3200,N_3065);
and U3556 (N_3556,N_3362,N_3476);
nor U3557 (N_3557,N_3083,N_3231);
and U3558 (N_3558,N_3274,N_3069);
or U3559 (N_3559,N_3186,N_3194);
nor U3560 (N_3560,N_3146,N_3070);
nand U3561 (N_3561,N_3010,N_3390);
nor U3562 (N_3562,N_3409,N_3103);
and U3563 (N_3563,N_3047,N_3486);
or U3564 (N_3564,N_3373,N_3392);
nand U3565 (N_3565,N_3408,N_3366);
or U3566 (N_3566,N_3437,N_3257);
nor U3567 (N_3567,N_3115,N_3395);
and U3568 (N_3568,N_3479,N_3023);
nand U3569 (N_3569,N_3433,N_3312);
and U3570 (N_3570,N_3079,N_3495);
nand U3571 (N_3571,N_3252,N_3240);
or U3572 (N_3572,N_3314,N_3220);
or U3573 (N_3573,N_3270,N_3379);
nand U3574 (N_3574,N_3062,N_3268);
and U3575 (N_3575,N_3067,N_3217);
and U3576 (N_3576,N_3185,N_3012);
nor U3577 (N_3577,N_3391,N_3426);
and U3578 (N_3578,N_3456,N_3162);
nor U3579 (N_3579,N_3402,N_3335);
nor U3580 (N_3580,N_3416,N_3230);
nand U3581 (N_3581,N_3499,N_3009);
nand U3582 (N_3582,N_3282,N_3277);
and U3583 (N_3583,N_3007,N_3283);
and U3584 (N_3584,N_3034,N_3417);
or U3585 (N_3585,N_3137,N_3280);
or U3586 (N_3586,N_3363,N_3255);
nand U3587 (N_3587,N_3128,N_3024);
nor U3588 (N_3588,N_3300,N_3149);
nor U3589 (N_3589,N_3262,N_3370);
nand U3590 (N_3590,N_3322,N_3036);
nand U3591 (N_3591,N_3439,N_3380);
and U3592 (N_3592,N_3097,N_3496);
or U3593 (N_3593,N_3251,N_3106);
and U3594 (N_3594,N_3291,N_3294);
and U3595 (N_3595,N_3474,N_3466);
or U3596 (N_3596,N_3250,N_3123);
or U3597 (N_3597,N_3292,N_3160);
nand U3598 (N_3598,N_3337,N_3396);
xor U3599 (N_3599,N_3243,N_3151);
and U3600 (N_3600,N_3144,N_3376);
or U3601 (N_3601,N_3472,N_3205);
nand U3602 (N_3602,N_3461,N_3317);
nand U3603 (N_3603,N_3060,N_3081);
or U3604 (N_3604,N_3059,N_3064);
nand U3605 (N_3605,N_3150,N_3385);
or U3606 (N_3606,N_3297,N_3030);
nand U3607 (N_3607,N_3339,N_3448);
nor U3608 (N_3608,N_3089,N_3253);
xnor U3609 (N_3609,N_3025,N_3279);
and U3610 (N_3610,N_3348,N_3236);
nand U3611 (N_3611,N_3126,N_3457);
and U3612 (N_3612,N_3313,N_3116);
nand U3613 (N_3613,N_3265,N_3038);
or U3614 (N_3614,N_3434,N_3428);
or U3615 (N_3615,N_3449,N_3367);
and U3616 (N_3616,N_3302,N_3206);
and U3617 (N_3617,N_3298,N_3438);
nand U3618 (N_3618,N_3074,N_3090);
xor U3619 (N_3619,N_3247,N_3491);
or U3620 (N_3620,N_3006,N_3254);
or U3621 (N_3621,N_3455,N_3133);
and U3622 (N_3622,N_3189,N_3343);
nor U3623 (N_3623,N_3035,N_3167);
nand U3624 (N_3624,N_3482,N_3102);
and U3625 (N_3625,N_3077,N_3497);
or U3626 (N_3626,N_3351,N_3349);
xor U3627 (N_3627,N_3080,N_3166);
and U3628 (N_3628,N_3469,N_3092);
nor U3629 (N_3629,N_3042,N_3244);
nor U3630 (N_3630,N_3301,N_3261);
nand U3631 (N_3631,N_3100,N_3068);
or U3632 (N_3632,N_3215,N_3287);
and U3633 (N_3633,N_3163,N_3316);
and U3634 (N_3634,N_3481,N_3204);
and U3635 (N_3635,N_3238,N_3487);
nor U3636 (N_3636,N_3141,N_3177);
and U3637 (N_3637,N_3052,N_3285);
nand U3638 (N_3638,N_3278,N_3152);
nand U3639 (N_3639,N_3330,N_3105);
nand U3640 (N_3640,N_3465,N_3422);
nand U3641 (N_3641,N_3161,N_3299);
or U3642 (N_3642,N_3353,N_3239);
nor U3643 (N_3643,N_3451,N_3397);
nor U3644 (N_3644,N_3181,N_3410);
or U3645 (N_3645,N_3094,N_3072);
or U3646 (N_3646,N_3490,N_3131);
and U3647 (N_3647,N_3415,N_3310);
or U3648 (N_3648,N_3435,N_3494);
or U3649 (N_3649,N_3147,N_3000);
nor U3650 (N_3650,N_3355,N_3369);
xnor U3651 (N_3651,N_3237,N_3224);
and U3652 (N_3652,N_3319,N_3443);
and U3653 (N_3653,N_3445,N_3411);
nand U3654 (N_3654,N_3228,N_3058);
nand U3655 (N_3655,N_3442,N_3400);
xor U3656 (N_3656,N_3488,N_3273);
and U3657 (N_3657,N_3331,N_3120);
nand U3658 (N_3658,N_3112,N_3338);
nor U3659 (N_3659,N_3127,N_3249);
nand U3660 (N_3660,N_3305,N_3306);
and U3661 (N_3661,N_3336,N_3117);
or U3662 (N_3662,N_3444,N_3329);
nor U3663 (N_3663,N_3429,N_3484);
nand U3664 (N_3664,N_3214,N_3130);
or U3665 (N_3665,N_3328,N_3078);
or U3666 (N_3666,N_3372,N_3304);
xnor U3667 (N_3667,N_3360,N_3387);
nor U3668 (N_3668,N_3158,N_3248);
or U3669 (N_3669,N_3191,N_3464);
or U3670 (N_3670,N_3423,N_3197);
nor U3671 (N_3671,N_3057,N_3179);
or U3672 (N_3672,N_3468,N_3119);
nand U3673 (N_3673,N_3404,N_3193);
nand U3674 (N_3674,N_3286,N_3475);
nand U3675 (N_3675,N_3108,N_3345);
xnor U3676 (N_3676,N_3212,N_3073);
xnor U3677 (N_3677,N_3086,N_3356);
nor U3678 (N_3678,N_3333,N_3104);
or U3679 (N_3679,N_3183,N_3096);
nand U3680 (N_3680,N_3266,N_3354);
nor U3681 (N_3681,N_3015,N_3008);
and U3682 (N_3682,N_3232,N_3180);
and U3683 (N_3683,N_3493,N_3165);
nand U3684 (N_3684,N_3170,N_3296);
or U3685 (N_3685,N_3066,N_3142);
nor U3686 (N_3686,N_3098,N_3383);
or U3687 (N_3687,N_3473,N_3210);
and U3688 (N_3688,N_3148,N_3401);
and U3689 (N_3689,N_3460,N_3281);
nand U3690 (N_3690,N_3216,N_3207);
nand U3691 (N_3691,N_3453,N_3199);
xor U3692 (N_3692,N_3110,N_3318);
xor U3693 (N_3693,N_3394,N_3087);
and U3694 (N_3694,N_3388,N_3386);
or U3695 (N_3695,N_3269,N_3046);
nand U3696 (N_3696,N_3145,N_3498);
and U3697 (N_3697,N_3211,N_3446);
and U3698 (N_3698,N_3016,N_3246);
nor U3699 (N_3699,N_3344,N_3393);
and U3700 (N_3700,N_3462,N_3226);
or U3701 (N_3701,N_3121,N_3027);
nor U3702 (N_3702,N_3368,N_3045);
nor U3703 (N_3703,N_3327,N_3459);
and U3704 (N_3704,N_3048,N_3458);
nand U3705 (N_3705,N_3414,N_3307);
nor U3706 (N_3706,N_3303,N_3471);
nand U3707 (N_3707,N_3403,N_3470);
nor U3708 (N_3708,N_3169,N_3091);
and U3709 (N_3709,N_3031,N_3190);
nand U3710 (N_3710,N_3051,N_3175);
nand U3711 (N_3711,N_3334,N_3028);
xor U3712 (N_3712,N_3381,N_3222);
xnor U3713 (N_3713,N_3093,N_3113);
or U3714 (N_3714,N_3056,N_3454);
or U3715 (N_3715,N_3412,N_3452);
or U3716 (N_3716,N_3138,N_3213);
or U3717 (N_3717,N_3267,N_3358);
nand U3718 (N_3718,N_3203,N_3014);
nand U3719 (N_3719,N_3477,N_3431);
nand U3720 (N_3720,N_3256,N_3143);
nand U3721 (N_3721,N_3424,N_3017);
nand U3722 (N_3722,N_3483,N_3050);
nor U3723 (N_3723,N_3139,N_3342);
nor U3724 (N_3724,N_3258,N_3340);
or U3725 (N_3725,N_3029,N_3359);
or U3726 (N_3726,N_3043,N_3463);
and U3727 (N_3727,N_3153,N_3275);
and U3728 (N_3728,N_3134,N_3002);
nor U3729 (N_3729,N_3159,N_3293);
or U3730 (N_3730,N_3227,N_3245);
nor U3731 (N_3731,N_3364,N_3332);
and U3732 (N_3732,N_3233,N_3063);
or U3733 (N_3733,N_3350,N_3235);
xor U3734 (N_3734,N_3323,N_3389);
nand U3735 (N_3735,N_3375,N_3082);
nand U3736 (N_3736,N_3173,N_3325);
nor U3737 (N_3737,N_3033,N_3377);
xor U3738 (N_3738,N_3202,N_3492);
nand U3739 (N_3739,N_3436,N_3184);
nor U3740 (N_3740,N_3111,N_3450);
and U3741 (N_3741,N_3114,N_3039);
nor U3742 (N_3742,N_3053,N_3107);
nand U3743 (N_3743,N_3209,N_3234);
nand U3744 (N_3744,N_3384,N_3044);
nor U3745 (N_3745,N_3288,N_3049);
or U3746 (N_3746,N_3071,N_3201);
nor U3747 (N_3747,N_3272,N_3430);
or U3748 (N_3748,N_3374,N_3347);
nor U3749 (N_3749,N_3290,N_3315);
nand U3750 (N_3750,N_3404,N_3367);
and U3751 (N_3751,N_3407,N_3318);
nor U3752 (N_3752,N_3295,N_3124);
and U3753 (N_3753,N_3107,N_3198);
xnor U3754 (N_3754,N_3435,N_3466);
and U3755 (N_3755,N_3145,N_3179);
nor U3756 (N_3756,N_3452,N_3446);
nor U3757 (N_3757,N_3402,N_3113);
or U3758 (N_3758,N_3147,N_3494);
and U3759 (N_3759,N_3298,N_3181);
nand U3760 (N_3760,N_3239,N_3204);
nand U3761 (N_3761,N_3213,N_3141);
nand U3762 (N_3762,N_3391,N_3077);
nor U3763 (N_3763,N_3123,N_3148);
and U3764 (N_3764,N_3298,N_3092);
nand U3765 (N_3765,N_3018,N_3487);
and U3766 (N_3766,N_3386,N_3053);
nand U3767 (N_3767,N_3000,N_3093);
or U3768 (N_3768,N_3101,N_3256);
nor U3769 (N_3769,N_3090,N_3394);
or U3770 (N_3770,N_3020,N_3155);
nor U3771 (N_3771,N_3203,N_3321);
nand U3772 (N_3772,N_3017,N_3077);
xnor U3773 (N_3773,N_3041,N_3284);
nand U3774 (N_3774,N_3004,N_3353);
nand U3775 (N_3775,N_3256,N_3222);
nor U3776 (N_3776,N_3102,N_3157);
and U3777 (N_3777,N_3468,N_3428);
nand U3778 (N_3778,N_3248,N_3082);
and U3779 (N_3779,N_3196,N_3467);
and U3780 (N_3780,N_3425,N_3343);
xnor U3781 (N_3781,N_3271,N_3397);
nor U3782 (N_3782,N_3068,N_3052);
nor U3783 (N_3783,N_3300,N_3269);
and U3784 (N_3784,N_3189,N_3243);
and U3785 (N_3785,N_3327,N_3051);
nor U3786 (N_3786,N_3033,N_3486);
nand U3787 (N_3787,N_3491,N_3443);
and U3788 (N_3788,N_3150,N_3302);
and U3789 (N_3789,N_3497,N_3255);
nand U3790 (N_3790,N_3035,N_3074);
or U3791 (N_3791,N_3497,N_3051);
nor U3792 (N_3792,N_3241,N_3183);
nand U3793 (N_3793,N_3113,N_3421);
and U3794 (N_3794,N_3371,N_3466);
nor U3795 (N_3795,N_3482,N_3245);
xnor U3796 (N_3796,N_3361,N_3066);
nand U3797 (N_3797,N_3010,N_3029);
xnor U3798 (N_3798,N_3483,N_3279);
nor U3799 (N_3799,N_3282,N_3442);
or U3800 (N_3800,N_3320,N_3134);
and U3801 (N_3801,N_3167,N_3306);
and U3802 (N_3802,N_3395,N_3361);
and U3803 (N_3803,N_3225,N_3442);
nand U3804 (N_3804,N_3006,N_3002);
or U3805 (N_3805,N_3360,N_3165);
or U3806 (N_3806,N_3257,N_3397);
and U3807 (N_3807,N_3434,N_3117);
nor U3808 (N_3808,N_3188,N_3257);
or U3809 (N_3809,N_3196,N_3354);
or U3810 (N_3810,N_3229,N_3244);
xnor U3811 (N_3811,N_3359,N_3215);
xnor U3812 (N_3812,N_3168,N_3154);
and U3813 (N_3813,N_3375,N_3423);
or U3814 (N_3814,N_3486,N_3198);
nor U3815 (N_3815,N_3358,N_3231);
xnor U3816 (N_3816,N_3378,N_3457);
xnor U3817 (N_3817,N_3449,N_3191);
nand U3818 (N_3818,N_3349,N_3348);
and U3819 (N_3819,N_3139,N_3059);
xnor U3820 (N_3820,N_3061,N_3025);
xor U3821 (N_3821,N_3126,N_3345);
or U3822 (N_3822,N_3466,N_3232);
nand U3823 (N_3823,N_3464,N_3019);
or U3824 (N_3824,N_3164,N_3341);
or U3825 (N_3825,N_3185,N_3127);
nor U3826 (N_3826,N_3093,N_3265);
and U3827 (N_3827,N_3164,N_3023);
and U3828 (N_3828,N_3322,N_3181);
or U3829 (N_3829,N_3029,N_3154);
and U3830 (N_3830,N_3090,N_3424);
or U3831 (N_3831,N_3064,N_3343);
or U3832 (N_3832,N_3115,N_3246);
nor U3833 (N_3833,N_3149,N_3241);
and U3834 (N_3834,N_3296,N_3370);
nor U3835 (N_3835,N_3364,N_3211);
and U3836 (N_3836,N_3224,N_3101);
nor U3837 (N_3837,N_3494,N_3189);
or U3838 (N_3838,N_3295,N_3380);
nand U3839 (N_3839,N_3307,N_3254);
nor U3840 (N_3840,N_3341,N_3124);
xor U3841 (N_3841,N_3463,N_3309);
nand U3842 (N_3842,N_3474,N_3256);
and U3843 (N_3843,N_3166,N_3152);
nor U3844 (N_3844,N_3109,N_3413);
nand U3845 (N_3845,N_3034,N_3281);
nor U3846 (N_3846,N_3116,N_3094);
nand U3847 (N_3847,N_3308,N_3351);
nor U3848 (N_3848,N_3059,N_3346);
xor U3849 (N_3849,N_3363,N_3127);
nand U3850 (N_3850,N_3450,N_3373);
xnor U3851 (N_3851,N_3449,N_3093);
and U3852 (N_3852,N_3392,N_3469);
xor U3853 (N_3853,N_3174,N_3248);
nand U3854 (N_3854,N_3327,N_3432);
nor U3855 (N_3855,N_3422,N_3316);
and U3856 (N_3856,N_3497,N_3135);
nand U3857 (N_3857,N_3183,N_3480);
or U3858 (N_3858,N_3190,N_3421);
and U3859 (N_3859,N_3187,N_3308);
or U3860 (N_3860,N_3254,N_3269);
and U3861 (N_3861,N_3311,N_3456);
or U3862 (N_3862,N_3089,N_3036);
or U3863 (N_3863,N_3233,N_3246);
or U3864 (N_3864,N_3490,N_3314);
and U3865 (N_3865,N_3407,N_3044);
nand U3866 (N_3866,N_3470,N_3201);
nand U3867 (N_3867,N_3017,N_3049);
nand U3868 (N_3868,N_3238,N_3249);
or U3869 (N_3869,N_3442,N_3160);
nor U3870 (N_3870,N_3245,N_3063);
and U3871 (N_3871,N_3462,N_3386);
and U3872 (N_3872,N_3388,N_3216);
nor U3873 (N_3873,N_3264,N_3153);
and U3874 (N_3874,N_3094,N_3092);
nor U3875 (N_3875,N_3386,N_3008);
nor U3876 (N_3876,N_3176,N_3022);
and U3877 (N_3877,N_3247,N_3297);
and U3878 (N_3878,N_3282,N_3415);
nand U3879 (N_3879,N_3087,N_3363);
nor U3880 (N_3880,N_3312,N_3290);
or U3881 (N_3881,N_3071,N_3123);
nand U3882 (N_3882,N_3429,N_3104);
nor U3883 (N_3883,N_3002,N_3126);
or U3884 (N_3884,N_3375,N_3204);
and U3885 (N_3885,N_3333,N_3161);
and U3886 (N_3886,N_3001,N_3091);
nor U3887 (N_3887,N_3125,N_3066);
xor U3888 (N_3888,N_3304,N_3332);
nand U3889 (N_3889,N_3188,N_3413);
or U3890 (N_3890,N_3145,N_3236);
and U3891 (N_3891,N_3394,N_3277);
nand U3892 (N_3892,N_3160,N_3208);
xnor U3893 (N_3893,N_3296,N_3302);
nor U3894 (N_3894,N_3348,N_3469);
and U3895 (N_3895,N_3455,N_3102);
and U3896 (N_3896,N_3413,N_3385);
or U3897 (N_3897,N_3057,N_3191);
or U3898 (N_3898,N_3186,N_3332);
nand U3899 (N_3899,N_3262,N_3254);
nor U3900 (N_3900,N_3474,N_3454);
or U3901 (N_3901,N_3290,N_3273);
nand U3902 (N_3902,N_3232,N_3205);
or U3903 (N_3903,N_3048,N_3289);
and U3904 (N_3904,N_3410,N_3351);
nand U3905 (N_3905,N_3157,N_3028);
nor U3906 (N_3906,N_3257,N_3212);
or U3907 (N_3907,N_3277,N_3461);
nor U3908 (N_3908,N_3201,N_3207);
nor U3909 (N_3909,N_3299,N_3074);
or U3910 (N_3910,N_3440,N_3001);
xor U3911 (N_3911,N_3465,N_3425);
or U3912 (N_3912,N_3008,N_3149);
and U3913 (N_3913,N_3223,N_3339);
or U3914 (N_3914,N_3232,N_3164);
nor U3915 (N_3915,N_3309,N_3453);
or U3916 (N_3916,N_3080,N_3465);
and U3917 (N_3917,N_3134,N_3060);
and U3918 (N_3918,N_3419,N_3259);
and U3919 (N_3919,N_3029,N_3367);
or U3920 (N_3920,N_3125,N_3417);
and U3921 (N_3921,N_3179,N_3014);
xor U3922 (N_3922,N_3009,N_3372);
nand U3923 (N_3923,N_3429,N_3279);
nor U3924 (N_3924,N_3273,N_3491);
or U3925 (N_3925,N_3056,N_3150);
and U3926 (N_3926,N_3444,N_3439);
nor U3927 (N_3927,N_3018,N_3127);
nand U3928 (N_3928,N_3333,N_3407);
or U3929 (N_3929,N_3306,N_3351);
nand U3930 (N_3930,N_3128,N_3131);
nor U3931 (N_3931,N_3357,N_3073);
and U3932 (N_3932,N_3034,N_3303);
or U3933 (N_3933,N_3404,N_3262);
and U3934 (N_3934,N_3308,N_3296);
nor U3935 (N_3935,N_3225,N_3246);
or U3936 (N_3936,N_3364,N_3282);
nand U3937 (N_3937,N_3417,N_3104);
and U3938 (N_3938,N_3477,N_3422);
and U3939 (N_3939,N_3346,N_3443);
and U3940 (N_3940,N_3183,N_3054);
and U3941 (N_3941,N_3095,N_3180);
or U3942 (N_3942,N_3357,N_3134);
nand U3943 (N_3943,N_3058,N_3284);
or U3944 (N_3944,N_3178,N_3400);
or U3945 (N_3945,N_3013,N_3245);
nand U3946 (N_3946,N_3123,N_3046);
or U3947 (N_3947,N_3397,N_3290);
or U3948 (N_3948,N_3132,N_3481);
nand U3949 (N_3949,N_3050,N_3113);
nand U3950 (N_3950,N_3220,N_3212);
nand U3951 (N_3951,N_3032,N_3477);
nand U3952 (N_3952,N_3236,N_3338);
and U3953 (N_3953,N_3288,N_3361);
or U3954 (N_3954,N_3017,N_3161);
nand U3955 (N_3955,N_3248,N_3218);
or U3956 (N_3956,N_3320,N_3186);
nand U3957 (N_3957,N_3458,N_3196);
nand U3958 (N_3958,N_3317,N_3375);
or U3959 (N_3959,N_3101,N_3336);
nand U3960 (N_3960,N_3319,N_3020);
nor U3961 (N_3961,N_3243,N_3074);
nor U3962 (N_3962,N_3224,N_3035);
or U3963 (N_3963,N_3492,N_3310);
nor U3964 (N_3964,N_3372,N_3116);
or U3965 (N_3965,N_3214,N_3149);
and U3966 (N_3966,N_3127,N_3414);
or U3967 (N_3967,N_3308,N_3243);
nand U3968 (N_3968,N_3241,N_3440);
or U3969 (N_3969,N_3376,N_3378);
and U3970 (N_3970,N_3026,N_3104);
xor U3971 (N_3971,N_3337,N_3206);
nand U3972 (N_3972,N_3376,N_3408);
or U3973 (N_3973,N_3064,N_3131);
and U3974 (N_3974,N_3278,N_3211);
nand U3975 (N_3975,N_3331,N_3130);
nand U3976 (N_3976,N_3198,N_3432);
nor U3977 (N_3977,N_3272,N_3047);
or U3978 (N_3978,N_3332,N_3166);
or U3979 (N_3979,N_3086,N_3447);
xor U3980 (N_3980,N_3260,N_3303);
nand U3981 (N_3981,N_3239,N_3207);
nor U3982 (N_3982,N_3408,N_3381);
and U3983 (N_3983,N_3345,N_3069);
and U3984 (N_3984,N_3289,N_3379);
and U3985 (N_3985,N_3370,N_3234);
and U3986 (N_3986,N_3446,N_3285);
nand U3987 (N_3987,N_3212,N_3296);
nand U3988 (N_3988,N_3322,N_3384);
nand U3989 (N_3989,N_3176,N_3118);
nor U3990 (N_3990,N_3330,N_3310);
nor U3991 (N_3991,N_3062,N_3421);
nand U3992 (N_3992,N_3055,N_3353);
xor U3993 (N_3993,N_3309,N_3336);
or U3994 (N_3994,N_3203,N_3355);
nor U3995 (N_3995,N_3441,N_3066);
and U3996 (N_3996,N_3163,N_3194);
or U3997 (N_3997,N_3283,N_3335);
nand U3998 (N_3998,N_3370,N_3497);
or U3999 (N_3999,N_3329,N_3041);
nor U4000 (N_4000,N_3569,N_3551);
and U4001 (N_4001,N_3736,N_3546);
nand U4002 (N_4002,N_3792,N_3828);
nor U4003 (N_4003,N_3872,N_3800);
or U4004 (N_4004,N_3525,N_3643);
nand U4005 (N_4005,N_3857,N_3819);
and U4006 (N_4006,N_3699,N_3501);
or U4007 (N_4007,N_3817,N_3747);
or U4008 (N_4008,N_3692,N_3612);
and U4009 (N_4009,N_3543,N_3632);
nand U4010 (N_4010,N_3676,N_3989);
nand U4011 (N_4011,N_3552,N_3767);
and U4012 (N_4012,N_3964,N_3658);
nor U4013 (N_4013,N_3944,N_3675);
nor U4014 (N_4014,N_3965,N_3926);
or U4015 (N_4015,N_3802,N_3861);
or U4016 (N_4016,N_3538,N_3743);
xnor U4017 (N_4017,N_3516,N_3687);
xnor U4018 (N_4018,N_3762,N_3704);
or U4019 (N_4019,N_3788,N_3834);
nor U4020 (N_4020,N_3639,N_3967);
and U4021 (N_4021,N_3672,N_3803);
nand U4022 (N_4022,N_3849,N_3642);
xor U4023 (N_4023,N_3850,N_3856);
nor U4024 (N_4024,N_3601,N_3727);
and U4025 (N_4025,N_3696,N_3522);
nor U4026 (N_4026,N_3689,N_3795);
xnor U4027 (N_4027,N_3983,N_3814);
nand U4028 (N_4028,N_3822,N_3905);
nand U4029 (N_4029,N_3674,N_3992);
nand U4030 (N_4030,N_3780,N_3877);
and U4031 (N_4031,N_3554,N_3997);
nand U4032 (N_4032,N_3726,N_3688);
or U4033 (N_4033,N_3793,N_3811);
and U4034 (N_4034,N_3994,N_3919);
and U4035 (N_4035,N_3592,N_3523);
and U4036 (N_4036,N_3591,N_3778);
and U4037 (N_4037,N_3644,N_3506);
nand U4038 (N_4038,N_3933,N_3535);
and U4039 (N_4039,N_3571,N_3627);
or U4040 (N_4040,N_3889,N_3904);
nor U4041 (N_4041,N_3786,N_3846);
nand U4042 (N_4042,N_3581,N_3930);
or U4043 (N_4043,N_3842,N_3827);
and U4044 (N_4044,N_3777,N_3716);
nor U4045 (N_4045,N_3695,N_3665);
and U4046 (N_4046,N_3691,N_3541);
or U4047 (N_4047,N_3991,N_3600);
and U4048 (N_4048,N_3745,N_3909);
xor U4049 (N_4049,N_3575,N_3621);
nand U4050 (N_4050,N_3536,N_3755);
and U4051 (N_4051,N_3680,N_3841);
xnor U4052 (N_4052,N_3902,N_3617);
nor U4053 (N_4053,N_3579,N_3661);
or U4054 (N_4054,N_3860,N_3911);
nor U4055 (N_4055,N_3609,N_3531);
or U4056 (N_4056,N_3830,N_3921);
and U4057 (N_4057,N_3999,N_3785);
nor U4058 (N_4058,N_3610,N_3720);
or U4059 (N_4059,N_3866,N_3836);
or U4060 (N_4060,N_3815,N_3844);
nand U4061 (N_4061,N_3570,N_3938);
and U4062 (N_4062,N_3995,N_3799);
and U4063 (N_4063,N_3611,N_3597);
nand U4064 (N_4064,N_3517,N_3824);
nor U4065 (N_4065,N_3553,N_3626);
nand U4066 (N_4066,N_3821,N_3813);
and U4067 (N_4067,N_3586,N_3532);
nor U4068 (N_4068,N_3787,N_3891);
and U4069 (N_4069,N_3895,N_3542);
or U4070 (N_4070,N_3721,N_3513);
nand U4071 (N_4071,N_3770,N_3763);
nor U4072 (N_4072,N_3764,N_3970);
and U4073 (N_4073,N_3556,N_3746);
or U4074 (N_4074,N_3550,N_3588);
nand U4075 (N_4075,N_3859,N_3594);
nand U4076 (N_4076,N_3577,N_3637);
and U4077 (N_4077,N_3843,N_3869);
or U4078 (N_4078,N_3740,N_3663);
nand U4079 (N_4079,N_3957,N_3707);
or U4080 (N_4080,N_3748,N_3684);
nand U4081 (N_4081,N_3858,N_3580);
and U4082 (N_4082,N_3718,N_3526);
nor U4083 (N_4083,N_3826,N_3972);
nor U4084 (N_4084,N_3664,N_3711);
nor U4085 (N_4085,N_3540,N_3947);
nor U4086 (N_4086,N_3982,N_3879);
or U4087 (N_4087,N_3629,N_3679);
or U4088 (N_4088,N_3912,N_3927);
and U4089 (N_4089,N_3710,N_3678);
and U4090 (N_4090,N_3503,N_3956);
nand U4091 (N_4091,N_3690,N_3880);
xor U4092 (N_4092,N_3724,N_3838);
or U4093 (N_4093,N_3804,N_3559);
nor U4094 (N_4094,N_3810,N_3515);
and U4095 (N_4095,N_3507,N_3761);
nand U4096 (N_4096,N_3700,N_3798);
nand U4097 (N_4097,N_3668,N_3511);
and U4098 (N_4098,N_3874,N_3568);
or U4099 (N_4099,N_3878,N_3618);
nor U4100 (N_4100,N_3654,N_3936);
xnor U4101 (N_4101,N_3774,N_3896);
xor U4102 (N_4102,N_3852,N_3922);
or U4103 (N_4103,N_3624,N_3607);
or U4104 (N_4104,N_3723,N_3741);
and U4105 (N_4105,N_3633,N_3809);
or U4106 (N_4106,N_3945,N_3766);
nand U4107 (N_4107,N_3835,N_3948);
nand U4108 (N_4108,N_3771,N_3587);
or U4109 (N_4109,N_3645,N_3693);
or U4110 (N_4110,N_3986,N_3660);
or U4111 (N_4111,N_3975,N_3980);
and U4112 (N_4112,N_3820,N_3722);
nor U4113 (N_4113,N_3705,N_3681);
nand U4114 (N_4114,N_3560,N_3833);
nand U4115 (N_4115,N_3653,N_3750);
or U4116 (N_4116,N_3988,N_3961);
nor U4117 (N_4117,N_3998,N_3518);
and U4118 (N_4118,N_3563,N_3537);
and U4119 (N_4119,N_3920,N_3502);
or U4120 (N_4120,N_3806,N_3595);
or U4121 (N_4121,N_3934,N_3655);
nor U4122 (N_4122,N_3840,N_3640);
and U4123 (N_4123,N_3558,N_3530);
and U4124 (N_4124,N_3873,N_3717);
nor U4125 (N_4125,N_3993,N_3925);
xor U4126 (N_4126,N_3625,N_3519);
nor U4127 (N_4127,N_3593,N_3818);
nand U4128 (N_4128,N_3590,N_3946);
and U4129 (N_4129,N_3702,N_3524);
and U4130 (N_4130,N_3776,N_3794);
or U4131 (N_4131,N_3968,N_3557);
or U4132 (N_4132,N_3917,N_3913);
and U4133 (N_4133,N_3529,N_3781);
or U4134 (N_4134,N_3737,N_3990);
and U4135 (N_4135,N_3508,N_3647);
xnor U4136 (N_4136,N_3953,N_3935);
nand U4137 (N_4137,N_3966,N_3751);
or U4138 (N_4138,N_3505,N_3574);
xnor U4139 (N_4139,N_3694,N_3918);
and U4140 (N_4140,N_3978,N_3728);
or U4141 (N_4141,N_3547,N_3709);
or U4142 (N_4142,N_3949,N_3862);
and U4143 (N_4143,N_3888,N_3883);
nor U4144 (N_4144,N_3744,N_3671);
nor U4145 (N_4145,N_3915,N_3662);
or U4146 (N_4146,N_3969,N_3510);
or U4147 (N_4147,N_3871,N_3686);
or U4148 (N_4148,N_3756,N_3562);
nor U4149 (N_4149,N_3730,N_3659);
xnor U4150 (N_4150,N_3753,N_3708);
and U4151 (N_4151,N_3954,N_3848);
nand U4152 (N_4152,N_3782,N_3649);
nor U4153 (N_4153,N_3719,N_3779);
and U4154 (N_4154,N_3976,N_3566);
nand U4155 (N_4155,N_3528,N_3853);
nand U4156 (N_4156,N_3725,N_3955);
nor U4157 (N_4157,N_3555,N_3548);
nand U4158 (N_4158,N_3876,N_3527);
or U4159 (N_4159,N_3772,N_3900);
or U4160 (N_4160,N_3666,N_3608);
or U4161 (N_4161,N_3646,N_3765);
nand U4162 (N_4162,N_3789,N_3942);
and U4163 (N_4163,N_3635,N_3735);
nor U4164 (N_4164,N_3619,N_3749);
and U4165 (N_4165,N_3738,N_3952);
and U4166 (N_4166,N_3573,N_3974);
and U4167 (N_4167,N_3549,N_3829);
nor U4168 (N_4168,N_3739,N_3882);
nand U4169 (N_4169,N_3604,N_3576);
and U4170 (N_4170,N_3996,N_3791);
and U4171 (N_4171,N_3931,N_3760);
xor U4172 (N_4172,N_3713,N_3939);
nand U4173 (N_4173,N_3729,N_3596);
nor U4174 (N_4174,N_3636,N_3582);
and U4175 (N_4175,N_3937,N_3837);
xor U4176 (N_4176,N_3768,N_3775);
nor U4177 (N_4177,N_3928,N_3685);
nand U4178 (N_4178,N_3545,N_3868);
nand U4179 (N_4179,N_3533,N_3539);
and U4180 (N_4180,N_3839,N_3697);
and U4181 (N_4181,N_3698,N_3941);
nand U4182 (N_4182,N_3914,N_3520);
nor U4183 (N_4183,N_3544,N_3894);
and U4184 (N_4184,N_3924,N_3583);
xnor U4185 (N_4185,N_3808,N_3784);
nand U4186 (N_4186,N_3863,N_3758);
nand U4187 (N_4187,N_3567,N_3881);
nor U4188 (N_4188,N_3669,N_3951);
nand U4189 (N_4189,N_3959,N_3855);
xnor U4190 (N_4190,N_3509,N_3977);
nand U4191 (N_4191,N_3682,N_3892);
xor U4192 (N_4192,N_3812,N_3534);
nand U4193 (N_4193,N_3500,N_3677);
and U4194 (N_4194,N_3932,N_3845);
and U4195 (N_4195,N_3823,N_3910);
nand U4196 (N_4196,N_3971,N_3870);
or U4197 (N_4197,N_3564,N_3790);
and U4198 (N_4198,N_3731,N_3732);
nand U4199 (N_4199,N_3923,N_3641);
nand U4200 (N_4200,N_3578,N_3648);
nand U4201 (N_4201,N_3963,N_3630);
nand U4202 (N_4202,N_3851,N_3907);
or U4203 (N_4203,N_3890,N_3985);
or U4204 (N_4204,N_3854,N_3634);
xnor U4205 (N_4205,N_3512,N_3701);
or U4206 (N_4206,N_3757,N_3514);
and U4207 (N_4207,N_3614,N_3801);
nor U4208 (N_4208,N_3950,N_3703);
xnor U4209 (N_4209,N_3589,N_3783);
nand U4210 (N_4210,N_3733,N_3906);
nand U4211 (N_4211,N_3638,N_3897);
or U4212 (N_4212,N_3885,N_3831);
xnor U4213 (N_4213,N_3807,N_3667);
or U4214 (N_4214,N_3984,N_3584);
nor U4215 (N_4215,N_3832,N_3613);
nor U4216 (N_4216,N_3901,N_3712);
or U4217 (N_4217,N_3887,N_3973);
nor U4218 (N_4218,N_3816,N_3865);
nor U4219 (N_4219,N_3884,N_3673);
nand U4220 (N_4220,N_3615,N_3960);
or U4221 (N_4221,N_3504,N_3652);
and U4222 (N_4222,N_3734,N_3521);
nand U4223 (N_4223,N_3979,N_3620);
nor U4224 (N_4224,N_3797,N_3623);
xnor U4225 (N_4225,N_3606,N_3940);
nand U4226 (N_4226,N_3670,N_3714);
xor U4227 (N_4227,N_3598,N_3706);
or U4228 (N_4228,N_3886,N_3864);
nor U4229 (N_4229,N_3759,N_3769);
or U4230 (N_4230,N_3603,N_3752);
nor U4231 (N_4231,N_3916,N_3943);
or U4232 (N_4232,N_3657,N_3867);
nand U4233 (N_4233,N_3898,N_3616);
nand U4234 (N_4234,N_3987,N_3599);
nand U4235 (N_4235,N_3715,N_3622);
or U4236 (N_4236,N_3754,N_3605);
nor U4237 (N_4237,N_3893,N_3908);
xnor U4238 (N_4238,N_3875,N_3561);
or U4239 (N_4239,N_3929,N_3572);
or U4240 (N_4240,N_3962,N_3585);
or U4241 (N_4241,N_3742,N_3656);
and U4242 (N_4242,N_3825,N_3650);
or U4243 (N_4243,N_3651,N_3628);
nand U4244 (N_4244,N_3796,N_3683);
nand U4245 (N_4245,N_3602,N_3631);
nand U4246 (N_4246,N_3903,N_3981);
and U4247 (N_4247,N_3899,N_3847);
nand U4248 (N_4248,N_3805,N_3958);
xor U4249 (N_4249,N_3565,N_3773);
nor U4250 (N_4250,N_3977,N_3610);
nor U4251 (N_4251,N_3570,N_3555);
or U4252 (N_4252,N_3994,N_3728);
nand U4253 (N_4253,N_3503,N_3738);
nor U4254 (N_4254,N_3531,N_3767);
nand U4255 (N_4255,N_3516,N_3576);
xor U4256 (N_4256,N_3718,N_3784);
or U4257 (N_4257,N_3693,N_3994);
xnor U4258 (N_4258,N_3931,N_3503);
or U4259 (N_4259,N_3609,N_3995);
and U4260 (N_4260,N_3574,N_3710);
or U4261 (N_4261,N_3941,N_3589);
nor U4262 (N_4262,N_3576,N_3682);
nor U4263 (N_4263,N_3902,N_3896);
nor U4264 (N_4264,N_3623,N_3851);
or U4265 (N_4265,N_3780,N_3901);
nor U4266 (N_4266,N_3745,N_3616);
or U4267 (N_4267,N_3770,N_3959);
or U4268 (N_4268,N_3886,N_3690);
xor U4269 (N_4269,N_3623,N_3624);
nand U4270 (N_4270,N_3745,N_3885);
or U4271 (N_4271,N_3832,N_3678);
nand U4272 (N_4272,N_3924,N_3935);
nor U4273 (N_4273,N_3524,N_3882);
and U4274 (N_4274,N_3900,N_3997);
and U4275 (N_4275,N_3521,N_3841);
or U4276 (N_4276,N_3644,N_3724);
nor U4277 (N_4277,N_3895,N_3861);
nand U4278 (N_4278,N_3556,N_3876);
or U4279 (N_4279,N_3540,N_3627);
xnor U4280 (N_4280,N_3860,N_3975);
or U4281 (N_4281,N_3656,N_3838);
and U4282 (N_4282,N_3953,N_3565);
or U4283 (N_4283,N_3983,N_3530);
nor U4284 (N_4284,N_3727,N_3909);
or U4285 (N_4285,N_3994,N_3569);
nor U4286 (N_4286,N_3853,N_3907);
nor U4287 (N_4287,N_3517,N_3815);
nand U4288 (N_4288,N_3887,N_3623);
nand U4289 (N_4289,N_3937,N_3827);
and U4290 (N_4290,N_3585,N_3621);
nor U4291 (N_4291,N_3833,N_3543);
nor U4292 (N_4292,N_3784,N_3774);
or U4293 (N_4293,N_3583,N_3903);
or U4294 (N_4294,N_3561,N_3719);
nor U4295 (N_4295,N_3914,N_3515);
nor U4296 (N_4296,N_3934,N_3712);
and U4297 (N_4297,N_3857,N_3748);
nand U4298 (N_4298,N_3795,N_3503);
and U4299 (N_4299,N_3793,N_3576);
and U4300 (N_4300,N_3679,N_3714);
or U4301 (N_4301,N_3992,N_3934);
or U4302 (N_4302,N_3579,N_3785);
and U4303 (N_4303,N_3561,N_3979);
nor U4304 (N_4304,N_3627,N_3546);
or U4305 (N_4305,N_3712,N_3897);
nand U4306 (N_4306,N_3839,N_3595);
or U4307 (N_4307,N_3638,N_3566);
or U4308 (N_4308,N_3751,N_3635);
or U4309 (N_4309,N_3883,N_3718);
nand U4310 (N_4310,N_3869,N_3723);
nand U4311 (N_4311,N_3836,N_3541);
and U4312 (N_4312,N_3850,N_3890);
and U4313 (N_4313,N_3623,N_3998);
nor U4314 (N_4314,N_3773,N_3746);
or U4315 (N_4315,N_3890,N_3829);
nor U4316 (N_4316,N_3730,N_3687);
nand U4317 (N_4317,N_3846,N_3947);
or U4318 (N_4318,N_3587,N_3744);
nor U4319 (N_4319,N_3683,N_3765);
and U4320 (N_4320,N_3857,N_3648);
and U4321 (N_4321,N_3978,N_3504);
nand U4322 (N_4322,N_3948,N_3714);
nor U4323 (N_4323,N_3866,N_3709);
nor U4324 (N_4324,N_3789,N_3720);
and U4325 (N_4325,N_3621,N_3750);
and U4326 (N_4326,N_3831,N_3783);
and U4327 (N_4327,N_3848,N_3731);
xor U4328 (N_4328,N_3871,N_3531);
and U4329 (N_4329,N_3871,N_3500);
or U4330 (N_4330,N_3997,N_3775);
or U4331 (N_4331,N_3575,N_3750);
nor U4332 (N_4332,N_3627,N_3962);
and U4333 (N_4333,N_3504,N_3900);
or U4334 (N_4334,N_3735,N_3959);
nand U4335 (N_4335,N_3826,N_3675);
and U4336 (N_4336,N_3701,N_3721);
and U4337 (N_4337,N_3814,N_3576);
nand U4338 (N_4338,N_3841,N_3588);
and U4339 (N_4339,N_3827,N_3948);
or U4340 (N_4340,N_3803,N_3914);
and U4341 (N_4341,N_3538,N_3981);
nand U4342 (N_4342,N_3994,N_3663);
and U4343 (N_4343,N_3933,N_3691);
nor U4344 (N_4344,N_3685,N_3740);
or U4345 (N_4345,N_3778,N_3763);
nand U4346 (N_4346,N_3857,N_3743);
nor U4347 (N_4347,N_3556,N_3608);
nand U4348 (N_4348,N_3949,N_3959);
xor U4349 (N_4349,N_3759,N_3878);
xor U4350 (N_4350,N_3987,N_3897);
or U4351 (N_4351,N_3667,N_3877);
and U4352 (N_4352,N_3990,N_3779);
nand U4353 (N_4353,N_3703,N_3817);
or U4354 (N_4354,N_3562,N_3525);
nor U4355 (N_4355,N_3619,N_3513);
nand U4356 (N_4356,N_3585,N_3527);
nand U4357 (N_4357,N_3715,N_3693);
nand U4358 (N_4358,N_3749,N_3937);
nor U4359 (N_4359,N_3658,N_3703);
nand U4360 (N_4360,N_3635,N_3815);
nand U4361 (N_4361,N_3550,N_3944);
or U4362 (N_4362,N_3951,N_3610);
nand U4363 (N_4363,N_3980,N_3696);
and U4364 (N_4364,N_3681,N_3628);
and U4365 (N_4365,N_3589,N_3983);
nand U4366 (N_4366,N_3838,N_3702);
xor U4367 (N_4367,N_3563,N_3529);
and U4368 (N_4368,N_3692,N_3673);
xnor U4369 (N_4369,N_3932,N_3806);
nor U4370 (N_4370,N_3590,N_3997);
nor U4371 (N_4371,N_3700,N_3626);
or U4372 (N_4372,N_3532,N_3681);
nand U4373 (N_4373,N_3753,N_3523);
nand U4374 (N_4374,N_3675,N_3520);
nor U4375 (N_4375,N_3827,N_3815);
nand U4376 (N_4376,N_3666,N_3691);
or U4377 (N_4377,N_3852,N_3860);
nor U4378 (N_4378,N_3837,N_3625);
and U4379 (N_4379,N_3797,N_3686);
nor U4380 (N_4380,N_3875,N_3978);
xnor U4381 (N_4381,N_3848,N_3953);
or U4382 (N_4382,N_3512,N_3749);
and U4383 (N_4383,N_3723,N_3899);
and U4384 (N_4384,N_3900,N_3985);
and U4385 (N_4385,N_3531,N_3639);
or U4386 (N_4386,N_3783,N_3600);
nor U4387 (N_4387,N_3601,N_3950);
nor U4388 (N_4388,N_3803,N_3810);
nand U4389 (N_4389,N_3549,N_3840);
or U4390 (N_4390,N_3829,N_3790);
or U4391 (N_4391,N_3857,N_3593);
or U4392 (N_4392,N_3692,N_3636);
nand U4393 (N_4393,N_3500,N_3616);
nand U4394 (N_4394,N_3922,N_3644);
or U4395 (N_4395,N_3851,N_3642);
or U4396 (N_4396,N_3689,N_3552);
or U4397 (N_4397,N_3704,N_3930);
nand U4398 (N_4398,N_3701,N_3801);
nor U4399 (N_4399,N_3862,N_3909);
nor U4400 (N_4400,N_3682,N_3865);
nand U4401 (N_4401,N_3676,N_3551);
nand U4402 (N_4402,N_3533,N_3653);
nand U4403 (N_4403,N_3758,N_3848);
and U4404 (N_4404,N_3955,N_3829);
or U4405 (N_4405,N_3977,N_3789);
or U4406 (N_4406,N_3813,N_3886);
nor U4407 (N_4407,N_3886,N_3507);
and U4408 (N_4408,N_3949,N_3936);
or U4409 (N_4409,N_3771,N_3584);
nand U4410 (N_4410,N_3964,N_3740);
nand U4411 (N_4411,N_3956,N_3964);
or U4412 (N_4412,N_3968,N_3706);
and U4413 (N_4413,N_3905,N_3834);
and U4414 (N_4414,N_3811,N_3540);
and U4415 (N_4415,N_3905,N_3807);
and U4416 (N_4416,N_3923,N_3971);
and U4417 (N_4417,N_3531,N_3593);
xnor U4418 (N_4418,N_3505,N_3565);
nand U4419 (N_4419,N_3845,N_3962);
or U4420 (N_4420,N_3595,N_3845);
nor U4421 (N_4421,N_3874,N_3857);
xor U4422 (N_4422,N_3706,N_3956);
nor U4423 (N_4423,N_3762,N_3881);
or U4424 (N_4424,N_3728,N_3642);
nand U4425 (N_4425,N_3737,N_3954);
and U4426 (N_4426,N_3613,N_3638);
nor U4427 (N_4427,N_3719,N_3786);
and U4428 (N_4428,N_3559,N_3536);
xnor U4429 (N_4429,N_3544,N_3608);
nor U4430 (N_4430,N_3575,N_3891);
and U4431 (N_4431,N_3687,N_3549);
and U4432 (N_4432,N_3720,N_3985);
nor U4433 (N_4433,N_3991,N_3839);
nand U4434 (N_4434,N_3542,N_3863);
nand U4435 (N_4435,N_3500,N_3539);
nand U4436 (N_4436,N_3620,N_3722);
nor U4437 (N_4437,N_3647,N_3862);
nand U4438 (N_4438,N_3819,N_3860);
and U4439 (N_4439,N_3870,N_3901);
and U4440 (N_4440,N_3824,N_3725);
or U4441 (N_4441,N_3947,N_3824);
nand U4442 (N_4442,N_3876,N_3770);
and U4443 (N_4443,N_3679,N_3767);
nand U4444 (N_4444,N_3615,N_3592);
and U4445 (N_4445,N_3542,N_3569);
nor U4446 (N_4446,N_3592,N_3529);
and U4447 (N_4447,N_3614,N_3743);
nor U4448 (N_4448,N_3905,N_3595);
nand U4449 (N_4449,N_3562,N_3869);
or U4450 (N_4450,N_3862,N_3916);
nor U4451 (N_4451,N_3867,N_3504);
and U4452 (N_4452,N_3679,N_3913);
and U4453 (N_4453,N_3976,N_3889);
or U4454 (N_4454,N_3768,N_3715);
or U4455 (N_4455,N_3866,N_3530);
nand U4456 (N_4456,N_3604,N_3592);
nor U4457 (N_4457,N_3601,N_3678);
or U4458 (N_4458,N_3904,N_3939);
nor U4459 (N_4459,N_3667,N_3628);
nand U4460 (N_4460,N_3788,N_3919);
or U4461 (N_4461,N_3604,N_3589);
or U4462 (N_4462,N_3697,N_3691);
nand U4463 (N_4463,N_3776,N_3914);
and U4464 (N_4464,N_3531,N_3529);
nand U4465 (N_4465,N_3778,N_3661);
nor U4466 (N_4466,N_3720,N_3742);
or U4467 (N_4467,N_3739,N_3559);
nor U4468 (N_4468,N_3888,N_3708);
and U4469 (N_4469,N_3775,N_3894);
nor U4470 (N_4470,N_3545,N_3827);
xnor U4471 (N_4471,N_3859,N_3537);
nor U4472 (N_4472,N_3787,N_3875);
and U4473 (N_4473,N_3724,N_3804);
nor U4474 (N_4474,N_3525,N_3707);
and U4475 (N_4475,N_3889,N_3594);
or U4476 (N_4476,N_3987,N_3546);
and U4477 (N_4477,N_3942,N_3830);
and U4478 (N_4478,N_3656,N_3936);
nor U4479 (N_4479,N_3882,N_3857);
xnor U4480 (N_4480,N_3676,N_3905);
nor U4481 (N_4481,N_3784,N_3782);
and U4482 (N_4482,N_3979,N_3522);
nor U4483 (N_4483,N_3591,N_3818);
nor U4484 (N_4484,N_3827,N_3656);
and U4485 (N_4485,N_3781,N_3904);
or U4486 (N_4486,N_3800,N_3540);
nor U4487 (N_4487,N_3625,N_3962);
xnor U4488 (N_4488,N_3643,N_3659);
or U4489 (N_4489,N_3791,N_3512);
nor U4490 (N_4490,N_3771,N_3911);
nor U4491 (N_4491,N_3993,N_3977);
or U4492 (N_4492,N_3917,N_3676);
nand U4493 (N_4493,N_3534,N_3872);
xnor U4494 (N_4494,N_3546,N_3513);
or U4495 (N_4495,N_3614,N_3809);
nor U4496 (N_4496,N_3808,N_3942);
nor U4497 (N_4497,N_3500,N_3940);
nor U4498 (N_4498,N_3573,N_3607);
or U4499 (N_4499,N_3658,N_3661);
nand U4500 (N_4500,N_4405,N_4327);
and U4501 (N_4501,N_4052,N_4152);
and U4502 (N_4502,N_4482,N_4045);
or U4503 (N_4503,N_4461,N_4436);
and U4504 (N_4504,N_4180,N_4046);
or U4505 (N_4505,N_4396,N_4392);
nor U4506 (N_4506,N_4384,N_4300);
nor U4507 (N_4507,N_4053,N_4109);
nand U4508 (N_4508,N_4126,N_4237);
nand U4509 (N_4509,N_4009,N_4273);
nor U4510 (N_4510,N_4067,N_4110);
xor U4511 (N_4511,N_4170,N_4194);
or U4512 (N_4512,N_4199,N_4441);
or U4513 (N_4513,N_4481,N_4262);
nand U4514 (N_4514,N_4062,N_4211);
or U4515 (N_4515,N_4411,N_4054);
nand U4516 (N_4516,N_4032,N_4279);
xor U4517 (N_4517,N_4129,N_4474);
or U4518 (N_4518,N_4426,N_4108);
nor U4519 (N_4519,N_4451,N_4242);
xnor U4520 (N_4520,N_4448,N_4388);
nor U4521 (N_4521,N_4358,N_4381);
nor U4522 (N_4522,N_4408,N_4316);
or U4523 (N_4523,N_4464,N_4489);
nand U4524 (N_4524,N_4150,N_4187);
nor U4525 (N_4525,N_4406,N_4167);
nor U4526 (N_4526,N_4035,N_4233);
nor U4527 (N_4527,N_4382,N_4287);
or U4528 (N_4528,N_4462,N_4076);
and U4529 (N_4529,N_4430,N_4257);
nor U4530 (N_4530,N_4278,N_4413);
xor U4531 (N_4531,N_4341,N_4143);
or U4532 (N_4532,N_4103,N_4339);
nor U4533 (N_4533,N_4386,N_4484);
nor U4534 (N_4534,N_4215,N_4330);
and U4535 (N_4535,N_4185,N_4420);
nand U4536 (N_4536,N_4146,N_4023);
or U4537 (N_4537,N_4348,N_4222);
nor U4538 (N_4538,N_4295,N_4352);
or U4539 (N_4539,N_4266,N_4440);
nand U4540 (N_4540,N_4007,N_4201);
nor U4541 (N_4541,N_4221,N_4228);
nor U4542 (N_4542,N_4059,N_4120);
xnor U4543 (N_4543,N_4472,N_4002);
nor U4544 (N_4544,N_4113,N_4213);
nor U4545 (N_4545,N_4250,N_4207);
and U4546 (N_4546,N_4486,N_4124);
and U4547 (N_4547,N_4027,N_4424);
or U4548 (N_4548,N_4463,N_4227);
and U4549 (N_4549,N_4097,N_4026);
and U4550 (N_4550,N_4226,N_4043);
and U4551 (N_4551,N_4077,N_4274);
and U4552 (N_4552,N_4333,N_4086);
xnor U4553 (N_4553,N_4105,N_4319);
and U4554 (N_4554,N_4323,N_4080);
or U4555 (N_4555,N_4265,N_4070);
and U4556 (N_4556,N_4286,N_4164);
or U4557 (N_4557,N_4219,N_4144);
or U4558 (N_4558,N_4299,N_4082);
or U4559 (N_4559,N_4303,N_4490);
or U4560 (N_4560,N_4181,N_4256);
nor U4561 (N_4561,N_4260,N_4000);
or U4562 (N_4562,N_4336,N_4049);
and U4563 (N_4563,N_4183,N_4083);
nand U4564 (N_4564,N_4387,N_4229);
and U4565 (N_4565,N_4241,N_4363);
nand U4566 (N_4566,N_4056,N_4239);
xor U4567 (N_4567,N_4313,N_4182);
nor U4568 (N_4568,N_4351,N_4141);
nand U4569 (N_4569,N_4494,N_4346);
or U4570 (N_4570,N_4485,N_4368);
or U4571 (N_4571,N_4473,N_4160);
nand U4572 (N_4572,N_4305,N_4453);
and U4573 (N_4573,N_4356,N_4131);
or U4574 (N_4574,N_4285,N_4444);
nor U4575 (N_4575,N_4337,N_4154);
or U4576 (N_4576,N_4499,N_4191);
nor U4577 (N_4577,N_4071,N_4263);
xnor U4578 (N_4578,N_4460,N_4409);
or U4579 (N_4579,N_4040,N_4459);
and U4580 (N_4580,N_4394,N_4497);
or U4581 (N_4581,N_4096,N_4163);
nor U4582 (N_4582,N_4362,N_4322);
or U4583 (N_4583,N_4369,N_4389);
and U4584 (N_4584,N_4024,N_4092);
and U4585 (N_4585,N_4085,N_4496);
xnor U4586 (N_4586,N_4304,N_4427);
or U4587 (N_4587,N_4470,N_4088);
xnor U4588 (N_4588,N_4118,N_4223);
or U4589 (N_4589,N_4335,N_4252);
nor U4590 (N_4590,N_4014,N_4471);
nor U4591 (N_4591,N_4331,N_4412);
xnor U4592 (N_4592,N_4188,N_4296);
nand U4593 (N_4593,N_4375,N_4030);
and U4594 (N_4594,N_4332,N_4061);
and U4595 (N_4595,N_4380,N_4399);
nand U4596 (N_4596,N_4370,N_4385);
nor U4597 (N_4597,N_4282,N_4364);
or U4598 (N_4598,N_4090,N_4031);
nand U4599 (N_4599,N_4224,N_4044);
or U4600 (N_4600,N_4458,N_4344);
or U4601 (N_4601,N_4443,N_4267);
nor U4602 (N_4602,N_4074,N_4102);
and U4603 (N_4603,N_4016,N_4048);
nand U4604 (N_4604,N_4438,N_4452);
or U4605 (N_4605,N_4217,N_4209);
or U4606 (N_4606,N_4039,N_4051);
or U4607 (N_4607,N_4421,N_4140);
nand U4608 (N_4608,N_4005,N_4317);
xor U4609 (N_4609,N_4477,N_4269);
or U4610 (N_4610,N_4121,N_4466);
and U4611 (N_4611,N_4376,N_4095);
and U4612 (N_4612,N_4145,N_4467);
and U4613 (N_4613,N_4135,N_4099);
nor U4614 (N_4614,N_4324,N_4218);
and U4615 (N_4615,N_4417,N_4010);
or U4616 (N_4616,N_4353,N_4243);
and U4617 (N_4617,N_4457,N_4345);
nand U4618 (N_4618,N_4259,N_4329);
nand U4619 (N_4619,N_4249,N_4136);
nor U4620 (N_4620,N_4210,N_4117);
and U4621 (N_4621,N_4360,N_4366);
nand U4622 (N_4622,N_4272,N_4383);
nand U4623 (N_4623,N_4123,N_4147);
or U4624 (N_4624,N_4310,N_4377);
or U4625 (N_4625,N_4315,N_4115);
nand U4626 (N_4626,N_4171,N_4177);
nor U4627 (N_4627,N_4491,N_4212);
or U4628 (N_4628,N_4042,N_4403);
and U4629 (N_4629,N_4078,N_4338);
or U4630 (N_4630,N_4404,N_4127);
or U4631 (N_4631,N_4400,N_4193);
and U4632 (N_4632,N_4214,N_4008);
and U4633 (N_4633,N_4320,N_4238);
nand U4634 (N_4634,N_4268,N_4200);
and U4635 (N_4635,N_4130,N_4186);
nand U4636 (N_4636,N_4166,N_4359);
or U4637 (N_4637,N_4240,N_4020);
or U4638 (N_4638,N_4419,N_4378);
and U4639 (N_4639,N_4068,N_4447);
or U4640 (N_4640,N_4433,N_4301);
nand U4641 (N_4641,N_4205,N_4246);
xor U4642 (N_4642,N_4232,N_4013);
and U4643 (N_4643,N_4373,N_4276);
nand U4644 (N_4644,N_4455,N_4401);
xor U4645 (N_4645,N_4493,N_4047);
nor U4646 (N_4646,N_4098,N_4176);
or U4647 (N_4647,N_4280,N_4283);
and U4648 (N_4648,N_4107,N_4410);
or U4649 (N_4649,N_4197,N_4089);
and U4650 (N_4650,N_4104,N_4060);
nand U4651 (N_4651,N_4153,N_4057);
or U4652 (N_4652,N_4206,N_4340);
nor U4653 (N_4653,N_4270,N_4175);
nor U4654 (N_4654,N_4001,N_4064);
and U4655 (N_4655,N_4137,N_4050);
and U4656 (N_4656,N_4101,N_4157);
nand U4657 (N_4657,N_4398,N_4407);
nor U4658 (N_4658,N_4432,N_4288);
and U4659 (N_4659,N_4036,N_4254);
or U4660 (N_4660,N_4365,N_4289);
or U4661 (N_4661,N_4314,N_4290);
nor U4662 (N_4662,N_4091,N_4343);
or U4663 (N_4663,N_4253,N_4195);
or U4664 (N_4664,N_4084,N_4087);
or U4665 (N_4665,N_4247,N_4367);
and U4666 (N_4666,N_4093,N_4372);
nand U4667 (N_4667,N_4311,N_4498);
or U4668 (N_4668,N_4012,N_4475);
or U4669 (N_4669,N_4423,N_4230);
nand U4670 (N_4670,N_4309,N_4018);
nor U4671 (N_4671,N_4066,N_4015);
and U4672 (N_4672,N_4058,N_4294);
and U4673 (N_4673,N_4255,N_4128);
or U4674 (N_4674,N_4142,N_4302);
xor U4675 (N_4675,N_4161,N_4179);
nand U4676 (N_4676,N_4435,N_4038);
or U4677 (N_4677,N_4029,N_4318);
nand U4678 (N_4678,N_4355,N_4198);
xor U4679 (N_4679,N_4292,N_4306);
nand U4680 (N_4680,N_4347,N_4075);
xnor U4681 (N_4681,N_4321,N_4431);
nand U4682 (N_4682,N_4122,N_4476);
or U4683 (N_4683,N_4468,N_4069);
xor U4684 (N_4684,N_4190,N_4133);
or U4685 (N_4685,N_4449,N_4244);
nor U4686 (N_4686,N_4231,N_4203);
nand U4687 (N_4687,N_4245,N_4202);
nand U4688 (N_4688,N_4132,N_4081);
or U4689 (N_4689,N_4326,N_4293);
or U4690 (N_4690,N_4487,N_4125);
and U4691 (N_4691,N_4418,N_4465);
or U4692 (N_4692,N_4437,N_4196);
nand U4693 (N_4693,N_4158,N_4297);
or U4694 (N_4694,N_4251,N_4445);
or U4695 (N_4695,N_4428,N_4155);
or U4696 (N_4696,N_4357,N_4450);
nor U4697 (N_4697,N_4371,N_4439);
xor U4698 (N_4698,N_4162,N_4139);
nand U4699 (N_4699,N_4172,N_4307);
nor U4700 (N_4700,N_4111,N_4151);
nand U4701 (N_4701,N_4033,N_4277);
nand U4702 (N_4702,N_4350,N_4425);
and U4703 (N_4703,N_4004,N_4034);
nand U4704 (N_4704,N_4192,N_4298);
or U4705 (N_4705,N_4173,N_4395);
nor U4706 (N_4706,N_4434,N_4281);
or U4707 (N_4707,N_4342,N_4479);
nor U4708 (N_4708,N_4422,N_4248);
nand U4709 (N_4709,N_4235,N_4414);
or U4710 (N_4710,N_4159,N_4079);
or U4711 (N_4711,N_4178,N_4165);
nor U4712 (N_4712,N_4119,N_4134);
or U4713 (N_4713,N_4361,N_4156);
or U4714 (N_4714,N_4379,N_4204);
or U4715 (N_4715,N_4374,N_4114);
or U4716 (N_4716,N_4429,N_4258);
nand U4717 (N_4717,N_4446,N_4174);
nor U4718 (N_4718,N_4236,N_4225);
and U4719 (N_4719,N_4011,N_4483);
and U4720 (N_4720,N_4334,N_4003);
xnor U4721 (N_4721,N_4168,N_4284);
and U4722 (N_4722,N_4234,N_4325);
nand U4723 (N_4723,N_4055,N_4492);
and U4724 (N_4724,N_4216,N_4264);
nor U4725 (N_4725,N_4041,N_4402);
xnor U4726 (N_4726,N_4148,N_4022);
and U4727 (N_4727,N_4328,N_4349);
and U4728 (N_4728,N_4100,N_4149);
or U4729 (N_4729,N_4019,N_4469);
nor U4730 (N_4730,N_4312,N_4072);
and U4731 (N_4731,N_4138,N_4189);
or U4732 (N_4732,N_4390,N_4495);
nor U4733 (N_4733,N_4112,N_4065);
nand U4734 (N_4734,N_4275,N_4106);
or U4735 (N_4735,N_4208,N_4456);
and U4736 (N_4736,N_4415,N_4488);
xnor U4737 (N_4737,N_4116,N_4354);
nand U4738 (N_4738,N_4480,N_4063);
nand U4739 (N_4739,N_4073,N_4442);
xor U4740 (N_4740,N_4271,N_4291);
xor U4741 (N_4741,N_4037,N_4393);
or U4742 (N_4742,N_4454,N_4184);
or U4743 (N_4743,N_4220,N_4017);
and U4744 (N_4744,N_4397,N_4261);
nand U4745 (N_4745,N_4478,N_4308);
or U4746 (N_4746,N_4021,N_4169);
nand U4747 (N_4747,N_4391,N_4025);
nand U4748 (N_4748,N_4416,N_4028);
nor U4749 (N_4749,N_4006,N_4094);
xor U4750 (N_4750,N_4094,N_4237);
nand U4751 (N_4751,N_4290,N_4249);
nand U4752 (N_4752,N_4274,N_4497);
nor U4753 (N_4753,N_4386,N_4075);
or U4754 (N_4754,N_4427,N_4457);
and U4755 (N_4755,N_4352,N_4378);
xor U4756 (N_4756,N_4343,N_4444);
and U4757 (N_4757,N_4088,N_4306);
and U4758 (N_4758,N_4441,N_4272);
and U4759 (N_4759,N_4146,N_4129);
nor U4760 (N_4760,N_4396,N_4256);
or U4761 (N_4761,N_4077,N_4197);
or U4762 (N_4762,N_4469,N_4171);
or U4763 (N_4763,N_4383,N_4030);
xnor U4764 (N_4764,N_4352,N_4254);
xor U4765 (N_4765,N_4029,N_4335);
xor U4766 (N_4766,N_4320,N_4079);
or U4767 (N_4767,N_4296,N_4412);
or U4768 (N_4768,N_4278,N_4137);
nand U4769 (N_4769,N_4498,N_4426);
nor U4770 (N_4770,N_4130,N_4387);
or U4771 (N_4771,N_4010,N_4427);
nand U4772 (N_4772,N_4064,N_4367);
nor U4773 (N_4773,N_4363,N_4483);
and U4774 (N_4774,N_4384,N_4127);
nand U4775 (N_4775,N_4071,N_4424);
nand U4776 (N_4776,N_4327,N_4452);
nor U4777 (N_4777,N_4194,N_4301);
nor U4778 (N_4778,N_4360,N_4393);
nor U4779 (N_4779,N_4001,N_4242);
nand U4780 (N_4780,N_4138,N_4224);
or U4781 (N_4781,N_4313,N_4494);
nand U4782 (N_4782,N_4433,N_4212);
nand U4783 (N_4783,N_4218,N_4168);
or U4784 (N_4784,N_4345,N_4430);
or U4785 (N_4785,N_4255,N_4471);
or U4786 (N_4786,N_4312,N_4071);
xnor U4787 (N_4787,N_4110,N_4298);
or U4788 (N_4788,N_4202,N_4206);
and U4789 (N_4789,N_4392,N_4488);
nor U4790 (N_4790,N_4287,N_4391);
nor U4791 (N_4791,N_4002,N_4478);
nand U4792 (N_4792,N_4079,N_4443);
nand U4793 (N_4793,N_4447,N_4099);
nand U4794 (N_4794,N_4071,N_4374);
nand U4795 (N_4795,N_4291,N_4184);
nor U4796 (N_4796,N_4021,N_4495);
nand U4797 (N_4797,N_4290,N_4338);
or U4798 (N_4798,N_4178,N_4122);
nand U4799 (N_4799,N_4328,N_4171);
and U4800 (N_4800,N_4297,N_4126);
xor U4801 (N_4801,N_4492,N_4325);
and U4802 (N_4802,N_4009,N_4280);
xor U4803 (N_4803,N_4325,N_4311);
nor U4804 (N_4804,N_4052,N_4412);
or U4805 (N_4805,N_4261,N_4124);
nor U4806 (N_4806,N_4273,N_4433);
and U4807 (N_4807,N_4240,N_4468);
or U4808 (N_4808,N_4305,N_4001);
nor U4809 (N_4809,N_4284,N_4140);
xor U4810 (N_4810,N_4355,N_4195);
or U4811 (N_4811,N_4316,N_4277);
nand U4812 (N_4812,N_4143,N_4348);
nor U4813 (N_4813,N_4458,N_4090);
xnor U4814 (N_4814,N_4312,N_4294);
and U4815 (N_4815,N_4376,N_4048);
and U4816 (N_4816,N_4065,N_4268);
or U4817 (N_4817,N_4240,N_4497);
nor U4818 (N_4818,N_4203,N_4063);
nand U4819 (N_4819,N_4292,N_4025);
nand U4820 (N_4820,N_4404,N_4403);
and U4821 (N_4821,N_4294,N_4240);
nor U4822 (N_4822,N_4156,N_4420);
nor U4823 (N_4823,N_4457,N_4364);
or U4824 (N_4824,N_4126,N_4473);
nand U4825 (N_4825,N_4105,N_4467);
nand U4826 (N_4826,N_4358,N_4251);
or U4827 (N_4827,N_4137,N_4494);
xnor U4828 (N_4828,N_4345,N_4011);
xor U4829 (N_4829,N_4219,N_4057);
xor U4830 (N_4830,N_4147,N_4232);
nor U4831 (N_4831,N_4297,N_4089);
nor U4832 (N_4832,N_4011,N_4138);
and U4833 (N_4833,N_4429,N_4371);
or U4834 (N_4834,N_4067,N_4416);
and U4835 (N_4835,N_4343,N_4227);
or U4836 (N_4836,N_4320,N_4138);
nor U4837 (N_4837,N_4221,N_4422);
nand U4838 (N_4838,N_4385,N_4259);
nand U4839 (N_4839,N_4340,N_4306);
nand U4840 (N_4840,N_4415,N_4315);
and U4841 (N_4841,N_4153,N_4409);
nor U4842 (N_4842,N_4373,N_4391);
nand U4843 (N_4843,N_4486,N_4043);
and U4844 (N_4844,N_4200,N_4186);
nor U4845 (N_4845,N_4021,N_4424);
or U4846 (N_4846,N_4333,N_4056);
nand U4847 (N_4847,N_4325,N_4354);
nand U4848 (N_4848,N_4391,N_4244);
or U4849 (N_4849,N_4332,N_4186);
or U4850 (N_4850,N_4058,N_4021);
xnor U4851 (N_4851,N_4081,N_4397);
or U4852 (N_4852,N_4096,N_4324);
or U4853 (N_4853,N_4453,N_4152);
or U4854 (N_4854,N_4395,N_4093);
xor U4855 (N_4855,N_4441,N_4227);
xor U4856 (N_4856,N_4117,N_4298);
nand U4857 (N_4857,N_4342,N_4403);
nor U4858 (N_4858,N_4343,N_4466);
nor U4859 (N_4859,N_4343,N_4339);
nor U4860 (N_4860,N_4311,N_4476);
xnor U4861 (N_4861,N_4165,N_4488);
and U4862 (N_4862,N_4202,N_4421);
nand U4863 (N_4863,N_4274,N_4218);
nor U4864 (N_4864,N_4419,N_4016);
nor U4865 (N_4865,N_4075,N_4141);
or U4866 (N_4866,N_4317,N_4201);
or U4867 (N_4867,N_4385,N_4468);
and U4868 (N_4868,N_4304,N_4474);
nor U4869 (N_4869,N_4420,N_4377);
and U4870 (N_4870,N_4250,N_4262);
nor U4871 (N_4871,N_4037,N_4211);
or U4872 (N_4872,N_4323,N_4068);
nand U4873 (N_4873,N_4385,N_4408);
or U4874 (N_4874,N_4305,N_4132);
nand U4875 (N_4875,N_4402,N_4150);
and U4876 (N_4876,N_4174,N_4471);
and U4877 (N_4877,N_4059,N_4341);
and U4878 (N_4878,N_4337,N_4378);
xnor U4879 (N_4879,N_4124,N_4052);
nor U4880 (N_4880,N_4227,N_4079);
or U4881 (N_4881,N_4193,N_4184);
and U4882 (N_4882,N_4131,N_4133);
and U4883 (N_4883,N_4319,N_4431);
and U4884 (N_4884,N_4139,N_4287);
nand U4885 (N_4885,N_4336,N_4461);
nand U4886 (N_4886,N_4211,N_4137);
nor U4887 (N_4887,N_4082,N_4352);
xor U4888 (N_4888,N_4176,N_4390);
xor U4889 (N_4889,N_4046,N_4243);
nor U4890 (N_4890,N_4367,N_4117);
and U4891 (N_4891,N_4474,N_4365);
and U4892 (N_4892,N_4028,N_4089);
or U4893 (N_4893,N_4109,N_4317);
or U4894 (N_4894,N_4190,N_4043);
nand U4895 (N_4895,N_4169,N_4028);
or U4896 (N_4896,N_4365,N_4482);
xor U4897 (N_4897,N_4349,N_4055);
or U4898 (N_4898,N_4027,N_4279);
nor U4899 (N_4899,N_4280,N_4258);
and U4900 (N_4900,N_4195,N_4378);
or U4901 (N_4901,N_4121,N_4314);
nor U4902 (N_4902,N_4319,N_4315);
or U4903 (N_4903,N_4119,N_4031);
nor U4904 (N_4904,N_4491,N_4184);
nand U4905 (N_4905,N_4156,N_4168);
or U4906 (N_4906,N_4325,N_4309);
and U4907 (N_4907,N_4256,N_4028);
and U4908 (N_4908,N_4363,N_4457);
nor U4909 (N_4909,N_4352,N_4348);
and U4910 (N_4910,N_4414,N_4046);
and U4911 (N_4911,N_4299,N_4135);
nor U4912 (N_4912,N_4466,N_4032);
and U4913 (N_4913,N_4285,N_4023);
or U4914 (N_4914,N_4238,N_4000);
nand U4915 (N_4915,N_4236,N_4016);
nor U4916 (N_4916,N_4018,N_4319);
or U4917 (N_4917,N_4203,N_4206);
nand U4918 (N_4918,N_4463,N_4039);
and U4919 (N_4919,N_4065,N_4280);
or U4920 (N_4920,N_4230,N_4265);
or U4921 (N_4921,N_4486,N_4016);
and U4922 (N_4922,N_4081,N_4068);
xor U4923 (N_4923,N_4254,N_4038);
or U4924 (N_4924,N_4109,N_4139);
and U4925 (N_4925,N_4229,N_4443);
or U4926 (N_4926,N_4150,N_4433);
nand U4927 (N_4927,N_4473,N_4325);
xnor U4928 (N_4928,N_4046,N_4388);
and U4929 (N_4929,N_4262,N_4132);
nor U4930 (N_4930,N_4352,N_4376);
and U4931 (N_4931,N_4263,N_4040);
nor U4932 (N_4932,N_4472,N_4333);
xnor U4933 (N_4933,N_4091,N_4264);
or U4934 (N_4934,N_4065,N_4094);
and U4935 (N_4935,N_4350,N_4434);
nand U4936 (N_4936,N_4452,N_4480);
nand U4937 (N_4937,N_4489,N_4437);
nor U4938 (N_4938,N_4253,N_4040);
or U4939 (N_4939,N_4043,N_4351);
nand U4940 (N_4940,N_4248,N_4049);
and U4941 (N_4941,N_4357,N_4488);
xor U4942 (N_4942,N_4071,N_4333);
or U4943 (N_4943,N_4346,N_4373);
and U4944 (N_4944,N_4267,N_4126);
and U4945 (N_4945,N_4131,N_4194);
nand U4946 (N_4946,N_4099,N_4386);
or U4947 (N_4947,N_4295,N_4161);
nand U4948 (N_4948,N_4327,N_4393);
and U4949 (N_4949,N_4023,N_4074);
nor U4950 (N_4950,N_4317,N_4087);
nand U4951 (N_4951,N_4197,N_4321);
or U4952 (N_4952,N_4348,N_4069);
nand U4953 (N_4953,N_4150,N_4434);
nand U4954 (N_4954,N_4293,N_4345);
and U4955 (N_4955,N_4195,N_4088);
nor U4956 (N_4956,N_4070,N_4495);
or U4957 (N_4957,N_4002,N_4163);
or U4958 (N_4958,N_4025,N_4367);
or U4959 (N_4959,N_4334,N_4182);
nor U4960 (N_4960,N_4011,N_4176);
nand U4961 (N_4961,N_4337,N_4090);
or U4962 (N_4962,N_4386,N_4058);
and U4963 (N_4963,N_4475,N_4453);
and U4964 (N_4964,N_4258,N_4105);
and U4965 (N_4965,N_4251,N_4151);
xor U4966 (N_4966,N_4277,N_4010);
and U4967 (N_4967,N_4419,N_4333);
nand U4968 (N_4968,N_4027,N_4076);
nand U4969 (N_4969,N_4011,N_4436);
nor U4970 (N_4970,N_4079,N_4153);
and U4971 (N_4971,N_4434,N_4100);
and U4972 (N_4972,N_4117,N_4354);
or U4973 (N_4973,N_4189,N_4333);
and U4974 (N_4974,N_4177,N_4002);
nor U4975 (N_4975,N_4481,N_4425);
or U4976 (N_4976,N_4057,N_4389);
nor U4977 (N_4977,N_4326,N_4227);
and U4978 (N_4978,N_4120,N_4224);
nor U4979 (N_4979,N_4396,N_4472);
and U4980 (N_4980,N_4378,N_4388);
and U4981 (N_4981,N_4108,N_4156);
nor U4982 (N_4982,N_4416,N_4499);
or U4983 (N_4983,N_4261,N_4205);
nor U4984 (N_4984,N_4247,N_4414);
nor U4985 (N_4985,N_4450,N_4484);
and U4986 (N_4986,N_4166,N_4489);
xnor U4987 (N_4987,N_4335,N_4108);
nand U4988 (N_4988,N_4118,N_4339);
nand U4989 (N_4989,N_4266,N_4100);
nor U4990 (N_4990,N_4275,N_4142);
nand U4991 (N_4991,N_4123,N_4462);
nor U4992 (N_4992,N_4131,N_4109);
and U4993 (N_4993,N_4217,N_4080);
or U4994 (N_4994,N_4100,N_4455);
and U4995 (N_4995,N_4153,N_4242);
and U4996 (N_4996,N_4210,N_4169);
or U4997 (N_4997,N_4260,N_4427);
nor U4998 (N_4998,N_4282,N_4324);
or U4999 (N_4999,N_4193,N_4499);
nor UO_0 (O_0,N_4709,N_4704);
or UO_1 (O_1,N_4945,N_4647);
nand UO_2 (O_2,N_4610,N_4719);
nand UO_3 (O_3,N_4726,N_4555);
nand UO_4 (O_4,N_4788,N_4768);
nor UO_5 (O_5,N_4894,N_4966);
and UO_6 (O_6,N_4955,N_4921);
nor UO_7 (O_7,N_4774,N_4986);
nor UO_8 (O_8,N_4531,N_4622);
nand UO_9 (O_9,N_4965,N_4889);
nor UO_10 (O_10,N_4918,N_4868);
nor UO_11 (O_11,N_4637,N_4938);
and UO_12 (O_12,N_4548,N_4526);
nand UO_13 (O_13,N_4642,N_4946);
and UO_14 (O_14,N_4716,N_4685);
or UO_15 (O_15,N_4663,N_4924);
xnor UO_16 (O_16,N_4883,N_4939);
and UO_17 (O_17,N_4739,N_4999);
or UO_18 (O_18,N_4944,N_4783);
nor UO_19 (O_19,N_4613,N_4862);
and UO_20 (O_20,N_4961,N_4780);
and UO_21 (O_21,N_4648,N_4640);
nor UO_22 (O_22,N_4651,N_4970);
or UO_23 (O_23,N_4718,N_4702);
and UO_24 (O_24,N_4627,N_4754);
or UO_25 (O_25,N_4933,N_4577);
nor UO_26 (O_26,N_4818,N_4821);
xnor UO_27 (O_27,N_4779,N_4776);
xnor UO_28 (O_28,N_4614,N_4811);
or UO_29 (O_29,N_4595,N_4512);
nand UO_30 (O_30,N_4993,N_4596);
nand UO_31 (O_31,N_4802,N_4520);
nor UO_32 (O_32,N_4517,N_4974);
xor UO_33 (O_33,N_4644,N_4529);
xnor UO_34 (O_34,N_4851,N_4571);
and UO_35 (O_35,N_4792,N_4837);
nand UO_36 (O_36,N_4757,N_4592);
xnor UO_37 (O_37,N_4748,N_4987);
nor UO_38 (O_38,N_4806,N_4952);
and UO_39 (O_39,N_4960,N_4675);
or UO_40 (O_40,N_4926,N_4925);
and UO_41 (O_41,N_4705,N_4735);
nor UO_42 (O_42,N_4805,N_4782);
xor UO_43 (O_43,N_4605,N_4988);
and UO_44 (O_44,N_4809,N_4803);
and UO_45 (O_45,N_4654,N_4764);
or UO_46 (O_46,N_4681,N_4971);
and UO_47 (O_47,N_4729,N_4917);
xor UO_48 (O_48,N_4597,N_4847);
nand UO_49 (O_49,N_4706,N_4752);
or UO_50 (O_50,N_4633,N_4701);
or UO_51 (O_51,N_4893,N_4948);
or UO_52 (O_52,N_4879,N_4601);
nand UO_53 (O_53,N_4690,N_4515);
and UO_54 (O_54,N_4852,N_4674);
and UO_55 (O_55,N_4725,N_4843);
nand UO_56 (O_56,N_4985,N_4968);
and UO_57 (O_57,N_4510,N_4677);
and UO_58 (O_58,N_4694,N_4907);
or UO_59 (O_59,N_4669,N_4877);
nand UO_60 (O_60,N_4858,N_4765);
nand UO_61 (O_61,N_4699,N_4972);
or UO_62 (O_62,N_4742,N_4934);
nor UO_63 (O_63,N_4861,N_4778);
nand UO_64 (O_64,N_4857,N_4874);
and UO_65 (O_65,N_4824,N_4813);
nand UO_66 (O_66,N_4591,N_4903);
or UO_67 (O_67,N_4682,N_4747);
and UO_68 (O_68,N_4902,N_4935);
and UO_69 (O_69,N_4579,N_4700);
xnor UO_70 (O_70,N_4880,N_4822);
xor UO_71 (O_71,N_4530,N_4814);
nand UO_72 (O_72,N_4562,N_4980);
or UO_73 (O_73,N_4570,N_4881);
nor UO_74 (O_74,N_4996,N_4745);
or UO_75 (O_75,N_4664,N_4661);
or UO_76 (O_76,N_4975,N_4582);
nand UO_77 (O_77,N_4528,N_4513);
and UO_78 (O_78,N_4932,N_4937);
and UO_79 (O_79,N_4667,N_4775);
xor UO_80 (O_80,N_4964,N_4626);
xnor UO_81 (O_81,N_4888,N_4798);
nand UO_82 (O_82,N_4770,N_4891);
nand UO_83 (O_83,N_4656,N_4947);
and UO_84 (O_84,N_4662,N_4679);
xor UO_85 (O_85,N_4636,N_4519);
and UO_86 (O_86,N_4741,N_4936);
and UO_87 (O_87,N_4619,N_4500);
nand UO_88 (O_88,N_4550,N_4635);
or UO_89 (O_89,N_4652,N_4722);
nor UO_90 (O_90,N_4542,N_4547);
nand UO_91 (O_91,N_4854,N_4624);
or UO_92 (O_92,N_4839,N_4749);
nand UO_93 (O_93,N_4866,N_4671);
and UO_94 (O_94,N_4557,N_4872);
or UO_95 (O_95,N_4816,N_4608);
or UO_96 (O_96,N_4695,N_4643);
nand UO_97 (O_97,N_4953,N_4620);
nand UO_98 (O_98,N_4958,N_4721);
or UO_99 (O_99,N_4501,N_4545);
nand UO_100 (O_100,N_4668,N_4766);
and UO_101 (O_101,N_4876,N_4537);
nor UO_102 (O_102,N_4929,N_4900);
nand UO_103 (O_103,N_4949,N_4587);
or UO_104 (O_104,N_4532,N_4767);
or UO_105 (O_105,N_4586,N_4518);
and UO_106 (O_106,N_4540,N_4576);
nor UO_107 (O_107,N_4559,N_4914);
or UO_108 (O_108,N_4732,N_4777);
or UO_109 (O_109,N_4896,N_4994);
or UO_110 (O_110,N_4838,N_4689);
or UO_111 (O_111,N_4680,N_4859);
nand UO_112 (O_112,N_4871,N_4919);
xor UO_113 (O_113,N_4713,N_4819);
and UO_114 (O_114,N_4808,N_4686);
nand UO_115 (O_115,N_4912,N_4621);
nand UO_116 (O_116,N_4503,N_4916);
nand UO_117 (O_117,N_4931,N_4940);
nand UO_118 (O_118,N_4920,N_4594);
or UO_119 (O_119,N_4790,N_4795);
or UO_120 (O_120,N_4556,N_4720);
or UO_121 (O_121,N_4533,N_4567);
or UO_122 (O_122,N_4524,N_4504);
nand UO_123 (O_123,N_4830,N_4717);
nand UO_124 (O_124,N_4575,N_4738);
xor UO_125 (O_125,N_4578,N_4962);
nor UO_126 (O_126,N_4554,N_4727);
or UO_127 (O_127,N_4590,N_4516);
or UO_128 (O_128,N_4864,N_4606);
or UO_129 (O_129,N_4923,N_4823);
and UO_130 (O_130,N_4616,N_4973);
and UO_131 (O_131,N_4801,N_4565);
nor UO_132 (O_132,N_4804,N_4740);
nor UO_133 (O_133,N_4511,N_4909);
nor UO_134 (O_134,N_4989,N_4631);
and UO_135 (O_135,N_4899,N_4525);
or UO_136 (O_136,N_4574,N_4760);
nand UO_137 (O_137,N_4885,N_4820);
nor UO_138 (O_138,N_4653,N_4855);
nand UO_139 (O_139,N_4981,N_4875);
and UO_140 (O_140,N_4698,N_4927);
nor UO_141 (O_141,N_4505,N_4826);
and UO_142 (O_142,N_4755,N_4956);
or UO_143 (O_143,N_4551,N_4743);
nor UO_144 (O_144,N_4672,N_4746);
nand UO_145 (O_145,N_4625,N_4734);
nand UO_146 (O_146,N_4865,N_4604);
nor UO_147 (O_147,N_4509,N_4673);
or UO_148 (O_148,N_4657,N_4645);
xnor UO_149 (O_149,N_4870,N_4541);
or UO_150 (O_150,N_4990,N_4609);
or UO_151 (O_151,N_4623,N_4585);
xor UO_152 (O_152,N_4997,N_4560);
nor UO_153 (O_153,N_4771,N_4794);
nand UO_154 (O_154,N_4791,N_4750);
or UO_155 (O_155,N_4841,N_4629);
and UO_156 (O_156,N_4569,N_4660);
or UO_157 (O_157,N_4963,N_4753);
nand UO_158 (O_158,N_4688,N_4723);
xnor UO_159 (O_159,N_4827,N_4632);
nor UO_160 (O_160,N_4611,N_4913);
and UO_161 (O_161,N_4762,N_4710);
nand UO_162 (O_162,N_4995,N_4976);
and UO_163 (O_163,N_4593,N_4763);
or UO_164 (O_164,N_4670,N_4853);
or UO_165 (O_165,N_4901,N_4712);
and UO_166 (O_166,N_4810,N_4869);
nand UO_167 (O_167,N_4967,N_4835);
nor UO_168 (O_168,N_4552,N_4845);
and UO_169 (O_169,N_4930,N_4897);
xnor UO_170 (O_170,N_4527,N_4915);
and UO_171 (O_171,N_4646,N_4544);
or UO_172 (O_172,N_4922,N_4737);
nand UO_173 (O_173,N_4507,N_4641);
nand UO_174 (O_174,N_4799,N_4807);
and UO_175 (O_175,N_4558,N_4583);
and UO_176 (O_176,N_4812,N_4584);
and UO_177 (O_177,N_4566,N_4756);
xor UO_178 (O_178,N_4856,N_4844);
nor UO_179 (O_179,N_4744,N_4772);
nor UO_180 (O_180,N_4957,N_4733);
nor UO_181 (O_181,N_4906,N_4508);
nand UO_182 (O_182,N_4886,N_4905);
nand UO_183 (O_183,N_4665,N_4607);
nand UO_184 (O_184,N_4815,N_4781);
nand UO_185 (O_185,N_4796,N_4829);
xor UO_186 (O_186,N_4943,N_4730);
and UO_187 (O_187,N_4834,N_4959);
or UO_188 (O_188,N_4860,N_4573);
nand UO_189 (O_189,N_4969,N_4724);
nor UO_190 (O_190,N_4867,N_4715);
nand UO_191 (O_191,N_4797,N_4534);
or UO_192 (O_192,N_4898,N_4836);
nand UO_193 (O_193,N_4840,N_4683);
and UO_194 (O_194,N_4785,N_4950);
nand UO_195 (O_195,N_4659,N_4884);
nor UO_196 (O_196,N_4800,N_4863);
nor UO_197 (O_197,N_4612,N_4979);
nor UO_198 (O_198,N_4758,N_4603);
or UO_199 (O_199,N_4588,N_4568);
xnor UO_200 (O_200,N_4638,N_4650);
or UO_201 (O_201,N_4696,N_4842);
nor UO_202 (O_202,N_4951,N_4983);
xor UO_203 (O_203,N_4506,N_4878);
and UO_204 (O_204,N_4954,N_4572);
or UO_205 (O_205,N_4546,N_4882);
nand UO_206 (O_206,N_4684,N_4848);
nor UO_207 (O_207,N_4887,N_4911);
and UO_208 (O_208,N_4978,N_4817);
nor UO_209 (O_209,N_4850,N_4666);
nand UO_210 (O_210,N_4536,N_4831);
xnor UO_211 (O_211,N_4543,N_4787);
nand UO_212 (O_212,N_4984,N_4890);
nand UO_213 (O_213,N_4761,N_4873);
and UO_214 (O_214,N_4703,N_4786);
nand UO_215 (O_215,N_4908,N_4580);
nand UO_216 (O_216,N_4904,N_4676);
xor UO_217 (O_217,N_4895,N_4617);
or UO_218 (O_218,N_4514,N_4849);
or UO_219 (O_219,N_4581,N_4692);
nand UO_220 (O_220,N_4521,N_4563);
nor UO_221 (O_221,N_4691,N_4649);
nand UO_222 (O_222,N_4564,N_4910);
nand UO_223 (O_223,N_4678,N_4832);
nor UO_224 (O_224,N_4553,N_4535);
or UO_225 (O_225,N_4707,N_4846);
nor UO_226 (O_226,N_4708,N_4991);
and UO_227 (O_227,N_4714,N_4634);
and UO_228 (O_228,N_4539,N_4825);
and UO_229 (O_229,N_4538,N_4784);
and UO_230 (O_230,N_4598,N_4828);
or UO_231 (O_231,N_4736,N_4589);
xnor UO_232 (O_232,N_4561,N_4618);
xnor UO_233 (O_233,N_4523,N_4693);
nand UO_234 (O_234,N_4769,N_4615);
nor UO_235 (O_235,N_4928,N_4982);
and UO_236 (O_236,N_4773,N_4711);
xor UO_237 (O_237,N_4751,N_4639);
nor UO_238 (O_238,N_4502,N_4942);
nor UO_239 (O_239,N_4977,N_4602);
nor UO_240 (O_240,N_4628,N_4892);
nand UO_241 (O_241,N_4599,N_4658);
nand UO_242 (O_242,N_4549,N_4687);
or UO_243 (O_243,N_4522,N_4759);
and UO_244 (O_244,N_4789,N_4793);
and UO_245 (O_245,N_4998,N_4833);
nand UO_246 (O_246,N_4728,N_4731);
nand UO_247 (O_247,N_4941,N_4992);
or UO_248 (O_248,N_4655,N_4697);
nor UO_249 (O_249,N_4600,N_4630);
xnor UO_250 (O_250,N_4733,N_4868);
and UO_251 (O_251,N_4790,N_4922);
xnor UO_252 (O_252,N_4987,N_4711);
and UO_253 (O_253,N_4927,N_4601);
nand UO_254 (O_254,N_4840,N_4686);
or UO_255 (O_255,N_4991,N_4574);
nand UO_256 (O_256,N_4880,N_4859);
and UO_257 (O_257,N_4839,N_4806);
and UO_258 (O_258,N_4807,N_4594);
xor UO_259 (O_259,N_4926,N_4538);
nor UO_260 (O_260,N_4784,N_4512);
or UO_261 (O_261,N_4971,N_4734);
nor UO_262 (O_262,N_4612,N_4654);
xnor UO_263 (O_263,N_4846,N_4977);
or UO_264 (O_264,N_4571,N_4830);
nand UO_265 (O_265,N_4951,N_4990);
and UO_266 (O_266,N_4897,N_4765);
xor UO_267 (O_267,N_4781,N_4674);
or UO_268 (O_268,N_4848,N_4933);
nor UO_269 (O_269,N_4793,N_4508);
or UO_270 (O_270,N_4501,N_4852);
and UO_271 (O_271,N_4879,N_4537);
and UO_272 (O_272,N_4755,N_4664);
nor UO_273 (O_273,N_4893,N_4600);
nand UO_274 (O_274,N_4541,N_4775);
nand UO_275 (O_275,N_4707,N_4991);
nand UO_276 (O_276,N_4922,N_4729);
or UO_277 (O_277,N_4770,N_4505);
and UO_278 (O_278,N_4604,N_4836);
and UO_279 (O_279,N_4965,N_4863);
or UO_280 (O_280,N_4631,N_4605);
and UO_281 (O_281,N_4636,N_4611);
nand UO_282 (O_282,N_4752,N_4866);
and UO_283 (O_283,N_4593,N_4552);
nand UO_284 (O_284,N_4709,N_4831);
nor UO_285 (O_285,N_4636,N_4873);
or UO_286 (O_286,N_4623,N_4722);
xnor UO_287 (O_287,N_4687,N_4737);
and UO_288 (O_288,N_4669,N_4545);
nand UO_289 (O_289,N_4901,N_4778);
nand UO_290 (O_290,N_4627,N_4577);
nor UO_291 (O_291,N_4825,N_4922);
or UO_292 (O_292,N_4516,N_4861);
or UO_293 (O_293,N_4594,N_4770);
nor UO_294 (O_294,N_4613,N_4893);
and UO_295 (O_295,N_4569,N_4675);
nor UO_296 (O_296,N_4991,N_4716);
or UO_297 (O_297,N_4548,N_4973);
nor UO_298 (O_298,N_4984,N_4628);
nor UO_299 (O_299,N_4597,N_4672);
nor UO_300 (O_300,N_4950,N_4510);
nand UO_301 (O_301,N_4502,N_4804);
and UO_302 (O_302,N_4884,N_4862);
nor UO_303 (O_303,N_4581,N_4753);
nand UO_304 (O_304,N_4757,N_4676);
nor UO_305 (O_305,N_4799,N_4923);
nand UO_306 (O_306,N_4651,N_4663);
and UO_307 (O_307,N_4502,N_4769);
or UO_308 (O_308,N_4670,N_4813);
and UO_309 (O_309,N_4996,N_4722);
nor UO_310 (O_310,N_4831,N_4705);
or UO_311 (O_311,N_4592,N_4761);
or UO_312 (O_312,N_4979,N_4850);
nand UO_313 (O_313,N_4671,N_4710);
or UO_314 (O_314,N_4984,N_4505);
and UO_315 (O_315,N_4867,N_4596);
nor UO_316 (O_316,N_4849,N_4529);
or UO_317 (O_317,N_4947,N_4969);
and UO_318 (O_318,N_4685,N_4809);
nor UO_319 (O_319,N_4996,N_4820);
nor UO_320 (O_320,N_4832,N_4609);
xor UO_321 (O_321,N_4960,N_4747);
nor UO_322 (O_322,N_4613,N_4780);
and UO_323 (O_323,N_4996,N_4943);
xnor UO_324 (O_324,N_4649,N_4785);
nand UO_325 (O_325,N_4776,N_4944);
or UO_326 (O_326,N_4730,N_4700);
nor UO_327 (O_327,N_4776,N_4898);
and UO_328 (O_328,N_4978,N_4782);
nor UO_329 (O_329,N_4983,N_4707);
or UO_330 (O_330,N_4858,N_4608);
xor UO_331 (O_331,N_4722,N_4594);
and UO_332 (O_332,N_4642,N_4756);
or UO_333 (O_333,N_4607,N_4937);
and UO_334 (O_334,N_4708,N_4511);
and UO_335 (O_335,N_4898,N_4665);
nand UO_336 (O_336,N_4883,N_4546);
or UO_337 (O_337,N_4684,N_4739);
nor UO_338 (O_338,N_4619,N_4972);
or UO_339 (O_339,N_4653,N_4627);
or UO_340 (O_340,N_4643,N_4915);
nand UO_341 (O_341,N_4990,N_4547);
and UO_342 (O_342,N_4671,N_4691);
xor UO_343 (O_343,N_4596,N_4919);
nand UO_344 (O_344,N_4653,N_4576);
nor UO_345 (O_345,N_4850,N_4746);
or UO_346 (O_346,N_4680,N_4932);
or UO_347 (O_347,N_4549,N_4660);
and UO_348 (O_348,N_4543,N_4801);
nand UO_349 (O_349,N_4729,N_4581);
nand UO_350 (O_350,N_4865,N_4927);
xnor UO_351 (O_351,N_4599,N_4558);
nand UO_352 (O_352,N_4869,N_4665);
and UO_353 (O_353,N_4977,N_4831);
or UO_354 (O_354,N_4505,N_4659);
and UO_355 (O_355,N_4990,N_4939);
nor UO_356 (O_356,N_4850,N_4571);
or UO_357 (O_357,N_4706,N_4749);
nand UO_358 (O_358,N_4889,N_4659);
nor UO_359 (O_359,N_4559,N_4666);
nor UO_360 (O_360,N_4741,N_4986);
nor UO_361 (O_361,N_4537,N_4506);
and UO_362 (O_362,N_4656,N_4865);
nand UO_363 (O_363,N_4679,N_4629);
nand UO_364 (O_364,N_4969,N_4719);
nand UO_365 (O_365,N_4513,N_4788);
or UO_366 (O_366,N_4517,N_4516);
nor UO_367 (O_367,N_4799,N_4969);
nor UO_368 (O_368,N_4716,N_4743);
and UO_369 (O_369,N_4577,N_4745);
or UO_370 (O_370,N_4557,N_4912);
and UO_371 (O_371,N_4697,N_4996);
nor UO_372 (O_372,N_4599,N_4502);
nor UO_373 (O_373,N_4501,N_4675);
or UO_374 (O_374,N_4740,N_4648);
and UO_375 (O_375,N_4754,N_4975);
nor UO_376 (O_376,N_4746,N_4996);
xnor UO_377 (O_377,N_4769,N_4720);
and UO_378 (O_378,N_4656,N_4963);
or UO_379 (O_379,N_4811,N_4843);
and UO_380 (O_380,N_4855,N_4518);
or UO_381 (O_381,N_4684,N_4672);
nor UO_382 (O_382,N_4991,N_4992);
and UO_383 (O_383,N_4987,N_4884);
nand UO_384 (O_384,N_4608,N_4926);
and UO_385 (O_385,N_4985,N_4866);
nor UO_386 (O_386,N_4772,N_4593);
and UO_387 (O_387,N_4690,N_4526);
nor UO_388 (O_388,N_4671,N_4887);
nor UO_389 (O_389,N_4840,N_4667);
or UO_390 (O_390,N_4834,N_4769);
and UO_391 (O_391,N_4757,N_4966);
xnor UO_392 (O_392,N_4692,N_4901);
nand UO_393 (O_393,N_4984,N_4596);
nand UO_394 (O_394,N_4705,N_4801);
xor UO_395 (O_395,N_4620,N_4732);
nor UO_396 (O_396,N_4658,N_4808);
nand UO_397 (O_397,N_4526,N_4897);
nor UO_398 (O_398,N_4954,N_4773);
nand UO_399 (O_399,N_4535,N_4675);
nor UO_400 (O_400,N_4755,N_4646);
nand UO_401 (O_401,N_4965,N_4755);
nand UO_402 (O_402,N_4552,N_4546);
xnor UO_403 (O_403,N_4749,N_4766);
nor UO_404 (O_404,N_4905,N_4767);
xnor UO_405 (O_405,N_4870,N_4861);
or UO_406 (O_406,N_4594,N_4850);
nor UO_407 (O_407,N_4768,N_4903);
nand UO_408 (O_408,N_4689,N_4984);
and UO_409 (O_409,N_4658,N_4639);
and UO_410 (O_410,N_4792,N_4960);
xnor UO_411 (O_411,N_4909,N_4689);
nand UO_412 (O_412,N_4509,N_4712);
and UO_413 (O_413,N_4868,N_4631);
nor UO_414 (O_414,N_4989,N_4566);
or UO_415 (O_415,N_4968,N_4807);
or UO_416 (O_416,N_4923,N_4895);
and UO_417 (O_417,N_4785,N_4772);
nand UO_418 (O_418,N_4544,N_4521);
nor UO_419 (O_419,N_4623,N_4965);
nor UO_420 (O_420,N_4672,N_4707);
nor UO_421 (O_421,N_4868,N_4706);
and UO_422 (O_422,N_4759,N_4859);
nor UO_423 (O_423,N_4956,N_4759);
nor UO_424 (O_424,N_4724,N_4753);
nor UO_425 (O_425,N_4694,N_4683);
and UO_426 (O_426,N_4735,N_4933);
xnor UO_427 (O_427,N_4518,N_4932);
or UO_428 (O_428,N_4972,N_4903);
and UO_429 (O_429,N_4788,N_4887);
xor UO_430 (O_430,N_4650,N_4657);
nor UO_431 (O_431,N_4584,N_4799);
nor UO_432 (O_432,N_4568,N_4728);
and UO_433 (O_433,N_4666,N_4501);
or UO_434 (O_434,N_4549,N_4878);
xor UO_435 (O_435,N_4579,N_4705);
nor UO_436 (O_436,N_4720,N_4896);
and UO_437 (O_437,N_4575,N_4550);
and UO_438 (O_438,N_4602,N_4937);
or UO_439 (O_439,N_4804,N_4913);
and UO_440 (O_440,N_4624,N_4514);
and UO_441 (O_441,N_4782,N_4596);
or UO_442 (O_442,N_4832,N_4837);
and UO_443 (O_443,N_4863,N_4923);
or UO_444 (O_444,N_4649,N_4585);
nand UO_445 (O_445,N_4531,N_4555);
or UO_446 (O_446,N_4561,N_4996);
nand UO_447 (O_447,N_4683,N_4661);
or UO_448 (O_448,N_4524,N_4841);
and UO_449 (O_449,N_4759,N_4908);
nor UO_450 (O_450,N_4588,N_4761);
or UO_451 (O_451,N_4550,N_4732);
and UO_452 (O_452,N_4510,N_4636);
nand UO_453 (O_453,N_4616,N_4527);
nor UO_454 (O_454,N_4641,N_4529);
or UO_455 (O_455,N_4665,N_4800);
and UO_456 (O_456,N_4975,N_4543);
nand UO_457 (O_457,N_4620,N_4750);
or UO_458 (O_458,N_4717,N_4581);
nor UO_459 (O_459,N_4559,N_4574);
and UO_460 (O_460,N_4937,N_4595);
nand UO_461 (O_461,N_4800,N_4964);
xor UO_462 (O_462,N_4688,N_4938);
or UO_463 (O_463,N_4712,N_4657);
or UO_464 (O_464,N_4929,N_4627);
or UO_465 (O_465,N_4523,N_4615);
nand UO_466 (O_466,N_4995,N_4541);
and UO_467 (O_467,N_4878,N_4900);
or UO_468 (O_468,N_4671,N_4888);
or UO_469 (O_469,N_4780,N_4528);
or UO_470 (O_470,N_4644,N_4612);
nand UO_471 (O_471,N_4716,N_4785);
or UO_472 (O_472,N_4810,N_4950);
xnor UO_473 (O_473,N_4998,N_4525);
or UO_474 (O_474,N_4921,N_4614);
nand UO_475 (O_475,N_4570,N_4599);
nand UO_476 (O_476,N_4983,N_4767);
nor UO_477 (O_477,N_4931,N_4786);
and UO_478 (O_478,N_4796,N_4972);
nor UO_479 (O_479,N_4551,N_4970);
nor UO_480 (O_480,N_4664,N_4932);
nand UO_481 (O_481,N_4977,N_4964);
and UO_482 (O_482,N_4847,N_4941);
nor UO_483 (O_483,N_4732,N_4505);
nor UO_484 (O_484,N_4834,N_4600);
nor UO_485 (O_485,N_4633,N_4803);
and UO_486 (O_486,N_4634,N_4823);
or UO_487 (O_487,N_4796,N_4802);
nand UO_488 (O_488,N_4794,N_4532);
nand UO_489 (O_489,N_4754,N_4534);
nand UO_490 (O_490,N_4927,N_4733);
and UO_491 (O_491,N_4519,N_4713);
nand UO_492 (O_492,N_4585,N_4804);
nor UO_493 (O_493,N_4740,N_4699);
or UO_494 (O_494,N_4758,N_4990);
nand UO_495 (O_495,N_4914,N_4798);
or UO_496 (O_496,N_4595,N_4730);
nand UO_497 (O_497,N_4632,N_4949);
nand UO_498 (O_498,N_4671,N_4551);
and UO_499 (O_499,N_4732,N_4855);
or UO_500 (O_500,N_4550,N_4910);
and UO_501 (O_501,N_4687,N_4758);
nand UO_502 (O_502,N_4911,N_4575);
nor UO_503 (O_503,N_4764,N_4547);
or UO_504 (O_504,N_4631,N_4571);
and UO_505 (O_505,N_4559,N_4602);
xor UO_506 (O_506,N_4610,N_4977);
or UO_507 (O_507,N_4806,N_4916);
xor UO_508 (O_508,N_4863,N_4540);
nand UO_509 (O_509,N_4583,N_4801);
and UO_510 (O_510,N_4618,N_4763);
or UO_511 (O_511,N_4954,N_4949);
nand UO_512 (O_512,N_4816,N_4574);
and UO_513 (O_513,N_4893,N_4508);
nor UO_514 (O_514,N_4785,N_4854);
xnor UO_515 (O_515,N_4856,N_4593);
and UO_516 (O_516,N_4960,N_4924);
nand UO_517 (O_517,N_4948,N_4667);
and UO_518 (O_518,N_4571,N_4918);
xnor UO_519 (O_519,N_4614,N_4827);
and UO_520 (O_520,N_4984,N_4811);
and UO_521 (O_521,N_4781,N_4543);
nor UO_522 (O_522,N_4763,N_4613);
nor UO_523 (O_523,N_4962,N_4888);
xor UO_524 (O_524,N_4522,N_4933);
and UO_525 (O_525,N_4597,N_4733);
nand UO_526 (O_526,N_4657,N_4900);
or UO_527 (O_527,N_4973,N_4708);
nand UO_528 (O_528,N_4803,N_4683);
and UO_529 (O_529,N_4655,N_4554);
nand UO_530 (O_530,N_4748,N_4689);
nand UO_531 (O_531,N_4905,N_4785);
or UO_532 (O_532,N_4772,N_4545);
and UO_533 (O_533,N_4983,N_4552);
and UO_534 (O_534,N_4910,N_4545);
and UO_535 (O_535,N_4778,N_4603);
nand UO_536 (O_536,N_4567,N_4676);
nor UO_537 (O_537,N_4993,N_4824);
and UO_538 (O_538,N_4702,N_4592);
nand UO_539 (O_539,N_4695,N_4657);
nor UO_540 (O_540,N_4677,N_4783);
and UO_541 (O_541,N_4975,N_4691);
and UO_542 (O_542,N_4651,N_4734);
nand UO_543 (O_543,N_4751,N_4714);
and UO_544 (O_544,N_4771,N_4791);
nor UO_545 (O_545,N_4848,N_4586);
nor UO_546 (O_546,N_4897,N_4984);
and UO_547 (O_547,N_4924,N_4530);
nor UO_548 (O_548,N_4844,N_4752);
xor UO_549 (O_549,N_4761,N_4862);
and UO_550 (O_550,N_4642,N_4528);
or UO_551 (O_551,N_4754,N_4727);
nand UO_552 (O_552,N_4831,N_4859);
nor UO_553 (O_553,N_4595,N_4783);
nand UO_554 (O_554,N_4602,N_4632);
nand UO_555 (O_555,N_4811,N_4846);
and UO_556 (O_556,N_4533,N_4603);
or UO_557 (O_557,N_4904,N_4908);
xnor UO_558 (O_558,N_4609,N_4724);
and UO_559 (O_559,N_4752,N_4731);
nor UO_560 (O_560,N_4935,N_4704);
and UO_561 (O_561,N_4761,N_4667);
nand UO_562 (O_562,N_4958,N_4678);
nand UO_563 (O_563,N_4732,N_4911);
or UO_564 (O_564,N_4762,N_4854);
or UO_565 (O_565,N_4966,N_4578);
nor UO_566 (O_566,N_4712,N_4552);
or UO_567 (O_567,N_4693,N_4676);
nor UO_568 (O_568,N_4602,N_4556);
nand UO_569 (O_569,N_4863,N_4996);
and UO_570 (O_570,N_4636,N_4925);
nand UO_571 (O_571,N_4568,N_4594);
nor UO_572 (O_572,N_4925,N_4530);
nor UO_573 (O_573,N_4890,N_4945);
nand UO_574 (O_574,N_4846,N_4550);
nor UO_575 (O_575,N_4698,N_4702);
nor UO_576 (O_576,N_4889,N_4529);
nor UO_577 (O_577,N_4723,N_4974);
nor UO_578 (O_578,N_4580,N_4762);
and UO_579 (O_579,N_4749,N_4748);
and UO_580 (O_580,N_4687,N_4578);
and UO_581 (O_581,N_4663,N_4740);
nand UO_582 (O_582,N_4910,N_4791);
nand UO_583 (O_583,N_4733,N_4727);
nor UO_584 (O_584,N_4716,N_4812);
and UO_585 (O_585,N_4523,N_4945);
and UO_586 (O_586,N_4570,N_4595);
and UO_587 (O_587,N_4912,N_4525);
nor UO_588 (O_588,N_4998,N_4574);
nor UO_589 (O_589,N_4595,N_4690);
and UO_590 (O_590,N_4618,N_4648);
nand UO_591 (O_591,N_4668,N_4531);
nor UO_592 (O_592,N_4743,N_4806);
or UO_593 (O_593,N_4806,N_4994);
nand UO_594 (O_594,N_4718,N_4771);
nor UO_595 (O_595,N_4645,N_4721);
nor UO_596 (O_596,N_4785,N_4938);
nor UO_597 (O_597,N_4866,N_4875);
nand UO_598 (O_598,N_4902,N_4783);
nand UO_599 (O_599,N_4804,N_4756);
or UO_600 (O_600,N_4622,N_4617);
or UO_601 (O_601,N_4944,N_4708);
and UO_602 (O_602,N_4944,N_4881);
nand UO_603 (O_603,N_4880,N_4631);
nor UO_604 (O_604,N_4684,N_4757);
nand UO_605 (O_605,N_4603,N_4991);
nor UO_606 (O_606,N_4633,N_4789);
nor UO_607 (O_607,N_4692,N_4892);
and UO_608 (O_608,N_4700,N_4942);
or UO_609 (O_609,N_4608,N_4901);
and UO_610 (O_610,N_4867,N_4903);
and UO_611 (O_611,N_4827,N_4530);
nand UO_612 (O_612,N_4996,N_4540);
nor UO_613 (O_613,N_4729,N_4907);
and UO_614 (O_614,N_4756,N_4763);
nand UO_615 (O_615,N_4890,N_4996);
and UO_616 (O_616,N_4566,N_4712);
nor UO_617 (O_617,N_4990,N_4869);
nand UO_618 (O_618,N_4820,N_4547);
or UO_619 (O_619,N_4747,N_4976);
or UO_620 (O_620,N_4587,N_4867);
nand UO_621 (O_621,N_4618,N_4866);
or UO_622 (O_622,N_4776,N_4666);
and UO_623 (O_623,N_4953,N_4784);
nand UO_624 (O_624,N_4528,N_4964);
or UO_625 (O_625,N_4913,N_4761);
and UO_626 (O_626,N_4795,N_4583);
xnor UO_627 (O_627,N_4527,N_4599);
and UO_628 (O_628,N_4740,N_4571);
or UO_629 (O_629,N_4705,N_4902);
nand UO_630 (O_630,N_4570,N_4527);
nand UO_631 (O_631,N_4789,N_4894);
and UO_632 (O_632,N_4518,N_4597);
and UO_633 (O_633,N_4639,N_4846);
nand UO_634 (O_634,N_4543,N_4966);
xor UO_635 (O_635,N_4627,N_4838);
or UO_636 (O_636,N_4738,N_4968);
nand UO_637 (O_637,N_4746,N_4776);
nand UO_638 (O_638,N_4931,N_4924);
and UO_639 (O_639,N_4583,N_4974);
nor UO_640 (O_640,N_4795,N_4944);
or UO_641 (O_641,N_4755,N_4913);
or UO_642 (O_642,N_4606,N_4504);
nor UO_643 (O_643,N_4596,N_4778);
or UO_644 (O_644,N_4609,N_4694);
or UO_645 (O_645,N_4721,N_4978);
and UO_646 (O_646,N_4511,N_4572);
or UO_647 (O_647,N_4982,N_4636);
nand UO_648 (O_648,N_4506,N_4937);
nand UO_649 (O_649,N_4575,N_4967);
nor UO_650 (O_650,N_4555,N_4678);
and UO_651 (O_651,N_4616,N_4744);
or UO_652 (O_652,N_4543,N_4699);
nand UO_653 (O_653,N_4840,N_4798);
nor UO_654 (O_654,N_4594,N_4566);
xor UO_655 (O_655,N_4661,N_4797);
or UO_656 (O_656,N_4929,N_4676);
and UO_657 (O_657,N_4567,N_4637);
and UO_658 (O_658,N_4560,N_4575);
nor UO_659 (O_659,N_4788,N_4907);
or UO_660 (O_660,N_4987,N_4687);
nand UO_661 (O_661,N_4987,N_4873);
and UO_662 (O_662,N_4956,N_4553);
and UO_663 (O_663,N_4973,N_4748);
nand UO_664 (O_664,N_4992,N_4823);
or UO_665 (O_665,N_4786,N_4876);
nand UO_666 (O_666,N_4614,N_4764);
nor UO_667 (O_667,N_4852,N_4966);
or UO_668 (O_668,N_4988,N_4509);
xor UO_669 (O_669,N_4674,N_4782);
xnor UO_670 (O_670,N_4989,N_4961);
xor UO_671 (O_671,N_4854,N_4948);
xor UO_672 (O_672,N_4794,N_4710);
or UO_673 (O_673,N_4849,N_4508);
or UO_674 (O_674,N_4923,N_4654);
or UO_675 (O_675,N_4682,N_4974);
and UO_676 (O_676,N_4993,N_4543);
xnor UO_677 (O_677,N_4766,N_4648);
xor UO_678 (O_678,N_4785,N_4506);
and UO_679 (O_679,N_4577,N_4684);
nor UO_680 (O_680,N_4895,N_4528);
nor UO_681 (O_681,N_4927,N_4730);
nand UO_682 (O_682,N_4673,N_4702);
nand UO_683 (O_683,N_4667,N_4535);
nor UO_684 (O_684,N_4870,N_4512);
nand UO_685 (O_685,N_4613,N_4759);
nor UO_686 (O_686,N_4927,N_4744);
or UO_687 (O_687,N_4831,N_4625);
xnor UO_688 (O_688,N_4774,N_4715);
or UO_689 (O_689,N_4668,N_4818);
or UO_690 (O_690,N_4911,N_4894);
or UO_691 (O_691,N_4931,N_4728);
and UO_692 (O_692,N_4940,N_4725);
nor UO_693 (O_693,N_4964,N_4817);
or UO_694 (O_694,N_4941,N_4714);
and UO_695 (O_695,N_4766,N_4889);
nand UO_696 (O_696,N_4700,N_4683);
nor UO_697 (O_697,N_4796,N_4726);
nand UO_698 (O_698,N_4730,N_4836);
and UO_699 (O_699,N_4987,N_4547);
and UO_700 (O_700,N_4758,N_4716);
nor UO_701 (O_701,N_4800,N_4779);
nand UO_702 (O_702,N_4966,N_4730);
nand UO_703 (O_703,N_4822,N_4671);
xnor UO_704 (O_704,N_4874,N_4831);
nand UO_705 (O_705,N_4874,N_4781);
nor UO_706 (O_706,N_4545,N_4633);
nor UO_707 (O_707,N_4592,N_4682);
nor UO_708 (O_708,N_4986,N_4730);
or UO_709 (O_709,N_4903,N_4548);
or UO_710 (O_710,N_4708,N_4994);
and UO_711 (O_711,N_4854,N_4511);
xor UO_712 (O_712,N_4971,N_4819);
or UO_713 (O_713,N_4858,N_4801);
or UO_714 (O_714,N_4910,N_4776);
xor UO_715 (O_715,N_4848,N_4824);
or UO_716 (O_716,N_4700,N_4618);
and UO_717 (O_717,N_4927,N_4812);
or UO_718 (O_718,N_4775,N_4826);
or UO_719 (O_719,N_4709,N_4618);
nor UO_720 (O_720,N_4719,N_4810);
and UO_721 (O_721,N_4510,N_4916);
nand UO_722 (O_722,N_4681,N_4606);
nor UO_723 (O_723,N_4734,N_4519);
nand UO_724 (O_724,N_4963,N_4789);
and UO_725 (O_725,N_4562,N_4983);
nand UO_726 (O_726,N_4997,N_4906);
and UO_727 (O_727,N_4581,N_4860);
and UO_728 (O_728,N_4600,N_4626);
nand UO_729 (O_729,N_4941,N_4820);
or UO_730 (O_730,N_4856,N_4789);
nor UO_731 (O_731,N_4964,N_4771);
nor UO_732 (O_732,N_4712,N_4731);
nor UO_733 (O_733,N_4663,N_4750);
and UO_734 (O_734,N_4546,N_4551);
nand UO_735 (O_735,N_4780,N_4960);
xor UO_736 (O_736,N_4707,N_4830);
nor UO_737 (O_737,N_4687,N_4862);
and UO_738 (O_738,N_4517,N_4609);
nor UO_739 (O_739,N_4504,N_4811);
nand UO_740 (O_740,N_4698,N_4544);
nand UO_741 (O_741,N_4778,N_4920);
and UO_742 (O_742,N_4751,N_4883);
nor UO_743 (O_743,N_4961,N_4756);
xor UO_744 (O_744,N_4712,N_4943);
nand UO_745 (O_745,N_4599,N_4826);
and UO_746 (O_746,N_4778,N_4512);
nor UO_747 (O_747,N_4726,N_4582);
or UO_748 (O_748,N_4702,N_4854);
nand UO_749 (O_749,N_4723,N_4857);
or UO_750 (O_750,N_4817,N_4838);
or UO_751 (O_751,N_4829,N_4587);
or UO_752 (O_752,N_4934,N_4750);
or UO_753 (O_753,N_4816,N_4814);
and UO_754 (O_754,N_4639,N_4757);
nor UO_755 (O_755,N_4512,N_4687);
and UO_756 (O_756,N_4613,N_4871);
and UO_757 (O_757,N_4940,N_4837);
or UO_758 (O_758,N_4705,N_4601);
nand UO_759 (O_759,N_4631,N_4513);
and UO_760 (O_760,N_4750,N_4971);
or UO_761 (O_761,N_4759,N_4937);
nand UO_762 (O_762,N_4527,N_4945);
nor UO_763 (O_763,N_4598,N_4513);
or UO_764 (O_764,N_4982,N_4964);
nand UO_765 (O_765,N_4664,N_4562);
nor UO_766 (O_766,N_4568,N_4599);
xnor UO_767 (O_767,N_4953,N_4859);
nand UO_768 (O_768,N_4978,N_4594);
nor UO_769 (O_769,N_4634,N_4715);
nor UO_770 (O_770,N_4970,N_4628);
or UO_771 (O_771,N_4705,N_4546);
or UO_772 (O_772,N_4919,N_4630);
or UO_773 (O_773,N_4972,N_4532);
nor UO_774 (O_774,N_4915,N_4888);
or UO_775 (O_775,N_4749,N_4586);
nand UO_776 (O_776,N_4878,N_4985);
or UO_777 (O_777,N_4632,N_4995);
or UO_778 (O_778,N_4871,N_4693);
nor UO_779 (O_779,N_4810,N_4750);
or UO_780 (O_780,N_4732,N_4859);
nand UO_781 (O_781,N_4500,N_4739);
and UO_782 (O_782,N_4840,N_4935);
nor UO_783 (O_783,N_4575,N_4665);
or UO_784 (O_784,N_4718,N_4829);
or UO_785 (O_785,N_4947,N_4844);
nand UO_786 (O_786,N_4913,N_4559);
and UO_787 (O_787,N_4569,N_4939);
xnor UO_788 (O_788,N_4647,N_4892);
or UO_789 (O_789,N_4910,N_4547);
nand UO_790 (O_790,N_4864,N_4573);
nor UO_791 (O_791,N_4895,N_4991);
or UO_792 (O_792,N_4520,N_4885);
nor UO_793 (O_793,N_4595,N_4992);
nand UO_794 (O_794,N_4776,N_4809);
and UO_795 (O_795,N_4583,N_4783);
and UO_796 (O_796,N_4629,N_4708);
and UO_797 (O_797,N_4755,N_4732);
or UO_798 (O_798,N_4616,N_4778);
and UO_799 (O_799,N_4548,N_4864);
nand UO_800 (O_800,N_4582,N_4908);
nor UO_801 (O_801,N_4961,N_4822);
nor UO_802 (O_802,N_4716,N_4615);
nand UO_803 (O_803,N_4650,N_4954);
xor UO_804 (O_804,N_4681,N_4927);
xor UO_805 (O_805,N_4818,N_4862);
or UO_806 (O_806,N_4926,N_4504);
or UO_807 (O_807,N_4545,N_4601);
or UO_808 (O_808,N_4865,N_4883);
and UO_809 (O_809,N_4948,N_4635);
nand UO_810 (O_810,N_4553,N_4679);
and UO_811 (O_811,N_4893,N_4670);
nand UO_812 (O_812,N_4613,N_4594);
nor UO_813 (O_813,N_4782,N_4813);
or UO_814 (O_814,N_4995,N_4913);
and UO_815 (O_815,N_4508,N_4676);
or UO_816 (O_816,N_4718,N_4850);
or UO_817 (O_817,N_4971,N_4660);
or UO_818 (O_818,N_4819,N_4771);
nand UO_819 (O_819,N_4784,N_4617);
nand UO_820 (O_820,N_4599,N_4950);
nand UO_821 (O_821,N_4886,N_4711);
or UO_822 (O_822,N_4548,N_4936);
and UO_823 (O_823,N_4857,N_4876);
nor UO_824 (O_824,N_4866,N_4625);
and UO_825 (O_825,N_4724,N_4646);
or UO_826 (O_826,N_4927,N_4591);
or UO_827 (O_827,N_4746,N_4887);
and UO_828 (O_828,N_4991,N_4990);
xor UO_829 (O_829,N_4780,N_4853);
and UO_830 (O_830,N_4810,N_4966);
nor UO_831 (O_831,N_4599,N_4549);
and UO_832 (O_832,N_4941,N_4630);
and UO_833 (O_833,N_4575,N_4519);
or UO_834 (O_834,N_4588,N_4502);
nand UO_835 (O_835,N_4671,N_4998);
or UO_836 (O_836,N_4786,N_4718);
and UO_837 (O_837,N_4513,N_4671);
and UO_838 (O_838,N_4913,N_4871);
xnor UO_839 (O_839,N_4921,N_4806);
nand UO_840 (O_840,N_4899,N_4532);
nand UO_841 (O_841,N_4755,N_4652);
or UO_842 (O_842,N_4993,N_4601);
or UO_843 (O_843,N_4920,N_4978);
nor UO_844 (O_844,N_4847,N_4790);
and UO_845 (O_845,N_4712,N_4638);
or UO_846 (O_846,N_4628,N_4616);
or UO_847 (O_847,N_4789,N_4565);
or UO_848 (O_848,N_4535,N_4814);
or UO_849 (O_849,N_4634,N_4998);
or UO_850 (O_850,N_4525,N_4955);
nor UO_851 (O_851,N_4768,N_4971);
nand UO_852 (O_852,N_4613,N_4774);
nor UO_853 (O_853,N_4647,N_4777);
or UO_854 (O_854,N_4702,N_4695);
nand UO_855 (O_855,N_4751,N_4753);
nand UO_856 (O_856,N_4768,N_4847);
nand UO_857 (O_857,N_4712,N_4887);
and UO_858 (O_858,N_4773,N_4579);
nand UO_859 (O_859,N_4982,N_4586);
nor UO_860 (O_860,N_4807,N_4866);
xnor UO_861 (O_861,N_4826,N_4901);
nor UO_862 (O_862,N_4509,N_4567);
nand UO_863 (O_863,N_4985,N_4989);
and UO_864 (O_864,N_4878,N_4544);
or UO_865 (O_865,N_4698,N_4587);
xnor UO_866 (O_866,N_4977,N_4752);
nor UO_867 (O_867,N_4870,N_4522);
nand UO_868 (O_868,N_4975,N_4627);
or UO_869 (O_869,N_4760,N_4766);
nand UO_870 (O_870,N_4568,N_4531);
nand UO_871 (O_871,N_4545,N_4514);
and UO_872 (O_872,N_4993,N_4797);
and UO_873 (O_873,N_4688,N_4872);
nor UO_874 (O_874,N_4922,N_4505);
nand UO_875 (O_875,N_4715,N_4927);
nor UO_876 (O_876,N_4864,N_4574);
xor UO_877 (O_877,N_4586,N_4933);
nand UO_878 (O_878,N_4766,N_4518);
and UO_879 (O_879,N_4590,N_4743);
or UO_880 (O_880,N_4852,N_4748);
or UO_881 (O_881,N_4982,N_4510);
and UO_882 (O_882,N_4643,N_4653);
or UO_883 (O_883,N_4922,N_4958);
nor UO_884 (O_884,N_4985,N_4923);
or UO_885 (O_885,N_4557,N_4927);
or UO_886 (O_886,N_4945,N_4742);
or UO_887 (O_887,N_4772,N_4595);
and UO_888 (O_888,N_4577,N_4898);
or UO_889 (O_889,N_4896,N_4750);
or UO_890 (O_890,N_4571,N_4760);
or UO_891 (O_891,N_4935,N_4752);
and UO_892 (O_892,N_4961,N_4962);
xnor UO_893 (O_893,N_4529,N_4651);
nand UO_894 (O_894,N_4615,N_4979);
or UO_895 (O_895,N_4998,N_4788);
and UO_896 (O_896,N_4629,N_4598);
nor UO_897 (O_897,N_4743,N_4603);
or UO_898 (O_898,N_4585,N_4923);
and UO_899 (O_899,N_4694,N_4598);
or UO_900 (O_900,N_4831,N_4547);
nor UO_901 (O_901,N_4614,N_4892);
or UO_902 (O_902,N_4520,N_4645);
nand UO_903 (O_903,N_4776,N_4860);
and UO_904 (O_904,N_4621,N_4870);
xor UO_905 (O_905,N_4926,N_4950);
and UO_906 (O_906,N_4552,N_4841);
nand UO_907 (O_907,N_4691,N_4563);
or UO_908 (O_908,N_4607,N_4639);
nor UO_909 (O_909,N_4695,N_4755);
or UO_910 (O_910,N_4959,N_4569);
nor UO_911 (O_911,N_4716,N_4879);
and UO_912 (O_912,N_4978,N_4888);
or UO_913 (O_913,N_4814,N_4616);
nand UO_914 (O_914,N_4985,N_4836);
nor UO_915 (O_915,N_4791,N_4921);
and UO_916 (O_916,N_4559,N_4645);
or UO_917 (O_917,N_4794,N_4540);
or UO_918 (O_918,N_4787,N_4528);
or UO_919 (O_919,N_4637,N_4638);
nor UO_920 (O_920,N_4970,N_4511);
nor UO_921 (O_921,N_4972,N_4656);
and UO_922 (O_922,N_4784,N_4922);
or UO_923 (O_923,N_4537,N_4953);
nand UO_924 (O_924,N_4904,N_4976);
nor UO_925 (O_925,N_4893,N_4632);
and UO_926 (O_926,N_4897,N_4719);
nor UO_927 (O_927,N_4622,N_4852);
or UO_928 (O_928,N_4960,N_4930);
nand UO_929 (O_929,N_4669,N_4586);
or UO_930 (O_930,N_4899,N_4859);
nand UO_931 (O_931,N_4756,N_4760);
nand UO_932 (O_932,N_4991,N_4651);
nor UO_933 (O_933,N_4590,N_4790);
nand UO_934 (O_934,N_4694,N_4624);
or UO_935 (O_935,N_4553,N_4797);
nor UO_936 (O_936,N_4659,N_4887);
nand UO_937 (O_937,N_4707,N_4814);
nor UO_938 (O_938,N_4527,N_4667);
or UO_939 (O_939,N_4757,N_4836);
nand UO_940 (O_940,N_4893,N_4991);
nand UO_941 (O_941,N_4596,N_4569);
nand UO_942 (O_942,N_4783,N_4691);
xnor UO_943 (O_943,N_4977,N_4973);
and UO_944 (O_944,N_4818,N_4662);
or UO_945 (O_945,N_4884,N_4878);
or UO_946 (O_946,N_4939,N_4533);
nand UO_947 (O_947,N_4765,N_4565);
or UO_948 (O_948,N_4776,N_4641);
nor UO_949 (O_949,N_4683,N_4754);
nor UO_950 (O_950,N_4562,N_4524);
nor UO_951 (O_951,N_4539,N_4822);
nor UO_952 (O_952,N_4967,N_4641);
and UO_953 (O_953,N_4824,N_4631);
and UO_954 (O_954,N_4832,N_4720);
nand UO_955 (O_955,N_4972,N_4919);
and UO_956 (O_956,N_4914,N_4643);
nor UO_957 (O_957,N_4979,N_4652);
nand UO_958 (O_958,N_4915,N_4668);
nand UO_959 (O_959,N_4504,N_4576);
and UO_960 (O_960,N_4992,N_4901);
nand UO_961 (O_961,N_4633,N_4975);
or UO_962 (O_962,N_4600,N_4688);
nand UO_963 (O_963,N_4537,N_4606);
nand UO_964 (O_964,N_4963,N_4511);
nand UO_965 (O_965,N_4945,N_4942);
nor UO_966 (O_966,N_4821,N_4589);
nor UO_967 (O_967,N_4796,N_4713);
xor UO_968 (O_968,N_4993,N_4903);
and UO_969 (O_969,N_4733,N_4942);
or UO_970 (O_970,N_4666,N_4900);
or UO_971 (O_971,N_4871,N_4514);
nor UO_972 (O_972,N_4813,N_4988);
xnor UO_973 (O_973,N_4916,N_4811);
and UO_974 (O_974,N_4776,N_4833);
nand UO_975 (O_975,N_4756,N_4548);
xnor UO_976 (O_976,N_4910,N_4681);
or UO_977 (O_977,N_4737,N_4989);
nand UO_978 (O_978,N_4912,N_4719);
and UO_979 (O_979,N_4635,N_4977);
nor UO_980 (O_980,N_4519,N_4708);
or UO_981 (O_981,N_4513,N_4889);
and UO_982 (O_982,N_4581,N_4601);
nand UO_983 (O_983,N_4903,N_4593);
nor UO_984 (O_984,N_4649,N_4819);
nand UO_985 (O_985,N_4620,N_4646);
or UO_986 (O_986,N_4582,N_4881);
nor UO_987 (O_987,N_4521,N_4754);
and UO_988 (O_988,N_4939,N_4523);
and UO_989 (O_989,N_4622,N_4591);
or UO_990 (O_990,N_4739,N_4769);
nand UO_991 (O_991,N_4510,N_4978);
and UO_992 (O_992,N_4769,N_4944);
nand UO_993 (O_993,N_4908,N_4621);
nand UO_994 (O_994,N_4931,N_4737);
and UO_995 (O_995,N_4970,N_4671);
nand UO_996 (O_996,N_4642,N_4664);
or UO_997 (O_997,N_4821,N_4702);
and UO_998 (O_998,N_4934,N_4545);
xnor UO_999 (O_999,N_4591,N_4677);
endmodule