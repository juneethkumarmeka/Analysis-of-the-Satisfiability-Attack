module basic_3000_30000_3500_20_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xor U0 (N_0,In_1726,In_876);
or U1 (N_1,In_1662,In_312);
xor U2 (N_2,In_1260,In_2676);
or U3 (N_3,In_2983,In_348);
nor U4 (N_4,In_2767,In_654);
xnor U5 (N_5,In_809,In_320);
and U6 (N_6,In_111,In_986);
and U7 (N_7,In_2683,In_2777);
xor U8 (N_8,In_1424,In_656);
nor U9 (N_9,In_881,In_2422);
nand U10 (N_10,In_1645,In_406);
or U11 (N_11,In_1030,In_2055);
xnor U12 (N_12,In_15,In_921);
xnor U13 (N_13,In_302,In_2465);
nand U14 (N_14,In_2090,In_1602);
and U15 (N_15,In_509,In_1788);
nand U16 (N_16,In_1512,In_2730);
xor U17 (N_17,In_698,In_559);
nor U18 (N_18,In_2343,In_2474);
nand U19 (N_19,In_431,In_2353);
and U20 (N_20,In_2540,In_27);
nor U21 (N_21,In_2697,In_2802);
nor U22 (N_22,In_379,In_1163);
nand U23 (N_23,In_2723,In_2989);
or U24 (N_24,In_1672,In_1896);
xor U25 (N_25,In_1061,In_361);
and U26 (N_26,In_1080,In_232);
nor U27 (N_27,In_852,In_1529);
xnor U28 (N_28,In_2986,In_2965);
or U29 (N_29,In_1173,In_1296);
nor U30 (N_30,In_1203,In_1874);
nand U31 (N_31,In_1263,In_2398);
and U32 (N_32,In_2503,In_2307);
and U33 (N_33,In_1346,In_86);
xor U34 (N_34,In_204,In_1687);
or U35 (N_35,In_249,In_1640);
and U36 (N_36,In_2289,In_223);
xor U37 (N_37,In_1057,In_1458);
xnor U38 (N_38,In_1714,In_554);
nand U39 (N_39,In_340,In_453);
xnor U40 (N_40,In_2991,In_1850);
nand U41 (N_41,In_2929,In_1973);
or U42 (N_42,In_888,In_478);
nor U43 (N_43,In_471,In_2102);
or U44 (N_44,In_1735,In_1913);
nand U45 (N_45,In_1768,In_1219);
xnor U46 (N_46,In_1097,In_893);
or U47 (N_47,In_141,In_2955);
nor U48 (N_48,In_2587,In_1832);
and U49 (N_49,In_1810,In_1326);
or U50 (N_50,In_129,In_2043);
xor U51 (N_51,In_174,In_2733);
nand U52 (N_52,In_1885,In_1237);
or U53 (N_53,In_2606,In_208);
and U54 (N_54,In_1839,In_1377);
and U55 (N_55,In_1270,In_1613);
xor U56 (N_56,In_507,In_1649);
xor U57 (N_57,In_2221,In_60);
or U58 (N_58,In_1635,In_868);
and U59 (N_59,In_607,In_1927);
nor U60 (N_60,In_952,In_518);
and U61 (N_61,In_1309,In_828);
nor U62 (N_62,In_1993,In_1611);
nor U63 (N_63,In_1781,In_2338);
nand U64 (N_64,In_2210,In_1794);
or U65 (N_65,In_2708,In_910);
nand U66 (N_66,In_2957,In_814);
nand U67 (N_67,In_1146,In_1614);
xnor U68 (N_68,In_551,In_874);
nand U69 (N_69,In_878,In_1158);
xor U70 (N_70,In_2887,In_1950);
nor U71 (N_71,In_100,In_2011);
xor U72 (N_72,In_1582,In_19);
or U73 (N_73,In_836,In_286);
and U74 (N_74,In_1289,In_900);
and U75 (N_75,In_366,In_711);
and U76 (N_76,In_310,In_1990);
xnor U77 (N_77,In_1059,In_822);
and U78 (N_78,In_190,In_2317);
or U79 (N_79,In_1807,In_109);
nor U80 (N_80,In_1510,In_132);
or U81 (N_81,In_1359,In_1052);
nand U82 (N_82,In_2114,In_84);
xnor U83 (N_83,In_964,In_1757);
nand U84 (N_84,In_1100,In_244);
xnor U85 (N_85,In_1713,In_2638);
and U86 (N_86,In_2452,In_501);
nor U87 (N_87,In_218,In_2566);
nor U88 (N_88,In_2926,In_1908);
or U89 (N_89,In_1540,In_181);
xnor U90 (N_90,In_2621,In_466);
nor U91 (N_91,In_323,In_2345);
xnor U92 (N_92,In_2180,In_265);
xor U93 (N_93,In_2968,In_1127);
and U94 (N_94,In_2260,In_1945);
and U95 (N_95,In_520,In_603);
nand U96 (N_96,In_1669,In_2899);
or U97 (N_97,In_942,In_1437);
or U98 (N_98,In_1806,In_2877);
xor U99 (N_99,In_527,In_301);
and U100 (N_100,In_2967,In_401);
xnor U101 (N_101,In_1084,In_2168);
or U102 (N_102,In_2220,In_679);
nor U103 (N_103,In_1200,In_1895);
or U104 (N_104,In_2495,In_623);
and U105 (N_105,In_395,In_572);
and U106 (N_106,In_760,In_1330);
xor U107 (N_107,In_1415,In_185);
nand U108 (N_108,In_1778,In_219);
nor U109 (N_109,In_975,In_782);
and U110 (N_110,In_1016,In_1968);
or U111 (N_111,In_2809,In_290);
nand U112 (N_112,In_1380,In_1678);
or U113 (N_113,In_2272,In_897);
or U114 (N_114,In_2848,In_1058);
nand U115 (N_115,In_1293,In_2882);
nand U116 (N_116,In_1533,In_176);
xor U117 (N_117,In_1576,In_544);
or U118 (N_118,In_1638,In_678);
and U119 (N_119,In_2753,In_30);
or U120 (N_120,In_745,In_552);
nand U121 (N_121,In_2508,In_1783);
nand U122 (N_122,In_69,In_1666);
nor U123 (N_123,In_1846,In_967);
nor U124 (N_124,In_2805,In_2065);
and U125 (N_125,In_2223,In_2513);
or U126 (N_126,In_1835,In_2254);
or U127 (N_127,In_414,In_2575);
xnor U128 (N_128,In_843,In_2190);
xnor U129 (N_129,In_2105,In_1621);
or U130 (N_130,In_1107,In_2379);
xor U131 (N_131,In_2564,In_925);
and U132 (N_132,In_2,In_410);
xor U133 (N_133,In_884,In_2467);
xor U134 (N_134,In_1776,In_2793);
nor U135 (N_135,In_2117,In_2921);
and U136 (N_136,In_765,In_546);
or U137 (N_137,In_2685,In_1563);
xor U138 (N_138,In_1938,In_1287);
xnor U139 (N_139,In_2814,In_1720);
nand U140 (N_140,In_1954,In_863);
or U141 (N_141,In_1251,In_2479);
or U142 (N_142,In_1855,In_251);
nand U143 (N_143,In_2721,In_2484);
nand U144 (N_144,In_1502,In_439);
nand U145 (N_145,In_2433,In_1024);
or U146 (N_146,In_1763,In_1965);
or U147 (N_147,In_1890,In_105);
nand U148 (N_148,In_1786,In_405);
or U149 (N_149,In_2292,In_432);
and U150 (N_150,In_2501,In_2219);
and U151 (N_151,In_1241,In_2532);
and U152 (N_152,In_1709,In_1356);
nand U153 (N_153,In_2021,In_1811);
nand U154 (N_154,In_1619,In_1469);
nand U155 (N_155,In_2731,In_160);
or U156 (N_156,In_1,In_2625);
and U157 (N_157,In_1616,In_1964);
nor U158 (N_158,In_2373,In_331);
and U159 (N_159,In_421,In_1281);
nor U160 (N_160,In_2188,In_832);
and U161 (N_161,In_1012,In_2537);
xnor U162 (N_162,In_2722,In_5);
nor U163 (N_163,In_1347,In_1498);
or U164 (N_164,In_52,In_602);
or U165 (N_165,In_1490,In_350);
nor U166 (N_166,In_1608,In_450);
nor U167 (N_167,In_508,In_1985);
xor U168 (N_168,In_1223,In_1104);
xor U169 (N_169,In_1130,In_2987);
nor U170 (N_170,In_926,In_169);
or U171 (N_171,In_1530,In_1474);
nand U172 (N_172,In_1836,In_152);
nor U173 (N_173,In_2944,In_1343);
nand U174 (N_174,In_2772,In_2547);
and U175 (N_175,In_474,In_2185);
or U176 (N_176,In_177,In_709);
xor U177 (N_177,In_1658,In_124);
xor U178 (N_178,In_2523,In_962);
and U179 (N_179,In_1489,In_1142);
nor U180 (N_180,In_461,In_2620);
nor U181 (N_181,In_1421,In_1222);
or U182 (N_182,In_1331,In_1144);
or U183 (N_183,In_248,In_1789);
xnor U184 (N_184,In_862,In_2486);
nor U185 (N_185,In_110,In_1884);
nor U186 (N_186,In_2633,In_2029);
and U187 (N_187,In_1006,In_598);
nor U188 (N_188,In_2641,In_2137);
nand U189 (N_189,In_2655,In_1160);
xnor U190 (N_190,In_212,In_791);
and U191 (N_191,In_1700,In_237);
nor U192 (N_192,In_1204,In_2992);
xnor U193 (N_193,In_2569,In_1093);
or U194 (N_194,In_2982,In_1663);
nor U195 (N_195,In_1949,In_1361);
nand U196 (N_196,In_2573,In_1573);
and U197 (N_197,In_1198,In_1842);
nor U198 (N_198,In_779,In_2781);
nand U199 (N_199,In_2460,In_708);
xnor U200 (N_200,In_2250,In_1169);
xor U201 (N_201,In_1370,In_752);
nor U202 (N_202,In_2834,In_699);
xnor U203 (N_203,In_1476,In_2860);
nor U204 (N_204,In_161,In_877);
and U205 (N_205,In_1499,In_903);
or U206 (N_206,In_1918,In_247);
nor U207 (N_207,In_2082,In_1017);
and U208 (N_208,In_400,In_269);
nand U209 (N_209,In_1622,In_2170);
nand U210 (N_210,In_2384,In_492);
nand U211 (N_211,In_590,In_264);
nor U212 (N_212,In_2096,In_1865);
nand U213 (N_213,In_948,In_436);
nand U214 (N_214,In_1053,In_1860);
nor U215 (N_215,In_1724,In_1979);
or U216 (N_216,In_1324,In_781);
nor U217 (N_217,In_1590,In_1078);
nand U218 (N_218,In_104,In_2365);
nand U219 (N_219,In_2006,In_992);
xor U220 (N_220,In_716,In_2959);
or U221 (N_221,In_1984,In_1322);
or U222 (N_222,In_2928,In_2129);
xnor U223 (N_223,In_337,In_1238);
and U224 (N_224,In_1653,In_275);
nand U225 (N_225,In_719,In_45);
or U226 (N_226,In_543,In_2195);
nand U227 (N_227,In_445,In_1577);
xor U228 (N_228,In_2897,In_1862);
xor U229 (N_229,In_305,In_1384);
and U230 (N_230,In_1205,In_2439);
and U231 (N_231,In_1420,In_2426);
nor U232 (N_232,In_506,In_575);
nor U233 (N_233,In_1725,In_1802);
or U234 (N_234,In_1628,In_1193);
or U235 (N_235,In_2825,In_2327);
and U236 (N_236,In_1126,In_2498);
nand U237 (N_237,In_2522,In_2624);
and U238 (N_238,In_615,In_2925);
or U239 (N_239,In_2788,In_963);
or U240 (N_240,In_61,In_123);
and U241 (N_241,In_2693,In_1961);
xnor U242 (N_242,In_2280,In_179);
nor U243 (N_243,In_1302,In_2357);
nand U244 (N_244,In_23,In_2387);
xor U245 (N_245,In_1374,In_12);
nand U246 (N_246,In_887,In_451);
nand U247 (N_247,In_135,In_2064);
or U248 (N_248,In_867,In_1026);
nor U249 (N_249,In_2405,In_1011);
or U250 (N_250,In_335,In_2397);
nand U251 (N_251,In_734,In_1857);
nor U252 (N_252,In_1069,In_1681);
xnor U253 (N_253,In_2165,In_1412);
xnor U254 (N_254,In_2670,In_2425);
nor U255 (N_255,In_566,In_2700);
and U256 (N_256,In_270,In_996);
xor U257 (N_257,In_2391,In_2674);
and U258 (N_258,In_180,In_1101);
nand U259 (N_259,In_2962,In_142);
nand U260 (N_260,In_1243,In_2661);
or U261 (N_261,In_776,In_936);
nand U262 (N_262,In_786,In_49);
nand U263 (N_263,In_2164,In_2702);
and U264 (N_264,In_2632,In_1817);
or U265 (N_265,In_701,In_2432);
nor U266 (N_266,In_458,In_1851);
and U267 (N_267,In_1680,In_1718);
nor U268 (N_268,In_2778,In_1830);
or U269 (N_269,In_1418,In_2418);
xor U270 (N_270,In_2110,In_1209);
nor U271 (N_271,In_594,In_2489);
nor U272 (N_272,In_668,In_1821);
xor U273 (N_273,In_2530,In_1320);
nor U274 (N_274,In_2429,In_829);
nor U275 (N_275,In_2823,In_1741);
xor U276 (N_276,In_844,In_1098);
and U277 (N_277,In_1578,In_1685);
nand U278 (N_278,In_1362,In_642);
nor U279 (N_279,In_2888,In_7);
xnor U280 (N_280,In_1038,In_1737);
nand U281 (N_281,In_1014,In_1937);
nand U282 (N_282,In_2504,In_263);
and U283 (N_283,In_589,In_2466);
nand U284 (N_284,In_2716,In_2647);
and U285 (N_285,In_1196,In_1917);
nand U286 (N_286,In_1230,In_2868);
nor U287 (N_287,In_799,In_1004);
nor U288 (N_288,In_523,In_1808);
nand U289 (N_289,In_2181,In_2175);
or U290 (N_290,In_899,In_2815);
xor U291 (N_291,In_1552,In_655);
nand U292 (N_292,In_847,In_2301);
nor U293 (N_293,In_1096,In_1119);
nand U294 (N_294,In_2966,In_2551);
xor U295 (N_295,In_1642,In_2328);
or U296 (N_296,In_1081,In_2738);
xnor U297 (N_297,In_2324,In_1708);
and U298 (N_298,In_1716,In_2146);
nand U299 (N_299,In_1704,In_404);
and U300 (N_300,In_1756,In_2619);
nand U301 (N_301,In_1790,In_2883);
xnor U302 (N_302,In_1513,In_1639);
xor U303 (N_303,In_120,In_1463);
or U304 (N_304,In_83,In_1934);
nand U305 (N_305,In_1800,In_1935);
or U306 (N_306,In_1311,In_2054);
and U307 (N_307,In_660,In_1166);
xor U308 (N_308,In_2889,In_487);
nand U309 (N_309,In_1665,In_556);
and U310 (N_310,In_2917,In_1515);
xnor U311 (N_311,In_833,In_1447);
and U312 (N_312,In_2818,In_483);
and U313 (N_313,In_1315,In_665);
xnor U314 (N_314,In_1020,In_1581);
and U315 (N_315,In_725,In_262);
and U316 (N_316,In_2378,In_363);
xnor U317 (N_317,In_1446,In_2933);
nand U318 (N_318,In_1803,In_2895);
or U319 (N_319,In_1702,In_412);
or U320 (N_320,In_2013,In_2584);
nor U321 (N_321,In_1998,In_2476);
nand U322 (N_322,In_502,In_637);
or U323 (N_323,In_1272,In_170);
nand U324 (N_324,In_2790,In_1395);
xnor U325 (N_325,In_664,In_297);
nor U326 (N_326,In_1240,In_1580);
xnor U327 (N_327,In_1970,In_2711);
and U328 (N_328,In_1345,In_2213);
or U329 (N_329,In_2320,In_256);
and U330 (N_330,In_2482,In_6);
and U331 (N_331,In_1609,In_2688);
nor U332 (N_332,In_2276,In_2281);
nor U333 (N_333,In_236,In_976);
and U334 (N_334,In_224,In_2845);
and U335 (N_335,In_1723,In_1487);
and U336 (N_336,In_606,In_754);
nand U337 (N_337,In_902,In_1245);
and U338 (N_338,In_1328,In_207);
xnor U339 (N_339,In_2060,In_1133);
nor U340 (N_340,In_226,In_672);
nand U341 (N_341,In_78,In_424);
nor U342 (N_342,In_1542,In_1083);
nor U343 (N_343,In_2528,In_1450);
xnor U344 (N_344,In_2867,In_2668);
nor U345 (N_345,In_1605,In_2994);
and U346 (N_346,In_2545,In_54);
xor U347 (N_347,In_1686,In_1536);
nor U348 (N_348,In_106,In_81);
or U349 (N_349,In_2509,In_2659);
nor U350 (N_350,In_333,In_2245);
and U351 (N_351,In_1001,In_2463);
and U352 (N_352,In_21,In_429);
and U353 (N_353,In_2812,In_2806);
nor U354 (N_354,In_1389,In_1792);
or U355 (N_355,In_2710,In_629);
or U356 (N_356,In_998,In_2757);
nand U357 (N_357,In_1094,In_1439);
xor U358 (N_358,In_2159,In_221);
or U359 (N_359,In_2748,In_2235);
nor U360 (N_360,In_562,In_553);
or U361 (N_361,In_1106,In_338);
nand U362 (N_362,In_1145,In_500);
xnor U363 (N_363,In_2061,In_2240);
or U364 (N_364,In_1115,In_2562);
and U365 (N_365,In_669,In_661);
or U366 (N_366,In_316,In_1462);
or U367 (N_367,In_582,In_1049);
or U368 (N_368,In_751,In_1572);
nor U369 (N_369,In_2207,In_2949);
or U370 (N_370,In_383,In_1300);
or U371 (N_371,In_1777,In_772);
nand U372 (N_372,In_2972,In_8);
and U373 (N_373,In_1838,In_1551);
and U374 (N_374,In_1199,In_2714);
nand U375 (N_375,In_2187,In_2843);
xor U376 (N_376,In_804,In_1693);
nor U377 (N_377,In_2340,In_666);
or U378 (N_378,In_1190,In_417);
nand U379 (N_379,In_2461,In_2577);
or U380 (N_380,In_724,In_20);
nand U381 (N_381,In_2667,In_1348);
and U382 (N_382,In_1863,In_1336);
nor U383 (N_383,In_1305,In_1618);
xnor U384 (N_384,In_524,In_2939);
and U385 (N_385,In_1705,In_260);
and U386 (N_386,In_1535,In_358);
xnor U387 (N_387,In_2924,In_614);
and U388 (N_388,In_1671,In_522);
and U389 (N_389,In_367,In_2666);
and U390 (N_390,In_1232,In_210);
nand U391 (N_391,In_1906,In_9);
nand U392 (N_392,In_1381,In_706);
xor U393 (N_393,In_1943,In_1912);
xnor U394 (N_394,In_596,In_851);
nand U395 (N_395,In_567,In_755);
nor U396 (N_396,In_1344,In_1285);
or U397 (N_397,In_209,In_2517);
and U398 (N_398,In_446,In_1910);
or U399 (N_399,In_2097,In_2367);
or U400 (N_400,In_1769,In_2447);
nor U401 (N_401,In_1698,In_2769);
xor U402 (N_402,In_2300,In_2763);
nand U403 (N_403,In_441,In_2483);
or U404 (N_404,In_1654,In_2464);
xor U405 (N_405,In_1556,In_1545);
nor U406 (N_406,In_610,In_139);
or U407 (N_407,In_2645,In_935);
nor U408 (N_408,In_1400,In_788);
xor U409 (N_409,In_29,In_1135);
nor U410 (N_410,In_1755,In_1168);
and U411 (N_411,In_1939,In_1368);
nor U412 (N_412,In_714,In_416);
nor U413 (N_413,In_2937,In_56);
xnor U414 (N_414,In_1335,In_532);
nor U415 (N_415,In_1366,In_1744);
nand U416 (N_416,In_1460,In_2617);
xnor U417 (N_417,In_908,In_736);
nor U418 (N_418,In_2291,In_2214);
and U419 (N_419,In_2256,In_1889);
nand U420 (N_420,In_274,In_749);
nor U421 (N_421,In_2492,In_703);
or U422 (N_422,In_2408,In_440);
or U423 (N_423,In_2368,In_2381);
and U424 (N_424,In_46,In_1275);
nor U425 (N_425,In_1172,In_1592);
xor U426 (N_426,In_2342,In_1997);
xor U427 (N_427,In_368,In_2016);
and U428 (N_428,In_2960,In_1712);
and U429 (N_429,In_2457,In_1604);
and U430 (N_430,In_1468,In_115);
or U431 (N_431,In_2827,In_1966);
or U432 (N_432,In_960,In_2001);
and U433 (N_433,In_2283,In_2062);
nand U434 (N_434,In_2971,In_2838);
and U435 (N_435,In_1449,In_993);
and U436 (N_436,In_2411,In_894);
nor U437 (N_437,In_2487,In_1833);
nand U438 (N_438,In_676,In_3);
nor U439 (N_439,In_1246,In_2184);
and U440 (N_440,In_1254,In_972);
nand U441 (N_441,In_341,In_980);
and U442 (N_442,In_381,In_1995);
nand U443 (N_443,In_2791,In_1719);
nand U444 (N_444,In_1774,In_1824);
and U445 (N_445,In_1153,In_1554);
or U446 (N_446,In_1559,In_1683);
nand U447 (N_447,In_1508,In_1099);
nor U448 (N_448,In_1549,In_1957);
nor U449 (N_449,In_382,In_1956);
and U450 (N_450,In_744,In_392);
and U451 (N_451,In_327,In_770);
or U452 (N_452,In_2125,In_842);
xnor U453 (N_453,In_682,In_1295);
or U454 (N_454,In_1282,In_1548);
nand U455 (N_455,In_1866,In_2347);
xnor U456 (N_456,In_2161,In_2401);
xnor U457 (N_457,In_2236,In_2735);
or U458 (N_458,In_1433,In_1387);
xnor U459 (N_459,In_1286,In_2525);
nor U460 (N_460,In_2747,In_2000);
xor U461 (N_461,In_1027,In_757);
nand U462 (N_462,In_1747,In_1044);
nor U463 (N_463,In_2796,In_2784);
nor U464 (N_464,In_2511,In_2044);
nand U465 (N_465,In_4,In_59);
nor U466 (N_466,In_1248,In_2063);
and U467 (N_467,In_717,In_1841);
nor U468 (N_468,In_2996,In_339);
nand U469 (N_469,In_2396,In_1070);
nand U470 (N_470,In_88,In_947);
nor U471 (N_471,In_2153,In_1626);
xnor U472 (N_472,In_2247,In_239);
and U473 (N_473,In_1459,In_2650);
and U474 (N_474,In_155,In_677);
nand U475 (N_475,In_2643,In_2741);
xor U476 (N_476,In_748,In_2973);
nor U477 (N_477,In_2521,In_838);
nand U478 (N_478,In_206,In_922);
nor U479 (N_479,In_138,In_396);
and U480 (N_480,In_2568,In_1929);
xnor U481 (N_481,In_2028,In_1480);
xor U482 (N_482,In_896,In_920);
or U483 (N_483,In_2576,In_229);
and U484 (N_484,In_634,In_1488);
xor U485 (N_485,In_2417,In_145);
nand U486 (N_486,In_2045,In_1699);
or U487 (N_487,In_2449,In_2718);
and U488 (N_488,In_1138,In_2085);
xnor U489 (N_489,In_203,In_1541);
xnor U490 (N_490,In_1211,In_192);
nor U491 (N_491,In_486,In_1073);
and U492 (N_492,In_600,In_571);
xor U493 (N_493,In_1603,In_2556);
or U494 (N_494,In_673,In_243);
and U495 (N_495,In_1484,In_1294);
and U496 (N_496,In_2392,In_2206);
or U497 (N_497,In_2154,In_2631);
or U498 (N_498,In_2360,In_497);
or U499 (N_499,In_435,In_101);
xor U500 (N_500,In_2279,In_1509);
or U501 (N_501,In_2896,In_773);
nand U502 (N_502,In_1063,In_1749);
nand U503 (N_503,In_2414,In_621);
xor U504 (N_504,In_1967,In_1583);
xor U505 (N_505,In_2009,In_73);
or U506 (N_506,In_2369,In_618);
nor U507 (N_507,In_318,In_2049);
nand U508 (N_508,In_2371,In_489);
and U509 (N_509,In_252,In_22);
xnor U510 (N_510,In_907,In_419);
xnor U511 (N_511,In_2592,In_173);
or U512 (N_512,In_2076,In_1338);
nor U513 (N_513,In_1132,In_2174);
xnor U514 (N_514,In_2402,In_1202);
xnor U515 (N_515,In_775,In_2069);
nand U516 (N_516,In_2040,In_28);
or U517 (N_517,In_1743,In_126);
and U518 (N_518,In_1497,In_730);
or U519 (N_519,In_299,In_2956);
or U520 (N_520,In_369,In_2329);
or U521 (N_521,In_1148,In_1731);
xor U522 (N_522,In_1175,In_1431);
nor U523 (N_523,In_2073,In_742);
nand U524 (N_524,In_1538,In_2554);
nor U525 (N_525,In_2998,In_2286);
xor U526 (N_526,In_783,In_2828);
xnor U527 (N_527,In_93,In_1877);
nor U528 (N_528,In_1771,In_785);
xnor U529 (N_529,In_2108,In_2092);
xor U530 (N_530,In_1717,In_1394);
nand U531 (N_531,In_2477,In_420);
and U532 (N_532,In_705,In_1633);
nor U533 (N_533,In_87,In_1813);
nor U534 (N_534,In_2902,In_2978);
or U535 (N_535,In_1991,In_2527);
nand U536 (N_536,In_1820,In_2022);
xnor U537 (N_537,In_871,In_1045);
nor U538 (N_538,In_2866,In_2293);
and U539 (N_539,In_1975,In_2990);
nor U540 (N_540,In_2166,In_2863);
xor U541 (N_541,In_1775,In_38);
or U542 (N_542,In_2014,In_1466);
nor U543 (N_543,In_1182,In_2037);
nand U544 (N_544,In_2680,In_2252);
nand U545 (N_545,In_1369,In_1650);
xor U546 (N_546,In_790,In_2382);
nand U547 (N_547,In_1594,In_1167);
nor U548 (N_548,In_2363,In_2273);
or U549 (N_549,In_75,In_2644);
nand U550 (N_550,In_584,In_1936);
and U551 (N_551,In_48,In_2941);
and U552 (N_552,In_415,In_153);
and U553 (N_553,In_1009,In_482);
and U554 (N_554,In_447,In_733);
or U555 (N_555,In_1430,In_840);
xor U556 (N_556,In_1478,In_625);
nand U557 (N_557,In_820,In_971);
nand U558 (N_558,In_216,In_870);
xnor U559 (N_559,In_2437,In_2017);
or U560 (N_560,In_955,In_854);
nor U561 (N_561,In_425,In_2261);
or U562 (N_562,In_858,In_1066);
xnor U563 (N_563,In_2842,In_2192);
xnor U564 (N_564,In_1740,In_2580);
nor U565 (N_565,In_1958,In_444);
xnor U566 (N_566,In_1562,In_317);
and U567 (N_567,In_1875,In_2754);
or U568 (N_568,In_214,In_230);
nand U569 (N_569,In_499,In_850);
nor U570 (N_570,In_2122,In_650);
and U571 (N_571,In_612,In_284);
xnor U572 (N_572,In_1473,In_2734);
or U573 (N_573,In_2052,In_1859);
nor U574 (N_574,In_402,In_780);
or U575 (N_575,In_2177,In_2927);
or U576 (N_576,In_2442,In_1407);
nor U577 (N_577,In_599,In_579);
nor U578 (N_578,In_1624,In_526);
xnor U579 (N_579,In_2226,In_1316);
and U580 (N_580,In_1464,In_2872);
nor U581 (N_581,In_1600,In_2669);
and U582 (N_582,In_2243,In_2563);
xor U583 (N_583,In_1754,In_495);
nand U584 (N_584,In_768,In_2309);
nand U585 (N_585,In_373,In_1647);
nor U586 (N_586,In_178,In_2189);
nor U587 (N_587,In_143,In_2098);
nand U588 (N_588,In_2331,In_2430);
xnor U589 (N_589,In_281,In_1451);
or U590 (N_590,In_2839,In_737);
nor U591 (N_591,In_2940,In_662);
xor U592 (N_592,In_2616,In_2648);
nand U593 (N_593,In_933,In_2890);
or U594 (N_594,In_1601,In_1008);
nand U595 (N_595,In_79,In_1785);
and U596 (N_596,In_2051,In_454);
and U597 (N_597,In_1746,In_2908);
nand U598 (N_598,In_2764,In_433);
or U599 (N_599,In_1812,In_2104);
and U600 (N_600,In_2275,In_1379);
or U601 (N_601,In_533,In_2266);
nor U602 (N_602,In_2421,In_491);
and U603 (N_603,In_2419,In_91);
or U604 (N_604,In_2262,In_898);
and U605 (N_605,In_2496,In_1894);
nor U606 (N_606,In_330,In_1472);
nor U607 (N_607,In_1994,In_1140);
nand U608 (N_608,In_2083,In_2010);
xnor U609 (N_609,In_24,In_1183);
or U610 (N_610,In_2087,In_426);
nand U611 (N_611,In_2552,In_1518);
nor U612 (N_612,In_2712,In_2520);
nor U613 (N_613,In_891,In_1085);
nand U614 (N_614,In_692,In_1504);
nand U615 (N_615,In_2561,In_743);
xnor U616 (N_616,In_94,In_329);
and U617 (N_617,In_1534,In_1983);
nor U618 (N_618,In_2251,In_2163);
nand U619 (N_619,In_2067,In_1531);
and U620 (N_620,In_31,In_1114);
nor U621 (N_621,In_103,In_923);
and U622 (N_622,In_1264,In_1150);
or U623 (N_623,In_2810,In_2270);
or U624 (N_624,In_2194,In_2582);
nand U625 (N_625,In_388,In_2543);
xnor U626 (N_626,In_939,In_96);
xor U627 (N_627,In_1341,In_1434);
and U628 (N_628,In_2871,In_1668);
or U629 (N_629,In_188,In_1881);
and U630 (N_630,In_2847,In_2765);
xnor U631 (N_631,In_2127,In_2149);
and U632 (N_632,In_2145,In_1095);
xnor U633 (N_633,In_200,In_2142);
and U634 (N_634,In_26,In_2229);
or U635 (N_635,In_1079,In_287);
or U636 (N_636,In_1089,In_1585);
and U637 (N_637,In_2844,In_55);
and U638 (N_638,In_456,In_739);
nand U639 (N_639,In_2770,In_427);
and U640 (N_640,In_1123,In_794);
xnor U641 (N_641,In_1999,In_393);
nor U642 (N_642,In_510,In_2977);
xnor U643 (N_643,In_2299,In_2830);
and U644 (N_644,In_2637,In_2393);
nor U645 (N_645,In_1350,In_1426);
nand U646 (N_646,In_2880,In_2231);
nor U647 (N_647,In_2837,In_2119);
and U648 (N_648,In_914,In_2930);
nand U649 (N_649,In_758,In_1891);
xor U650 (N_650,In_2002,In_2657);
and U651 (N_651,In_1299,In_403);
nand U652 (N_652,In_2759,In_950);
nand U653 (N_653,In_1226,In_2824);
nand U654 (N_654,In_2970,In_308);
and U655 (N_655,In_2094,In_784);
nor U656 (N_656,In_25,In_797);
nand U657 (N_657,In_1926,In_2230);
and U658 (N_658,In_1974,In_1442);
nor U659 (N_659,In_2725,In_102);
and U660 (N_660,In_2135,In_2756);
and U661 (N_661,In_825,In_1503);
and U662 (N_662,In_76,In_2332);
and U663 (N_663,In_1767,In_2599);
or U664 (N_664,In_555,In_57);
or U665 (N_665,In_517,In_2948);
xor U666 (N_666,In_2658,In_2779);
xnor U667 (N_667,In_1445,In_2018);
nor U668 (N_668,In_2535,In_1766);
and U669 (N_669,In_1516,In_171);
nor U670 (N_670,In_1567,In_538);
or U671 (N_671,In_2677,In_928);
and U672 (N_672,In_2480,In_2036);
xor U673 (N_673,In_117,In_2707);
xor U674 (N_674,In_1088,In_681);
nand U675 (N_675,In_2359,In_1564);
nor U676 (N_676,In_1697,In_328);
or U677 (N_677,In_480,In_513);
and U678 (N_678,In_1634,In_2789);
or U679 (N_679,In_2330,In_720);
and U680 (N_680,In_2947,In_1306);
xnor U681 (N_681,In_1423,In_1491);
or U682 (N_682,In_531,In_2894);
xnor U683 (N_683,In_2395,In_1852);
xor U684 (N_684,In_1630,In_815);
nand U685 (N_685,In_2541,In_1404);
or U686 (N_686,In_702,In_1869);
xnor U687 (N_687,In_1122,In_892);
and U688 (N_688,In_2356,In_1759);
xnor U689 (N_689,In_2325,In_1715);
xnor U690 (N_690,In_1631,In_2816);
or U691 (N_691,In_991,In_354);
and U692 (N_692,In_118,In_953);
nand U693 (N_693,In_688,In_630);
or U694 (N_694,In_674,In_2819);
xnor U695 (N_695,In_2435,In_2074);
nor U696 (N_696,In_2578,In_2740);
xnor U697 (N_697,In_1417,In_2350);
or U698 (N_698,In_2413,In_2446);
or U699 (N_699,In_1041,In_718);
nand U700 (N_700,In_817,In_1461);
or U701 (N_701,In_1854,In_1050);
or U702 (N_702,In_1651,In_864);
xor U703 (N_703,In_1188,In_2719);
nand U704 (N_704,In_467,In_2334);
nand U705 (N_705,In_1332,In_805);
or U706 (N_706,In_32,In_498);
xnor U707 (N_707,In_1197,In_2056);
nor U708 (N_708,In_254,In_324);
nand U709 (N_709,In_2415,In_2822);
nor U710 (N_710,In_1925,In_74);
nor U711 (N_711,In_2726,In_547);
nor U712 (N_712,In_11,In_70);
xnor U713 (N_713,In_1179,In_2416);
nand U714 (N_714,In_407,In_2720);
nor U715 (N_715,In_1235,In_2409);
and U716 (N_716,In_2783,In_2200);
xnor U717 (N_717,In_1612,In_1514);
or U718 (N_718,In_2248,In_1818);
nand U719 (N_719,In_1087,In_332);
or U720 (N_720,In_1397,In_1221);
nor U721 (N_721,In_157,In_2954);
nor U722 (N_722,In_837,In_2958);
or U723 (N_723,In_1452,In_159);
nand U724 (N_724,In_1055,In_595);
nand U725 (N_725,In_587,In_2820);
or U726 (N_726,In_1023,In_1082);
or U727 (N_727,In_1729,In_2512);
and U728 (N_728,In_233,In_1124);
xor U729 (N_729,In_1102,In_2033);
nand U730 (N_730,In_165,In_1892);
and U731 (N_731,In_2023,In_2086);
and U732 (N_732,In_2212,In_292);
nor U733 (N_733,In_647,In_1177);
or U734 (N_734,In_1919,In_789);
or U735 (N_735,In_1517,In_2351);
and U736 (N_736,In_807,In_1448);
or U737 (N_737,In_2202,In_2035);
and U738 (N_738,In_2800,In_1677);
or U739 (N_739,In_460,In_375);
and U740 (N_740,In_1268,In_1561);
nor U741 (N_741,In_1482,In_597);
and U742 (N_742,In_389,In_1987);
and U743 (N_743,In_715,In_90);
nand U744 (N_744,In_723,In_1780);
nand U745 (N_745,In_1826,In_272);
or U746 (N_746,In_1118,In_1217);
nor U747 (N_747,In_2172,In_1035);
or U748 (N_748,In_2068,In_516);
or U749 (N_749,In_2821,In_694);
xnor U750 (N_750,In_2403,In_384);
nand U751 (N_751,In_1481,In_747);
and U752 (N_752,In_2798,In_1401);
or U753 (N_753,In_994,In_2015);
or U754 (N_754,In_235,In_1701);
nor U755 (N_755,In_376,In_2242);
xnor U756 (N_756,In_1477,In_1823);
and U757 (N_757,In_2323,In_380);
and U758 (N_758,In_462,In_731);
and U759 (N_759,In_2290,In_707);
xor U760 (N_760,In_1738,In_2608);
xnor U761 (N_761,In_1455,In_872);
nand U762 (N_762,In_2203,In_774);
nor U763 (N_763,In_2869,In_2390);
and U764 (N_764,In_1040,In_2386);
or U765 (N_765,In_285,In_1128);
and U766 (N_766,In_2792,In_1372);
or U767 (N_767,In_470,In_1643);
and U768 (N_768,In_2053,In_2077);
and U769 (N_769,In_1224,In_485);
or U770 (N_770,In_1034,In_1750);
or U771 (N_771,In_541,In_2746);
and U772 (N_772,In_2529,In_2443);
and U773 (N_773,In_2634,In_1596);
nand U774 (N_774,In_1928,In_1876);
and U775 (N_775,In_1191,In_1325);
and U776 (N_776,In_154,In_2969);
and U777 (N_777,In_2348,In_853);
nor U778 (N_778,In_1840,In_901);
and U779 (N_779,In_1234,In_515);
nand U780 (N_780,In_601,In_1406);
xnor U781 (N_781,In_2081,In_182);
or U782 (N_782,In_1156,In_2558);
nand U783 (N_783,In_423,In_371);
and U784 (N_784,In_2804,In_477);
or U785 (N_785,In_675,In_2436);
nor U786 (N_786,In_2760,In_2876);
xor U787 (N_787,In_2361,In_732);
xnor U788 (N_788,In_2349,In_2886);
or U789 (N_789,In_1676,In_835);
nor U790 (N_790,In_1111,In_372);
and U791 (N_791,In_2901,In_2295);
and U792 (N_792,In_222,In_2458);
nand U793 (N_793,In_1727,In_738);
nor U794 (N_794,In_1276,In_684);
nand U795 (N_795,In_2656,In_1511);
and U796 (N_796,In_1684,In_2553);
and U797 (N_797,In_1402,In_777);
or U798 (N_798,In_1539,In_811);
and U799 (N_799,In_2864,In_1456);
and U800 (N_800,In_1354,In_311);
nor U801 (N_801,In_2107,In_1154);
or U802 (N_802,In_2704,In_2284);
nand U803 (N_803,In_2136,In_2080);
and U804 (N_804,In_2628,In_296);
and U805 (N_805,In_2407,In_1732);
nand U806 (N_806,In_1252,In_2453);
xor U807 (N_807,In_1779,In_360);
and U808 (N_808,In_2198,In_133);
or U809 (N_809,In_2728,In_1526);
or U810 (N_810,In_535,In_2019);
or U811 (N_811,In_1844,In_2651);
or U812 (N_812,In_632,In_191);
and U813 (N_813,In_1942,In_1247);
nor U814 (N_814,In_2178,In_2150);
nor U815 (N_815,In_2201,In_2271);
nor U816 (N_816,In_1228,In_2639);
xnor U817 (N_817,In_2774,In_995);
nand U818 (N_818,In_2923,In_1265);
nor U819 (N_819,In_2100,In_1758);
and U820 (N_820,In_2399,In_2911);
or U821 (N_821,In_1946,In_2865);
nand U822 (N_822,In_2618,In_2516);
nand U823 (N_823,In_1664,In_608);
nand U824 (N_824,In_2629,In_378);
xor U825 (N_825,In_917,In_561);
xor U826 (N_826,In_496,In_1279);
nand U827 (N_827,In_795,In_988);
nor U828 (N_828,In_1721,In_1745);
nand U829 (N_829,In_1816,In_80);
nor U830 (N_830,In_349,In_1827);
nand U831 (N_831,In_2319,In_1000);
or U832 (N_832,In_307,In_1955);
nor U833 (N_833,In_2539,In_2470);
and U834 (N_834,In_640,In_1170);
or U835 (N_835,In_1868,In_2233);
nor U836 (N_836,In_906,In_2167);
nor U837 (N_837,In_2315,In_2640);
nor U838 (N_838,In_529,In_114);
xor U839 (N_839,In_2101,In_2609);
xor U840 (N_840,In_2287,In_1659);
nand U841 (N_841,In_1483,In_639);
and U842 (N_842,In_573,In_2311);
nand U843 (N_843,In_2066,In_464);
or U844 (N_844,In_150,In_457);
or U845 (N_845,In_1814,In_58);
or U846 (N_846,In_121,In_1382);
or U847 (N_847,In_912,In_2542);
and U848 (N_848,In_2854,In_298);
nand U849 (N_849,In_17,In_620);
nand U850 (N_850,In_2833,In_2383);
nor U851 (N_851,In_576,In_643);
nor U852 (N_852,In_1086,In_394);
and U853 (N_853,In_1303,In_2505);
xnor U854 (N_854,In_1787,In_2109);
nand U855 (N_855,In_2027,In_2758);
nand U856 (N_856,In_865,In_2116);
and U857 (N_857,In_839,In_240);
or U858 (N_858,In_2910,In_2604);
nand U859 (N_859,In_72,In_127);
or U860 (N_860,In_961,In_1164);
nor U861 (N_861,In_1365,In_205);
xnor U862 (N_862,In_2481,In_728);
nand U863 (N_863,In_2622,In_77);
nor U864 (N_864,In_1550,In_1465);
and U865 (N_865,In_2905,In_2485);
nand U866 (N_866,In_1028,In_2047);
and U867 (N_867,In_2690,In_271);
nand U868 (N_868,In_2218,In_2596);
or U869 (N_869,In_1229,In_539);
nand U870 (N_870,In_437,In_2518);
or U871 (N_871,In_479,In_1334);
nor U872 (N_872,In_2428,In_488);
nand U873 (N_873,In_2589,In_2884);
nand U874 (N_874,In_2642,In_753);
xor U875 (N_875,In_983,In_1218);
xor U876 (N_876,In_413,In_2682);
nor U877 (N_877,In_2900,In_2246);
nor U878 (N_878,In_1184,In_2445);
xnor U879 (N_879,In_1292,In_442);
nand U880 (N_880,In_116,In_2468);
or U881 (N_881,In_2298,In_2737);
or U882 (N_882,In_1988,In_1652);
nor U883 (N_883,In_2199,In_1155);
nor U884 (N_884,In_89,In_2831);
and U885 (N_885,In_1920,In_1524);
nor U886 (N_886,In_1784,In_196);
or U887 (N_887,In_558,In_2811);
xor U888 (N_888,In_2269,In_1953);
nand U889 (N_889,In_1304,In_1470);
nand U890 (N_890,In_2879,In_1213);
and U891 (N_891,In_1736,In_1900);
nor U892 (N_892,In_2103,In_1385);
nand U893 (N_893,In_2255,In_796);
xor U894 (N_894,In_646,In_1249);
and U895 (N_895,In_1003,In_636);
nor U896 (N_896,In_1259,In_512);
xnor U897 (N_897,In_570,In_68);
nand U898 (N_898,In_198,In_2424);
or U899 (N_899,In_1318,In_1689);
and U900 (N_900,In_1392,In_766);
or U901 (N_901,In_2951,In_2776);
xor U902 (N_902,In_2120,In_580);
nor U903 (N_903,In_2030,In_1856);
nor U904 (N_904,In_2727,In_889);
xor U905 (N_905,In_294,In_924);
and U906 (N_906,In_756,In_1923);
nand U907 (N_907,In_586,In_2611);
xor U908 (N_908,In_1244,In_2689);
and U909 (N_909,In_574,In_1185);
and U910 (N_910,In_2151,In_549);
nor U911 (N_911,In_362,In_849);
and U912 (N_912,In_140,In_2936);
nand U913 (N_913,In_2358,In_1216);
nand U914 (N_914,In_1625,In_1728);
and U915 (N_915,In_1632,In_1091);
xnor U916 (N_916,In_315,In_2341);
and U917 (N_917,In_63,In_1734);
or U918 (N_918,In_2026,In_268);
nand U919 (N_919,In_2038,In_680);
nor U920 (N_920,In_149,In_2183);
or U921 (N_921,In_542,In_1523);
and U922 (N_922,In_36,In_283);
or U923 (N_923,In_2603,In_616);
nor U924 (N_924,In_2873,In_521);
xor U925 (N_925,In_2623,In_2186);
xor U926 (N_926,In_1706,In_2588);
or U927 (N_927,In_1125,In_693);
or U928 (N_928,In_1284,In_1575);
nand U929 (N_929,In_2222,In_593);
or U930 (N_930,In_459,In_1948);
and U931 (N_931,In_183,In_33);
or U932 (N_932,In_1753,In_511);
or U933 (N_933,In_2787,In_151);
and U934 (N_934,In_721,In_2239);
nor U935 (N_935,In_848,In_82);
or U936 (N_936,In_2132,In_2138);
and U937 (N_937,In_2434,In_2613);
or U938 (N_938,In_658,In_937);
nor U939 (N_939,In_2953,In_13);
xor U940 (N_940,In_1312,In_1569);
nand U941 (N_941,In_391,In_1210);
nor U942 (N_942,In_2858,In_1339);
nor U943 (N_943,In_2209,In_2071);
nor U944 (N_944,In_810,In_882);
and U945 (N_945,In_1815,In_1262);
nand U946 (N_946,In_1340,In_469);
or U947 (N_947,In_1570,In_1062);
nand U948 (N_948,In_16,In_2713);
nor U949 (N_949,In_1636,In_2630);
and U950 (N_950,In_2491,In_2519);
nor U951 (N_951,In_364,In_2773);
nor U952 (N_952,In_1360,In_671);
or U953 (N_953,In_2420,In_2431);
xor U954 (N_954,In_2258,In_885);
or U955 (N_955,In_2326,In_359);
nand U956 (N_956,In_1108,In_1962);
and U957 (N_957,In_1637,In_2514);
xor U958 (N_958,In_2717,In_2366);
nand U959 (N_959,In_965,In_2472);
nand U960 (N_960,In_1007,In_2020);
nand U961 (N_961,In_1441,In_649);
nor U962 (N_962,In_1301,In_812);
nor U963 (N_963,In_304,In_2985);
xor U964 (N_964,In_1588,In_1911);
and U965 (N_965,In_279,In_1670);
or U966 (N_966,In_969,In_2922);
or U967 (N_967,In_2600,In_956);
nand U968 (N_968,In_1599,In_2736);
and U969 (N_969,In_1002,In_1454);
nand U970 (N_970,In_514,In_1710);
nor U971 (N_971,In_946,In_1342);
nand U972 (N_972,In_215,In_504);
nor U973 (N_973,In_2380,In_2997);
nor U974 (N_974,In_345,In_1887);
xnor U975 (N_975,In_1907,In_1969);
and U976 (N_976,In_1931,In_228);
nand U977 (N_977,In_545,In_2034);
nor U978 (N_978,In_1212,In_282);
xnor U979 (N_979,In_1208,In_890);
nand U980 (N_980,In_2438,In_2410);
and U981 (N_981,In_2197,In_1932);
nand U982 (N_982,In_2963,In_619);
or U983 (N_983,In_347,In_1136);
and U984 (N_984,In_2857,In_148);
or U985 (N_985,In_651,In_186);
nor U986 (N_986,In_2355,In_2550);
or U987 (N_987,In_1795,In_158);
nor U988 (N_988,In_2585,In_968);
xnor U989 (N_989,In_691,In_2913);
nor U990 (N_990,In_2952,In_1485);
xor U991 (N_991,In_1770,In_2475);
nand U992 (N_992,In_2211,In_1250);
or U993 (N_993,In_1924,In_2673);
xor U994 (N_994,In_1703,In_1617);
and U995 (N_995,In_1432,In_2158);
and U996 (N_996,In_2500,In_2915);
xor U997 (N_997,In_2448,In_1453);
and U998 (N_998,In_1598,In_2441);
xor U999 (N_999,In_918,In_2684);
nor U1000 (N_1000,In_136,In_2698);
and U1001 (N_1001,In_1479,In_2400);
nor U1002 (N_1002,In_537,In_1105);
and U1003 (N_1003,In_1809,In_472);
and U1004 (N_1004,In_2084,In_2652);
nand U1005 (N_1005,In_949,In_943);
and U1006 (N_1006,In_1595,In_156);
or U1007 (N_1007,In_764,In_1909);
nor U1008 (N_1008,In_1915,In_1799);
or U1009 (N_1009,In_1644,In_2976);
xor U1010 (N_1010,In_2354,In_534);
nor U1011 (N_1011,In_696,In_1187);
xor U1012 (N_1012,In_1329,In_119);
nor U1013 (N_1013,In_2362,In_2454);
nor U1014 (N_1014,In_107,In_2593);
or U1015 (N_1015,In_984,In_1116);
nand U1016 (N_1016,In_2878,In_657);
or U1017 (N_1017,In_187,In_1355);
nand U1018 (N_1018,In_2179,In_2627);
and U1019 (N_1019,In_686,In_2316);
or U1020 (N_1020,In_957,In_2861);
nand U1021 (N_1021,In_1501,In_1266);
nand U1022 (N_1022,In_1711,In_966);
xnor U1023 (N_1023,In_1139,In_144);
nand U1024 (N_1024,In_808,In_2920);
xor U1025 (N_1025,In_351,In_1610);
or U1026 (N_1026,In_2099,In_1521);
xor U1027 (N_1027,In_408,In_1178);
nand U1028 (N_1028,In_2612,In_2590);
nor U1029 (N_1029,In_357,In_64);
nand U1030 (N_1030,In_1443,In_50);
nand U1031 (N_1031,In_2574,In_954);
and U1032 (N_1032,In_1989,In_2602);
nor U1033 (N_1033,In_1831,In_1878);
xor U1034 (N_1034,In_2565,In_1733);
nor U1035 (N_1035,In_2840,In_1586);
xnor U1036 (N_1036,In_2302,In_1358);
nand U1037 (N_1037,In_1072,In_128);
nor U1038 (N_1038,In_2891,In_990);
nand U1039 (N_1039,In_1317,In_1039);
and U1040 (N_1040,In_689,In_1162);
nor U1041 (N_1041,In_1761,In_1399);
xnor U1042 (N_1042,In_2768,In_2304);
and U1043 (N_1043,In_2841,In_746);
nand U1044 (N_1044,In_1422,In_869);
nor U1045 (N_1045,In_827,In_659);
xnor U1046 (N_1046,In_927,In_1593);
nor U1047 (N_1047,In_2058,In_2507);
xnor U1048 (N_1048,In_2143,In_2404);
and U1049 (N_1049,In_321,In_2548);
or U1050 (N_1050,In_940,In_1043);
nor U1051 (N_1051,In_1742,In_147);
nand U1052 (N_1052,In_2601,In_741);
xnor U1053 (N_1053,In_628,In_1277);
or U1054 (N_1054,In_2932,In_568);
nor U1055 (N_1055,In_2364,In_313);
and U1056 (N_1056,In_2935,In_2274);
and U1057 (N_1057,In_2745,In_793);
nor U1058 (N_1058,In_2130,In_974);
xnor U1059 (N_1059,In_944,In_2856);
nor U1060 (N_1060,In_1897,In_2140);
nor U1061 (N_1061,In_1880,In_325);
xor U1062 (N_1062,In_2494,In_2870);
or U1063 (N_1063,In_2265,In_638);
or U1064 (N_1064,In_2306,In_1560);
or U1065 (N_1065,In_1904,In_1547);
and U1066 (N_1066,In_1688,In_1791);
nand U1067 (N_1067,In_879,In_1149);
xor U1068 (N_1068,In_2663,In_819);
and U1069 (N_1069,In_1797,In_1373);
and U1070 (N_1070,In_2662,In_40);
nand U1071 (N_1071,In_2715,In_342);
and U1072 (N_1072,In_1901,In_2134);
or U1073 (N_1073,In_2993,In_1077);
nor U1074 (N_1074,In_1390,In_1930);
or U1075 (N_1075,In_2832,In_1398);
and U1076 (N_1076,In_1764,In_189);
xor U1077 (N_1077,In_2335,In_697);
and U1078 (N_1078,In_353,In_411);
xnor U1079 (N_1079,In_609,In_343);
and U1080 (N_1080,In_1152,In_1413);
nor U1081 (N_1081,In_2257,In_1033);
and U1082 (N_1082,In_2699,In_1321);
xor U1083 (N_1083,In_2692,In_873);
nor U1084 (N_1084,In_1215,In_2909);
and U1085 (N_1085,In_2296,In_1117);
and U1086 (N_1086,In_759,In_2152);
and U1087 (N_1087,In_399,In_97);
nor U1088 (N_1088,In_14,In_1367);
or U1089 (N_1089,In_2471,In_1822);
xor U1090 (N_1090,In_336,In_1546);
nor U1091 (N_1091,In_1532,In_565);
or U1092 (N_1092,In_246,In_167);
nand U1093 (N_1093,In_1682,In_1307);
and U1094 (N_1094,In_2228,In_592);
nor U1095 (N_1095,In_2352,In_2455);
or U1096 (N_1096,In_1391,In_1707);
or U1097 (N_1097,In_2336,In_2907);
xor U1098 (N_1098,In_979,In_2238);
and U1099 (N_1099,In_2859,In_2314);
nand U1100 (N_1100,In_2559,In_1870);
xnor U1101 (N_1101,In_2337,In_2635);
nor U1102 (N_1102,In_1314,In_1071);
nor U1103 (N_1103,In_2088,In_2123);
nand U1104 (N_1104,In_2128,In_1843);
or U1105 (N_1105,In_267,In_2462);
xor U1106 (N_1106,In_1137,In_1274);
or U1107 (N_1107,In_2526,In_945);
and U1108 (N_1108,In_1032,In_2742);
or U1109 (N_1109,In_1440,In_2732);
xor U1110 (N_1110,In_1267,In_1290);
and U1111 (N_1111,In_803,In_1971);
or U1112 (N_1112,In_293,In_1914);
or U1113 (N_1113,In_1506,In_398);
nor U1114 (N_1114,In_1858,In_1239);
or U1115 (N_1115,In_42,In_1022);
or U1116 (N_1116,In_1819,In_2115);
nand U1117 (N_1117,In_1065,In_85);
nor U1118 (N_1118,In_1493,In_2807);
xor U1119 (N_1119,In_771,In_2945);
and U1120 (N_1120,In_2456,In_43);
or U1121 (N_1121,In_1386,In_710);
and U1122 (N_1122,In_1679,In_2148);
or U1123 (N_1123,In_2237,In_1436);
and U1124 (N_1124,In_1952,In_62);
and U1125 (N_1125,In_1765,In_2916);
and U1126 (N_1126,In_1978,In_1192);
nor U1127 (N_1127,In_1467,In_2893);
and U1128 (N_1128,In_1186,In_35);
nand U1129 (N_1129,In_47,In_1591);
xnor U1130 (N_1130,In_787,In_422);
or U1131 (N_1131,In_2310,In_2961);
nor U1132 (N_1132,In_2739,In_1371);
xnor U1133 (N_1133,In_2785,In_1667);
nand U1134 (N_1134,In_2605,In_277);
or U1135 (N_1135,In_1963,In_2024);
nor U1136 (N_1136,In_1425,In_2898);
and U1137 (N_1137,In_1495,In_2942);
or U1138 (N_1138,In_2169,In_1655);
nor U1139 (N_1139,In_2615,In_1051);
xor U1140 (N_1140,In_1253,In_856);
xor U1141 (N_1141,In_2524,In_261);
or U1142 (N_1142,In_2216,In_1319);
xnor U1143 (N_1143,In_564,In_1047);
or U1144 (N_1144,In_2078,In_792);
or U1145 (N_1145,In_2946,In_627);
nand U1146 (N_1146,In_2705,In_1557);
nor U1147 (N_1147,In_2703,In_1793);
nand U1148 (N_1148,In_1574,In_37);
and U1149 (N_1149,In_211,In_1976);
and U1150 (N_1150,In_2089,In_604);
nor U1151 (N_1151,In_941,In_550);
or U1152 (N_1152,In_41,In_2488);
xnor U1153 (N_1153,In_1147,In_2118);
nand U1154 (N_1154,In_2752,In_300);
or U1155 (N_1155,In_2995,In_1494);
xor U1156 (N_1156,In_970,In_2694);
and U1157 (N_1157,In_2046,In_1351);
xor U1158 (N_1158,In_1507,In_1134);
or U1159 (N_1159,In_611,In_1471);
xnor U1160 (N_1160,In_2836,In_452);
nor U1161 (N_1161,In_1013,In_2282);
nand U1162 (N_1162,In_806,In_112);
nor U1163 (N_1163,In_434,In_1848);
nand U1164 (N_1164,In_1333,In_1435);
and U1165 (N_1165,In_1313,In_2156);
xnor U1166 (N_1166,In_71,In_1195);
or U1167 (N_1167,In_195,In_2984);
nand U1168 (N_1168,In_1327,In_306);
nand U1169 (N_1169,In_1427,In_2131);
nand U1170 (N_1170,In_722,In_2675);
nand U1171 (N_1171,In_1256,In_2224);
and U1172 (N_1172,In_727,In_982);
xor U1173 (N_1173,In_2534,In_438);
xor U1174 (N_1174,In_2057,In_217);
and U1175 (N_1175,In_641,In_44);
xor U1176 (N_1176,In_981,In_2493);
nand U1177 (N_1177,In_2313,In_930);
or U1178 (N_1178,In_2729,In_1233);
nand U1179 (N_1179,In_2225,In_2654);
xor U1180 (N_1180,In_2755,In_2849);
nor U1181 (N_1181,In_370,In_635);
xor U1182 (N_1182,In_1109,In_1828);
xnor U1183 (N_1183,In_213,In_2444);
or U1184 (N_1184,In_1227,In_2934);
or U1185 (N_1185,In_1527,In_1054);
xor U1186 (N_1186,In_2144,In_39);
nand U1187 (N_1187,In_1206,In_2249);
nand U1188 (N_1188,In_1629,In_2162);
xor U1189 (N_1189,In_184,In_915);
xnor U1190 (N_1190,In_476,In_987);
or U1191 (N_1191,In_735,In_355);
xnor U1192 (N_1192,In_137,In_1597);
nor U1193 (N_1193,In_276,In_1825);
nand U1194 (N_1194,In_2406,In_2598);
or U1195 (N_1195,In_295,In_465);
and U1196 (N_1196,In_18,In_418);
nand U1197 (N_1197,In_2892,In_2048);
or U1198 (N_1198,In_255,In_245);
nand U1199 (N_1199,In_1067,In_2297);
or U1200 (N_1200,In_2263,In_1690);
xnor U1201 (N_1201,In_1291,In_845);
xnor U1202 (N_1202,In_2999,In_2232);
nand U1203 (N_1203,In_1537,In_2032);
and U1204 (N_1204,In_2571,In_2506);
nand U1205 (N_1205,In_131,In_1037);
nor U1206 (N_1206,In_99,In_2322);
and U1207 (N_1207,In_326,In_1695);
or U1208 (N_1208,In_1378,In_463);
or U1209 (N_1209,In_1113,In_563);
and U1210 (N_1210,In_875,In_1201);
and U1211 (N_1211,In_1261,In_2075);
nand U1212 (N_1212,In_605,In_1589);
or U1213 (N_1213,In_1048,In_2182);
nand U1214 (N_1214,In_1353,In_2093);
or U1215 (N_1215,In_1607,In_2155);
nand U1216 (N_1216,In_1568,In_1762);
xor U1217 (N_1217,In_1899,In_824);
or U1218 (N_1218,In_303,In_2005);
or U1219 (N_1219,In_1558,In_1231);
or U1220 (N_1220,In_2268,In_700);
xor U1221 (N_1221,In_904,In_2581);
nor U1222 (N_1222,In_857,In_2208);
nor U1223 (N_1223,In_2817,In_2706);
xor U1224 (N_1224,In_2751,In_53);
nor U1225 (N_1225,In_490,In_1519);
xnor U1226 (N_1226,In_1176,In_2835);
or U1227 (N_1227,In_2173,In_2636);
nor U1228 (N_1228,In_2308,In_1092);
and U1229 (N_1229,In_227,In_2377);
nand U1230 (N_1230,In_1396,In_1879);
xor U1231 (N_1231,In_2041,In_834);
and U1232 (N_1232,In_1940,In_528);
and U1233 (N_1233,In_2003,In_92);
nor U1234 (N_1234,In_280,In_481);
xor U1235 (N_1235,In_385,In_1019);
nor U1236 (N_1236,In_823,In_1751);
and U1237 (N_1237,In_1225,In_2259);
xor U1238 (N_1238,In_0,In_818);
nand U1239 (N_1239,In_1873,In_1403);
and U1240 (N_1240,In_763,In_2906);
xor U1241 (N_1241,In_2007,In_1414);
nor U1242 (N_1242,In_2862,In_2288);
nor U1243 (N_1243,In_493,In_2607);
nor U1244 (N_1244,In_1376,In_377);
nand U1245 (N_1245,In_1722,In_2570);
nand U1246 (N_1246,In_653,In_830);
xor U1247 (N_1247,In_1352,In_1883);
and U1248 (N_1248,In_2191,In_1103);
nor U1249 (N_1249,In_846,In_1120);
nand U1250 (N_1250,In_1804,In_193);
nor U1251 (N_1251,In_2294,In_648);
or U1252 (N_1252,In_2473,In_2091);
xnor U1253 (N_1253,In_932,In_201);
nand U1254 (N_1254,In_613,In_2502);
xor U1255 (N_1255,In_1056,In_2124);
nor U1256 (N_1256,In_1357,In_1060);
nand U1257 (N_1257,In_2375,In_2875);
or U1258 (N_1258,In_365,In_2780);
and U1259 (N_1259,In_1980,In_2012);
nor U1260 (N_1260,In_2008,In_2775);
xnor U1261 (N_1261,In_2594,In_289);
xnor U1262 (N_1262,In_2686,In_855);
nor U1263 (N_1263,In_670,In_1269);
nor U1264 (N_1264,In_2797,In_687);
and U1265 (N_1265,In_2370,In_409);
and U1266 (N_1266,In_1871,In_1090);
nor U1267 (N_1267,In_250,In_2799);
nor U1268 (N_1268,In_1129,In_1375);
nor U1269 (N_1269,In_1673,In_2244);
nor U1270 (N_1270,In_1565,In_475);
and U1271 (N_1271,In_1641,In_813);
and U1272 (N_1272,In_1805,In_729);
nor U1273 (N_1273,In_2039,In_1174);
and U1274 (N_1274,In_1438,In_2095);
nand U1275 (N_1275,In_397,In_2557);
nor U1276 (N_1276,In_1308,In_2160);
nand U1277 (N_1277,In_931,In_1064);
and U1278 (N_1278,In_1220,In_1349);
xnor U1279 (N_1279,In_1143,In_2829);
or U1280 (N_1280,In_2709,In_1886);
xnor U1281 (N_1281,In_1773,In_278);
xnor U1282 (N_1282,In_997,In_2346);
and U1283 (N_1283,In_390,In_2070);
nand U1284 (N_1284,In_2943,In_726);
nor U1285 (N_1285,In_583,In_769);
nand U1286 (N_1286,In_2931,In_2389);
and U1287 (N_1287,In_309,In_2515);
or U1288 (N_1288,In_258,In_2531);
nand U1289 (N_1289,In_2450,In_2285);
nand U1290 (N_1290,In_2671,In_1068);
or U1291 (N_1291,In_1500,In_344);
or U1292 (N_1292,In_1475,In_1782);
and U1293 (N_1293,In_65,In_2478);
nor U1294 (N_1294,In_1739,In_2885);
and U1295 (N_1295,In_1992,In_1410);
nand U1296 (N_1296,In_978,In_443);
nand U1297 (N_1297,In_1772,In_1656);
xor U1298 (N_1298,In_1520,In_762);
nor U1299 (N_1299,In_2215,In_2579);
or U1300 (N_1300,In_2312,In_951);
xnor U1301 (N_1301,In_2544,In_1834);
xnor U1302 (N_1302,In_1337,In_374);
and U1303 (N_1303,In_2277,In_916);
or U1304 (N_1304,In_2451,In_2646);
nand U1305 (N_1305,In_2560,In_288);
xor U1306 (N_1306,In_1310,In_1584);
nand U1307 (N_1307,In_2388,In_585);
nand U1308 (N_1308,In_319,In_2808);
xnor U1309 (N_1309,In_2749,In_1258);
or U1310 (N_1310,In_2204,In_2025);
nand U1311 (N_1311,In_2914,In_778);
xnor U1312 (N_1312,In_125,In_617);
or U1313 (N_1313,In_386,In_1921);
xor U1314 (N_1314,In_1853,In_1075);
xor U1315 (N_1315,In_2813,In_1363);
or U1316 (N_1316,In_2660,In_557);
nor U1317 (N_1317,In_259,In_113);
xor U1318 (N_1318,In_2975,In_2850);
and U1319 (N_1319,In_1161,In_663);
and U1320 (N_1320,In_1021,In_2546);
xor U1321 (N_1321,In_2133,In_2591);
xor U1322 (N_1322,In_1393,In_816);
or U1323 (N_1323,In_2059,In_494);
nor U1324 (N_1324,In_2691,In_1566);
xor U1325 (N_1325,In_2072,In_2801);
nand U1326 (N_1326,In_1416,In_241);
or U1327 (N_1327,In_1864,In_2112);
and U1328 (N_1328,In_2881,In_2851);
nand U1329 (N_1329,In_2227,In_164);
nor U1330 (N_1330,In_2385,In_1847);
nand U1331 (N_1331,In_231,In_866);
or U1332 (N_1332,In_704,In_1660);
nor U1333 (N_1333,In_2533,In_2572);
xnor U1334 (N_1334,In_2903,In_1486);
and U1335 (N_1335,In_1207,In_2344);
xnor U1336 (N_1336,In_1444,In_1121);
xor U1337 (N_1337,In_2374,In_1141);
xor U1338 (N_1338,In_1555,In_569);
or U1339 (N_1339,In_242,In_1615);
and U1340 (N_1340,In_2241,In_322);
nor U1341 (N_1341,In_802,In_578);
nor U1342 (N_1342,In_2469,In_683);
nor U1343 (N_1343,In_2724,In_468);
xnor U1344 (N_1344,In_886,In_2653);
nand U1345 (N_1345,In_95,In_761);
and U1346 (N_1346,In_1903,In_2555);
and U1347 (N_1347,In_66,In_1760);
nor U1348 (N_1348,In_1553,In_2234);
nor U1349 (N_1349,In_168,In_1905);
or U1350 (N_1350,In_220,In_973);
nand U1351 (N_1351,In_1236,In_861);
or U1352 (N_1352,In_1110,In_2141);
xnor U1353 (N_1353,In_1941,In_1025);
and U1354 (N_1354,In_1587,In_798);
and U1355 (N_1355,In_831,In_2855);
or U1356 (N_1356,In_199,In_577);
or U1357 (N_1357,In_2766,In_1898);
and U1358 (N_1358,In_1010,In_1982);
nand U1359 (N_1359,In_695,In_197);
nor U1360 (N_1360,In_525,In_2803);
nand U1361 (N_1361,In_2695,In_750);
nor U1362 (N_1362,In_1951,In_1661);
and U1363 (N_1363,In_2171,In_314);
nand U1364 (N_1364,In_172,In_938);
nand U1365 (N_1365,In_667,In_2614);
xor U1366 (N_1366,In_2510,In_2372);
and U1367 (N_1367,In_2278,In_1189);
nand U1368 (N_1368,In_130,In_1752);
xnor U1369 (N_1369,In_1159,In_346);
and U1370 (N_1370,In_1888,In_1323);
xnor U1371 (N_1371,In_1242,In_234);
and U1372 (N_1372,In_536,In_2853);
nor U1373 (N_1373,In_1872,In_712);
or U1374 (N_1374,In_2305,In_1005);
or U1375 (N_1375,In_2031,In_2771);
and U1376 (N_1376,In_1280,In_1181);
xor U1377 (N_1377,In_624,In_2980);
and U1378 (N_1378,In_1675,In_859);
nor U1379 (N_1379,In_2919,In_588);
and U1380 (N_1380,In_10,In_266);
nor U1381 (N_1381,In_1018,In_1916);
nand U1382 (N_1382,In_2610,In_162);
xor U1383 (N_1383,In_626,In_905);
nand U1384 (N_1384,In_2681,In_880);
nand U1385 (N_1385,In_2846,In_591);
xnor U1386 (N_1386,In_291,In_1165);
and U1387 (N_1387,In_1364,In_1046);
or U1388 (N_1388,In_1429,In_2497);
or U1389 (N_1389,In_633,In_473);
nor U1390 (N_1390,In_1411,In_225);
nand U1391 (N_1391,In_2664,In_1646);
and U1392 (N_1392,In_1798,In_2196);
nor U1393 (N_1393,In_740,In_1674);
or U1394 (N_1394,In_1867,In_146);
and U1395 (N_1395,In_1405,In_2217);
and U1396 (N_1396,In_1543,In_1042);
nor U1397 (N_1397,In_1076,In_645);
and U1398 (N_1398,In_1544,In_2157);
nor U1399 (N_1399,In_2538,In_2744);
or U1400 (N_1400,In_1571,In_2264);
and U1401 (N_1401,In_2701,In_2794);
nor U1402 (N_1402,In_1692,In_505);
xor U1403 (N_1403,In_1297,In_2874);
nand U1404 (N_1404,In_1960,In_1944);
and U1405 (N_1405,In_913,In_1528);
and U1406 (N_1406,In_2988,In_2795);
nor U1407 (N_1407,In_352,In_2696);
or U1408 (N_1408,In_1977,In_2440);
nand U1409 (N_1409,In_1257,In_2950);
xor U1410 (N_1410,In_977,In_826);
nand U1411 (N_1411,In_2412,In_1383);
and U1412 (N_1412,In_1388,In_800);
nand U1413 (N_1413,In_2678,In_1801);
nor U1414 (N_1414,In_2672,In_985);
xor U1415 (N_1415,In_2567,In_2147);
or U1416 (N_1416,In_2499,In_1271);
and U1417 (N_1417,In_1171,In_1408);
nand U1418 (N_1418,In_1837,In_108);
nor U1419 (N_1419,In_2626,In_2303);
nand U1420 (N_1420,In_560,In_2321);
and U1421 (N_1421,In_2394,In_2267);
nand U1422 (N_1422,In_2536,In_1947);
nor U1423 (N_1423,In_2333,In_257);
nor U1424 (N_1424,In_449,In_1298);
xor U1425 (N_1425,In_1409,In_1933);
nor U1426 (N_1426,In_67,In_2904);
and U1427 (N_1427,In_2761,In_1902);
xnor U1428 (N_1428,In_2649,In_1730);
or U1429 (N_1429,In_2583,In_581);
or U1430 (N_1430,In_1428,In_1522);
and U1431 (N_1431,In_2938,In_2762);
xor U1432 (N_1432,In_911,In_503);
or U1433 (N_1433,In_1288,In_1180);
nor U1434 (N_1434,In_2918,In_1972);
nor U1435 (N_1435,In_652,In_484);
nor U1436 (N_1436,In_1620,In_801);
nand U1437 (N_1437,In_2339,In_2750);
xor U1438 (N_1438,In_122,In_1131);
or U1439 (N_1439,In_2964,In_519);
or U1440 (N_1440,In_2595,In_1657);
nor U1441 (N_1441,In_2974,In_1648);
xor U1442 (N_1442,In_1157,In_356);
nand U1443 (N_1443,In_51,In_2679);
nor U1444 (N_1444,In_334,In_166);
and U1445 (N_1445,In_622,In_253);
nor U1446 (N_1446,In_2113,In_989);
nand U1447 (N_1447,In_2786,In_1029);
nor U1448 (N_1448,In_202,In_2852);
xor U1449 (N_1449,In_98,In_1882);
xor U1450 (N_1450,In_540,In_2318);
xor U1451 (N_1451,In_2111,In_2743);
and U1452 (N_1452,In_2826,In_34);
and U1453 (N_1453,In_1623,In_690);
xnor U1454 (N_1454,In_2549,In_2042);
xnor U1455 (N_1455,In_194,In_1151);
nor U1456 (N_1456,In_1255,In_1845);
nand U1457 (N_1457,In_2176,In_1457);
nor U1458 (N_1458,In_2253,In_883);
or U1459 (N_1459,In_644,In_1214);
nand U1460 (N_1460,In_713,In_175);
or U1461 (N_1461,In_1015,In_1849);
and U1462 (N_1462,In_2912,In_919);
nor U1463 (N_1463,In_1496,In_1959);
and U1464 (N_1464,In_2597,In_1283);
nor U1465 (N_1465,In_1981,In_2106);
nand U1466 (N_1466,In_448,In_909);
and U1467 (N_1467,In_685,In_1691);
and U1468 (N_1468,In_1273,In_428);
and U1469 (N_1469,In_163,In_2665);
and U1470 (N_1470,In_895,In_2139);
nor U1471 (N_1471,In_1074,In_2423);
nand U1472 (N_1472,In_387,In_2205);
or U1473 (N_1473,In_1694,In_2979);
nand U1474 (N_1474,In_2050,In_2687);
xnor U1475 (N_1475,In_1505,In_1492);
or U1476 (N_1476,In_1525,In_2490);
nor U1477 (N_1477,In_238,In_1036);
xor U1478 (N_1478,In_2376,In_2193);
or U1479 (N_1479,In_1606,In_1579);
and U1480 (N_1480,In_2079,In_1861);
nand U1481 (N_1481,In_273,In_999);
xnor U1482 (N_1482,In_430,In_767);
nor U1483 (N_1483,In_1986,In_1893);
or U1484 (N_1484,In_929,In_1748);
and U1485 (N_1485,In_959,In_631);
and U1486 (N_1486,In_2459,In_1696);
or U1487 (N_1487,In_2126,In_1278);
xnor U1488 (N_1488,In_1922,In_841);
nand U1489 (N_1489,In_2981,In_1627);
and U1490 (N_1490,In_821,In_958);
nor U1491 (N_1491,In_134,In_1031);
and U1492 (N_1492,In_1194,In_2004);
nand U1493 (N_1493,In_934,In_1419);
nor U1494 (N_1494,In_2586,In_2782);
or U1495 (N_1495,In_2427,In_1829);
or U1496 (N_1496,In_455,In_548);
nand U1497 (N_1497,In_1996,In_530);
or U1498 (N_1498,In_860,In_2121);
and U1499 (N_1499,In_1112,In_1796);
and U1500 (N_1500,N_869,N_315);
nand U1501 (N_1501,N_1293,N_812);
or U1502 (N_1502,N_1274,N_875);
or U1503 (N_1503,N_48,N_239);
nand U1504 (N_1504,N_549,N_957);
and U1505 (N_1505,N_1211,N_660);
nor U1506 (N_1506,N_606,N_1305);
xnor U1507 (N_1507,N_510,N_1080);
or U1508 (N_1508,N_543,N_357);
and U1509 (N_1509,N_876,N_884);
and U1510 (N_1510,N_803,N_1038);
or U1511 (N_1511,N_777,N_1046);
and U1512 (N_1512,N_72,N_1434);
and U1513 (N_1513,N_1258,N_847);
or U1514 (N_1514,N_587,N_1150);
nand U1515 (N_1515,N_753,N_503);
nand U1516 (N_1516,N_711,N_1246);
and U1517 (N_1517,N_1403,N_976);
or U1518 (N_1518,N_0,N_1317);
and U1519 (N_1519,N_317,N_71);
nand U1520 (N_1520,N_52,N_313);
and U1521 (N_1521,N_1360,N_348);
xor U1522 (N_1522,N_681,N_1433);
nor U1523 (N_1523,N_915,N_894);
and U1524 (N_1524,N_7,N_1320);
nand U1525 (N_1525,N_1342,N_696);
nand U1526 (N_1526,N_1260,N_18);
and U1527 (N_1527,N_656,N_1435);
nand U1528 (N_1528,N_1271,N_1257);
and U1529 (N_1529,N_1102,N_1376);
or U1530 (N_1530,N_972,N_1371);
nand U1531 (N_1531,N_436,N_728);
nor U1532 (N_1532,N_330,N_1338);
or U1533 (N_1533,N_708,N_1157);
or U1534 (N_1534,N_163,N_1066);
or U1535 (N_1535,N_467,N_493);
nor U1536 (N_1536,N_987,N_598);
nand U1537 (N_1537,N_199,N_128);
or U1538 (N_1538,N_478,N_862);
nand U1539 (N_1539,N_588,N_505);
nand U1540 (N_1540,N_437,N_789);
and U1541 (N_1541,N_462,N_902);
or U1542 (N_1542,N_1440,N_557);
or U1543 (N_1543,N_1334,N_1057);
nand U1544 (N_1544,N_608,N_1343);
xor U1545 (N_1545,N_1365,N_565);
xnor U1546 (N_1546,N_887,N_912);
or U1547 (N_1547,N_1359,N_922);
nor U1548 (N_1548,N_146,N_1228);
nand U1549 (N_1549,N_1111,N_225);
xnor U1550 (N_1550,N_531,N_118);
nor U1551 (N_1551,N_817,N_1491);
and U1552 (N_1552,N_1350,N_1352);
or U1553 (N_1553,N_1424,N_794);
and U1554 (N_1554,N_202,N_1485);
or U1555 (N_1555,N_1286,N_102);
nand U1556 (N_1556,N_1421,N_1177);
nor U1557 (N_1557,N_204,N_1128);
or U1558 (N_1558,N_29,N_1105);
or U1559 (N_1559,N_104,N_953);
and U1560 (N_1560,N_157,N_1010);
and U1561 (N_1561,N_300,N_375);
xor U1562 (N_1562,N_558,N_126);
or U1563 (N_1563,N_756,N_1112);
nand U1564 (N_1564,N_535,N_734);
xnor U1565 (N_1565,N_729,N_779);
or U1566 (N_1566,N_270,N_672);
xnor U1567 (N_1567,N_1268,N_1234);
nor U1568 (N_1568,N_466,N_371);
nand U1569 (N_1569,N_217,N_476);
nand U1570 (N_1570,N_1070,N_1292);
nand U1571 (N_1571,N_422,N_715);
or U1572 (N_1572,N_230,N_122);
nor U1573 (N_1573,N_56,N_109);
and U1574 (N_1574,N_120,N_1156);
xnor U1575 (N_1575,N_627,N_27);
or U1576 (N_1576,N_295,N_1084);
or U1577 (N_1577,N_162,N_364);
xnor U1578 (N_1578,N_99,N_1461);
nand U1579 (N_1579,N_117,N_488);
nor U1580 (N_1580,N_964,N_1226);
nand U1581 (N_1581,N_1022,N_207);
nor U1582 (N_1582,N_1071,N_905);
nand U1583 (N_1583,N_489,N_1074);
or U1584 (N_1584,N_759,N_554);
and U1585 (N_1585,N_31,N_630);
and U1586 (N_1586,N_159,N_242);
nand U1587 (N_1587,N_917,N_5);
or U1588 (N_1588,N_487,N_358);
nand U1589 (N_1589,N_1129,N_444);
nand U1590 (N_1590,N_215,N_216);
xnor U1591 (N_1591,N_797,N_622);
nor U1592 (N_1592,N_890,N_1390);
and U1593 (N_1593,N_147,N_1396);
nand U1594 (N_1594,N_368,N_1470);
nand U1595 (N_1595,N_1155,N_405);
and U1596 (N_1596,N_267,N_433);
or U1597 (N_1597,N_552,N_465);
nand U1598 (N_1598,N_376,N_322);
or U1599 (N_1599,N_106,N_124);
xor U1600 (N_1600,N_1007,N_30);
and U1601 (N_1601,N_663,N_634);
nand U1602 (N_1602,N_604,N_423);
xnor U1603 (N_1603,N_25,N_1458);
nand U1604 (N_1604,N_1327,N_865);
and U1605 (N_1605,N_365,N_702);
and U1606 (N_1606,N_1487,N_572);
or U1607 (N_1607,N_463,N_509);
and U1608 (N_1608,N_1017,N_1459);
and U1609 (N_1609,N_1207,N_1197);
and U1610 (N_1610,N_1263,N_537);
and U1611 (N_1611,N_532,N_1291);
xnor U1612 (N_1612,N_1180,N_151);
or U1613 (N_1613,N_114,N_568);
nand U1614 (N_1614,N_200,N_757);
nand U1615 (N_1615,N_500,N_533);
and U1616 (N_1616,N_1230,N_539);
nand U1617 (N_1617,N_982,N_551);
nand U1618 (N_1618,N_1096,N_827);
xnor U1619 (N_1619,N_1166,N_1313);
nand U1620 (N_1620,N_567,N_281);
nand U1621 (N_1621,N_599,N_921);
nor U1622 (N_1622,N_1368,N_158);
and U1623 (N_1623,N_981,N_1452);
or U1624 (N_1624,N_1489,N_62);
nor U1625 (N_1625,N_440,N_282);
nand U1626 (N_1626,N_713,N_331);
and U1627 (N_1627,N_623,N_652);
nor U1628 (N_1628,N_1020,N_1418);
or U1629 (N_1629,N_635,N_1181);
or U1630 (N_1630,N_939,N_274);
nand U1631 (N_1631,N_195,N_805);
xnor U1632 (N_1632,N_137,N_188);
nand U1633 (N_1633,N_1040,N_996);
nand U1634 (N_1634,N_1450,N_787);
and U1635 (N_1635,N_798,N_990);
nand U1636 (N_1636,N_717,N_142);
or U1637 (N_1637,N_1205,N_1034);
or U1638 (N_1638,N_1321,N_522);
and U1639 (N_1639,N_534,N_859);
nor U1640 (N_1640,N_633,N_576);
or U1641 (N_1641,N_889,N_700);
nand U1642 (N_1642,N_1233,N_748);
xnor U1643 (N_1643,N_193,N_885);
xor U1644 (N_1644,N_473,N_457);
or U1645 (N_1645,N_1389,N_1428);
or U1646 (N_1646,N_886,N_924);
nor U1647 (N_1647,N_1044,N_946);
or U1648 (N_1648,N_1499,N_989);
or U1649 (N_1649,N_1179,N_666);
or U1650 (N_1650,N_942,N_143);
xnor U1651 (N_1651,N_1219,N_1358);
or U1652 (N_1652,N_1451,N_479);
or U1653 (N_1653,N_454,N_742);
or U1654 (N_1654,N_1134,N_998);
xor U1655 (N_1655,N_297,N_398);
and U1656 (N_1656,N_1152,N_910);
or U1657 (N_1657,N_625,N_832);
and U1658 (N_1658,N_545,N_1107);
nand U1659 (N_1659,N_1151,N_920);
nor U1660 (N_1660,N_1160,N_424);
nor U1661 (N_1661,N_1168,N_836);
nor U1662 (N_1662,N_373,N_825);
nand U1663 (N_1663,N_723,N_82);
nand U1664 (N_1664,N_718,N_716);
and U1665 (N_1665,N_1106,N_1138);
nor U1666 (N_1666,N_712,N_302);
nand U1667 (N_1667,N_764,N_95);
xor U1668 (N_1668,N_1063,N_1280);
or U1669 (N_1669,N_888,N_196);
nor U1670 (N_1670,N_309,N_526);
and U1671 (N_1671,N_1273,N_1486);
xor U1672 (N_1672,N_1279,N_1462);
nand U1673 (N_1673,N_1484,N_1130);
and U1674 (N_1674,N_645,N_1131);
nand U1675 (N_1675,N_596,N_1231);
and U1676 (N_1676,N_471,N_932);
or U1677 (N_1677,N_737,N_1182);
or U1678 (N_1678,N_359,N_1079);
nand U1679 (N_1679,N_342,N_513);
and U1680 (N_1680,N_459,N_1149);
or U1681 (N_1681,N_1314,N_1185);
nor U1682 (N_1682,N_1319,N_192);
and U1683 (N_1683,N_1229,N_388);
and U1684 (N_1684,N_291,N_1052);
nand U1685 (N_1685,N_321,N_1206);
xor U1686 (N_1686,N_1032,N_928);
nor U1687 (N_1687,N_1266,N_1223);
and U1688 (N_1688,N_1409,N_1097);
or U1689 (N_1689,N_840,N_1221);
nand U1690 (N_1690,N_977,N_863);
nand U1691 (N_1691,N_986,N_307);
nand U1692 (N_1692,N_907,N_582);
nor U1693 (N_1693,N_1239,N_324);
or U1694 (N_1694,N_186,N_272);
and U1695 (N_1695,N_592,N_1361);
nor U1696 (N_1696,N_67,N_1391);
xnor U1697 (N_1697,N_450,N_39);
and U1698 (N_1698,N_1225,N_853);
or U1699 (N_1699,N_1113,N_822);
nor U1700 (N_1700,N_265,N_900);
xor U1701 (N_1701,N_741,N_185);
or U1702 (N_1702,N_59,N_133);
and U1703 (N_1703,N_1411,N_175);
nor U1704 (N_1704,N_1460,N_129);
and U1705 (N_1705,N_1384,N_1426);
xnor U1706 (N_1706,N_941,N_1000);
nand U1707 (N_1707,N_835,N_439);
xnor U1708 (N_1708,N_895,N_1423);
nand U1709 (N_1709,N_994,N_969);
nor U1710 (N_1710,N_1407,N_516);
nand U1711 (N_1711,N_332,N_36);
and U1712 (N_1712,N_447,N_721);
nand U1713 (N_1713,N_1090,N_1457);
and U1714 (N_1714,N_451,N_856);
nand U1715 (N_1715,N_542,N_394);
xor U1716 (N_1716,N_1132,N_289);
nand U1717 (N_1717,N_1165,N_738);
xor U1718 (N_1718,N_1146,N_937);
nand U1719 (N_1719,N_1029,N_481);
or U1720 (N_1720,N_792,N_893);
nand U1721 (N_1721,N_1203,N_1100);
nor U1722 (N_1722,N_1495,N_287);
and U1723 (N_1723,N_949,N_1255);
xor U1724 (N_1724,N_1023,N_1159);
and U1725 (N_1725,N_130,N_1043);
nand U1726 (N_1726,N_775,N_233);
and U1727 (N_1727,N_821,N_1281);
or U1728 (N_1728,N_670,N_1312);
or U1729 (N_1729,N_768,N_1171);
or U1730 (N_1730,N_898,N_40);
nor U1731 (N_1731,N_1088,N_1250);
xor U1732 (N_1732,N_148,N_10);
nand U1733 (N_1733,N_1340,N_303);
or U1734 (N_1734,N_24,N_897);
nand U1735 (N_1735,N_1235,N_418);
xor U1736 (N_1736,N_564,N_784);
and U1737 (N_1737,N_257,N_1133);
xnor U1738 (N_1738,N_201,N_1099);
and U1739 (N_1739,N_134,N_569);
xor U1740 (N_1740,N_44,N_349);
or U1741 (N_1741,N_1008,N_38);
and U1742 (N_1742,N_399,N_94);
nand U1743 (N_1743,N_92,N_1215);
nand U1744 (N_1744,N_1049,N_1476);
and U1745 (N_1745,N_563,N_908);
or U1746 (N_1746,N_494,N_793);
xor U1747 (N_1747,N_1363,N_212);
and U1748 (N_1748,N_570,N_732);
nor U1749 (N_1749,N_919,N_690);
and U1750 (N_1750,N_879,N_662);
xor U1751 (N_1751,N_786,N_527);
nor U1752 (N_1752,N_1309,N_745);
xnor U1753 (N_1753,N_801,N_584);
nand U1754 (N_1754,N_26,N_766);
xor U1755 (N_1755,N_618,N_385);
or U1756 (N_1756,N_947,N_621);
nor U1757 (N_1757,N_1011,N_54);
xnor U1758 (N_1758,N_1075,N_640);
xor U1759 (N_1759,N_1441,N_308);
xor U1760 (N_1760,N_452,N_1158);
and U1761 (N_1761,N_55,N_1037);
xnor U1762 (N_1762,N_968,N_173);
and U1763 (N_1763,N_88,N_1101);
nand U1764 (N_1764,N_1078,N_111);
nor U1765 (N_1765,N_783,N_1035);
nand U1766 (N_1766,N_286,N_773);
nor U1767 (N_1767,N_1393,N_284);
or U1768 (N_1768,N_1209,N_538);
nor U1769 (N_1769,N_860,N_425);
nand U1770 (N_1770,N_442,N_579);
nor U1771 (N_1771,N_19,N_566);
nor U1772 (N_1772,N_746,N_160);
nand U1773 (N_1773,N_639,N_1253);
nand U1774 (N_1774,N_1399,N_730);
xnor U1775 (N_1775,N_1265,N_1167);
or U1776 (N_1776,N_1238,N_704);
nor U1777 (N_1777,N_562,N_273);
and U1778 (N_1778,N_1392,N_1194);
and U1779 (N_1779,N_555,N_1013);
nor U1780 (N_1780,N_1410,N_400);
and U1781 (N_1781,N_410,N_791);
and U1782 (N_1782,N_1061,N_203);
or U1783 (N_1783,N_1243,N_1304);
or U1784 (N_1784,N_844,N_416);
xor U1785 (N_1785,N_892,N_1042);
xnor U1786 (N_1786,N_1222,N_1184);
nor U1787 (N_1787,N_1076,N_991);
nor U1788 (N_1788,N_1148,N_1269);
and U1789 (N_1789,N_1432,N_432);
xor U1790 (N_1790,N_1251,N_682);
and U1791 (N_1791,N_316,N_508);
xor U1792 (N_1792,N_641,N_1244);
xor U1793 (N_1793,N_1115,N_586);
xnor U1794 (N_1794,N_170,N_1296);
nor U1795 (N_1795,N_1436,N_736);
nor U1796 (N_1796,N_49,N_854);
or U1797 (N_1797,N_430,N_218);
or U1798 (N_1798,N_1164,N_1357);
nand U1799 (N_1799,N_98,N_387);
and U1800 (N_1800,N_268,N_1287);
xnor U1801 (N_1801,N_81,N_1439);
and U1802 (N_1802,N_1086,N_119);
or U1803 (N_1803,N_1002,N_809);
or U1804 (N_1804,N_664,N_115);
xor U1805 (N_1805,N_1416,N_988);
xor U1806 (N_1806,N_41,N_1443);
nand U1807 (N_1807,N_1375,N_253);
nor U1808 (N_1808,N_395,N_918);
nor U1809 (N_1809,N_413,N_849);
nor U1810 (N_1810,N_680,N_156);
nor U1811 (N_1811,N_352,N_8);
xor U1812 (N_1812,N_356,N_1103);
nand U1813 (N_1813,N_610,N_426);
nand U1814 (N_1814,N_1387,N_731);
and U1815 (N_1815,N_210,N_389);
nand U1816 (N_1816,N_1003,N_1329);
nand U1817 (N_1817,N_1475,N_1366);
nor U1818 (N_1818,N_278,N_1082);
nor U1819 (N_1819,N_758,N_1204);
nand U1820 (N_1820,N_259,N_765);
nor U1821 (N_1821,N_34,N_1404);
xor U1822 (N_1822,N_1402,N_280);
nor U1823 (N_1823,N_392,N_420);
nand U1824 (N_1824,N_524,N_149);
xnor U1825 (N_1825,N_402,N_1298);
nand U1826 (N_1826,N_11,N_927);
or U1827 (N_1827,N_1142,N_396);
xnor U1828 (N_1828,N_880,N_100);
nor U1829 (N_1829,N_1333,N_1009);
nand U1830 (N_1830,N_227,N_699);
xor U1831 (N_1831,N_589,N_1483);
and U1832 (N_1832,N_751,N_518);
or U1833 (N_1833,N_811,N_1069);
nor U1834 (N_1834,N_1021,N_153);
nand U1835 (N_1835,N_1378,N_112);
xnor U1836 (N_1836,N_829,N_57);
or U1837 (N_1837,N_950,N_523);
nor U1838 (N_1838,N_429,N_1162);
nand U1839 (N_1839,N_1062,N_978);
xnor U1840 (N_1840,N_1153,N_914);
xnor U1841 (N_1841,N_1245,N_1473);
nor U1842 (N_1842,N_602,N_370);
and U1843 (N_1843,N_179,N_1444);
xor U1844 (N_1844,N_979,N_1144);
or U1845 (N_1845,N_512,N_1449);
nand U1846 (N_1846,N_810,N_1303);
nand U1847 (N_1847,N_261,N_826);
or U1848 (N_1848,N_1218,N_601);
nor U1849 (N_1849,N_1001,N_823);
nand U1850 (N_1850,N_675,N_279);
xnor U1851 (N_1851,N_658,N_483);
xnor U1852 (N_1852,N_245,N_896);
nand U1853 (N_1853,N_644,N_1122);
nor U1854 (N_1854,N_28,N_674);
xnor U1855 (N_1855,N_161,N_726);
and U1856 (N_1856,N_1455,N_1172);
and U1857 (N_1857,N_1469,N_382);
or U1858 (N_1858,N_852,N_288);
xor U1859 (N_1859,N_310,N_511);
nor U1860 (N_1860,N_911,N_1004);
nand U1861 (N_1861,N_930,N_69);
xnor U1862 (N_1862,N_1060,N_1104);
or U1863 (N_1863,N_340,N_1417);
nand U1864 (N_1864,N_1379,N_616);
xnor U1865 (N_1865,N_577,N_497);
or U1866 (N_1866,N_181,N_66);
and U1867 (N_1867,N_266,N_35);
and U1868 (N_1868,N_677,N_1195);
nor U1869 (N_1869,N_714,N_1412);
nor U1870 (N_1870,N_1200,N_850);
and U1871 (N_1871,N_653,N_472);
nor U1872 (N_1872,N_956,N_1341);
nor U1873 (N_1873,N_255,N_206);
xor U1874 (N_1874,N_1169,N_1326);
and U1875 (N_1875,N_1154,N_529);
nand U1876 (N_1876,N_1118,N_632);
nor U1877 (N_1877,N_727,N_933);
or U1878 (N_1878,N_150,N_1479);
nor U1879 (N_1879,N_325,N_857);
or U1880 (N_1880,N_1490,N_431);
nand U1881 (N_1881,N_1064,N_458);
nand U1882 (N_1882,N_1488,N_1249);
xor U1883 (N_1883,N_830,N_776);
and U1884 (N_1884,N_269,N_1300);
or U1885 (N_1885,N_241,N_1247);
nor U1886 (N_1886,N_1224,N_406);
xor U1887 (N_1887,N_695,N_232);
nor U1888 (N_1888,N_2,N_299);
or U1889 (N_1889,N_1331,N_1496);
nor U1890 (N_1890,N_1237,N_1302);
nor U1891 (N_1891,N_1477,N_1285);
nor U1892 (N_1892,N_1398,N_1236);
nor U1893 (N_1893,N_834,N_305);
or U1894 (N_1894,N_390,N_995);
xor U1895 (N_1895,N_999,N_53);
xor U1896 (N_1896,N_848,N_223);
and U1897 (N_1897,N_899,N_1447);
and U1898 (N_1898,N_744,N_1137);
nor U1899 (N_1899,N_254,N_1147);
xor U1900 (N_1900,N_103,N_14);
and U1901 (N_1901,N_294,N_1031);
or U1902 (N_1902,N_1039,N_1463);
nand U1903 (N_1903,N_1311,N_1337);
and U1904 (N_1904,N_993,N_362);
and U1905 (N_1905,N_1126,N_724);
nor U1906 (N_1906,N_83,N_818);
or U1907 (N_1907,N_593,N_1098);
nand U1908 (N_1908,N_407,N_1119);
or U1909 (N_1909,N_1033,N_1380);
nand U1910 (N_1910,N_446,N_397);
xor U1911 (N_1911,N_971,N_1308);
xnor U1912 (N_1912,N_460,N_314);
xor U1913 (N_1913,N_747,N_631);
xnor U1914 (N_1914,N_1307,N_845);
xnor U1915 (N_1915,N_329,N_417);
and U1916 (N_1916,N_131,N_578);
and U1917 (N_1917,N_248,N_1494);
xnor U1918 (N_1918,N_60,N_614);
or U1919 (N_1919,N_229,N_461);
and U1920 (N_1920,N_1026,N_354);
nor U1921 (N_1921,N_1109,N_45);
xnor U1922 (N_1922,N_17,N_401);
or U1923 (N_1923,N_1498,N_1466);
and U1924 (N_1924,N_581,N_689);
nand U1925 (N_1925,N_943,N_962);
nor U1926 (N_1926,N_182,N_1383);
or U1927 (N_1927,N_228,N_1216);
nand U1928 (N_1928,N_867,N_750);
and U1929 (N_1929,N_781,N_141);
nor U1930 (N_1930,N_948,N_1425);
xor U1931 (N_1931,N_221,N_209);
nand U1932 (N_1932,N_1056,N_683);
and U1933 (N_1933,N_575,N_292);
nand U1934 (N_1934,N_763,N_64);
nand U1935 (N_1935,N_363,N_403);
or U1936 (N_1936,N_719,N_251);
xor U1937 (N_1937,N_1089,N_624);
and U1938 (N_1938,N_1480,N_1478);
xor U1939 (N_1939,N_468,N_760);
and U1940 (N_1940,N_1186,N_1430);
nor U1941 (N_1941,N_553,N_136);
or U1942 (N_1942,N_33,N_1045);
or U1943 (N_1943,N_165,N_46);
or U1944 (N_1944,N_1429,N_1370);
nor U1945 (N_1945,N_1356,N_983);
or U1946 (N_1946,N_521,N_164);
nor U1947 (N_1947,N_1306,N_344);
nor U1948 (N_1948,N_620,N_506);
or U1949 (N_1949,N_37,N_68);
nor U1950 (N_1950,N_603,N_219);
and U1951 (N_1951,N_796,N_1065);
nor U1952 (N_1952,N_372,N_694);
nor U1953 (N_1953,N_76,N_722);
nand U1954 (N_1954,N_89,N_1114);
nor U1955 (N_1955,N_247,N_380);
xor U1956 (N_1956,N_32,N_168);
nand U1957 (N_1957,N_813,N_1068);
and U1958 (N_1958,N_491,N_184);
and U1959 (N_1959,N_484,N_108);
and U1960 (N_1960,N_1217,N_367);
or U1961 (N_1961,N_679,N_1220);
xnor U1962 (N_1962,N_123,N_1339);
or U1963 (N_1963,N_1212,N_263);
or U1964 (N_1964,N_1136,N_561);
or U1965 (N_1965,N_1014,N_1427);
xnor U1966 (N_1966,N_613,N_965);
nor U1967 (N_1967,N_1362,N_1170);
nand U1968 (N_1968,N_1214,N_1272);
or U1969 (N_1969,N_246,N_1369);
nand U1970 (N_1970,N_421,N_1406);
nor U1971 (N_1971,N_668,N_492);
nand U1972 (N_1972,N_1335,N_877);
xnor U1973 (N_1973,N_1240,N_767);
nor U1974 (N_1974,N_936,N_1005);
and U1975 (N_1975,N_720,N_1242);
and U1976 (N_1976,N_1422,N_311);
nor U1977 (N_1977,N_1213,N_550);
or U1978 (N_1978,N_409,N_1019);
nand U1979 (N_1979,N_1227,N_480);
and U1980 (N_1980,N_654,N_1454);
nand U1981 (N_1981,N_617,N_1067);
or U1982 (N_1982,N_871,N_967);
nor U1983 (N_1983,N_138,N_772);
nor U1984 (N_1984,N_778,N_183);
nand U1985 (N_1985,N_1054,N_1353);
and U1986 (N_1986,N_1453,N_328);
or U1987 (N_1987,N_691,N_501);
and U1988 (N_1988,N_1108,N_698);
and U1989 (N_1989,N_1058,N_1275);
nand U1990 (N_1990,N_445,N_1301);
or U1991 (N_1991,N_113,N_975);
xnor U1992 (N_1992,N_20,N_252);
xnor U1993 (N_1993,N_327,N_612);
nand U1994 (N_1994,N_1474,N_125);
or U1995 (N_1995,N_966,N_960);
nand U1996 (N_1996,N_1413,N_600);
and U1997 (N_1997,N_774,N_735);
xor U1998 (N_1998,N_205,N_846);
xor U1999 (N_1999,N_815,N_951);
nand U2000 (N_2000,N_298,N_546);
nand U2001 (N_2001,N_336,N_408);
or U2002 (N_2002,N_1201,N_455);
xor U2003 (N_2003,N_301,N_642);
or U2004 (N_2004,N_96,N_350);
or U2005 (N_2005,N_180,N_1318);
nor U2006 (N_2006,N_1085,N_944);
or U2007 (N_2007,N_337,N_673);
nand U2008 (N_2008,N_547,N_235);
xor U2009 (N_2009,N_304,N_1471);
or U2010 (N_2010,N_9,N_955);
nor U2011 (N_2011,N_761,N_13);
or U2012 (N_2012,N_1355,N_121);
or U2013 (N_2013,N_178,N_1264);
nand U2014 (N_2014,N_1414,N_619);
nor U2015 (N_2015,N_1140,N_1161);
or U2016 (N_2016,N_1123,N_739);
nor U2017 (N_2017,N_667,N_1394);
nand U2018 (N_2018,N_1232,N_75);
or U2019 (N_2019,N_1431,N_23);
and U2020 (N_2020,N_323,N_434);
nand U2021 (N_2021,N_499,N_688);
nor U2022 (N_2022,N_819,N_980);
and U2023 (N_2023,N_1482,N_482);
and U2024 (N_2024,N_244,N_1497);
nand U2025 (N_2025,N_271,N_50);
xor U2026 (N_2026,N_780,N_636);
and U2027 (N_2027,N_140,N_486);
or U2028 (N_2028,N_290,N_70);
xnor U2029 (N_2029,N_954,N_1016);
and U2030 (N_2030,N_671,N_293);
and U2031 (N_2031,N_1288,N_906);
or U2032 (N_2032,N_646,N_843);
nor U2033 (N_2033,N_1322,N_974);
and U2034 (N_2034,N_1377,N_306);
xnor U2035 (N_2035,N_684,N_243);
nand U2036 (N_2036,N_1467,N_1006);
nand U2037 (N_2037,N_1120,N_1053);
nor U2038 (N_2038,N_1256,N_1187);
or U2039 (N_2039,N_934,N_961);
or U2040 (N_2040,N_238,N_1262);
xnor U2041 (N_2041,N_116,N_1178);
xnor U2042 (N_2042,N_609,N_507);
or U2043 (N_2043,N_909,N_1041);
xor U2044 (N_2044,N_105,N_992);
and U2045 (N_2045,N_1437,N_790);
and U2046 (N_2046,N_1401,N_441);
and U2047 (N_2047,N_1139,N_498);
nand U2048 (N_2048,N_709,N_63);
nand U2049 (N_2049,N_277,N_958);
or U2050 (N_2050,N_1289,N_913);
or U2051 (N_2051,N_1027,N_1192);
nand U2052 (N_2052,N_172,N_1199);
xor U2053 (N_2053,N_851,N_237);
or U2054 (N_2054,N_800,N_814);
or U2055 (N_2055,N_374,N_743);
xnor U2056 (N_2056,N_47,N_806);
nor U2057 (N_2057,N_1092,N_864);
xnor U2058 (N_2058,N_580,N_339);
nor U2059 (N_2059,N_970,N_167);
nor U2060 (N_2060,N_931,N_548);
or U2061 (N_2061,N_1254,N_807);
nor U2062 (N_2062,N_615,N_657);
xnor U2063 (N_2063,N_187,N_1330);
nor U2064 (N_2064,N_1083,N_214);
nor U2065 (N_2065,N_256,N_377);
xor U2066 (N_2066,N_1198,N_1174);
or U2067 (N_2067,N_449,N_540);
nand U2068 (N_2068,N_91,N_456);
nor U2069 (N_2069,N_882,N_1316);
and U2070 (N_2070,N_1493,N_366);
nor U2071 (N_2071,N_171,N_1278);
nand U2072 (N_2072,N_762,N_1252);
nor U2073 (N_2073,N_296,N_648);
xor U2074 (N_2074,N_504,N_1382);
nor U2075 (N_2075,N_595,N_938);
nor U2076 (N_2076,N_379,N_144);
and U2077 (N_2077,N_1468,N_1191);
and U2078 (N_2078,N_669,N_984);
and U2079 (N_2079,N_1297,N_785);
and U2080 (N_2080,N_701,N_264);
or U2081 (N_2081,N_404,N_831);
or U2082 (N_2082,N_355,N_393);
and U2083 (N_2083,N_517,N_883);
and U2084 (N_2084,N_923,N_872);
xnor U2085 (N_2085,N_378,N_275);
and U2086 (N_2086,N_594,N_1442);
nand U2087 (N_2087,N_904,N_226);
nor U2088 (N_2088,N_16,N_661);
nand U2089 (N_2089,N_1445,N_1028);
nor U2090 (N_2090,N_85,N_496);
nand U2091 (N_2091,N_191,N_234);
or U2092 (N_2092,N_929,N_222);
nor U2093 (N_2093,N_107,N_353);
or U2094 (N_2094,N_590,N_525);
nand U2095 (N_2095,N_249,N_319);
xor U2096 (N_2096,N_1176,N_1055);
nor U2097 (N_2097,N_1270,N_692);
nor U2098 (N_2098,N_51,N_665);
and U2099 (N_2099,N_369,N_655);
xnor U2100 (N_2100,N_1284,N_1124);
or U2101 (N_2101,N_176,N_515);
or U2102 (N_2102,N_84,N_749);
or U2103 (N_2103,N_1295,N_1464);
nand U2104 (N_2104,N_1354,N_1091);
xnor U2105 (N_2105,N_1397,N_1492);
and U2106 (N_2106,N_502,N_448);
nand U2107 (N_2107,N_833,N_607);
or U2108 (N_2108,N_1081,N_15);
nand U2109 (N_2109,N_1408,N_326);
and U2110 (N_2110,N_345,N_475);
xor U2111 (N_2111,N_190,N_412);
or U2112 (N_2112,N_1420,N_676);
nor U2113 (N_2113,N_725,N_769);
nand U2114 (N_2114,N_470,N_1290);
nand U2115 (N_2115,N_360,N_231);
or U2116 (N_2116,N_583,N_795);
or U2117 (N_2117,N_649,N_152);
and U2118 (N_2118,N_87,N_65);
or U2119 (N_2119,N_1351,N_1135);
or U2120 (N_2120,N_771,N_571);
and U2121 (N_2121,N_985,N_629);
nand U2122 (N_2122,N_428,N_560);
nand U2123 (N_2123,N_1419,N_343);
or U2124 (N_2124,N_643,N_870);
xor U2125 (N_2125,N_1283,N_816);
or U2126 (N_2126,N_520,N_1125);
nand U2127 (N_2127,N_419,N_707);
and U2128 (N_2128,N_1036,N_1294);
nand U2129 (N_2129,N_1015,N_1323);
or U2130 (N_2130,N_194,N_820);
nand U2131 (N_2131,N_997,N_808);
xnor U2132 (N_2132,N_438,N_464);
nand U2133 (N_2133,N_1087,N_443);
nor U2134 (N_2134,N_1388,N_647);
and U2135 (N_2135,N_338,N_1299);
or U2136 (N_2136,N_1095,N_127);
or U2137 (N_2137,N_1047,N_211);
or U2138 (N_2138,N_628,N_536);
and U2139 (N_2139,N_1241,N_935);
nand U2140 (N_2140,N_386,N_333);
xnor U2141 (N_2141,N_1117,N_110);
or U2142 (N_2142,N_903,N_1324);
or U2143 (N_2143,N_1077,N_1093);
nand U2144 (N_2144,N_611,N_901);
xor U2145 (N_2145,N_1415,N_208);
nand U2146 (N_2146,N_1094,N_959);
or U2147 (N_2147,N_706,N_693);
or U2148 (N_2148,N_1059,N_651);
or U2149 (N_2149,N_637,N_1051);
nor U2150 (N_2150,N_58,N_155);
and U2151 (N_2151,N_320,N_236);
nand U2152 (N_2152,N_782,N_838);
nor U2153 (N_2153,N_858,N_42);
nor U2154 (N_2154,N_1344,N_101);
xnor U2155 (N_2155,N_1348,N_250);
and U2156 (N_2156,N_139,N_740);
nor U2157 (N_2157,N_427,N_469);
or U2158 (N_2158,N_1018,N_1189);
xnor U2159 (N_2159,N_837,N_1282);
nand U2160 (N_2160,N_1395,N_659);
and U2161 (N_2161,N_78,N_1175);
nand U2162 (N_2162,N_1190,N_1405);
nor U2163 (N_2163,N_1141,N_855);
or U2164 (N_2164,N_1030,N_559);
and U2165 (N_2165,N_240,N_73);
or U2166 (N_2166,N_154,N_891);
or U2167 (N_2167,N_262,N_145);
and U2168 (N_2168,N_973,N_519);
nor U2169 (N_2169,N_346,N_415);
and U2170 (N_2170,N_485,N_61);
or U2171 (N_2171,N_952,N_1267);
or U2172 (N_2172,N_4,N_1110);
nand U2173 (N_2173,N_1364,N_1347);
xnor U2174 (N_2174,N_585,N_1367);
and U2175 (N_2175,N_1196,N_1073);
or U2176 (N_2176,N_1,N_414);
nor U2177 (N_2177,N_1193,N_945);
xnor U2178 (N_2178,N_80,N_1386);
and U2179 (N_2179,N_132,N_703);
nor U2180 (N_2180,N_687,N_312);
or U2181 (N_2181,N_1373,N_318);
nor U2182 (N_2182,N_1208,N_1202);
xor U2183 (N_2183,N_285,N_874);
xor U2184 (N_2184,N_381,N_1183);
xnor U2185 (N_2185,N_605,N_43);
nand U2186 (N_2186,N_334,N_490);
xnor U2187 (N_2187,N_733,N_541);
nand U2188 (N_2188,N_514,N_283);
nor U2189 (N_2189,N_1116,N_866);
and U2190 (N_2190,N_1188,N_1336);
and U2191 (N_2191,N_828,N_90);
xnor U2192 (N_2192,N_1332,N_788);
xnor U2193 (N_2193,N_754,N_341);
nor U2194 (N_2194,N_213,N_224);
nor U2195 (N_2195,N_1048,N_804);
and U2196 (N_2196,N_1448,N_22);
nor U2197 (N_2197,N_1248,N_1261);
or U2198 (N_2198,N_705,N_1127);
or U2199 (N_2199,N_335,N_678);
nor U2200 (N_2200,N_435,N_411);
xnor U2201 (N_2201,N_351,N_1024);
or U2202 (N_2202,N_6,N_474);
xnor U2203 (N_2203,N_530,N_1315);
xnor U2204 (N_2204,N_79,N_963);
and U2205 (N_2205,N_1121,N_925);
nand U2206 (N_2206,N_12,N_1346);
nor U2207 (N_2207,N_574,N_1349);
nand U2208 (N_2208,N_1374,N_74);
nand U2209 (N_2209,N_1372,N_868);
nor U2210 (N_2210,N_544,N_1163);
nor U2211 (N_2211,N_1259,N_1143);
nand U2212 (N_2212,N_802,N_86);
nand U2213 (N_2213,N_495,N_169);
nor U2214 (N_2214,N_174,N_3);
nand U2215 (N_2215,N_1210,N_347);
nand U2216 (N_2216,N_697,N_198);
xnor U2217 (N_2217,N_1465,N_638);
or U2218 (N_2218,N_166,N_220);
or U2219 (N_2219,N_770,N_799);
or U2220 (N_2220,N_916,N_626);
and U2221 (N_2221,N_650,N_1446);
or U2222 (N_2222,N_528,N_841);
and U2223 (N_2223,N_1276,N_710);
nand U2224 (N_2224,N_135,N_556);
nor U2225 (N_2225,N_1481,N_1072);
xnor U2226 (N_2226,N_1381,N_1310);
and U2227 (N_2227,N_1456,N_361);
and U2228 (N_2228,N_177,N_477);
or U2229 (N_2229,N_573,N_873);
and U2230 (N_2230,N_881,N_1400);
nand U2231 (N_2231,N_276,N_189);
and U2232 (N_2232,N_597,N_453);
or U2233 (N_2233,N_752,N_1472);
and U2234 (N_2234,N_21,N_755);
nor U2235 (N_2235,N_686,N_1277);
nor U2236 (N_2236,N_685,N_77);
nand U2237 (N_2237,N_1173,N_391);
nand U2238 (N_2238,N_878,N_197);
nand U2239 (N_2239,N_1050,N_258);
nand U2240 (N_2240,N_93,N_824);
xor U2241 (N_2241,N_383,N_384);
nor U2242 (N_2242,N_260,N_97);
xor U2243 (N_2243,N_1025,N_940);
nand U2244 (N_2244,N_1345,N_842);
or U2245 (N_2245,N_861,N_926);
xor U2246 (N_2246,N_1012,N_1328);
nor U2247 (N_2247,N_839,N_1438);
nand U2248 (N_2248,N_1385,N_1325);
and U2249 (N_2249,N_1145,N_591);
and U2250 (N_2250,N_719,N_283);
xnor U2251 (N_2251,N_539,N_318);
xor U2252 (N_2252,N_161,N_1181);
nand U2253 (N_2253,N_990,N_1347);
nor U2254 (N_2254,N_1343,N_1118);
nand U2255 (N_2255,N_408,N_552);
nor U2256 (N_2256,N_715,N_953);
and U2257 (N_2257,N_829,N_530);
or U2258 (N_2258,N_469,N_917);
xor U2259 (N_2259,N_429,N_1418);
or U2260 (N_2260,N_296,N_590);
xor U2261 (N_2261,N_378,N_282);
nand U2262 (N_2262,N_1121,N_577);
nor U2263 (N_2263,N_453,N_686);
or U2264 (N_2264,N_1052,N_248);
and U2265 (N_2265,N_589,N_1361);
nor U2266 (N_2266,N_1452,N_1278);
or U2267 (N_2267,N_445,N_1275);
and U2268 (N_2268,N_841,N_566);
xnor U2269 (N_2269,N_877,N_989);
xor U2270 (N_2270,N_69,N_1016);
or U2271 (N_2271,N_33,N_377);
xnor U2272 (N_2272,N_1247,N_22);
nand U2273 (N_2273,N_738,N_829);
and U2274 (N_2274,N_56,N_112);
or U2275 (N_2275,N_1390,N_79);
nor U2276 (N_2276,N_1053,N_623);
xor U2277 (N_2277,N_1060,N_392);
or U2278 (N_2278,N_1331,N_915);
and U2279 (N_2279,N_569,N_1192);
nand U2280 (N_2280,N_1428,N_324);
xor U2281 (N_2281,N_839,N_284);
nor U2282 (N_2282,N_1415,N_1479);
xnor U2283 (N_2283,N_1259,N_1174);
nand U2284 (N_2284,N_1349,N_344);
nand U2285 (N_2285,N_1307,N_91);
and U2286 (N_2286,N_471,N_1221);
nand U2287 (N_2287,N_1411,N_678);
nor U2288 (N_2288,N_1373,N_953);
nor U2289 (N_2289,N_853,N_267);
xnor U2290 (N_2290,N_1452,N_324);
nor U2291 (N_2291,N_1409,N_1056);
xnor U2292 (N_2292,N_912,N_866);
and U2293 (N_2293,N_423,N_1330);
nor U2294 (N_2294,N_809,N_442);
nand U2295 (N_2295,N_797,N_1257);
or U2296 (N_2296,N_842,N_677);
xnor U2297 (N_2297,N_1047,N_277);
and U2298 (N_2298,N_838,N_1215);
nor U2299 (N_2299,N_327,N_1052);
nor U2300 (N_2300,N_285,N_483);
nor U2301 (N_2301,N_883,N_547);
nor U2302 (N_2302,N_1317,N_895);
and U2303 (N_2303,N_368,N_1365);
or U2304 (N_2304,N_291,N_1443);
or U2305 (N_2305,N_1096,N_391);
or U2306 (N_2306,N_451,N_976);
and U2307 (N_2307,N_1207,N_750);
or U2308 (N_2308,N_990,N_1466);
nand U2309 (N_2309,N_578,N_1296);
nor U2310 (N_2310,N_463,N_1047);
or U2311 (N_2311,N_308,N_1406);
or U2312 (N_2312,N_1360,N_1270);
xnor U2313 (N_2313,N_1483,N_1434);
nor U2314 (N_2314,N_1358,N_731);
and U2315 (N_2315,N_1475,N_1373);
and U2316 (N_2316,N_27,N_1347);
nand U2317 (N_2317,N_1407,N_874);
xor U2318 (N_2318,N_1406,N_980);
or U2319 (N_2319,N_904,N_1164);
nand U2320 (N_2320,N_208,N_867);
nor U2321 (N_2321,N_112,N_9);
xor U2322 (N_2322,N_1318,N_219);
nor U2323 (N_2323,N_184,N_792);
and U2324 (N_2324,N_71,N_1129);
xnor U2325 (N_2325,N_361,N_66);
nand U2326 (N_2326,N_733,N_369);
and U2327 (N_2327,N_1490,N_357);
nand U2328 (N_2328,N_165,N_1441);
xor U2329 (N_2329,N_1377,N_1410);
nand U2330 (N_2330,N_124,N_1296);
xor U2331 (N_2331,N_651,N_437);
nor U2332 (N_2332,N_951,N_1394);
xor U2333 (N_2333,N_182,N_665);
and U2334 (N_2334,N_1200,N_987);
and U2335 (N_2335,N_1012,N_472);
nor U2336 (N_2336,N_435,N_1414);
or U2337 (N_2337,N_45,N_250);
nor U2338 (N_2338,N_328,N_1282);
xnor U2339 (N_2339,N_1392,N_1124);
xnor U2340 (N_2340,N_1301,N_395);
and U2341 (N_2341,N_1364,N_51);
or U2342 (N_2342,N_1339,N_247);
or U2343 (N_2343,N_1196,N_1135);
nand U2344 (N_2344,N_690,N_1276);
xor U2345 (N_2345,N_1050,N_205);
nor U2346 (N_2346,N_418,N_30);
nor U2347 (N_2347,N_221,N_597);
nand U2348 (N_2348,N_276,N_920);
and U2349 (N_2349,N_690,N_563);
nor U2350 (N_2350,N_339,N_554);
nand U2351 (N_2351,N_835,N_954);
and U2352 (N_2352,N_946,N_661);
xnor U2353 (N_2353,N_360,N_1042);
nand U2354 (N_2354,N_397,N_1087);
and U2355 (N_2355,N_45,N_105);
nand U2356 (N_2356,N_694,N_466);
xor U2357 (N_2357,N_507,N_1357);
nand U2358 (N_2358,N_1443,N_422);
nor U2359 (N_2359,N_83,N_1198);
and U2360 (N_2360,N_1109,N_69);
nand U2361 (N_2361,N_1395,N_538);
nor U2362 (N_2362,N_926,N_1138);
or U2363 (N_2363,N_690,N_754);
or U2364 (N_2364,N_1443,N_921);
or U2365 (N_2365,N_486,N_1355);
xnor U2366 (N_2366,N_1364,N_115);
xor U2367 (N_2367,N_837,N_730);
xnor U2368 (N_2368,N_1451,N_250);
and U2369 (N_2369,N_1144,N_1137);
and U2370 (N_2370,N_69,N_695);
nand U2371 (N_2371,N_764,N_948);
nand U2372 (N_2372,N_1479,N_99);
nor U2373 (N_2373,N_996,N_816);
or U2374 (N_2374,N_741,N_1331);
nor U2375 (N_2375,N_1486,N_1003);
and U2376 (N_2376,N_864,N_938);
or U2377 (N_2377,N_1287,N_856);
and U2378 (N_2378,N_1495,N_113);
xor U2379 (N_2379,N_362,N_752);
nand U2380 (N_2380,N_1309,N_727);
or U2381 (N_2381,N_630,N_1072);
nor U2382 (N_2382,N_853,N_1066);
nand U2383 (N_2383,N_1126,N_1115);
xnor U2384 (N_2384,N_955,N_1441);
or U2385 (N_2385,N_502,N_1386);
nor U2386 (N_2386,N_1210,N_770);
and U2387 (N_2387,N_687,N_648);
and U2388 (N_2388,N_95,N_1391);
nand U2389 (N_2389,N_667,N_980);
nand U2390 (N_2390,N_572,N_284);
xnor U2391 (N_2391,N_633,N_418);
and U2392 (N_2392,N_88,N_375);
and U2393 (N_2393,N_1245,N_856);
and U2394 (N_2394,N_139,N_1346);
nor U2395 (N_2395,N_729,N_106);
xnor U2396 (N_2396,N_1123,N_87);
xor U2397 (N_2397,N_529,N_471);
nand U2398 (N_2398,N_1395,N_344);
or U2399 (N_2399,N_469,N_1344);
and U2400 (N_2400,N_1373,N_398);
nor U2401 (N_2401,N_865,N_928);
nand U2402 (N_2402,N_361,N_1402);
xor U2403 (N_2403,N_631,N_1307);
or U2404 (N_2404,N_1314,N_1474);
or U2405 (N_2405,N_1435,N_1388);
or U2406 (N_2406,N_708,N_292);
or U2407 (N_2407,N_230,N_1338);
nand U2408 (N_2408,N_1214,N_370);
nand U2409 (N_2409,N_643,N_994);
nand U2410 (N_2410,N_342,N_1276);
nand U2411 (N_2411,N_811,N_20);
nor U2412 (N_2412,N_673,N_851);
nand U2413 (N_2413,N_648,N_1215);
nor U2414 (N_2414,N_146,N_1276);
nand U2415 (N_2415,N_209,N_1487);
xnor U2416 (N_2416,N_1496,N_660);
xnor U2417 (N_2417,N_434,N_974);
and U2418 (N_2418,N_759,N_1415);
nand U2419 (N_2419,N_1083,N_1010);
nor U2420 (N_2420,N_961,N_809);
xor U2421 (N_2421,N_563,N_808);
xnor U2422 (N_2422,N_1039,N_761);
and U2423 (N_2423,N_767,N_191);
or U2424 (N_2424,N_1240,N_654);
xnor U2425 (N_2425,N_421,N_1463);
nor U2426 (N_2426,N_715,N_932);
nand U2427 (N_2427,N_1407,N_1148);
nor U2428 (N_2428,N_52,N_1063);
xor U2429 (N_2429,N_603,N_1112);
xor U2430 (N_2430,N_285,N_509);
nor U2431 (N_2431,N_1278,N_38);
nor U2432 (N_2432,N_507,N_586);
and U2433 (N_2433,N_443,N_245);
and U2434 (N_2434,N_333,N_664);
nor U2435 (N_2435,N_1143,N_931);
and U2436 (N_2436,N_1109,N_958);
and U2437 (N_2437,N_1268,N_823);
nand U2438 (N_2438,N_1204,N_709);
nor U2439 (N_2439,N_401,N_25);
nor U2440 (N_2440,N_253,N_17);
nand U2441 (N_2441,N_223,N_450);
nand U2442 (N_2442,N_1050,N_164);
and U2443 (N_2443,N_1496,N_425);
nand U2444 (N_2444,N_1376,N_1124);
or U2445 (N_2445,N_1066,N_1047);
xor U2446 (N_2446,N_1286,N_1315);
nand U2447 (N_2447,N_591,N_1463);
or U2448 (N_2448,N_1101,N_1374);
nand U2449 (N_2449,N_665,N_498);
xnor U2450 (N_2450,N_1040,N_72);
xnor U2451 (N_2451,N_1269,N_391);
and U2452 (N_2452,N_1061,N_1383);
or U2453 (N_2453,N_828,N_327);
nand U2454 (N_2454,N_287,N_570);
or U2455 (N_2455,N_949,N_408);
and U2456 (N_2456,N_1408,N_809);
nand U2457 (N_2457,N_1035,N_120);
nand U2458 (N_2458,N_1244,N_1098);
and U2459 (N_2459,N_672,N_550);
or U2460 (N_2460,N_479,N_473);
nor U2461 (N_2461,N_155,N_695);
nor U2462 (N_2462,N_1235,N_240);
xnor U2463 (N_2463,N_638,N_194);
or U2464 (N_2464,N_1442,N_36);
or U2465 (N_2465,N_819,N_565);
and U2466 (N_2466,N_754,N_1380);
or U2467 (N_2467,N_954,N_613);
or U2468 (N_2468,N_824,N_1160);
and U2469 (N_2469,N_341,N_1348);
and U2470 (N_2470,N_1443,N_176);
and U2471 (N_2471,N_1297,N_65);
or U2472 (N_2472,N_805,N_844);
and U2473 (N_2473,N_1342,N_557);
or U2474 (N_2474,N_709,N_1015);
xor U2475 (N_2475,N_594,N_885);
nor U2476 (N_2476,N_1455,N_87);
or U2477 (N_2477,N_849,N_232);
xor U2478 (N_2478,N_1485,N_742);
or U2479 (N_2479,N_353,N_1112);
and U2480 (N_2480,N_1484,N_1430);
nand U2481 (N_2481,N_662,N_83);
nand U2482 (N_2482,N_1051,N_1370);
xnor U2483 (N_2483,N_693,N_10);
or U2484 (N_2484,N_460,N_643);
nand U2485 (N_2485,N_1032,N_638);
and U2486 (N_2486,N_1247,N_1330);
nor U2487 (N_2487,N_1168,N_1212);
nand U2488 (N_2488,N_1313,N_472);
nand U2489 (N_2489,N_89,N_1048);
xor U2490 (N_2490,N_519,N_59);
nor U2491 (N_2491,N_43,N_1061);
nor U2492 (N_2492,N_506,N_357);
nand U2493 (N_2493,N_1468,N_620);
or U2494 (N_2494,N_160,N_545);
nor U2495 (N_2495,N_842,N_745);
and U2496 (N_2496,N_146,N_1496);
xor U2497 (N_2497,N_104,N_1352);
nand U2498 (N_2498,N_1151,N_1407);
xor U2499 (N_2499,N_1484,N_109);
nand U2500 (N_2500,N_1343,N_1135);
nor U2501 (N_2501,N_118,N_936);
and U2502 (N_2502,N_588,N_885);
xor U2503 (N_2503,N_1410,N_1458);
and U2504 (N_2504,N_998,N_288);
nand U2505 (N_2505,N_848,N_331);
nor U2506 (N_2506,N_670,N_427);
or U2507 (N_2507,N_1347,N_1260);
xnor U2508 (N_2508,N_965,N_57);
nand U2509 (N_2509,N_12,N_1091);
and U2510 (N_2510,N_637,N_167);
nor U2511 (N_2511,N_1392,N_352);
nand U2512 (N_2512,N_688,N_180);
nor U2513 (N_2513,N_547,N_563);
or U2514 (N_2514,N_1249,N_1371);
and U2515 (N_2515,N_13,N_956);
nand U2516 (N_2516,N_946,N_1003);
nand U2517 (N_2517,N_71,N_396);
or U2518 (N_2518,N_782,N_955);
xor U2519 (N_2519,N_568,N_149);
or U2520 (N_2520,N_780,N_1222);
and U2521 (N_2521,N_187,N_1423);
xor U2522 (N_2522,N_786,N_1126);
and U2523 (N_2523,N_423,N_1169);
xnor U2524 (N_2524,N_738,N_793);
nor U2525 (N_2525,N_647,N_1313);
xor U2526 (N_2526,N_852,N_531);
and U2527 (N_2527,N_1249,N_115);
xnor U2528 (N_2528,N_282,N_771);
xor U2529 (N_2529,N_550,N_838);
xnor U2530 (N_2530,N_897,N_492);
nand U2531 (N_2531,N_1050,N_1048);
and U2532 (N_2532,N_1260,N_672);
and U2533 (N_2533,N_613,N_1473);
and U2534 (N_2534,N_574,N_127);
or U2535 (N_2535,N_747,N_891);
nand U2536 (N_2536,N_1251,N_1284);
nand U2537 (N_2537,N_449,N_1159);
nor U2538 (N_2538,N_580,N_967);
and U2539 (N_2539,N_193,N_657);
nand U2540 (N_2540,N_993,N_1140);
and U2541 (N_2541,N_407,N_878);
or U2542 (N_2542,N_625,N_590);
xnor U2543 (N_2543,N_1443,N_639);
or U2544 (N_2544,N_938,N_840);
xor U2545 (N_2545,N_69,N_398);
nand U2546 (N_2546,N_1032,N_1162);
nand U2547 (N_2547,N_723,N_801);
or U2548 (N_2548,N_1005,N_308);
nor U2549 (N_2549,N_605,N_600);
or U2550 (N_2550,N_130,N_985);
and U2551 (N_2551,N_1053,N_1392);
nor U2552 (N_2552,N_1467,N_462);
and U2553 (N_2553,N_339,N_1024);
nand U2554 (N_2554,N_741,N_1310);
xor U2555 (N_2555,N_450,N_644);
nand U2556 (N_2556,N_1386,N_690);
or U2557 (N_2557,N_1317,N_580);
and U2558 (N_2558,N_983,N_450);
and U2559 (N_2559,N_533,N_1061);
xnor U2560 (N_2560,N_400,N_1349);
and U2561 (N_2561,N_79,N_1316);
and U2562 (N_2562,N_678,N_1286);
xor U2563 (N_2563,N_1412,N_1480);
nor U2564 (N_2564,N_419,N_385);
nand U2565 (N_2565,N_133,N_1139);
xor U2566 (N_2566,N_1041,N_0);
and U2567 (N_2567,N_69,N_751);
nand U2568 (N_2568,N_1162,N_579);
and U2569 (N_2569,N_538,N_1253);
nand U2570 (N_2570,N_987,N_1233);
or U2571 (N_2571,N_371,N_191);
nand U2572 (N_2572,N_59,N_379);
nand U2573 (N_2573,N_440,N_960);
xor U2574 (N_2574,N_201,N_641);
nand U2575 (N_2575,N_196,N_576);
or U2576 (N_2576,N_719,N_1143);
nor U2577 (N_2577,N_1182,N_356);
and U2578 (N_2578,N_854,N_194);
xnor U2579 (N_2579,N_734,N_775);
nor U2580 (N_2580,N_710,N_1396);
or U2581 (N_2581,N_1245,N_443);
nand U2582 (N_2582,N_36,N_100);
nand U2583 (N_2583,N_219,N_661);
nor U2584 (N_2584,N_1473,N_1114);
nor U2585 (N_2585,N_1303,N_35);
xnor U2586 (N_2586,N_1496,N_807);
or U2587 (N_2587,N_988,N_920);
nand U2588 (N_2588,N_364,N_675);
xnor U2589 (N_2589,N_569,N_885);
xnor U2590 (N_2590,N_370,N_281);
nor U2591 (N_2591,N_153,N_460);
nand U2592 (N_2592,N_221,N_390);
or U2593 (N_2593,N_1266,N_977);
or U2594 (N_2594,N_1256,N_417);
xor U2595 (N_2595,N_939,N_138);
nor U2596 (N_2596,N_1086,N_1346);
nor U2597 (N_2597,N_1114,N_741);
nand U2598 (N_2598,N_1429,N_686);
nor U2599 (N_2599,N_634,N_717);
xnor U2600 (N_2600,N_855,N_80);
xnor U2601 (N_2601,N_819,N_990);
xor U2602 (N_2602,N_1452,N_846);
nor U2603 (N_2603,N_846,N_416);
nor U2604 (N_2604,N_295,N_1453);
and U2605 (N_2605,N_322,N_1069);
or U2606 (N_2606,N_1365,N_1429);
xor U2607 (N_2607,N_149,N_479);
nor U2608 (N_2608,N_999,N_919);
or U2609 (N_2609,N_1139,N_424);
and U2610 (N_2610,N_1148,N_826);
xor U2611 (N_2611,N_1178,N_773);
nor U2612 (N_2612,N_615,N_551);
xnor U2613 (N_2613,N_1407,N_1482);
nor U2614 (N_2614,N_92,N_1206);
nand U2615 (N_2615,N_3,N_776);
nand U2616 (N_2616,N_872,N_359);
and U2617 (N_2617,N_239,N_33);
or U2618 (N_2618,N_868,N_1160);
or U2619 (N_2619,N_1194,N_655);
nand U2620 (N_2620,N_451,N_977);
or U2621 (N_2621,N_132,N_1248);
or U2622 (N_2622,N_1264,N_55);
or U2623 (N_2623,N_805,N_1187);
xnor U2624 (N_2624,N_513,N_77);
nor U2625 (N_2625,N_1188,N_864);
nor U2626 (N_2626,N_255,N_1189);
nand U2627 (N_2627,N_140,N_325);
or U2628 (N_2628,N_175,N_632);
and U2629 (N_2629,N_1069,N_695);
or U2630 (N_2630,N_331,N_1443);
and U2631 (N_2631,N_302,N_208);
nor U2632 (N_2632,N_1418,N_237);
xor U2633 (N_2633,N_894,N_279);
nor U2634 (N_2634,N_1428,N_29);
and U2635 (N_2635,N_1151,N_1115);
nor U2636 (N_2636,N_19,N_87);
nor U2637 (N_2637,N_573,N_866);
nor U2638 (N_2638,N_793,N_1204);
and U2639 (N_2639,N_941,N_557);
or U2640 (N_2640,N_612,N_1137);
or U2641 (N_2641,N_169,N_670);
nand U2642 (N_2642,N_1329,N_418);
nand U2643 (N_2643,N_1362,N_21);
and U2644 (N_2644,N_1033,N_1447);
and U2645 (N_2645,N_1429,N_581);
and U2646 (N_2646,N_762,N_592);
nand U2647 (N_2647,N_627,N_575);
nor U2648 (N_2648,N_146,N_1378);
nand U2649 (N_2649,N_1434,N_893);
nor U2650 (N_2650,N_1018,N_858);
or U2651 (N_2651,N_625,N_339);
nand U2652 (N_2652,N_527,N_448);
nand U2653 (N_2653,N_1262,N_329);
or U2654 (N_2654,N_385,N_1232);
nor U2655 (N_2655,N_599,N_1294);
or U2656 (N_2656,N_46,N_1027);
nand U2657 (N_2657,N_1018,N_1068);
and U2658 (N_2658,N_1376,N_188);
and U2659 (N_2659,N_848,N_951);
nor U2660 (N_2660,N_1417,N_597);
nor U2661 (N_2661,N_1382,N_53);
or U2662 (N_2662,N_1067,N_230);
nor U2663 (N_2663,N_530,N_732);
and U2664 (N_2664,N_1265,N_425);
nand U2665 (N_2665,N_1265,N_1259);
nor U2666 (N_2666,N_1020,N_1176);
nand U2667 (N_2667,N_456,N_1006);
xnor U2668 (N_2668,N_1025,N_491);
and U2669 (N_2669,N_663,N_1277);
nand U2670 (N_2670,N_529,N_1296);
nor U2671 (N_2671,N_846,N_1456);
and U2672 (N_2672,N_294,N_811);
and U2673 (N_2673,N_61,N_1451);
nor U2674 (N_2674,N_926,N_1291);
nand U2675 (N_2675,N_1373,N_1138);
nor U2676 (N_2676,N_517,N_921);
nor U2677 (N_2677,N_946,N_1135);
xor U2678 (N_2678,N_1358,N_833);
and U2679 (N_2679,N_237,N_518);
nand U2680 (N_2680,N_538,N_184);
and U2681 (N_2681,N_895,N_343);
xor U2682 (N_2682,N_838,N_468);
xor U2683 (N_2683,N_786,N_358);
nand U2684 (N_2684,N_438,N_847);
nand U2685 (N_2685,N_1158,N_937);
and U2686 (N_2686,N_1188,N_1398);
xor U2687 (N_2687,N_1028,N_42);
nand U2688 (N_2688,N_519,N_669);
or U2689 (N_2689,N_821,N_1026);
nand U2690 (N_2690,N_1168,N_308);
or U2691 (N_2691,N_93,N_42);
and U2692 (N_2692,N_170,N_114);
nor U2693 (N_2693,N_44,N_732);
xor U2694 (N_2694,N_314,N_449);
or U2695 (N_2695,N_846,N_1488);
xnor U2696 (N_2696,N_123,N_608);
xnor U2697 (N_2697,N_1409,N_645);
xnor U2698 (N_2698,N_833,N_309);
or U2699 (N_2699,N_686,N_1469);
and U2700 (N_2700,N_1148,N_585);
or U2701 (N_2701,N_571,N_87);
nor U2702 (N_2702,N_997,N_445);
nor U2703 (N_2703,N_133,N_1091);
nand U2704 (N_2704,N_1311,N_177);
nor U2705 (N_2705,N_924,N_936);
or U2706 (N_2706,N_1199,N_102);
nor U2707 (N_2707,N_1253,N_1201);
nor U2708 (N_2708,N_1225,N_959);
nand U2709 (N_2709,N_613,N_1023);
nand U2710 (N_2710,N_654,N_1402);
nand U2711 (N_2711,N_1068,N_1345);
xnor U2712 (N_2712,N_958,N_301);
xnor U2713 (N_2713,N_214,N_1392);
xnor U2714 (N_2714,N_122,N_1037);
xnor U2715 (N_2715,N_833,N_976);
nor U2716 (N_2716,N_502,N_552);
xnor U2717 (N_2717,N_1313,N_696);
xor U2718 (N_2718,N_381,N_159);
or U2719 (N_2719,N_762,N_939);
and U2720 (N_2720,N_744,N_266);
and U2721 (N_2721,N_623,N_1268);
and U2722 (N_2722,N_1255,N_10);
xor U2723 (N_2723,N_966,N_1044);
xnor U2724 (N_2724,N_400,N_1306);
nand U2725 (N_2725,N_307,N_807);
and U2726 (N_2726,N_592,N_274);
or U2727 (N_2727,N_423,N_762);
xor U2728 (N_2728,N_1369,N_895);
nand U2729 (N_2729,N_434,N_1265);
nand U2730 (N_2730,N_138,N_1179);
and U2731 (N_2731,N_1045,N_1380);
nor U2732 (N_2732,N_316,N_966);
nand U2733 (N_2733,N_192,N_240);
or U2734 (N_2734,N_1249,N_550);
or U2735 (N_2735,N_805,N_905);
nand U2736 (N_2736,N_302,N_544);
and U2737 (N_2737,N_315,N_1415);
and U2738 (N_2738,N_228,N_75);
nand U2739 (N_2739,N_1491,N_1321);
and U2740 (N_2740,N_913,N_440);
nor U2741 (N_2741,N_44,N_1396);
xor U2742 (N_2742,N_1201,N_471);
nor U2743 (N_2743,N_255,N_791);
xor U2744 (N_2744,N_1477,N_92);
or U2745 (N_2745,N_99,N_588);
or U2746 (N_2746,N_1423,N_1139);
xor U2747 (N_2747,N_222,N_1226);
and U2748 (N_2748,N_1325,N_1073);
and U2749 (N_2749,N_171,N_638);
and U2750 (N_2750,N_1289,N_682);
nand U2751 (N_2751,N_509,N_723);
nand U2752 (N_2752,N_1331,N_1273);
nor U2753 (N_2753,N_608,N_1149);
xnor U2754 (N_2754,N_355,N_1012);
nand U2755 (N_2755,N_358,N_1141);
xnor U2756 (N_2756,N_771,N_1210);
or U2757 (N_2757,N_210,N_1137);
nor U2758 (N_2758,N_1056,N_1098);
nand U2759 (N_2759,N_345,N_775);
and U2760 (N_2760,N_1220,N_1164);
nand U2761 (N_2761,N_9,N_1334);
or U2762 (N_2762,N_246,N_406);
or U2763 (N_2763,N_524,N_1327);
or U2764 (N_2764,N_526,N_152);
or U2765 (N_2765,N_951,N_858);
nor U2766 (N_2766,N_69,N_1283);
and U2767 (N_2767,N_184,N_1270);
nor U2768 (N_2768,N_1075,N_1016);
and U2769 (N_2769,N_900,N_1285);
and U2770 (N_2770,N_572,N_1373);
xor U2771 (N_2771,N_502,N_308);
or U2772 (N_2772,N_702,N_527);
xnor U2773 (N_2773,N_1361,N_1345);
nand U2774 (N_2774,N_1220,N_255);
nor U2775 (N_2775,N_1381,N_1189);
or U2776 (N_2776,N_600,N_731);
xor U2777 (N_2777,N_81,N_1468);
nor U2778 (N_2778,N_623,N_1123);
and U2779 (N_2779,N_151,N_859);
xnor U2780 (N_2780,N_887,N_1269);
and U2781 (N_2781,N_553,N_36);
nor U2782 (N_2782,N_347,N_32);
xor U2783 (N_2783,N_1009,N_1303);
nor U2784 (N_2784,N_973,N_1323);
or U2785 (N_2785,N_429,N_1342);
nand U2786 (N_2786,N_660,N_675);
and U2787 (N_2787,N_284,N_929);
and U2788 (N_2788,N_971,N_13);
or U2789 (N_2789,N_740,N_7);
and U2790 (N_2790,N_1286,N_880);
and U2791 (N_2791,N_572,N_841);
nand U2792 (N_2792,N_518,N_680);
and U2793 (N_2793,N_1194,N_1298);
nand U2794 (N_2794,N_1223,N_666);
xor U2795 (N_2795,N_1464,N_645);
xor U2796 (N_2796,N_535,N_34);
or U2797 (N_2797,N_177,N_682);
nor U2798 (N_2798,N_804,N_1166);
xor U2799 (N_2799,N_809,N_998);
or U2800 (N_2800,N_417,N_572);
xor U2801 (N_2801,N_6,N_423);
or U2802 (N_2802,N_73,N_369);
and U2803 (N_2803,N_152,N_484);
nand U2804 (N_2804,N_830,N_265);
and U2805 (N_2805,N_211,N_1122);
nand U2806 (N_2806,N_392,N_630);
and U2807 (N_2807,N_1145,N_1073);
nand U2808 (N_2808,N_423,N_74);
and U2809 (N_2809,N_668,N_966);
xor U2810 (N_2810,N_261,N_1482);
and U2811 (N_2811,N_139,N_1047);
xnor U2812 (N_2812,N_1440,N_446);
nand U2813 (N_2813,N_34,N_1040);
nor U2814 (N_2814,N_695,N_1131);
nand U2815 (N_2815,N_380,N_494);
nand U2816 (N_2816,N_259,N_653);
xor U2817 (N_2817,N_1483,N_441);
or U2818 (N_2818,N_1269,N_1401);
or U2819 (N_2819,N_282,N_879);
xnor U2820 (N_2820,N_304,N_718);
and U2821 (N_2821,N_475,N_988);
and U2822 (N_2822,N_250,N_630);
xnor U2823 (N_2823,N_634,N_417);
xor U2824 (N_2824,N_127,N_1411);
nand U2825 (N_2825,N_178,N_1105);
nor U2826 (N_2826,N_1150,N_1469);
or U2827 (N_2827,N_985,N_162);
nand U2828 (N_2828,N_140,N_575);
and U2829 (N_2829,N_1180,N_628);
and U2830 (N_2830,N_1436,N_58);
nor U2831 (N_2831,N_485,N_380);
and U2832 (N_2832,N_899,N_626);
nand U2833 (N_2833,N_270,N_519);
and U2834 (N_2834,N_185,N_961);
nor U2835 (N_2835,N_746,N_423);
xnor U2836 (N_2836,N_124,N_848);
nand U2837 (N_2837,N_594,N_1085);
nand U2838 (N_2838,N_750,N_401);
xor U2839 (N_2839,N_772,N_375);
xor U2840 (N_2840,N_1346,N_691);
nand U2841 (N_2841,N_485,N_186);
nor U2842 (N_2842,N_801,N_836);
nor U2843 (N_2843,N_1474,N_1204);
and U2844 (N_2844,N_832,N_747);
and U2845 (N_2845,N_654,N_958);
xor U2846 (N_2846,N_651,N_1002);
or U2847 (N_2847,N_136,N_693);
nand U2848 (N_2848,N_1371,N_250);
or U2849 (N_2849,N_444,N_107);
xor U2850 (N_2850,N_1345,N_1447);
nand U2851 (N_2851,N_610,N_1129);
and U2852 (N_2852,N_1200,N_361);
and U2853 (N_2853,N_133,N_75);
xor U2854 (N_2854,N_428,N_986);
nor U2855 (N_2855,N_492,N_1279);
nand U2856 (N_2856,N_247,N_570);
or U2857 (N_2857,N_1450,N_585);
nand U2858 (N_2858,N_1021,N_1335);
nand U2859 (N_2859,N_630,N_923);
nor U2860 (N_2860,N_1016,N_139);
nand U2861 (N_2861,N_1120,N_136);
and U2862 (N_2862,N_1256,N_489);
nand U2863 (N_2863,N_744,N_1440);
xor U2864 (N_2864,N_943,N_576);
and U2865 (N_2865,N_734,N_7);
and U2866 (N_2866,N_13,N_361);
and U2867 (N_2867,N_1113,N_1066);
and U2868 (N_2868,N_481,N_388);
nor U2869 (N_2869,N_1415,N_229);
or U2870 (N_2870,N_173,N_1025);
xnor U2871 (N_2871,N_1150,N_1225);
or U2872 (N_2872,N_1470,N_727);
xor U2873 (N_2873,N_806,N_621);
and U2874 (N_2874,N_47,N_660);
nand U2875 (N_2875,N_1457,N_1431);
nor U2876 (N_2876,N_436,N_847);
nor U2877 (N_2877,N_64,N_143);
and U2878 (N_2878,N_728,N_232);
or U2879 (N_2879,N_1036,N_224);
and U2880 (N_2880,N_655,N_887);
or U2881 (N_2881,N_480,N_885);
nor U2882 (N_2882,N_125,N_553);
or U2883 (N_2883,N_1227,N_1384);
or U2884 (N_2884,N_186,N_1199);
nand U2885 (N_2885,N_1478,N_755);
nand U2886 (N_2886,N_488,N_942);
or U2887 (N_2887,N_315,N_1219);
nand U2888 (N_2888,N_908,N_1316);
and U2889 (N_2889,N_1444,N_1032);
nand U2890 (N_2890,N_1372,N_756);
xnor U2891 (N_2891,N_219,N_493);
and U2892 (N_2892,N_560,N_1308);
nand U2893 (N_2893,N_19,N_965);
and U2894 (N_2894,N_1425,N_1274);
and U2895 (N_2895,N_1425,N_228);
nand U2896 (N_2896,N_1440,N_403);
xnor U2897 (N_2897,N_5,N_98);
nand U2898 (N_2898,N_384,N_899);
xnor U2899 (N_2899,N_1291,N_66);
nand U2900 (N_2900,N_1077,N_310);
and U2901 (N_2901,N_1037,N_607);
nand U2902 (N_2902,N_1101,N_161);
and U2903 (N_2903,N_1495,N_452);
nand U2904 (N_2904,N_799,N_934);
xnor U2905 (N_2905,N_42,N_86);
nor U2906 (N_2906,N_1411,N_287);
nand U2907 (N_2907,N_567,N_390);
xor U2908 (N_2908,N_1168,N_247);
xnor U2909 (N_2909,N_1431,N_1427);
xor U2910 (N_2910,N_79,N_985);
or U2911 (N_2911,N_54,N_1015);
and U2912 (N_2912,N_1473,N_239);
nor U2913 (N_2913,N_1299,N_1260);
or U2914 (N_2914,N_687,N_1035);
nor U2915 (N_2915,N_879,N_128);
xnor U2916 (N_2916,N_70,N_1263);
xor U2917 (N_2917,N_1119,N_1428);
xnor U2918 (N_2918,N_46,N_796);
nand U2919 (N_2919,N_654,N_46);
xor U2920 (N_2920,N_81,N_916);
and U2921 (N_2921,N_254,N_509);
nor U2922 (N_2922,N_907,N_1316);
xor U2923 (N_2923,N_1237,N_1473);
and U2924 (N_2924,N_192,N_203);
nand U2925 (N_2925,N_612,N_207);
nor U2926 (N_2926,N_526,N_188);
or U2927 (N_2927,N_1252,N_421);
xnor U2928 (N_2928,N_167,N_206);
or U2929 (N_2929,N_87,N_534);
nand U2930 (N_2930,N_873,N_217);
xnor U2931 (N_2931,N_849,N_1094);
nor U2932 (N_2932,N_113,N_325);
and U2933 (N_2933,N_901,N_503);
and U2934 (N_2934,N_346,N_886);
nor U2935 (N_2935,N_357,N_727);
xor U2936 (N_2936,N_50,N_499);
nand U2937 (N_2937,N_66,N_332);
xor U2938 (N_2938,N_660,N_1114);
nand U2939 (N_2939,N_1490,N_410);
or U2940 (N_2940,N_1191,N_365);
and U2941 (N_2941,N_1023,N_1008);
xor U2942 (N_2942,N_1160,N_131);
and U2943 (N_2943,N_789,N_355);
and U2944 (N_2944,N_912,N_1097);
nor U2945 (N_2945,N_36,N_385);
or U2946 (N_2946,N_1177,N_863);
or U2947 (N_2947,N_120,N_1088);
xnor U2948 (N_2948,N_1446,N_852);
or U2949 (N_2949,N_1205,N_273);
xor U2950 (N_2950,N_276,N_363);
and U2951 (N_2951,N_117,N_858);
nor U2952 (N_2952,N_1282,N_1163);
xnor U2953 (N_2953,N_1431,N_1179);
and U2954 (N_2954,N_963,N_1031);
xor U2955 (N_2955,N_356,N_1439);
xnor U2956 (N_2956,N_895,N_122);
xor U2957 (N_2957,N_66,N_555);
nor U2958 (N_2958,N_1436,N_824);
nand U2959 (N_2959,N_1073,N_1354);
or U2960 (N_2960,N_814,N_1125);
and U2961 (N_2961,N_489,N_680);
xnor U2962 (N_2962,N_940,N_1340);
xnor U2963 (N_2963,N_830,N_393);
or U2964 (N_2964,N_522,N_1303);
and U2965 (N_2965,N_802,N_49);
nand U2966 (N_2966,N_1376,N_279);
or U2967 (N_2967,N_1118,N_628);
and U2968 (N_2968,N_1387,N_86);
xor U2969 (N_2969,N_224,N_577);
nor U2970 (N_2970,N_1357,N_1088);
nor U2971 (N_2971,N_873,N_636);
xor U2972 (N_2972,N_166,N_177);
and U2973 (N_2973,N_919,N_292);
nand U2974 (N_2974,N_262,N_1384);
or U2975 (N_2975,N_1231,N_1470);
nor U2976 (N_2976,N_1499,N_659);
or U2977 (N_2977,N_1025,N_1484);
nor U2978 (N_2978,N_849,N_1437);
nand U2979 (N_2979,N_1405,N_481);
and U2980 (N_2980,N_91,N_1206);
and U2981 (N_2981,N_1274,N_491);
xnor U2982 (N_2982,N_1470,N_1121);
and U2983 (N_2983,N_1362,N_909);
and U2984 (N_2984,N_398,N_400);
nor U2985 (N_2985,N_218,N_1149);
nand U2986 (N_2986,N_853,N_1218);
nor U2987 (N_2987,N_1045,N_1145);
nand U2988 (N_2988,N_1353,N_55);
or U2989 (N_2989,N_700,N_913);
nand U2990 (N_2990,N_1154,N_677);
xor U2991 (N_2991,N_818,N_1406);
xnor U2992 (N_2992,N_625,N_1012);
or U2993 (N_2993,N_611,N_449);
xnor U2994 (N_2994,N_337,N_817);
or U2995 (N_2995,N_817,N_1019);
or U2996 (N_2996,N_373,N_1144);
nand U2997 (N_2997,N_78,N_1425);
nor U2998 (N_2998,N_1152,N_47);
and U2999 (N_2999,N_1324,N_341);
and U3000 (N_3000,N_1616,N_2782);
and U3001 (N_3001,N_2112,N_2804);
nand U3002 (N_3002,N_1786,N_2096);
or U3003 (N_3003,N_2010,N_2329);
xnor U3004 (N_3004,N_2526,N_2139);
nor U3005 (N_3005,N_2473,N_1799);
nand U3006 (N_3006,N_1985,N_1706);
xor U3007 (N_3007,N_2753,N_1612);
xor U3008 (N_3008,N_2118,N_2882);
nand U3009 (N_3009,N_2244,N_2859);
and U3010 (N_3010,N_2805,N_2016);
and U3011 (N_3011,N_2463,N_2959);
nand U3012 (N_3012,N_1641,N_2320);
nor U3013 (N_3013,N_1816,N_2190);
or U3014 (N_3014,N_1746,N_2057);
nor U3015 (N_3015,N_1865,N_2348);
xnor U3016 (N_3016,N_2440,N_2145);
xnor U3017 (N_3017,N_1782,N_1956);
or U3018 (N_3018,N_2628,N_1548);
nor U3019 (N_3019,N_1827,N_1769);
nor U3020 (N_3020,N_2484,N_1747);
or U3021 (N_3021,N_2087,N_1589);
xor U3022 (N_3022,N_2012,N_2925);
xor U3023 (N_3023,N_2779,N_2806);
nand U3024 (N_3024,N_2441,N_1748);
nor U3025 (N_3025,N_1707,N_2266);
and U3026 (N_3026,N_1951,N_1656);
and U3027 (N_3027,N_1536,N_2319);
xnor U3028 (N_3028,N_1726,N_2129);
nor U3029 (N_3029,N_2454,N_2234);
or U3030 (N_3030,N_2910,N_2227);
nand U3031 (N_3031,N_2342,N_2403);
or U3032 (N_3032,N_2969,N_2801);
nor U3033 (N_3033,N_2477,N_2379);
nand U3034 (N_3034,N_2604,N_2461);
xor U3035 (N_3035,N_2887,N_2412);
xor U3036 (N_3036,N_1744,N_2174);
or U3037 (N_3037,N_1849,N_2014);
nor U3038 (N_3038,N_1884,N_2549);
or U3039 (N_3039,N_1636,N_2920);
nor U3040 (N_3040,N_2027,N_2019);
nor U3041 (N_3041,N_1540,N_2563);
and U3042 (N_3042,N_1648,N_1962);
nand U3043 (N_3043,N_1992,N_1917);
nand U3044 (N_3044,N_2817,N_1960);
nor U3045 (N_3045,N_2942,N_2172);
or U3046 (N_3046,N_2094,N_2072);
xor U3047 (N_3047,N_1520,N_1991);
and U3048 (N_3048,N_1561,N_2991);
and U3049 (N_3049,N_1879,N_2229);
and U3050 (N_3050,N_2772,N_2207);
nand U3051 (N_3051,N_2562,N_2356);
nor U3052 (N_3052,N_2392,N_1547);
xor U3053 (N_3053,N_1607,N_2505);
nand U3054 (N_3054,N_2049,N_2247);
or U3055 (N_3055,N_1683,N_2273);
nand U3056 (N_3056,N_2109,N_2789);
and U3057 (N_3057,N_1899,N_2545);
or U3058 (N_3058,N_1688,N_2040);
and U3059 (N_3059,N_2557,N_1659);
or U3060 (N_3060,N_2099,N_1657);
or U3061 (N_3061,N_1929,N_2203);
nand U3062 (N_3062,N_2961,N_2922);
and U3063 (N_3063,N_2659,N_1949);
nor U3064 (N_3064,N_1701,N_2693);
or U3065 (N_3065,N_2586,N_1768);
xor U3066 (N_3066,N_2200,N_2485);
xnor U3067 (N_3067,N_2107,N_1613);
or U3068 (N_3068,N_2464,N_2359);
or U3069 (N_3069,N_1761,N_1762);
nor U3070 (N_3070,N_2222,N_1982);
and U3071 (N_3071,N_2582,N_2799);
xnor U3072 (N_3072,N_1663,N_1564);
nor U3073 (N_3073,N_1878,N_1546);
or U3074 (N_3074,N_2666,N_1605);
nor U3075 (N_3075,N_2315,N_1753);
xnor U3076 (N_3076,N_1594,N_2541);
nand U3077 (N_3077,N_1802,N_1886);
nand U3078 (N_3078,N_2085,N_2343);
xor U3079 (N_3079,N_2818,N_2990);
or U3080 (N_3080,N_2766,N_2381);
or U3081 (N_3081,N_2089,N_2154);
nand U3082 (N_3082,N_2603,N_2930);
xnor U3083 (N_3083,N_2377,N_1711);
nand U3084 (N_3084,N_2785,N_1887);
nand U3085 (N_3085,N_2728,N_1972);
and U3086 (N_3086,N_2559,N_1759);
nand U3087 (N_3087,N_2147,N_1506);
and U3088 (N_3088,N_2214,N_1981);
and U3089 (N_3089,N_2476,N_2896);
nor U3090 (N_3090,N_1731,N_2593);
xnor U3091 (N_3091,N_2974,N_2909);
and U3092 (N_3092,N_1674,N_2196);
nor U3093 (N_3093,N_2899,N_2550);
xor U3094 (N_3094,N_2372,N_2796);
nand U3095 (N_3095,N_2385,N_2626);
nor U3096 (N_3096,N_2439,N_1596);
nor U3097 (N_3097,N_2965,N_1534);
nand U3098 (N_3098,N_2544,N_2836);
nor U3099 (N_3099,N_1932,N_2369);
xnor U3100 (N_3100,N_1653,N_2687);
and U3101 (N_3101,N_2396,N_1790);
nor U3102 (N_3102,N_2904,N_1999);
nand U3103 (N_3103,N_2043,N_2050);
nand U3104 (N_3104,N_2652,N_2455);
nand U3105 (N_3105,N_2890,N_1647);
and U3106 (N_3106,N_2187,N_2707);
nor U3107 (N_3107,N_2558,N_2434);
nand U3108 (N_3108,N_2255,N_2475);
nor U3109 (N_3109,N_1687,N_2765);
nand U3110 (N_3110,N_2722,N_2824);
and U3111 (N_3111,N_2345,N_2560);
or U3112 (N_3112,N_2325,N_2422);
and U3113 (N_3113,N_2729,N_1888);
nand U3114 (N_3114,N_1758,N_2474);
and U3115 (N_3115,N_1832,N_1538);
xor U3116 (N_3116,N_1697,N_1939);
nand U3117 (N_3117,N_1915,N_2192);
or U3118 (N_3118,N_2781,N_2250);
and U3119 (N_3119,N_2000,N_1974);
nand U3120 (N_3120,N_2874,N_1576);
and U3121 (N_3121,N_2240,N_1639);
nor U3122 (N_3122,N_1608,N_1535);
nor U3123 (N_3123,N_2860,N_2996);
nor U3124 (N_3124,N_2185,N_1692);
xnor U3125 (N_3125,N_1842,N_1825);
and U3126 (N_3126,N_2274,N_2408);
nor U3127 (N_3127,N_2931,N_2241);
xnor U3128 (N_3128,N_1791,N_1959);
or U3129 (N_3129,N_1710,N_2142);
xor U3130 (N_3130,N_2522,N_1785);
or U3131 (N_3131,N_2703,N_1812);
and U3132 (N_3132,N_2637,N_2960);
nand U3133 (N_3133,N_2872,N_2847);
nor U3134 (N_3134,N_2238,N_2326);
and U3135 (N_3135,N_2862,N_2378);
nand U3136 (N_3136,N_1515,N_2675);
nor U3137 (N_3137,N_2483,N_2606);
or U3138 (N_3138,N_1723,N_2263);
nand U3139 (N_3139,N_2973,N_2022);
xor U3140 (N_3140,N_1914,N_1783);
nand U3141 (N_3141,N_2173,N_2365);
nand U3142 (N_3142,N_2084,N_1655);
nand U3143 (N_3143,N_1779,N_2747);
and U3144 (N_3144,N_2748,N_1580);
and U3145 (N_3145,N_1621,N_2540);
xor U3146 (N_3146,N_2720,N_1798);
nand U3147 (N_3147,N_2144,N_2656);
or U3148 (N_3148,N_2865,N_1752);
and U3149 (N_3149,N_2776,N_2391);
xor U3150 (N_3150,N_2199,N_1642);
nor U3151 (N_3151,N_2008,N_1863);
or U3152 (N_3152,N_2823,N_2808);
nand U3153 (N_3153,N_2283,N_1821);
nor U3154 (N_3154,N_2984,N_2225);
and U3155 (N_3155,N_2394,N_2625);
xnor U3156 (N_3156,N_2082,N_2884);
or U3157 (N_3157,N_2067,N_2528);
nand U3158 (N_3158,N_2682,N_2253);
or U3159 (N_3159,N_2344,N_1504);
and U3160 (N_3160,N_2695,N_2148);
and U3161 (N_3161,N_2055,N_1780);
nor U3162 (N_3162,N_2955,N_1893);
nand U3163 (N_3163,N_1591,N_1989);
and U3164 (N_3164,N_2193,N_1619);
nor U3165 (N_3165,N_1807,N_2061);
xnor U3166 (N_3166,N_2009,N_2617);
xnor U3167 (N_3167,N_1852,N_2797);
xor U3168 (N_3168,N_1528,N_2376);
xor U3169 (N_3169,N_2191,N_2683);
nand U3170 (N_3170,N_2355,N_1850);
nor U3171 (N_3171,N_2104,N_2023);
nand U3172 (N_3172,N_2878,N_2332);
xor U3173 (N_3173,N_1705,N_2533);
nor U3174 (N_3174,N_2845,N_1671);
nor U3175 (N_3175,N_2709,N_1599);
nand U3176 (N_3176,N_2135,N_2171);
nor U3177 (N_3177,N_2945,N_2843);
or U3178 (N_3178,N_1637,N_2065);
nand U3179 (N_3179,N_2764,N_2224);
xor U3180 (N_3180,N_1730,N_2598);
or U3181 (N_3181,N_2654,N_2091);
nand U3182 (N_3182,N_1900,N_2001);
or U3183 (N_3183,N_2892,N_1675);
or U3184 (N_3184,N_1595,N_2948);
or U3185 (N_3185,N_2246,N_2552);
xor U3186 (N_3186,N_2197,N_2432);
nor U3187 (N_3187,N_1664,N_2727);
xnor U3188 (N_3188,N_2641,N_2854);
and U3189 (N_3189,N_1524,N_2844);
nand U3190 (N_3190,N_2730,N_2803);
nor U3191 (N_3191,N_2795,N_2750);
and U3192 (N_3192,N_2731,N_2116);
xor U3193 (N_3193,N_1623,N_2302);
xnor U3194 (N_3194,N_2208,N_2855);
or U3195 (N_3195,N_2100,N_2151);
xnor U3196 (N_3196,N_2223,N_2968);
xnor U3197 (N_3197,N_2964,N_1829);
nor U3198 (N_3198,N_2269,N_1502);
nand U3199 (N_3199,N_2608,N_2346);
or U3200 (N_3200,N_1615,N_2630);
nand U3201 (N_3201,N_1880,N_2062);
xor U3202 (N_3202,N_1976,N_2600);
and U3203 (N_3203,N_2431,N_1885);
and U3204 (N_3204,N_1874,N_1630);
xnor U3205 (N_3205,N_1715,N_2259);
or U3206 (N_3206,N_2835,N_2128);
nor U3207 (N_3207,N_2627,N_2577);
xnor U3208 (N_3208,N_2068,N_2827);
nor U3209 (N_3209,N_2839,N_2537);
xnor U3210 (N_3210,N_2678,N_2640);
nor U3211 (N_3211,N_1679,N_2815);
nand U3212 (N_3212,N_1570,N_2936);
or U3213 (N_3213,N_2251,N_2987);
and U3214 (N_3214,N_2140,N_2021);
or U3215 (N_3215,N_2445,N_2900);
nand U3216 (N_3216,N_2364,N_2609);
and U3217 (N_3217,N_2066,N_1892);
or U3218 (N_3218,N_2168,N_2673);
and U3219 (N_3219,N_2424,N_2689);
or U3220 (N_3220,N_1864,N_2712);
or U3221 (N_3221,N_1559,N_2778);
nand U3222 (N_3222,N_1704,N_2902);
nor U3223 (N_3223,N_2306,N_2571);
nand U3224 (N_3224,N_1517,N_2733);
nand U3225 (N_3225,N_1530,N_2405);
and U3226 (N_3226,N_2481,N_2363);
nor U3227 (N_3227,N_2327,N_1624);
nand U3228 (N_3228,N_2773,N_1733);
and U3229 (N_3229,N_1658,N_2696);
nor U3230 (N_3230,N_1954,N_2447);
nor U3231 (N_3231,N_2536,N_2256);
and U3232 (N_3232,N_2397,N_1646);
nor U3233 (N_3233,N_1720,N_1582);
nand U3234 (N_3234,N_2108,N_2032);
or U3235 (N_3235,N_2525,N_2449);
nor U3236 (N_3236,N_2740,N_2003);
or U3237 (N_3237,N_2460,N_1618);
and U3238 (N_3238,N_1795,N_2267);
and U3239 (N_3239,N_2122,N_2233);
nand U3240 (N_3240,N_1562,N_2771);
or U3241 (N_3241,N_2458,N_1940);
nor U3242 (N_3242,N_2162,N_2569);
xnor U3243 (N_3243,N_2794,N_2564);
and U3244 (N_3244,N_1877,N_1708);
or U3245 (N_3245,N_1567,N_2573);
or U3246 (N_3246,N_2868,N_1862);
xnor U3247 (N_3247,N_2383,N_1859);
xor U3248 (N_3248,N_2894,N_2056);
nor U3249 (N_3249,N_2702,N_2430);
and U3250 (N_3250,N_2311,N_2366);
nand U3251 (N_3251,N_2442,N_2111);
xnor U3252 (N_3252,N_1776,N_2098);
and U3253 (N_3253,N_2195,N_2752);
and U3254 (N_3254,N_2788,N_2787);
xor U3255 (N_3255,N_2914,N_2141);
and U3256 (N_3256,N_1691,N_1539);
nand U3257 (N_3257,N_1818,N_2851);
and U3258 (N_3258,N_1550,N_2530);
nor U3259 (N_3259,N_2982,N_2534);
nor U3260 (N_3260,N_1926,N_2388);
xor U3261 (N_3261,N_2301,N_2287);
nor U3262 (N_3262,N_1660,N_1868);
nand U3263 (N_3263,N_2706,N_1871);
nand U3264 (N_3264,N_2024,N_2998);
or U3265 (N_3265,N_1728,N_2456);
and U3266 (N_3266,N_2239,N_2264);
xnor U3267 (N_3267,N_2946,N_1967);
or U3268 (N_3268,N_2840,N_2158);
and U3269 (N_3269,N_2038,N_2331);
xnor U3270 (N_3270,N_2286,N_2482);
or U3271 (N_3271,N_1794,N_2828);
and U3272 (N_3272,N_2755,N_2680);
or U3273 (N_3273,N_1512,N_2163);
nor U3274 (N_3274,N_2888,N_1627);
or U3275 (N_3275,N_2291,N_1916);
or U3276 (N_3276,N_1853,N_1604);
or U3277 (N_3277,N_1973,N_1765);
xor U3278 (N_3278,N_2967,N_1668);
or U3279 (N_3279,N_2511,N_2030);
xnor U3280 (N_3280,N_1793,N_2212);
or U3281 (N_3281,N_2188,N_2210);
or U3282 (N_3282,N_2206,N_2318);
xor U3283 (N_3283,N_2143,N_1797);
xnor U3284 (N_3284,N_2113,N_1650);
and U3285 (N_3285,N_2837,N_1652);
nand U3286 (N_3286,N_2903,N_2940);
and U3287 (N_3287,N_2471,N_1993);
nor U3288 (N_3288,N_1609,N_2048);
nand U3289 (N_3289,N_2334,N_2452);
xor U3290 (N_3290,N_2323,N_1775);
nand U3291 (N_3291,N_2181,N_1597);
nand U3292 (N_3292,N_2417,N_2723);
nand U3293 (N_3293,N_2531,N_1680);
or U3294 (N_3294,N_2711,N_2047);
or U3295 (N_3295,N_2226,N_2036);
nor U3296 (N_3296,N_2347,N_2297);
nor U3297 (N_3297,N_2947,N_1695);
nor U3298 (N_3298,N_2176,N_2130);
nand U3299 (N_3299,N_2125,N_1840);
nand U3300 (N_3300,N_1774,N_1861);
nor U3301 (N_3301,N_2700,N_2653);
xor U3302 (N_3302,N_1667,N_2951);
and U3303 (N_3303,N_2595,N_2086);
and U3304 (N_3304,N_1883,N_2761);
and U3305 (N_3305,N_2262,N_1971);
xor U3306 (N_3306,N_2167,N_1945);
xnor U3307 (N_3307,N_2136,N_2127);
nand U3308 (N_3308,N_2491,N_2891);
nand U3309 (N_3309,N_2917,N_1645);
or U3310 (N_3310,N_2419,N_1507);
or U3311 (N_3311,N_2395,N_2415);
nand U3312 (N_3312,N_1537,N_2303);
nor U3313 (N_3313,N_2514,N_2426);
nand U3314 (N_3314,N_2261,N_2005);
and U3315 (N_3315,N_1523,N_1770);
xnor U3316 (N_3316,N_1923,N_2290);
or U3317 (N_3317,N_1633,N_1568);
nor U3318 (N_3318,N_1727,N_2590);
or U3319 (N_3319,N_2852,N_2978);
nand U3320 (N_3320,N_2769,N_2293);
and U3321 (N_3321,N_2390,N_1846);
nor U3322 (N_3322,N_2179,N_2893);
nand U3323 (N_3323,N_2927,N_2393);
nand U3324 (N_3324,N_2970,N_1970);
nor U3325 (N_3325,N_2619,N_2184);
or U3326 (N_3326,N_1845,N_1709);
nor U3327 (N_3327,N_2800,N_2101);
nor U3328 (N_3328,N_1577,N_1751);
or U3329 (N_3329,N_2863,N_1778);
nand U3330 (N_3330,N_2280,N_2639);
nand U3331 (N_3331,N_2074,N_1684);
and U3332 (N_3332,N_2643,N_1978);
xnor U3333 (N_3333,N_2983,N_1673);
or U3334 (N_3334,N_2416,N_2219);
and U3335 (N_3335,N_2919,N_2295);
nand U3336 (N_3336,N_2749,N_2042);
nor U3337 (N_3337,N_1743,N_2739);
xor U3338 (N_3338,N_2592,N_1532);
nor U3339 (N_3339,N_2596,N_1928);
and U3340 (N_3340,N_1854,N_2398);
or U3341 (N_3341,N_2153,N_2258);
and U3342 (N_3342,N_2816,N_2493);
nand U3343 (N_3343,N_2202,N_2017);
xnor U3344 (N_3344,N_1844,N_1957);
or U3345 (N_3345,N_2849,N_1558);
and U3346 (N_3346,N_2133,N_2532);
and U3347 (N_3347,N_2612,N_2883);
or U3348 (N_3348,N_2205,N_2809);
or U3349 (N_3349,N_2581,N_2567);
or U3350 (N_3350,N_2825,N_1702);
nor U3351 (N_3351,N_1651,N_2490);
xnor U3352 (N_3352,N_2307,N_2985);
or U3353 (N_3353,N_2324,N_1964);
nand U3354 (N_3354,N_1766,N_2513);
or U3355 (N_3355,N_2620,N_1937);
and U3356 (N_3356,N_1822,N_2438);
nor U3357 (N_3357,N_2611,N_2102);
and U3358 (N_3358,N_2811,N_2830);
or U3359 (N_3359,N_2688,N_1529);
and U3360 (N_3360,N_2516,N_2367);
and U3361 (N_3361,N_2076,N_1969);
xnor U3362 (N_3362,N_2570,N_2783);
xor U3363 (N_3363,N_2155,N_1904);
or U3364 (N_3364,N_2252,N_1631);
and U3365 (N_3365,N_1541,N_1511);
nor U3366 (N_3366,N_1551,N_2648);
and U3367 (N_3367,N_2160,N_1866);
and U3368 (N_3368,N_1736,N_2907);
nor U3369 (N_3369,N_2236,N_1872);
xnor U3370 (N_3370,N_1942,N_2124);
or U3371 (N_3371,N_1737,N_2999);
nor U3372 (N_3372,N_2615,N_2183);
nand U3373 (N_3373,N_1533,N_2131);
xor U3374 (N_3374,N_2686,N_1741);
or U3375 (N_3375,N_2953,N_1677);
nand U3376 (N_3376,N_1620,N_2770);
or U3377 (N_3377,N_2336,N_1689);
nand U3378 (N_3378,N_2235,N_2231);
nand U3379 (N_3379,N_1514,N_2864);
xnor U3380 (N_3380,N_2069,N_2576);
nand U3381 (N_3381,N_2508,N_2822);
or U3382 (N_3382,N_1943,N_2446);
xor U3383 (N_3383,N_1920,N_2885);
nor U3384 (N_3384,N_2157,N_2833);
or U3385 (N_3385,N_2480,N_2333);
or U3386 (N_3386,N_2995,N_2052);
or U3387 (N_3387,N_2046,N_1738);
xnor U3388 (N_3388,N_1955,N_2501);
xnor U3389 (N_3389,N_2725,N_1950);
xnor U3390 (N_3390,N_2362,N_2025);
xnor U3391 (N_3391,N_1724,N_1958);
and U3392 (N_3392,N_2813,N_2243);
xnor U3393 (N_3393,N_2414,N_2044);
nor U3394 (N_3394,N_2121,N_2360);
nor U3395 (N_3395,N_2605,N_1681);
xnor U3396 (N_3396,N_2309,N_1760);
nand U3397 (N_3397,N_2340,N_1921);
xnor U3398 (N_3398,N_2736,N_2510);
or U3399 (N_3399,N_1555,N_1781);
nand U3400 (N_3400,N_2775,N_2499);
or U3401 (N_3401,N_1544,N_2175);
or U3402 (N_3402,N_2992,N_1686);
and U3403 (N_3403,N_2715,N_1834);
xor U3404 (N_3404,N_1699,N_2591);
nor U3405 (N_3405,N_2034,N_2095);
and U3406 (N_3406,N_2507,N_2186);
and U3407 (N_3407,N_2786,N_1771);
nand U3408 (N_3408,N_2589,N_1573);
and U3409 (N_3409,N_1767,N_1755);
or U3410 (N_3410,N_2539,N_1732);
xor U3411 (N_3411,N_1830,N_2404);
or U3412 (N_3412,N_2583,N_2245);
nor U3413 (N_3413,N_2691,N_2088);
nor U3414 (N_3414,N_2138,N_2704);
or U3415 (N_3415,N_2632,N_2956);
nand U3416 (N_3416,N_2759,N_1610);
nor U3417 (N_3417,N_1581,N_2103);
xor U3418 (N_3418,N_2838,N_2807);
nor U3419 (N_3419,N_2368,N_1997);
xnor U3420 (N_3420,N_2667,N_1526);
and U3421 (N_3421,N_1678,N_2895);
or U3422 (N_3422,N_1763,N_1784);
xnor U3423 (N_3423,N_1870,N_1856);
nor U3424 (N_3424,N_2486,N_2300);
nor U3425 (N_3425,N_2784,N_2421);
and U3426 (N_3426,N_2658,N_2875);
or U3427 (N_3427,N_1841,N_2672);
nor U3428 (N_3428,N_2018,N_2923);
or U3429 (N_3429,N_2879,N_2081);
and U3430 (N_3430,N_1585,N_2798);
nor U3431 (N_3431,N_1666,N_2543);
nor U3432 (N_3432,N_2646,N_2926);
nor U3433 (N_3433,N_2793,N_2436);
nand U3434 (N_3434,N_2270,N_2738);
and U3435 (N_3435,N_2670,N_2734);
and U3436 (N_3436,N_1953,N_2977);
nor U3437 (N_3437,N_2380,N_2556);
nand U3438 (N_3438,N_2232,N_2073);
xor U3439 (N_3439,N_2314,N_1662);
nand U3440 (N_3440,N_2399,N_2650);
or U3441 (N_3441,N_1948,N_2834);
or U3442 (N_3442,N_2468,N_1556);
xor U3443 (N_3443,N_2459,N_2848);
nand U3444 (N_3444,N_1661,N_2497);
and U3445 (N_3445,N_1603,N_1819);
or U3446 (N_3446,N_2466,N_1922);
and U3447 (N_3447,N_2039,N_1516);
and U3448 (N_3448,N_2819,N_1882);
and U3449 (N_3449,N_2580,N_1936);
and U3450 (N_3450,N_2880,N_1890);
or U3451 (N_3451,N_1907,N_2370);
nor U3452 (N_3452,N_2305,N_2120);
xnor U3453 (N_3453,N_2520,N_2349);
xnor U3454 (N_3454,N_1503,N_2915);
and U3455 (N_3455,N_2745,N_2943);
and U3456 (N_3456,N_1895,N_2515);
and U3457 (N_3457,N_2821,N_2685);
or U3458 (N_3458,N_2897,N_2437);
and U3459 (N_3459,N_2189,N_1806);
nor U3460 (N_3460,N_2870,N_1961);
nand U3461 (N_3461,N_2401,N_2448);
and U3462 (N_3462,N_2294,N_1898);
and U3463 (N_3463,N_2754,N_2029);
xnor U3464 (N_3464,N_2166,N_1975);
xnor U3465 (N_3465,N_2002,N_2092);
and U3466 (N_3466,N_1754,N_2519);
nor U3467 (N_3467,N_2535,N_2861);
xnor U3468 (N_3468,N_2792,N_2150);
or U3469 (N_3469,N_2007,N_2677);
xnor U3470 (N_3470,N_1810,N_1788);
and U3471 (N_3471,N_2699,N_1734);
xnor U3472 (N_3472,N_2435,N_2413);
and U3473 (N_3473,N_2972,N_2574);
or U3474 (N_3474,N_2070,N_2976);
and U3475 (N_3475,N_2674,N_1601);
xor U3476 (N_3476,N_2271,N_2777);
or U3477 (N_3477,N_1833,N_1977);
or U3478 (N_3478,N_2209,N_2607);
nand U3479 (N_3479,N_1946,N_2767);
or U3480 (N_3480,N_2676,N_2724);
and U3481 (N_3481,N_2737,N_2820);
and U3482 (N_3482,N_2791,N_1569);
nor U3483 (N_3483,N_2033,N_2935);
xor U3484 (N_3484,N_1944,N_2279);
nor U3485 (N_3485,N_1625,N_2020);
nor U3486 (N_3486,N_2518,N_2117);
or U3487 (N_3487,N_2554,N_2579);
nor U3488 (N_3488,N_2928,N_2975);
nand U3489 (N_3489,N_2994,N_1897);
xor U3490 (N_3490,N_1518,N_1682);
or U3491 (N_3491,N_2751,N_2906);
or U3492 (N_3492,N_1965,N_2644);
nand U3493 (N_3493,N_1789,N_1593);
nand U3494 (N_3494,N_2826,N_1716);
nor U3495 (N_3495,N_1531,N_2054);
and U3496 (N_3496,N_2555,N_2097);
and U3497 (N_3497,N_2106,N_2420);
nand U3498 (N_3498,N_2374,N_2812);
xnor U3499 (N_3499,N_2078,N_2871);
or U3500 (N_3500,N_2886,N_1519);
and U3501 (N_3501,N_1773,N_1501);
and U3502 (N_3502,N_2502,N_2763);
xnor U3503 (N_3503,N_2450,N_2265);
and U3504 (N_3504,N_1930,N_1764);
or U3505 (N_3505,N_2159,N_1719);
and U3506 (N_3506,N_2743,N_1934);
nor U3507 (N_3507,N_2407,N_1891);
or U3508 (N_3508,N_2866,N_2433);
and U3509 (N_3509,N_1574,N_1557);
or U3510 (N_3510,N_1903,N_2944);
and U3511 (N_3511,N_2004,N_2857);
and U3512 (N_3512,N_2277,N_1722);
or U3513 (N_3513,N_2498,N_2064);
or U3514 (N_3514,N_2913,N_2829);
or U3515 (N_3515,N_2134,N_2911);
nor U3516 (N_3516,N_1740,N_2624);
nor U3517 (N_3517,N_1598,N_1602);
or U3518 (N_3518,N_2547,N_1800);
nand U3519 (N_3519,N_2832,N_2802);
xnor U3520 (N_3520,N_2993,N_2308);
nor U3521 (N_3521,N_2217,N_2671);
and U3522 (N_3522,N_1805,N_2929);
nand U3523 (N_3523,N_2523,N_1521);
nand U3524 (N_3524,N_2952,N_2105);
or U3525 (N_3525,N_1925,N_1698);
and U3526 (N_3526,N_2714,N_1729);
or U3527 (N_3527,N_2869,N_2979);
xor U3528 (N_3528,N_2713,N_1966);
nand U3529 (N_3529,N_1909,N_2846);
or U3530 (N_3530,N_2079,N_1912);
nand U3531 (N_3531,N_1685,N_2694);
nand U3532 (N_3532,N_1858,N_2338);
xor U3533 (N_3533,N_1565,N_2981);
and U3534 (N_3534,N_2119,N_2220);
xor U3535 (N_3535,N_1838,N_2517);
xnor U3536 (N_3536,N_1839,N_2758);
xor U3537 (N_3537,N_2410,N_1665);
or U3538 (N_3538,N_1614,N_2180);
and U3539 (N_3539,N_1809,N_2889);
xor U3540 (N_3540,N_1979,N_1983);
xor U3541 (N_3541,N_1587,N_1542);
and U3542 (N_3542,N_1980,N_2623);
xor U3543 (N_3543,N_2500,N_2177);
or U3544 (N_3544,N_2651,N_1906);
nand U3545 (N_3545,N_2469,N_2351);
nor U3546 (N_3546,N_2877,N_2661);
xnor U3547 (N_3547,N_2488,N_2585);
nor U3548 (N_3548,N_2288,N_1996);
xnor U3549 (N_3549,N_2170,N_2506);
xnor U3550 (N_3550,N_1693,N_2698);
nor U3551 (N_3551,N_2566,N_1813);
nor U3552 (N_3552,N_1938,N_2735);
and U3553 (N_3553,N_1919,N_1575);
nor U3554 (N_3554,N_1995,N_2282);
or U3555 (N_3555,N_2411,N_1984);
or U3556 (N_3556,N_2873,N_2921);
nor U3557 (N_3557,N_2527,N_2165);
and U3558 (N_3558,N_2645,N_2588);
nor U3559 (N_3559,N_1994,N_2853);
xor U3560 (N_3560,N_2912,N_2281);
xor U3561 (N_3561,N_1756,N_2152);
or U3562 (N_3562,N_1632,N_2132);
or U3563 (N_3563,N_1654,N_2053);
and U3564 (N_3564,N_1824,N_1509);
and U3565 (N_3565,N_2215,N_1745);
nor U3566 (N_3566,N_2313,N_2575);
nand U3567 (N_3567,N_2831,N_1968);
or U3568 (N_3568,N_2489,N_2492);
and U3569 (N_3569,N_1713,N_2924);
xor U3570 (N_3570,N_2322,N_2429);
nor U3571 (N_3571,N_2697,N_2059);
or U3572 (N_3572,N_1670,N_2939);
and U3573 (N_3573,N_2402,N_2289);
xor U3574 (N_3574,N_2453,N_2842);
or U3575 (N_3575,N_2237,N_2932);
xor U3576 (N_3576,N_1635,N_2668);
nor U3577 (N_3577,N_1835,N_2657);
and U3578 (N_3578,N_2741,N_1777);
and U3579 (N_3579,N_2898,N_2182);
nand U3580 (N_3580,N_2756,N_2478);
nor U3581 (N_3581,N_1644,N_2705);
nor U3582 (N_3582,N_1643,N_1560);
xor U3583 (N_3583,N_2963,N_1963);
nor U3584 (N_3584,N_2642,N_1947);
and U3585 (N_3585,N_1588,N_2013);
nand U3586 (N_3586,N_2718,N_2512);
nand U3587 (N_3587,N_2260,N_2298);
nand U3588 (N_3588,N_1811,N_1628);
and U3589 (N_3589,N_1606,N_2710);
or U3590 (N_3590,N_2548,N_2938);
xnor U3591 (N_3591,N_2080,N_2529);
nor U3592 (N_3592,N_2169,N_1629);
nor U3593 (N_3593,N_1831,N_1703);
nor U3594 (N_3594,N_2660,N_2503);
or U3595 (N_3595,N_1590,N_2856);
nand U3596 (N_3596,N_1500,N_2958);
xnor U3597 (N_3597,N_2123,N_1843);
xor U3598 (N_3598,N_2341,N_2934);
xnor U3599 (N_3599,N_2425,N_1600);
nor U3600 (N_3600,N_1649,N_2353);
nor U3601 (N_3601,N_1796,N_2071);
nor U3602 (N_3602,N_2962,N_2249);
nand U3603 (N_3603,N_1584,N_2093);
xnor U3604 (N_3604,N_2876,N_1714);
nand U3605 (N_3605,N_2521,N_2638);
xnor U3606 (N_3606,N_1987,N_2578);
or U3607 (N_3607,N_1622,N_2622);
and U3608 (N_3608,N_2810,N_2479);
xnor U3609 (N_3609,N_2916,N_1712);
nand U3610 (N_3610,N_2204,N_1739);
and U3611 (N_3611,N_2462,N_1857);
nand U3612 (N_3612,N_2285,N_2649);
nor U3613 (N_3613,N_2375,N_2634);
or U3614 (N_3614,N_1543,N_2768);
and U3615 (N_3615,N_2387,N_2495);
nand U3616 (N_3616,N_2774,N_2470);
nor U3617 (N_3617,N_1552,N_2409);
and U3618 (N_3618,N_1803,N_1847);
or U3619 (N_3619,N_1896,N_2382);
or U3620 (N_3620,N_1572,N_1611);
nand U3621 (N_3621,N_1690,N_1554);
or U3622 (N_3622,N_2218,N_2602);
nor U3623 (N_3623,N_1505,N_1676);
nand U3624 (N_3624,N_2337,N_1749);
nand U3625 (N_3625,N_2744,N_2164);
nor U3626 (N_3626,N_2597,N_2035);
or U3627 (N_3627,N_1988,N_1757);
xor U3628 (N_3628,N_2358,N_1817);
nand U3629 (N_3629,N_1527,N_2561);
or U3630 (N_3630,N_2966,N_2278);
nand U3631 (N_3631,N_1881,N_1931);
nand U3632 (N_3632,N_1808,N_2354);
xnor U3633 (N_3633,N_2971,N_1820);
nand U3634 (N_3634,N_2568,N_1583);
xor U3635 (N_3635,N_2601,N_2504);
nor U3636 (N_3636,N_1894,N_2386);
xor U3637 (N_3637,N_2051,N_2268);
nor U3638 (N_3638,N_2933,N_2284);
xor U3639 (N_3639,N_2352,N_2681);
and U3640 (N_3640,N_2198,N_1586);
nor U3641 (N_3641,N_2406,N_1814);
nor U3642 (N_3642,N_2228,N_2716);
and U3643 (N_3643,N_2565,N_2663);
xor U3644 (N_3644,N_2467,N_2257);
nand U3645 (N_3645,N_1901,N_2616);
or U3646 (N_3646,N_1941,N_1694);
nor U3647 (N_3647,N_2664,N_2717);
or U3648 (N_3648,N_1549,N_2941);
and U3649 (N_3649,N_2427,N_2330);
xnor U3650 (N_3650,N_2679,N_1855);
nand U3651 (N_3651,N_2321,N_1823);
or U3652 (N_3652,N_1735,N_1869);
and U3653 (N_3653,N_1787,N_2028);
or U3654 (N_3654,N_2814,N_2780);
nand U3655 (N_3655,N_2443,N_1860);
nor U3656 (N_3656,N_2692,N_2418);
nand U3657 (N_3657,N_2310,N_2614);
xor U3658 (N_3658,N_1578,N_1828);
nor U3659 (N_3659,N_1902,N_1617);
and U3660 (N_3660,N_1889,N_2254);
nor U3661 (N_3661,N_1669,N_2350);
nor U3662 (N_3662,N_2746,N_2918);
nor U3663 (N_3663,N_1717,N_2149);
or U3664 (N_3664,N_1910,N_2465);
xor U3665 (N_3665,N_2584,N_2721);
nand U3666 (N_3666,N_2451,N_1933);
and U3667 (N_3667,N_1579,N_2719);
or U3668 (N_3668,N_2496,N_1525);
xor U3669 (N_3669,N_1672,N_2077);
nor U3670 (N_3670,N_2633,N_1836);
or U3671 (N_3671,N_1545,N_2272);
nand U3672 (N_3672,N_1837,N_1986);
xor U3673 (N_3673,N_2201,N_2509);
nand U3674 (N_3674,N_2156,N_1571);
and U3675 (N_3675,N_2618,N_2684);
and U3676 (N_3676,N_1563,N_2328);
and U3677 (N_3677,N_2037,N_1522);
and U3678 (N_3678,N_2316,N_2587);
or U3679 (N_3679,N_2317,N_2949);
and U3680 (N_3680,N_2242,N_2146);
or U3681 (N_3681,N_2045,N_1908);
xnor U3682 (N_3682,N_2790,N_2621);
nand U3683 (N_3683,N_2841,N_2060);
nor U3684 (N_3684,N_2400,N_2762);
nand U3685 (N_3685,N_2075,N_1867);
nor U3686 (N_3686,N_2850,N_2194);
and U3687 (N_3687,N_2058,N_2757);
and U3688 (N_3688,N_1952,N_1927);
and U3689 (N_3689,N_1638,N_2126);
nand U3690 (N_3690,N_2275,N_1510);
nand U3691 (N_3691,N_2980,N_2708);
nand U3692 (N_3692,N_2090,N_2161);
nor U3693 (N_3693,N_2292,N_2950);
or U3694 (N_3694,N_2742,N_1876);
xor U3695 (N_3695,N_1826,N_2542);
or U3696 (N_3696,N_2553,N_2732);
nand U3697 (N_3697,N_2083,N_1913);
nand U3698 (N_3698,N_2011,N_2015);
xor U3699 (N_3699,N_2997,N_2110);
nand U3700 (N_3700,N_1873,N_2538);
and U3701 (N_3701,N_1848,N_2361);
xor U3702 (N_3702,N_2304,N_2551);
xor U3703 (N_3703,N_2954,N_2216);
and U3704 (N_3704,N_2026,N_2957);
or U3705 (N_3705,N_1725,N_2901);
and U3706 (N_3706,N_2690,N_2178);
or U3707 (N_3707,N_2655,N_2248);
xnor U3708 (N_3708,N_2114,N_2665);
xnor U3709 (N_3709,N_2339,N_2063);
or U3710 (N_3710,N_2629,N_1721);
nor U3711 (N_3711,N_2221,N_2457);
and U3712 (N_3712,N_1792,N_2905);
nand U3713 (N_3713,N_2335,N_2631);
nor U3714 (N_3714,N_1935,N_1911);
xnor U3715 (N_3715,N_1696,N_1634);
xnor U3716 (N_3716,N_1553,N_2389);
and U3717 (N_3717,N_2572,N_2701);
nor U3718 (N_3718,N_1513,N_2524);
and U3719 (N_3719,N_2373,N_2299);
nand U3720 (N_3720,N_2989,N_1700);
nand U3721 (N_3721,N_2357,N_2881);
nor U3722 (N_3722,N_1640,N_2296);
or U3723 (N_3723,N_2371,N_2384);
and U3724 (N_3724,N_2662,N_2312);
and U3725 (N_3725,N_2867,N_1804);
nand U3726 (N_3726,N_1924,N_1566);
xnor U3727 (N_3727,N_2635,N_1905);
xnor U3728 (N_3728,N_2211,N_2472);
xor U3729 (N_3729,N_2137,N_2594);
xnor U3730 (N_3730,N_1998,N_2669);
and U3731 (N_3731,N_2636,N_2213);
nand U3732 (N_3732,N_2760,N_2610);
nand U3733 (N_3733,N_2937,N_2444);
nand U3734 (N_3734,N_1918,N_1772);
xnor U3735 (N_3735,N_1851,N_1815);
nand U3736 (N_3736,N_2858,N_2423);
nand U3737 (N_3737,N_2006,N_2494);
or U3738 (N_3738,N_1750,N_1875);
and U3739 (N_3739,N_1990,N_1742);
nand U3740 (N_3740,N_2988,N_2276);
nor U3741 (N_3741,N_2428,N_2726);
xnor U3742 (N_3742,N_2613,N_2041);
nor U3743 (N_3743,N_2986,N_1508);
nor U3744 (N_3744,N_2546,N_2908);
xnor U3745 (N_3745,N_2115,N_1592);
or U3746 (N_3746,N_2487,N_1718);
nand U3747 (N_3747,N_2647,N_1626);
nor U3748 (N_3748,N_2599,N_1801);
nor U3749 (N_3749,N_2031,N_2230);
nor U3750 (N_3750,N_2329,N_2515);
or U3751 (N_3751,N_2133,N_2806);
and U3752 (N_3752,N_2480,N_1604);
and U3753 (N_3753,N_1577,N_1558);
nor U3754 (N_3754,N_2975,N_2476);
and U3755 (N_3755,N_2420,N_1820);
and U3756 (N_3756,N_2741,N_1766);
xnor U3757 (N_3757,N_1970,N_1763);
nor U3758 (N_3758,N_2275,N_2107);
nor U3759 (N_3759,N_2985,N_2639);
and U3760 (N_3760,N_2216,N_2817);
nor U3761 (N_3761,N_2308,N_2424);
and U3762 (N_3762,N_2574,N_2254);
xor U3763 (N_3763,N_2757,N_2077);
nor U3764 (N_3764,N_2151,N_2295);
nor U3765 (N_3765,N_2721,N_2291);
xor U3766 (N_3766,N_2188,N_2428);
or U3767 (N_3767,N_2252,N_1987);
nand U3768 (N_3768,N_2492,N_2173);
or U3769 (N_3769,N_2153,N_2121);
xnor U3770 (N_3770,N_1512,N_2573);
and U3771 (N_3771,N_1708,N_2940);
nor U3772 (N_3772,N_2753,N_2389);
and U3773 (N_3773,N_2691,N_1669);
nand U3774 (N_3774,N_2325,N_2036);
nor U3775 (N_3775,N_1643,N_1983);
nor U3776 (N_3776,N_1991,N_2652);
nor U3777 (N_3777,N_2332,N_2267);
nand U3778 (N_3778,N_2197,N_2475);
and U3779 (N_3779,N_1674,N_1749);
or U3780 (N_3780,N_1842,N_2897);
or U3781 (N_3781,N_2039,N_2933);
or U3782 (N_3782,N_1732,N_1866);
xnor U3783 (N_3783,N_2785,N_2306);
nand U3784 (N_3784,N_2524,N_1747);
or U3785 (N_3785,N_2458,N_1509);
or U3786 (N_3786,N_2449,N_2099);
or U3787 (N_3787,N_2961,N_1618);
nand U3788 (N_3788,N_1859,N_1896);
and U3789 (N_3789,N_2706,N_2627);
nor U3790 (N_3790,N_2053,N_1707);
xnor U3791 (N_3791,N_2024,N_1751);
and U3792 (N_3792,N_2712,N_2312);
or U3793 (N_3793,N_1601,N_2386);
and U3794 (N_3794,N_2361,N_2876);
nor U3795 (N_3795,N_1765,N_2875);
or U3796 (N_3796,N_2159,N_1692);
nand U3797 (N_3797,N_2839,N_1525);
or U3798 (N_3798,N_1962,N_2252);
nand U3799 (N_3799,N_1816,N_1756);
xor U3800 (N_3800,N_2909,N_2114);
xor U3801 (N_3801,N_2487,N_2079);
or U3802 (N_3802,N_2258,N_2367);
and U3803 (N_3803,N_2430,N_2352);
xor U3804 (N_3804,N_2081,N_2922);
xor U3805 (N_3805,N_1837,N_1708);
and U3806 (N_3806,N_2091,N_2999);
nor U3807 (N_3807,N_2205,N_2675);
nand U3808 (N_3808,N_1818,N_2986);
or U3809 (N_3809,N_2059,N_2565);
nor U3810 (N_3810,N_2736,N_2453);
xnor U3811 (N_3811,N_2530,N_2036);
and U3812 (N_3812,N_2289,N_1688);
nand U3813 (N_3813,N_2451,N_1977);
and U3814 (N_3814,N_2782,N_2180);
nor U3815 (N_3815,N_1902,N_1996);
xnor U3816 (N_3816,N_2666,N_2603);
xor U3817 (N_3817,N_2010,N_1679);
or U3818 (N_3818,N_2956,N_2099);
nor U3819 (N_3819,N_2694,N_2635);
xor U3820 (N_3820,N_1810,N_2637);
or U3821 (N_3821,N_1993,N_2022);
xor U3822 (N_3822,N_1818,N_2554);
nor U3823 (N_3823,N_2502,N_2401);
or U3824 (N_3824,N_1969,N_2403);
or U3825 (N_3825,N_2365,N_2158);
and U3826 (N_3826,N_2141,N_1937);
or U3827 (N_3827,N_2240,N_1647);
nand U3828 (N_3828,N_2089,N_2400);
and U3829 (N_3829,N_2087,N_2215);
or U3830 (N_3830,N_2188,N_2912);
nor U3831 (N_3831,N_1609,N_1748);
and U3832 (N_3832,N_2099,N_2359);
nand U3833 (N_3833,N_2120,N_2506);
or U3834 (N_3834,N_2811,N_2066);
and U3835 (N_3835,N_1568,N_2317);
or U3836 (N_3836,N_2298,N_1687);
xor U3837 (N_3837,N_2222,N_1584);
nor U3838 (N_3838,N_2020,N_1538);
and U3839 (N_3839,N_2860,N_2641);
xnor U3840 (N_3840,N_2331,N_2517);
nor U3841 (N_3841,N_2392,N_1916);
xor U3842 (N_3842,N_1707,N_1702);
nand U3843 (N_3843,N_2557,N_1852);
nor U3844 (N_3844,N_2877,N_2201);
nor U3845 (N_3845,N_2276,N_2998);
xor U3846 (N_3846,N_2396,N_2780);
or U3847 (N_3847,N_2870,N_1837);
or U3848 (N_3848,N_2483,N_2225);
or U3849 (N_3849,N_2821,N_1994);
xnor U3850 (N_3850,N_2717,N_1768);
xor U3851 (N_3851,N_1751,N_1524);
xnor U3852 (N_3852,N_1915,N_2791);
or U3853 (N_3853,N_2368,N_1695);
or U3854 (N_3854,N_1908,N_2607);
or U3855 (N_3855,N_2436,N_1626);
nor U3856 (N_3856,N_2228,N_2668);
xor U3857 (N_3857,N_1922,N_1951);
or U3858 (N_3858,N_2976,N_2762);
nand U3859 (N_3859,N_2744,N_2410);
or U3860 (N_3860,N_2656,N_1561);
and U3861 (N_3861,N_2923,N_1871);
or U3862 (N_3862,N_2952,N_2554);
or U3863 (N_3863,N_2646,N_2699);
and U3864 (N_3864,N_1865,N_1658);
and U3865 (N_3865,N_2652,N_1620);
nand U3866 (N_3866,N_2593,N_2409);
and U3867 (N_3867,N_2368,N_1774);
or U3868 (N_3868,N_2367,N_2399);
xnor U3869 (N_3869,N_2199,N_1988);
xnor U3870 (N_3870,N_2150,N_2379);
nor U3871 (N_3871,N_2331,N_2032);
or U3872 (N_3872,N_1612,N_1691);
nand U3873 (N_3873,N_2593,N_2879);
nand U3874 (N_3874,N_2323,N_2981);
and U3875 (N_3875,N_1695,N_2123);
or U3876 (N_3876,N_1611,N_2942);
xor U3877 (N_3877,N_1739,N_2092);
and U3878 (N_3878,N_1744,N_2406);
and U3879 (N_3879,N_1782,N_1973);
nor U3880 (N_3880,N_1733,N_1692);
nor U3881 (N_3881,N_2994,N_2704);
and U3882 (N_3882,N_2361,N_2921);
or U3883 (N_3883,N_2644,N_2909);
xnor U3884 (N_3884,N_1940,N_2390);
xnor U3885 (N_3885,N_2413,N_1846);
nor U3886 (N_3886,N_2416,N_1881);
or U3887 (N_3887,N_1764,N_2513);
and U3888 (N_3888,N_2945,N_1844);
and U3889 (N_3889,N_2420,N_2800);
nor U3890 (N_3890,N_2411,N_1658);
nor U3891 (N_3891,N_2740,N_2454);
and U3892 (N_3892,N_1543,N_2015);
xnor U3893 (N_3893,N_2102,N_2458);
nor U3894 (N_3894,N_1599,N_2914);
nor U3895 (N_3895,N_2934,N_2782);
and U3896 (N_3896,N_1736,N_1745);
and U3897 (N_3897,N_2151,N_2930);
and U3898 (N_3898,N_1993,N_2305);
nor U3899 (N_3899,N_2764,N_1613);
xor U3900 (N_3900,N_2432,N_2150);
and U3901 (N_3901,N_2803,N_2478);
xnor U3902 (N_3902,N_1839,N_2696);
nand U3903 (N_3903,N_1869,N_2466);
nand U3904 (N_3904,N_1678,N_1551);
nor U3905 (N_3905,N_2080,N_2978);
nor U3906 (N_3906,N_1546,N_2898);
and U3907 (N_3907,N_2222,N_1853);
nand U3908 (N_3908,N_1780,N_2260);
xor U3909 (N_3909,N_1930,N_2772);
nor U3910 (N_3910,N_2825,N_2207);
nand U3911 (N_3911,N_2566,N_2978);
or U3912 (N_3912,N_2806,N_1652);
and U3913 (N_3913,N_1526,N_1955);
xor U3914 (N_3914,N_2557,N_2396);
or U3915 (N_3915,N_2072,N_2361);
or U3916 (N_3916,N_2306,N_1555);
nor U3917 (N_3917,N_2657,N_2327);
or U3918 (N_3918,N_2310,N_1540);
nand U3919 (N_3919,N_1962,N_2817);
or U3920 (N_3920,N_1718,N_1926);
nand U3921 (N_3921,N_2725,N_2457);
and U3922 (N_3922,N_2949,N_1768);
nor U3923 (N_3923,N_2717,N_1926);
xnor U3924 (N_3924,N_1508,N_2855);
nor U3925 (N_3925,N_2051,N_1593);
and U3926 (N_3926,N_2835,N_2037);
or U3927 (N_3927,N_2169,N_2070);
nand U3928 (N_3928,N_2756,N_2121);
and U3929 (N_3929,N_2470,N_2214);
xor U3930 (N_3930,N_1726,N_2400);
nor U3931 (N_3931,N_1603,N_2957);
and U3932 (N_3932,N_1769,N_2079);
nor U3933 (N_3933,N_2816,N_2458);
and U3934 (N_3934,N_2825,N_2536);
nand U3935 (N_3935,N_2101,N_1868);
xor U3936 (N_3936,N_2151,N_2810);
and U3937 (N_3937,N_2471,N_1803);
or U3938 (N_3938,N_2660,N_2510);
or U3939 (N_3939,N_2294,N_1601);
nor U3940 (N_3940,N_2999,N_2480);
nand U3941 (N_3941,N_1512,N_2868);
or U3942 (N_3942,N_1772,N_1707);
nand U3943 (N_3943,N_2865,N_1616);
and U3944 (N_3944,N_2571,N_1790);
nand U3945 (N_3945,N_1645,N_2496);
nand U3946 (N_3946,N_2181,N_2638);
or U3947 (N_3947,N_1647,N_2864);
xor U3948 (N_3948,N_1551,N_2630);
xor U3949 (N_3949,N_1604,N_1652);
or U3950 (N_3950,N_2202,N_2439);
and U3951 (N_3951,N_2482,N_1646);
nand U3952 (N_3952,N_2044,N_1954);
nand U3953 (N_3953,N_2880,N_2700);
and U3954 (N_3954,N_2541,N_1609);
or U3955 (N_3955,N_2289,N_2507);
nand U3956 (N_3956,N_2802,N_2926);
nor U3957 (N_3957,N_2918,N_1787);
nor U3958 (N_3958,N_2213,N_1873);
nand U3959 (N_3959,N_2914,N_2333);
nor U3960 (N_3960,N_1710,N_2654);
or U3961 (N_3961,N_1853,N_1708);
and U3962 (N_3962,N_2811,N_2583);
nand U3963 (N_3963,N_2353,N_2324);
xnor U3964 (N_3964,N_2099,N_1636);
xnor U3965 (N_3965,N_2436,N_2048);
and U3966 (N_3966,N_2698,N_1759);
and U3967 (N_3967,N_1788,N_2057);
or U3968 (N_3968,N_1663,N_1918);
nand U3969 (N_3969,N_2311,N_2706);
or U3970 (N_3970,N_2229,N_1502);
or U3971 (N_3971,N_2281,N_2277);
or U3972 (N_3972,N_1744,N_2049);
and U3973 (N_3973,N_1565,N_2779);
or U3974 (N_3974,N_2449,N_1907);
xor U3975 (N_3975,N_2149,N_2180);
and U3976 (N_3976,N_2125,N_2280);
nor U3977 (N_3977,N_2777,N_2472);
nor U3978 (N_3978,N_2564,N_1823);
and U3979 (N_3979,N_1822,N_1645);
and U3980 (N_3980,N_2776,N_2158);
or U3981 (N_3981,N_1564,N_1536);
and U3982 (N_3982,N_2777,N_2346);
xnor U3983 (N_3983,N_2039,N_2488);
xnor U3984 (N_3984,N_2957,N_2062);
xor U3985 (N_3985,N_2638,N_2603);
and U3986 (N_3986,N_2204,N_2335);
nor U3987 (N_3987,N_2308,N_2404);
xnor U3988 (N_3988,N_2106,N_1573);
and U3989 (N_3989,N_2948,N_2864);
nand U3990 (N_3990,N_1571,N_1791);
nor U3991 (N_3991,N_2422,N_2946);
or U3992 (N_3992,N_2178,N_2209);
xor U3993 (N_3993,N_2860,N_2269);
and U3994 (N_3994,N_2713,N_2209);
nor U3995 (N_3995,N_1748,N_1576);
xor U3996 (N_3996,N_2575,N_1864);
nor U3997 (N_3997,N_2677,N_1786);
nor U3998 (N_3998,N_1727,N_1794);
and U3999 (N_3999,N_2830,N_1701);
nor U4000 (N_4000,N_2561,N_1770);
and U4001 (N_4001,N_2949,N_1793);
nor U4002 (N_4002,N_2488,N_2371);
xnor U4003 (N_4003,N_2701,N_2708);
or U4004 (N_4004,N_1982,N_2164);
and U4005 (N_4005,N_2954,N_2493);
or U4006 (N_4006,N_2235,N_2876);
xor U4007 (N_4007,N_2380,N_2185);
nor U4008 (N_4008,N_2896,N_1565);
or U4009 (N_4009,N_2857,N_2334);
nand U4010 (N_4010,N_1646,N_2364);
xnor U4011 (N_4011,N_2593,N_2602);
nand U4012 (N_4012,N_2238,N_2306);
xnor U4013 (N_4013,N_2482,N_2352);
or U4014 (N_4014,N_2198,N_2891);
nand U4015 (N_4015,N_2467,N_2415);
xor U4016 (N_4016,N_2711,N_2796);
nor U4017 (N_4017,N_2447,N_2524);
or U4018 (N_4018,N_2971,N_1930);
or U4019 (N_4019,N_2927,N_2143);
nor U4020 (N_4020,N_2045,N_2294);
xor U4021 (N_4021,N_2809,N_2610);
and U4022 (N_4022,N_1607,N_2312);
or U4023 (N_4023,N_2187,N_2591);
nand U4024 (N_4024,N_1624,N_1997);
and U4025 (N_4025,N_2979,N_2983);
xor U4026 (N_4026,N_2929,N_1736);
nor U4027 (N_4027,N_2982,N_1750);
and U4028 (N_4028,N_1744,N_2899);
and U4029 (N_4029,N_2740,N_2563);
nor U4030 (N_4030,N_2190,N_2274);
nand U4031 (N_4031,N_2200,N_2247);
or U4032 (N_4032,N_2303,N_1748);
nand U4033 (N_4033,N_2445,N_1585);
nand U4034 (N_4034,N_1991,N_1901);
nand U4035 (N_4035,N_2548,N_2039);
and U4036 (N_4036,N_2871,N_2172);
and U4037 (N_4037,N_2135,N_2266);
nand U4038 (N_4038,N_2910,N_2310);
and U4039 (N_4039,N_2050,N_2188);
or U4040 (N_4040,N_2834,N_1815);
xnor U4041 (N_4041,N_2413,N_2760);
and U4042 (N_4042,N_2038,N_2072);
or U4043 (N_4043,N_2626,N_1745);
and U4044 (N_4044,N_2175,N_1546);
and U4045 (N_4045,N_1607,N_2628);
nor U4046 (N_4046,N_2282,N_1680);
and U4047 (N_4047,N_2716,N_2608);
or U4048 (N_4048,N_2185,N_2045);
or U4049 (N_4049,N_2618,N_2122);
and U4050 (N_4050,N_2582,N_2709);
or U4051 (N_4051,N_1836,N_2864);
xnor U4052 (N_4052,N_2924,N_2144);
xor U4053 (N_4053,N_1724,N_1819);
and U4054 (N_4054,N_2879,N_1777);
xnor U4055 (N_4055,N_2874,N_2700);
nand U4056 (N_4056,N_1714,N_1626);
nor U4057 (N_4057,N_2960,N_1746);
nand U4058 (N_4058,N_2990,N_1786);
xnor U4059 (N_4059,N_2438,N_2646);
nor U4060 (N_4060,N_2225,N_2308);
or U4061 (N_4061,N_2069,N_2570);
and U4062 (N_4062,N_2084,N_1562);
or U4063 (N_4063,N_1603,N_2419);
or U4064 (N_4064,N_1724,N_2325);
and U4065 (N_4065,N_2271,N_2049);
nand U4066 (N_4066,N_2307,N_2816);
nand U4067 (N_4067,N_2827,N_2381);
nor U4068 (N_4068,N_2500,N_2093);
and U4069 (N_4069,N_2343,N_1573);
nand U4070 (N_4070,N_2262,N_2988);
and U4071 (N_4071,N_1646,N_1971);
or U4072 (N_4072,N_2032,N_2756);
nor U4073 (N_4073,N_2368,N_2454);
or U4074 (N_4074,N_1992,N_2728);
or U4075 (N_4075,N_2123,N_2308);
and U4076 (N_4076,N_2509,N_2587);
nand U4077 (N_4077,N_2703,N_1969);
and U4078 (N_4078,N_2265,N_1909);
nor U4079 (N_4079,N_2686,N_2758);
or U4080 (N_4080,N_2396,N_2812);
and U4081 (N_4081,N_2593,N_2967);
nor U4082 (N_4082,N_1543,N_2942);
xor U4083 (N_4083,N_1534,N_2011);
and U4084 (N_4084,N_2850,N_2676);
and U4085 (N_4085,N_2590,N_1590);
xnor U4086 (N_4086,N_1802,N_2380);
nor U4087 (N_4087,N_2522,N_2989);
or U4088 (N_4088,N_2009,N_2514);
and U4089 (N_4089,N_1976,N_1697);
nor U4090 (N_4090,N_1547,N_2992);
nand U4091 (N_4091,N_2421,N_1912);
xnor U4092 (N_4092,N_1786,N_2117);
nor U4093 (N_4093,N_1887,N_2057);
and U4094 (N_4094,N_2250,N_2772);
or U4095 (N_4095,N_2661,N_2093);
and U4096 (N_4096,N_1966,N_2308);
and U4097 (N_4097,N_2952,N_2042);
xnor U4098 (N_4098,N_1556,N_2200);
nor U4099 (N_4099,N_2538,N_2273);
or U4100 (N_4100,N_2706,N_2645);
or U4101 (N_4101,N_2920,N_2549);
xnor U4102 (N_4102,N_2015,N_2995);
nand U4103 (N_4103,N_2732,N_2894);
or U4104 (N_4104,N_2870,N_1846);
nand U4105 (N_4105,N_2735,N_2589);
xnor U4106 (N_4106,N_2636,N_2429);
nor U4107 (N_4107,N_2349,N_2178);
or U4108 (N_4108,N_2663,N_2331);
or U4109 (N_4109,N_2428,N_2707);
nand U4110 (N_4110,N_1743,N_2736);
nor U4111 (N_4111,N_1866,N_1828);
nor U4112 (N_4112,N_2437,N_2523);
xor U4113 (N_4113,N_1675,N_1546);
or U4114 (N_4114,N_2603,N_2816);
xor U4115 (N_4115,N_2092,N_2171);
nor U4116 (N_4116,N_2017,N_2218);
or U4117 (N_4117,N_1846,N_2433);
xnor U4118 (N_4118,N_1771,N_2430);
xor U4119 (N_4119,N_2704,N_2827);
nand U4120 (N_4120,N_1570,N_1673);
nor U4121 (N_4121,N_2663,N_1994);
nor U4122 (N_4122,N_2303,N_2849);
xnor U4123 (N_4123,N_2086,N_2796);
nand U4124 (N_4124,N_2176,N_1517);
xor U4125 (N_4125,N_2241,N_2917);
nand U4126 (N_4126,N_2283,N_2418);
xnor U4127 (N_4127,N_2990,N_2316);
or U4128 (N_4128,N_2113,N_2990);
or U4129 (N_4129,N_1509,N_1559);
or U4130 (N_4130,N_2509,N_1835);
nor U4131 (N_4131,N_2238,N_2278);
nand U4132 (N_4132,N_2289,N_2197);
xnor U4133 (N_4133,N_2013,N_1907);
nand U4134 (N_4134,N_1967,N_2042);
xor U4135 (N_4135,N_2747,N_2962);
and U4136 (N_4136,N_2822,N_2671);
nor U4137 (N_4137,N_1735,N_2840);
nand U4138 (N_4138,N_2708,N_2152);
or U4139 (N_4139,N_2593,N_1644);
or U4140 (N_4140,N_1813,N_2666);
and U4141 (N_4141,N_1987,N_1747);
and U4142 (N_4142,N_2013,N_1892);
or U4143 (N_4143,N_2841,N_2375);
xor U4144 (N_4144,N_1848,N_2999);
and U4145 (N_4145,N_2509,N_1563);
or U4146 (N_4146,N_1833,N_2128);
xnor U4147 (N_4147,N_2880,N_1712);
xnor U4148 (N_4148,N_2300,N_2343);
or U4149 (N_4149,N_1712,N_2456);
nand U4150 (N_4150,N_1620,N_2727);
or U4151 (N_4151,N_2210,N_1830);
and U4152 (N_4152,N_2516,N_2923);
xor U4153 (N_4153,N_1927,N_2213);
xor U4154 (N_4154,N_1955,N_2829);
or U4155 (N_4155,N_2972,N_2748);
xor U4156 (N_4156,N_1900,N_2604);
xnor U4157 (N_4157,N_2844,N_1513);
or U4158 (N_4158,N_2498,N_1621);
xnor U4159 (N_4159,N_1647,N_2484);
and U4160 (N_4160,N_2381,N_2443);
nand U4161 (N_4161,N_2790,N_1749);
and U4162 (N_4162,N_1775,N_2165);
or U4163 (N_4163,N_2597,N_1724);
and U4164 (N_4164,N_2175,N_2598);
or U4165 (N_4165,N_2719,N_2962);
and U4166 (N_4166,N_2380,N_1991);
xnor U4167 (N_4167,N_1942,N_2637);
and U4168 (N_4168,N_2165,N_1862);
nor U4169 (N_4169,N_2739,N_2191);
xor U4170 (N_4170,N_2629,N_2742);
xor U4171 (N_4171,N_2541,N_2293);
xor U4172 (N_4172,N_2231,N_2636);
xnor U4173 (N_4173,N_2009,N_2262);
and U4174 (N_4174,N_1553,N_1980);
xor U4175 (N_4175,N_1523,N_2249);
and U4176 (N_4176,N_1734,N_1865);
and U4177 (N_4177,N_2925,N_2432);
nor U4178 (N_4178,N_2710,N_1980);
nand U4179 (N_4179,N_1834,N_2437);
or U4180 (N_4180,N_2667,N_2896);
xnor U4181 (N_4181,N_2755,N_2820);
nor U4182 (N_4182,N_2743,N_2319);
xnor U4183 (N_4183,N_2013,N_1723);
or U4184 (N_4184,N_2746,N_2151);
nor U4185 (N_4185,N_1614,N_2500);
and U4186 (N_4186,N_2933,N_2101);
xor U4187 (N_4187,N_2184,N_2114);
xor U4188 (N_4188,N_1681,N_2023);
nor U4189 (N_4189,N_2921,N_1723);
nor U4190 (N_4190,N_1956,N_1666);
and U4191 (N_4191,N_1535,N_1941);
nand U4192 (N_4192,N_2584,N_1784);
nor U4193 (N_4193,N_2352,N_2767);
and U4194 (N_4194,N_1912,N_2170);
xnor U4195 (N_4195,N_1963,N_2792);
or U4196 (N_4196,N_1558,N_2740);
and U4197 (N_4197,N_1763,N_1615);
and U4198 (N_4198,N_2922,N_2257);
nand U4199 (N_4199,N_2964,N_2492);
xor U4200 (N_4200,N_2425,N_2412);
nor U4201 (N_4201,N_2394,N_2711);
nand U4202 (N_4202,N_1778,N_1781);
nand U4203 (N_4203,N_1942,N_2535);
and U4204 (N_4204,N_1529,N_1519);
nor U4205 (N_4205,N_1768,N_2171);
xnor U4206 (N_4206,N_2375,N_1541);
or U4207 (N_4207,N_2027,N_1997);
or U4208 (N_4208,N_2951,N_2396);
and U4209 (N_4209,N_2800,N_2176);
xnor U4210 (N_4210,N_2165,N_1813);
and U4211 (N_4211,N_2333,N_2238);
or U4212 (N_4212,N_2740,N_2768);
nor U4213 (N_4213,N_2035,N_2247);
nand U4214 (N_4214,N_1860,N_1833);
and U4215 (N_4215,N_2382,N_1959);
or U4216 (N_4216,N_1794,N_2257);
nor U4217 (N_4217,N_2901,N_1921);
and U4218 (N_4218,N_2166,N_1528);
xnor U4219 (N_4219,N_1611,N_1629);
or U4220 (N_4220,N_2813,N_2970);
or U4221 (N_4221,N_2879,N_2370);
xnor U4222 (N_4222,N_2525,N_2252);
xor U4223 (N_4223,N_2990,N_1711);
or U4224 (N_4224,N_2031,N_2215);
and U4225 (N_4225,N_2566,N_2506);
nor U4226 (N_4226,N_2559,N_1880);
nor U4227 (N_4227,N_2903,N_1823);
xor U4228 (N_4228,N_2692,N_2001);
nand U4229 (N_4229,N_1598,N_2663);
xnor U4230 (N_4230,N_2848,N_2782);
nor U4231 (N_4231,N_2500,N_2756);
nand U4232 (N_4232,N_2411,N_1551);
nand U4233 (N_4233,N_2935,N_2678);
and U4234 (N_4234,N_2707,N_2209);
and U4235 (N_4235,N_1518,N_1981);
or U4236 (N_4236,N_2315,N_2179);
nor U4237 (N_4237,N_1907,N_2638);
nand U4238 (N_4238,N_1511,N_2170);
xor U4239 (N_4239,N_1922,N_1520);
nor U4240 (N_4240,N_1550,N_2546);
nand U4241 (N_4241,N_1697,N_2252);
nor U4242 (N_4242,N_1571,N_1839);
and U4243 (N_4243,N_2541,N_2061);
nand U4244 (N_4244,N_1597,N_2998);
or U4245 (N_4245,N_1871,N_2804);
or U4246 (N_4246,N_2515,N_1617);
or U4247 (N_4247,N_1612,N_2955);
nor U4248 (N_4248,N_1978,N_1706);
nand U4249 (N_4249,N_1744,N_2649);
nand U4250 (N_4250,N_2847,N_2570);
nor U4251 (N_4251,N_2070,N_1657);
and U4252 (N_4252,N_1786,N_1935);
and U4253 (N_4253,N_2996,N_1530);
xor U4254 (N_4254,N_1980,N_2637);
nand U4255 (N_4255,N_2418,N_2847);
and U4256 (N_4256,N_2140,N_2861);
or U4257 (N_4257,N_2697,N_2644);
or U4258 (N_4258,N_2998,N_2805);
nand U4259 (N_4259,N_2497,N_1815);
xnor U4260 (N_4260,N_2571,N_1649);
nand U4261 (N_4261,N_2364,N_1576);
nor U4262 (N_4262,N_2689,N_2337);
nor U4263 (N_4263,N_1584,N_1908);
nand U4264 (N_4264,N_1760,N_2226);
xor U4265 (N_4265,N_1674,N_2393);
nand U4266 (N_4266,N_2650,N_1607);
nor U4267 (N_4267,N_1589,N_2469);
nand U4268 (N_4268,N_2579,N_2532);
nor U4269 (N_4269,N_1829,N_2665);
and U4270 (N_4270,N_2900,N_1738);
nand U4271 (N_4271,N_1777,N_2118);
nor U4272 (N_4272,N_1588,N_2499);
and U4273 (N_4273,N_2597,N_2387);
nor U4274 (N_4274,N_2030,N_1645);
nand U4275 (N_4275,N_2882,N_1826);
or U4276 (N_4276,N_2935,N_2190);
xnor U4277 (N_4277,N_1885,N_2066);
xnor U4278 (N_4278,N_1708,N_2527);
and U4279 (N_4279,N_1974,N_1551);
or U4280 (N_4280,N_2840,N_2167);
nand U4281 (N_4281,N_2679,N_1857);
xor U4282 (N_4282,N_1770,N_2663);
and U4283 (N_4283,N_2635,N_2460);
xnor U4284 (N_4284,N_2037,N_2910);
nor U4285 (N_4285,N_2117,N_2700);
xor U4286 (N_4286,N_2500,N_2309);
or U4287 (N_4287,N_2515,N_2258);
nor U4288 (N_4288,N_1649,N_1729);
and U4289 (N_4289,N_2037,N_2704);
nor U4290 (N_4290,N_1834,N_2432);
nor U4291 (N_4291,N_1985,N_2422);
and U4292 (N_4292,N_1916,N_2489);
nor U4293 (N_4293,N_1503,N_1554);
or U4294 (N_4294,N_2650,N_2118);
nor U4295 (N_4295,N_2175,N_2781);
nand U4296 (N_4296,N_2563,N_2592);
and U4297 (N_4297,N_2170,N_2255);
nand U4298 (N_4298,N_2422,N_1963);
xor U4299 (N_4299,N_2935,N_2867);
nor U4300 (N_4300,N_2491,N_1877);
nor U4301 (N_4301,N_1611,N_1754);
nand U4302 (N_4302,N_1532,N_2953);
xor U4303 (N_4303,N_2729,N_1848);
nand U4304 (N_4304,N_2857,N_2808);
xnor U4305 (N_4305,N_2419,N_2333);
and U4306 (N_4306,N_2151,N_1592);
nor U4307 (N_4307,N_2918,N_1729);
or U4308 (N_4308,N_2142,N_1760);
or U4309 (N_4309,N_2869,N_2574);
xor U4310 (N_4310,N_2427,N_2351);
xnor U4311 (N_4311,N_2231,N_2458);
or U4312 (N_4312,N_2456,N_2861);
nor U4313 (N_4313,N_1557,N_1851);
nand U4314 (N_4314,N_2534,N_2179);
or U4315 (N_4315,N_2078,N_2600);
xnor U4316 (N_4316,N_2433,N_2916);
xnor U4317 (N_4317,N_1922,N_2619);
xnor U4318 (N_4318,N_2567,N_1614);
nor U4319 (N_4319,N_2861,N_2587);
xor U4320 (N_4320,N_2690,N_1729);
and U4321 (N_4321,N_1546,N_1723);
nor U4322 (N_4322,N_2873,N_2772);
and U4323 (N_4323,N_2668,N_2416);
xnor U4324 (N_4324,N_2795,N_2242);
nand U4325 (N_4325,N_2342,N_2034);
or U4326 (N_4326,N_2618,N_2620);
or U4327 (N_4327,N_2286,N_2797);
or U4328 (N_4328,N_2059,N_2003);
xor U4329 (N_4329,N_1792,N_2952);
xnor U4330 (N_4330,N_1834,N_2352);
nor U4331 (N_4331,N_1617,N_2338);
and U4332 (N_4332,N_1636,N_2675);
and U4333 (N_4333,N_2796,N_2469);
and U4334 (N_4334,N_1892,N_2153);
and U4335 (N_4335,N_2136,N_1893);
or U4336 (N_4336,N_2124,N_1714);
xor U4337 (N_4337,N_2827,N_2081);
and U4338 (N_4338,N_1536,N_2646);
xor U4339 (N_4339,N_2658,N_2196);
nand U4340 (N_4340,N_1868,N_2974);
xnor U4341 (N_4341,N_2349,N_1651);
nor U4342 (N_4342,N_2080,N_2161);
or U4343 (N_4343,N_2847,N_1663);
or U4344 (N_4344,N_1753,N_2860);
and U4345 (N_4345,N_2836,N_1615);
nand U4346 (N_4346,N_1612,N_2482);
and U4347 (N_4347,N_2655,N_1593);
and U4348 (N_4348,N_2727,N_2147);
or U4349 (N_4349,N_2032,N_2272);
xor U4350 (N_4350,N_2734,N_2020);
nand U4351 (N_4351,N_2420,N_2187);
and U4352 (N_4352,N_1762,N_2554);
nand U4353 (N_4353,N_2232,N_2014);
and U4354 (N_4354,N_2859,N_1861);
xor U4355 (N_4355,N_2204,N_1968);
and U4356 (N_4356,N_2743,N_2401);
nand U4357 (N_4357,N_2943,N_2242);
nor U4358 (N_4358,N_2683,N_2966);
nor U4359 (N_4359,N_2609,N_1741);
xor U4360 (N_4360,N_1836,N_2229);
xnor U4361 (N_4361,N_2036,N_1509);
nand U4362 (N_4362,N_2191,N_1538);
xnor U4363 (N_4363,N_2388,N_2572);
nand U4364 (N_4364,N_1856,N_1560);
xor U4365 (N_4365,N_2257,N_1887);
and U4366 (N_4366,N_2286,N_1770);
or U4367 (N_4367,N_2723,N_2383);
and U4368 (N_4368,N_2662,N_2416);
and U4369 (N_4369,N_2808,N_2550);
or U4370 (N_4370,N_2584,N_2393);
nand U4371 (N_4371,N_1586,N_2716);
nand U4372 (N_4372,N_2454,N_2854);
nor U4373 (N_4373,N_1936,N_1892);
and U4374 (N_4374,N_2650,N_1567);
and U4375 (N_4375,N_2978,N_2764);
xnor U4376 (N_4376,N_1641,N_2580);
nand U4377 (N_4377,N_1704,N_2230);
nor U4378 (N_4378,N_2697,N_1787);
or U4379 (N_4379,N_2308,N_2644);
or U4380 (N_4380,N_2617,N_1668);
xor U4381 (N_4381,N_2181,N_2288);
xnor U4382 (N_4382,N_1720,N_2669);
xnor U4383 (N_4383,N_2328,N_2762);
nor U4384 (N_4384,N_1500,N_2211);
and U4385 (N_4385,N_2402,N_2444);
xor U4386 (N_4386,N_1979,N_2171);
xnor U4387 (N_4387,N_2708,N_1962);
and U4388 (N_4388,N_2830,N_1570);
nand U4389 (N_4389,N_1951,N_2345);
nand U4390 (N_4390,N_2225,N_2466);
nor U4391 (N_4391,N_2579,N_1706);
or U4392 (N_4392,N_1618,N_1815);
nand U4393 (N_4393,N_2887,N_2531);
nor U4394 (N_4394,N_2509,N_1686);
or U4395 (N_4395,N_2642,N_2074);
nor U4396 (N_4396,N_1966,N_1986);
and U4397 (N_4397,N_1987,N_2391);
xor U4398 (N_4398,N_2076,N_1709);
or U4399 (N_4399,N_2634,N_1762);
and U4400 (N_4400,N_2529,N_1675);
nor U4401 (N_4401,N_1546,N_2814);
or U4402 (N_4402,N_2482,N_2744);
and U4403 (N_4403,N_2203,N_2734);
and U4404 (N_4404,N_2181,N_2084);
xor U4405 (N_4405,N_2915,N_1556);
and U4406 (N_4406,N_1834,N_1754);
nor U4407 (N_4407,N_2379,N_1824);
xor U4408 (N_4408,N_1543,N_1869);
nor U4409 (N_4409,N_2888,N_1825);
nor U4410 (N_4410,N_2084,N_2249);
xor U4411 (N_4411,N_2223,N_2585);
xnor U4412 (N_4412,N_1650,N_1753);
and U4413 (N_4413,N_2303,N_2331);
or U4414 (N_4414,N_1549,N_1581);
or U4415 (N_4415,N_1985,N_2278);
nor U4416 (N_4416,N_2664,N_2586);
nor U4417 (N_4417,N_2813,N_2166);
nor U4418 (N_4418,N_2210,N_2651);
xnor U4419 (N_4419,N_2197,N_2476);
or U4420 (N_4420,N_1906,N_1500);
nor U4421 (N_4421,N_2548,N_1590);
xor U4422 (N_4422,N_1680,N_1849);
nand U4423 (N_4423,N_1828,N_2805);
nand U4424 (N_4424,N_2935,N_1867);
nor U4425 (N_4425,N_2870,N_1897);
nand U4426 (N_4426,N_2595,N_1579);
and U4427 (N_4427,N_2949,N_1503);
or U4428 (N_4428,N_2868,N_2138);
and U4429 (N_4429,N_1595,N_1696);
xor U4430 (N_4430,N_1561,N_2148);
nand U4431 (N_4431,N_2032,N_2800);
nor U4432 (N_4432,N_2054,N_2256);
nor U4433 (N_4433,N_2404,N_2209);
or U4434 (N_4434,N_2930,N_2278);
nor U4435 (N_4435,N_2984,N_2001);
and U4436 (N_4436,N_2655,N_2019);
or U4437 (N_4437,N_2350,N_2512);
nand U4438 (N_4438,N_1532,N_1619);
and U4439 (N_4439,N_2715,N_2690);
and U4440 (N_4440,N_1949,N_1893);
nor U4441 (N_4441,N_2410,N_2731);
nor U4442 (N_4442,N_1900,N_2210);
nor U4443 (N_4443,N_1954,N_2411);
and U4444 (N_4444,N_2043,N_2895);
nor U4445 (N_4445,N_2259,N_2842);
or U4446 (N_4446,N_2928,N_1549);
or U4447 (N_4447,N_1861,N_1894);
or U4448 (N_4448,N_2815,N_1919);
nand U4449 (N_4449,N_1803,N_2942);
nand U4450 (N_4450,N_2959,N_2592);
xor U4451 (N_4451,N_2064,N_2885);
nor U4452 (N_4452,N_1574,N_2136);
nand U4453 (N_4453,N_2143,N_2990);
xnor U4454 (N_4454,N_2996,N_1869);
xor U4455 (N_4455,N_2607,N_2036);
and U4456 (N_4456,N_2971,N_2872);
xnor U4457 (N_4457,N_2152,N_2366);
or U4458 (N_4458,N_2037,N_2865);
and U4459 (N_4459,N_1617,N_1700);
nand U4460 (N_4460,N_2596,N_1791);
and U4461 (N_4461,N_2174,N_1532);
nand U4462 (N_4462,N_2968,N_2581);
nor U4463 (N_4463,N_2884,N_2236);
or U4464 (N_4464,N_2483,N_2227);
or U4465 (N_4465,N_2681,N_2764);
nand U4466 (N_4466,N_2187,N_2763);
xnor U4467 (N_4467,N_2128,N_2168);
nor U4468 (N_4468,N_1692,N_2211);
nor U4469 (N_4469,N_2533,N_2216);
nand U4470 (N_4470,N_2035,N_2955);
nor U4471 (N_4471,N_2810,N_2280);
xor U4472 (N_4472,N_2995,N_2048);
or U4473 (N_4473,N_2494,N_1751);
and U4474 (N_4474,N_2625,N_2302);
and U4475 (N_4475,N_2495,N_1679);
xnor U4476 (N_4476,N_2424,N_2482);
nor U4477 (N_4477,N_2303,N_1618);
and U4478 (N_4478,N_1794,N_2596);
or U4479 (N_4479,N_2704,N_1552);
xor U4480 (N_4480,N_1743,N_2806);
nor U4481 (N_4481,N_1585,N_2267);
nor U4482 (N_4482,N_2493,N_2492);
nor U4483 (N_4483,N_1946,N_2807);
xnor U4484 (N_4484,N_1640,N_2755);
nand U4485 (N_4485,N_1516,N_2768);
xnor U4486 (N_4486,N_2559,N_1727);
nand U4487 (N_4487,N_2956,N_1932);
or U4488 (N_4488,N_2979,N_1634);
or U4489 (N_4489,N_2368,N_1938);
xor U4490 (N_4490,N_1869,N_2195);
or U4491 (N_4491,N_2219,N_2671);
nor U4492 (N_4492,N_2392,N_2703);
nor U4493 (N_4493,N_1570,N_2460);
or U4494 (N_4494,N_2600,N_2327);
and U4495 (N_4495,N_2270,N_2549);
and U4496 (N_4496,N_2275,N_1897);
xnor U4497 (N_4497,N_1530,N_1508);
xnor U4498 (N_4498,N_2299,N_1712);
nor U4499 (N_4499,N_2419,N_2024);
nand U4500 (N_4500,N_4460,N_4495);
or U4501 (N_4501,N_4413,N_3299);
or U4502 (N_4502,N_4210,N_3432);
xor U4503 (N_4503,N_3198,N_3298);
xnor U4504 (N_4504,N_3871,N_3827);
xnor U4505 (N_4505,N_3025,N_3194);
or U4506 (N_4506,N_3884,N_3407);
nor U4507 (N_4507,N_4160,N_3764);
and U4508 (N_4508,N_4230,N_4079);
or U4509 (N_4509,N_4251,N_4362);
or U4510 (N_4510,N_3197,N_4162);
nand U4511 (N_4511,N_3689,N_3623);
xnor U4512 (N_4512,N_4120,N_3000);
or U4513 (N_4513,N_4365,N_4307);
or U4514 (N_4514,N_4014,N_4201);
nand U4515 (N_4515,N_3115,N_4467);
or U4516 (N_4516,N_3011,N_3383);
and U4517 (N_4517,N_4206,N_3727);
nand U4518 (N_4518,N_3139,N_3931);
nand U4519 (N_4519,N_4414,N_4324);
nand U4520 (N_4520,N_3347,N_3962);
nor U4521 (N_4521,N_4381,N_3789);
xnor U4522 (N_4522,N_3022,N_4056);
and U4523 (N_4523,N_4109,N_3142);
and U4524 (N_4524,N_4075,N_3122);
and U4525 (N_4525,N_3326,N_3862);
xnor U4526 (N_4526,N_4156,N_3223);
and U4527 (N_4527,N_3105,N_3372);
nand U4528 (N_4528,N_4435,N_4137);
nand U4529 (N_4529,N_4057,N_3163);
or U4530 (N_4530,N_4419,N_4353);
or U4531 (N_4531,N_4148,N_3265);
or U4532 (N_4532,N_3874,N_3553);
and U4533 (N_4533,N_3751,N_3189);
xor U4534 (N_4534,N_4333,N_4484);
or U4535 (N_4535,N_4012,N_3945);
nand U4536 (N_4536,N_4022,N_3597);
nor U4537 (N_4537,N_4047,N_4299);
and U4538 (N_4538,N_3877,N_4217);
xor U4539 (N_4539,N_3604,N_3841);
nor U4540 (N_4540,N_3733,N_3636);
xor U4541 (N_4541,N_3208,N_3692);
nand U4542 (N_4542,N_4440,N_3735);
and U4543 (N_4543,N_3626,N_3232);
nand U4544 (N_4544,N_3296,N_3001);
nor U4545 (N_4545,N_4049,N_3499);
nor U4546 (N_4546,N_4011,N_4347);
and U4547 (N_4547,N_3271,N_3805);
and U4548 (N_4548,N_3571,N_3206);
xor U4549 (N_4549,N_3849,N_4025);
xnor U4550 (N_4550,N_3095,N_4354);
or U4551 (N_4551,N_4262,N_3450);
or U4552 (N_4552,N_4383,N_3737);
and U4553 (N_4553,N_4259,N_3882);
xnor U4554 (N_4554,N_4301,N_4402);
nand U4555 (N_4555,N_4281,N_4039);
nor U4556 (N_4556,N_4260,N_4395);
nand U4557 (N_4557,N_4078,N_3681);
and U4558 (N_4558,N_3759,N_3244);
nor U4559 (N_4559,N_4265,N_4096);
and U4560 (N_4560,N_3104,N_4300);
or U4561 (N_4561,N_3131,N_3821);
nand U4562 (N_4562,N_3948,N_3778);
xor U4563 (N_4563,N_3595,N_3472);
xor U4564 (N_4564,N_3508,N_3312);
xnor U4565 (N_4565,N_4010,N_3077);
xor U4566 (N_4566,N_3483,N_3140);
and U4567 (N_4567,N_3979,N_3520);
nor U4568 (N_4568,N_3099,N_3182);
xnor U4569 (N_4569,N_3837,N_4352);
or U4570 (N_4570,N_3766,N_4184);
nand U4571 (N_4571,N_4093,N_4181);
nor U4572 (N_4572,N_4406,N_3656);
nand U4573 (N_4573,N_4430,N_4149);
or U4574 (N_4574,N_3944,N_4042);
nand U4575 (N_4575,N_4007,N_3224);
or U4576 (N_4576,N_3678,N_3707);
xor U4577 (N_4577,N_3728,N_3536);
and U4578 (N_4578,N_3988,N_3010);
and U4579 (N_4579,N_3091,N_3240);
xnor U4580 (N_4580,N_3763,N_3101);
and U4581 (N_4581,N_4214,N_4222);
and U4582 (N_4582,N_3014,N_3594);
nor U4583 (N_4583,N_4199,N_3990);
and U4584 (N_4584,N_4094,N_3580);
nor U4585 (N_4585,N_3467,N_3797);
and U4586 (N_4586,N_4375,N_3263);
nor U4587 (N_4587,N_3693,N_3869);
nor U4588 (N_4588,N_3982,N_3034);
nor U4589 (N_4589,N_3523,N_4164);
or U4590 (N_4590,N_4015,N_4297);
nand U4591 (N_4591,N_4445,N_3422);
and U4592 (N_4592,N_4188,N_3225);
and U4593 (N_4593,N_3791,N_4028);
or U4594 (N_4594,N_3270,N_3804);
nand U4595 (N_4595,N_3532,N_3507);
nor U4596 (N_4596,N_3799,N_4331);
nor U4597 (N_4597,N_4397,N_4417);
or U4598 (N_4598,N_4461,N_4146);
nor U4599 (N_4599,N_3753,N_3607);
nand U4600 (N_4600,N_3331,N_3645);
and U4601 (N_4601,N_3284,N_3583);
or U4602 (N_4602,N_4292,N_4338);
nor U4603 (N_4603,N_3860,N_3592);
nor U4604 (N_4604,N_3441,N_3795);
nand U4605 (N_4605,N_3167,N_4437);
nor U4606 (N_4606,N_4498,N_4153);
or U4607 (N_4607,N_4062,N_3842);
or U4608 (N_4608,N_3466,N_3016);
nor U4609 (N_4609,N_4227,N_3458);
nand U4610 (N_4610,N_4169,N_4315);
xnor U4611 (N_4611,N_3309,N_3878);
xnor U4612 (N_4612,N_3713,N_3921);
and U4613 (N_4613,N_3866,N_4104);
nand U4614 (N_4614,N_4409,N_3582);
xnor U4615 (N_4615,N_3323,N_4212);
or U4616 (N_4616,N_3491,N_3541);
nand U4617 (N_4617,N_4316,N_3412);
and U4618 (N_4618,N_4434,N_3625);
nand U4619 (N_4619,N_4091,N_3500);
xor U4620 (N_4620,N_3913,N_3730);
nor U4621 (N_4621,N_3086,N_4166);
xor U4622 (N_4622,N_3694,N_3999);
nand U4623 (N_4623,N_4085,N_3457);
nand U4624 (N_4624,N_3932,N_3983);
and U4625 (N_4625,N_4083,N_4418);
nand U4626 (N_4626,N_4245,N_3629);
xor U4627 (N_4627,N_3285,N_4111);
nor U4628 (N_4628,N_3596,N_4134);
nor U4629 (N_4629,N_3494,N_3665);
xor U4630 (N_4630,N_3202,N_3239);
or U4631 (N_4631,N_3069,N_3120);
nor U4632 (N_4632,N_3760,N_4373);
or U4633 (N_4633,N_3885,N_4102);
or U4634 (N_4634,N_3828,N_3984);
or U4635 (N_4635,N_3961,N_4043);
nor U4636 (N_4636,N_3712,N_3647);
nand U4637 (N_4637,N_3661,N_3745);
xor U4638 (N_4638,N_3369,N_4155);
xor U4639 (N_4639,N_3565,N_3551);
nor U4640 (N_4640,N_4275,N_3406);
nand U4641 (N_4641,N_4340,N_3251);
nand U4642 (N_4642,N_3590,N_3262);
xor U4643 (N_4643,N_3776,N_4186);
nand U4644 (N_4644,N_3168,N_3709);
and U4645 (N_4645,N_4038,N_4220);
or U4646 (N_4646,N_3004,N_3610);
and U4647 (N_4647,N_3429,N_3910);
xor U4648 (N_4648,N_4432,N_3639);
and U4649 (N_4649,N_3030,N_3835);
nor U4650 (N_4650,N_4098,N_3471);
and U4651 (N_4651,N_3688,N_3447);
or U4652 (N_4652,N_3575,N_3855);
or U4653 (N_4653,N_3445,N_4462);
nor U4654 (N_4654,N_3315,N_3181);
or U4655 (N_4655,N_4205,N_3598);
or U4656 (N_4656,N_3492,N_3676);
and U4657 (N_4657,N_3686,N_3246);
or U4658 (N_4658,N_3854,N_4341);
nand U4659 (N_4659,N_3840,N_3859);
nand U4660 (N_4660,N_4448,N_4399);
xnor U4661 (N_4661,N_4369,N_4097);
and U4662 (N_4662,N_3336,N_4031);
or U4663 (N_4663,N_3761,N_3079);
or U4664 (N_4664,N_3547,N_3677);
or U4665 (N_4665,N_3515,N_3964);
or U4666 (N_4666,N_3416,N_3375);
or U4667 (N_4667,N_3527,N_3937);
and U4668 (N_4668,N_4326,N_4150);
xnor U4669 (N_4669,N_4232,N_4286);
or U4670 (N_4670,N_3305,N_3072);
xnor U4671 (N_4671,N_3810,N_3734);
nor U4672 (N_4672,N_3192,N_3891);
or U4673 (N_4673,N_3083,N_3358);
or U4674 (N_4674,N_4284,N_3762);
and U4675 (N_4675,N_3098,N_3679);
nor U4676 (N_4676,N_4351,N_3972);
nor U4677 (N_4677,N_4191,N_3635);
and U4678 (N_4678,N_3749,N_4368);
nor U4679 (N_4679,N_3672,N_3915);
nor U4680 (N_4680,N_3599,N_3478);
xnor U4681 (N_4681,N_3070,N_3360);
and U4682 (N_4682,N_4327,N_3825);
xnor U4683 (N_4683,N_3390,N_4185);
nand U4684 (N_4684,N_4264,N_4363);
and U4685 (N_4685,N_3497,N_3865);
nor U4686 (N_4686,N_3129,N_3603);
or U4687 (N_4687,N_3785,N_3744);
xor U4688 (N_4688,N_4189,N_3411);
or U4689 (N_4689,N_3529,N_4266);
and U4690 (N_4690,N_3796,N_4380);
nor U4691 (N_4691,N_3180,N_3555);
or U4692 (N_4692,N_3593,N_3558);
xor U4693 (N_4693,N_3769,N_3046);
or U4694 (N_4694,N_4103,N_3930);
nor U4695 (N_4695,N_3824,N_3047);
nor U4696 (N_4696,N_3637,N_3158);
or U4697 (N_4697,N_4170,N_3107);
nand U4698 (N_4698,N_4303,N_3027);
or U4699 (N_4699,N_4016,N_3338);
nor U4700 (N_4700,N_4026,N_3628);
nand U4701 (N_4701,N_3489,N_3159);
nand U4702 (N_4702,N_3550,N_3718);
nand U4703 (N_4703,N_3516,N_4329);
nand U4704 (N_4704,N_3442,N_3616);
xor U4705 (N_4705,N_3188,N_3459);
or U4706 (N_4706,N_3666,N_3473);
nor U4707 (N_4707,N_4429,N_3184);
or U4708 (N_4708,N_3461,N_3687);
and U4709 (N_4709,N_4309,N_3266);
xnor U4710 (N_4710,N_3577,N_3738);
nand U4711 (N_4711,N_3278,N_4306);
and U4712 (N_4712,N_3183,N_3141);
nand U4713 (N_4713,N_3370,N_3585);
and U4714 (N_4714,N_3396,N_3199);
nand U4715 (N_4715,N_3094,N_3248);
or U4716 (N_4716,N_4172,N_3886);
and U4717 (N_4717,N_3798,N_4036);
nor U4718 (N_4718,N_3160,N_3684);
nand U4719 (N_4719,N_3916,N_3844);
nor U4720 (N_4720,N_4479,N_3024);
or U4721 (N_4721,N_4377,N_4425);
or U4722 (N_4722,N_3469,N_3561);
nand U4723 (N_4723,N_3235,N_3228);
or U4724 (N_4724,N_3381,N_3674);
nand U4725 (N_4725,N_4229,N_3780);
or U4726 (N_4726,N_3815,N_3301);
xor U4727 (N_4727,N_4051,N_3029);
and U4728 (N_4728,N_3451,N_3905);
nor U4729 (N_4729,N_4454,N_3464);
xor U4730 (N_4730,N_3588,N_4133);
nand U4731 (N_4731,N_3531,N_3090);
xor U4732 (N_4732,N_3272,N_3777);
nor U4733 (N_4733,N_4140,N_4465);
xor U4734 (N_4734,N_4276,N_3956);
or U4735 (N_4735,N_3950,N_3820);
or U4736 (N_4736,N_4261,N_3978);
xor U4737 (N_4737,N_4318,N_4357);
nor U4738 (N_4738,N_3330,N_4482);
nor U4739 (N_4739,N_4001,N_3377);
nand U4740 (N_4740,N_3949,N_3439);
xnor U4741 (N_4741,N_3559,N_4335);
or U4742 (N_4742,N_3606,N_3848);
and U4743 (N_4743,N_3876,N_3624);
and U4744 (N_4744,N_3917,N_3682);
xnor U4745 (N_4745,N_3619,N_3993);
xnor U4746 (N_4746,N_3981,N_3430);
nand U4747 (N_4747,N_3770,N_3426);
or U4748 (N_4748,N_3943,N_3031);
nand U4749 (N_4749,N_4058,N_4302);
and U4750 (N_4750,N_4408,N_4213);
nand U4751 (N_4751,N_4470,N_3229);
or U4752 (N_4752,N_4055,N_3087);
xor U4753 (N_4753,N_3242,N_3097);
or U4754 (N_4754,N_4250,N_3048);
nor U4755 (N_4755,N_4426,N_3307);
nor U4756 (N_4756,N_3273,N_3490);
nand U4757 (N_4757,N_4280,N_3890);
xor U4758 (N_4758,N_3161,N_3925);
and U4759 (N_4759,N_3287,N_3608);
or U4760 (N_4760,N_3379,N_3108);
xnor U4761 (N_4761,N_4438,N_3057);
nor U4762 (N_4762,N_3125,N_3935);
and U4763 (N_4763,N_3843,N_3026);
nor U4764 (N_4764,N_3126,N_3893);
and U4765 (N_4765,N_4486,N_4107);
nor U4766 (N_4766,N_4428,N_3773);
xor U4767 (N_4767,N_3758,N_3234);
xor U4768 (N_4768,N_3657,N_3059);
and U4769 (N_4769,N_4171,N_3190);
nor U4770 (N_4770,N_4138,N_4499);
nand U4771 (N_4771,N_3690,N_3704);
nand U4772 (N_4772,N_3393,N_4494);
and U4773 (N_4773,N_4290,N_4143);
and U4774 (N_4774,N_3040,N_4411);
nor U4775 (N_4775,N_3252,N_3018);
and U4776 (N_4776,N_3389,N_4378);
and U4777 (N_4777,N_4200,N_3186);
nand U4778 (N_4778,N_3339,N_3652);
nor U4779 (N_4779,N_4480,N_3802);
and U4780 (N_4780,N_3264,N_3067);
nand U4781 (N_4781,N_3801,N_4325);
nand U4782 (N_4782,N_3781,N_4060);
nor U4783 (N_4783,N_3172,N_3035);
xor U4784 (N_4784,N_3659,N_3517);
nor U4785 (N_4785,N_3053,N_3669);
or U4786 (N_4786,N_3084,N_4089);
and U4787 (N_4787,N_4223,N_3076);
nand U4788 (N_4788,N_3513,N_4246);
or U4789 (N_4789,N_3443,N_4045);
and U4790 (N_4790,N_3373,N_3038);
nand U4791 (N_4791,N_3691,N_3997);
xnor U4792 (N_4792,N_4456,N_4034);
and U4793 (N_4793,N_3431,N_3554);
or U4794 (N_4794,N_4008,N_3648);
xnor U4795 (N_4795,N_3258,N_4469);
or U4796 (N_4796,N_4219,N_3992);
nor U4797 (N_4797,N_4433,N_3280);
xor U4798 (N_4798,N_3552,N_4404);
xor U4799 (N_4799,N_3775,N_4053);
and U4800 (N_4800,N_3174,N_4044);
nor U4801 (N_4801,N_4386,N_4032);
and U4802 (N_4802,N_4361,N_3415);
nor U4803 (N_4803,N_3498,N_3237);
nand U4804 (N_4804,N_3870,N_3293);
nor U4805 (N_4805,N_3214,N_3875);
and U4806 (N_4806,N_3570,N_4289);
and U4807 (N_4807,N_4348,N_3348);
and U4808 (N_4808,N_3311,N_4350);
nor U4809 (N_4809,N_3154,N_3060);
and U4810 (N_4810,N_3774,N_3427);
and U4811 (N_4811,N_4084,N_4431);
nor U4812 (N_4812,N_4311,N_4124);
xor U4813 (N_4813,N_4203,N_3813);
or U4814 (N_4814,N_4288,N_4236);
xor U4815 (N_4815,N_3574,N_3933);
nand U4816 (N_4816,N_4033,N_4115);
nor U4817 (N_4817,N_3261,N_3725);
or U4818 (N_4818,N_3663,N_3455);
nor U4819 (N_4819,N_4127,N_4447);
xnor U4820 (N_4820,N_4048,N_3465);
or U4821 (N_4821,N_3941,N_3023);
or U4822 (N_4822,N_3642,N_3951);
nor U4823 (N_4823,N_3589,N_4345);
or U4824 (N_4824,N_3534,N_3319);
xor U4825 (N_4825,N_3452,N_3123);
or U4826 (N_4826,N_3146,N_4030);
and U4827 (N_4827,N_4080,N_3542);
nand U4828 (N_4828,N_3392,N_3468);
and U4829 (N_4829,N_3425,N_4403);
nand U4830 (N_4830,N_3936,N_3519);
or U4831 (N_4831,N_3892,N_3074);
nand U4832 (N_4832,N_3803,N_3039);
nand U4833 (N_4833,N_3880,N_3966);
or U4834 (N_4834,N_3327,N_3291);
and U4835 (N_4835,N_4197,N_4215);
nand U4836 (N_4836,N_3852,N_3581);
nor U4837 (N_4837,N_3817,N_3811);
nand U4838 (N_4838,N_3128,N_3446);
xor U4839 (N_4839,N_3524,N_3867);
nor U4840 (N_4840,N_3320,N_3722);
nand U4841 (N_4841,N_3408,N_3740);
nand U4842 (N_4842,N_4196,N_3719);
and U4843 (N_4843,N_3924,N_4393);
and U4844 (N_4844,N_3404,N_3147);
nand U4845 (N_4845,N_3005,N_3476);
xor U4846 (N_4846,N_3475,N_3236);
and U4847 (N_4847,N_4019,N_3349);
xnor U4848 (N_4848,N_3260,N_4366);
xnor U4849 (N_4849,N_4455,N_3721);
nand U4850 (N_4850,N_4151,N_3658);
nor U4851 (N_4851,N_4141,N_3403);
nand U4852 (N_4852,N_4439,N_3112);
or U4853 (N_4853,N_3250,N_3401);
or U4854 (N_4854,N_3012,N_4020);
nand U4855 (N_4855,N_3627,N_3667);
and U4856 (N_4856,N_3953,N_4382);
or U4857 (N_4857,N_4180,N_3479);
nand U4858 (N_4858,N_3530,N_3434);
xor U4859 (N_4859,N_3814,N_4407);
and U4860 (N_4860,N_3217,N_3175);
or U4861 (N_4861,N_3346,N_4334);
or U4862 (N_4862,N_3253,N_3858);
nand U4863 (N_4863,N_4475,N_3153);
xor U4864 (N_4864,N_3711,N_4310);
nor U4865 (N_4865,N_4427,N_3906);
nand U4866 (N_4866,N_4391,N_4167);
nand U4867 (N_4867,N_3831,N_4235);
nand U4868 (N_4868,N_4077,N_3985);
nor U4869 (N_4869,N_3909,N_4464);
or U4870 (N_4870,N_3433,N_3899);
xor U4871 (N_4871,N_3539,N_3103);
nor U4872 (N_4872,N_3958,N_3850);
nor U4873 (N_4873,N_3081,N_3883);
or U4874 (N_4874,N_4194,N_3952);
or U4875 (N_4875,N_4076,N_3823);
nor U4876 (N_4876,N_3423,N_4002);
nand U4877 (N_4877,N_4142,N_3371);
nor U4878 (N_4878,N_3238,N_3093);
nor U4879 (N_4879,N_3474,N_3643);
nand U4880 (N_4880,N_3337,N_3509);
xor U4881 (N_4881,N_4054,N_3367);
and U4882 (N_4882,N_3600,N_3605);
nor U4883 (N_4883,N_4018,N_3230);
or U4884 (N_4884,N_3213,N_3151);
and U4885 (N_4885,N_3673,N_3901);
nor U4886 (N_4886,N_4061,N_3328);
or U4887 (N_4887,N_3556,N_3826);
and U4888 (N_4888,N_3685,N_4446);
nand U4889 (N_4889,N_3792,N_3397);
xor U4890 (N_4890,N_3568,N_3080);
xor U4891 (N_4891,N_3548,N_3856);
nand U4892 (N_4892,N_4123,N_3051);
xnor U4893 (N_4893,N_3481,N_3942);
nor U4894 (N_4894,N_3545,N_3706);
and U4895 (N_4895,N_4270,N_3402);
or U4896 (N_4896,N_3630,N_3382);
nand U4897 (N_4897,N_4256,N_4072);
nand U4898 (N_4898,N_4165,N_3698);
and U4899 (N_4899,N_3839,N_3912);
xnor U4900 (N_4900,N_4394,N_3788);
xor U4901 (N_4901,N_3193,N_3454);
nor U4902 (N_4902,N_3960,N_3584);
nor U4903 (N_4903,N_4159,N_3638);
nand U4904 (N_4904,N_4086,N_4081);
nand U4905 (N_4905,N_3991,N_3655);
nand U4906 (N_4906,N_4005,N_3680);
nand U4907 (N_4907,N_3329,N_3152);
and U4908 (N_4908,N_3830,N_3670);
and U4909 (N_4909,N_4122,N_3954);
nor U4910 (N_4910,N_3365,N_4116);
and U4911 (N_4911,N_3008,N_3085);
or U4912 (N_4912,N_3634,N_3058);
or U4913 (N_4913,N_3286,N_4294);
nor U4914 (N_4914,N_3276,N_3748);
nor U4915 (N_4915,N_3746,N_3487);
xor U4916 (N_4916,N_3613,N_4356);
nor U4917 (N_4917,N_3611,N_3353);
xor U4918 (N_4918,N_3247,N_3340);
nand U4919 (N_4919,N_3173,N_3222);
nand U4920 (N_4920,N_3203,N_3109);
and U4921 (N_4921,N_4332,N_4234);
nand U4922 (N_4922,N_3512,N_3290);
nor U4923 (N_4923,N_4224,N_4412);
and U4924 (N_4924,N_3233,N_3768);
or U4925 (N_4925,N_3926,N_3049);
and U4926 (N_4926,N_4457,N_3786);
and U4927 (N_4927,N_3695,N_4496);
and U4928 (N_4928,N_3563,N_4105);
nand U4929 (N_4929,N_3050,N_3488);
nor U4930 (N_4930,N_4342,N_3310);
nand U4931 (N_4931,N_3259,N_3853);
xor U4932 (N_4932,N_3646,N_4163);
or U4933 (N_4933,N_3662,N_4073);
and U4934 (N_4934,N_4242,N_4070);
nand U4935 (N_4935,N_4291,N_4064);
and U4936 (N_4936,N_3054,N_3755);
or U4937 (N_4937,N_3818,N_4466);
nand U4938 (N_4938,N_3526,N_4158);
or U4939 (N_4939,N_4065,N_3731);
and U4940 (N_4940,N_3480,N_3904);
nand U4941 (N_4941,N_3352,N_4263);
or U4942 (N_4942,N_3650,N_4052);
nor U4943 (N_4943,N_3361,N_3205);
xnor U4944 (N_4944,N_4204,N_4364);
nand U4945 (N_4945,N_3812,N_4313);
nand U4946 (N_4946,N_3052,N_4449);
or U4947 (N_4947,N_3887,N_3207);
nand U4948 (N_4948,N_3649,N_3171);
nor U4949 (N_4949,N_3968,N_3255);
xor U4950 (N_4950,N_4379,N_3573);
and U4951 (N_4951,N_3345,N_4021);
xor U4952 (N_4952,N_3410,N_3089);
and U4953 (N_4953,N_3576,N_3110);
and U4954 (N_4954,N_3918,N_4145);
xnor U4955 (N_4955,N_4237,N_3378);
and U4956 (N_4956,N_4279,N_3946);
or U4957 (N_4957,N_3133,N_3897);
nand U4958 (N_4958,N_3622,N_4257);
and U4959 (N_4959,N_3388,N_4177);
xor U4960 (N_4960,N_3363,N_3518);
xor U4961 (N_4961,N_4241,N_3033);
xnor U4962 (N_4962,N_4240,N_3697);
or U4963 (N_4963,N_3342,N_3021);
or U4964 (N_4964,N_3664,N_3056);
or U4965 (N_4965,N_3137,N_4390);
or U4966 (N_4966,N_4004,N_4298);
or U4967 (N_4967,N_3460,N_4491);
or U4968 (N_4968,N_3463,N_4450);
nand U4969 (N_4969,N_3136,N_3994);
and U4970 (N_4970,N_4385,N_3249);
and U4971 (N_4971,N_3864,N_4154);
nand U4972 (N_4972,N_3438,N_4321);
or U4973 (N_4973,N_4320,N_3861);
nor U4974 (N_4974,N_3975,N_4218);
nor U4975 (N_4975,N_3297,N_3295);
or U4976 (N_4976,N_3809,N_4283);
or U4977 (N_4977,N_4463,N_4040);
and U4978 (N_4978,N_4067,N_4176);
or U4979 (N_4979,N_3782,N_3503);
and U4980 (N_4980,N_3771,N_3394);
or U4981 (N_4981,N_4488,N_3601);
xnor U4982 (N_4982,N_4359,N_3165);
nor U4983 (N_4983,N_3144,N_3857);
nand U4984 (N_4984,N_4175,N_3325);
nand U4985 (N_4985,N_3767,N_3380);
nor U4986 (N_4986,N_3633,N_4346);
and U4987 (N_4987,N_3036,N_4131);
or U4988 (N_4988,N_3088,N_3710);
and U4989 (N_4989,N_4023,N_3341);
nor U4990 (N_4990,N_4211,N_4221);
nand U4991 (N_4991,N_3364,N_3569);
nand U4992 (N_4992,N_4287,N_3176);
or U4993 (N_4993,N_3279,N_3836);
and U4994 (N_4994,N_3743,N_3387);
nand U4995 (N_4995,N_3929,N_3609);
and U4996 (N_4996,N_3113,N_3164);
nand U4997 (N_4997,N_3359,N_4243);
and U4998 (N_4998,N_4187,N_3741);
or U4999 (N_4999,N_3437,N_3787);
nand U5000 (N_5000,N_3567,N_3453);
nor U5001 (N_5001,N_4095,N_3417);
nand U5002 (N_5002,N_4443,N_4207);
and U5003 (N_5003,N_3243,N_3914);
and U5004 (N_5004,N_3169,N_3620);
or U5005 (N_5005,N_4228,N_4349);
or U5006 (N_5006,N_4066,N_3845);
and U5007 (N_5007,N_4136,N_3927);
nor U5008 (N_5008,N_3418,N_3963);
or U5009 (N_5009,N_4247,N_3566);
nand U5010 (N_5010,N_3724,N_3132);
nand U5011 (N_5011,N_3671,N_4490);
nand U5012 (N_5012,N_4305,N_3538);
nor U5013 (N_5013,N_3277,N_3334);
nand U5014 (N_5014,N_3700,N_3544);
or U5015 (N_5015,N_4493,N_3986);
xnor U5016 (N_5016,N_3654,N_4029);
nor U5017 (N_5017,N_3424,N_3409);
and U5018 (N_5018,N_3374,N_3201);
nand U5019 (N_5019,N_4139,N_4147);
and U5020 (N_5020,N_4152,N_3708);
nand U5021 (N_5021,N_4035,N_3391);
and U5022 (N_5022,N_3703,N_3216);
xnor U5023 (N_5023,N_3134,N_4336);
nor U5024 (N_5024,N_3400,N_4144);
nand U5025 (N_5025,N_4238,N_3356);
nor U5026 (N_5026,N_3484,N_4249);
nand U5027 (N_5027,N_3732,N_3324);
nor U5028 (N_5028,N_3449,N_3618);
and U5029 (N_5029,N_3641,N_4476);
xnor U5030 (N_5030,N_4129,N_3384);
or U5031 (N_5031,N_4190,N_3300);
nor U5032 (N_5032,N_3354,N_3332);
or U5033 (N_5033,N_3241,N_3998);
nor U5034 (N_5034,N_4202,N_4339);
or U5035 (N_5035,N_3838,N_3501);
or U5036 (N_5036,N_3579,N_4453);
nand U5037 (N_5037,N_4119,N_3100);
or U5038 (N_5038,N_3267,N_4372);
xnor U5039 (N_5039,N_4239,N_3282);
nor U5040 (N_5040,N_4027,N_4444);
xor U5041 (N_5041,N_4392,N_3974);
and U5042 (N_5042,N_3148,N_4328);
nor U5043 (N_5043,N_3195,N_3533);
nor U5044 (N_5044,N_4082,N_3075);
or U5045 (N_5045,N_3281,N_3042);
or U5046 (N_5046,N_3631,N_4254);
or U5047 (N_5047,N_3955,N_3355);
xor U5048 (N_5048,N_3614,N_3421);
xnor U5049 (N_5049,N_4420,N_4087);
and U5050 (N_5050,N_3398,N_3525);
nand U5051 (N_5051,N_4209,N_3414);
or U5052 (N_5052,N_3834,N_3227);
xnor U5053 (N_5053,N_4135,N_3779);
nor U5054 (N_5054,N_3114,N_3292);
nor U5055 (N_5055,N_3562,N_3226);
nand U5056 (N_5056,N_3902,N_3032);
or U5057 (N_5057,N_4252,N_3940);
xor U5058 (N_5058,N_4273,N_3477);
and U5059 (N_5059,N_3068,N_3510);
or U5060 (N_5060,N_3756,N_3977);
nor U5061 (N_5061,N_3889,N_4225);
nor U5062 (N_5062,N_3017,N_4074);
nor U5063 (N_5063,N_3557,N_3177);
nor U5064 (N_5064,N_3055,N_3683);
and U5065 (N_5065,N_4168,N_3702);
nor U5066 (N_5066,N_3254,N_4106);
or U5067 (N_5067,N_4416,N_3846);
xor U5068 (N_5068,N_4009,N_3969);
xnor U5069 (N_5069,N_4358,N_3313);
or U5070 (N_5070,N_3395,N_4398);
and U5071 (N_5071,N_3747,N_4000);
xor U5072 (N_5072,N_3283,N_4110);
nand U5073 (N_5073,N_4322,N_3757);
nor U5074 (N_5074,N_3653,N_3894);
nor U5075 (N_5075,N_3895,N_4355);
or U5076 (N_5076,N_4489,N_3816);
and U5077 (N_5077,N_4118,N_4013);
and U5078 (N_5078,N_3294,N_3651);
xnor U5079 (N_5079,N_3335,N_3162);
and U5080 (N_5080,N_4126,N_3947);
xnor U5081 (N_5081,N_3317,N_3970);
xor U5082 (N_5082,N_3428,N_4485);
nand U5083 (N_5083,N_3521,N_3420);
xnor U5084 (N_5084,N_4003,N_3275);
and U5085 (N_5085,N_4293,N_4068);
nand U5086 (N_5086,N_3967,N_3806);
nand U5087 (N_5087,N_3037,N_4319);
xor U5088 (N_5088,N_4253,N_3316);
and U5089 (N_5089,N_3485,N_4132);
or U5090 (N_5090,N_3868,N_3019);
nand U5091 (N_5091,N_4088,N_3919);
nor U5092 (N_5092,N_3121,N_4248);
nor U5093 (N_5093,N_3204,N_3833);
and U5094 (N_5094,N_4192,N_3350);
nand U5095 (N_5095,N_3268,N_3435);
or U5096 (N_5096,N_4183,N_4090);
or U5097 (N_5097,N_4268,N_3896);
xnor U5098 (N_5098,N_3179,N_3191);
nor U5099 (N_5099,N_3220,N_3495);
and U5100 (N_5100,N_3211,N_4415);
nor U5101 (N_5101,N_4193,N_4226);
or U5102 (N_5102,N_3765,N_3119);
or U5103 (N_5103,N_3959,N_4312);
nor U5104 (N_5104,N_4474,N_3082);
xor U5105 (N_5105,N_3219,N_3965);
nor U5106 (N_5106,N_3462,N_3288);
nand U5107 (N_5107,N_4125,N_3543);
nand U5108 (N_5108,N_3980,N_4472);
xnor U5109 (N_5109,N_4063,N_4451);
nor U5110 (N_5110,N_3493,N_3009);
nor U5111 (N_5111,N_3822,N_3496);
or U5112 (N_5112,N_3957,N_4244);
xnor U5113 (N_5113,N_4121,N_3602);
or U5114 (N_5114,N_4337,N_3071);
nor U5115 (N_5115,N_3045,N_4317);
nand U5116 (N_5116,N_3092,N_3314);
and U5117 (N_5117,N_3750,N_3898);
or U5118 (N_5118,N_4017,N_3726);
nand U5119 (N_5119,N_3343,N_3696);
and U5120 (N_5120,N_3448,N_3130);
nand U5121 (N_5121,N_3736,N_3578);
or U5122 (N_5122,N_3911,N_3701);
and U5123 (N_5123,N_4113,N_3209);
and U5124 (N_5124,N_3135,N_3705);
nor U5125 (N_5125,N_4216,N_3118);
nor U5126 (N_5126,N_3007,N_4128);
nand U5127 (N_5127,N_3308,N_3073);
nand U5128 (N_5128,N_3020,N_3989);
or U5129 (N_5129,N_3720,N_3399);
nand U5130 (N_5130,N_3043,N_4092);
xor U5131 (N_5131,N_3405,N_3546);
and U5132 (N_5132,N_4304,N_3143);
nor U5133 (N_5133,N_4258,N_3714);
nor U5134 (N_5134,N_4006,N_4272);
and U5135 (N_5135,N_3934,N_3504);
and U5136 (N_5136,N_3549,N_4278);
nand U5137 (N_5137,N_3257,N_4182);
xor U5138 (N_5138,N_3061,N_4400);
or U5139 (N_5139,N_3987,N_3028);
nor U5140 (N_5140,N_4046,N_3540);
or U5141 (N_5141,N_3807,N_3729);
and U5142 (N_5142,N_3514,N_3615);
nand U5143 (N_5143,N_4389,N_3752);
and U5144 (N_5144,N_4376,N_3502);
or U5145 (N_5145,N_3231,N_4423);
nand U5146 (N_5146,N_4492,N_4344);
or U5147 (N_5147,N_3586,N_4101);
nand U5148 (N_5148,N_3863,N_4396);
nand U5149 (N_5149,N_3881,N_3772);
xor U5150 (N_5150,N_4497,N_4360);
nand U5151 (N_5151,N_3304,N_3170);
nand U5152 (N_5152,N_4037,N_3215);
and U5153 (N_5153,N_3888,N_3922);
xor U5154 (N_5154,N_3385,N_3587);
nand U5155 (N_5155,N_3535,N_3715);
nor U5156 (N_5156,N_3939,N_3591);
and U5157 (N_5157,N_3218,N_4388);
nand U5158 (N_5158,N_3794,N_3344);
or U5159 (N_5159,N_4442,N_4459);
and U5160 (N_5160,N_4231,N_3716);
xor U5161 (N_5161,N_4114,N_3907);
or U5162 (N_5162,N_3138,N_3187);
nand U5163 (N_5163,N_3908,N_4477);
or U5164 (N_5164,N_3200,N_3564);
nand U5165 (N_5165,N_4130,N_3819);
and U5166 (N_5166,N_4296,N_4099);
xnor U5167 (N_5167,N_3973,N_3790);
nor U5168 (N_5168,N_3995,N_3063);
xnor U5169 (N_5169,N_3617,N_4255);
and U5170 (N_5170,N_3212,N_3366);
nor U5171 (N_5171,N_3928,N_3376);
nor U5172 (N_5172,N_3274,N_4069);
nand U5173 (N_5173,N_3245,N_3413);
and U5174 (N_5174,N_4405,N_4441);
nor U5175 (N_5175,N_3196,N_3872);
nand U5176 (N_5176,N_3302,N_3116);
xor U5177 (N_5177,N_4371,N_3644);
or U5178 (N_5178,N_4282,N_3511);
or U5179 (N_5179,N_4233,N_3318);
or U5180 (N_5180,N_4174,N_4401);
nor U5181 (N_5181,N_4487,N_3166);
or U5182 (N_5182,N_3124,N_3668);
and U5183 (N_5183,N_3640,N_3793);
and U5184 (N_5184,N_4452,N_3621);
or U5185 (N_5185,N_3436,N_4410);
xor U5186 (N_5186,N_3808,N_3632);
and U5187 (N_5187,N_3041,N_4059);
or U5188 (N_5188,N_4071,N_4050);
or U5189 (N_5189,N_3127,N_3879);
xor U5190 (N_5190,N_3096,N_3013);
xnor U5191 (N_5191,N_4370,N_3221);
nand U5192 (N_5192,N_4269,N_3322);
or U5193 (N_5193,N_3111,N_3783);
xor U5194 (N_5194,N_3155,N_3470);
and U5195 (N_5195,N_3351,N_4367);
and U5196 (N_5196,N_3900,N_3178);
nor U5197 (N_5197,N_4473,N_3537);
or U5198 (N_5198,N_3723,N_4271);
and U5199 (N_5199,N_3976,N_3742);
nor U5200 (N_5200,N_3800,N_4471);
nor U5201 (N_5201,N_4173,N_4208);
nand U5202 (N_5202,N_3066,N_3002);
xnor U5203 (N_5203,N_3362,N_3306);
and U5204 (N_5204,N_3106,N_3660);
nor U5205 (N_5205,N_4330,N_3572);
nor U5206 (N_5206,N_3754,N_3784);
or U5207 (N_5207,N_3185,N_4468);
nand U5208 (N_5208,N_3150,N_3157);
or U5209 (N_5209,N_4108,N_4308);
or U5210 (N_5210,N_4483,N_3612);
or U5211 (N_5211,N_3971,N_3996);
nand U5212 (N_5212,N_3444,N_3333);
xor U5213 (N_5213,N_4436,N_4295);
nor U5214 (N_5214,N_4157,N_4117);
nor U5215 (N_5215,N_3873,N_4421);
nor U5216 (N_5216,N_3015,N_3506);
xnor U5217 (N_5217,N_4100,N_4179);
or U5218 (N_5218,N_4267,N_3832);
nand U5219 (N_5219,N_3102,N_3699);
or U5220 (N_5220,N_3357,N_3923);
or U5221 (N_5221,N_3847,N_3269);
nor U5222 (N_5222,N_4285,N_3065);
xnor U5223 (N_5223,N_3851,N_3062);
and U5224 (N_5224,N_3560,N_4478);
xor U5225 (N_5225,N_3044,N_3078);
nor U5226 (N_5226,N_3003,N_3419);
and U5227 (N_5227,N_3289,N_4458);
nand U5228 (N_5228,N_4112,N_3739);
and U5229 (N_5229,N_3006,N_3321);
nor U5230 (N_5230,N_4387,N_3117);
and U5231 (N_5231,N_3156,N_3903);
nor U5232 (N_5232,N_4314,N_3528);
or U5233 (N_5233,N_4374,N_3829);
nand U5234 (N_5234,N_3440,N_3386);
nor U5235 (N_5235,N_4422,N_3256);
or U5236 (N_5236,N_3717,N_3210);
nand U5237 (N_5237,N_4481,N_3303);
nand U5238 (N_5238,N_3920,N_3675);
or U5239 (N_5239,N_3522,N_4274);
xnor U5240 (N_5240,N_4323,N_3505);
nand U5241 (N_5241,N_3486,N_4041);
nand U5242 (N_5242,N_4178,N_4198);
and U5243 (N_5243,N_3456,N_4024);
xor U5244 (N_5244,N_3149,N_4424);
nor U5245 (N_5245,N_3145,N_3482);
and U5246 (N_5246,N_4384,N_4161);
or U5247 (N_5247,N_3064,N_3368);
xor U5248 (N_5248,N_4195,N_3938);
nor U5249 (N_5249,N_4343,N_4277);
nor U5250 (N_5250,N_4412,N_4289);
or U5251 (N_5251,N_3888,N_4030);
or U5252 (N_5252,N_3263,N_3486);
and U5253 (N_5253,N_4330,N_3543);
nor U5254 (N_5254,N_3268,N_3523);
xnor U5255 (N_5255,N_4344,N_3748);
nand U5256 (N_5256,N_4118,N_3490);
nor U5257 (N_5257,N_3229,N_3896);
and U5258 (N_5258,N_3004,N_3723);
xnor U5259 (N_5259,N_3247,N_4424);
xnor U5260 (N_5260,N_3726,N_3802);
nor U5261 (N_5261,N_4097,N_3719);
xor U5262 (N_5262,N_4327,N_3097);
nor U5263 (N_5263,N_3611,N_3471);
and U5264 (N_5264,N_4255,N_3012);
and U5265 (N_5265,N_4074,N_3096);
and U5266 (N_5266,N_4091,N_3221);
xor U5267 (N_5267,N_3024,N_3896);
and U5268 (N_5268,N_4476,N_3863);
nand U5269 (N_5269,N_4269,N_4218);
and U5270 (N_5270,N_3646,N_3682);
xnor U5271 (N_5271,N_3262,N_4087);
xor U5272 (N_5272,N_3959,N_4320);
nor U5273 (N_5273,N_3136,N_3820);
nand U5274 (N_5274,N_3697,N_3403);
xnor U5275 (N_5275,N_3146,N_3665);
nor U5276 (N_5276,N_3777,N_3468);
or U5277 (N_5277,N_3628,N_3979);
and U5278 (N_5278,N_3466,N_3675);
and U5279 (N_5279,N_3834,N_3296);
nand U5280 (N_5280,N_4216,N_3308);
nor U5281 (N_5281,N_3166,N_3200);
nor U5282 (N_5282,N_3875,N_3251);
xor U5283 (N_5283,N_4195,N_3053);
or U5284 (N_5284,N_3838,N_4410);
or U5285 (N_5285,N_3639,N_4038);
nand U5286 (N_5286,N_3392,N_4320);
nand U5287 (N_5287,N_3951,N_4440);
or U5288 (N_5288,N_3292,N_4313);
nor U5289 (N_5289,N_3415,N_3675);
and U5290 (N_5290,N_3609,N_4242);
nor U5291 (N_5291,N_3420,N_4032);
or U5292 (N_5292,N_3605,N_3505);
xor U5293 (N_5293,N_3314,N_3148);
xnor U5294 (N_5294,N_3448,N_3843);
xor U5295 (N_5295,N_3147,N_3432);
xor U5296 (N_5296,N_3099,N_4416);
or U5297 (N_5297,N_3510,N_3626);
or U5298 (N_5298,N_3167,N_3778);
nor U5299 (N_5299,N_3707,N_4185);
or U5300 (N_5300,N_3280,N_4272);
xnor U5301 (N_5301,N_3615,N_4030);
nand U5302 (N_5302,N_4293,N_3419);
xor U5303 (N_5303,N_3989,N_4109);
nor U5304 (N_5304,N_4119,N_4147);
nor U5305 (N_5305,N_3418,N_3010);
and U5306 (N_5306,N_3828,N_4060);
nor U5307 (N_5307,N_3861,N_3569);
xor U5308 (N_5308,N_4113,N_3770);
xor U5309 (N_5309,N_3157,N_3424);
or U5310 (N_5310,N_3414,N_3380);
or U5311 (N_5311,N_3965,N_4065);
nand U5312 (N_5312,N_3066,N_4278);
nor U5313 (N_5313,N_4143,N_3937);
or U5314 (N_5314,N_3827,N_3208);
xnor U5315 (N_5315,N_3955,N_3404);
nand U5316 (N_5316,N_3322,N_3032);
and U5317 (N_5317,N_3511,N_3179);
or U5318 (N_5318,N_3699,N_3523);
or U5319 (N_5319,N_4027,N_4012);
and U5320 (N_5320,N_3715,N_3579);
and U5321 (N_5321,N_3409,N_3630);
or U5322 (N_5322,N_3280,N_4135);
nor U5323 (N_5323,N_3220,N_3830);
nor U5324 (N_5324,N_4366,N_4367);
or U5325 (N_5325,N_3741,N_3274);
or U5326 (N_5326,N_3179,N_3600);
and U5327 (N_5327,N_3032,N_3877);
nor U5328 (N_5328,N_3143,N_3267);
nand U5329 (N_5329,N_4336,N_3260);
and U5330 (N_5330,N_3763,N_3422);
xor U5331 (N_5331,N_3601,N_3284);
xor U5332 (N_5332,N_3859,N_3590);
nand U5333 (N_5333,N_3059,N_4066);
nand U5334 (N_5334,N_4438,N_3314);
or U5335 (N_5335,N_4435,N_3614);
xor U5336 (N_5336,N_3727,N_3506);
nand U5337 (N_5337,N_3489,N_3493);
nor U5338 (N_5338,N_3586,N_3433);
nand U5339 (N_5339,N_4055,N_4196);
or U5340 (N_5340,N_3518,N_4324);
nor U5341 (N_5341,N_4139,N_3633);
xor U5342 (N_5342,N_3264,N_3913);
or U5343 (N_5343,N_3330,N_3494);
or U5344 (N_5344,N_3805,N_4439);
xnor U5345 (N_5345,N_4426,N_3814);
xor U5346 (N_5346,N_3436,N_3167);
nand U5347 (N_5347,N_3032,N_3335);
xnor U5348 (N_5348,N_3285,N_3876);
nand U5349 (N_5349,N_4359,N_4200);
or U5350 (N_5350,N_4382,N_3204);
or U5351 (N_5351,N_3900,N_4485);
or U5352 (N_5352,N_4466,N_3399);
nor U5353 (N_5353,N_3456,N_4243);
and U5354 (N_5354,N_4039,N_3089);
nand U5355 (N_5355,N_3656,N_3350);
nor U5356 (N_5356,N_4195,N_3683);
and U5357 (N_5357,N_3351,N_4046);
nor U5358 (N_5358,N_3907,N_3915);
nand U5359 (N_5359,N_3774,N_4231);
nand U5360 (N_5360,N_3182,N_3519);
and U5361 (N_5361,N_3492,N_3099);
xnor U5362 (N_5362,N_3670,N_3521);
or U5363 (N_5363,N_4227,N_3620);
and U5364 (N_5364,N_4031,N_4480);
xnor U5365 (N_5365,N_3101,N_4498);
nand U5366 (N_5366,N_3442,N_3095);
and U5367 (N_5367,N_4123,N_3164);
or U5368 (N_5368,N_4212,N_4476);
nor U5369 (N_5369,N_4493,N_3593);
or U5370 (N_5370,N_3834,N_4481);
nor U5371 (N_5371,N_3914,N_4254);
nor U5372 (N_5372,N_3030,N_4435);
and U5373 (N_5373,N_3280,N_3573);
nor U5374 (N_5374,N_4375,N_3432);
nor U5375 (N_5375,N_4028,N_4003);
nand U5376 (N_5376,N_4361,N_4466);
xnor U5377 (N_5377,N_3219,N_3108);
xor U5378 (N_5378,N_4491,N_4029);
nand U5379 (N_5379,N_3027,N_3420);
or U5380 (N_5380,N_3165,N_3870);
nor U5381 (N_5381,N_3446,N_3333);
and U5382 (N_5382,N_4471,N_3889);
nand U5383 (N_5383,N_3964,N_3300);
or U5384 (N_5384,N_4179,N_3338);
xnor U5385 (N_5385,N_3169,N_4092);
or U5386 (N_5386,N_3061,N_3915);
xor U5387 (N_5387,N_3790,N_3898);
nand U5388 (N_5388,N_4392,N_3325);
nor U5389 (N_5389,N_4006,N_3583);
and U5390 (N_5390,N_3587,N_4124);
and U5391 (N_5391,N_4152,N_4431);
or U5392 (N_5392,N_4469,N_3394);
and U5393 (N_5393,N_3186,N_3722);
xor U5394 (N_5394,N_3547,N_4087);
xor U5395 (N_5395,N_4135,N_4412);
and U5396 (N_5396,N_3397,N_4035);
and U5397 (N_5397,N_3384,N_4198);
and U5398 (N_5398,N_3277,N_4022);
and U5399 (N_5399,N_4118,N_3374);
xor U5400 (N_5400,N_4263,N_4356);
nor U5401 (N_5401,N_4402,N_4459);
nand U5402 (N_5402,N_4233,N_3429);
xor U5403 (N_5403,N_3594,N_3920);
and U5404 (N_5404,N_4173,N_4037);
nor U5405 (N_5405,N_3177,N_4168);
nor U5406 (N_5406,N_3755,N_3916);
xor U5407 (N_5407,N_3443,N_4430);
and U5408 (N_5408,N_4000,N_4156);
and U5409 (N_5409,N_3485,N_3821);
nand U5410 (N_5410,N_3006,N_3261);
and U5411 (N_5411,N_4227,N_4024);
or U5412 (N_5412,N_3345,N_3013);
or U5413 (N_5413,N_3446,N_3411);
nand U5414 (N_5414,N_3869,N_3487);
nand U5415 (N_5415,N_3795,N_3679);
nand U5416 (N_5416,N_3034,N_3281);
nand U5417 (N_5417,N_3506,N_3154);
or U5418 (N_5418,N_4297,N_3853);
nand U5419 (N_5419,N_3149,N_3323);
nand U5420 (N_5420,N_4099,N_3898);
or U5421 (N_5421,N_3203,N_4065);
nand U5422 (N_5422,N_3619,N_4152);
nor U5423 (N_5423,N_3447,N_4129);
xnor U5424 (N_5424,N_3790,N_3072);
nand U5425 (N_5425,N_3339,N_3510);
or U5426 (N_5426,N_3047,N_3512);
and U5427 (N_5427,N_3220,N_3899);
nor U5428 (N_5428,N_3059,N_4016);
and U5429 (N_5429,N_4441,N_4348);
nor U5430 (N_5430,N_3908,N_3720);
or U5431 (N_5431,N_3773,N_3471);
nor U5432 (N_5432,N_4436,N_3188);
xor U5433 (N_5433,N_3746,N_3760);
and U5434 (N_5434,N_4368,N_3052);
nand U5435 (N_5435,N_4057,N_3071);
xor U5436 (N_5436,N_3042,N_3151);
xor U5437 (N_5437,N_4010,N_3518);
nor U5438 (N_5438,N_3740,N_3483);
nor U5439 (N_5439,N_3916,N_3607);
nand U5440 (N_5440,N_3740,N_3984);
xor U5441 (N_5441,N_3361,N_4094);
nor U5442 (N_5442,N_3661,N_3667);
xnor U5443 (N_5443,N_3035,N_4489);
nand U5444 (N_5444,N_3200,N_3493);
and U5445 (N_5445,N_4109,N_3554);
and U5446 (N_5446,N_3990,N_3850);
nor U5447 (N_5447,N_3849,N_4152);
nor U5448 (N_5448,N_3639,N_3855);
and U5449 (N_5449,N_3280,N_4278);
or U5450 (N_5450,N_4368,N_3527);
or U5451 (N_5451,N_3584,N_4239);
and U5452 (N_5452,N_4260,N_4455);
and U5453 (N_5453,N_3042,N_4344);
nand U5454 (N_5454,N_3405,N_4062);
nor U5455 (N_5455,N_4066,N_3362);
nand U5456 (N_5456,N_3365,N_3473);
nand U5457 (N_5457,N_4377,N_3516);
nand U5458 (N_5458,N_4021,N_3985);
or U5459 (N_5459,N_3269,N_3550);
and U5460 (N_5460,N_3041,N_4190);
xnor U5461 (N_5461,N_3159,N_3573);
nand U5462 (N_5462,N_4357,N_3447);
or U5463 (N_5463,N_3858,N_4107);
nor U5464 (N_5464,N_3032,N_3149);
or U5465 (N_5465,N_4127,N_4008);
nand U5466 (N_5466,N_3902,N_4090);
or U5467 (N_5467,N_3492,N_4118);
xnor U5468 (N_5468,N_3908,N_4242);
xnor U5469 (N_5469,N_3535,N_4200);
or U5470 (N_5470,N_3763,N_4140);
or U5471 (N_5471,N_3532,N_4424);
and U5472 (N_5472,N_3739,N_4421);
nor U5473 (N_5473,N_3260,N_4153);
nor U5474 (N_5474,N_3849,N_4465);
or U5475 (N_5475,N_3448,N_3437);
xor U5476 (N_5476,N_3706,N_3991);
nand U5477 (N_5477,N_4421,N_4160);
xor U5478 (N_5478,N_3249,N_4002);
nand U5479 (N_5479,N_3084,N_3766);
nand U5480 (N_5480,N_3398,N_4234);
or U5481 (N_5481,N_4140,N_3948);
xnor U5482 (N_5482,N_3256,N_4063);
xnor U5483 (N_5483,N_4057,N_4202);
or U5484 (N_5484,N_4186,N_3712);
and U5485 (N_5485,N_3270,N_3662);
nor U5486 (N_5486,N_4337,N_4344);
nand U5487 (N_5487,N_3512,N_3426);
or U5488 (N_5488,N_3929,N_4180);
or U5489 (N_5489,N_3481,N_3523);
and U5490 (N_5490,N_3165,N_3645);
or U5491 (N_5491,N_3217,N_3253);
or U5492 (N_5492,N_3764,N_4381);
nand U5493 (N_5493,N_4369,N_3384);
xnor U5494 (N_5494,N_3090,N_3426);
nor U5495 (N_5495,N_3358,N_3424);
and U5496 (N_5496,N_3718,N_4324);
and U5497 (N_5497,N_4447,N_3506);
xnor U5498 (N_5498,N_4238,N_4422);
or U5499 (N_5499,N_3677,N_3843);
nand U5500 (N_5500,N_3707,N_4458);
nor U5501 (N_5501,N_4332,N_4285);
or U5502 (N_5502,N_3979,N_4366);
xor U5503 (N_5503,N_3692,N_4327);
or U5504 (N_5504,N_3709,N_3518);
xor U5505 (N_5505,N_3124,N_4126);
xnor U5506 (N_5506,N_3602,N_3765);
and U5507 (N_5507,N_4167,N_4441);
or U5508 (N_5508,N_3641,N_4230);
xnor U5509 (N_5509,N_3569,N_3250);
nand U5510 (N_5510,N_3937,N_3343);
xor U5511 (N_5511,N_3029,N_4245);
nand U5512 (N_5512,N_4290,N_4332);
and U5513 (N_5513,N_3365,N_3848);
or U5514 (N_5514,N_4174,N_4395);
nor U5515 (N_5515,N_4258,N_3405);
or U5516 (N_5516,N_3088,N_3095);
or U5517 (N_5517,N_3505,N_3827);
xnor U5518 (N_5518,N_3259,N_3756);
nor U5519 (N_5519,N_3799,N_3495);
xor U5520 (N_5520,N_4044,N_3348);
nor U5521 (N_5521,N_4342,N_3283);
nand U5522 (N_5522,N_3382,N_4419);
or U5523 (N_5523,N_3184,N_3660);
nand U5524 (N_5524,N_3094,N_3851);
nand U5525 (N_5525,N_3841,N_4187);
or U5526 (N_5526,N_3006,N_3185);
xnor U5527 (N_5527,N_3354,N_3216);
and U5528 (N_5528,N_3583,N_3451);
or U5529 (N_5529,N_3912,N_3204);
nand U5530 (N_5530,N_4399,N_3919);
nor U5531 (N_5531,N_3274,N_4051);
nand U5532 (N_5532,N_4042,N_3779);
and U5533 (N_5533,N_4006,N_4473);
and U5534 (N_5534,N_3378,N_3043);
and U5535 (N_5535,N_3088,N_4054);
nor U5536 (N_5536,N_3029,N_3490);
nor U5537 (N_5537,N_4046,N_3828);
and U5538 (N_5538,N_3757,N_4177);
xor U5539 (N_5539,N_3120,N_3067);
or U5540 (N_5540,N_3196,N_3528);
or U5541 (N_5541,N_3499,N_3674);
nor U5542 (N_5542,N_3656,N_3401);
xor U5543 (N_5543,N_3377,N_3560);
and U5544 (N_5544,N_3027,N_3992);
or U5545 (N_5545,N_3449,N_3632);
xor U5546 (N_5546,N_3113,N_4099);
nor U5547 (N_5547,N_3545,N_3229);
xnor U5548 (N_5548,N_4209,N_4483);
nand U5549 (N_5549,N_3908,N_3300);
and U5550 (N_5550,N_3648,N_3430);
and U5551 (N_5551,N_4329,N_3509);
nand U5552 (N_5552,N_3317,N_3493);
or U5553 (N_5553,N_3454,N_3934);
or U5554 (N_5554,N_4403,N_3305);
and U5555 (N_5555,N_3358,N_3888);
and U5556 (N_5556,N_4148,N_3880);
nor U5557 (N_5557,N_3149,N_4216);
nor U5558 (N_5558,N_3901,N_3411);
and U5559 (N_5559,N_4390,N_4430);
nand U5560 (N_5560,N_3304,N_3102);
or U5561 (N_5561,N_3084,N_4171);
nor U5562 (N_5562,N_3630,N_3112);
and U5563 (N_5563,N_3234,N_3005);
nor U5564 (N_5564,N_3069,N_3111);
nand U5565 (N_5565,N_4489,N_3160);
nand U5566 (N_5566,N_4455,N_3963);
nor U5567 (N_5567,N_3468,N_4277);
xnor U5568 (N_5568,N_3599,N_3304);
or U5569 (N_5569,N_4453,N_4004);
nand U5570 (N_5570,N_4052,N_4339);
xor U5571 (N_5571,N_4187,N_3369);
and U5572 (N_5572,N_4402,N_4167);
xor U5573 (N_5573,N_3831,N_3642);
xor U5574 (N_5574,N_3017,N_4437);
nand U5575 (N_5575,N_4007,N_3722);
and U5576 (N_5576,N_4022,N_3214);
nand U5577 (N_5577,N_3088,N_3017);
xor U5578 (N_5578,N_4113,N_3134);
or U5579 (N_5579,N_3976,N_4387);
or U5580 (N_5580,N_3924,N_4332);
or U5581 (N_5581,N_3215,N_4460);
and U5582 (N_5582,N_3737,N_3577);
nor U5583 (N_5583,N_3493,N_4136);
and U5584 (N_5584,N_3450,N_3249);
or U5585 (N_5585,N_3470,N_3432);
nor U5586 (N_5586,N_4499,N_4052);
nand U5587 (N_5587,N_3921,N_3972);
and U5588 (N_5588,N_3487,N_3199);
nor U5589 (N_5589,N_3201,N_4098);
or U5590 (N_5590,N_4088,N_4112);
and U5591 (N_5591,N_3279,N_4351);
nor U5592 (N_5592,N_4173,N_3723);
xor U5593 (N_5593,N_4310,N_3059);
and U5594 (N_5594,N_4408,N_3044);
and U5595 (N_5595,N_3316,N_4334);
and U5596 (N_5596,N_3819,N_3303);
nor U5597 (N_5597,N_4357,N_3005);
xnor U5598 (N_5598,N_3369,N_4308);
and U5599 (N_5599,N_3718,N_3811);
or U5600 (N_5600,N_3881,N_3792);
or U5601 (N_5601,N_4324,N_3528);
and U5602 (N_5602,N_3683,N_3503);
nand U5603 (N_5603,N_4172,N_3977);
nand U5604 (N_5604,N_4077,N_4011);
and U5605 (N_5605,N_4262,N_4083);
and U5606 (N_5606,N_4418,N_3005);
and U5607 (N_5607,N_3019,N_3797);
or U5608 (N_5608,N_4145,N_4362);
nand U5609 (N_5609,N_3493,N_3531);
and U5610 (N_5610,N_4207,N_3974);
and U5611 (N_5611,N_3015,N_3082);
nand U5612 (N_5612,N_3226,N_3412);
xor U5613 (N_5613,N_4093,N_4368);
nand U5614 (N_5614,N_4389,N_3830);
nor U5615 (N_5615,N_4368,N_3978);
nand U5616 (N_5616,N_4436,N_4169);
nand U5617 (N_5617,N_3350,N_3900);
nor U5618 (N_5618,N_3358,N_3192);
nor U5619 (N_5619,N_3143,N_3056);
nor U5620 (N_5620,N_4003,N_3941);
nand U5621 (N_5621,N_3310,N_4318);
and U5622 (N_5622,N_3654,N_3656);
nand U5623 (N_5623,N_4282,N_3930);
and U5624 (N_5624,N_3605,N_3611);
xnor U5625 (N_5625,N_4000,N_3956);
nand U5626 (N_5626,N_3466,N_3364);
nand U5627 (N_5627,N_4496,N_3108);
nor U5628 (N_5628,N_3397,N_3769);
nand U5629 (N_5629,N_3347,N_3769);
or U5630 (N_5630,N_3942,N_4390);
xor U5631 (N_5631,N_3708,N_3110);
xnor U5632 (N_5632,N_3646,N_3339);
and U5633 (N_5633,N_3203,N_3837);
nand U5634 (N_5634,N_3582,N_3030);
and U5635 (N_5635,N_3788,N_3781);
nand U5636 (N_5636,N_3612,N_3040);
nand U5637 (N_5637,N_4186,N_3933);
and U5638 (N_5638,N_3851,N_4272);
nand U5639 (N_5639,N_3336,N_3647);
or U5640 (N_5640,N_3729,N_3401);
or U5641 (N_5641,N_3026,N_3512);
or U5642 (N_5642,N_4187,N_4169);
and U5643 (N_5643,N_3232,N_3168);
or U5644 (N_5644,N_4436,N_4049);
and U5645 (N_5645,N_3103,N_3040);
nor U5646 (N_5646,N_3407,N_4303);
xor U5647 (N_5647,N_3919,N_3190);
xnor U5648 (N_5648,N_3053,N_3825);
or U5649 (N_5649,N_3964,N_3861);
xnor U5650 (N_5650,N_3048,N_4229);
nor U5651 (N_5651,N_3177,N_3643);
nand U5652 (N_5652,N_3812,N_3036);
or U5653 (N_5653,N_4173,N_4445);
xor U5654 (N_5654,N_3436,N_4098);
nand U5655 (N_5655,N_4011,N_3158);
xor U5656 (N_5656,N_4445,N_3989);
nand U5657 (N_5657,N_3094,N_3005);
nor U5658 (N_5658,N_3164,N_3096);
nand U5659 (N_5659,N_4364,N_3776);
nor U5660 (N_5660,N_3150,N_4361);
or U5661 (N_5661,N_3332,N_4352);
and U5662 (N_5662,N_3794,N_3401);
or U5663 (N_5663,N_3187,N_3949);
nand U5664 (N_5664,N_3912,N_4073);
or U5665 (N_5665,N_4489,N_3443);
xnor U5666 (N_5666,N_3634,N_3670);
nand U5667 (N_5667,N_3082,N_3588);
nand U5668 (N_5668,N_3324,N_4350);
nor U5669 (N_5669,N_3525,N_3891);
or U5670 (N_5670,N_4333,N_3071);
and U5671 (N_5671,N_3759,N_4401);
nor U5672 (N_5672,N_3822,N_3226);
nor U5673 (N_5673,N_3490,N_4351);
nor U5674 (N_5674,N_4070,N_3130);
or U5675 (N_5675,N_3338,N_3775);
nand U5676 (N_5676,N_3980,N_3920);
nor U5677 (N_5677,N_3419,N_3290);
or U5678 (N_5678,N_3754,N_4424);
and U5679 (N_5679,N_3532,N_3669);
nand U5680 (N_5680,N_3439,N_4216);
nand U5681 (N_5681,N_4316,N_3563);
xor U5682 (N_5682,N_4139,N_3598);
xnor U5683 (N_5683,N_3831,N_3931);
nor U5684 (N_5684,N_3659,N_3658);
or U5685 (N_5685,N_3992,N_3531);
or U5686 (N_5686,N_3169,N_3035);
nand U5687 (N_5687,N_3923,N_3822);
or U5688 (N_5688,N_4310,N_3549);
nor U5689 (N_5689,N_3117,N_3637);
or U5690 (N_5690,N_3046,N_3059);
nor U5691 (N_5691,N_3324,N_3274);
and U5692 (N_5692,N_4168,N_3086);
nor U5693 (N_5693,N_4391,N_4042);
nor U5694 (N_5694,N_3180,N_3953);
nand U5695 (N_5695,N_4477,N_3898);
xor U5696 (N_5696,N_3344,N_4289);
xnor U5697 (N_5697,N_3454,N_3357);
nand U5698 (N_5698,N_4327,N_3186);
nor U5699 (N_5699,N_3244,N_4284);
xor U5700 (N_5700,N_3776,N_3815);
or U5701 (N_5701,N_3079,N_3310);
nor U5702 (N_5702,N_4100,N_4325);
nand U5703 (N_5703,N_3146,N_4369);
nor U5704 (N_5704,N_3303,N_4313);
or U5705 (N_5705,N_4020,N_4153);
and U5706 (N_5706,N_3089,N_3095);
and U5707 (N_5707,N_3706,N_3481);
nand U5708 (N_5708,N_3852,N_4238);
nand U5709 (N_5709,N_4173,N_3154);
nand U5710 (N_5710,N_4463,N_4357);
or U5711 (N_5711,N_3442,N_3921);
or U5712 (N_5712,N_3864,N_4415);
nand U5713 (N_5713,N_4069,N_3980);
and U5714 (N_5714,N_3648,N_3336);
and U5715 (N_5715,N_4059,N_4284);
nand U5716 (N_5716,N_3574,N_4266);
or U5717 (N_5717,N_3128,N_3844);
nand U5718 (N_5718,N_3396,N_3138);
nand U5719 (N_5719,N_3385,N_3934);
xor U5720 (N_5720,N_3834,N_4092);
nand U5721 (N_5721,N_4066,N_3075);
xnor U5722 (N_5722,N_3118,N_3973);
nor U5723 (N_5723,N_4202,N_3654);
or U5724 (N_5724,N_3433,N_3888);
xor U5725 (N_5725,N_4246,N_3505);
xnor U5726 (N_5726,N_3691,N_3950);
and U5727 (N_5727,N_3746,N_4197);
or U5728 (N_5728,N_3012,N_3900);
nor U5729 (N_5729,N_3540,N_3870);
xnor U5730 (N_5730,N_4327,N_3377);
or U5731 (N_5731,N_3526,N_4180);
xnor U5732 (N_5732,N_4223,N_3899);
xnor U5733 (N_5733,N_4212,N_3508);
or U5734 (N_5734,N_3541,N_4256);
xnor U5735 (N_5735,N_3753,N_3168);
or U5736 (N_5736,N_3495,N_3176);
nor U5737 (N_5737,N_4103,N_3627);
xor U5738 (N_5738,N_4364,N_4046);
and U5739 (N_5739,N_3623,N_3804);
or U5740 (N_5740,N_4342,N_3402);
nor U5741 (N_5741,N_3290,N_4432);
and U5742 (N_5742,N_3996,N_4486);
nand U5743 (N_5743,N_4402,N_3022);
and U5744 (N_5744,N_3862,N_3473);
nor U5745 (N_5745,N_4495,N_4312);
and U5746 (N_5746,N_4363,N_3377);
and U5747 (N_5747,N_4375,N_3780);
xnor U5748 (N_5748,N_3361,N_3003);
xnor U5749 (N_5749,N_3152,N_3637);
or U5750 (N_5750,N_3264,N_3883);
and U5751 (N_5751,N_3539,N_3117);
and U5752 (N_5752,N_4342,N_3568);
or U5753 (N_5753,N_3907,N_3561);
xnor U5754 (N_5754,N_4469,N_4423);
nand U5755 (N_5755,N_3682,N_4225);
nand U5756 (N_5756,N_4108,N_3293);
nor U5757 (N_5757,N_4158,N_3888);
and U5758 (N_5758,N_4265,N_4019);
nand U5759 (N_5759,N_3065,N_3055);
nor U5760 (N_5760,N_4183,N_4068);
xor U5761 (N_5761,N_4288,N_4183);
nor U5762 (N_5762,N_4053,N_3958);
nand U5763 (N_5763,N_3407,N_3457);
and U5764 (N_5764,N_3858,N_3023);
nor U5765 (N_5765,N_3619,N_4437);
and U5766 (N_5766,N_4425,N_4133);
and U5767 (N_5767,N_3983,N_3326);
and U5768 (N_5768,N_3894,N_4095);
or U5769 (N_5769,N_3543,N_4179);
nand U5770 (N_5770,N_4111,N_3583);
or U5771 (N_5771,N_4097,N_3843);
nand U5772 (N_5772,N_4036,N_4431);
nand U5773 (N_5773,N_3674,N_4201);
nand U5774 (N_5774,N_3124,N_4135);
nor U5775 (N_5775,N_3862,N_3810);
nor U5776 (N_5776,N_3266,N_4336);
nand U5777 (N_5777,N_4190,N_3234);
xnor U5778 (N_5778,N_4443,N_3121);
nand U5779 (N_5779,N_3242,N_3180);
nor U5780 (N_5780,N_4310,N_3698);
or U5781 (N_5781,N_4480,N_4319);
nor U5782 (N_5782,N_3397,N_3483);
and U5783 (N_5783,N_3645,N_4094);
nand U5784 (N_5784,N_3891,N_4405);
xor U5785 (N_5785,N_4050,N_4438);
and U5786 (N_5786,N_3840,N_3110);
xnor U5787 (N_5787,N_4325,N_3590);
nor U5788 (N_5788,N_3063,N_3613);
or U5789 (N_5789,N_4374,N_4235);
or U5790 (N_5790,N_3114,N_3402);
nor U5791 (N_5791,N_3380,N_4025);
nand U5792 (N_5792,N_3093,N_4471);
or U5793 (N_5793,N_4004,N_4016);
xor U5794 (N_5794,N_3310,N_3622);
and U5795 (N_5795,N_4177,N_4488);
nor U5796 (N_5796,N_4014,N_3226);
nor U5797 (N_5797,N_3608,N_3239);
nand U5798 (N_5798,N_3174,N_4067);
xnor U5799 (N_5799,N_3689,N_3513);
and U5800 (N_5800,N_3171,N_4366);
or U5801 (N_5801,N_3824,N_3360);
nand U5802 (N_5802,N_3943,N_3905);
nor U5803 (N_5803,N_4184,N_3972);
or U5804 (N_5804,N_4103,N_4183);
nor U5805 (N_5805,N_3084,N_3650);
xnor U5806 (N_5806,N_3980,N_4269);
or U5807 (N_5807,N_4353,N_3732);
and U5808 (N_5808,N_3051,N_4306);
nor U5809 (N_5809,N_4298,N_3188);
or U5810 (N_5810,N_4426,N_3044);
or U5811 (N_5811,N_3465,N_4049);
and U5812 (N_5812,N_4245,N_4411);
nand U5813 (N_5813,N_3858,N_4229);
nand U5814 (N_5814,N_3687,N_4221);
or U5815 (N_5815,N_3562,N_3037);
and U5816 (N_5816,N_4090,N_3259);
nor U5817 (N_5817,N_3624,N_3270);
and U5818 (N_5818,N_3088,N_4254);
xnor U5819 (N_5819,N_3936,N_3001);
xnor U5820 (N_5820,N_4312,N_4065);
or U5821 (N_5821,N_3669,N_3117);
xnor U5822 (N_5822,N_3760,N_4091);
xnor U5823 (N_5823,N_3470,N_4441);
nor U5824 (N_5824,N_3846,N_3931);
xnor U5825 (N_5825,N_3224,N_3337);
or U5826 (N_5826,N_3967,N_3096);
nor U5827 (N_5827,N_4064,N_4358);
nand U5828 (N_5828,N_3002,N_3444);
nor U5829 (N_5829,N_3368,N_3782);
or U5830 (N_5830,N_3835,N_3207);
nand U5831 (N_5831,N_3509,N_3952);
nand U5832 (N_5832,N_3809,N_3737);
nor U5833 (N_5833,N_4090,N_3274);
nand U5834 (N_5834,N_3806,N_3247);
or U5835 (N_5835,N_4275,N_3750);
and U5836 (N_5836,N_4307,N_3036);
and U5837 (N_5837,N_3463,N_3251);
or U5838 (N_5838,N_4232,N_3702);
xor U5839 (N_5839,N_4432,N_3495);
nor U5840 (N_5840,N_3212,N_3684);
xnor U5841 (N_5841,N_3461,N_3137);
or U5842 (N_5842,N_3124,N_3896);
xor U5843 (N_5843,N_4062,N_3107);
or U5844 (N_5844,N_3521,N_3780);
and U5845 (N_5845,N_4238,N_3040);
xnor U5846 (N_5846,N_3778,N_3659);
and U5847 (N_5847,N_4365,N_3774);
or U5848 (N_5848,N_4028,N_4170);
nand U5849 (N_5849,N_3750,N_3534);
nor U5850 (N_5850,N_3016,N_3867);
nand U5851 (N_5851,N_3087,N_3478);
nand U5852 (N_5852,N_3434,N_4078);
nor U5853 (N_5853,N_3192,N_4161);
nor U5854 (N_5854,N_3067,N_3040);
and U5855 (N_5855,N_3482,N_3532);
or U5856 (N_5856,N_4121,N_4233);
and U5857 (N_5857,N_3253,N_4386);
and U5858 (N_5858,N_3807,N_3270);
nor U5859 (N_5859,N_4355,N_3614);
or U5860 (N_5860,N_3221,N_3293);
or U5861 (N_5861,N_4273,N_3790);
xnor U5862 (N_5862,N_3985,N_3143);
and U5863 (N_5863,N_3645,N_3221);
nor U5864 (N_5864,N_3332,N_3616);
or U5865 (N_5865,N_3232,N_3107);
nand U5866 (N_5866,N_4228,N_3493);
and U5867 (N_5867,N_4323,N_3674);
and U5868 (N_5868,N_4223,N_3021);
nand U5869 (N_5869,N_3595,N_4117);
or U5870 (N_5870,N_4207,N_3809);
nor U5871 (N_5871,N_4208,N_3510);
and U5872 (N_5872,N_4305,N_4047);
xor U5873 (N_5873,N_4132,N_4025);
nand U5874 (N_5874,N_3695,N_4475);
xnor U5875 (N_5875,N_3065,N_3592);
xnor U5876 (N_5876,N_4331,N_3335);
nor U5877 (N_5877,N_3530,N_3462);
xnor U5878 (N_5878,N_4291,N_3759);
xnor U5879 (N_5879,N_3436,N_3935);
xnor U5880 (N_5880,N_4128,N_4099);
nor U5881 (N_5881,N_3852,N_3164);
or U5882 (N_5882,N_4030,N_4193);
or U5883 (N_5883,N_4136,N_4265);
and U5884 (N_5884,N_3257,N_3941);
nor U5885 (N_5885,N_3838,N_3895);
and U5886 (N_5886,N_3574,N_4094);
nor U5887 (N_5887,N_4235,N_3827);
nand U5888 (N_5888,N_3328,N_3537);
or U5889 (N_5889,N_4464,N_4050);
xnor U5890 (N_5890,N_3334,N_3736);
and U5891 (N_5891,N_3877,N_3681);
nand U5892 (N_5892,N_4056,N_3875);
nand U5893 (N_5893,N_4384,N_3509);
or U5894 (N_5894,N_3166,N_4003);
and U5895 (N_5895,N_4086,N_4116);
nor U5896 (N_5896,N_3393,N_4188);
xnor U5897 (N_5897,N_4255,N_3927);
nand U5898 (N_5898,N_3113,N_4029);
or U5899 (N_5899,N_3340,N_4445);
nand U5900 (N_5900,N_4422,N_3005);
xor U5901 (N_5901,N_3886,N_3115);
and U5902 (N_5902,N_3302,N_3363);
nor U5903 (N_5903,N_3801,N_4002);
nand U5904 (N_5904,N_3178,N_4136);
and U5905 (N_5905,N_3507,N_3264);
nand U5906 (N_5906,N_3808,N_3684);
nor U5907 (N_5907,N_4225,N_3200);
or U5908 (N_5908,N_4414,N_3269);
or U5909 (N_5909,N_4107,N_4132);
and U5910 (N_5910,N_3689,N_3934);
nand U5911 (N_5911,N_4495,N_3693);
and U5912 (N_5912,N_3332,N_3637);
and U5913 (N_5913,N_3034,N_3633);
or U5914 (N_5914,N_3282,N_4339);
and U5915 (N_5915,N_3095,N_3059);
nor U5916 (N_5916,N_3807,N_4429);
nand U5917 (N_5917,N_3660,N_4231);
xor U5918 (N_5918,N_3752,N_3511);
nand U5919 (N_5919,N_4068,N_3890);
or U5920 (N_5920,N_3722,N_3607);
nand U5921 (N_5921,N_4259,N_3491);
xor U5922 (N_5922,N_3052,N_3479);
and U5923 (N_5923,N_4048,N_3307);
xnor U5924 (N_5924,N_3751,N_3089);
nor U5925 (N_5925,N_3608,N_3741);
and U5926 (N_5926,N_3854,N_4388);
nor U5927 (N_5927,N_3813,N_4300);
xor U5928 (N_5928,N_3701,N_3041);
xor U5929 (N_5929,N_3747,N_3756);
nor U5930 (N_5930,N_3732,N_4093);
or U5931 (N_5931,N_4295,N_4335);
xnor U5932 (N_5932,N_4042,N_3595);
nor U5933 (N_5933,N_3374,N_3699);
or U5934 (N_5934,N_4094,N_4119);
nand U5935 (N_5935,N_3208,N_4408);
nand U5936 (N_5936,N_4068,N_3910);
nand U5937 (N_5937,N_4024,N_3901);
or U5938 (N_5938,N_3090,N_3334);
or U5939 (N_5939,N_4098,N_3293);
and U5940 (N_5940,N_4064,N_4464);
and U5941 (N_5941,N_3618,N_3977);
xnor U5942 (N_5942,N_3267,N_4146);
nor U5943 (N_5943,N_4143,N_3374);
or U5944 (N_5944,N_3340,N_4217);
nor U5945 (N_5945,N_3664,N_3512);
or U5946 (N_5946,N_3532,N_3873);
nor U5947 (N_5947,N_3841,N_3977);
or U5948 (N_5948,N_4402,N_4228);
xor U5949 (N_5949,N_3952,N_3092);
nor U5950 (N_5950,N_3862,N_3759);
nor U5951 (N_5951,N_3436,N_3281);
nor U5952 (N_5952,N_3628,N_4013);
nand U5953 (N_5953,N_4053,N_4084);
xor U5954 (N_5954,N_3937,N_3957);
xor U5955 (N_5955,N_3968,N_4023);
and U5956 (N_5956,N_3005,N_3920);
nor U5957 (N_5957,N_3150,N_3305);
nand U5958 (N_5958,N_4275,N_3359);
and U5959 (N_5959,N_3265,N_3128);
and U5960 (N_5960,N_3213,N_3176);
nor U5961 (N_5961,N_3901,N_3352);
and U5962 (N_5962,N_4368,N_3167);
xnor U5963 (N_5963,N_3693,N_3169);
nand U5964 (N_5964,N_3761,N_4340);
xor U5965 (N_5965,N_4233,N_4062);
or U5966 (N_5966,N_3398,N_4182);
and U5967 (N_5967,N_3942,N_3999);
or U5968 (N_5968,N_3706,N_3170);
or U5969 (N_5969,N_4266,N_4318);
nand U5970 (N_5970,N_4123,N_4324);
xor U5971 (N_5971,N_3793,N_4054);
nor U5972 (N_5972,N_4185,N_4455);
or U5973 (N_5973,N_4375,N_3039);
or U5974 (N_5974,N_3004,N_3973);
or U5975 (N_5975,N_3943,N_3196);
nand U5976 (N_5976,N_4193,N_3282);
nor U5977 (N_5977,N_3437,N_3832);
xor U5978 (N_5978,N_3457,N_4013);
nor U5979 (N_5979,N_4236,N_3291);
and U5980 (N_5980,N_3381,N_3629);
or U5981 (N_5981,N_3888,N_3212);
nor U5982 (N_5982,N_3806,N_3735);
nor U5983 (N_5983,N_4383,N_4249);
or U5984 (N_5984,N_4214,N_3657);
and U5985 (N_5985,N_3745,N_3513);
and U5986 (N_5986,N_4139,N_3416);
nor U5987 (N_5987,N_4191,N_4135);
nor U5988 (N_5988,N_3048,N_3684);
nor U5989 (N_5989,N_4363,N_3822);
nand U5990 (N_5990,N_3554,N_3930);
nand U5991 (N_5991,N_3200,N_3112);
or U5992 (N_5992,N_3216,N_3111);
nor U5993 (N_5993,N_4125,N_4069);
xnor U5994 (N_5994,N_4069,N_3966);
nor U5995 (N_5995,N_3010,N_4237);
nor U5996 (N_5996,N_3462,N_3887);
nor U5997 (N_5997,N_3434,N_3400);
and U5998 (N_5998,N_4220,N_3159);
nand U5999 (N_5999,N_3429,N_4448);
xor U6000 (N_6000,N_5198,N_4887);
nand U6001 (N_6001,N_5270,N_5734);
and U6002 (N_6002,N_5737,N_5772);
xor U6003 (N_6003,N_5941,N_5799);
nor U6004 (N_6004,N_4706,N_5306);
nand U6005 (N_6005,N_5447,N_4515);
or U6006 (N_6006,N_5070,N_5411);
nor U6007 (N_6007,N_4611,N_4879);
xnor U6008 (N_6008,N_4597,N_5190);
nand U6009 (N_6009,N_5197,N_5653);
and U6010 (N_6010,N_5573,N_5612);
and U6011 (N_6011,N_4541,N_4538);
nand U6012 (N_6012,N_5714,N_4516);
and U6013 (N_6013,N_5843,N_5425);
or U6014 (N_6014,N_5648,N_5549);
or U6015 (N_6015,N_5251,N_5485);
or U6016 (N_6016,N_5615,N_5798);
nand U6017 (N_6017,N_5422,N_5309);
nand U6018 (N_6018,N_5862,N_4874);
nor U6019 (N_6019,N_5252,N_5462);
nor U6020 (N_6020,N_5598,N_5167);
and U6021 (N_6021,N_5933,N_5357);
nor U6022 (N_6022,N_5189,N_5666);
and U6023 (N_6023,N_4907,N_5906);
nand U6024 (N_6024,N_4758,N_4625);
or U6025 (N_6025,N_5311,N_5542);
or U6026 (N_6026,N_4579,N_4634);
or U6027 (N_6027,N_5592,N_5876);
or U6028 (N_6028,N_5032,N_5302);
or U6029 (N_6029,N_5443,N_5509);
nand U6030 (N_6030,N_5572,N_4821);
and U6031 (N_6031,N_5345,N_5238);
nor U6032 (N_6032,N_5579,N_5661);
xor U6033 (N_6033,N_4975,N_5668);
or U6034 (N_6034,N_5724,N_4995);
xor U6035 (N_6035,N_4877,N_4735);
nor U6036 (N_6036,N_5313,N_4923);
xnor U6037 (N_6037,N_5092,N_5670);
and U6038 (N_6038,N_4782,N_5466);
xnor U6039 (N_6039,N_5013,N_5107);
and U6040 (N_6040,N_5526,N_5452);
or U6041 (N_6041,N_5828,N_5684);
nor U6042 (N_6042,N_4826,N_5488);
nor U6043 (N_6043,N_5529,N_4937);
nand U6044 (N_6044,N_5335,N_5209);
nand U6045 (N_6045,N_5300,N_5434);
and U6046 (N_6046,N_5704,N_5791);
nand U6047 (N_6047,N_5649,N_5676);
nand U6048 (N_6048,N_5176,N_5701);
xor U6049 (N_6049,N_5654,N_4551);
xnor U6050 (N_6050,N_4891,N_4674);
or U6051 (N_6051,N_4765,N_5894);
nor U6052 (N_6052,N_5548,N_5562);
xnor U6053 (N_6053,N_5363,N_5959);
and U6054 (N_6054,N_5312,N_5587);
xnor U6055 (N_6055,N_4615,N_5545);
and U6056 (N_6056,N_4702,N_5338);
and U6057 (N_6057,N_5492,N_4829);
or U6058 (N_6058,N_5680,N_4637);
and U6059 (N_6059,N_4521,N_5420);
xnor U6060 (N_6060,N_4948,N_4562);
and U6061 (N_6061,N_4980,N_5928);
or U6062 (N_6062,N_5128,N_5203);
nor U6063 (N_6063,N_5387,N_4575);
nor U6064 (N_6064,N_5867,N_4942);
nand U6065 (N_6065,N_5984,N_4746);
nor U6066 (N_6066,N_5178,N_5632);
nor U6067 (N_6067,N_5046,N_5374);
nand U6068 (N_6068,N_5228,N_5860);
nand U6069 (N_6069,N_4685,N_5308);
nor U6070 (N_6070,N_5504,N_4853);
nand U6071 (N_6071,N_5564,N_5097);
nand U6072 (N_6072,N_5813,N_5002);
and U6073 (N_6073,N_4664,N_5410);
xnor U6074 (N_6074,N_5179,N_5428);
nor U6075 (N_6075,N_4622,N_4857);
and U6076 (N_6076,N_4508,N_5890);
nor U6077 (N_6077,N_5267,N_5191);
xnor U6078 (N_6078,N_5929,N_5534);
and U6079 (N_6079,N_5405,N_5379);
nor U6080 (N_6080,N_5872,N_4546);
nand U6081 (N_6081,N_5682,N_4741);
or U6082 (N_6082,N_4987,N_5431);
nor U6083 (N_6083,N_5138,N_5570);
nand U6084 (N_6084,N_5738,N_5815);
nand U6085 (N_6085,N_5976,N_5433);
xor U6086 (N_6086,N_5142,N_4695);
nor U6087 (N_6087,N_5038,N_4881);
nor U6088 (N_6088,N_4900,N_5050);
nand U6089 (N_6089,N_4639,N_5625);
and U6090 (N_6090,N_5842,N_5963);
xor U6091 (N_6091,N_5494,N_5557);
nand U6092 (N_6092,N_5574,N_4592);
nand U6093 (N_6093,N_4527,N_4965);
xnor U6094 (N_6094,N_5322,N_5160);
nor U6095 (N_6095,N_4960,N_4729);
xor U6096 (N_6096,N_4828,N_5200);
xnor U6097 (N_6097,N_4982,N_4563);
xnor U6098 (N_6098,N_5973,N_4819);
nand U6099 (N_6099,N_5459,N_5827);
nor U6100 (N_6100,N_4889,N_5435);
and U6101 (N_6101,N_4860,N_5911);
or U6102 (N_6102,N_5851,N_4607);
and U6103 (N_6103,N_5997,N_5939);
or U6104 (N_6104,N_4773,N_4967);
or U6105 (N_6105,N_4809,N_5717);
nor U6106 (N_6106,N_5151,N_5691);
and U6107 (N_6107,N_4750,N_4623);
and U6108 (N_6108,N_5458,N_5773);
nor U6109 (N_6109,N_5848,N_4940);
and U6110 (N_6110,N_4897,N_5499);
or U6111 (N_6111,N_5871,N_5878);
and U6112 (N_6112,N_5027,N_5328);
or U6113 (N_6113,N_5817,N_5465);
and U6114 (N_6114,N_5541,N_5419);
nor U6115 (N_6115,N_5109,N_5879);
or U6116 (N_6116,N_4918,N_5366);
or U6117 (N_6117,N_4545,N_4529);
nand U6118 (N_6118,N_4689,N_5825);
and U6119 (N_6119,N_5518,N_5993);
or U6120 (N_6120,N_5750,N_4552);
xor U6121 (N_6121,N_4864,N_5715);
nand U6122 (N_6122,N_4818,N_4973);
nand U6123 (N_6123,N_5693,N_5547);
nand U6124 (N_6124,N_4501,N_5152);
nand U6125 (N_6125,N_5216,N_4598);
or U6126 (N_6126,N_4752,N_5613);
and U6127 (N_6127,N_5165,N_4757);
and U6128 (N_6128,N_4831,N_5482);
nand U6129 (N_6129,N_4703,N_5644);
nor U6130 (N_6130,N_5657,N_5507);
nor U6131 (N_6131,N_5173,N_4616);
nor U6132 (N_6132,N_4715,N_5861);
nor U6133 (N_6133,N_5158,N_4600);
nor U6134 (N_6134,N_5175,N_5427);
nor U6135 (N_6135,N_5273,N_5346);
nor U6136 (N_6136,N_5728,N_4657);
and U6137 (N_6137,N_5282,N_4548);
or U6138 (N_6138,N_5789,N_5761);
xor U6139 (N_6139,N_5351,N_5709);
nor U6140 (N_6140,N_5729,N_5414);
nand U6141 (N_6141,N_5040,N_5120);
and U6142 (N_6142,N_4935,N_5600);
nand U6143 (N_6143,N_5093,N_5469);
xnor U6144 (N_6144,N_5826,N_5486);
nand U6145 (N_6145,N_4558,N_4537);
or U6146 (N_6146,N_5088,N_5225);
nand U6147 (N_6147,N_4949,N_5636);
or U6148 (N_6148,N_5025,N_5051);
and U6149 (N_6149,N_5902,N_4908);
and U6150 (N_6150,N_5368,N_4512);
or U6151 (N_6151,N_5586,N_4500);
and U6152 (N_6152,N_5919,N_5697);
nand U6153 (N_6153,N_5855,N_5974);
nand U6154 (N_6154,N_5857,N_4793);
or U6155 (N_6155,N_4614,N_5936);
nand U6156 (N_6156,N_5490,N_5089);
or U6157 (N_6157,N_4720,N_5082);
or U6158 (N_6158,N_5725,N_5117);
xnor U6159 (N_6159,N_4756,N_5161);
and U6160 (N_6160,N_4903,N_5667);
nand U6161 (N_6161,N_5767,N_5819);
and U6162 (N_6162,N_5930,N_5400);
nand U6163 (N_6163,N_5588,N_5449);
or U6164 (N_6164,N_5009,N_4930);
nand U6165 (N_6165,N_4928,N_5525);
or U6166 (N_6166,N_5188,N_5145);
xor U6167 (N_6167,N_5455,N_5629);
and U6168 (N_6168,N_4636,N_4768);
nand U6169 (N_6169,N_4730,N_4963);
nand U6170 (N_6170,N_4784,N_4693);
and U6171 (N_6171,N_5177,N_4862);
or U6172 (N_6172,N_5155,N_4876);
nand U6173 (N_6173,N_5818,N_4882);
nor U6174 (N_6174,N_5192,N_5266);
nand U6175 (N_6175,N_4704,N_5533);
or U6176 (N_6176,N_5365,N_4909);
nor U6177 (N_6177,N_5949,N_5806);
xnor U6178 (N_6178,N_5268,N_4912);
xor U6179 (N_6179,N_5515,N_5426);
nand U6180 (N_6180,N_4854,N_5491);
xor U6181 (N_6181,N_4904,N_4760);
or U6182 (N_6182,N_5836,N_5550);
nand U6183 (N_6183,N_4599,N_4550);
nor U6184 (N_6184,N_4847,N_5000);
xor U6185 (N_6185,N_5640,N_5917);
nor U6186 (N_6186,N_5147,N_5141);
and U6187 (N_6187,N_5164,N_5703);
xor U6188 (N_6188,N_4531,N_5227);
nand U6189 (N_6189,N_5100,N_5982);
or U6190 (N_6190,N_4823,N_5336);
nand U6191 (N_6191,N_5333,N_5927);
nor U6192 (N_6192,N_5344,N_5217);
and U6193 (N_6193,N_4796,N_5679);
or U6194 (N_6194,N_5620,N_4711);
nand U6195 (N_6195,N_5133,N_5501);
and U6196 (N_6196,N_4858,N_5039);
and U6197 (N_6197,N_4941,N_5619);
nand U6198 (N_6198,N_5575,N_4751);
nand U6199 (N_6199,N_5430,N_4986);
nand U6200 (N_6200,N_5972,N_4865);
or U6201 (N_6201,N_5677,N_4662);
nand U6202 (N_6202,N_5403,N_5742);
xnor U6203 (N_6203,N_5539,N_4885);
and U6204 (N_6204,N_5240,N_5054);
and U6205 (N_6205,N_4565,N_4691);
and U6206 (N_6206,N_5638,N_4656);
nor U6207 (N_6207,N_4806,N_5977);
xnor U6208 (N_6208,N_5886,N_5904);
or U6209 (N_6209,N_4671,N_4884);
and U6210 (N_6210,N_5187,N_5370);
or U6211 (N_6211,N_5681,N_5477);
or U6212 (N_6212,N_5066,N_5237);
nor U6213 (N_6213,N_4966,N_4601);
xor U6214 (N_6214,N_5776,N_4766);
nor U6215 (N_6215,N_5135,N_5249);
xnor U6216 (N_6216,N_4856,N_5678);
nand U6217 (N_6217,N_5394,N_4920);
or U6218 (N_6218,N_5912,N_5845);
and U6219 (N_6219,N_5528,N_4839);
nand U6220 (N_6220,N_5956,N_5988);
or U6221 (N_6221,N_4716,N_4540);
nand U6222 (N_6222,N_5323,N_5095);
xnor U6223 (N_6223,N_5075,N_5398);
or U6224 (N_6224,N_5630,N_4898);
nor U6225 (N_6225,N_4996,N_5213);
nand U6226 (N_6226,N_5388,N_4506);
nor U6227 (N_6227,N_5569,N_5891);
or U6228 (N_6228,N_4810,N_4841);
xor U6229 (N_6229,N_4754,N_5204);
nand U6230 (N_6230,N_4635,N_5146);
nand U6231 (N_6231,N_5162,N_5994);
nor U6232 (N_6232,N_5017,N_5086);
or U6233 (N_6233,N_5830,N_5766);
nor U6234 (N_6234,N_4547,N_5108);
nor U6235 (N_6235,N_4787,N_4571);
or U6236 (N_6236,N_5360,N_5865);
and U6237 (N_6237,N_4762,N_5800);
or U6238 (N_6238,N_5256,N_5236);
xor U6239 (N_6239,N_5775,N_4910);
xor U6240 (N_6240,N_5608,N_4713);
nand U6241 (N_6241,N_5012,N_5473);
nor U6242 (N_6242,N_5663,N_5418);
and U6243 (N_6243,N_5016,N_4699);
nand U6244 (N_6244,N_5617,N_5372);
nor U6245 (N_6245,N_4916,N_4872);
xnor U6246 (N_6246,N_5711,N_4728);
nand U6247 (N_6247,N_4732,N_4914);
nand U6248 (N_6248,N_5467,N_5659);
and U6249 (N_6249,N_4804,N_5597);
xnor U6250 (N_6250,N_5429,N_4777);
xnor U6251 (N_6251,N_5856,N_5645);
or U6252 (N_6252,N_5153,N_5081);
and U6253 (N_6253,N_4525,N_4619);
xnor U6254 (N_6254,N_5321,N_5220);
and U6255 (N_6255,N_5790,N_5348);
nand U6256 (N_6256,N_5290,N_4648);
nand U6257 (N_6257,N_5674,N_5055);
or U6258 (N_6258,N_4605,N_4740);
and U6259 (N_6259,N_4725,N_5445);
and U6260 (N_6260,N_5373,N_5812);
or U6261 (N_6261,N_4800,N_5713);
or U6262 (N_6262,N_4582,N_5331);
nand U6263 (N_6263,N_4507,N_5646);
nor U6264 (N_6264,N_5683,N_4526);
nor U6265 (N_6265,N_4924,N_5866);
xnor U6266 (N_6266,N_4712,N_5870);
and U6267 (N_6267,N_4669,N_5740);
or U6268 (N_6268,N_4859,N_5537);
nor U6269 (N_6269,N_5457,N_5087);
nor U6270 (N_6270,N_4985,N_4532);
xor U6271 (N_6271,N_5883,N_5578);
and U6272 (N_6272,N_5234,N_5299);
nand U6273 (N_6273,N_4846,N_5859);
nand U6274 (N_6274,N_4644,N_5609);
nand U6275 (N_6275,N_5544,N_5523);
nor U6276 (N_6276,N_5361,N_5448);
and U6277 (N_6277,N_4667,N_5942);
or U6278 (N_6278,N_4927,N_4799);
or U6279 (N_6279,N_5786,N_5705);
and U6280 (N_6280,N_5397,N_4992);
nand U6281 (N_6281,N_5222,N_5258);
nor U6282 (N_6282,N_5126,N_4604);
and U6283 (N_6283,N_5156,N_5074);
nand U6284 (N_6284,N_4666,N_5257);
or U6285 (N_6285,N_4700,N_4697);
nand U6286 (N_6286,N_5030,N_4951);
nand U6287 (N_6287,N_4845,N_5310);
or U6288 (N_6288,N_4807,N_5495);
and U6289 (N_6289,N_4961,N_5937);
or U6290 (N_6290,N_4707,N_5888);
or U6291 (N_6291,N_5985,N_5487);
nor U6292 (N_6292,N_4922,N_5552);
nand U6293 (N_6293,N_5062,N_4913);
xor U6294 (N_6294,N_4947,N_5957);
or U6295 (N_6295,N_5854,N_5780);
or U6296 (N_6296,N_4931,N_5036);
or U6297 (N_6297,N_4997,N_4663);
and U6298 (N_6298,N_4917,N_5926);
nor U6299 (N_6299,N_5496,N_4549);
or U6300 (N_6300,N_4812,N_4833);
nand U6301 (N_6301,N_5546,N_4629);
nor U6302 (N_6302,N_5049,N_4983);
and U6303 (N_6303,N_5837,N_5987);
nor U6304 (N_6304,N_5034,N_5205);
nor U6305 (N_6305,N_5960,N_5771);
and U6306 (N_6306,N_5444,N_5858);
xor U6307 (N_6307,N_5978,N_4843);
nor U6308 (N_6308,N_5923,N_5530);
or U6309 (N_6309,N_4934,N_5139);
nand U6310 (N_6310,N_4613,N_5456);
and U6311 (N_6311,N_5764,N_5895);
or U6312 (N_6312,N_5924,N_4677);
nor U6313 (N_6313,N_4559,N_4755);
or U6314 (N_6314,N_5053,N_5384);
nor U6315 (N_6315,N_5364,N_5626);
nand U6316 (N_6316,N_5889,N_4640);
nor U6317 (N_6317,N_5900,N_5755);
and U6318 (N_6318,N_5409,N_5011);
nor U6319 (N_6319,N_4813,N_4871);
and U6320 (N_6320,N_5787,N_5820);
nand U6321 (N_6321,N_5353,N_4785);
nor U6322 (N_6322,N_5698,N_4791);
nor U6323 (N_6323,N_5367,N_5702);
and U6324 (N_6324,N_5281,N_5446);
and U6325 (N_6325,N_4668,N_4722);
nand U6326 (N_6326,N_5271,N_5639);
nor U6327 (N_6327,N_5424,N_5127);
or U6328 (N_6328,N_5568,N_4971);
nor U6329 (N_6329,N_4737,N_4676);
and U6330 (N_6330,N_4645,N_5741);
nand U6331 (N_6331,N_5059,N_5932);
and U6332 (N_6332,N_5315,N_4727);
nor U6333 (N_6333,N_4993,N_5159);
or U6334 (N_6334,N_4647,N_5736);
nor U6335 (N_6335,N_5358,N_5134);
or U6336 (N_6336,N_5967,N_5603);
and U6337 (N_6337,N_5324,N_4781);
and U6338 (N_6338,N_5349,N_5968);
or U6339 (N_6339,N_4519,N_5882);
nor U6340 (N_6340,N_4717,N_5849);
or U6341 (N_6341,N_4984,N_5280);
nor U6342 (N_6342,N_4905,N_5833);
nand U6343 (N_6343,N_5915,N_5295);
nor U6344 (N_6344,N_5201,N_5314);
xor U6345 (N_6345,N_5685,N_5814);
xor U6346 (N_6346,N_4701,N_5005);
and U6347 (N_6347,N_5407,N_4771);
xor U6348 (N_6348,N_5850,N_5047);
or U6349 (N_6349,N_5934,N_5792);
nand U6350 (N_6350,N_5058,N_5606);
or U6351 (N_6351,N_5706,N_5964);
or U6352 (N_6352,N_5390,N_4679);
and U6353 (N_6353,N_4588,N_5413);
nand U6354 (N_6354,N_5244,N_5327);
nand U6355 (N_6355,N_4788,N_5747);
and U6356 (N_6356,N_4564,N_4544);
nor U6357 (N_6357,N_5946,N_4632);
xnor U6358 (N_6358,N_5264,N_5686);
or U6359 (N_6359,N_5334,N_5226);
nand U6360 (N_6360,N_4710,N_5503);
xor U6361 (N_6361,N_5010,N_5788);
nor U6362 (N_6362,N_5991,N_4553);
xor U6363 (N_6363,N_4950,N_4590);
xnor U6364 (N_6364,N_5060,N_5130);
and U6365 (N_6365,N_5821,N_5745);
nand U6366 (N_6366,N_5642,N_5149);
nand U6367 (N_6367,N_5292,N_5277);
nand U6368 (N_6368,N_5041,N_5621);
and U6369 (N_6369,N_5535,N_4926);
and U6370 (N_6370,N_4817,N_4684);
xnor U6371 (N_6371,N_4581,N_4836);
or U6372 (N_6372,N_4682,N_5064);
nand U6373 (N_6373,N_4683,N_5901);
nor U6374 (N_6374,N_4567,N_5451);
nor U6375 (N_6375,N_5938,N_5710);
nand U6376 (N_6376,N_5008,N_5248);
or U6377 (N_6377,N_4504,N_5952);
xor U6378 (N_6378,N_5877,N_5382);
xor U6379 (N_6379,N_5031,N_5920);
or U6380 (N_6380,N_5950,N_4936);
xor U6381 (N_6381,N_5359,N_4834);
and U6382 (N_6382,N_4998,N_4816);
nand U6383 (N_6383,N_5514,N_5660);
xnor U6384 (N_6384,N_5898,N_4822);
nand U6385 (N_6385,N_5184,N_5463);
or U6386 (N_6386,N_5563,N_5071);
or U6387 (N_6387,N_5098,N_5880);
xnor U6388 (N_6388,N_5996,N_5947);
nand U6389 (N_6389,N_5576,N_5981);
xnor U6390 (N_6390,N_4628,N_5869);
and U6391 (N_6391,N_5555,N_5084);
xor U6392 (N_6392,N_5406,N_4994);
xor U6393 (N_6393,N_4911,N_5520);
nand U6394 (N_6394,N_4850,N_5633);
or U6395 (N_6395,N_5591,N_5415);
and U6396 (N_6396,N_4851,N_5399);
nor U6397 (N_6397,N_4867,N_5594);
nor U6398 (N_6398,N_5986,N_5412);
or U6399 (N_6399,N_5521,N_5671);
xnor U6400 (N_6400,N_5777,N_4863);
and U6401 (N_6401,N_4795,N_4972);
nor U6402 (N_6402,N_4901,N_4658);
xnor U6403 (N_6403,N_5230,N_4838);
nand U6404 (N_6404,N_5181,N_5905);
xnor U6405 (N_6405,N_4543,N_4554);
nor U6406 (N_6406,N_5832,N_5332);
nand U6407 (N_6407,N_5199,N_4583);
nor U6408 (N_6408,N_5498,N_5692);
or U6409 (N_6409,N_5834,N_5749);
xnor U6410 (N_6410,N_5069,N_4830);
nand U6411 (N_6411,N_5718,N_4568);
nor U6412 (N_6412,N_5132,N_5369);
and U6413 (N_6413,N_5185,N_5675);
nand U6414 (N_6414,N_5122,N_5553);
nor U6415 (N_6415,N_4946,N_4724);
or U6416 (N_6416,N_5512,N_5722);
xor U6417 (N_6417,N_5913,N_4578);
and U6418 (N_6418,N_4630,N_5899);
and U6419 (N_6419,N_5182,N_5532);
xnor U6420 (N_6420,N_5720,N_5940);
nor U6421 (N_6421,N_5739,N_5506);
nand U6422 (N_6422,N_4719,N_5085);
and U6423 (N_6423,N_4759,N_5805);
and U6424 (N_6424,N_5975,N_5762);
nand U6425 (N_6425,N_5206,N_5339);
or U6426 (N_6426,N_5057,N_5948);
or U6427 (N_6427,N_5247,N_4692);
nand U6428 (N_6428,N_5752,N_5885);
nand U6429 (N_6429,N_5091,N_5116);
nor U6430 (N_6430,N_4820,N_4919);
nand U6431 (N_6431,N_4849,N_5171);
and U6432 (N_6432,N_5567,N_5090);
xor U6433 (N_6433,N_5768,N_4533);
xnor U6434 (N_6434,N_5042,N_4938);
nor U6435 (N_6435,N_4591,N_5634);
nor U6436 (N_6436,N_4510,N_5774);
xor U6437 (N_6437,N_5538,N_5440);
xor U6438 (N_6438,N_5536,N_4690);
or U6439 (N_6439,N_5481,N_5078);
nand U6440 (N_6440,N_5916,N_4848);
xnor U6441 (N_6441,N_5371,N_5840);
nand U6442 (N_6442,N_5026,N_5647);
nor U6443 (N_6443,N_5246,N_4962);
xnor U6444 (N_6444,N_5242,N_5195);
and U6445 (N_6445,N_4573,N_5391);
nor U6446 (N_6446,N_5115,N_5753);
nand U6447 (N_6447,N_5483,N_4783);
or U6448 (N_6448,N_5637,N_4959);
xnor U6449 (N_6449,N_5080,N_4844);
nand U6450 (N_6450,N_5381,N_5875);
or U6451 (N_6451,N_4815,N_4535);
nor U6452 (N_6452,N_5272,N_5297);
nand U6453 (N_6453,N_4958,N_5873);
xnor U6454 (N_6454,N_4566,N_4620);
and U6455 (N_6455,N_4873,N_4572);
nand U6456 (N_6456,N_5232,N_5999);
xnor U6457 (N_6457,N_5610,N_4811);
xnor U6458 (N_6458,N_5795,N_5453);
xor U6459 (N_6459,N_4522,N_5112);
or U6460 (N_6460,N_5694,N_5493);
or U6461 (N_6461,N_5961,N_5196);
and U6462 (N_6462,N_4659,N_4921);
nand U6463 (N_6463,N_4779,N_5980);
or U6464 (N_6464,N_5186,N_5293);
or U6465 (N_6465,N_5695,N_5918);
xor U6466 (N_6466,N_5223,N_5325);
nor U6467 (N_6467,N_5992,N_5241);
nand U6468 (N_6468,N_4868,N_4569);
nor U6469 (N_6469,N_4557,N_5669);
nand U6470 (N_6470,N_5438,N_4523);
xnor U6471 (N_6471,N_5807,N_4866);
nor U6472 (N_6472,N_5278,N_5760);
nand U6473 (N_6473,N_4520,N_5914);
xnor U6474 (N_6474,N_5565,N_4837);
nand U6475 (N_6475,N_5001,N_5500);
xnor U6476 (N_6476,N_5835,N_4824);
xor U6477 (N_6477,N_5154,N_4585);
xnor U6478 (N_6478,N_4978,N_5037);
xor U6479 (N_6479,N_5170,N_5073);
nand U6480 (N_6480,N_5377,N_5925);
nor U6481 (N_6481,N_5423,N_5044);
and U6482 (N_6482,N_5782,N_4767);
and U6483 (N_6483,N_4772,N_4803);
or U6484 (N_6484,N_4832,N_5735);
nand U6485 (N_6485,N_5472,N_5470);
nor U6486 (N_6486,N_5708,N_5931);
xnor U6487 (N_6487,N_4952,N_4738);
xnor U6488 (N_6488,N_5589,N_5380);
and U6489 (N_6489,N_5590,N_5831);
and U6490 (N_6490,N_5383,N_5021);
nor U6491 (N_6491,N_5436,N_4840);
or U6492 (N_6492,N_5604,N_4956);
nand U6493 (N_6493,N_4652,N_4915);
and U6494 (N_6494,N_4624,N_5519);
and U6495 (N_6495,N_5104,N_4610);
or U6496 (N_6496,N_5696,N_5551);
xnor U6497 (N_6497,N_5759,N_4749);
or U6498 (N_6498,N_5556,N_4718);
xor U6499 (N_6499,N_5983,N_5262);
and U6500 (N_6500,N_5275,N_5224);
or U6501 (N_6501,N_5125,N_5096);
or U6502 (N_6502,N_4627,N_5700);
nor U6503 (N_6503,N_5285,N_4555);
and U6504 (N_6504,N_5392,N_5793);
nor U6505 (N_6505,N_5131,N_5194);
nand U6506 (N_6506,N_5595,N_4776);
or U6507 (N_6507,N_5770,N_5471);
nand U6508 (N_6508,N_4786,N_5350);
and U6509 (N_6509,N_5072,N_4748);
and U6510 (N_6510,N_4753,N_5953);
nor U6511 (N_6511,N_5816,N_4649);
and U6512 (N_6512,N_5319,N_4888);
and U6513 (N_6513,N_4842,N_5721);
nand U6514 (N_6514,N_5943,N_4778);
and U6515 (N_6515,N_5829,N_5144);
and U6516 (N_6516,N_5099,N_5137);
nand U6517 (N_6517,N_5602,N_5022);
nand U6518 (N_6518,N_4855,N_5307);
nand U6519 (N_6519,N_4665,N_4709);
xnor U6520 (N_6520,N_4705,N_4686);
xor U6521 (N_6521,N_5094,N_5454);
or U6522 (N_6522,N_5076,N_5015);
nand U6523 (N_6523,N_5652,N_5110);
nand U6524 (N_6524,N_5219,N_5884);
nand U6525 (N_6525,N_5970,N_5824);
nand U6526 (N_6526,N_5375,N_5847);
nand U6527 (N_6527,N_5690,N_4954);
or U6528 (N_6528,N_5045,N_4835);
or U6529 (N_6529,N_4883,N_5396);
nor U6530 (N_6530,N_5113,N_5111);
nor U6531 (N_6531,N_5221,N_5067);
and U6532 (N_6532,N_5823,N_5174);
nand U6533 (N_6533,N_4745,N_5317);
or U6534 (N_6534,N_4991,N_4694);
or U6535 (N_6535,N_4617,N_4852);
xnor U6536 (N_6536,N_4939,N_5731);
or U6537 (N_6537,N_4618,N_5231);
xnor U6538 (N_6538,N_5580,N_5303);
nand U6539 (N_6539,N_4503,N_4764);
or U6540 (N_6540,N_5352,N_5183);
nor U6541 (N_6541,N_5254,N_5497);
xor U6542 (N_6542,N_5763,N_4633);
and U6543 (N_6543,N_4528,N_4505);
and U6544 (N_6544,N_4641,N_5035);
xor U6545 (N_6545,N_5294,N_4661);
xor U6546 (N_6546,N_4653,N_4736);
nand U6547 (N_6547,N_5643,N_4513);
xnor U6548 (N_6548,N_4688,N_5118);
and U6549 (N_6549,N_5079,N_5260);
or U6550 (N_6550,N_4721,N_5635);
xor U6551 (N_6551,N_4654,N_5468);
and U6552 (N_6552,N_5007,N_5616);
nor U6553 (N_6553,N_5907,N_5356);
xor U6554 (N_6554,N_4586,N_5347);
nor U6555 (N_6555,N_5801,N_5839);
xnor U6556 (N_6556,N_5540,N_5461);
nand U6557 (N_6557,N_4517,N_4989);
and U6558 (N_6558,N_5516,N_5605);
and U6559 (N_6559,N_5979,N_4957);
and U6560 (N_6560,N_5558,N_5607);
xor U6561 (N_6561,N_4769,N_4589);
nand U6562 (N_6562,N_5502,N_4990);
xnor U6563 (N_6563,N_5505,N_4814);
nor U6564 (N_6564,N_5316,N_5475);
nor U6565 (N_6565,N_5784,N_5235);
xnor U6566 (N_6566,N_5618,N_5255);
nand U6567 (N_6567,N_4650,N_4642);
nor U6568 (N_6568,N_4609,N_5148);
nor U6569 (N_6569,N_4638,N_5121);
or U6570 (N_6570,N_5655,N_5326);
nand U6571 (N_6571,N_5781,N_4945);
nor U6572 (N_6572,N_5962,N_5474);
and U6573 (N_6573,N_5802,N_4631);
nand U6574 (N_6574,N_5751,N_5510);
and U6575 (N_6575,N_5601,N_5043);
xnor U6576 (N_6576,N_5385,N_5210);
xnor U6577 (N_6577,N_5892,N_5665);
or U6578 (N_6578,N_5990,N_5376);
and U6579 (N_6579,N_5887,N_4933);
nand U6580 (N_6580,N_5945,N_5921);
or U6581 (N_6581,N_4678,N_5897);
or U6582 (N_6582,N_5593,N_4999);
xor U6583 (N_6583,N_5301,N_5864);
nor U6584 (N_6584,N_5658,N_4536);
and U6585 (N_6585,N_5014,N_5757);
nor U6586 (N_6586,N_5508,N_5157);
and U6587 (N_6587,N_4672,N_5935);
xnor U6588 (N_6588,N_5531,N_5136);
or U6589 (N_6589,N_5688,N_5441);
or U6590 (N_6590,N_5803,N_5672);
nor U6591 (N_6591,N_4825,N_4955);
and U6592 (N_6592,N_5279,N_5386);
nand U6593 (N_6593,N_4511,N_4890);
nand U6594 (N_6594,N_4502,N_5522);
nand U6595 (N_6595,N_4680,N_5291);
nand U6596 (N_6596,N_4708,N_5754);
nand U6597 (N_6597,N_5284,N_5006);
nor U6598 (N_6598,N_4602,N_5239);
xnor U6599 (N_6599,N_5758,N_5863);
nand U6600 (N_6600,N_5298,N_5614);
xor U6601 (N_6601,N_4577,N_4761);
xnor U6602 (N_6602,N_5378,N_4988);
nand U6603 (N_6603,N_5852,N_4790);
nand U6604 (N_6604,N_5583,N_5908);
nor U6605 (N_6605,N_4801,N_5218);
and U6606 (N_6606,N_5476,N_5105);
and U6607 (N_6607,N_5489,N_5163);
xor U6608 (N_6608,N_4892,N_4808);
nand U6609 (N_6609,N_4587,N_5896);
nor U6610 (N_6610,N_5746,N_4518);
or U6611 (N_6611,N_4780,N_5582);
xnor U6612 (N_6612,N_5129,N_5061);
or U6613 (N_6613,N_4802,N_5169);
xnor U6614 (N_6614,N_5903,N_5250);
or U6615 (N_6615,N_5641,N_5796);
and U6616 (N_6616,N_5101,N_4805);
nor U6617 (N_6617,N_5401,N_4576);
nor U6618 (N_6618,N_5362,N_5874);
nand U6619 (N_6619,N_4742,N_5511);
and U6620 (N_6620,N_5207,N_5211);
xor U6621 (N_6621,N_4970,N_5342);
or U6622 (N_6622,N_5804,N_5337);
nand U6623 (N_6623,N_5288,N_5664);
xor U6624 (N_6624,N_5868,N_5662);
or U6625 (N_6625,N_5028,N_5408);
nor U6626 (N_6626,N_5123,N_4539);
or U6627 (N_6627,N_5554,N_5102);
nor U6628 (N_6628,N_4561,N_5286);
nor U6629 (N_6629,N_4580,N_4714);
or U6630 (N_6630,N_5846,N_5719);
nand U6631 (N_6631,N_4925,N_4899);
xor U6632 (N_6632,N_5106,N_5744);
and U6633 (N_6633,N_4670,N_5460);
and U6634 (N_6634,N_4875,N_5727);
nand U6635 (N_6635,N_5150,N_5778);
nand U6636 (N_6636,N_4556,N_5029);
nor U6637 (N_6637,N_4675,N_4655);
xor U6638 (N_6638,N_5743,N_5673);
or U6639 (N_6639,N_4968,N_5969);
nor U6640 (N_6640,N_5881,N_5723);
xor U6641 (N_6641,N_5305,N_5822);
nor U6642 (N_6642,N_4621,N_4608);
xor U6643 (N_6643,N_4895,N_5417);
and U6644 (N_6644,N_4827,N_4880);
nor U6645 (N_6645,N_5432,N_5421);
nor U6646 (N_6646,N_5783,N_4774);
nand U6647 (N_6647,N_5627,N_5048);
nand U6648 (N_6648,N_5951,N_4739);
or U6649 (N_6649,N_5631,N_4595);
and U6650 (N_6650,N_5330,N_5656);
nand U6651 (N_6651,N_4861,N_4596);
or U6652 (N_6652,N_5215,N_5003);
and U6653 (N_6653,N_4534,N_5585);
nand U6654 (N_6654,N_5561,N_4651);
nor U6655 (N_6655,N_5958,N_4953);
nand U6656 (N_6656,N_4570,N_5318);
nand U6657 (N_6657,N_4775,N_5212);
nand U6658 (N_6658,N_5596,N_5622);
xnor U6659 (N_6659,N_5730,N_5966);
nand U6660 (N_6660,N_5922,N_5243);
and U6661 (N_6661,N_4932,N_4681);
and U6662 (N_6662,N_4981,N_5699);
xnor U6663 (N_6663,N_5765,N_5442);
and U6664 (N_6664,N_5056,N_5995);
xnor U6665 (N_6665,N_5114,N_5395);
xor U6666 (N_6666,N_5944,N_5543);
and U6667 (N_6667,N_5954,N_5143);
and U6668 (N_6668,N_5732,N_5393);
and U6669 (N_6669,N_5748,N_5261);
nand U6670 (N_6670,N_5304,N_5560);
xnor U6671 (N_6671,N_5168,N_4646);
xor U6672 (N_6672,N_5794,N_5214);
or U6673 (N_6673,N_5527,N_5265);
or U6674 (N_6674,N_5083,N_5276);
nor U6675 (N_6675,N_5517,N_5726);
nor U6676 (N_6676,N_5584,N_4878);
nand U6677 (N_6677,N_4698,N_4902);
or U6678 (N_6678,N_4886,N_5998);
and U6679 (N_6679,N_5624,N_5844);
and U6680 (N_6680,N_4943,N_5320);
or U6681 (N_6681,N_5052,N_5769);
or U6682 (N_6682,N_5269,N_4944);
nand U6683 (N_6683,N_4542,N_5811);
nand U6684 (N_6684,N_4643,N_5808);
nand U6685 (N_6685,N_5229,N_4964);
or U6686 (N_6686,N_4524,N_4514);
or U6687 (N_6687,N_5004,N_5611);
nand U6688 (N_6688,N_5259,N_5478);
and U6689 (N_6689,N_5809,N_4603);
xor U6690 (N_6690,N_5651,N_5989);
nor U6691 (N_6691,N_5402,N_5566);
nor U6692 (N_6692,N_5416,N_5893);
nand U6693 (N_6693,N_4894,N_4979);
or U6694 (N_6694,N_5599,N_5065);
or U6695 (N_6695,N_5341,N_5733);
xnor U6696 (N_6696,N_5779,N_5797);
or U6697 (N_6697,N_5623,N_5464);
xor U6698 (N_6698,N_4723,N_5329);
nor U6699 (N_6699,N_5202,N_4789);
and U6700 (N_6700,N_5479,N_5581);
or U6701 (N_6701,N_4763,N_4893);
and U6702 (N_6702,N_4734,N_5193);
xor U6703 (N_6703,N_5571,N_4584);
or U6704 (N_6704,N_4744,N_4687);
nor U6705 (N_6705,N_5233,N_4870);
xor U6706 (N_6706,N_4976,N_5389);
xnor U6707 (N_6707,N_5245,N_5343);
nor U6708 (N_6708,N_5140,N_5263);
nand U6709 (N_6709,N_5253,N_5909);
xor U6710 (N_6710,N_4594,N_5971);
xor U6711 (N_6711,N_5450,N_5785);
xor U6712 (N_6712,N_5068,N_5172);
xor U6713 (N_6713,N_4593,N_5077);
nand U6714 (N_6714,N_4726,N_5023);
and U6715 (N_6715,N_5716,N_4794);
nand U6716 (N_6716,N_5289,N_5103);
nand U6717 (N_6717,N_5559,N_5853);
nor U6718 (N_6718,N_5340,N_5484);
and U6719 (N_6719,N_5955,N_4798);
or U6720 (N_6720,N_5712,N_4743);
xor U6721 (N_6721,N_4606,N_5687);
or U6722 (N_6722,N_4696,N_4574);
xnor U6723 (N_6723,N_5480,N_5033);
nand U6724 (N_6724,N_5296,N_4673);
nand U6725 (N_6725,N_5689,N_5180);
xnor U6726 (N_6726,N_5020,N_5650);
or U6727 (N_6727,N_5756,N_4906);
nor U6728 (N_6728,N_5287,N_4869);
or U6729 (N_6729,N_4626,N_4509);
and U6730 (N_6730,N_4974,N_5274);
nand U6731 (N_6731,N_5404,N_5355);
or U6732 (N_6732,N_4896,N_4969);
or U6733 (N_6733,N_5838,N_5354);
or U6734 (N_6734,N_4797,N_5841);
xor U6735 (N_6735,N_5283,N_5018);
or U6736 (N_6736,N_4792,N_4770);
or U6737 (N_6737,N_5124,N_5577);
or U6738 (N_6738,N_4560,N_5810);
nand U6739 (N_6739,N_5513,N_5208);
or U6740 (N_6740,N_5524,N_5439);
or U6741 (N_6741,N_4731,N_5166);
nor U6742 (N_6742,N_4929,N_5965);
nand U6743 (N_6743,N_5707,N_4977);
or U6744 (N_6744,N_4530,N_5437);
nor U6745 (N_6745,N_5019,N_5063);
and U6746 (N_6746,N_4660,N_5910);
nand U6747 (N_6747,N_5119,N_4612);
and U6748 (N_6748,N_4733,N_5628);
nor U6749 (N_6749,N_4747,N_5024);
xor U6750 (N_6750,N_5567,N_4806);
nand U6751 (N_6751,N_5629,N_5493);
xor U6752 (N_6752,N_5055,N_4741);
xnor U6753 (N_6753,N_5006,N_5277);
nand U6754 (N_6754,N_4946,N_4985);
nor U6755 (N_6755,N_5546,N_4513);
and U6756 (N_6756,N_5405,N_5868);
or U6757 (N_6757,N_5120,N_4662);
nand U6758 (N_6758,N_5117,N_5354);
nand U6759 (N_6759,N_4842,N_5514);
nor U6760 (N_6760,N_5807,N_5016);
nor U6761 (N_6761,N_5759,N_4980);
and U6762 (N_6762,N_5981,N_5739);
nand U6763 (N_6763,N_4880,N_4740);
or U6764 (N_6764,N_4832,N_4583);
and U6765 (N_6765,N_5943,N_5381);
or U6766 (N_6766,N_5411,N_4684);
and U6767 (N_6767,N_5552,N_4760);
nand U6768 (N_6768,N_4915,N_5797);
xnor U6769 (N_6769,N_4933,N_4770);
xor U6770 (N_6770,N_5049,N_5120);
xnor U6771 (N_6771,N_5158,N_4724);
nor U6772 (N_6772,N_4995,N_5108);
or U6773 (N_6773,N_5741,N_5506);
xor U6774 (N_6774,N_4629,N_5813);
nor U6775 (N_6775,N_5072,N_4895);
and U6776 (N_6776,N_5972,N_5251);
and U6777 (N_6777,N_4923,N_5086);
xnor U6778 (N_6778,N_5987,N_5826);
and U6779 (N_6779,N_5867,N_5643);
or U6780 (N_6780,N_5220,N_4992);
and U6781 (N_6781,N_5835,N_4740);
nand U6782 (N_6782,N_5380,N_5176);
or U6783 (N_6783,N_5343,N_5185);
and U6784 (N_6784,N_4799,N_5985);
nand U6785 (N_6785,N_5226,N_5408);
and U6786 (N_6786,N_5178,N_5912);
nor U6787 (N_6787,N_5171,N_5334);
nand U6788 (N_6788,N_5031,N_5855);
nand U6789 (N_6789,N_5339,N_4726);
nand U6790 (N_6790,N_5242,N_4744);
nor U6791 (N_6791,N_4860,N_4532);
nor U6792 (N_6792,N_4973,N_4705);
and U6793 (N_6793,N_4997,N_4634);
or U6794 (N_6794,N_5921,N_5116);
or U6795 (N_6795,N_4766,N_5279);
or U6796 (N_6796,N_4855,N_4953);
or U6797 (N_6797,N_4548,N_4870);
or U6798 (N_6798,N_4626,N_4652);
nand U6799 (N_6799,N_5330,N_5565);
or U6800 (N_6800,N_5086,N_5538);
nand U6801 (N_6801,N_5627,N_5223);
xnor U6802 (N_6802,N_4946,N_4941);
nand U6803 (N_6803,N_5407,N_4575);
or U6804 (N_6804,N_4883,N_5286);
xor U6805 (N_6805,N_5777,N_5112);
and U6806 (N_6806,N_5007,N_5458);
nor U6807 (N_6807,N_5828,N_5075);
xor U6808 (N_6808,N_5491,N_5217);
nor U6809 (N_6809,N_5866,N_5939);
xnor U6810 (N_6810,N_5305,N_5412);
and U6811 (N_6811,N_4963,N_4871);
nand U6812 (N_6812,N_5829,N_4813);
nor U6813 (N_6813,N_5713,N_4623);
xnor U6814 (N_6814,N_5129,N_5143);
and U6815 (N_6815,N_5331,N_4577);
nor U6816 (N_6816,N_4526,N_4675);
nand U6817 (N_6817,N_5442,N_5471);
nor U6818 (N_6818,N_5392,N_5076);
or U6819 (N_6819,N_4548,N_5402);
nor U6820 (N_6820,N_4998,N_5968);
nand U6821 (N_6821,N_4658,N_5421);
and U6822 (N_6822,N_4633,N_5337);
or U6823 (N_6823,N_5506,N_4505);
nand U6824 (N_6824,N_5975,N_5732);
or U6825 (N_6825,N_5833,N_5538);
nand U6826 (N_6826,N_5273,N_5378);
nand U6827 (N_6827,N_4788,N_4898);
or U6828 (N_6828,N_5088,N_5492);
nor U6829 (N_6829,N_5272,N_5426);
nand U6830 (N_6830,N_4854,N_4946);
and U6831 (N_6831,N_4780,N_5474);
nand U6832 (N_6832,N_5887,N_5095);
or U6833 (N_6833,N_5573,N_5218);
and U6834 (N_6834,N_5611,N_5479);
nor U6835 (N_6835,N_5349,N_5519);
xnor U6836 (N_6836,N_4925,N_4525);
nor U6837 (N_6837,N_5167,N_5362);
xor U6838 (N_6838,N_5861,N_5546);
or U6839 (N_6839,N_5829,N_4606);
nor U6840 (N_6840,N_5331,N_5379);
nand U6841 (N_6841,N_4611,N_5395);
or U6842 (N_6842,N_5834,N_4712);
or U6843 (N_6843,N_5484,N_4797);
nand U6844 (N_6844,N_5273,N_4637);
or U6845 (N_6845,N_5832,N_5882);
nand U6846 (N_6846,N_5829,N_5666);
or U6847 (N_6847,N_5799,N_4880);
and U6848 (N_6848,N_4915,N_5155);
nor U6849 (N_6849,N_5964,N_5306);
nand U6850 (N_6850,N_5582,N_4978);
nor U6851 (N_6851,N_4678,N_4751);
nor U6852 (N_6852,N_4547,N_5328);
nor U6853 (N_6853,N_5289,N_5756);
xnor U6854 (N_6854,N_4634,N_5023);
xor U6855 (N_6855,N_5599,N_5388);
xnor U6856 (N_6856,N_5970,N_4743);
nand U6857 (N_6857,N_5602,N_5931);
or U6858 (N_6858,N_5624,N_4582);
nor U6859 (N_6859,N_4703,N_5836);
xor U6860 (N_6860,N_5527,N_5308);
or U6861 (N_6861,N_5922,N_4903);
nand U6862 (N_6862,N_5142,N_4662);
nand U6863 (N_6863,N_5529,N_5169);
xor U6864 (N_6864,N_5202,N_5628);
nand U6865 (N_6865,N_5780,N_5601);
nand U6866 (N_6866,N_4699,N_4646);
and U6867 (N_6867,N_4584,N_4907);
or U6868 (N_6868,N_5186,N_4859);
nand U6869 (N_6869,N_4821,N_4982);
nand U6870 (N_6870,N_4527,N_5733);
nand U6871 (N_6871,N_5479,N_4666);
nand U6872 (N_6872,N_5244,N_5624);
or U6873 (N_6873,N_5697,N_5799);
or U6874 (N_6874,N_5408,N_5749);
and U6875 (N_6875,N_4894,N_5554);
xor U6876 (N_6876,N_4909,N_5204);
xor U6877 (N_6877,N_5197,N_5030);
and U6878 (N_6878,N_4991,N_4739);
nor U6879 (N_6879,N_5039,N_5921);
or U6880 (N_6880,N_5298,N_5346);
or U6881 (N_6881,N_5275,N_5406);
or U6882 (N_6882,N_5367,N_4577);
or U6883 (N_6883,N_5258,N_5185);
and U6884 (N_6884,N_4935,N_5217);
and U6885 (N_6885,N_4583,N_5165);
nand U6886 (N_6886,N_5314,N_5867);
nand U6887 (N_6887,N_5199,N_5444);
or U6888 (N_6888,N_5704,N_4563);
nand U6889 (N_6889,N_4625,N_5151);
nor U6890 (N_6890,N_5158,N_4835);
and U6891 (N_6891,N_5911,N_5891);
xnor U6892 (N_6892,N_4511,N_5950);
nor U6893 (N_6893,N_4851,N_5846);
and U6894 (N_6894,N_5393,N_5985);
or U6895 (N_6895,N_4834,N_5757);
xor U6896 (N_6896,N_4567,N_5954);
or U6897 (N_6897,N_5580,N_5115);
nand U6898 (N_6898,N_5477,N_5708);
xor U6899 (N_6899,N_4548,N_5715);
xor U6900 (N_6900,N_4926,N_5312);
or U6901 (N_6901,N_5268,N_5616);
or U6902 (N_6902,N_5374,N_5461);
nand U6903 (N_6903,N_4830,N_5238);
nor U6904 (N_6904,N_5404,N_5933);
nand U6905 (N_6905,N_4893,N_4757);
or U6906 (N_6906,N_5022,N_4743);
nor U6907 (N_6907,N_4766,N_5710);
nand U6908 (N_6908,N_4759,N_5227);
nor U6909 (N_6909,N_4681,N_4878);
nor U6910 (N_6910,N_5302,N_4996);
nand U6911 (N_6911,N_5190,N_5653);
nand U6912 (N_6912,N_5242,N_5307);
nor U6913 (N_6913,N_5220,N_4545);
or U6914 (N_6914,N_4847,N_5962);
or U6915 (N_6915,N_5465,N_5307);
or U6916 (N_6916,N_4599,N_5597);
nor U6917 (N_6917,N_5191,N_5240);
or U6918 (N_6918,N_5227,N_4696);
nand U6919 (N_6919,N_5950,N_4699);
xnor U6920 (N_6920,N_5821,N_5911);
or U6921 (N_6921,N_5855,N_5706);
nand U6922 (N_6922,N_4986,N_5239);
xnor U6923 (N_6923,N_5184,N_5640);
nor U6924 (N_6924,N_5140,N_5572);
nor U6925 (N_6925,N_5708,N_5048);
nor U6926 (N_6926,N_5884,N_5570);
xor U6927 (N_6927,N_5057,N_5195);
nor U6928 (N_6928,N_4871,N_5383);
xor U6929 (N_6929,N_5594,N_4523);
and U6930 (N_6930,N_5448,N_4882);
nand U6931 (N_6931,N_5516,N_5991);
nor U6932 (N_6932,N_5190,N_4828);
nor U6933 (N_6933,N_5814,N_5908);
xor U6934 (N_6934,N_5755,N_5228);
and U6935 (N_6935,N_4773,N_5966);
nand U6936 (N_6936,N_5693,N_4731);
and U6937 (N_6937,N_5104,N_5312);
nand U6938 (N_6938,N_4543,N_5234);
nor U6939 (N_6939,N_4627,N_5946);
and U6940 (N_6940,N_5560,N_5635);
nand U6941 (N_6941,N_4872,N_5670);
xnor U6942 (N_6942,N_5693,N_5422);
xor U6943 (N_6943,N_5550,N_5651);
nand U6944 (N_6944,N_4760,N_4859);
or U6945 (N_6945,N_5932,N_5861);
and U6946 (N_6946,N_4972,N_5638);
nor U6947 (N_6947,N_5415,N_4547);
or U6948 (N_6948,N_4571,N_4964);
or U6949 (N_6949,N_5914,N_5605);
nor U6950 (N_6950,N_5107,N_5229);
nand U6951 (N_6951,N_5739,N_4919);
nand U6952 (N_6952,N_5269,N_5586);
nor U6953 (N_6953,N_4929,N_5154);
xnor U6954 (N_6954,N_5591,N_4868);
xor U6955 (N_6955,N_5153,N_5669);
nand U6956 (N_6956,N_5885,N_5874);
and U6957 (N_6957,N_5833,N_5906);
xor U6958 (N_6958,N_4561,N_5133);
and U6959 (N_6959,N_5300,N_5628);
or U6960 (N_6960,N_5532,N_5225);
xor U6961 (N_6961,N_4834,N_5575);
and U6962 (N_6962,N_5675,N_4741);
nand U6963 (N_6963,N_5735,N_5663);
xnor U6964 (N_6964,N_5335,N_5398);
and U6965 (N_6965,N_5472,N_5005);
or U6966 (N_6966,N_5014,N_4541);
xor U6967 (N_6967,N_5832,N_5149);
xnor U6968 (N_6968,N_4729,N_4653);
nand U6969 (N_6969,N_4753,N_5154);
and U6970 (N_6970,N_5670,N_5957);
and U6971 (N_6971,N_5823,N_5034);
nand U6972 (N_6972,N_5836,N_4610);
xnor U6973 (N_6973,N_5531,N_5325);
nand U6974 (N_6974,N_5745,N_4568);
and U6975 (N_6975,N_5730,N_4758);
nand U6976 (N_6976,N_5197,N_5363);
nand U6977 (N_6977,N_5776,N_5742);
nand U6978 (N_6978,N_5412,N_5967);
and U6979 (N_6979,N_4977,N_5945);
and U6980 (N_6980,N_4636,N_4917);
and U6981 (N_6981,N_5322,N_5966);
xnor U6982 (N_6982,N_4653,N_5975);
xnor U6983 (N_6983,N_4687,N_4940);
xnor U6984 (N_6984,N_5713,N_4828);
nor U6985 (N_6985,N_5587,N_5209);
nor U6986 (N_6986,N_4727,N_5414);
nand U6987 (N_6987,N_5114,N_4875);
and U6988 (N_6988,N_5618,N_4681);
nor U6989 (N_6989,N_4600,N_4725);
or U6990 (N_6990,N_4664,N_4593);
nor U6991 (N_6991,N_4970,N_4917);
nand U6992 (N_6992,N_5532,N_5608);
or U6993 (N_6993,N_5674,N_4861);
or U6994 (N_6994,N_5692,N_5390);
and U6995 (N_6995,N_5343,N_4643);
nor U6996 (N_6996,N_5248,N_5240);
or U6997 (N_6997,N_5427,N_5115);
xnor U6998 (N_6998,N_5416,N_4615);
nor U6999 (N_6999,N_4641,N_5399);
xnor U7000 (N_7000,N_4606,N_5656);
xnor U7001 (N_7001,N_5901,N_4866);
xor U7002 (N_7002,N_5158,N_5570);
nand U7003 (N_7003,N_5363,N_5819);
and U7004 (N_7004,N_5284,N_5433);
xnor U7005 (N_7005,N_5500,N_5536);
nand U7006 (N_7006,N_5997,N_5946);
nand U7007 (N_7007,N_4863,N_4550);
or U7008 (N_7008,N_5140,N_4757);
nor U7009 (N_7009,N_4902,N_5366);
nor U7010 (N_7010,N_5995,N_4688);
nor U7011 (N_7011,N_5384,N_4981);
or U7012 (N_7012,N_4956,N_5500);
nand U7013 (N_7013,N_4697,N_5088);
or U7014 (N_7014,N_4627,N_4714);
or U7015 (N_7015,N_4907,N_5051);
nand U7016 (N_7016,N_5896,N_4927);
and U7017 (N_7017,N_5567,N_5695);
xnor U7018 (N_7018,N_5757,N_5151);
nand U7019 (N_7019,N_4820,N_4642);
or U7020 (N_7020,N_5397,N_5252);
xnor U7021 (N_7021,N_5926,N_5711);
xor U7022 (N_7022,N_4860,N_5212);
or U7023 (N_7023,N_5369,N_4887);
xnor U7024 (N_7024,N_4561,N_5326);
or U7025 (N_7025,N_5664,N_5481);
or U7026 (N_7026,N_5301,N_4666);
and U7027 (N_7027,N_5589,N_5465);
and U7028 (N_7028,N_5778,N_4928);
and U7029 (N_7029,N_5730,N_5773);
and U7030 (N_7030,N_5874,N_5570);
nor U7031 (N_7031,N_5597,N_4537);
or U7032 (N_7032,N_5874,N_5359);
xnor U7033 (N_7033,N_4946,N_5902);
and U7034 (N_7034,N_5302,N_4678);
or U7035 (N_7035,N_5418,N_5445);
and U7036 (N_7036,N_4717,N_4860);
nor U7037 (N_7037,N_4526,N_5883);
nor U7038 (N_7038,N_4538,N_5327);
or U7039 (N_7039,N_5403,N_4623);
xnor U7040 (N_7040,N_5044,N_5325);
or U7041 (N_7041,N_4605,N_4534);
and U7042 (N_7042,N_5262,N_4694);
or U7043 (N_7043,N_4582,N_5822);
xnor U7044 (N_7044,N_4556,N_5026);
nor U7045 (N_7045,N_5737,N_5184);
xnor U7046 (N_7046,N_4660,N_5887);
nor U7047 (N_7047,N_4665,N_5143);
or U7048 (N_7048,N_5515,N_5028);
and U7049 (N_7049,N_5620,N_5266);
nand U7050 (N_7050,N_4610,N_5509);
xnor U7051 (N_7051,N_4926,N_5019);
xor U7052 (N_7052,N_4885,N_4896);
xor U7053 (N_7053,N_5819,N_4655);
xnor U7054 (N_7054,N_4905,N_5963);
and U7055 (N_7055,N_4736,N_5959);
nor U7056 (N_7056,N_5087,N_5514);
nor U7057 (N_7057,N_5947,N_5418);
or U7058 (N_7058,N_5770,N_4805);
xnor U7059 (N_7059,N_4642,N_5621);
xnor U7060 (N_7060,N_5312,N_5660);
or U7061 (N_7061,N_4546,N_5532);
and U7062 (N_7062,N_5234,N_5288);
xor U7063 (N_7063,N_4720,N_5219);
nor U7064 (N_7064,N_5749,N_4904);
xnor U7065 (N_7065,N_5635,N_5521);
nand U7066 (N_7066,N_4512,N_4698);
or U7067 (N_7067,N_5757,N_4955);
nand U7068 (N_7068,N_5171,N_5089);
nand U7069 (N_7069,N_5361,N_5238);
nand U7070 (N_7070,N_5896,N_5985);
or U7071 (N_7071,N_5101,N_4988);
or U7072 (N_7072,N_5783,N_5689);
nand U7073 (N_7073,N_4535,N_5908);
xnor U7074 (N_7074,N_5042,N_5560);
xor U7075 (N_7075,N_4996,N_4795);
or U7076 (N_7076,N_5029,N_5430);
xnor U7077 (N_7077,N_5871,N_5965);
nor U7078 (N_7078,N_5527,N_5103);
and U7079 (N_7079,N_4592,N_4630);
nand U7080 (N_7080,N_5315,N_4813);
nor U7081 (N_7081,N_5826,N_5224);
nor U7082 (N_7082,N_4603,N_4566);
xor U7083 (N_7083,N_5970,N_5835);
and U7084 (N_7084,N_4768,N_5081);
and U7085 (N_7085,N_5867,N_5082);
and U7086 (N_7086,N_5332,N_5768);
and U7087 (N_7087,N_5964,N_5528);
and U7088 (N_7088,N_4924,N_5993);
nor U7089 (N_7089,N_5571,N_5589);
xor U7090 (N_7090,N_5959,N_5922);
nand U7091 (N_7091,N_4542,N_5505);
nand U7092 (N_7092,N_4555,N_5709);
nor U7093 (N_7093,N_5578,N_4701);
or U7094 (N_7094,N_5025,N_5826);
and U7095 (N_7095,N_5481,N_5983);
or U7096 (N_7096,N_5411,N_4858);
and U7097 (N_7097,N_4941,N_5316);
xnor U7098 (N_7098,N_4978,N_5616);
nor U7099 (N_7099,N_5246,N_4779);
or U7100 (N_7100,N_4800,N_5390);
nor U7101 (N_7101,N_4727,N_5159);
xnor U7102 (N_7102,N_5168,N_4658);
nor U7103 (N_7103,N_5251,N_5899);
nand U7104 (N_7104,N_4968,N_4924);
nand U7105 (N_7105,N_4525,N_5939);
and U7106 (N_7106,N_5795,N_5402);
xor U7107 (N_7107,N_5593,N_5476);
and U7108 (N_7108,N_4576,N_4514);
nor U7109 (N_7109,N_5001,N_5343);
and U7110 (N_7110,N_5458,N_4830);
and U7111 (N_7111,N_5625,N_5813);
or U7112 (N_7112,N_5979,N_5786);
nor U7113 (N_7113,N_4938,N_5584);
xor U7114 (N_7114,N_4935,N_4607);
nor U7115 (N_7115,N_5642,N_5605);
and U7116 (N_7116,N_5127,N_5988);
xor U7117 (N_7117,N_5509,N_5307);
nor U7118 (N_7118,N_5962,N_5612);
and U7119 (N_7119,N_5120,N_5159);
or U7120 (N_7120,N_5114,N_5605);
or U7121 (N_7121,N_5729,N_4519);
xnor U7122 (N_7122,N_5421,N_5114);
xnor U7123 (N_7123,N_4998,N_4986);
xor U7124 (N_7124,N_5485,N_4936);
and U7125 (N_7125,N_4715,N_4838);
nand U7126 (N_7126,N_4919,N_4534);
and U7127 (N_7127,N_5653,N_4803);
nand U7128 (N_7128,N_4777,N_5304);
xnor U7129 (N_7129,N_5465,N_5073);
nand U7130 (N_7130,N_5155,N_5883);
nand U7131 (N_7131,N_5329,N_5524);
and U7132 (N_7132,N_5298,N_5420);
nand U7133 (N_7133,N_5535,N_5272);
xor U7134 (N_7134,N_5230,N_5533);
and U7135 (N_7135,N_5240,N_5257);
or U7136 (N_7136,N_4724,N_5991);
or U7137 (N_7137,N_5170,N_5651);
and U7138 (N_7138,N_5651,N_5646);
or U7139 (N_7139,N_5936,N_5158);
xor U7140 (N_7140,N_4564,N_5513);
nand U7141 (N_7141,N_4942,N_5095);
or U7142 (N_7142,N_5058,N_5154);
nand U7143 (N_7143,N_5184,N_4840);
xor U7144 (N_7144,N_5387,N_5465);
and U7145 (N_7145,N_5571,N_5568);
xor U7146 (N_7146,N_5467,N_5655);
and U7147 (N_7147,N_5200,N_4654);
nor U7148 (N_7148,N_4953,N_5594);
and U7149 (N_7149,N_4683,N_5943);
or U7150 (N_7150,N_5224,N_5088);
and U7151 (N_7151,N_4852,N_5569);
xor U7152 (N_7152,N_5454,N_5042);
nand U7153 (N_7153,N_4931,N_4991);
nand U7154 (N_7154,N_5507,N_4971);
xor U7155 (N_7155,N_4729,N_5406);
nor U7156 (N_7156,N_5187,N_4547);
xnor U7157 (N_7157,N_4838,N_5418);
nor U7158 (N_7158,N_5360,N_5533);
nor U7159 (N_7159,N_5032,N_5875);
or U7160 (N_7160,N_5591,N_4790);
nand U7161 (N_7161,N_4707,N_4713);
nor U7162 (N_7162,N_5702,N_4801);
nand U7163 (N_7163,N_5029,N_4667);
xnor U7164 (N_7164,N_5046,N_5213);
xor U7165 (N_7165,N_4618,N_5591);
xnor U7166 (N_7166,N_5807,N_5099);
nand U7167 (N_7167,N_5197,N_5324);
nor U7168 (N_7168,N_4606,N_5324);
and U7169 (N_7169,N_5547,N_5097);
nor U7170 (N_7170,N_5328,N_5777);
and U7171 (N_7171,N_4594,N_5514);
nand U7172 (N_7172,N_5999,N_4626);
xor U7173 (N_7173,N_5554,N_5505);
nor U7174 (N_7174,N_5070,N_5506);
nor U7175 (N_7175,N_4606,N_5832);
nor U7176 (N_7176,N_4621,N_4546);
and U7177 (N_7177,N_5964,N_5609);
and U7178 (N_7178,N_5029,N_5974);
xor U7179 (N_7179,N_4777,N_4663);
nor U7180 (N_7180,N_4809,N_5181);
and U7181 (N_7181,N_4580,N_5252);
and U7182 (N_7182,N_5975,N_5331);
xnor U7183 (N_7183,N_5293,N_4524);
xnor U7184 (N_7184,N_4971,N_5609);
nor U7185 (N_7185,N_5715,N_4999);
or U7186 (N_7186,N_4885,N_4624);
and U7187 (N_7187,N_5780,N_5093);
or U7188 (N_7188,N_5435,N_5560);
and U7189 (N_7189,N_5180,N_5938);
xnor U7190 (N_7190,N_5212,N_4965);
nand U7191 (N_7191,N_4808,N_4773);
nor U7192 (N_7192,N_4674,N_4974);
nor U7193 (N_7193,N_4794,N_5398);
and U7194 (N_7194,N_5320,N_5922);
and U7195 (N_7195,N_5086,N_5280);
xor U7196 (N_7196,N_4520,N_5113);
nor U7197 (N_7197,N_5249,N_4520);
or U7198 (N_7198,N_5764,N_5917);
xor U7199 (N_7199,N_5932,N_5512);
xor U7200 (N_7200,N_4818,N_4605);
and U7201 (N_7201,N_5613,N_4792);
nor U7202 (N_7202,N_4944,N_5850);
nor U7203 (N_7203,N_5287,N_4924);
xnor U7204 (N_7204,N_5636,N_5663);
nand U7205 (N_7205,N_5758,N_5587);
nor U7206 (N_7206,N_5690,N_4646);
nand U7207 (N_7207,N_5804,N_4886);
xor U7208 (N_7208,N_4794,N_5792);
xor U7209 (N_7209,N_5752,N_5032);
xnor U7210 (N_7210,N_4505,N_5348);
nand U7211 (N_7211,N_4795,N_4612);
nor U7212 (N_7212,N_4678,N_5143);
nand U7213 (N_7213,N_4941,N_5197);
or U7214 (N_7214,N_5566,N_5848);
nor U7215 (N_7215,N_5913,N_5525);
xnor U7216 (N_7216,N_4966,N_5407);
or U7217 (N_7217,N_5639,N_4806);
xnor U7218 (N_7218,N_5570,N_5392);
and U7219 (N_7219,N_5932,N_5829);
and U7220 (N_7220,N_4656,N_4935);
and U7221 (N_7221,N_5460,N_5684);
nand U7222 (N_7222,N_5785,N_4736);
nor U7223 (N_7223,N_5380,N_4965);
xnor U7224 (N_7224,N_5529,N_4539);
nor U7225 (N_7225,N_5538,N_4956);
nand U7226 (N_7226,N_5521,N_5395);
or U7227 (N_7227,N_5399,N_5977);
or U7228 (N_7228,N_5017,N_5989);
nor U7229 (N_7229,N_5646,N_4657);
nand U7230 (N_7230,N_4954,N_5986);
xnor U7231 (N_7231,N_5802,N_5418);
xor U7232 (N_7232,N_4980,N_5775);
and U7233 (N_7233,N_5671,N_5900);
and U7234 (N_7234,N_5981,N_5946);
and U7235 (N_7235,N_5311,N_5651);
xnor U7236 (N_7236,N_5273,N_5646);
or U7237 (N_7237,N_4707,N_5252);
and U7238 (N_7238,N_5961,N_5997);
nand U7239 (N_7239,N_5242,N_4741);
and U7240 (N_7240,N_5530,N_5421);
xnor U7241 (N_7241,N_5526,N_5209);
xor U7242 (N_7242,N_5827,N_5091);
xnor U7243 (N_7243,N_4898,N_4965);
nand U7244 (N_7244,N_5137,N_4809);
nor U7245 (N_7245,N_5011,N_5154);
nand U7246 (N_7246,N_5098,N_5741);
nand U7247 (N_7247,N_5887,N_5723);
nand U7248 (N_7248,N_4722,N_5044);
or U7249 (N_7249,N_5949,N_4997);
nor U7250 (N_7250,N_4777,N_5627);
nor U7251 (N_7251,N_5303,N_5088);
nor U7252 (N_7252,N_5536,N_5800);
xor U7253 (N_7253,N_5177,N_5234);
nand U7254 (N_7254,N_5123,N_4653);
nand U7255 (N_7255,N_5236,N_5808);
nand U7256 (N_7256,N_4786,N_5856);
and U7257 (N_7257,N_4856,N_5129);
and U7258 (N_7258,N_5915,N_5447);
or U7259 (N_7259,N_5289,N_4712);
and U7260 (N_7260,N_5628,N_5145);
and U7261 (N_7261,N_5933,N_5937);
and U7262 (N_7262,N_5734,N_5812);
and U7263 (N_7263,N_5641,N_5542);
nand U7264 (N_7264,N_5871,N_5945);
xor U7265 (N_7265,N_5848,N_4941);
nand U7266 (N_7266,N_4877,N_5556);
xnor U7267 (N_7267,N_5685,N_5549);
and U7268 (N_7268,N_4867,N_4719);
nand U7269 (N_7269,N_5843,N_5848);
and U7270 (N_7270,N_4749,N_5845);
xnor U7271 (N_7271,N_4768,N_5888);
nor U7272 (N_7272,N_5141,N_5854);
nand U7273 (N_7273,N_5740,N_5303);
xnor U7274 (N_7274,N_4996,N_5950);
and U7275 (N_7275,N_5746,N_5505);
and U7276 (N_7276,N_5447,N_5939);
nor U7277 (N_7277,N_5803,N_5038);
xnor U7278 (N_7278,N_4593,N_4851);
xnor U7279 (N_7279,N_5395,N_5636);
nor U7280 (N_7280,N_4945,N_4595);
or U7281 (N_7281,N_5779,N_4613);
and U7282 (N_7282,N_5515,N_5926);
or U7283 (N_7283,N_5499,N_4505);
nand U7284 (N_7284,N_5471,N_5681);
xnor U7285 (N_7285,N_4837,N_4540);
xor U7286 (N_7286,N_5049,N_4816);
nand U7287 (N_7287,N_4666,N_5120);
xnor U7288 (N_7288,N_4781,N_4632);
and U7289 (N_7289,N_5882,N_5403);
or U7290 (N_7290,N_5772,N_5594);
and U7291 (N_7291,N_5109,N_5218);
or U7292 (N_7292,N_5872,N_5885);
and U7293 (N_7293,N_5150,N_4841);
xor U7294 (N_7294,N_5464,N_5068);
nand U7295 (N_7295,N_5570,N_5251);
and U7296 (N_7296,N_5750,N_4891);
or U7297 (N_7297,N_5252,N_5263);
nand U7298 (N_7298,N_5728,N_5655);
nor U7299 (N_7299,N_4671,N_4729);
xnor U7300 (N_7300,N_5087,N_4710);
nor U7301 (N_7301,N_5336,N_4635);
and U7302 (N_7302,N_4672,N_4507);
xor U7303 (N_7303,N_5484,N_5634);
xor U7304 (N_7304,N_5913,N_5868);
nor U7305 (N_7305,N_4604,N_4861);
nand U7306 (N_7306,N_5387,N_5041);
nand U7307 (N_7307,N_4915,N_5286);
xor U7308 (N_7308,N_5889,N_5148);
and U7309 (N_7309,N_5182,N_5786);
or U7310 (N_7310,N_5761,N_5865);
nand U7311 (N_7311,N_4524,N_5251);
nor U7312 (N_7312,N_5518,N_4836);
or U7313 (N_7313,N_5043,N_5274);
nand U7314 (N_7314,N_5285,N_5398);
xor U7315 (N_7315,N_5228,N_4693);
or U7316 (N_7316,N_5415,N_5025);
nand U7317 (N_7317,N_4898,N_5650);
nand U7318 (N_7318,N_5384,N_5376);
xor U7319 (N_7319,N_5348,N_5600);
nand U7320 (N_7320,N_5771,N_4728);
nor U7321 (N_7321,N_5167,N_5048);
and U7322 (N_7322,N_5102,N_4662);
or U7323 (N_7323,N_4624,N_5148);
nand U7324 (N_7324,N_5524,N_4674);
nand U7325 (N_7325,N_5306,N_5149);
xor U7326 (N_7326,N_5951,N_5223);
and U7327 (N_7327,N_5489,N_5209);
nand U7328 (N_7328,N_4543,N_5623);
nand U7329 (N_7329,N_5671,N_5339);
nor U7330 (N_7330,N_5935,N_5583);
nor U7331 (N_7331,N_4577,N_5516);
nand U7332 (N_7332,N_4558,N_5324);
or U7333 (N_7333,N_4938,N_5667);
nand U7334 (N_7334,N_5711,N_4767);
nand U7335 (N_7335,N_4784,N_5182);
nand U7336 (N_7336,N_5078,N_4846);
nor U7337 (N_7337,N_5987,N_5041);
nor U7338 (N_7338,N_4554,N_5680);
and U7339 (N_7339,N_4930,N_5570);
xnor U7340 (N_7340,N_4584,N_5944);
or U7341 (N_7341,N_5829,N_5527);
and U7342 (N_7342,N_5218,N_5552);
nand U7343 (N_7343,N_5963,N_4571);
xnor U7344 (N_7344,N_5658,N_5257);
nand U7345 (N_7345,N_4865,N_4598);
xor U7346 (N_7346,N_4894,N_5131);
xnor U7347 (N_7347,N_5079,N_5147);
or U7348 (N_7348,N_5751,N_5694);
nand U7349 (N_7349,N_5947,N_5841);
or U7350 (N_7350,N_5316,N_5821);
or U7351 (N_7351,N_5759,N_5693);
nand U7352 (N_7352,N_4849,N_5985);
xnor U7353 (N_7353,N_5920,N_4612);
or U7354 (N_7354,N_5400,N_5155);
nor U7355 (N_7355,N_5584,N_5175);
xnor U7356 (N_7356,N_5827,N_4637);
or U7357 (N_7357,N_4873,N_4833);
nand U7358 (N_7358,N_4733,N_5858);
xnor U7359 (N_7359,N_4814,N_4795);
xor U7360 (N_7360,N_5553,N_4873);
xnor U7361 (N_7361,N_5291,N_5670);
xnor U7362 (N_7362,N_5098,N_4551);
nor U7363 (N_7363,N_4637,N_5106);
nand U7364 (N_7364,N_4514,N_5441);
and U7365 (N_7365,N_5990,N_5746);
and U7366 (N_7366,N_5885,N_5951);
nor U7367 (N_7367,N_5217,N_5546);
nand U7368 (N_7368,N_5783,N_5185);
or U7369 (N_7369,N_5236,N_5070);
and U7370 (N_7370,N_5673,N_5330);
nor U7371 (N_7371,N_5071,N_4762);
xor U7372 (N_7372,N_4555,N_4757);
nand U7373 (N_7373,N_5863,N_5233);
or U7374 (N_7374,N_5878,N_5722);
xor U7375 (N_7375,N_5801,N_5022);
and U7376 (N_7376,N_4986,N_5297);
nor U7377 (N_7377,N_5072,N_4912);
and U7378 (N_7378,N_5982,N_5712);
nor U7379 (N_7379,N_5568,N_5413);
nand U7380 (N_7380,N_4646,N_5550);
nor U7381 (N_7381,N_5327,N_5937);
nand U7382 (N_7382,N_4954,N_5890);
xnor U7383 (N_7383,N_4885,N_4716);
and U7384 (N_7384,N_5699,N_5645);
xor U7385 (N_7385,N_5934,N_5860);
nand U7386 (N_7386,N_4514,N_5767);
nand U7387 (N_7387,N_5152,N_5610);
and U7388 (N_7388,N_5449,N_5304);
nand U7389 (N_7389,N_5079,N_5825);
or U7390 (N_7390,N_5665,N_5031);
xnor U7391 (N_7391,N_5086,N_4596);
nor U7392 (N_7392,N_4589,N_5856);
and U7393 (N_7393,N_4717,N_4989);
xnor U7394 (N_7394,N_5927,N_5804);
nor U7395 (N_7395,N_4687,N_5732);
nand U7396 (N_7396,N_5960,N_5494);
and U7397 (N_7397,N_5768,N_5909);
xnor U7398 (N_7398,N_4867,N_4699);
or U7399 (N_7399,N_5717,N_5686);
xnor U7400 (N_7400,N_5188,N_4681);
xor U7401 (N_7401,N_4531,N_5243);
and U7402 (N_7402,N_5841,N_4536);
and U7403 (N_7403,N_4845,N_5531);
and U7404 (N_7404,N_5063,N_5626);
nand U7405 (N_7405,N_5093,N_4885);
or U7406 (N_7406,N_5757,N_4967);
or U7407 (N_7407,N_5378,N_4706);
nand U7408 (N_7408,N_4763,N_4507);
nand U7409 (N_7409,N_5502,N_5927);
and U7410 (N_7410,N_5332,N_5183);
or U7411 (N_7411,N_5321,N_5179);
xor U7412 (N_7412,N_5983,N_5938);
and U7413 (N_7413,N_5201,N_4626);
xnor U7414 (N_7414,N_5043,N_4696);
nand U7415 (N_7415,N_5713,N_5816);
nand U7416 (N_7416,N_5837,N_4944);
or U7417 (N_7417,N_4670,N_5635);
nand U7418 (N_7418,N_5932,N_5979);
or U7419 (N_7419,N_5278,N_4787);
nand U7420 (N_7420,N_5373,N_5732);
xor U7421 (N_7421,N_5891,N_5822);
or U7422 (N_7422,N_5518,N_4741);
xor U7423 (N_7423,N_4629,N_5769);
and U7424 (N_7424,N_4952,N_5921);
or U7425 (N_7425,N_4533,N_4706);
and U7426 (N_7426,N_5364,N_5255);
nor U7427 (N_7427,N_5982,N_4548);
nand U7428 (N_7428,N_4726,N_4518);
nor U7429 (N_7429,N_4696,N_5495);
nand U7430 (N_7430,N_5138,N_5121);
and U7431 (N_7431,N_5300,N_4922);
xnor U7432 (N_7432,N_5515,N_5761);
nor U7433 (N_7433,N_5600,N_5056);
xnor U7434 (N_7434,N_5319,N_5467);
xnor U7435 (N_7435,N_5397,N_5963);
nand U7436 (N_7436,N_5764,N_5855);
xnor U7437 (N_7437,N_4757,N_5006);
nand U7438 (N_7438,N_4985,N_5064);
nand U7439 (N_7439,N_5841,N_5303);
and U7440 (N_7440,N_5111,N_5275);
nand U7441 (N_7441,N_5743,N_5176);
xor U7442 (N_7442,N_5132,N_4981);
nor U7443 (N_7443,N_5691,N_5462);
nand U7444 (N_7444,N_5400,N_5755);
nor U7445 (N_7445,N_4942,N_5931);
nor U7446 (N_7446,N_4883,N_4846);
nand U7447 (N_7447,N_5475,N_5191);
nor U7448 (N_7448,N_5832,N_4621);
or U7449 (N_7449,N_4500,N_4777);
nand U7450 (N_7450,N_5101,N_5780);
or U7451 (N_7451,N_4811,N_5991);
nand U7452 (N_7452,N_5663,N_5256);
nor U7453 (N_7453,N_5978,N_5817);
and U7454 (N_7454,N_5979,N_5435);
nand U7455 (N_7455,N_5520,N_5521);
xnor U7456 (N_7456,N_5179,N_5239);
xor U7457 (N_7457,N_4797,N_5456);
nand U7458 (N_7458,N_5573,N_5060);
nand U7459 (N_7459,N_4974,N_4580);
xnor U7460 (N_7460,N_4920,N_5409);
nand U7461 (N_7461,N_5289,N_5158);
or U7462 (N_7462,N_5839,N_4612);
nand U7463 (N_7463,N_4973,N_5210);
nor U7464 (N_7464,N_4814,N_5404);
nand U7465 (N_7465,N_5683,N_5352);
and U7466 (N_7466,N_5394,N_5666);
nand U7467 (N_7467,N_5657,N_5223);
and U7468 (N_7468,N_5577,N_4684);
and U7469 (N_7469,N_4509,N_5836);
xnor U7470 (N_7470,N_4581,N_4719);
or U7471 (N_7471,N_4656,N_4527);
nand U7472 (N_7472,N_4648,N_5262);
xnor U7473 (N_7473,N_5429,N_5148);
nand U7474 (N_7474,N_5819,N_5471);
and U7475 (N_7475,N_5483,N_4605);
and U7476 (N_7476,N_4865,N_5474);
nand U7477 (N_7477,N_5823,N_5651);
and U7478 (N_7478,N_5748,N_4970);
xor U7479 (N_7479,N_5709,N_4687);
xnor U7480 (N_7480,N_4680,N_4909);
xnor U7481 (N_7481,N_4982,N_4798);
xnor U7482 (N_7482,N_4519,N_5332);
xor U7483 (N_7483,N_4771,N_5043);
and U7484 (N_7484,N_5939,N_4789);
nand U7485 (N_7485,N_4541,N_5947);
and U7486 (N_7486,N_5229,N_5684);
nand U7487 (N_7487,N_5090,N_5710);
or U7488 (N_7488,N_5373,N_4755);
nand U7489 (N_7489,N_5165,N_4542);
nor U7490 (N_7490,N_5135,N_5525);
nand U7491 (N_7491,N_5354,N_4574);
nand U7492 (N_7492,N_4986,N_5050);
and U7493 (N_7493,N_5069,N_4771);
or U7494 (N_7494,N_4643,N_4689);
or U7495 (N_7495,N_5238,N_5862);
or U7496 (N_7496,N_5291,N_5802);
or U7497 (N_7497,N_5160,N_5305);
nand U7498 (N_7498,N_5004,N_4930);
and U7499 (N_7499,N_5965,N_5489);
nor U7500 (N_7500,N_6305,N_6535);
and U7501 (N_7501,N_6204,N_7258);
xor U7502 (N_7502,N_6183,N_7067);
and U7503 (N_7503,N_6439,N_7059);
nand U7504 (N_7504,N_6530,N_6415);
and U7505 (N_7505,N_7307,N_7194);
nor U7506 (N_7506,N_6723,N_6128);
xnor U7507 (N_7507,N_7010,N_6505);
or U7508 (N_7508,N_6539,N_6832);
or U7509 (N_7509,N_7265,N_7152);
xor U7510 (N_7510,N_7309,N_6162);
xnor U7511 (N_7511,N_6501,N_6947);
and U7512 (N_7512,N_7123,N_7174);
or U7513 (N_7513,N_7373,N_7208);
or U7514 (N_7514,N_6679,N_6036);
and U7515 (N_7515,N_6536,N_6447);
or U7516 (N_7516,N_6508,N_7132);
nand U7517 (N_7517,N_6798,N_6796);
xor U7518 (N_7518,N_7320,N_6902);
nand U7519 (N_7519,N_7427,N_6895);
nand U7520 (N_7520,N_6084,N_6690);
and U7521 (N_7521,N_6281,N_6239);
xor U7522 (N_7522,N_6253,N_7481);
or U7523 (N_7523,N_6569,N_6233);
xnor U7524 (N_7524,N_6836,N_6152);
and U7525 (N_7525,N_6790,N_6694);
or U7526 (N_7526,N_7392,N_7256);
or U7527 (N_7527,N_6019,N_6748);
xor U7528 (N_7528,N_6781,N_6333);
xor U7529 (N_7529,N_6026,N_7379);
and U7530 (N_7530,N_7070,N_7149);
xor U7531 (N_7531,N_6698,N_6753);
or U7532 (N_7532,N_7031,N_6481);
xor U7533 (N_7533,N_7122,N_6572);
nand U7534 (N_7534,N_6038,N_7326);
nand U7535 (N_7535,N_7316,N_6802);
nor U7536 (N_7536,N_7173,N_6440);
and U7537 (N_7537,N_6990,N_7482);
and U7538 (N_7538,N_6489,N_6358);
nand U7539 (N_7539,N_6526,N_6755);
and U7540 (N_7540,N_6774,N_7297);
nor U7541 (N_7541,N_6692,N_7022);
xnor U7542 (N_7542,N_6100,N_6403);
or U7543 (N_7543,N_7211,N_7124);
nor U7544 (N_7544,N_7156,N_6289);
xnor U7545 (N_7545,N_6394,N_7428);
and U7546 (N_7546,N_6719,N_6455);
xor U7547 (N_7547,N_7065,N_7319);
and U7548 (N_7548,N_7414,N_6938);
nor U7549 (N_7549,N_6966,N_6971);
nor U7550 (N_7550,N_7252,N_7417);
or U7551 (N_7551,N_6376,N_7113);
or U7552 (N_7552,N_6012,N_6915);
nand U7553 (N_7553,N_7232,N_6490);
nor U7554 (N_7554,N_6568,N_6127);
or U7555 (N_7555,N_6854,N_7290);
xnor U7556 (N_7556,N_6261,N_7391);
xnor U7557 (N_7557,N_6903,N_6046);
or U7558 (N_7558,N_7011,N_7176);
xor U7559 (N_7559,N_7412,N_6430);
or U7560 (N_7560,N_7255,N_6845);
xnor U7561 (N_7561,N_7160,N_6906);
nor U7562 (N_7562,N_6103,N_7293);
nor U7563 (N_7563,N_7244,N_6782);
nand U7564 (N_7564,N_7418,N_6766);
and U7565 (N_7565,N_6635,N_7085);
or U7566 (N_7566,N_7469,N_6093);
nor U7567 (N_7567,N_7462,N_7197);
or U7568 (N_7568,N_6512,N_6863);
or U7569 (N_7569,N_6543,N_6744);
xnor U7570 (N_7570,N_6070,N_7451);
nor U7571 (N_7571,N_6951,N_6434);
or U7572 (N_7572,N_6094,N_6384);
nor U7573 (N_7573,N_6637,N_6106);
or U7574 (N_7574,N_7029,N_6463);
nor U7575 (N_7575,N_6112,N_6701);
xor U7576 (N_7576,N_6130,N_6979);
nand U7577 (N_7577,N_6914,N_6867);
xor U7578 (N_7578,N_7014,N_6329);
or U7579 (N_7579,N_6303,N_6920);
and U7580 (N_7580,N_6378,N_6123);
and U7581 (N_7581,N_6764,N_7329);
nor U7582 (N_7582,N_6461,N_7179);
or U7583 (N_7583,N_7177,N_6677);
xnor U7584 (N_7584,N_6482,N_6628);
nor U7585 (N_7585,N_6874,N_7322);
and U7586 (N_7586,N_6797,N_6085);
and U7587 (N_7587,N_6274,N_6353);
or U7588 (N_7588,N_6150,N_6087);
or U7589 (N_7589,N_7060,N_7088);
and U7590 (N_7590,N_6860,N_6761);
or U7591 (N_7591,N_6980,N_6785);
and U7592 (N_7592,N_6777,N_7380);
or U7593 (N_7593,N_6059,N_6264);
or U7594 (N_7594,N_6187,N_7157);
xor U7595 (N_7595,N_6339,N_6007);
and U7596 (N_7596,N_7477,N_6504);
nand U7597 (N_7597,N_6667,N_7277);
nor U7598 (N_7598,N_6423,N_6205);
nand U7599 (N_7599,N_6418,N_7443);
xnor U7600 (N_7600,N_7220,N_6402);
nand U7601 (N_7601,N_6483,N_7386);
nor U7602 (N_7602,N_6315,N_7366);
xor U7603 (N_7603,N_7476,N_6148);
or U7604 (N_7604,N_7050,N_6312);
xor U7605 (N_7605,N_6617,N_7049);
xnor U7606 (N_7606,N_7433,N_6165);
or U7607 (N_7607,N_6081,N_6562);
nand U7608 (N_7608,N_6927,N_6842);
or U7609 (N_7609,N_6018,N_7158);
or U7610 (N_7610,N_6567,N_6578);
xnor U7611 (N_7611,N_6086,N_6426);
nor U7612 (N_7612,N_6533,N_6346);
nor U7613 (N_7613,N_6944,N_6754);
or U7614 (N_7614,N_6642,N_6843);
and U7615 (N_7615,N_7151,N_6886);
nand U7616 (N_7616,N_6214,N_6293);
xnor U7617 (N_7617,N_7448,N_6209);
and U7618 (N_7618,N_6844,N_7004);
xor U7619 (N_7619,N_6928,N_6869);
or U7620 (N_7620,N_6275,N_6338);
xor U7621 (N_7621,N_7042,N_6215);
nor U7622 (N_7622,N_6509,N_7155);
and U7623 (N_7623,N_6283,N_6976);
nor U7624 (N_7624,N_6221,N_7037);
or U7625 (N_7625,N_6138,N_6288);
nor U7626 (N_7626,N_7096,N_7215);
nand U7627 (N_7627,N_6424,N_6699);
and U7628 (N_7628,N_6905,N_7402);
and U7629 (N_7629,N_6089,N_7394);
xor U7630 (N_7630,N_6243,N_6257);
nand U7631 (N_7631,N_7259,N_7278);
nand U7632 (N_7632,N_6973,N_6219);
xnor U7633 (N_7633,N_6357,N_6776);
or U7634 (N_7634,N_6479,N_7036);
nand U7635 (N_7635,N_6270,N_6140);
xor U7636 (N_7636,N_7304,N_6669);
nor U7637 (N_7637,N_6682,N_6803);
or U7638 (N_7638,N_6657,N_6220);
and U7639 (N_7639,N_6736,N_6088);
or U7640 (N_7640,N_6466,N_7321);
xor U7641 (N_7641,N_6039,N_6950);
nor U7642 (N_7642,N_7193,N_6580);
nand U7643 (N_7643,N_6111,N_7487);
xor U7644 (N_7644,N_6188,N_7110);
xor U7645 (N_7645,N_6573,N_6815);
xor U7646 (N_7646,N_6948,N_6672);
nand U7647 (N_7647,N_6320,N_6325);
nor U7648 (N_7648,N_6210,N_6704);
xnor U7649 (N_7649,N_6640,N_7337);
nand U7650 (N_7650,N_6666,N_7350);
nand U7651 (N_7651,N_7361,N_6406);
and U7652 (N_7652,N_7311,N_7114);
nand U7653 (N_7653,N_6593,N_6620);
nand U7654 (N_7654,N_7352,N_6160);
xor U7655 (N_7655,N_7239,N_6276);
or U7656 (N_7656,N_7013,N_6115);
and U7657 (N_7657,N_6476,N_6465);
nand U7658 (N_7658,N_6155,N_6826);
nor U7659 (N_7659,N_7463,N_6784);
xor U7660 (N_7660,N_7040,N_6622);
or U7661 (N_7661,N_7466,N_7214);
xnor U7662 (N_7662,N_6726,N_6853);
nor U7663 (N_7663,N_6175,N_7198);
nand U7664 (N_7664,N_6011,N_6082);
nor U7665 (N_7665,N_6134,N_6374);
or U7666 (N_7666,N_7057,N_6592);
or U7667 (N_7667,N_6818,N_7238);
xor U7668 (N_7668,N_7263,N_6208);
nor U7669 (N_7669,N_6519,N_6992);
nor U7670 (N_7670,N_6201,N_6960);
nor U7671 (N_7671,N_6416,N_6090);
xor U7672 (N_7672,N_7133,N_7415);
nand U7673 (N_7673,N_7136,N_6232);
and U7674 (N_7674,N_6662,N_6549);
and U7675 (N_7675,N_6189,N_6331);
or U7676 (N_7676,N_6297,N_7204);
and U7677 (N_7677,N_6043,N_6225);
nand U7678 (N_7678,N_7456,N_7295);
nand U7679 (N_7679,N_7430,N_7161);
or U7680 (N_7680,N_7461,N_6145);
xor U7681 (N_7681,N_7112,N_7353);
nor U7682 (N_7682,N_7076,N_6433);
and U7683 (N_7683,N_7184,N_6008);
or U7684 (N_7684,N_6332,N_6459);
and U7685 (N_7685,N_6805,N_6627);
xor U7686 (N_7686,N_7262,N_6684);
and U7687 (N_7687,N_6213,N_7368);
xor U7688 (N_7688,N_6054,N_6300);
xor U7689 (N_7689,N_7474,N_6299);
xnor U7690 (N_7690,N_7400,N_6733);
and U7691 (N_7691,N_6449,N_6752);
xor U7692 (N_7692,N_6249,N_7356);
nor U7693 (N_7693,N_7219,N_7413);
xor U7694 (N_7694,N_7016,N_7073);
nor U7695 (N_7695,N_6269,N_6993);
nand U7696 (N_7696,N_7494,N_7387);
xor U7697 (N_7697,N_6323,N_6142);
or U7698 (N_7698,N_7328,N_6639);
nor U7699 (N_7699,N_7478,N_7213);
nand U7700 (N_7700,N_6584,N_6837);
or U7701 (N_7701,N_6069,N_7331);
nor U7702 (N_7702,N_6136,N_7245);
nor U7703 (N_7703,N_6872,N_7121);
xnor U7704 (N_7704,N_6551,N_7475);
and U7705 (N_7705,N_6922,N_6661);
xnor U7706 (N_7706,N_6453,N_6711);
xor U7707 (N_7707,N_6073,N_6460);
xor U7708 (N_7708,N_6027,N_7334);
nand U7709 (N_7709,N_7175,N_6045);
or U7710 (N_7710,N_6196,N_6946);
and U7711 (N_7711,N_6675,N_6859);
nand U7712 (N_7712,N_7131,N_6751);
and U7713 (N_7713,N_6387,N_7118);
and U7714 (N_7714,N_6240,N_7496);
or U7715 (N_7715,N_7008,N_7183);
xor U7716 (N_7716,N_6643,N_6404);
xnor U7717 (N_7717,N_6819,N_7127);
nand U7718 (N_7718,N_6885,N_6500);
or U7719 (N_7719,N_6010,N_7484);
nor U7720 (N_7720,N_6603,N_6884);
nand U7721 (N_7721,N_6840,N_6255);
or U7722 (N_7722,N_6646,N_7336);
xnor U7723 (N_7723,N_6560,N_7148);
nand U7724 (N_7724,N_6427,N_7281);
xor U7725 (N_7725,N_6147,N_7495);
or U7726 (N_7726,N_7374,N_6817);
nor U7727 (N_7727,N_7468,N_6231);
nor U7728 (N_7728,N_7341,N_7228);
and U7729 (N_7729,N_6907,N_6982);
xnor U7730 (N_7730,N_6095,N_6097);
xnor U7731 (N_7731,N_6534,N_6282);
and U7732 (N_7732,N_6480,N_6912);
nand U7733 (N_7733,N_6149,N_6858);
and U7734 (N_7734,N_6623,N_6779);
and U7735 (N_7735,N_6924,N_6795);
xnor U7736 (N_7736,N_7288,N_6926);
nand U7737 (N_7737,N_7426,N_7143);
or U7738 (N_7738,N_6290,N_7492);
xor U7739 (N_7739,N_6203,N_7075);
nor U7740 (N_7740,N_6350,N_6961);
or U7741 (N_7741,N_7438,N_7066);
xnor U7742 (N_7742,N_7128,N_6049);
nand U7743 (N_7743,N_6999,N_6379);
nand U7744 (N_7744,N_6173,N_6197);
and U7745 (N_7745,N_6322,N_7250);
and U7746 (N_7746,N_6890,N_6120);
nor U7747 (N_7747,N_6185,N_6464);
xor U7748 (N_7748,N_6848,N_7335);
and U7749 (N_7749,N_6435,N_7223);
or U7750 (N_7750,N_7384,N_6892);
nand U7751 (N_7751,N_6941,N_6822);
and U7752 (N_7752,N_6607,N_7453);
and U7753 (N_7753,N_6484,N_7165);
nand U7754 (N_7754,N_6780,N_7276);
nor U7755 (N_7755,N_6141,N_7490);
nor U7756 (N_7756,N_7362,N_6362);
or U7757 (N_7757,N_6746,N_7312);
and U7758 (N_7758,N_6577,N_6117);
or U7759 (N_7759,N_6491,N_6473);
and U7760 (N_7760,N_6878,N_6137);
or U7761 (N_7761,N_7126,N_6234);
xor U7762 (N_7762,N_6119,N_6688);
or U7763 (N_7763,N_7190,N_6436);
or U7764 (N_7764,N_6241,N_7333);
nor U7765 (N_7765,N_7188,N_6388);
xor U7766 (N_7766,N_6532,N_6756);
nor U7767 (N_7767,N_6347,N_6718);
xnor U7768 (N_7768,N_6556,N_7455);
xnor U7769 (N_7769,N_6548,N_7452);
nor U7770 (N_7770,N_7420,N_7437);
xnor U7771 (N_7771,N_6077,N_6262);
and U7772 (N_7772,N_7306,N_6864);
nor U7773 (N_7773,N_6053,N_6172);
or U7774 (N_7774,N_6277,N_6507);
and U7775 (N_7775,N_6495,N_7163);
nand U7776 (N_7776,N_6601,N_7226);
nor U7777 (N_7777,N_6652,N_6887);
xor U7778 (N_7778,N_6349,N_6184);
xor U7779 (N_7779,N_6816,N_6105);
and U7780 (N_7780,N_6870,N_6177);
nor U7781 (N_7781,N_7377,N_7038);
and U7782 (N_7782,N_6061,N_6468);
or U7783 (N_7783,N_7497,N_6135);
xnor U7784 (N_7784,N_7272,N_6066);
and U7785 (N_7785,N_7358,N_6023);
xnor U7786 (N_7786,N_6831,N_6943);
nand U7787 (N_7787,N_6381,N_7162);
and U7788 (N_7788,N_6099,N_7376);
or U7789 (N_7789,N_6207,N_7167);
nor U7790 (N_7790,N_6621,N_6064);
and U7791 (N_7791,N_7308,N_6908);
or U7792 (N_7792,N_7129,N_7144);
nor U7793 (N_7793,N_6032,N_6079);
and U7794 (N_7794,N_6498,N_6326);
nand U7795 (N_7795,N_6918,N_6037);
xor U7796 (N_7796,N_7283,N_6740);
nor U7797 (N_7797,N_7091,N_6686);
xnor U7798 (N_7798,N_6492,N_7317);
nor U7799 (N_7799,N_7235,N_6348);
and U7800 (N_7800,N_6762,N_6367);
and U7801 (N_7801,N_6625,N_6398);
nand U7802 (N_7802,N_6366,N_6898);
nor U7803 (N_7803,N_6681,N_6132);
xnor U7804 (N_7804,N_6113,N_6013);
nor U7805 (N_7805,N_7241,N_6442);
nor U7806 (N_7806,N_7485,N_6995);
or U7807 (N_7807,N_6389,N_6502);
or U7808 (N_7808,N_6773,N_6820);
or U7809 (N_7809,N_7111,N_6707);
or U7810 (N_7810,N_7480,N_6810);
nor U7811 (N_7811,N_6553,N_6644);
nor U7812 (N_7812,N_6865,N_6952);
and U7813 (N_7813,N_6563,N_6517);
nand U7814 (N_7814,N_6737,N_7315);
and U7815 (N_7815,N_6983,N_6585);
and U7816 (N_7816,N_6361,N_7222);
nor U7817 (N_7817,N_6396,N_6048);
nand U7818 (N_7818,N_6687,N_7007);
nor U7819 (N_7819,N_7388,N_7185);
or U7820 (N_7820,N_7166,N_6044);
nor U7821 (N_7821,N_7360,N_6015);
nand U7822 (N_7822,N_7488,N_7172);
nor U7823 (N_7823,N_7472,N_6497);
nand U7824 (N_7824,N_6009,N_7498);
nor U7825 (N_7825,N_7125,N_6454);
and U7826 (N_7826,N_6636,N_7052);
xnor U7827 (N_7827,N_7369,N_6448);
or U7828 (N_7828,N_6765,N_6179);
and U7829 (N_7829,N_6000,N_6986);
and U7830 (N_7830,N_7090,N_6334);
nand U7831 (N_7831,N_6020,N_6899);
nand U7832 (N_7832,N_6917,N_6629);
xor U7833 (N_7833,N_7225,N_7429);
nor U7834 (N_7834,N_6072,N_6581);
or U7835 (N_7835,N_6963,N_6407);
nand U7836 (N_7836,N_6359,N_6741);
nor U7837 (N_7837,N_7314,N_6713);
xor U7838 (N_7838,N_7457,N_6352);
and U7839 (N_7839,N_6956,N_6850);
nand U7840 (N_7840,N_7145,N_7460);
nand U7841 (N_7841,N_6472,N_6558);
xnor U7842 (N_7842,N_6862,N_7001);
xnor U7843 (N_7843,N_6763,N_7318);
xnor U7844 (N_7844,N_6031,N_6630);
xor U7845 (N_7845,N_6594,N_6217);
xor U7846 (N_7846,N_6739,N_6178);
xor U7847 (N_7847,N_6934,N_6056);
and U7848 (N_7848,N_6324,N_6597);
nand U7849 (N_7849,N_7063,N_7401);
nand U7850 (N_7850,N_6005,N_6583);
nor U7851 (N_7851,N_6432,N_7382);
and U7852 (N_7852,N_6868,N_6876);
and U7853 (N_7853,N_7324,N_6488);
nor U7854 (N_7854,N_6146,N_7154);
or U7855 (N_7855,N_6586,N_6709);
nand U7856 (N_7856,N_7086,N_6058);
nand U7857 (N_7857,N_6298,N_6871);
nor U7858 (N_7858,N_6170,N_6645);
nand U7859 (N_7859,N_7195,N_7459);
and U7860 (N_7860,N_7261,N_6540);
xor U7861 (N_7861,N_6827,N_7275);
nand U7862 (N_7862,N_7491,N_6608);
nor U7863 (N_7863,N_6485,N_6311);
or U7864 (N_7864,N_6997,N_7146);
or U7865 (N_7865,N_6561,N_6144);
or U7866 (N_7866,N_6372,N_6919);
nand U7867 (N_7867,N_6028,N_7270);
nand U7868 (N_7868,N_6405,N_6857);
xnor U7869 (N_7869,N_7233,N_6571);
nor U7870 (N_7870,N_6550,N_6953);
nand U7871 (N_7871,N_6789,N_7021);
nor U7872 (N_7872,N_6697,N_6904);
xor U7873 (N_7873,N_6354,N_6096);
nand U7874 (N_7874,N_7248,N_6921);
nor U7875 (N_7875,N_6942,N_6579);
nand U7876 (N_7876,N_7139,N_7499);
nand U7877 (N_7877,N_6002,N_6957);
and U7878 (N_7878,N_7323,N_6431);
nor U7879 (N_7879,N_7473,N_6450);
nor U7880 (N_7880,N_7093,N_7104);
xnor U7881 (N_7881,N_6846,N_7440);
nand U7882 (N_7882,N_7030,N_6273);
and U7883 (N_7883,N_7051,N_6588);
and U7884 (N_7884,N_6937,N_7039);
or U7885 (N_7885,N_7141,N_6098);
or U7886 (N_7886,N_7349,N_6683);
and U7887 (N_7887,N_6531,N_6768);
nand U7888 (N_7888,N_7169,N_7027);
nor U7889 (N_7889,N_7363,N_6808);
and U7890 (N_7890,N_6198,N_6291);
xor U7891 (N_7891,N_6109,N_6286);
nand U7892 (N_7892,N_6566,N_7483);
and U7893 (N_7893,N_7273,N_7072);
xor U7894 (N_7894,N_7168,N_6457);
or U7895 (N_7895,N_7002,N_6589);
nand U7896 (N_7896,N_6771,N_7058);
and U7897 (N_7897,N_6655,N_6373);
nor U7898 (N_7898,N_6911,N_6057);
nor U7899 (N_7899,N_6778,N_7130);
nand U7900 (N_7900,N_6749,N_7449);
xor U7901 (N_7901,N_7105,N_6658);
xor U7902 (N_7902,N_7330,N_6245);
or U7903 (N_7903,N_6606,N_7340);
or U7904 (N_7904,N_6954,N_7431);
xnor U7905 (N_7905,N_7000,N_6757);
and U7906 (N_7906,N_7303,N_6268);
or U7907 (N_7907,N_6981,N_7383);
and U7908 (N_7908,N_6546,N_7009);
xnor U7909 (N_7909,N_7447,N_6962);
nor U7910 (N_7910,N_6877,N_6564);
xor U7911 (N_7911,N_6246,N_6659);
or U7912 (N_7912,N_6164,N_6462);
or U7913 (N_7913,N_6494,N_6368);
or U7914 (N_7914,N_7043,N_6309);
or U7915 (N_7915,N_6725,N_6122);
xnor U7916 (N_7916,N_6823,N_7097);
nand U7917 (N_7917,N_7257,N_7117);
or U7918 (N_7918,N_6720,N_6344);
nand U7919 (N_7919,N_6716,N_6247);
and U7920 (N_7920,N_7397,N_6668);
or U7921 (N_7921,N_7302,N_6158);
nand U7922 (N_7922,N_6156,N_6799);
and U7923 (N_7923,N_6835,N_6118);
xnor U7924 (N_7924,N_7062,N_7054);
or U7925 (N_7925,N_6619,N_7355);
nor U7926 (N_7926,N_6345,N_6614);
nor U7927 (N_7927,N_6665,N_6511);
xor U7928 (N_7928,N_6318,N_7260);
and U7929 (N_7929,N_6412,N_6306);
or U7930 (N_7930,N_6024,N_6590);
nand U7931 (N_7931,N_6316,N_7403);
nor U7932 (N_7932,N_6397,N_7237);
nand U7933 (N_7933,N_7061,N_7458);
xor U7934 (N_7934,N_7053,N_6055);
xnor U7935 (N_7935,N_6244,N_6596);
xnor U7936 (N_7936,N_6104,N_6861);
or U7937 (N_7937,N_6166,N_7253);
or U7938 (N_7938,N_7365,N_6191);
and U7939 (N_7939,N_6445,N_6991);
nand U7940 (N_7940,N_6913,N_6342);
nor U7941 (N_7941,N_6626,N_7134);
xor U7942 (N_7942,N_6852,N_6419);
nand U7943 (N_7943,N_7017,N_7092);
or U7944 (N_7944,N_7285,N_6794);
xor U7945 (N_7945,N_6458,N_7342);
nand U7946 (N_7946,N_6545,N_6080);
nand U7947 (N_7947,N_7035,N_7434);
and U7948 (N_7948,N_6313,N_6897);
xnor U7949 (N_7949,N_6994,N_7221);
nand U7950 (N_7950,N_6775,N_7227);
and U7951 (N_7951,N_6839,N_6356);
and U7952 (N_7952,N_7446,N_6143);
xor U7953 (N_7953,N_7299,N_6351);
nand U7954 (N_7954,N_6295,N_6236);
and U7955 (N_7955,N_6071,N_6801);
nor U7956 (N_7956,N_6654,N_6758);
xnor U7957 (N_7957,N_7095,N_6615);
and U7958 (N_7958,N_7298,N_6211);
nand U7959 (N_7959,N_6408,N_7102);
xor U7960 (N_7960,N_6499,N_7422);
nand U7961 (N_7961,N_6428,N_6182);
xnor U7962 (N_7962,N_6518,N_6451);
nand U7963 (N_7963,N_7206,N_7234);
nand U7964 (N_7964,N_6266,N_6260);
xor U7965 (N_7965,N_6310,N_7019);
xnor U7966 (N_7966,N_7381,N_7364);
nand U7967 (N_7967,N_7189,N_6824);
nor U7968 (N_7968,N_7243,N_6633);
and U7969 (N_7969,N_7064,N_6989);
xor U7970 (N_7970,N_7291,N_6841);
or U7971 (N_7971,N_6515,N_6278);
or U7972 (N_7972,N_6769,N_6194);
xor U7973 (N_7973,N_7003,N_7347);
xor U7974 (N_7974,N_6847,N_7089);
and U7975 (N_7975,N_7313,N_6399);
and U7976 (N_7976,N_7406,N_7294);
xor U7977 (N_7977,N_6163,N_6154);
nand U7978 (N_7978,N_6228,N_7182);
and U7979 (N_7979,N_6930,N_6734);
xor U7980 (N_7980,N_6017,N_6900);
nand U7981 (N_7981,N_7147,N_6851);
nand U7982 (N_7982,N_6248,N_6503);
and U7983 (N_7983,N_7068,N_6896);
nand U7984 (N_7984,N_6939,N_7109);
xnor U7985 (N_7985,N_7367,N_6267);
xnor U7986 (N_7986,N_7399,N_6304);
nand U7987 (N_7987,N_6237,N_6727);
nor U7988 (N_7988,N_6663,N_6557);
and U7989 (N_7989,N_6881,N_6474);
nand U7990 (N_7990,N_6074,N_6591);
nand U7991 (N_7991,N_7325,N_7209);
nor U7992 (N_7992,N_6833,N_6559);
nor U7993 (N_7993,N_6949,N_6516);
nor U7994 (N_7994,N_6493,N_6041);
nand U7995 (N_7995,N_7047,N_7249);
nor U7996 (N_7996,N_6092,N_7470);
nor U7997 (N_7997,N_6216,N_6714);
and U7998 (N_7998,N_7180,N_6029);
or U7999 (N_7999,N_6696,N_7419);
nor U8000 (N_8000,N_7486,N_6722);
nor U8001 (N_8001,N_7271,N_7266);
and U8002 (N_8002,N_6307,N_6383);
nor U8003 (N_8003,N_6369,N_7018);
or U8004 (N_8004,N_6014,N_6308);
and U8005 (N_8005,N_6855,N_6582);
xor U8006 (N_8006,N_6238,N_7108);
nand U8007 (N_8007,N_7231,N_6856);
or U8008 (N_8008,N_6967,N_6730);
xnor U8009 (N_8009,N_6471,N_6265);
xnor U8010 (N_8010,N_6047,N_7207);
and U8011 (N_8011,N_7216,N_6226);
nor U8012 (N_8012,N_6972,N_6883);
or U8013 (N_8013,N_6964,N_7408);
nor U8014 (N_8014,N_6616,N_6783);
nand U8015 (N_8015,N_6417,N_6343);
or U8016 (N_8016,N_6108,N_7300);
nand U8017 (N_8017,N_6806,N_7116);
nand U8018 (N_8018,N_6385,N_6574);
and U8019 (N_8019,N_6259,N_6610);
nor U8020 (N_8020,N_7267,N_7398);
nor U8021 (N_8021,N_6958,N_6728);
nor U8022 (N_8022,N_7083,N_6478);
and U8023 (N_8023,N_7348,N_7395);
or U8024 (N_8024,N_6068,N_6016);
nor U8025 (N_8025,N_6169,N_6319);
xor U8026 (N_8026,N_7024,N_7153);
nand U8027 (N_8027,N_7192,N_6167);
xor U8028 (N_8028,N_6252,N_6377);
xor U8029 (N_8029,N_6541,N_6676);
nor U8030 (N_8030,N_7025,N_6674);
and U8031 (N_8031,N_6793,N_6067);
or U8032 (N_8032,N_6287,N_6422);
nor U8033 (N_8033,N_7404,N_7251);
xor U8034 (N_8034,N_7450,N_7201);
nor U8035 (N_8035,N_6370,N_7236);
nor U8036 (N_8036,N_7170,N_7033);
or U8037 (N_8037,N_6202,N_6116);
xor U8038 (N_8038,N_6280,N_7407);
or U8039 (N_8039,N_6786,N_6506);
or U8040 (N_8040,N_6602,N_7409);
and U8041 (N_8041,N_6708,N_6302);
nand U8042 (N_8042,N_6258,N_6425);
nand U8043 (N_8043,N_6738,N_6651);
and U8044 (N_8044,N_7218,N_7028);
xnor U8045 (N_8045,N_7454,N_6528);
or U8046 (N_8046,N_7301,N_7099);
or U8047 (N_8047,N_6955,N_6732);
or U8048 (N_8048,N_7048,N_6882);
nor U8049 (N_8049,N_7138,N_6624);
xnor U8050 (N_8050,N_7087,N_6413);
nor U8051 (N_8051,N_7026,N_6742);
xor U8052 (N_8052,N_6552,N_6410);
nor U8053 (N_8053,N_6599,N_6161);
and U8054 (N_8054,N_6968,N_6200);
and U8055 (N_8055,N_6125,N_6129);
nand U8056 (N_8056,N_6706,N_6171);
and U8057 (N_8057,N_6604,N_6970);
nor U8058 (N_8058,N_7055,N_6371);
and U8059 (N_8059,N_6174,N_7378);
nand U8060 (N_8060,N_6632,N_6409);
xnor U8061 (N_8061,N_6218,N_7274);
and U8062 (N_8062,N_7435,N_7005);
xor U8063 (N_8063,N_7150,N_6363);
nor U8064 (N_8064,N_6242,N_6375);
and U8065 (N_8065,N_6724,N_6469);
nand U8066 (N_8066,N_7071,N_6695);
or U8067 (N_8067,N_6811,N_6660);
nor U8068 (N_8068,N_6042,N_7186);
or U8069 (N_8069,N_6486,N_6446);
xor U8070 (N_8070,N_7212,N_6294);
xnor U8071 (N_8071,N_6712,N_7135);
or U8072 (N_8072,N_6284,N_6444);
nor U8073 (N_8073,N_7202,N_6618);
nand U8074 (N_8074,N_7346,N_6829);
or U8075 (N_8075,N_6555,N_6925);
xor U8076 (N_8076,N_6717,N_7345);
and U8077 (N_8077,N_6996,N_6030);
or U8078 (N_8078,N_6025,N_6969);
nor U8079 (N_8079,N_7375,N_7079);
xor U8080 (N_8080,N_6916,N_6487);
nand U8081 (N_8081,N_6702,N_7140);
or U8082 (N_8082,N_6965,N_6974);
and U8083 (N_8083,N_6159,N_6875);
and U8084 (N_8084,N_6788,N_7247);
and U8085 (N_8085,N_6729,N_6513);
nand U8086 (N_8086,N_7115,N_7012);
or U8087 (N_8087,N_6544,N_6671);
nand U8088 (N_8088,N_6747,N_6401);
nand U8089 (N_8089,N_7246,N_6542);
nor U8090 (N_8090,N_6075,N_7411);
nor U8091 (N_8091,N_6514,N_6078);
xor U8092 (N_8092,N_7344,N_6650);
and U8093 (N_8093,N_6033,N_7041);
and U8094 (N_8094,N_6812,N_6664);
xnor U8095 (N_8095,N_6595,N_6576);
xor U8096 (N_8096,N_6429,N_6656);
and U8097 (N_8097,N_6673,N_7044);
nor U8098 (N_8098,N_7416,N_6301);
xor U8099 (N_8099,N_6263,N_7254);
and U8100 (N_8100,N_6467,N_7191);
and U8101 (N_8101,N_6124,N_6022);
or U8102 (N_8102,N_7081,N_6392);
or U8103 (N_8103,N_7310,N_6003);
or U8104 (N_8104,N_6570,N_6587);
and U8105 (N_8105,N_6206,N_7200);
nand U8106 (N_8106,N_6341,N_6554);
and U8107 (N_8107,N_7390,N_7441);
nor U8108 (N_8108,N_6390,N_6648);
nand U8109 (N_8109,N_7015,N_6977);
or U8110 (N_8110,N_6452,N_6959);
or U8111 (N_8111,N_6529,N_6051);
and U8112 (N_8112,N_7217,N_7119);
or U8113 (N_8113,N_6834,N_7142);
nand U8114 (N_8114,N_6693,N_7354);
xor U8115 (N_8115,N_7296,N_6382);
xnor U8116 (N_8116,N_7436,N_6443);
or U8117 (N_8117,N_6121,N_6735);
and U8118 (N_8118,N_6400,N_7101);
or U8119 (N_8119,N_7078,N_6441);
xnor U8120 (N_8120,N_6975,N_6910);
nand U8121 (N_8121,N_7465,N_6527);
or U8122 (N_8122,N_6653,N_6750);
and U8123 (N_8123,N_6229,N_6894);
nand U8124 (N_8124,N_6849,N_6411);
and U8125 (N_8125,N_6420,N_7103);
nand U8126 (N_8126,N_7280,N_6828);
xor U8127 (N_8127,N_6678,N_7371);
nor U8128 (N_8128,N_7351,N_6110);
xor U8129 (N_8129,N_6613,N_6364);
xor U8130 (N_8130,N_6101,N_6770);
and U8131 (N_8131,N_7372,N_7084);
xnor U8132 (N_8132,N_7289,N_6767);
and U8133 (N_8133,N_7240,N_7230);
and U8134 (N_8134,N_6223,N_6804);
xor U8135 (N_8135,N_7100,N_6314);
nor U8136 (N_8136,N_6114,N_7046);
and U8137 (N_8137,N_6760,N_7137);
or U8138 (N_8138,N_6609,N_6649);
nor U8139 (N_8139,N_6800,N_7357);
nor U8140 (N_8140,N_6929,N_6745);
nor U8141 (N_8141,N_6224,N_6279);
and U8142 (N_8142,N_6131,N_6933);
or U8143 (N_8143,N_7439,N_7205);
nor U8144 (N_8144,N_7292,N_7196);
and U8145 (N_8145,N_6888,N_6292);
nand U8146 (N_8146,N_6195,N_6985);
and U8147 (N_8147,N_7425,N_6879);
nor U8148 (N_8148,N_7287,N_6522);
and U8149 (N_8149,N_6133,N_6932);
nor U8150 (N_8150,N_6759,N_6792);
and U8151 (N_8151,N_6525,N_6062);
nand U8152 (N_8152,N_6988,N_7444);
nor U8153 (N_8153,N_6076,N_6336);
xnor U8154 (N_8154,N_6251,N_6360);
nand U8155 (N_8155,N_6889,N_7032);
nor U8156 (N_8156,N_6821,N_7445);
nand U8157 (N_8157,N_7269,N_6605);
xnor U8158 (N_8158,N_7107,N_6670);
nor U8159 (N_8159,N_7098,N_6139);
nor U8160 (N_8160,N_7268,N_6296);
xor U8161 (N_8161,N_6063,N_7359);
xor U8162 (N_8162,N_6193,N_7424);
and U8163 (N_8163,N_6190,N_6126);
nor U8164 (N_8164,N_6250,N_6523);
nand U8165 (N_8165,N_7489,N_7284);
nor U8166 (N_8166,N_6456,N_7077);
nand U8167 (N_8167,N_7464,N_7229);
nand U8168 (N_8168,N_6330,N_7467);
and U8169 (N_8169,N_6035,N_6691);
xnor U8170 (N_8170,N_7187,N_6380);
and U8171 (N_8171,N_7332,N_6321);
nor U8172 (N_8172,N_6940,N_6157);
and U8173 (N_8173,N_6510,N_7479);
or U8174 (N_8174,N_6317,N_6931);
nor U8175 (N_8175,N_7056,N_6340);
nor U8176 (N_8176,N_6520,N_6873);
nand U8177 (N_8177,N_6705,N_6945);
xnor U8178 (N_8178,N_7343,N_7423);
xnor U8179 (N_8179,N_6477,N_6703);
and U8180 (N_8180,N_6715,N_7094);
nor U8181 (N_8181,N_7421,N_6181);
or U8182 (N_8182,N_6328,N_7082);
or U8183 (N_8183,N_7178,N_6052);
and U8184 (N_8184,N_7106,N_6638);
xnor U8185 (N_8185,N_6600,N_7210);
or U8186 (N_8186,N_6365,N_7471);
nor U8187 (N_8187,N_6337,N_7396);
nand U8188 (N_8188,N_6538,N_6153);
nand U8189 (N_8189,N_6475,N_6612);
or U8190 (N_8190,N_6978,N_6634);
xor U8191 (N_8191,N_6180,N_6987);
nand U8192 (N_8192,N_6598,N_6391);
xnor U8193 (N_8193,N_6271,N_6230);
xnor U8194 (N_8194,N_6787,N_6791);
xnor U8195 (N_8195,N_6731,N_6936);
nor U8196 (N_8196,N_6168,N_7023);
and U8197 (N_8197,N_6813,N_6700);
nand U8198 (N_8198,N_6935,N_6631);
nor U8199 (N_8199,N_7224,N_6830);
xnor U8200 (N_8200,N_6901,N_7410);
nand U8201 (N_8201,N_7389,N_7442);
xnor U8202 (N_8202,N_6227,N_7286);
xnor U8203 (N_8203,N_6524,N_6001);
nor U8204 (N_8204,N_6395,N_6199);
nor U8205 (N_8205,N_7242,N_7405);
and U8206 (N_8206,N_7080,N_6437);
nor U8207 (N_8207,N_6102,N_7493);
nand U8208 (N_8208,N_6192,N_7370);
or U8209 (N_8209,N_6006,N_6004);
nand U8210 (N_8210,N_7181,N_7006);
nor U8211 (N_8211,N_6923,N_6470);
or U8212 (N_8212,N_6891,N_6421);
nor U8213 (N_8213,N_7339,N_6021);
or U8214 (N_8214,N_7282,N_6880);
or U8215 (N_8215,N_6060,N_6814);
nand U8216 (N_8216,N_6254,N_6807);
or U8217 (N_8217,N_7034,N_6040);
nor U8218 (N_8218,N_6825,N_6327);
xnor U8219 (N_8219,N_6438,N_6641);
and U8220 (N_8220,N_7069,N_6647);
xor U8221 (N_8221,N_7045,N_6083);
nand U8222 (N_8222,N_6547,N_7279);
nand U8223 (N_8223,N_7120,N_6186);
and U8224 (N_8224,N_6537,N_7327);
nor U8225 (N_8225,N_6107,N_7171);
or U8226 (N_8226,N_6680,N_7385);
or U8227 (N_8227,N_7393,N_6575);
nand U8228 (N_8228,N_6909,N_6998);
xor U8229 (N_8229,N_7305,N_7159);
nand U8230 (N_8230,N_6611,N_6050);
nor U8231 (N_8231,N_6743,N_6893);
and U8232 (N_8232,N_6335,N_6984);
or U8233 (N_8233,N_6866,N_6393);
nor U8234 (N_8234,N_6256,N_6176);
nand U8235 (N_8235,N_7264,N_6521);
nor U8236 (N_8236,N_6091,N_6386);
xnor U8237 (N_8237,N_6151,N_6689);
or U8238 (N_8238,N_6235,N_7164);
and U8239 (N_8239,N_6721,N_7074);
and U8240 (N_8240,N_6710,N_6355);
or U8241 (N_8241,N_6212,N_7199);
and U8242 (N_8242,N_6034,N_6838);
or U8243 (N_8243,N_6496,N_6565);
or U8244 (N_8244,N_6414,N_7432);
or U8245 (N_8245,N_7338,N_6685);
xnor U8246 (N_8246,N_6222,N_6809);
or U8247 (N_8247,N_6772,N_7203);
and U8248 (N_8248,N_6285,N_6065);
nand U8249 (N_8249,N_6272,N_7020);
nor U8250 (N_8250,N_6527,N_6908);
nand U8251 (N_8251,N_6667,N_6178);
nand U8252 (N_8252,N_6778,N_6673);
or U8253 (N_8253,N_7384,N_6359);
nand U8254 (N_8254,N_6465,N_7275);
xnor U8255 (N_8255,N_6019,N_6886);
xor U8256 (N_8256,N_6685,N_7472);
nand U8257 (N_8257,N_6898,N_6421);
xnor U8258 (N_8258,N_7202,N_7154);
nand U8259 (N_8259,N_7136,N_6134);
nand U8260 (N_8260,N_6081,N_6482);
nor U8261 (N_8261,N_6781,N_7196);
and U8262 (N_8262,N_7395,N_7156);
nor U8263 (N_8263,N_6590,N_6011);
and U8264 (N_8264,N_7311,N_6697);
nor U8265 (N_8265,N_6975,N_7106);
and U8266 (N_8266,N_7218,N_6039);
and U8267 (N_8267,N_7497,N_7042);
nand U8268 (N_8268,N_6855,N_6190);
and U8269 (N_8269,N_6434,N_6775);
and U8270 (N_8270,N_6077,N_7074);
nand U8271 (N_8271,N_6159,N_7264);
nor U8272 (N_8272,N_6613,N_7066);
or U8273 (N_8273,N_6749,N_7402);
or U8274 (N_8274,N_6519,N_6871);
nand U8275 (N_8275,N_6558,N_7232);
xor U8276 (N_8276,N_6025,N_7384);
xor U8277 (N_8277,N_6876,N_6349);
xnor U8278 (N_8278,N_6801,N_7177);
nor U8279 (N_8279,N_6123,N_6140);
or U8280 (N_8280,N_6606,N_7397);
nand U8281 (N_8281,N_6613,N_6000);
xnor U8282 (N_8282,N_6779,N_6990);
nand U8283 (N_8283,N_6460,N_7114);
nor U8284 (N_8284,N_7162,N_6784);
nor U8285 (N_8285,N_7292,N_6013);
and U8286 (N_8286,N_6585,N_6950);
and U8287 (N_8287,N_6027,N_6670);
and U8288 (N_8288,N_6808,N_6869);
nor U8289 (N_8289,N_6461,N_6283);
nand U8290 (N_8290,N_6394,N_7027);
nor U8291 (N_8291,N_7194,N_6982);
or U8292 (N_8292,N_7190,N_7131);
xor U8293 (N_8293,N_6567,N_6088);
nor U8294 (N_8294,N_7108,N_6369);
and U8295 (N_8295,N_6815,N_6007);
nand U8296 (N_8296,N_6486,N_6560);
nand U8297 (N_8297,N_6812,N_7152);
nor U8298 (N_8298,N_6399,N_6491);
nand U8299 (N_8299,N_6098,N_6050);
or U8300 (N_8300,N_6943,N_6384);
nand U8301 (N_8301,N_6255,N_6224);
and U8302 (N_8302,N_6570,N_6567);
nand U8303 (N_8303,N_6089,N_6173);
nor U8304 (N_8304,N_6788,N_7039);
and U8305 (N_8305,N_6778,N_7001);
and U8306 (N_8306,N_6075,N_6373);
xnor U8307 (N_8307,N_6542,N_6103);
nor U8308 (N_8308,N_7212,N_6220);
and U8309 (N_8309,N_6307,N_7320);
xnor U8310 (N_8310,N_6198,N_6946);
xor U8311 (N_8311,N_7216,N_6372);
nand U8312 (N_8312,N_6079,N_7479);
nor U8313 (N_8313,N_6613,N_6407);
nand U8314 (N_8314,N_7221,N_6490);
and U8315 (N_8315,N_6777,N_6078);
or U8316 (N_8316,N_7180,N_6519);
xor U8317 (N_8317,N_7002,N_7059);
nor U8318 (N_8318,N_7210,N_6779);
nor U8319 (N_8319,N_6631,N_7083);
xor U8320 (N_8320,N_6916,N_7020);
nand U8321 (N_8321,N_6504,N_6781);
and U8322 (N_8322,N_6063,N_7189);
nand U8323 (N_8323,N_7465,N_6868);
xnor U8324 (N_8324,N_6660,N_6032);
nor U8325 (N_8325,N_6380,N_6397);
xnor U8326 (N_8326,N_6502,N_6677);
xor U8327 (N_8327,N_7410,N_6228);
and U8328 (N_8328,N_6494,N_6522);
and U8329 (N_8329,N_6803,N_7193);
nand U8330 (N_8330,N_7308,N_6491);
nand U8331 (N_8331,N_6716,N_6417);
and U8332 (N_8332,N_6468,N_7472);
nor U8333 (N_8333,N_6042,N_7028);
xnor U8334 (N_8334,N_6299,N_6058);
nand U8335 (N_8335,N_7377,N_6088);
nor U8336 (N_8336,N_7360,N_6403);
or U8337 (N_8337,N_6982,N_6973);
xor U8338 (N_8338,N_6920,N_6617);
and U8339 (N_8339,N_6191,N_6461);
or U8340 (N_8340,N_7257,N_6539);
nor U8341 (N_8341,N_6133,N_6063);
xor U8342 (N_8342,N_7204,N_6962);
or U8343 (N_8343,N_6364,N_7006);
nand U8344 (N_8344,N_6926,N_6780);
or U8345 (N_8345,N_6729,N_6086);
and U8346 (N_8346,N_7297,N_6893);
xnor U8347 (N_8347,N_6293,N_6117);
and U8348 (N_8348,N_6369,N_7457);
nand U8349 (N_8349,N_7455,N_6956);
nand U8350 (N_8350,N_7193,N_7155);
nor U8351 (N_8351,N_6410,N_7493);
nand U8352 (N_8352,N_6015,N_6914);
and U8353 (N_8353,N_7080,N_7399);
xor U8354 (N_8354,N_7040,N_6143);
xor U8355 (N_8355,N_7325,N_6828);
and U8356 (N_8356,N_7452,N_6155);
nand U8357 (N_8357,N_6675,N_7259);
and U8358 (N_8358,N_6965,N_6057);
nor U8359 (N_8359,N_7460,N_6348);
nand U8360 (N_8360,N_6313,N_6468);
xor U8361 (N_8361,N_6559,N_6847);
xnor U8362 (N_8362,N_6544,N_7222);
nor U8363 (N_8363,N_6336,N_6579);
xor U8364 (N_8364,N_7349,N_6927);
and U8365 (N_8365,N_7207,N_6319);
xor U8366 (N_8366,N_6508,N_7176);
or U8367 (N_8367,N_6226,N_7009);
or U8368 (N_8368,N_6327,N_7152);
nand U8369 (N_8369,N_6049,N_6065);
nand U8370 (N_8370,N_6012,N_7261);
nor U8371 (N_8371,N_6481,N_6464);
and U8372 (N_8372,N_6594,N_7033);
or U8373 (N_8373,N_7000,N_6522);
and U8374 (N_8374,N_6656,N_6857);
xnor U8375 (N_8375,N_6084,N_6171);
nand U8376 (N_8376,N_7065,N_7451);
nand U8377 (N_8377,N_6558,N_7017);
xnor U8378 (N_8378,N_7160,N_6564);
xor U8379 (N_8379,N_7033,N_6751);
nand U8380 (N_8380,N_6788,N_6990);
xnor U8381 (N_8381,N_6634,N_7308);
nor U8382 (N_8382,N_7283,N_6390);
nor U8383 (N_8383,N_6971,N_6681);
nand U8384 (N_8384,N_6672,N_6020);
nand U8385 (N_8385,N_6822,N_7081);
and U8386 (N_8386,N_7144,N_7079);
and U8387 (N_8387,N_7212,N_7405);
xnor U8388 (N_8388,N_7193,N_6851);
nor U8389 (N_8389,N_6759,N_7345);
nand U8390 (N_8390,N_6303,N_6487);
xor U8391 (N_8391,N_6137,N_6059);
nand U8392 (N_8392,N_7027,N_6429);
and U8393 (N_8393,N_6409,N_7219);
and U8394 (N_8394,N_7326,N_6187);
nor U8395 (N_8395,N_7451,N_6378);
nand U8396 (N_8396,N_7086,N_6504);
and U8397 (N_8397,N_6757,N_6377);
xnor U8398 (N_8398,N_7182,N_6822);
nand U8399 (N_8399,N_6832,N_7039);
nor U8400 (N_8400,N_6949,N_6761);
nor U8401 (N_8401,N_6667,N_7221);
nand U8402 (N_8402,N_6102,N_6886);
xnor U8403 (N_8403,N_7365,N_6277);
xor U8404 (N_8404,N_6388,N_6949);
nand U8405 (N_8405,N_6359,N_7254);
xor U8406 (N_8406,N_7115,N_6291);
xor U8407 (N_8407,N_6225,N_6070);
nand U8408 (N_8408,N_6976,N_7084);
xor U8409 (N_8409,N_6278,N_6644);
or U8410 (N_8410,N_6235,N_6781);
or U8411 (N_8411,N_6528,N_6837);
and U8412 (N_8412,N_6456,N_6489);
nand U8413 (N_8413,N_7273,N_6083);
and U8414 (N_8414,N_6521,N_6601);
and U8415 (N_8415,N_7248,N_6387);
or U8416 (N_8416,N_6270,N_7298);
nor U8417 (N_8417,N_6426,N_6199);
xnor U8418 (N_8418,N_6138,N_7150);
or U8419 (N_8419,N_6713,N_6715);
and U8420 (N_8420,N_7375,N_6259);
or U8421 (N_8421,N_6760,N_7182);
nor U8422 (N_8422,N_6716,N_6283);
and U8423 (N_8423,N_6934,N_7167);
xor U8424 (N_8424,N_7115,N_6879);
nor U8425 (N_8425,N_6258,N_7295);
xor U8426 (N_8426,N_6486,N_6518);
nand U8427 (N_8427,N_6410,N_6840);
xor U8428 (N_8428,N_6579,N_6037);
nor U8429 (N_8429,N_6834,N_6296);
and U8430 (N_8430,N_7275,N_7227);
or U8431 (N_8431,N_6992,N_7003);
xor U8432 (N_8432,N_6853,N_7120);
or U8433 (N_8433,N_6936,N_7424);
and U8434 (N_8434,N_7157,N_6349);
nor U8435 (N_8435,N_6759,N_7204);
or U8436 (N_8436,N_7053,N_6126);
nor U8437 (N_8437,N_6796,N_6280);
xor U8438 (N_8438,N_6219,N_6039);
xnor U8439 (N_8439,N_6868,N_7359);
nor U8440 (N_8440,N_7091,N_6515);
xnor U8441 (N_8441,N_6018,N_6601);
nor U8442 (N_8442,N_6914,N_6289);
xor U8443 (N_8443,N_7078,N_7050);
nor U8444 (N_8444,N_6109,N_7459);
nand U8445 (N_8445,N_6592,N_6184);
nand U8446 (N_8446,N_6602,N_6772);
or U8447 (N_8447,N_7462,N_7038);
or U8448 (N_8448,N_6159,N_6444);
xnor U8449 (N_8449,N_7224,N_6163);
nand U8450 (N_8450,N_6606,N_7207);
nand U8451 (N_8451,N_6896,N_6804);
nand U8452 (N_8452,N_6813,N_6308);
and U8453 (N_8453,N_7464,N_7195);
xor U8454 (N_8454,N_6059,N_6363);
nand U8455 (N_8455,N_7350,N_6631);
xnor U8456 (N_8456,N_6935,N_6122);
nor U8457 (N_8457,N_7305,N_6826);
nor U8458 (N_8458,N_6873,N_7390);
xnor U8459 (N_8459,N_7363,N_7468);
xnor U8460 (N_8460,N_7148,N_6023);
nand U8461 (N_8461,N_6361,N_6121);
nor U8462 (N_8462,N_7453,N_6885);
nand U8463 (N_8463,N_6752,N_6078);
or U8464 (N_8464,N_6504,N_6867);
xnor U8465 (N_8465,N_6865,N_7180);
xnor U8466 (N_8466,N_7330,N_6367);
or U8467 (N_8467,N_6170,N_7284);
and U8468 (N_8468,N_6770,N_6774);
or U8469 (N_8469,N_6689,N_6330);
or U8470 (N_8470,N_6605,N_6397);
or U8471 (N_8471,N_6947,N_6629);
and U8472 (N_8472,N_6798,N_6751);
nor U8473 (N_8473,N_6276,N_6953);
and U8474 (N_8474,N_6582,N_7328);
xor U8475 (N_8475,N_6175,N_7200);
nand U8476 (N_8476,N_6041,N_7279);
and U8477 (N_8477,N_7308,N_6436);
and U8478 (N_8478,N_6307,N_6478);
and U8479 (N_8479,N_6746,N_7391);
xnor U8480 (N_8480,N_6606,N_7076);
nand U8481 (N_8481,N_6178,N_6077);
nand U8482 (N_8482,N_7415,N_6437);
or U8483 (N_8483,N_6083,N_6003);
and U8484 (N_8484,N_6162,N_7388);
nand U8485 (N_8485,N_7411,N_6910);
xor U8486 (N_8486,N_6901,N_7207);
nor U8487 (N_8487,N_6726,N_7244);
nor U8488 (N_8488,N_6636,N_6323);
nor U8489 (N_8489,N_6358,N_6277);
xor U8490 (N_8490,N_6571,N_6544);
xnor U8491 (N_8491,N_7074,N_6061);
nor U8492 (N_8492,N_7072,N_6019);
nand U8493 (N_8493,N_7206,N_6545);
nor U8494 (N_8494,N_7375,N_6594);
nor U8495 (N_8495,N_7434,N_7417);
xor U8496 (N_8496,N_7242,N_6659);
and U8497 (N_8497,N_7389,N_6559);
xnor U8498 (N_8498,N_6513,N_7173);
nand U8499 (N_8499,N_6625,N_6729);
and U8500 (N_8500,N_6001,N_6275);
xor U8501 (N_8501,N_7047,N_6579);
nand U8502 (N_8502,N_7294,N_7077);
or U8503 (N_8503,N_7085,N_7116);
xor U8504 (N_8504,N_6410,N_6405);
xor U8505 (N_8505,N_6592,N_6975);
nor U8506 (N_8506,N_7286,N_6563);
and U8507 (N_8507,N_7028,N_7132);
nand U8508 (N_8508,N_6023,N_6565);
nor U8509 (N_8509,N_7048,N_6777);
or U8510 (N_8510,N_6721,N_6187);
or U8511 (N_8511,N_6545,N_6652);
and U8512 (N_8512,N_7075,N_6280);
nor U8513 (N_8513,N_7261,N_6841);
and U8514 (N_8514,N_6805,N_6230);
nor U8515 (N_8515,N_6349,N_6242);
nor U8516 (N_8516,N_6500,N_7390);
xnor U8517 (N_8517,N_7000,N_7209);
nand U8518 (N_8518,N_6880,N_6527);
or U8519 (N_8519,N_6927,N_6902);
xor U8520 (N_8520,N_6500,N_7353);
nor U8521 (N_8521,N_6526,N_7047);
nand U8522 (N_8522,N_6845,N_7175);
nor U8523 (N_8523,N_6659,N_6628);
xnor U8524 (N_8524,N_7432,N_6307);
or U8525 (N_8525,N_7405,N_7417);
and U8526 (N_8526,N_6987,N_6323);
nor U8527 (N_8527,N_7364,N_6868);
xnor U8528 (N_8528,N_6990,N_6251);
or U8529 (N_8529,N_6192,N_7338);
or U8530 (N_8530,N_7392,N_7457);
and U8531 (N_8531,N_6552,N_6474);
xor U8532 (N_8532,N_6521,N_6842);
and U8533 (N_8533,N_7111,N_6719);
xnor U8534 (N_8534,N_6646,N_6959);
xor U8535 (N_8535,N_6890,N_6988);
nor U8536 (N_8536,N_7439,N_6457);
xor U8537 (N_8537,N_7104,N_6977);
xor U8538 (N_8538,N_6648,N_6750);
or U8539 (N_8539,N_6893,N_6457);
or U8540 (N_8540,N_6990,N_6069);
and U8541 (N_8541,N_7294,N_7013);
nor U8542 (N_8542,N_6442,N_6521);
or U8543 (N_8543,N_6265,N_7481);
xor U8544 (N_8544,N_7462,N_7040);
or U8545 (N_8545,N_6997,N_6370);
nor U8546 (N_8546,N_6904,N_7277);
nand U8547 (N_8547,N_6490,N_6784);
nand U8548 (N_8548,N_6734,N_7022);
nand U8549 (N_8549,N_7093,N_7486);
or U8550 (N_8550,N_7315,N_6651);
xor U8551 (N_8551,N_6138,N_6092);
xor U8552 (N_8552,N_6528,N_6331);
or U8553 (N_8553,N_6119,N_6132);
and U8554 (N_8554,N_6037,N_6797);
xor U8555 (N_8555,N_7095,N_6535);
nor U8556 (N_8556,N_7403,N_6480);
and U8557 (N_8557,N_6679,N_7345);
and U8558 (N_8558,N_6732,N_7422);
nor U8559 (N_8559,N_6200,N_6080);
or U8560 (N_8560,N_6647,N_6324);
xnor U8561 (N_8561,N_6548,N_6741);
and U8562 (N_8562,N_6705,N_6928);
and U8563 (N_8563,N_6015,N_6901);
xnor U8564 (N_8564,N_6412,N_6907);
or U8565 (N_8565,N_6585,N_6427);
nand U8566 (N_8566,N_7192,N_7315);
nor U8567 (N_8567,N_6671,N_7413);
nor U8568 (N_8568,N_6049,N_6040);
and U8569 (N_8569,N_6367,N_6480);
nand U8570 (N_8570,N_7025,N_6403);
and U8571 (N_8571,N_7317,N_6248);
and U8572 (N_8572,N_6399,N_6712);
and U8573 (N_8573,N_7435,N_6997);
and U8574 (N_8574,N_7095,N_6998);
or U8575 (N_8575,N_7044,N_6254);
nor U8576 (N_8576,N_6417,N_7488);
nand U8577 (N_8577,N_7379,N_6770);
nor U8578 (N_8578,N_7355,N_7108);
nor U8579 (N_8579,N_7189,N_7030);
and U8580 (N_8580,N_7215,N_7067);
xnor U8581 (N_8581,N_6124,N_6121);
xor U8582 (N_8582,N_6843,N_6077);
nand U8583 (N_8583,N_7406,N_6896);
and U8584 (N_8584,N_6930,N_7066);
nor U8585 (N_8585,N_6552,N_7346);
nor U8586 (N_8586,N_6100,N_6577);
nor U8587 (N_8587,N_6863,N_6708);
nand U8588 (N_8588,N_6309,N_7130);
and U8589 (N_8589,N_6061,N_6236);
or U8590 (N_8590,N_6111,N_6844);
or U8591 (N_8591,N_7109,N_7096);
nor U8592 (N_8592,N_6326,N_7207);
nor U8593 (N_8593,N_6838,N_7135);
nand U8594 (N_8594,N_6090,N_7259);
nor U8595 (N_8595,N_7416,N_6523);
nand U8596 (N_8596,N_6951,N_6406);
and U8597 (N_8597,N_6770,N_7286);
xor U8598 (N_8598,N_6752,N_6193);
nor U8599 (N_8599,N_7338,N_6419);
nand U8600 (N_8600,N_7476,N_6765);
or U8601 (N_8601,N_6768,N_6154);
xnor U8602 (N_8602,N_7415,N_6902);
nand U8603 (N_8603,N_7090,N_6554);
and U8604 (N_8604,N_7456,N_6289);
or U8605 (N_8605,N_7166,N_7276);
nor U8606 (N_8606,N_6627,N_6695);
nor U8607 (N_8607,N_7432,N_7426);
xor U8608 (N_8608,N_7302,N_6225);
nand U8609 (N_8609,N_6275,N_7292);
or U8610 (N_8610,N_7016,N_7332);
nand U8611 (N_8611,N_6875,N_6773);
and U8612 (N_8612,N_7186,N_7145);
or U8613 (N_8613,N_6872,N_7415);
nor U8614 (N_8614,N_7055,N_7476);
nor U8615 (N_8615,N_6224,N_7056);
or U8616 (N_8616,N_6144,N_6303);
or U8617 (N_8617,N_7363,N_7404);
and U8618 (N_8618,N_7466,N_6511);
nor U8619 (N_8619,N_6964,N_6670);
or U8620 (N_8620,N_6271,N_7104);
nand U8621 (N_8621,N_6822,N_6294);
and U8622 (N_8622,N_6501,N_7053);
nand U8623 (N_8623,N_6441,N_6522);
xor U8624 (N_8624,N_7066,N_6476);
xor U8625 (N_8625,N_7342,N_6041);
and U8626 (N_8626,N_6611,N_6422);
nor U8627 (N_8627,N_7131,N_6918);
nand U8628 (N_8628,N_7366,N_6548);
nand U8629 (N_8629,N_6931,N_7071);
nor U8630 (N_8630,N_7343,N_6566);
xor U8631 (N_8631,N_6967,N_7129);
or U8632 (N_8632,N_6041,N_6848);
nand U8633 (N_8633,N_6461,N_6167);
nor U8634 (N_8634,N_7165,N_6061);
xnor U8635 (N_8635,N_6980,N_6513);
xnor U8636 (N_8636,N_6797,N_6069);
and U8637 (N_8637,N_7345,N_7176);
and U8638 (N_8638,N_6632,N_6525);
or U8639 (N_8639,N_6664,N_6380);
xnor U8640 (N_8640,N_6504,N_7180);
xor U8641 (N_8641,N_7252,N_6918);
xnor U8642 (N_8642,N_7076,N_6937);
or U8643 (N_8643,N_7439,N_6611);
nor U8644 (N_8644,N_6655,N_6052);
nor U8645 (N_8645,N_6420,N_7351);
xnor U8646 (N_8646,N_7067,N_7453);
and U8647 (N_8647,N_6958,N_6377);
and U8648 (N_8648,N_6047,N_7401);
or U8649 (N_8649,N_6205,N_6317);
or U8650 (N_8650,N_6310,N_6786);
nand U8651 (N_8651,N_7499,N_6648);
or U8652 (N_8652,N_6071,N_6165);
xnor U8653 (N_8653,N_6256,N_7031);
nor U8654 (N_8654,N_6866,N_7465);
and U8655 (N_8655,N_6556,N_7202);
nor U8656 (N_8656,N_6262,N_6397);
or U8657 (N_8657,N_6405,N_6144);
nor U8658 (N_8658,N_7267,N_7015);
or U8659 (N_8659,N_7167,N_6627);
and U8660 (N_8660,N_6089,N_6492);
or U8661 (N_8661,N_7203,N_6987);
and U8662 (N_8662,N_7000,N_6645);
nor U8663 (N_8663,N_7265,N_7154);
nor U8664 (N_8664,N_7329,N_7193);
or U8665 (N_8665,N_6030,N_6626);
xnor U8666 (N_8666,N_7115,N_6598);
xor U8667 (N_8667,N_7258,N_6695);
nor U8668 (N_8668,N_7230,N_6362);
xnor U8669 (N_8669,N_6524,N_6760);
xnor U8670 (N_8670,N_7341,N_6526);
xnor U8671 (N_8671,N_6604,N_7158);
and U8672 (N_8672,N_6867,N_6706);
or U8673 (N_8673,N_6890,N_6035);
nor U8674 (N_8674,N_6819,N_6199);
nor U8675 (N_8675,N_7468,N_7207);
xnor U8676 (N_8676,N_7318,N_6145);
nor U8677 (N_8677,N_6116,N_6218);
xor U8678 (N_8678,N_6689,N_6448);
or U8679 (N_8679,N_6517,N_7149);
and U8680 (N_8680,N_6129,N_6806);
xor U8681 (N_8681,N_7122,N_6345);
and U8682 (N_8682,N_6025,N_6852);
xnor U8683 (N_8683,N_6139,N_6280);
or U8684 (N_8684,N_6470,N_7338);
nor U8685 (N_8685,N_6568,N_7496);
nand U8686 (N_8686,N_6525,N_6673);
and U8687 (N_8687,N_6000,N_7409);
nand U8688 (N_8688,N_6154,N_7059);
or U8689 (N_8689,N_7245,N_7474);
or U8690 (N_8690,N_6226,N_6643);
xor U8691 (N_8691,N_6490,N_6615);
and U8692 (N_8692,N_6593,N_6826);
or U8693 (N_8693,N_6116,N_7026);
nand U8694 (N_8694,N_6452,N_6413);
or U8695 (N_8695,N_7009,N_7487);
or U8696 (N_8696,N_6872,N_6995);
and U8697 (N_8697,N_7116,N_6702);
nor U8698 (N_8698,N_7314,N_7383);
or U8699 (N_8699,N_6300,N_6970);
nor U8700 (N_8700,N_6153,N_6516);
nand U8701 (N_8701,N_7405,N_7110);
or U8702 (N_8702,N_7430,N_6510);
nand U8703 (N_8703,N_6187,N_6592);
xnor U8704 (N_8704,N_7205,N_6096);
nor U8705 (N_8705,N_7412,N_6575);
nor U8706 (N_8706,N_7147,N_7252);
nor U8707 (N_8707,N_6633,N_6094);
and U8708 (N_8708,N_6668,N_6555);
and U8709 (N_8709,N_6410,N_6512);
or U8710 (N_8710,N_6616,N_6032);
or U8711 (N_8711,N_6421,N_6591);
nand U8712 (N_8712,N_6333,N_6594);
and U8713 (N_8713,N_6445,N_6848);
xnor U8714 (N_8714,N_7280,N_7441);
or U8715 (N_8715,N_6475,N_6889);
or U8716 (N_8716,N_7485,N_6139);
or U8717 (N_8717,N_6288,N_7049);
or U8718 (N_8718,N_6473,N_6591);
or U8719 (N_8719,N_6384,N_6617);
nor U8720 (N_8720,N_7116,N_7318);
xor U8721 (N_8721,N_6168,N_6270);
or U8722 (N_8722,N_7145,N_6365);
or U8723 (N_8723,N_7349,N_7165);
xor U8724 (N_8724,N_6206,N_6569);
xnor U8725 (N_8725,N_7451,N_6272);
or U8726 (N_8726,N_6473,N_7193);
or U8727 (N_8727,N_6610,N_7147);
nor U8728 (N_8728,N_6882,N_6982);
xnor U8729 (N_8729,N_6861,N_7331);
xor U8730 (N_8730,N_7298,N_6290);
and U8731 (N_8731,N_6799,N_6494);
nor U8732 (N_8732,N_7050,N_7055);
xnor U8733 (N_8733,N_7029,N_7301);
nand U8734 (N_8734,N_6273,N_6769);
xor U8735 (N_8735,N_7426,N_6753);
or U8736 (N_8736,N_7241,N_7030);
xor U8737 (N_8737,N_6710,N_6281);
nand U8738 (N_8738,N_7064,N_6913);
and U8739 (N_8739,N_6727,N_6648);
and U8740 (N_8740,N_7238,N_6220);
nor U8741 (N_8741,N_6849,N_6098);
or U8742 (N_8742,N_6367,N_6518);
nor U8743 (N_8743,N_6327,N_7235);
and U8744 (N_8744,N_6169,N_7251);
nand U8745 (N_8745,N_6199,N_7253);
nor U8746 (N_8746,N_6437,N_6800);
xor U8747 (N_8747,N_6885,N_7215);
nand U8748 (N_8748,N_7003,N_6854);
nor U8749 (N_8749,N_7299,N_6499);
nor U8750 (N_8750,N_6525,N_6213);
nor U8751 (N_8751,N_6469,N_6413);
or U8752 (N_8752,N_6716,N_6199);
nand U8753 (N_8753,N_6117,N_7458);
or U8754 (N_8754,N_7235,N_7389);
nor U8755 (N_8755,N_6274,N_7032);
xor U8756 (N_8756,N_6647,N_6061);
and U8757 (N_8757,N_6554,N_7092);
nand U8758 (N_8758,N_6242,N_6936);
nor U8759 (N_8759,N_6478,N_7292);
xor U8760 (N_8760,N_6398,N_7447);
and U8761 (N_8761,N_7068,N_6022);
nand U8762 (N_8762,N_6182,N_7406);
and U8763 (N_8763,N_7062,N_7377);
or U8764 (N_8764,N_6786,N_7450);
and U8765 (N_8765,N_6515,N_7157);
nor U8766 (N_8766,N_7194,N_7413);
or U8767 (N_8767,N_6311,N_6806);
or U8768 (N_8768,N_6153,N_6101);
nand U8769 (N_8769,N_7026,N_7076);
xor U8770 (N_8770,N_6700,N_6025);
nand U8771 (N_8771,N_6612,N_6226);
and U8772 (N_8772,N_7296,N_6853);
nor U8773 (N_8773,N_7083,N_7424);
and U8774 (N_8774,N_6850,N_6277);
and U8775 (N_8775,N_6830,N_6826);
and U8776 (N_8776,N_7218,N_7017);
and U8777 (N_8777,N_7364,N_7149);
xor U8778 (N_8778,N_6269,N_7302);
nor U8779 (N_8779,N_7153,N_7417);
nand U8780 (N_8780,N_7409,N_7128);
nor U8781 (N_8781,N_6161,N_6227);
nand U8782 (N_8782,N_6250,N_7206);
nor U8783 (N_8783,N_6096,N_7154);
xor U8784 (N_8784,N_7263,N_6413);
and U8785 (N_8785,N_6847,N_6065);
nand U8786 (N_8786,N_6797,N_7461);
or U8787 (N_8787,N_6029,N_6753);
nor U8788 (N_8788,N_6462,N_6721);
xnor U8789 (N_8789,N_7189,N_6003);
nand U8790 (N_8790,N_7129,N_7361);
nand U8791 (N_8791,N_6932,N_7484);
or U8792 (N_8792,N_6503,N_6971);
nor U8793 (N_8793,N_6322,N_6485);
or U8794 (N_8794,N_6490,N_7149);
xnor U8795 (N_8795,N_6272,N_6678);
nor U8796 (N_8796,N_7183,N_6915);
xnor U8797 (N_8797,N_6470,N_6071);
or U8798 (N_8798,N_7103,N_7183);
and U8799 (N_8799,N_6244,N_6842);
nand U8800 (N_8800,N_6922,N_6321);
nor U8801 (N_8801,N_6395,N_6051);
and U8802 (N_8802,N_6929,N_7261);
and U8803 (N_8803,N_6238,N_7166);
nor U8804 (N_8804,N_7409,N_6530);
nor U8805 (N_8805,N_7087,N_6373);
and U8806 (N_8806,N_6522,N_6902);
xnor U8807 (N_8807,N_7221,N_6500);
and U8808 (N_8808,N_7279,N_7048);
and U8809 (N_8809,N_6756,N_7318);
or U8810 (N_8810,N_6198,N_6190);
nor U8811 (N_8811,N_7127,N_6963);
xnor U8812 (N_8812,N_7167,N_6755);
and U8813 (N_8813,N_6869,N_7187);
nand U8814 (N_8814,N_7032,N_7060);
xor U8815 (N_8815,N_6671,N_6734);
nor U8816 (N_8816,N_7260,N_6221);
nand U8817 (N_8817,N_6450,N_6697);
xnor U8818 (N_8818,N_6745,N_6911);
nand U8819 (N_8819,N_6405,N_6968);
nor U8820 (N_8820,N_6138,N_6857);
or U8821 (N_8821,N_6065,N_7325);
nand U8822 (N_8822,N_6265,N_6817);
nor U8823 (N_8823,N_7313,N_7234);
and U8824 (N_8824,N_7359,N_6148);
and U8825 (N_8825,N_6486,N_7011);
nor U8826 (N_8826,N_6243,N_6163);
nand U8827 (N_8827,N_7482,N_6582);
xor U8828 (N_8828,N_7239,N_6999);
and U8829 (N_8829,N_7429,N_7132);
nand U8830 (N_8830,N_7385,N_6250);
nand U8831 (N_8831,N_6784,N_6889);
nand U8832 (N_8832,N_6967,N_6910);
or U8833 (N_8833,N_6623,N_7276);
or U8834 (N_8834,N_6865,N_7317);
nor U8835 (N_8835,N_6419,N_7413);
nor U8836 (N_8836,N_6814,N_7376);
nor U8837 (N_8837,N_6059,N_6691);
nand U8838 (N_8838,N_6088,N_6145);
or U8839 (N_8839,N_6411,N_6227);
nand U8840 (N_8840,N_6985,N_7157);
and U8841 (N_8841,N_7259,N_7157);
or U8842 (N_8842,N_7432,N_6634);
and U8843 (N_8843,N_6665,N_7457);
xnor U8844 (N_8844,N_7128,N_6875);
nand U8845 (N_8845,N_7497,N_7178);
xnor U8846 (N_8846,N_6156,N_7348);
nand U8847 (N_8847,N_6687,N_6079);
or U8848 (N_8848,N_6734,N_6906);
nor U8849 (N_8849,N_7238,N_6668);
nor U8850 (N_8850,N_7024,N_7312);
nor U8851 (N_8851,N_6730,N_6748);
xnor U8852 (N_8852,N_6796,N_6229);
and U8853 (N_8853,N_7328,N_6877);
nand U8854 (N_8854,N_7237,N_6569);
or U8855 (N_8855,N_6419,N_6109);
and U8856 (N_8856,N_6863,N_7472);
nor U8857 (N_8857,N_6509,N_6845);
nand U8858 (N_8858,N_6862,N_6134);
nand U8859 (N_8859,N_6631,N_7298);
nor U8860 (N_8860,N_6740,N_7263);
xor U8861 (N_8861,N_6124,N_7076);
and U8862 (N_8862,N_6076,N_7439);
and U8863 (N_8863,N_7486,N_6124);
and U8864 (N_8864,N_7277,N_6715);
xnor U8865 (N_8865,N_6699,N_7398);
nand U8866 (N_8866,N_7240,N_6711);
nor U8867 (N_8867,N_6542,N_6438);
nand U8868 (N_8868,N_7307,N_6279);
and U8869 (N_8869,N_6837,N_6635);
xnor U8870 (N_8870,N_6710,N_6164);
nand U8871 (N_8871,N_6643,N_7155);
and U8872 (N_8872,N_6280,N_7457);
or U8873 (N_8873,N_6118,N_7110);
xnor U8874 (N_8874,N_6806,N_6497);
nand U8875 (N_8875,N_6284,N_7327);
and U8876 (N_8876,N_7361,N_6297);
and U8877 (N_8877,N_6857,N_6940);
or U8878 (N_8878,N_6290,N_6469);
nand U8879 (N_8879,N_7085,N_6241);
and U8880 (N_8880,N_6260,N_6884);
nand U8881 (N_8881,N_6401,N_6001);
xor U8882 (N_8882,N_7125,N_6638);
nand U8883 (N_8883,N_6287,N_6567);
nor U8884 (N_8884,N_7034,N_7032);
or U8885 (N_8885,N_6576,N_6197);
and U8886 (N_8886,N_6609,N_6752);
or U8887 (N_8887,N_6972,N_7194);
nand U8888 (N_8888,N_7182,N_7228);
or U8889 (N_8889,N_7288,N_6523);
xor U8890 (N_8890,N_6792,N_6693);
and U8891 (N_8891,N_7459,N_6498);
xor U8892 (N_8892,N_6933,N_7435);
xnor U8893 (N_8893,N_6865,N_7176);
xnor U8894 (N_8894,N_7397,N_6821);
and U8895 (N_8895,N_6296,N_7380);
or U8896 (N_8896,N_7410,N_7295);
nand U8897 (N_8897,N_6820,N_6066);
xor U8898 (N_8898,N_6880,N_6249);
xor U8899 (N_8899,N_6533,N_6449);
and U8900 (N_8900,N_6525,N_6422);
nand U8901 (N_8901,N_7335,N_7278);
or U8902 (N_8902,N_7267,N_7325);
nand U8903 (N_8903,N_7021,N_7214);
and U8904 (N_8904,N_6643,N_6670);
nand U8905 (N_8905,N_6153,N_7061);
nor U8906 (N_8906,N_6222,N_6391);
or U8907 (N_8907,N_6219,N_6831);
nor U8908 (N_8908,N_6517,N_6019);
nor U8909 (N_8909,N_7464,N_6571);
xor U8910 (N_8910,N_7145,N_7138);
and U8911 (N_8911,N_6098,N_7402);
xor U8912 (N_8912,N_7239,N_7201);
xnor U8913 (N_8913,N_6635,N_6030);
nor U8914 (N_8914,N_7446,N_6089);
or U8915 (N_8915,N_6331,N_6178);
nand U8916 (N_8916,N_6646,N_6914);
and U8917 (N_8917,N_6424,N_6378);
nand U8918 (N_8918,N_6754,N_7413);
xor U8919 (N_8919,N_6815,N_6038);
or U8920 (N_8920,N_7368,N_6337);
nand U8921 (N_8921,N_7080,N_6712);
nor U8922 (N_8922,N_7202,N_6013);
or U8923 (N_8923,N_6899,N_7485);
or U8924 (N_8924,N_6976,N_6478);
or U8925 (N_8925,N_6508,N_6511);
nand U8926 (N_8926,N_6847,N_7050);
or U8927 (N_8927,N_6084,N_7207);
or U8928 (N_8928,N_6343,N_6371);
or U8929 (N_8929,N_6170,N_6158);
xnor U8930 (N_8930,N_6401,N_7341);
or U8931 (N_8931,N_6754,N_6698);
xor U8932 (N_8932,N_7448,N_6295);
nor U8933 (N_8933,N_6596,N_7467);
or U8934 (N_8934,N_7366,N_6212);
or U8935 (N_8935,N_7178,N_6679);
nand U8936 (N_8936,N_7100,N_6475);
nor U8937 (N_8937,N_7443,N_6276);
xor U8938 (N_8938,N_7380,N_6374);
nand U8939 (N_8939,N_7410,N_6664);
or U8940 (N_8940,N_6937,N_6932);
nand U8941 (N_8941,N_6448,N_6837);
nor U8942 (N_8942,N_6104,N_6677);
or U8943 (N_8943,N_6053,N_7341);
nor U8944 (N_8944,N_6282,N_6416);
nor U8945 (N_8945,N_7454,N_7091);
xor U8946 (N_8946,N_6942,N_6832);
and U8947 (N_8947,N_6464,N_7130);
xnor U8948 (N_8948,N_6487,N_6098);
or U8949 (N_8949,N_6987,N_6313);
or U8950 (N_8950,N_6574,N_7258);
nand U8951 (N_8951,N_7118,N_7119);
nor U8952 (N_8952,N_6583,N_6438);
xor U8953 (N_8953,N_6600,N_6072);
or U8954 (N_8954,N_6949,N_6981);
and U8955 (N_8955,N_7214,N_7432);
or U8956 (N_8956,N_6721,N_6264);
and U8957 (N_8957,N_7051,N_6904);
xnor U8958 (N_8958,N_6494,N_7034);
or U8959 (N_8959,N_6686,N_7302);
or U8960 (N_8960,N_6588,N_6956);
nor U8961 (N_8961,N_6164,N_6778);
nor U8962 (N_8962,N_6421,N_7145);
xor U8963 (N_8963,N_7327,N_6860);
xor U8964 (N_8964,N_6940,N_6328);
xor U8965 (N_8965,N_6407,N_6277);
xor U8966 (N_8966,N_6647,N_6296);
and U8967 (N_8967,N_6193,N_6679);
nand U8968 (N_8968,N_6092,N_6625);
nor U8969 (N_8969,N_7211,N_7038);
nand U8970 (N_8970,N_6708,N_6114);
xnor U8971 (N_8971,N_7021,N_6208);
nand U8972 (N_8972,N_6384,N_6240);
or U8973 (N_8973,N_7329,N_6972);
nor U8974 (N_8974,N_7444,N_6494);
nand U8975 (N_8975,N_6312,N_6454);
nor U8976 (N_8976,N_6193,N_6471);
xnor U8977 (N_8977,N_7249,N_6583);
nand U8978 (N_8978,N_6528,N_6775);
xor U8979 (N_8979,N_6724,N_7199);
nor U8980 (N_8980,N_7283,N_6123);
xnor U8981 (N_8981,N_6170,N_6293);
or U8982 (N_8982,N_7324,N_6183);
xnor U8983 (N_8983,N_6692,N_7207);
xnor U8984 (N_8984,N_6275,N_7061);
nand U8985 (N_8985,N_7189,N_7444);
nor U8986 (N_8986,N_6331,N_6075);
xor U8987 (N_8987,N_6857,N_6504);
nor U8988 (N_8988,N_7065,N_6399);
and U8989 (N_8989,N_6470,N_7191);
nor U8990 (N_8990,N_7065,N_6940);
nor U8991 (N_8991,N_6796,N_6302);
or U8992 (N_8992,N_7447,N_7015);
and U8993 (N_8993,N_7063,N_6851);
nand U8994 (N_8994,N_6540,N_7315);
nor U8995 (N_8995,N_6320,N_6246);
or U8996 (N_8996,N_7292,N_6969);
xor U8997 (N_8997,N_7401,N_7411);
or U8998 (N_8998,N_7026,N_6884);
and U8999 (N_8999,N_7453,N_6741);
nor U9000 (N_9000,N_7511,N_7649);
xor U9001 (N_9001,N_7739,N_8390);
or U9002 (N_9002,N_8149,N_7898);
xnor U9003 (N_9003,N_8179,N_7573);
and U9004 (N_9004,N_8858,N_7697);
xor U9005 (N_9005,N_8355,N_8927);
nor U9006 (N_9006,N_7987,N_7748);
xnor U9007 (N_9007,N_8679,N_8518);
or U9008 (N_9008,N_7607,N_7947);
nor U9009 (N_9009,N_8926,N_7976);
or U9010 (N_9010,N_7938,N_8134);
nand U9011 (N_9011,N_8370,N_8048);
nor U9012 (N_9012,N_7841,N_8563);
xor U9013 (N_9013,N_8972,N_8878);
nor U9014 (N_9014,N_8405,N_7879);
xor U9015 (N_9015,N_7978,N_8908);
nand U9016 (N_9016,N_8816,N_8107);
nand U9017 (N_9017,N_8553,N_7889);
or U9018 (N_9018,N_8730,N_7711);
xor U9019 (N_9019,N_8865,N_7811);
nor U9020 (N_9020,N_8766,N_8975);
nor U9021 (N_9021,N_7535,N_8546);
and U9022 (N_9022,N_7679,N_8812);
nor U9023 (N_9023,N_8308,N_7634);
xor U9024 (N_9024,N_8891,N_8254);
nor U9025 (N_9025,N_8354,N_8519);
and U9026 (N_9026,N_8960,N_8172);
nor U9027 (N_9027,N_7916,N_7720);
nor U9028 (N_9028,N_8080,N_7895);
and U9029 (N_9029,N_7771,N_8826);
xor U9030 (N_9030,N_8316,N_7866);
and U9031 (N_9031,N_8260,N_7543);
xor U9032 (N_9032,N_8430,N_8132);
or U9033 (N_9033,N_8871,N_8980);
and U9034 (N_9034,N_7981,N_8581);
and U9035 (N_9035,N_8702,N_7730);
xnor U9036 (N_9036,N_8846,N_8221);
nand U9037 (N_9037,N_8995,N_7865);
nor U9038 (N_9038,N_7683,N_7927);
nor U9039 (N_9039,N_8326,N_7997);
and U9040 (N_9040,N_8018,N_8177);
nand U9041 (N_9041,N_7501,N_8231);
xor U9042 (N_9042,N_8947,N_8763);
and U9043 (N_9043,N_8073,N_8005);
and U9044 (N_9044,N_7521,N_8218);
and U9045 (N_9045,N_8567,N_8450);
nor U9046 (N_9046,N_7819,N_7961);
or U9047 (N_9047,N_8038,N_8569);
nand U9048 (N_9048,N_7763,N_8304);
nand U9049 (N_9049,N_8590,N_8401);
and U9050 (N_9050,N_8717,N_8618);
nand U9051 (N_9051,N_8566,N_7738);
nand U9052 (N_9052,N_7877,N_7685);
nor U9053 (N_9053,N_8297,N_8209);
and U9054 (N_9054,N_8464,N_7958);
xnor U9055 (N_9055,N_7655,N_8731);
xor U9056 (N_9056,N_8406,N_7853);
nor U9057 (N_9057,N_8629,N_8537);
or U9058 (N_9058,N_8637,N_7876);
nor U9059 (N_9059,N_7658,N_7974);
or U9060 (N_9060,N_7552,N_8901);
or U9061 (N_9061,N_8822,N_8071);
and U9062 (N_9062,N_8914,N_7827);
or U9063 (N_9063,N_8930,N_8797);
xnor U9064 (N_9064,N_8351,N_7859);
or U9065 (N_9065,N_8420,N_7681);
nand U9066 (N_9066,N_8558,N_8002);
nor U9067 (N_9067,N_7572,N_8769);
and U9068 (N_9068,N_7537,N_8216);
or U9069 (N_9069,N_8950,N_8695);
and U9070 (N_9070,N_7509,N_8491);
xnor U9071 (N_9071,N_8051,N_8396);
and U9072 (N_9072,N_8873,N_8157);
or U9073 (N_9073,N_7656,N_7937);
nor U9074 (N_9074,N_8715,N_7903);
nand U9075 (N_9075,N_8727,N_8565);
and U9076 (N_9076,N_8530,N_8597);
or U9077 (N_9077,N_8916,N_8887);
nor U9078 (N_9078,N_8014,N_8800);
or U9079 (N_9079,N_7642,N_8900);
nand U9080 (N_9080,N_8793,N_7992);
nand U9081 (N_9081,N_7957,N_8965);
or U9082 (N_9082,N_7684,N_7709);
and U9083 (N_9083,N_7868,N_8076);
nand U9084 (N_9084,N_7792,N_8448);
nand U9085 (N_9085,N_7631,N_8986);
nand U9086 (N_9086,N_8659,N_8239);
or U9087 (N_9087,N_7527,N_7528);
nand U9088 (N_9088,N_8199,N_8761);
xor U9089 (N_9089,N_8647,N_8643);
nor U9090 (N_9090,N_8976,N_8755);
and U9091 (N_9091,N_8840,N_8295);
or U9092 (N_9092,N_7963,N_7670);
xor U9093 (N_9093,N_8009,N_8658);
and U9094 (N_9094,N_7773,N_8875);
nand U9095 (N_9095,N_8620,N_7694);
nand U9096 (N_9096,N_8831,N_8968);
and U9097 (N_9097,N_8582,N_8333);
xnor U9098 (N_9098,N_7904,N_8056);
xor U9099 (N_9099,N_7575,N_8286);
and U9100 (N_9100,N_8161,N_8952);
xnor U9101 (N_9101,N_8317,N_8140);
xnor U9102 (N_9102,N_7640,N_7675);
and U9103 (N_9103,N_8278,N_8290);
and U9104 (N_9104,N_8810,N_8625);
and U9105 (N_9105,N_7596,N_7836);
nor U9106 (N_9106,N_8890,N_7909);
nand U9107 (N_9107,N_8981,N_8455);
or U9108 (N_9108,N_8327,N_8245);
nand U9109 (N_9109,N_7969,N_7783);
xnor U9110 (N_9110,N_7614,N_7775);
nand U9111 (N_9111,N_8714,N_8735);
nand U9112 (N_9112,N_8380,N_8229);
xnor U9113 (N_9113,N_8501,N_8392);
nand U9114 (N_9114,N_8917,N_7691);
nand U9115 (N_9115,N_8446,N_8570);
xor U9116 (N_9116,N_8603,N_7822);
nor U9117 (N_9117,N_8441,N_7837);
and U9118 (N_9118,N_7885,N_8109);
nor U9119 (N_9119,N_8599,N_7673);
xnor U9120 (N_9120,N_8827,N_8824);
nand U9121 (N_9121,N_8361,N_8206);
or U9122 (N_9122,N_8021,N_7627);
and U9123 (N_9123,N_8589,N_7786);
nor U9124 (N_9124,N_7599,N_8269);
or U9125 (N_9125,N_7531,N_8374);
nor U9126 (N_9126,N_8527,N_8693);
nor U9127 (N_9127,N_8262,N_8024);
nor U9128 (N_9128,N_8288,N_8505);
and U9129 (N_9129,N_8811,N_7516);
or U9130 (N_9130,N_8306,N_7584);
nand U9131 (N_9131,N_8939,N_7547);
nor U9132 (N_9132,N_8749,N_7559);
and U9133 (N_9133,N_7831,N_8204);
xnor U9134 (N_9134,N_8468,N_8334);
nand U9135 (N_9135,N_8640,N_8750);
and U9136 (N_9136,N_7979,N_8435);
or U9137 (N_9137,N_7556,N_8608);
nor U9138 (N_9138,N_8895,N_7973);
nand U9139 (N_9139,N_8985,N_8862);
and U9140 (N_9140,N_8594,N_8884);
nor U9141 (N_9141,N_7776,N_8801);
nor U9142 (N_9142,N_8743,N_8185);
xnor U9143 (N_9143,N_8632,N_8232);
and U9144 (N_9144,N_8561,N_8915);
nor U9145 (N_9145,N_8495,N_8384);
xor U9146 (N_9146,N_8694,N_7849);
nor U9147 (N_9147,N_7870,N_8851);
nor U9148 (N_9148,N_8809,N_8772);
or U9149 (N_9149,N_8186,N_7812);
nand U9150 (N_9150,N_7581,N_8789);
and U9151 (N_9151,N_7561,N_8685);
nor U9152 (N_9152,N_8310,N_8634);
and U9153 (N_9153,N_8805,N_8686);
and U9154 (N_9154,N_7918,N_8487);
nand U9155 (N_9155,N_8961,N_7712);
nor U9156 (N_9156,N_7660,N_8258);
and U9157 (N_9157,N_7637,N_7619);
nor U9158 (N_9158,N_7566,N_7839);
and U9159 (N_9159,N_8322,N_7793);
and U9160 (N_9160,N_8174,N_7817);
or U9161 (N_9161,N_8711,N_7603);
xor U9162 (N_9162,N_8284,N_8166);
or U9163 (N_9163,N_8742,N_7980);
nor U9164 (N_9164,N_7678,N_8545);
xnor U9165 (N_9165,N_8087,N_7504);
and U9166 (N_9166,N_7648,N_8765);
nor U9167 (N_9167,N_8114,N_8825);
nand U9168 (N_9168,N_8378,N_8301);
or U9169 (N_9169,N_8841,N_7750);
or U9170 (N_9170,N_8549,N_8358);
or U9171 (N_9171,N_7624,N_8692);
nor U9172 (N_9172,N_7816,N_7695);
nor U9173 (N_9173,N_7884,N_8339);
and U9174 (N_9174,N_7540,N_8838);
nand U9175 (N_9175,N_8399,N_8320);
nor U9176 (N_9176,N_7514,N_8135);
xnor U9177 (N_9177,N_8243,N_8525);
nor U9178 (N_9178,N_8323,N_8662);
xor U9179 (N_9179,N_8959,N_8540);
nand U9180 (N_9180,N_7911,N_7565);
and U9181 (N_9181,N_7705,N_8194);
nand U9182 (N_9182,N_8543,N_8493);
nor U9183 (N_9183,N_8385,N_7990);
nand U9184 (N_9184,N_8906,N_7715);
or U9185 (N_9185,N_8195,N_8585);
or U9186 (N_9186,N_8515,N_7782);
and U9187 (N_9187,N_7882,N_8630);
nand U9188 (N_9188,N_8214,N_8661);
nor U9189 (N_9189,N_8207,N_7743);
and U9190 (N_9190,N_8723,N_7662);
nand U9191 (N_9191,N_7668,N_7864);
nand U9192 (N_9192,N_7784,N_8422);
nand U9193 (N_9193,N_8604,N_8188);
and U9194 (N_9194,N_7588,N_7688);
or U9195 (N_9195,N_8829,N_8780);
nor U9196 (N_9196,N_7828,N_8413);
xor U9197 (N_9197,N_8744,N_7731);
nand U9198 (N_9198,N_8270,N_8181);
or U9199 (N_9199,N_8854,N_8646);
and U9200 (N_9200,N_8303,N_8756);
nand U9201 (N_9201,N_8595,N_8432);
nand U9202 (N_9202,N_8069,N_8434);
and U9203 (N_9203,N_8237,N_8752);
or U9204 (N_9204,N_7671,N_8423);
nand U9205 (N_9205,N_7677,N_7805);
or U9206 (N_9206,N_8047,N_8803);
or U9207 (N_9207,N_8880,N_7570);
nand U9208 (N_9208,N_8760,N_8667);
xnor U9209 (N_9209,N_8918,N_7626);
or U9210 (N_9210,N_8870,N_8377);
and U9211 (N_9211,N_8781,N_8145);
nor U9212 (N_9212,N_7567,N_7534);
and U9213 (N_9213,N_8642,N_8097);
and U9214 (N_9214,N_7910,N_8654);
xor U9215 (N_9215,N_8408,N_7644);
xnor U9216 (N_9216,N_7861,N_7966);
nor U9217 (N_9217,N_8298,N_8050);
nor U9218 (N_9218,N_7753,N_8718);
nand U9219 (N_9219,N_8987,N_8032);
nor U9220 (N_9220,N_8799,N_8782);
and U9221 (N_9221,N_8777,N_7667);
nand U9222 (N_9222,N_7777,N_7574);
nor U9223 (N_9223,N_7506,N_8101);
xnor U9224 (N_9224,N_8510,N_8176);
nand U9225 (N_9225,N_7690,N_7999);
or U9226 (N_9226,N_8293,N_8342);
and U9227 (N_9227,N_8485,N_8256);
or U9228 (N_9228,N_8480,N_7700);
and U9229 (N_9229,N_8592,N_7718);
nand U9230 (N_9230,N_7800,N_8118);
nor U9231 (N_9231,N_7721,N_7878);
nor U9232 (N_9232,N_8808,N_8834);
nand U9233 (N_9233,N_8211,N_8224);
nand U9234 (N_9234,N_7794,N_8287);
xnor U9235 (N_9235,N_8967,N_8279);
or U9236 (N_9236,N_8559,N_7914);
nand U9237 (N_9237,N_7576,N_7647);
xor U9238 (N_9238,N_8294,N_8063);
and U9239 (N_9239,N_8283,N_8276);
xnor U9240 (N_9240,N_8746,N_8249);
xnor U9241 (N_9241,N_7965,N_8119);
xor U9242 (N_9242,N_8117,N_8191);
xnor U9243 (N_9243,N_7842,N_8657);
nor U9244 (N_9244,N_8285,N_8259);
or U9245 (N_9245,N_7716,N_8219);
and U9246 (N_9246,N_8412,N_8652);
xnor U9247 (N_9247,N_7915,N_8183);
nand U9248 (N_9248,N_8886,N_8261);
and U9249 (N_9249,N_7922,N_7809);
nand U9250 (N_9250,N_8645,N_8335);
xor U9251 (N_9251,N_8672,N_7850);
or U9252 (N_9252,N_8226,N_8321);
or U9253 (N_9253,N_8210,N_8669);
and U9254 (N_9254,N_8180,N_7845);
or U9255 (N_9255,N_8639,N_7995);
and U9256 (N_9256,N_7944,N_7558);
nand U9257 (N_9257,N_7867,N_8196);
and U9258 (N_9258,N_8273,N_8644);
xor U9259 (N_9259,N_7931,N_8470);
and U9260 (N_9260,N_7863,N_8150);
and U9261 (N_9261,N_8167,N_7757);
or U9262 (N_9262,N_8362,N_8504);
nand U9263 (N_9263,N_8990,N_7761);
or U9264 (N_9264,N_8302,N_8579);
or U9265 (N_9265,N_8612,N_8163);
nand U9266 (N_9266,N_8153,N_7893);
nor U9267 (N_9267,N_7900,N_7740);
and U9268 (N_9268,N_8500,N_8331);
xor U9269 (N_9269,N_8758,N_8542);
nand U9270 (N_9270,N_8820,N_7989);
and U9271 (N_9271,N_8458,N_8966);
xnor U9272 (N_9272,N_8792,N_7796);
and U9273 (N_9273,N_7577,N_8934);
xnor U9274 (N_9274,N_7956,N_8614);
xnor U9275 (N_9275,N_8475,N_7769);
xor U9276 (N_9276,N_8275,N_7830);
and U9277 (N_9277,N_8416,N_7682);
xor U9278 (N_9278,N_8709,N_7808);
nor U9279 (N_9279,N_8061,N_8757);
or U9280 (N_9280,N_7610,N_8085);
xnor U9281 (N_9281,N_7536,N_8409);
or U9282 (N_9282,N_8400,N_7546);
xor U9283 (N_9283,N_8187,N_8190);
nand U9284 (N_9284,N_8856,N_8978);
or U9285 (N_9285,N_8452,N_7797);
or U9286 (N_9286,N_7747,N_7650);
or U9287 (N_9287,N_8739,N_8607);
or U9288 (N_9288,N_7928,N_8786);
and U9289 (N_9289,N_8095,N_8318);
or U9290 (N_9290,N_8600,N_8555);
or U9291 (N_9291,N_7703,N_7874);
nor U9292 (N_9292,N_7829,N_7825);
or U9293 (N_9293,N_8837,N_8282);
or U9294 (N_9294,N_8876,N_8931);
or U9295 (N_9295,N_8712,N_7620);
and U9296 (N_9296,N_8424,N_7636);
or U9297 (N_9297,N_8359,N_8775);
or U9298 (N_9298,N_7563,N_8954);
and U9299 (N_9299,N_8668,N_8855);
nor U9300 (N_9300,N_7994,N_8690);
or U9301 (N_9301,N_8902,N_7781);
and U9302 (N_9302,N_8921,N_8911);
xnor U9303 (N_9303,N_7657,N_8689);
or U9304 (N_9304,N_8996,N_8120);
or U9305 (N_9305,N_7933,N_8957);
and U9306 (N_9306,N_8687,N_7512);
nand U9307 (N_9307,N_7926,N_8748);
or U9308 (N_9308,N_8688,N_8872);
or U9309 (N_9309,N_7526,N_8465);
or U9310 (N_9310,N_8200,N_8139);
xnor U9311 (N_9311,N_8473,N_8088);
nand U9312 (N_9312,N_8705,N_8116);
nor U9313 (N_9313,N_8235,N_8513);
or U9314 (N_9314,N_7666,N_8857);
or U9315 (N_9315,N_8098,N_7801);
and U9316 (N_9316,N_8007,N_8492);
nand U9317 (N_9317,N_8713,N_8853);
or U9318 (N_9318,N_8779,N_8090);
nor U9319 (N_9319,N_8049,N_7632);
xnor U9320 (N_9320,N_8881,N_8751);
nand U9321 (N_9321,N_7815,N_7701);
or U9322 (N_9322,N_8674,N_8057);
nor U9323 (N_9323,N_8832,N_8268);
and U9324 (N_9324,N_8460,N_8587);
nand U9325 (N_9325,N_8389,N_8263);
and U9326 (N_9326,N_7635,N_8729);
and U9327 (N_9327,N_7766,N_8238);
xor U9328 (N_9328,N_8576,N_8255);
and U9329 (N_9329,N_8813,N_8523);
xnor U9330 (N_9330,N_8305,N_8111);
nor U9331 (N_9331,N_7772,N_7606);
nand U9332 (N_9332,N_7846,N_8676);
xor U9333 (N_9333,N_8201,N_7665);
nand U9334 (N_9334,N_7959,N_7734);
xnor U9335 (N_9335,N_8535,N_8205);
or U9336 (N_9336,N_8830,N_8146);
nor U9337 (N_9337,N_8212,N_7948);
nand U9338 (N_9338,N_7719,N_7615);
and U9339 (N_9339,N_8814,N_8324);
xnor U9340 (N_9340,N_8806,N_8251);
or U9341 (N_9341,N_7618,N_8478);
xnor U9342 (N_9342,N_8598,N_8319);
nand U9343 (N_9343,N_8343,N_7600);
or U9344 (N_9344,N_8708,N_8538);
nor U9345 (N_9345,N_7545,N_8125);
nand U9346 (N_9346,N_8074,N_8591);
and U9347 (N_9347,N_7851,N_8184);
nand U9348 (N_9348,N_8337,N_7741);
nand U9349 (N_9349,N_7823,N_7951);
nand U9350 (N_9350,N_8850,N_7736);
nand U9351 (N_9351,N_8017,N_8223);
nor U9352 (N_9352,N_8175,N_7892);
nand U9353 (N_9353,N_8019,N_8747);
and U9354 (N_9354,N_8601,N_8866);
nand U9355 (N_9355,N_8113,N_8393);
xnor U9356 (N_9356,N_7722,N_8086);
and U9357 (N_9357,N_8796,N_8707);
xnor U9358 (N_9358,N_8022,N_8469);
xor U9359 (N_9359,N_8020,N_8681);
and U9360 (N_9360,N_8068,N_8722);
nand U9361 (N_9361,N_8999,N_8903);
xnor U9362 (N_9362,N_8889,N_8363);
nand U9363 (N_9363,N_8030,N_8764);
xor U9364 (N_9364,N_7977,N_8483);
and U9365 (N_9365,N_7806,N_8586);
nor U9366 (N_9366,N_8953,N_8008);
nand U9367 (N_9367,N_8557,N_8497);
nand U9368 (N_9368,N_8615,N_8964);
or U9369 (N_9369,N_8461,N_8828);
and U9370 (N_9370,N_7663,N_8015);
nand U9371 (N_9371,N_8536,N_8064);
nand U9372 (N_9372,N_8035,N_8474);
or U9373 (N_9373,N_7522,N_7686);
and U9374 (N_9374,N_8867,N_7770);
and U9375 (N_9375,N_8045,N_8158);
xor U9376 (N_9376,N_8445,N_8281);
and U9377 (N_9377,N_7983,N_7661);
xnor U9378 (N_9378,N_8457,N_8471);
and U9379 (N_9379,N_8171,N_8443);
nand U9380 (N_9380,N_8753,N_8577);
and U9381 (N_9381,N_8266,N_7713);
nand U9382 (N_9382,N_7824,N_7953);
and U9383 (N_9383,N_7945,N_7592);
xor U9384 (N_9384,N_7733,N_7896);
nor U9385 (N_9385,N_7840,N_7970);
xnor U9386 (N_9386,N_8197,N_8381);
or U9387 (N_9387,N_8128,N_7856);
and U9388 (N_9388,N_8054,N_7518);
and U9389 (N_9389,N_8041,N_7723);
nor U9390 (N_9390,N_8453,N_8108);
and U9391 (N_9391,N_8998,N_8202);
nor U9392 (N_9392,N_8033,N_8888);
or U9393 (N_9393,N_7706,N_8821);
nand U9394 (N_9394,N_8092,N_7891);
nor U9395 (N_9395,N_8861,N_7887);
nand U9396 (N_9396,N_7803,N_8250);
and U9397 (N_9397,N_8421,N_8271);
nor U9398 (N_9398,N_8449,N_8459);
and U9399 (N_9399,N_8058,N_7996);
nand U9400 (N_9400,N_8039,N_7548);
nand U9401 (N_9401,N_7569,N_8932);
or U9402 (N_9402,N_7590,N_8849);
and U9403 (N_9403,N_8622,N_8371);
nand U9404 (N_9404,N_8716,N_8904);
and U9405 (N_9405,N_7932,N_8230);
nand U9406 (N_9406,N_8949,N_8368);
and U9407 (N_9407,N_7943,N_8367);
xnor U9408 (N_9408,N_8564,N_8332);
nand U9409 (N_9409,N_7756,N_8697);
and U9410 (N_9410,N_8635,N_8913);
or U9411 (N_9411,N_8588,N_8403);
and U9412 (N_9412,N_8307,N_8127);
and U9413 (N_9413,N_7985,N_7550);
or U9414 (N_9414,N_8847,N_8943);
nor U9415 (N_9415,N_8842,N_8833);
nor U9416 (N_9416,N_7638,N_8706);
nor U9417 (N_9417,N_8733,N_8843);
xor U9418 (N_9418,N_7609,N_8394);
nor U9419 (N_9419,N_8539,N_8313);
nor U9420 (N_9420,N_7873,N_8664);
nor U9421 (N_9421,N_7855,N_7993);
xnor U9422 (N_9422,N_8144,N_7854);
nand U9423 (N_9423,N_8490,N_8454);
xnor U9424 (N_9424,N_8340,N_7586);
xnor U9425 (N_9425,N_8924,N_7710);
nand U9426 (N_9426,N_8920,N_8126);
and U9427 (N_9427,N_8839,N_8628);
or U9428 (N_9428,N_8971,N_7986);
and U9429 (N_9429,N_7826,N_8933);
and U9430 (N_9430,N_8192,N_8509);
and U9431 (N_9431,N_8883,N_7539);
and U9432 (N_9432,N_7871,N_8198);
or U9433 (N_9433,N_7833,N_7551);
and U9434 (N_9434,N_7982,N_7848);
nor U9435 (N_9435,N_8240,N_7758);
nor U9436 (N_9436,N_8438,N_7964);
xor U9437 (N_9437,N_8962,N_8675);
or U9438 (N_9438,N_8350,N_8511);
nand U9439 (N_9439,N_7962,N_8000);
nand U9440 (N_9440,N_7862,N_7802);
xor U9441 (N_9441,N_8869,N_8466);
nand U9442 (N_9442,N_8141,N_8574);
xnor U9443 (N_9443,N_8072,N_8548);
xor U9444 (N_9444,N_7901,N_8155);
xnor U9445 (N_9445,N_8152,N_8521);
nor U9446 (N_9446,N_8512,N_8698);
nor U9447 (N_9447,N_8143,N_8330);
or U9448 (N_9448,N_7894,N_7813);
and U9449 (N_9449,N_7704,N_8463);
and U9450 (N_9450,N_8696,N_8514);
nand U9451 (N_9451,N_8958,N_8103);
nor U9452 (N_9452,N_7768,N_8060);
xnor U9453 (N_9453,N_7519,N_7939);
or U9454 (N_9454,N_7905,N_7639);
or U9455 (N_9455,N_8344,N_8044);
and U9456 (N_9456,N_8070,N_7886);
nor U9457 (N_9457,N_8462,N_8554);
nor U9458 (N_9458,N_8955,N_8624);
nand U9459 (N_9459,N_8583,N_8345);
nand U9460 (N_9460,N_8426,N_8787);
nor U9461 (N_9461,N_8383,N_7544);
and U9462 (N_9462,N_8397,N_7787);
xnor U9463 (N_9463,N_7968,N_7680);
and U9464 (N_9464,N_7858,N_7617);
nand U9465 (N_9465,N_8874,N_7594);
nor U9466 (N_9466,N_8724,N_7625);
and U9467 (N_9467,N_8252,N_7595);
and U9468 (N_9468,N_8164,N_7669);
nand U9469 (N_9469,N_7717,N_8124);
and U9470 (N_9470,N_8165,N_7643);
xnor U9471 (N_9471,N_7532,N_8447);
nand U9472 (N_9472,N_8738,N_8894);
and U9473 (N_9473,N_8376,N_8817);
nor U9474 (N_9474,N_8879,N_7517);
and U9475 (N_9475,N_8928,N_7912);
nor U9476 (N_9476,N_8402,N_8885);
or U9477 (N_9477,N_7674,N_8028);
xnor U9478 (N_9478,N_8770,N_8541);
nor U9479 (N_9479,N_7897,N_7920);
xnor U9480 (N_9480,N_8488,N_7696);
xor U9481 (N_9481,N_8524,N_8479);
xor U9482 (N_9482,N_8759,N_8925);
and U9483 (N_9483,N_7538,N_7560);
nand U9484 (N_9484,N_8673,N_7835);
xor U9485 (N_9485,N_7754,N_8573);
or U9486 (N_9486,N_8062,N_7742);
or U9487 (N_9487,N_7799,N_7875);
and U9488 (N_9488,N_8671,N_8993);
xor U9489 (N_9489,N_7923,N_7908);
xor U9490 (N_9490,N_8100,N_8067);
nor U9491 (N_9491,N_8228,N_8531);
and U9492 (N_9492,N_8868,N_8936);
nor U9493 (N_9493,N_8774,N_8234);
nand U9494 (N_9494,N_8666,N_8575);
nor U9495 (N_9495,N_8942,N_8027);
nand U9496 (N_9496,N_7525,N_7707);
and U9497 (N_9497,N_7557,N_8220);
and U9498 (N_9498,N_8771,N_8043);
nor U9499 (N_9499,N_8649,N_8300);
nand U9500 (N_9500,N_8807,N_8528);
or U9501 (N_9501,N_8336,N_7542);
nand U9502 (N_9502,N_8776,N_8055);
and U9503 (N_9503,N_8507,N_8677);
nand U9504 (N_9504,N_8636,N_8026);
nand U9505 (N_9505,N_8631,N_8083);
nor U9506 (N_9506,N_8802,N_8762);
nand U9507 (N_9507,N_8233,N_7689);
or U9508 (N_9508,N_8929,N_8701);
or U9509 (N_9509,N_8948,N_8836);
or U9510 (N_9510,N_8526,N_8105);
or U9511 (N_9511,N_7533,N_8225);
nor U9512 (N_9512,N_8012,N_8241);
nand U9513 (N_9513,N_8905,N_8042);
or U9514 (N_9514,N_7745,N_7724);
nand U9515 (N_9515,N_7751,N_8935);
and U9516 (N_9516,N_8414,N_7737);
xor U9517 (N_9517,N_7633,N_8123);
or U9518 (N_9518,N_7984,N_8973);
xor U9519 (N_9519,N_8946,N_7578);
or U9520 (N_9520,N_8481,N_7628);
xor U9521 (N_9521,N_8503,N_8859);
and U9522 (N_9522,N_8977,N_8439);
nor U9523 (N_9523,N_7820,N_8571);
or U9524 (N_9524,N_8348,N_8138);
or U9525 (N_9525,N_8940,N_8919);
xor U9526 (N_9526,N_8277,N_8265);
xor U9527 (N_9527,N_8721,N_7530);
and U9528 (N_9528,N_8023,N_8272);
nand U9529 (N_9529,N_8616,N_7692);
and U9530 (N_9530,N_8997,N_8467);
nand U9531 (N_9531,N_8863,N_8506);
nor U9532 (N_9532,N_7975,N_8398);
nor U9533 (N_9533,N_8395,N_8845);
or U9534 (N_9534,N_7752,N_8626);
xor U9535 (N_9535,N_7843,N_8352);
or U9536 (N_9536,N_8096,N_8819);
and U9537 (N_9537,N_8795,N_8115);
and U9538 (N_9538,N_7579,N_7929);
nor U9539 (N_9539,N_7698,N_8078);
nand U9540 (N_9540,N_7608,N_8684);
or U9541 (N_9541,N_8922,N_8791);
nand U9542 (N_9542,N_8937,N_7708);
or U9543 (N_9543,N_8079,N_8325);
nand U9544 (N_9544,N_8016,N_7729);
nand U9545 (N_9545,N_7946,N_7529);
nand U9546 (N_9546,N_7759,N_8522);
or U9547 (N_9547,N_7907,N_8773);
nand U9548 (N_9548,N_7834,N_8292);
xor U9549 (N_9549,N_8754,N_7764);
nor U9550 (N_9550,N_8349,N_8989);
nand U9551 (N_9551,N_7622,N_8444);
xor U9552 (N_9552,N_8720,N_8623);
and U9553 (N_9553,N_8882,N_7587);
xnor U9554 (N_9554,N_8683,N_8941);
nand U9555 (N_9555,N_7934,N_8663);
nor U9556 (N_9556,N_7591,N_8788);
nand U9557 (N_9557,N_8142,N_7941);
nor U9558 (N_9558,N_8703,N_8160);
nor U9559 (N_9559,N_8898,N_7583);
nor U9560 (N_9560,N_7503,N_8477);
nand U9561 (N_9561,N_7844,N_8341);
xor U9562 (N_9562,N_8173,N_7919);
xnor U9563 (N_9563,N_7888,N_8670);
xor U9564 (N_9564,N_8499,N_8893);
and U9565 (N_9565,N_7693,N_8338);
nor U9566 (N_9566,N_7883,N_7925);
nand U9567 (N_9567,N_7621,N_7510);
xor U9568 (N_9568,N_8433,N_8372);
and U9569 (N_9569,N_8373,N_8011);
xor U9570 (N_9570,N_7629,N_8619);
nand U9571 (N_9571,N_8208,N_8094);
nor U9572 (N_9572,N_8159,N_8852);
nor U9573 (N_9573,N_8311,N_8992);
nor U9574 (N_9574,N_8248,N_7899);
xor U9575 (N_9575,N_8605,N_7972);
xor U9576 (N_9576,N_8168,N_8036);
or U9577 (N_9577,N_8328,N_8899);
nand U9578 (N_9578,N_7791,N_8728);
nor U9579 (N_9579,N_7902,N_7880);
and U9580 (N_9580,N_8736,N_7623);
or U9581 (N_9581,N_8299,N_8162);
xnor U9582 (N_9582,N_7935,N_8296);
nand U9583 (N_9583,N_7950,N_8081);
xor U9584 (N_9584,N_7804,N_8641);
xor U9585 (N_9585,N_7988,N_8029);
and U9586 (N_9586,N_8602,N_8844);
nand U9587 (N_9587,N_8486,N_8147);
nand U9588 (N_9588,N_8482,N_7760);
nand U9589 (N_9589,N_8429,N_8745);
and U9590 (N_9590,N_8665,N_8596);
xnor U9591 (N_9591,N_8082,N_7554);
or U9592 (N_9592,N_7832,N_8215);
or U9593 (N_9593,N_8387,N_7582);
or U9594 (N_9594,N_8236,N_7857);
nor U9595 (N_9595,N_8923,N_7818);
or U9596 (N_9596,N_8737,N_8442);
or U9597 (N_9597,N_8785,N_8551);
or U9598 (N_9598,N_8835,N_8909);
nand U9599 (N_9599,N_8544,N_7762);
and U9600 (N_9600,N_8077,N_7676);
xnor U9601 (N_9601,N_8741,N_8956);
and U9602 (N_9602,N_8609,N_8451);
nand U9603 (N_9603,N_8419,N_7780);
nor U9604 (N_9604,N_7651,N_7645);
nand U9605 (N_9605,N_8193,N_8534);
nand U9606 (N_9606,N_8508,N_7714);
nand U9607 (N_9607,N_7604,N_8106);
nor U9608 (N_9608,N_8312,N_8386);
nor U9609 (N_9609,N_8133,N_8650);
nor U9610 (N_9610,N_8734,N_7971);
nand U9611 (N_9611,N_8991,N_8818);
xor U9612 (N_9612,N_8314,N_8003);
nor U9613 (N_9613,N_8578,N_7872);
nor U9614 (N_9614,N_8938,N_7702);
nand U9615 (N_9615,N_7921,N_8365);
xnor U9616 (N_9616,N_8375,N_8267);
nor U9617 (N_9617,N_8004,N_8994);
nand U9618 (N_9618,N_8031,N_8170);
xor U9619 (N_9619,N_8912,N_8053);
nand U9620 (N_9620,N_8346,N_7630);
xor U9621 (N_9621,N_8790,N_8617);
nor U9622 (N_9622,N_7541,N_8691);
nor U9623 (N_9623,N_7821,N_8732);
and U9624 (N_9624,N_8892,N_8651);
and U9625 (N_9625,N_7611,N_8982);
nor U9626 (N_9626,N_8489,N_8415);
or U9627 (N_9627,N_7798,N_8472);
or U9628 (N_9628,N_8529,N_7940);
or U9629 (N_9629,N_7659,N_8476);
xnor U9630 (N_9630,N_8169,N_7520);
or U9631 (N_9631,N_7788,N_8006);
nand U9632 (N_9632,N_7807,N_8648);
nor U9633 (N_9633,N_8110,N_7641);
nor U9634 (N_9634,N_8227,N_8606);
nand U9635 (N_9635,N_8794,N_8502);
or U9636 (N_9636,N_8156,N_7502);
xor U9637 (N_9637,N_8700,N_8610);
xor U9638 (N_9638,N_8963,N_8010);
nand U9639 (N_9639,N_8678,N_8264);
and U9640 (N_9640,N_7699,N_7616);
nand U9641 (N_9641,N_8593,N_8613);
xor U9642 (N_9642,N_8066,N_8257);
and U9643 (N_9643,N_7814,N_7913);
or U9644 (N_9644,N_8075,N_8768);
or U9645 (N_9645,N_8550,N_8568);
nand U9646 (N_9646,N_7653,N_7942);
or U9647 (N_9647,N_8633,N_8726);
nor U9648 (N_9648,N_8222,N_8130);
nand U9649 (N_9649,N_8065,N_8494);
and U9650 (N_9650,N_8740,N_8516);
nor U9651 (N_9651,N_8089,N_8112);
nor U9652 (N_9652,N_8001,N_8203);
nand U9653 (N_9653,N_8046,N_7917);
nor U9654 (N_9654,N_7513,N_7597);
nor U9655 (N_9655,N_7767,N_8517);
nor U9656 (N_9656,N_8877,N_8391);
xnor U9657 (N_9657,N_8428,N_7553);
xnor U9658 (N_9658,N_8572,N_8860);
xor U9659 (N_9659,N_7906,N_8660);
nand U9660 (N_9660,N_8407,N_8556);
nor U9661 (N_9661,N_7589,N_7991);
nor U9662 (N_9662,N_8154,N_8823);
nand U9663 (N_9663,N_8347,N_8246);
nand U9664 (N_9664,N_7652,N_7778);
xor U9665 (N_9665,N_8725,N_8767);
or U9666 (N_9666,N_8710,N_8848);
nor U9667 (N_9667,N_8784,N_8136);
or U9668 (N_9668,N_7555,N_8456);
nor U9669 (N_9669,N_7869,N_8182);
xnor U9670 (N_9670,N_8437,N_7727);
or U9671 (N_9671,N_8034,N_8052);
nor U9672 (N_9672,N_7613,N_7795);
nor U9673 (N_9673,N_8896,N_8411);
nand U9674 (N_9674,N_7605,N_8621);
nor U9675 (N_9675,N_8983,N_8356);
nand U9676 (N_9676,N_8244,N_8353);
and U9677 (N_9677,N_8360,N_8309);
or U9678 (N_9678,N_7664,N_8151);
nand U9679 (N_9679,N_8484,N_8366);
nor U9680 (N_9680,N_7507,N_8611);
xnor U9681 (N_9681,N_7598,N_7746);
or U9682 (N_9682,N_8804,N_7728);
and U9683 (N_9683,N_7726,N_8242);
nor U9684 (N_9684,N_8783,N_7508);
nor U9685 (N_9685,N_7646,N_7955);
or U9686 (N_9686,N_8013,N_8025);
nand U9687 (N_9687,N_8655,N_7954);
or U9688 (N_9688,N_8974,N_8580);
nand U9689 (N_9689,N_8533,N_7735);
nand U9690 (N_9690,N_8404,N_7785);
or U9691 (N_9691,N_7930,N_8638);
or U9692 (N_9692,N_7860,N_7765);
nand U9693 (N_9693,N_8656,N_8410);
and U9694 (N_9694,N_8369,N_8148);
or U9695 (N_9695,N_7500,N_7687);
and U9696 (N_9696,N_7838,N_8418);
nor U9697 (N_9697,N_8121,N_8137);
or U9698 (N_9698,N_7998,N_7779);
nand U9699 (N_9699,N_7725,N_8274);
and U9700 (N_9700,N_7890,N_7960);
or U9701 (N_9701,N_8864,N_8969);
and U9702 (N_9702,N_7790,N_8584);
xnor U9703 (N_9703,N_7924,N_7732);
nor U9704 (N_9704,N_7571,N_7949);
nand U9705 (N_9705,N_8436,N_8379);
nor U9706 (N_9706,N_8357,N_8547);
xnor U9707 (N_9707,N_8907,N_7585);
xor U9708 (N_9708,N_8440,N_8280);
nor U9709 (N_9709,N_7523,N_7602);
nor U9710 (N_9710,N_8037,N_8560);
and U9711 (N_9711,N_8552,N_8178);
nor U9712 (N_9712,N_8122,N_8093);
nand U9713 (N_9713,N_8291,N_7755);
and U9714 (N_9714,N_8719,N_8253);
and U9715 (N_9715,N_7672,N_7505);
nand U9716 (N_9716,N_8417,N_8498);
and U9717 (N_9717,N_8988,N_8364);
xnor U9718 (N_9718,N_7936,N_8562);
nor U9719 (N_9719,N_8329,N_8798);
nor U9720 (N_9720,N_7593,N_8680);
xnor U9721 (N_9721,N_8315,N_7568);
nor U9722 (N_9722,N_7601,N_7749);
nand U9723 (N_9723,N_8289,N_7952);
and U9724 (N_9724,N_7580,N_8979);
nor U9725 (N_9725,N_7774,N_7881);
and U9726 (N_9726,N_7515,N_7564);
or U9727 (N_9727,N_8084,N_8388);
nand U9728 (N_9728,N_7967,N_8217);
or U9729 (N_9729,N_8627,N_8425);
nor U9730 (N_9730,N_8102,N_7612);
or U9731 (N_9731,N_8104,N_7562);
and U9732 (N_9732,N_8189,N_8247);
and U9733 (N_9733,N_8091,N_8213);
nor U9734 (N_9734,N_7524,N_8945);
xnor U9735 (N_9735,N_7852,N_8778);
xor U9736 (N_9736,N_8040,N_8520);
and U9737 (N_9737,N_7789,N_8951);
nand U9738 (N_9738,N_8815,N_7744);
xor U9739 (N_9739,N_8129,N_8970);
nand U9740 (N_9740,N_8059,N_7847);
xnor U9741 (N_9741,N_8099,N_8431);
and U9742 (N_9742,N_8653,N_7654);
nor U9743 (N_9743,N_7549,N_7810);
xnor U9744 (N_9744,N_8496,N_8944);
and U9745 (N_9745,N_8699,N_8427);
xnor U9746 (N_9746,N_8382,N_8532);
or U9747 (N_9747,N_8704,N_8984);
and U9748 (N_9748,N_8910,N_8682);
or U9749 (N_9749,N_8131,N_8897);
or U9750 (N_9750,N_8607,N_8110);
nor U9751 (N_9751,N_7635,N_8843);
nor U9752 (N_9752,N_7762,N_7618);
nand U9753 (N_9753,N_7888,N_8306);
or U9754 (N_9754,N_8604,N_8814);
and U9755 (N_9755,N_8317,N_8536);
or U9756 (N_9756,N_8728,N_7940);
xor U9757 (N_9757,N_7623,N_8576);
nand U9758 (N_9758,N_8109,N_8299);
and U9759 (N_9759,N_8511,N_7872);
or U9760 (N_9760,N_8737,N_8500);
nand U9761 (N_9761,N_8311,N_8538);
nand U9762 (N_9762,N_8635,N_8374);
and U9763 (N_9763,N_8027,N_8040);
nor U9764 (N_9764,N_8200,N_7648);
xor U9765 (N_9765,N_8898,N_8608);
and U9766 (N_9766,N_7707,N_8259);
xor U9767 (N_9767,N_8580,N_8489);
and U9768 (N_9768,N_8707,N_8056);
nand U9769 (N_9769,N_8482,N_8727);
xor U9770 (N_9770,N_8181,N_8806);
nand U9771 (N_9771,N_8773,N_7664);
and U9772 (N_9772,N_7547,N_8966);
nor U9773 (N_9773,N_8587,N_7955);
nor U9774 (N_9774,N_7782,N_7883);
nand U9775 (N_9775,N_8128,N_8567);
xnor U9776 (N_9776,N_7882,N_7828);
and U9777 (N_9777,N_7669,N_7685);
and U9778 (N_9778,N_7952,N_8190);
or U9779 (N_9779,N_8333,N_8802);
or U9780 (N_9780,N_7742,N_8665);
nor U9781 (N_9781,N_8226,N_7932);
or U9782 (N_9782,N_7629,N_7680);
xor U9783 (N_9783,N_8855,N_8734);
xor U9784 (N_9784,N_8193,N_7850);
or U9785 (N_9785,N_8251,N_7599);
nand U9786 (N_9786,N_8134,N_8731);
or U9787 (N_9787,N_7507,N_7733);
nand U9788 (N_9788,N_8635,N_7719);
nand U9789 (N_9789,N_8428,N_7636);
and U9790 (N_9790,N_8022,N_8389);
nor U9791 (N_9791,N_7539,N_8669);
nor U9792 (N_9792,N_8957,N_8309);
xor U9793 (N_9793,N_8221,N_8137);
and U9794 (N_9794,N_8948,N_7918);
and U9795 (N_9795,N_7795,N_7625);
or U9796 (N_9796,N_8670,N_8248);
and U9797 (N_9797,N_8543,N_8443);
nor U9798 (N_9798,N_8400,N_7588);
nor U9799 (N_9799,N_7876,N_7971);
or U9800 (N_9800,N_8235,N_8453);
or U9801 (N_9801,N_8442,N_8997);
or U9802 (N_9802,N_8542,N_8574);
and U9803 (N_9803,N_8784,N_7960);
nor U9804 (N_9804,N_8825,N_8022);
nand U9805 (N_9805,N_8003,N_8702);
nor U9806 (N_9806,N_7863,N_8122);
xor U9807 (N_9807,N_8767,N_8220);
nor U9808 (N_9808,N_8235,N_8783);
or U9809 (N_9809,N_8446,N_8387);
nor U9810 (N_9810,N_8271,N_8326);
nor U9811 (N_9811,N_7775,N_8389);
or U9812 (N_9812,N_8478,N_8838);
xnor U9813 (N_9813,N_8276,N_7555);
nor U9814 (N_9814,N_8002,N_8175);
nand U9815 (N_9815,N_8953,N_8449);
nand U9816 (N_9816,N_7938,N_8441);
nor U9817 (N_9817,N_8838,N_7936);
xor U9818 (N_9818,N_8407,N_8373);
nand U9819 (N_9819,N_7683,N_8132);
and U9820 (N_9820,N_7749,N_8444);
nor U9821 (N_9821,N_8643,N_8451);
or U9822 (N_9822,N_8377,N_8299);
xor U9823 (N_9823,N_8275,N_7906);
xor U9824 (N_9824,N_7633,N_7851);
nand U9825 (N_9825,N_7721,N_8460);
nand U9826 (N_9826,N_8123,N_8186);
nand U9827 (N_9827,N_7749,N_7666);
nand U9828 (N_9828,N_8055,N_8116);
and U9829 (N_9829,N_8316,N_8463);
xnor U9830 (N_9830,N_7994,N_8260);
xor U9831 (N_9831,N_8406,N_8588);
nor U9832 (N_9832,N_7511,N_7824);
or U9833 (N_9833,N_8041,N_8118);
nand U9834 (N_9834,N_8850,N_8551);
xor U9835 (N_9835,N_7769,N_8784);
and U9836 (N_9836,N_8594,N_7882);
nand U9837 (N_9837,N_8780,N_8873);
or U9838 (N_9838,N_7532,N_7606);
or U9839 (N_9839,N_8989,N_8756);
and U9840 (N_9840,N_7921,N_8612);
xnor U9841 (N_9841,N_7845,N_8192);
nand U9842 (N_9842,N_7679,N_8433);
and U9843 (N_9843,N_8117,N_7755);
nand U9844 (N_9844,N_8570,N_8444);
xor U9845 (N_9845,N_8036,N_7579);
nand U9846 (N_9846,N_8060,N_8453);
and U9847 (N_9847,N_8668,N_7888);
and U9848 (N_9848,N_7692,N_7521);
or U9849 (N_9849,N_7603,N_8493);
nor U9850 (N_9850,N_8320,N_7795);
xor U9851 (N_9851,N_7526,N_8161);
nor U9852 (N_9852,N_8973,N_8142);
nor U9853 (N_9853,N_8077,N_8855);
nand U9854 (N_9854,N_8657,N_8706);
or U9855 (N_9855,N_8524,N_8292);
xor U9856 (N_9856,N_8645,N_8950);
and U9857 (N_9857,N_7878,N_8803);
nor U9858 (N_9858,N_8639,N_7651);
or U9859 (N_9859,N_8952,N_8167);
or U9860 (N_9860,N_8314,N_8509);
xnor U9861 (N_9861,N_8617,N_8192);
xnor U9862 (N_9862,N_8436,N_7547);
or U9863 (N_9863,N_7847,N_8927);
or U9864 (N_9864,N_8333,N_8165);
xnor U9865 (N_9865,N_8028,N_7625);
or U9866 (N_9866,N_8119,N_7707);
and U9867 (N_9867,N_8614,N_7789);
and U9868 (N_9868,N_8126,N_8325);
xnor U9869 (N_9869,N_7601,N_8429);
nor U9870 (N_9870,N_7980,N_8974);
or U9871 (N_9871,N_8717,N_7688);
xor U9872 (N_9872,N_8051,N_8455);
and U9873 (N_9873,N_8311,N_8675);
xnor U9874 (N_9874,N_8761,N_8492);
nand U9875 (N_9875,N_8304,N_8436);
nor U9876 (N_9876,N_8282,N_8351);
xor U9877 (N_9877,N_8992,N_7724);
xor U9878 (N_9878,N_8066,N_7865);
xor U9879 (N_9879,N_8054,N_8278);
nor U9880 (N_9880,N_8193,N_8282);
xor U9881 (N_9881,N_8625,N_8985);
xnor U9882 (N_9882,N_8110,N_8178);
or U9883 (N_9883,N_8492,N_8658);
nand U9884 (N_9884,N_8051,N_7836);
or U9885 (N_9885,N_7919,N_7750);
xor U9886 (N_9886,N_8202,N_7637);
nor U9887 (N_9887,N_8994,N_8710);
xnor U9888 (N_9888,N_8171,N_8273);
xnor U9889 (N_9889,N_8098,N_7854);
xnor U9890 (N_9890,N_8682,N_8257);
nand U9891 (N_9891,N_7761,N_8007);
nand U9892 (N_9892,N_8331,N_7912);
nand U9893 (N_9893,N_8961,N_8738);
xnor U9894 (N_9894,N_8465,N_8412);
nor U9895 (N_9895,N_8937,N_7693);
nor U9896 (N_9896,N_7783,N_7838);
xnor U9897 (N_9897,N_8628,N_7629);
nor U9898 (N_9898,N_7823,N_8838);
and U9899 (N_9899,N_7729,N_8641);
or U9900 (N_9900,N_7765,N_8129);
or U9901 (N_9901,N_7989,N_8868);
or U9902 (N_9902,N_7509,N_7805);
xor U9903 (N_9903,N_8090,N_7760);
nor U9904 (N_9904,N_7801,N_8869);
xor U9905 (N_9905,N_7984,N_7626);
or U9906 (N_9906,N_8354,N_8532);
or U9907 (N_9907,N_8299,N_8704);
xnor U9908 (N_9908,N_7838,N_8599);
or U9909 (N_9909,N_8291,N_8281);
nor U9910 (N_9910,N_8416,N_8280);
and U9911 (N_9911,N_8224,N_7727);
or U9912 (N_9912,N_8356,N_7662);
xnor U9913 (N_9913,N_7882,N_8064);
nand U9914 (N_9914,N_8619,N_7670);
xnor U9915 (N_9915,N_8107,N_7664);
and U9916 (N_9916,N_7650,N_8555);
nor U9917 (N_9917,N_7757,N_7854);
nor U9918 (N_9918,N_8432,N_7773);
nand U9919 (N_9919,N_8455,N_8764);
or U9920 (N_9920,N_7942,N_8702);
xnor U9921 (N_9921,N_8985,N_7597);
xnor U9922 (N_9922,N_7737,N_8685);
nor U9923 (N_9923,N_8207,N_7561);
and U9924 (N_9924,N_8717,N_7754);
or U9925 (N_9925,N_7657,N_8509);
nor U9926 (N_9926,N_8409,N_7927);
xnor U9927 (N_9927,N_8073,N_8411);
nor U9928 (N_9928,N_7562,N_8858);
nor U9929 (N_9929,N_8917,N_8992);
xor U9930 (N_9930,N_8145,N_7560);
and U9931 (N_9931,N_8551,N_7887);
xnor U9932 (N_9932,N_7842,N_8489);
xnor U9933 (N_9933,N_8202,N_8183);
nand U9934 (N_9934,N_8321,N_7876);
or U9935 (N_9935,N_7822,N_8405);
and U9936 (N_9936,N_8518,N_8459);
xnor U9937 (N_9937,N_7659,N_7866);
nand U9938 (N_9938,N_8392,N_8076);
nand U9939 (N_9939,N_8929,N_8817);
or U9940 (N_9940,N_8497,N_8737);
nand U9941 (N_9941,N_8390,N_8711);
xor U9942 (N_9942,N_8778,N_8840);
nand U9943 (N_9943,N_8785,N_8375);
and U9944 (N_9944,N_8126,N_8185);
or U9945 (N_9945,N_7747,N_8216);
nand U9946 (N_9946,N_8251,N_7757);
xnor U9947 (N_9947,N_8161,N_7809);
or U9948 (N_9948,N_8937,N_8527);
nand U9949 (N_9949,N_8516,N_8024);
nor U9950 (N_9950,N_8650,N_7861);
and U9951 (N_9951,N_7950,N_8538);
and U9952 (N_9952,N_8401,N_8971);
nand U9953 (N_9953,N_8149,N_8610);
or U9954 (N_9954,N_8644,N_8224);
nand U9955 (N_9955,N_7931,N_8124);
and U9956 (N_9956,N_8064,N_7975);
or U9957 (N_9957,N_7824,N_8532);
or U9958 (N_9958,N_8733,N_8845);
nand U9959 (N_9959,N_8630,N_8729);
nand U9960 (N_9960,N_8449,N_8331);
nand U9961 (N_9961,N_8254,N_8111);
and U9962 (N_9962,N_8355,N_8715);
xor U9963 (N_9963,N_8226,N_8495);
xnor U9964 (N_9964,N_7583,N_7785);
or U9965 (N_9965,N_8846,N_8943);
and U9966 (N_9966,N_8887,N_7766);
nand U9967 (N_9967,N_7704,N_8977);
or U9968 (N_9968,N_8488,N_8754);
and U9969 (N_9969,N_7843,N_8595);
nor U9970 (N_9970,N_8010,N_8965);
nor U9971 (N_9971,N_7564,N_8467);
xor U9972 (N_9972,N_8423,N_7880);
nor U9973 (N_9973,N_8916,N_8917);
nor U9974 (N_9974,N_8610,N_8143);
nand U9975 (N_9975,N_8893,N_8096);
nand U9976 (N_9976,N_8319,N_8890);
nand U9977 (N_9977,N_8459,N_8385);
nand U9978 (N_9978,N_8217,N_8893);
nor U9979 (N_9979,N_8895,N_8331);
xnor U9980 (N_9980,N_7690,N_8506);
and U9981 (N_9981,N_7564,N_8418);
or U9982 (N_9982,N_8224,N_7906);
and U9983 (N_9983,N_8572,N_8666);
or U9984 (N_9984,N_8517,N_7675);
xor U9985 (N_9985,N_7852,N_8740);
and U9986 (N_9986,N_8679,N_8998);
xor U9987 (N_9987,N_8467,N_8734);
or U9988 (N_9988,N_7783,N_8687);
nor U9989 (N_9989,N_8672,N_8423);
or U9990 (N_9990,N_8550,N_8112);
and U9991 (N_9991,N_7807,N_8854);
xor U9992 (N_9992,N_8217,N_8487);
xor U9993 (N_9993,N_8423,N_8636);
or U9994 (N_9994,N_8143,N_7739);
or U9995 (N_9995,N_7890,N_8395);
xnor U9996 (N_9996,N_8060,N_8562);
or U9997 (N_9997,N_7850,N_7600);
nor U9998 (N_9998,N_8742,N_8143);
or U9999 (N_9999,N_8993,N_8791);
and U10000 (N_10000,N_8469,N_8445);
or U10001 (N_10001,N_8403,N_7774);
or U10002 (N_10002,N_8980,N_7703);
or U10003 (N_10003,N_7751,N_7530);
xnor U10004 (N_10004,N_7516,N_8653);
and U10005 (N_10005,N_8753,N_8661);
and U10006 (N_10006,N_8646,N_7666);
nor U10007 (N_10007,N_8774,N_8214);
and U10008 (N_10008,N_8409,N_8462);
or U10009 (N_10009,N_8500,N_7789);
or U10010 (N_10010,N_8901,N_8589);
xnor U10011 (N_10011,N_8960,N_7862);
xor U10012 (N_10012,N_8065,N_7777);
and U10013 (N_10013,N_8613,N_8352);
and U10014 (N_10014,N_7510,N_7862);
and U10015 (N_10015,N_7688,N_8687);
or U10016 (N_10016,N_8304,N_8148);
nor U10017 (N_10017,N_7681,N_8525);
nand U10018 (N_10018,N_7805,N_8511);
nand U10019 (N_10019,N_8788,N_8130);
xnor U10020 (N_10020,N_7541,N_8223);
or U10021 (N_10021,N_7991,N_7501);
nor U10022 (N_10022,N_8807,N_8145);
and U10023 (N_10023,N_8674,N_8992);
nor U10024 (N_10024,N_8480,N_7933);
nand U10025 (N_10025,N_7775,N_8036);
nor U10026 (N_10026,N_8935,N_7725);
xor U10027 (N_10027,N_7772,N_8982);
nor U10028 (N_10028,N_8551,N_8957);
and U10029 (N_10029,N_7826,N_8529);
nand U10030 (N_10030,N_8351,N_8907);
and U10031 (N_10031,N_8932,N_8635);
or U10032 (N_10032,N_8659,N_7708);
and U10033 (N_10033,N_7649,N_8388);
or U10034 (N_10034,N_8038,N_7855);
and U10035 (N_10035,N_7761,N_8835);
nor U10036 (N_10036,N_8501,N_7882);
nand U10037 (N_10037,N_8863,N_8354);
nor U10038 (N_10038,N_8614,N_7812);
and U10039 (N_10039,N_7566,N_8899);
and U10040 (N_10040,N_8866,N_8204);
xor U10041 (N_10041,N_8668,N_8871);
and U10042 (N_10042,N_8450,N_8587);
nand U10043 (N_10043,N_8112,N_8667);
xnor U10044 (N_10044,N_8327,N_8989);
nor U10045 (N_10045,N_8548,N_7501);
nand U10046 (N_10046,N_8903,N_8944);
and U10047 (N_10047,N_7935,N_7933);
nor U10048 (N_10048,N_8265,N_8666);
xor U10049 (N_10049,N_7909,N_8628);
or U10050 (N_10050,N_7724,N_7861);
and U10051 (N_10051,N_8771,N_7767);
or U10052 (N_10052,N_7718,N_8405);
and U10053 (N_10053,N_8160,N_7569);
nor U10054 (N_10054,N_8801,N_8221);
and U10055 (N_10055,N_8419,N_8899);
and U10056 (N_10056,N_8967,N_8272);
xor U10057 (N_10057,N_7569,N_8181);
and U10058 (N_10058,N_8847,N_8055);
nor U10059 (N_10059,N_7641,N_8105);
xnor U10060 (N_10060,N_8285,N_8996);
nand U10061 (N_10061,N_8336,N_8850);
xnor U10062 (N_10062,N_7741,N_7520);
xor U10063 (N_10063,N_7987,N_8895);
nand U10064 (N_10064,N_8625,N_8506);
xnor U10065 (N_10065,N_8998,N_8860);
or U10066 (N_10066,N_8647,N_8564);
nand U10067 (N_10067,N_7887,N_8101);
or U10068 (N_10068,N_7857,N_8317);
xor U10069 (N_10069,N_7965,N_7535);
or U10070 (N_10070,N_7960,N_8762);
and U10071 (N_10071,N_7558,N_8018);
xnor U10072 (N_10072,N_7945,N_8805);
nand U10073 (N_10073,N_8229,N_8216);
nand U10074 (N_10074,N_7808,N_8172);
nand U10075 (N_10075,N_7801,N_7845);
nor U10076 (N_10076,N_7687,N_7789);
nor U10077 (N_10077,N_7959,N_8338);
xor U10078 (N_10078,N_8157,N_8977);
or U10079 (N_10079,N_8530,N_8441);
nand U10080 (N_10080,N_7694,N_8883);
xnor U10081 (N_10081,N_8326,N_7543);
and U10082 (N_10082,N_7640,N_7873);
nand U10083 (N_10083,N_7865,N_8508);
xor U10084 (N_10084,N_7743,N_8666);
nor U10085 (N_10085,N_8046,N_8419);
or U10086 (N_10086,N_8328,N_8124);
xnor U10087 (N_10087,N_7800,N_7852);
and U10088 (N_10088,N_8675,N_8313);
xnor U10089 (N_10089,N_7529,N_8166);
nor U10090 (N_10090,N_8236,N_7696);
xor U10091 (N_10091,N_8429,N_8196);
or U10092 (N_10092,N_7611,N_8193);
xor U10093 (N_10093,N_7973,N_8425);
nand U10094 (N_10094,N_8838,N_8283);
nand U10095 (N_10095,N_8206,N_8723);
nand U10096 (N_10096,N_8532,N_7784);
and U10097 (N_10097,N_8027,N_8650);
or U10098 (N_10098,N_7659,N_8114);
and U10099 (N_10099,N_8745,N_8203);
or U10100 (N_10100,N_8960,N_8458);
nor U10101 (N_10101,N_8789,N_8114);
nand U10102 (N_10102,N_7523,N_8858);
nor U10103 (N_10103,N_7711,N_8708);
or U10104 (N_10104,N_7664,N_8258);
nor U10105 (N_10105,N_7902,N_8108);
nor U10106 (N_10106,N_8936,N_8206);
nor U10107 (N_10107,N_7733,N_8678);
nand U10108 (N_10108,N_8104,N_8384);
xnor U10109 (N_10109,N_8430,N_8627);
nor U10110 (N_10110,N_8832,N_8709);
xor U10111 (N_10111,N_8537,N_8726);
or U10112 (N_10112,N_8964,N_8254);
and U10113 (N_10113,N_8093,N_8148);
and U10114 (N_10114,N_8694,N_8527);
and U10115 (N_10115,N_8316,N_8232);
nor U10116 (N_10116,N_8532,N_8038);
nor U10117 (N_10117,N_8242,N_8741);
xor U10118 (N_10118,N_7929,N_7999);
or U10119 (N_10119,N_8442,N_7537);
nand U10120 (N_10120,N_8499,N_8697);
and U10121 (N_10121,N_8327,N_7511);
or U10122 (N_10122,N_8452,N_8405);
and U10123 (N_10123,N_8431,N_8354);
or U10124 (N_10124,N_8800,N_8857);
nor U10125 (N_10125,N_8555,N_8984);
or U10126 (N_10126,N_8289,N_8657);
xor U10127 (N_10127,N_7555,N_7557);
and U10128 (N_10128,N_8033,N_8548);
xor U10129 (N_10129,N_8431,N_8753);
nand U10130 (N_10130,N_8574,N_8698);
nand U10131 (N_10131,N_7635,N_7977);
nand U10132 (N_10132,N_8946,N_8741);
or U10133 (N_10133,N_8245,N_8160);
xor U10134 (N_10134,N_8902,N_7578);
and U10135 (N_10135,N_8212,N_8645);
or U10136 (N_10136,N_8220,N_8781);
xnor U10137 (N_10137,N_7996,N_8595);
or U10138 (N_10138,N_8887,N_8970);
xnor U10139 (N_10139,N_7962,N_8589);
or U10140 (N_10140,N_7680,N_7639);
and U10141 (N_10141,N_7949,N_8283);
and U10142 (N_10142,N_8655,N_8553);
xor U10143 (N_10143,N_7809,N_8550);
or U10144 (N_10144,N_8699,N_7734);
and U10145 (N_10145,N_8355,N_8406);
nor U10146 (N_10146,N_8467,N_7954);
nand U10147 (N_10147,N_7525,N_8188);
nor U10148 (N_10148,N_8392,N_8560);
xor U10149 (N_10149,N_8372,N_8534);
and U10150 (N_10150,N_8896,N_7620);
and U10151 (N_10151,N_8888,N_8872);
nor U10152 (N_10152,N_8505,N_7781);
nor U10153 (N_10153,N_8227,N_8601);
nor U10154 (N_10154,N_8182,N_8542);
and U10155 (N_10155,N_8228,N_8383);
nand U10156 (N_10156,N_8642,N_8329);
nor U10157 (N_10157,N_7758,N_8203);
xnor U10158 (N_10158,N_8878,N_8859);
nand U10159 (N_10159,N_7664,N_8361);
nand U10160 (N_10160,N_8513,N_8012);
nor U10161 (N_10161,N_8250,N_7724);
nor U10162 (N_10162,N_8804,N_8428);
nand U10163 (N_10163,N_8839,N_8060);
nor U10164 (N_10164,N_8363,N_7968);
xor U10165 (N_10165,N_8980,N_8684);
nor U10166 (N_10166,N_8680,N_8631);
or U10167 (N_10167,N_7843,N_7507);
or U10168 (N_10168,N_8930,N_7786);
nand U10169 (N_10169,N_8399,N_7600);
xor U10170 (N_10170,N_8003,N_8817);
nand U10171 (N_10171,N_7673,N_7915);
and U10172 (N_10172,N_7528,N_8125);
or U10173 (N_10173,N_8650,N_8564);
xnor U10174 (N_10174,N_8887,N_8931);
nor U10175 (N_10175,N_7926,N_8347);
or U10176 (N_10176,N_7644,N_7794);
xor U10177 (N_10177,N_8341,N_7956);
nor U10178 (N_10178,N_7746,N_8907);
nand U10179 (N_10179,N_8164,N_7689);
xor U10180 (N_10180,N_8583,N_8708);
nand U10181 (N_10181,N_8939,N_7988);
or U10182 (N_10182,N_8597,N_8403);
xor U10183 (N_10183,N_8108,N_8567);
or U10184 (N_10184,N_7763,N_8984);
and U10185 (N_10185,N_8641,N_7501);
or U10186 (N_10186,N_7932,N_8973);
and U10187 (N_10187,N_7634,N_7733);
nand U10188 (N_10188,N_7564,N_7626);
and U10189 (N_10189,N_8697,N_8019);
xnor U10190 (N_10190,N_8105,N_7741);
or U10191 (N_10191,N_7890,N_7779);
xnor U10192 (N_10192,N_7827,N_7704);
xor U10193 (N_10193,N_8429,N_8716);
or U10194 (N_10194,N_7883,N_7650);
and U10195 (N_10195,N_8769,N_7915);
or U10196 (N_10196,N_7624,N_8999);
and U10197 (N_10197,N_8290,N_7823);
and U10198 (N_10198,N_8335,N_8960);
or U10199 (N_10199,N_8999,N_8964);
nand U10200 (N_10200,N_7510,N_8784);
xnor U10201 (N_10201,N_8176,N_8823);
or U10202 (N_10202,N_8525,N_7774);
or U10203 (N_10203,N_8164,N_8825);
or U10204 (N_10204,N_7873,N_8483);
nor U10205 (N_10205,N_8125,N_7759);
and U10206 (N_10206,N_7789,N_8255);
and U10207 (N_10207,N_8830,N_8207);
and U10208 (N_10208,N_8289,N_7674);
nand U10209 (N_10209,N_8975,N_8930);
nor U10210 (N_10210,N_8350,N_7622);
nor U10211 (N_10211,N_8923,N_8322);
nor U10212 (N_10212,N_7638,N_8555);
xor U10213 (N_10213,N_7574,N_8163);
or U10214 (N_10214,N_8589,N_8033);
or U10215 (N_10215,N_8921,N_7620);
and U10216 (N_10216,N_7665,N_7756);
and U10217 (N_10217,N_8020,N_8206);
xnor U10218 (N_10218,N_7587,N_8796);
xor U10219 (N_10219,N_8455,N_8315);
nand U10220 (N_10220,N_8520,N_7709);
nand U10221 (N_10221,N_7884,N_7741);
and U10222 (N_10222,N_8820,N_8749);
xor U10223 (N_10223,N_8347,N_8262);
xor U10224 (N_10224,N_8567,N_8248);
or U10225 (N_10225,N_8207,N_8506);
and U10226 (N_10226,N_7665,N_7856);
or U10227 (N_10227,N_8791,N_8756);
nand U10228 (N_10228,N_7749,N_8844);
nand U10229 (N_10229,N_8464,N_8568);
or U10230 (N_10230,N_8008,N_8276);
xnor U10231 (N_10231,N_7991,N_8694);
nor U10232 (N_10232,N_8929,N_8421);
and U10233 (N_10233,N_7673,N_8501);
nor U10234 (N_10234,N_8520,N_8325);
nor U10235 (N_10235,N_7689,N_8876);
and U10236 (N_10236,N_8262,N_8894);
and U10237 (N_10237,N_8604,N_8339);
or U10238 (N_10238,N_8112,N_8858);
or U10239 (N_10239,N_7529,N_7646);
and U10240 (N_10240,N_7518,N_7772);
xnor U10241 (N_10241,N_8038,N_8300);
nor U10242 (N_10242,N_8523,N_7596);
or U10243 (N_10243,N_8167,N_8536);
and U10244 (N_10244,N_8481,N_8332);
or U10245 (N_10245,N_8938,N_8093);
or U10246 (N_10246,N_8202,N_7690);
nor U10247 (N_10247,N_8792,N_8011);
nor U10248 (N_10248,N_8748,N_7827);
or U10249 (N_10249,N_7974,N_7911);
nor U10250 (N_10250,N_8802,N_8651);
xnor U10251 (N_10251,N_8178,N_7570);
or U10252 (N_10252,N_8588,N_8006);
nand U10253 (N_10253,N_8142,N_8475);
xnor U10254 (N_10254,N_8025,N_8915);
or U10255 (N_10255,N_8315,N_8449);
nand U10256 (N_10256,N_8528,N_7926);
or U10257 (N_10257,N_8520,N_8971);
xor U10258 (N_10258,N_7936,N_7838);
nand U10259 (N_10259,N_8309,N_8968);
and U10260 (N_10260,N_7851,N_8268);
xnor U10261 (N_10261,N_7698,N_7954);
nor U10262 (N_10262,N_8209,N_8710);
nand U10263 (N_10263,N_8603,N_8524);
nor U10264 (N_10264,N_7715,N_8434);
nand U10265 (N_10265,N_7526,N_7764);
nand U10266 (N_10266,N_7974,N_7604);
nor U10267 (N_10267,N_8357,N_8982);
or U10268 (N_10268,N_7842,N_8859);
and U10269 (N_10269,N_7613,N_8626);
and U10270 (N_10270,N_7623,N_8058);
xor U10271 (N_10271,N_7542,N_7697);
or U10272 (N_10272,N_8227,N_8454);
xnor U10273 (N_10273,N_7858,N_8963);
nor U10274 (N_10274,N_8338,N_7780);
xnor U10275 (N_10275,N_7666,N_8589);
nor U10276 (N_10276,N_7554,N_8217);
or U10277 (N_10277,N_7636,N_7531);
nand U10278 (N_10278,N_7646,N_8876);
and U10279 (N_10279,N_8965,N_8767);
xor U10280 (N_10280,N_8494,N_7949);
or U10281 (N_10281,N_8468,N_8046);
nand U10282 (N_10282,N_7625,N_8359);
nor U10283 (N_10283,N_8232,N_8714);
nor U10284 (N_10284,N_7782,N_7564);
xor U10285 (N_10285,N_8448,N_8879);
nand U10286 (N_10286,N_8030,N_8593);
or U10287 (N_10287,N_8689,N_7690);
nand U10288 (N_10288,N_7948,N_7862);
and U10289 (N_10289,N_8542,N_8600);
xnor U10290 (N_10290,N_8920,N_8549);
or U10291 (N_10291,N_8675,N_8818);
or U10292 (N_10292,N_7989,N_7759);
nand U10293 (N_10293,N_8303,N_7641);
nor U10294 (N_10294,N_7796,N_8880);
nand U10295 (N_10295,N_8484,N_8950);
and U10296 (N_10296,N_8991,N_7549);
and U10297 (N_10297,N_8917,N_8477);
xnor U10298 (N_10298,N_8187,N_7506);
nand U10299 (N_10299,N_8976,N_8591);
and U10300 (N_10300,N_7860,N_8473);
nand U10301 (N_10301,N_8634,N_8188);
nand U10302 (N_10302,N_8137,N_7501);
nand U10303 (N_10303,N_8710,N_7956);
nand U10304 (N_10304,N_8066,N_7668);
nor U10305 (N_10305,N_8327,N_7842);
nor U10306 (N_10306,N_8290,N_8933);
xor U10307 (N_10307,N_8780,N_8235);
nor U10308 (N_10308,N_8587,N_8535);
nand U10309 (N_10309,N_7819,N_7953);
or U10310 (N_10310,N_7773,N_8852);
and U10311 (N_10311,N_8848,N_7715);
and U10312 (N_10312,N_7612,N_7887);
and U10313 (N_10313,N_7807,N_8263);
nand U10314 (N_10314,N_7987,N_8955);
or U10315 (N_10315,N_8102,N_8038);
or U10316 (N_10316,N_8391,N_8754);
xnor U10317 (N_10317,N_8394,N_8888);
xnor U10318 (N_10318,N_8414,N_8285);
or U10319 (N_10319,N_8474,N_8922);
nor U10320 (N_10320,N_8935,N_8125);
and U10321 (N_10321,N_8776,N_7756);
or U10322 (N_10322,N_8835,N_8857);
or U10323 (N_10323,N_8778,N_7758);
nand U10324 (N_10324,N_7900,N_8805);
or U10325 (N_10325,N_8639,N_8862);
xor U10326 (N_10326,N_7653,N_8840);
and U10327 (N_10327,N_8428,N_8536);
xor U10328 (N_10328,N_8606,N_8882);
xor U10329 (N_10329,N_8771,N_8438);
or U10330 (N_10330,N_7793,N_8642);
or U10331 (N_10331,N_8756,N_8310);
and U10332 (N_10332,N_7647,N_7939);
xor U10333 (N_10333,N_8398,N_8747);
xor U10334 (N_10334,N_8685,N_8168);
nor U10335 (N_10335,N_8221,N_8768);
xor U10336 (N_10336,N_8239,N_8006);
or U10337 (N_10337,N_7562,N_8686);
nor U10338 (N_10338,N_8458,N_8589);
nor U10339 (N_10339,N_8922,N_7847);
or U10340 (N_10340,N_8067,N_8395);
nand U10341 (N_10341,N_8094,N_8602);
xnor U10342 (N_10342,N_8136,N_8510);
xor U10343 (N_10343,N_8203,N_8508);
and U10344 (N_10344,N_8311,N_7547);
nor U10345 (N_10345,N_8565,N_8652);
or U10346 (N_10346,N_8198,N_7866);
nor U10347 (N_10347,N_7950,N_8074);
or U10348 (N_10348,N_7675,N_8460);
or U10349 (N_10349,N_7715,N_8593);
xor U10350 (N_10350,N_7649,N_8983);
and U10351 (N_10351,N_7822,N_7724);
nand U10352 (N_10352,N_7864,N_7654);
and U10353 (N_10353,N_8181,N_7785);
xnor U10354 (N_10354,N_7631,N_8542);
or U10355 (N_10355,N_8458,N_7527);
or U10356 (N_10356,N_7655,N_7543);
or U10357 (N_10357,N_8028,N_7897);
and U10358 (N_10358,N_7964,N_8853);
xnor U10359 (N_10359,N_8179,N_8673);
and U10360 (N_10360,N_8624,N_7777);
xnor U10361 (N_10361,N_8272,N_8548);
and U10362 (N_10362,N_8151,N_8248);
or U10363 (N_10363,N_7518,N_8422);
or U10364 (N_10364,N_7781,N_8303);
xor U10365 (N_10365,N_8510,N_7913);
or U10366 (N_10366,N_7750,N_8844);
and U10367 (N_10367,N_8362,N_8570);
nand U10368 (N_10368,N_7658,N_8488);
nand U10369 (N_10369,N_8975,N_8046);
nand U10370 (N_10370,N_8388,N_8323);
nand U10371 (N_10371,N_8383,N_8504);
nand U10372 (N_10372,N_8792,N_8500);
nor U10373 (N_10373,N_8827,N_7762);
nand U10374 (N_10374,N_7532,N_8513);
and U10375 (N_10375,N_8151,N_8075);
and U10376 (N_10376,N_8098,N_7985);
and U10377 (N_10377,N_7767,N_7875);
and U10378 (N_10378,N_7943,N_8652);
and U10379 (N_10379,N_8217,N_8107);
nor U10380 (N_10380,N_7932,N_8452);
or U10381 (N_10381,N_8868,N_8464);
xnor U10382 (N_10382,N_8778,N_8025);
xnor U10383 (N_10383,N_8327,N_8983);
and U10384 (N_10384,N_8716,N_8561);
xnor U10385 (N_10385,N_8267,N_7696);
nor U10386 (N_10386,N_8527,N_8562);
xor U10387 (N_10387,N_7593,N_8515);
xor U10388 (N_10388,N_8770,N_8768);
nor U10389 (N_10389,N_8189,N_8596);
or U10390 (N_10390,N_7675,N_7524);
or U10391 (N_10391,N_8956,N_8545);
or U10392 (N_10392,N_7512,N_7782);
and U10393 (N_10393,N_8800,N_8767);
xnor U10394 (N_10394,N_7727,N_7549);
nor U10395 (N_10395,N_7723,N_8628);
nand U10396 (N_10396,N_8668,N_8866);
and U10397 (N_10397,N_8732,N_7797);
xnor U10398 (N_10398,N_8174,N_8584);
nor U10399 (N_10399,N_8545,N_8248);
and U10400 (N_10400,N_7806,N_7912);
and U10401 (N_10401,N_8032,N_7880);
nand U10402 (N_10402,N_8740,N_8934);
or U10403 (N_10403,N_7954,N_7818);
or U10404 (N_10404,N_8269,N_8235);
or U10405 (N_10405,N_8618,N_8120);
nand U10406 (N_10406,N_8908,N_8812);
nor U10407 (N_10407,N_8684,N_8521);
and U10408 (N_10408,N_8366,N_8779);
or U10409 (N_10409,N_7763,N_8893);
nor U10410 (N_10410,N_8133,N_7718);
or U10411 (N_10411,N_8422,N_7508);
nand U10412 (N_10412,N_7637,N_7823);
nor U10413 (N_10413,N_7672,N_8941);
and U10414 (N_10414,N_7653,N_8607);
and U10415 (N_10415,N_8862,N_8614);
and U10416 (N_10416,N_8636,N_8264);
nand U10417 (N_10417,N_8283,N_7915);
and U10418 (N_10418,N_8272,N_8624);
nor U10419 (N_10419,N_8593,N_7696);
or U10420 (N_10420,N_7665,N_8502);
xor U10421 (N_10421,N_7899,N_8808);
and U10422 (N_10422,N_8754,N_8644);
and U10423 (N_10423,N_7966,N_8597);
nor U10424 (N_10424,N_8004,N_7938);
or U10425 (N_10425,N_8210,N_8769);
and U10426 (N_10426,N_8586,N_8502);
nand U10427 (N_10427,N_7955,N_7615);
and U10428 (N_10428,N_8952,N_8083);
xnor U10429 (N_10429,N_7937,N_7714);
xnor U10430 (N_10430,N_8786,N_7991);
nor U10431 (N_10431,N_8134,N_7635);
nor U10432 (N_10432,N_7677,N_8759);
xor U10433 (N_10433,N_7575,N_7782);
xnor U10434 (N_10434,N_8056,N_7518);
xnor U10435 (N_10435,N_8021,N_8145);
and U10436 (N_10436,N_7526,N_8407);
or U10437 (N_10437,N_8688,N_8590);
nand U10438 (N_10438,N_8143,N_8843);
nand U10439 (N_10439,N_8346,N_8897);
and U10440 (N_10440,N_7757,N_7855);
or U10441 (N_10441,N_8838,N_8134);
nor U10442 (N_10442,N_8609,N_8356);
and U10443 (N_10443,N_7601,N_8010);
nor U10444 (N_10444,N_8832,N_8689);
or U10445 (N_10445,N_8940,N_7712);
and U10446 (N_10446,N_8889,N_8500);
nand U10447 (N_10447,N_8150,N_8617);
or U10448 (N_10448,N_8886,N_8961);
or U10449 (N_10449,N_7811,N_8569);
and U10450 (N_10450,N_7864,N_8251);
xnor U10451 (N_10451,N_7922,N_8796);
nor U10452 (N_10452,N_8807,N_7609);
nand U10453 (N_10453,N_8766,N_7651);
and U10454 (N_10454,N_7796,N_8957);
and U10455 (N_10455,N_7816,N_8195);
xnor U10456 (N_10456,N_8335,N_8968);
or U10457 (N_10457,N_7574,N_8651);
nand U10458 (N_10458,N_8726,N_8256);
xor U10459 (N_10459,N_7552,N_8270);
and U10460 (N_10460,N_8599,N_7855);
nand U10461 (N_10461,N_7989,N_8796);
and U10462 (N_10462,N_7560,N_8928);
and U10463 (N_10463,N_8314,N_7970);
nor U10464 (N_10464,N_7943,N_7950);
nor U10465 (N_10465,N_7755,N_8892);
nand U10466 (N_10466,N_7888,N_7703);
and U10467 (N_10467,N_7747,N_8367);
and U10468 (N_10468,N_8183,N_7658);
nor U10469 (N_10469,N_8184,N_7901);
nand U10470 (N_10470,N_8362,N_8024);
or U10471 (N_10471,N_8376,N_7789);
nand U10472 (N_10472,N_8356,N_8660);
nand U10473 (N_10473,N_8296,N_7784);
nor U10474 (N_10474,N_8356,N_7811);
nor U10475 (N_10475,N_8135,N_8446);
or U10476 (N_10476,N_7682,N_8633);
or U10477 (N_10477,N_8560,N_8256);
nand U10478 (N_10478,N_8987,N_8091);
xnor U10479 (N_10479,N_8445,N_7520);
nor U10480 (N_10480,N_8376,N_8855);
and U10481 (N_10481,N_8120,N_8846);
nand U10482 (N_10482,N_7794,N_8033);
or U10483 (N_10483,N_8204,N_7511);
and U10484 (N_10484,N_8820,N_8619);
nand U10485 (N_10485,N_8065,N_8256);
nand U10486 (N_10486,N_8377,N_8769);
and U10487 (N_10487,N_8529,N_8512);
and U10488 (N_10488,N_8168,N_8727);
nor U10489 (N_10489,N_8686,N_8309);
xor U10490 (N_10490,N_7756,N_8786);
nor U10491 (N_10491,N_8711,N_7951);
or U10492 (N_10492,N_8757,N_7620);
and U10493 (N_10493,N_8639,N_8876);
nand U10494 (N_10494,N_8518,N_8308);
nand U10495 (N_10495,N_8209,N_8164);
or U10496 (N_10496,N_8612,N_8957);
or U10497 (N_10497,N_8233,N_8880);
and U10498 (N_10498,N_8388,N_7793);
nor U10499 (N_10499,N_8435,N_8623);
xnor U10500 (N_10500,N_9670,N_9638);
and U10501 (N_10501,N_10001,N_9515);
and U10502 (N_10502,N_9088,N_9754);
and U10503 (N_10503,N_9265,N_9955);
or U10504 (N_10504,N_9220,N_10106);
or U10505 (N_10505,N_9390,N_9616);
or U10506 (N_10506,N_9486,N_10299);
or U10507 (N_10507,N_9214,N_9467);
nor U10508 (N_10508,N_9983,N_9854);
xor U10509 (N_10509,N_10103,N_10034);
or U10510 (N_10510,N_9816,N_10082);
nand U10511 (N_10511,N_9419,N_10029);
xnor U10512 (N_10512,N_9328,N_9618);
or U10513 (N_10513,N_9764,N_9026);
xor U10514 (N_10514,N_10204,N_9911);
or U10515 (N_10515,N_9239,N_9921);
or U10516 (N_10516,N_9685,N_9741);
and U10517 (N_10517,N_10014,N_9292);
or U10518 (N_10518,N_10385,N_9534);
and U10519 (N_10519,N_9510,N_9468);
nor U10520 (N_10520,N_9182,N_9123);
or U10521 (N_10521,N_10165,N_9868);
nor U10522 (N_10522,N_9080,N_9284);
and U10523 (N_10523,N_9682,N_10364);
nor U10524 (N_10524,N_9283,N_9811);
nor U10525 (N_10525,N_9228,N_9382);
and U10526 (N_10526,N_9938,N_10116);
or U10527 (N_10527,N_10188,N_9025);
nor U10528 (N_10528,N_9307,N_9386);
or U10529 (N_10529,N_10187,N_10419);
xnor U10530 (N_10530,N_9491,N_9998);
nand U10531 (N_10531,N_9936,N_9312);
nor U10532 (N_10532,N_9321,N_10412);
and U10533 (N_10533,N_10448,N_9412);
xor U10534 (N_10534,N_9848,N_10214);
or U10535 (N_10535,N_9801,N_10073);
xor U10536 (N_10536,N_9232,N_10338);
xnor U10537 (N_10537,N_10157,N_10417);
and U10538 (N_10538,N_9069,N_9314);
or U10539 (N_10539,N_10233,N_9769);
xor U10540 (N_10540,N_10046,N_9859);
nand U10541 (N_10541,N_9442,N_9432);
or U10542 (N_10542,N_9999,N_9969);
nand U10543 (N_10543,N_10362,N_9315);
xnor U10544 (N_10544,N_10420,N_9574);
or U10545 (N_10545,N_10413,N_10167);
and U10546 (N_10546,N_9610,N_9603);
or U10547 (N_10547,N_9406,N_9222);
xnor U10548 (N_10548,N_9558,N_10217);
nor U10549 (N_10549,N_10372,N_9941);
and U10550 (N_10550,N_10485,N_10063);
or U10551 (N_10551,N_9950,N_9247);
and U10552 (N_10552,N_9774,N_10440);
nor U10553 (N_10553,N_9600,N_10451);
and U10554 (N_10554,N_10269,N_9932);
nor U10555 (N_10555,N_9575,N_9837);
nor U10556 (N_10556,N_9330,N_10126);
or U10557 (N_10557,N_10345,N_9378);
xor U10558 (N_10558,N_9789,N_9552);
xor U10559 (N_10559,N_9466,N_10291);
and U10560 (N_10560,N_9579,N_9503);
nor U10561 (N_10561,N_10382,N_9150);
nand U10562 (N_10562,N_10471,N_9179);
nand U10563 (N_10563,N_9267,N_9633);
nand U10564 (N_10564,N_9186,N_9093);
or U10565 (N_10565,N_10323,N_9359);
nand U10566 (N_10566,N_9607,N_9210);
nor U10567 (N_10567,N_9641,N_9187);
and U10568 (N_10568,N_9876,N_9216);
and U10569 (N_10569,N_9734,N_10093);
nand U10570 (N_10570,N_9438,N_10488);
nand U10571 (N_10571,N_9061,N_9826);
nand U10572 (N_10572,N_10480,N_9821);
xnor U10573 (N_10573,N_9007,N_9286);
nand U10574 (N_10574,N_10322,N_9391);
nand U10575 (N_10575,N_9892,N_10139);
or U10576 (N_10576,N_9016,N_9248);
and U10577 (N_10577,N_9110,N_9383);
or U10578 (N_10578,N_9869,N_9049);
or U10579 (N_10579,N_9213,N_9522);
nor U10580 (N_10580,N_9853,N_10251);
and U10581 (N_10581,N_9287,N_10404);
xor U10582 (N_10582,N_10184,N_9925);
nor U10583 (N_10583,N_10215,N_9352);
or U10584 (N_10584,N_9835,N_9151);
nand U10585 (N_10585,N_9174,N_9626);
nand U10586 (N_10586,N_10499,N_9772);
xnor U10587 (N_10587,N_9096,N_10429);
xor U10588 (N_10588,N_9116,N_9430);
nor U10589 (N_10589,N_9591,N_9797);
or U10590 (N_10590,N_9608,N_9800);
and U10591 (N_10591,N_9855,N_10314);
nand U10592 (N_10592,N_9888,N_9875);
nand U10593 (N_10593,N_10444,N_9071);
nor U10594 (N_10594,N_10386,N_9254);
and U10595 (N_10595,N_10361,N_9237);
xnor U10596 (N_10596,N_10181,N_9379);
or U10597 (N_10597,N_9554,N_9846);
nor U10598 (N_10598,N_9528,N_10459);
or U10599 (N_10599,N_9565,N_9631);
xnor U10600 (N_10600,N_9022,N_9326);
nor U10601 (N_10601,N_9251,N_10381);
nand U10602 (N_10602,N_10324,N_10307);
xnor U10603 (N_10603,N_9327,N_9738);
and U10604 (N_10604,N_9740,N_10434);
xnor U10605 (N_10605,N_9481,N_10258);
xor U10606 (N_10606,N_9792,N_9578);
nand U10607 (N_10607,N_9423,N_9995);
nor U10608 (N_10608,N_10278,N_10332);
nand U10609 (N_10609,N_10042,N_9289);
nand U10610 (N_10610,N_10030,N_9097);
xor U10611 (N_10611,N_9172,N_9725);
and U10612 (N_10612,N_9744,N_9648);
xor U10613 (N_10613,N_9791,N_9297);
xor U10614 (N_10614,N_10170,N_10473);
xor U10615 (N_10615,N_9871,N_9862);
xor U10616 (N_10616,N_10153,N_9303);
xnor U10617 (N_10617,N_10067,N_9877);
and U10618 (N_10618,N_10129,N_9490);
nor U10619 (N_10619,N_9465,N_10221);
or U10620 (N_10620,N_10032,N_9593);
nand U10621 (N_10621,N_9394,N_9900);
nand U10622 (N_10622,N_10334,N_9006);
nand U10623 (N_10623,N_9884,N_10186);
nand U10624 (N_10624,N_9523,N_9996);
xor U10625 (N_10625,N_10293,N_10262);
and U10626 (N_10626,N_9913,N_10430);
and U10627 (N_10627,N_9197,N_10218);
or U10628 (N_10628,N_9700,N_9380);
xor U10629 (N_10629,N_10271,N_9191);
and U10630 (N_10630,N_10422,N_10131);
nor U10631 (N_10631,N_10344,N_9422);
or U10632 (N_10632,N_10267,N_10497);
and U10633 (N_10633,N_9569,N_9505);
or U10634 (N_10634,N_10354,N_9677);
or U10635 (N_10635,N_9958,N_9278);
nor U10636 (N_10636,N_9674,N_9873);
nand U10637 (N_10637,N_10283,N_9985);
nor U10638 (N_10638,N_10239,N_9949);
or U10639 (N_10639,N_9680,N_10149);
nand U10640 (N_10640,N_9755,N_9189);
nand U10641 (N_10641,N_10398,N_10077);
nor U10642 (N_10642,N_9144,N_9780);
or U10643 (N_10643,N_9167,N_9098);
xor U10644 (N_10644,N_9008,N_9389);
or U10645 (N_10645,N_9269,N_9227);
nor U10646 (N_10646,N_9033,N_9953);
or U10647 (N_10647,N_10246,N_9375);
nand U10648 (N_10648,N_9890,N_10424);
nor U10649 (N_10649,N_10125,N_10015);
and U10650 (N_10650,N_9400,N_9601);
or U10651 (N_10651,N_9904,N_10016);
nand U10652 (N_10652,N_9839,N_10260);
and U10653 (N_10653,N_10368,N_9332);
and U10654 (N_10654,N_9537,N_10486);
nor U10655 (N_10655,N_10189,N_9899);
nor U10656 (N_10656,N_9847,N_9403);
nand U10657 (N_10657,N_9479,N_9739);
or U10658 (N_10658,N_10020,N_9489);
or U10659 (N_10659,N_9166,N_10257);
and U10660 (N_10660,N_9895,N_9517);
or U10661 (N_10661,N_9605,N_9188);
nand U10662 (N_10662,N_9735,N_9291);
nand U10663 (N_10663,N_10004,N_9122);
and U10664 (N_10664,N_9543,N_9094);
and U10665 (N_10665,N_9912,N_9253);
and U10666 (N_10666,N_9689,N_9067);
nand U10667 (N_10667,N_10238,N_9243);
xnor U10668 (N_10668,N_10357,N_10330);
or U10669 (N_10669,N_9842,N_9850);
xnor U10670 (N_10670,N_9681,N_9134);
xnor U10671 (N_10671,N_9437,N_9924);
and U10672 (N_10672,N_9429,N_9849);
and U10673 (N_10673,N_9145,N_9852);
xor U10674 (N_10674,N_9997,N_9050);
nor U10675 (N_10675,N_9066,N_9015);
nand U10676 (N_10676,N_9162,N_10273);
and U10677 (N_10677,N_9181,N_9632);
nor U10678 (N_10678,N_9562,N_9651);
or U10679 (N_10679,N_9812,N_10219);
nand U10680 (N_10680,N_9054,N_9018);
xnor U10681 (N_10681,N_10234,N_10027);
and U10682 (N_10682,N_10250,N_10152);
or U10683 (N_10683,N_9087,N_10377);
nor U10684 (N_10684,N_9365,N_10370);
nand U10685 (N_10685,N_9190,N_9915);
and U10686 (N_10686,N_9539,N_9665);
and U10687 (N_10687,N_9663,N_10007);
xnor U10688 (N_10688,N_9456,N_9336);
xor U10689 (N_10689,N_9635,N_10491);
or U10690 (N_10690,N_9477,N_9952);
xor U10691 (N_10691,N_9079,N_10158);
or U10692 (N_10692,N_9559,N_9957);
nand U10693 (N_10693,N_10064,N_10247);
or U10694 (N_10694,N_9266,N_9337);
nand U10695 (N_10695,N_10208,N_10242);
nor U10696 (N_10696,N_9502,N_9991);
nor U10697 (N_10697,N_9546,N_9003);
and U10698 (N_10698,N_9860,N_9547);
xnor U10699 (N_10699,N_10328,N_9930);
or U10700 (N_10700,N_9787,N_9541);
and U10701 (N_10701,N_9751,N_9258);
nand U10702 (N_10702,N_10037,N_10353);
nor U10703 (N_10703,N_9160,N_9420);
nor U10704 (N_10704,N_10320,N_9447);
nand U10705 (N_10705,N_9139,N_9360);
nand U10706 (N_10706,N_9555,N_9777);
xor U10707 (N_10707,N_9760,N_10403);
nor U10708 (N_10708,N_9034,N_10099);
or U10709 (N_10709,N_9679,N_9310);
nor U10710 (N_10710,N_10384,N_9418);
or U10711 (N_10711,N_9200,N_9459);
or U10712 (N_10712,N_9927,N_9727);
nor U10713 (N_10713,N_10366,N_10498);
xor U10714 (N_10714,N_10285,N_9010);
and U10715 (N_10715,N_10365,N_10178);
and U10716 (N_10716,N_10155,N_9115);
or U10717 (N_10717,N_9225,N_9937);
nand U10718 (N_10718,N_9673,N_9343);
nor U10719 (N_10719,N_10468,N_10450);
nor U10720 (N_10720,N_10095,N_9730);
nor U10721 (N_10721,N_9961,N_9410);
or U10722 (N_10722,N_9276,N_9833);
nand U10723 (N_10723,N_9047,N_9105);
and U10724 (N_10724,N_10347,N_9393);
and U10725 (N_10725,N_9717,N_9401);
and U10726 (N_10726,N_9594,N_9453);
and U10727 (N_10727,N_9756,N_9678);
nor U10728 (N_10728,N_10472,N_9652);
and U10729 (N_10729,N_10150,N_9926);
nor U10730 (N_10730,N_9268,N_10091);
or U10731 (N_10731,N_9036,N_9142);
nor U10732 (N_10732,N_9712,N_9973);
or U10733 (N_10733,N_9604,N_9290);
or U10734 (N_10734,N_10484,N_9806);
nor U10735 (N_10735,N_9704,N_9940);
or U10736 (N_10736,N_10400,N_10389);
nand U10737 (N_10737,N_9507,N_10223);
or U10738 (N_10738,N_9100,N_9175);
xor U10739 (N_10739,N_9439,N_10475);
nor U10740 (N_10740,N_9907,N_9170);
or U10741 (N_10741,N_10261,N_9282);
xnor U10742 (N_10742,N_9550,N_9485);
nand U10743 (N_10743,N_9318,N_10454);
nor U10744 (N_10744,N_10296,N_9385);
and U10745 (N_10745,N_9732,N_10481);
nor U10746 (N_10746,N_9701,N_9211);
nand U10747 (N_10747,N_9989,N_9788);
and U10748 (N_10748,N_10142,N_10080);
xor U10749 (N_10749,N_9690,N_9300);
xor U10750 (N_10750,N_9639,N_9830);
and U10751 (N_10751,N_9970,N_9843);
xnor U10752 (N_10752,N_9514,N_9667);
nand U10753 (N_10753,N_9295,N_9325);
nand U10754 (N_10754,N_9082,N_9729);
nand U10755 (N_10755,N_9874,N_9368);
nand U10756 (N_10756,N_9138,N_10349);
or U10757 (N_10757,N_9392,N_9688);
nand U10758 (N_10758,N_9234,N_9250);
nand U10759 (N_10759,N_9346,N_10495);
nand U10760 (N_10760,N_10012,N_9135);
nor U10761 (N_10761,N_10105,N_10405);
or U10762 (N_10762,N_9630,N_9815);
nand U10763 (N_10763,N_10363,N_10199);
nor U10764 (N_10764,N_9834,N_9553);
and U10765 (N_10765,N_9260,N_9357);
or U10766 (N_10766,N_9778,N_9664);
or U10767 (N_10767,N_9526,N_9060);
or U10768 (N_10768,N_9484,N_10193);
or U10769 (N_10769,N_9919,N_9469);
nand U10770 (N_10770,N_9993,N_9118);
or U10771 (N_10771,N_9770,N_9095);
nor U10772 (N_10772,N_10297,N_10248);
nand U10773 (N_10773,N_10308,N_9715);
xor U10774 (N_10774,N_9982,N_9657);
xor U10775 (N_10775,N_9722,N_10263);
nor U10776 (N_10776,N_9563,N_9818);
nor U10777 (N_10777,N_9301,N_9277);
xnor U10778 (N_10778,N_9598,N_9158);
nand U10779 (N_10779,N_10051,N_9596);
nor U10780 (N_10780,N_9045,N_9500);
nor U10781 (N_10781,N_10089,N_9513);
xnor U10782 (N_10782,N_10092,N_10447);
and U10783 (N_10783,N_9345,N_9977);
nor U10784 (N_10784,N_9582,N_9483);
and U10785 (N_10785,N_9647,N_9051);
or U10786 (N_10786,N_9195,N_9387);
and U10787 (N_10787,N_9832,N_9446);
xor U10788 (N_10788,N_10036,N_9910);
xor U10789 (N_10789,N_9137,N_10043);
or U10790 (N_10790,N_10425,N_9793);
and U10791 (N_10791,N_10375,N_9627);
xnor U10792 (N_10792,N_9473,N_10060);
or U10793 (N_10793,N_9411,N_10207);
nand U10794 (N_10794,N_10453,N_9542);
and U10795 (N_10795,N_9226,N_9521);
nand U10796 (N_10796,N_9299,N_10478);
or U10797 (N_10797,N_9572,N_9173);
or U10798 (N_10798,N_9767,N_10058);
xor U10799 (N_10799,N_9714,N_9384);
or U10800 (N_10800,N_9027,N_9779);
xor U10801 (N_10801,N_9658,N_9339);
or U10802 (N_10802,N_9471,N_10226);
or U10803 (N_10803,N_9043,N_10394);
nand U10804 (N_10804,N_10418,N_10115);
nor U10805 (N_10805,N_10121,N_10339);
nand U10806 (N_10806,N_10411,N_9721);
xor U10807 (N_10807,N_9068,N_9408);
nor U10808 (N_10808,N_10492,N_9140);
nand U10809 (N_10809,N_9462,N_9568);
and U10810 (N_10810,N_9896,N_9235);
xor U10811 (N_10811,N_9205,N_10176);
nor U10812 (N_10812,N_10230,N_10331);
xnor U10813 (N_10813,N_9032,N_9723);
nand U10814 (N_10814,N_9646,N_9245);
nor U10815 (N_10815,N_9802,N_10410);
nor U10816 (N_10816,N_9595,N_10210);
nor U10817 (N_10817,N_9799,N_9076);
or U10818 (N_10818,N_10083,N_9750);
and U10819 (N_10819,N_9246,N_9693);
or U10820 (N_10820,N_9785,N_10018);
nor U10821 (N_10821,N_10359,N_10071);
nor U10822 (N_10822,N_9012,N_10062);
xor U10823 (N_10823,N_9883,N_9341);
nand U10824 (N_10824,N_10138,N_9240);
or U10825 (N_10825,N_9255,N_9388);
or U10826 (N_10826,N_10079,N_9057);
or U10827 (N_10827,N_9156,N_9091);
and U10828 (N_10828,N_9274,N_10433);
and U10829 (N_10829,N_9544,N_10168);
nand U10830 (N_10830,N_9586,N_10458);
xnor U10831 (N_10831,N_10216,N_9795);
xnor U10832 (N_10832,N_9692,N_10108);
and U10833 (N_10833,N_10387,N_9966);
xnor U10834 (N_10834,N_10346,N_10240);
nand U10835 (N_10835,N_9333,N_9203);
nor U10836 (N_10836,N_10052,N_9441);
and U10837 (N_10837,N_9407,N_10084);
xor U10838 (N_10838,N_10351,N_10054);
nor U10839 (N_10839,N_9427,N_9649);
xnor U10840 (N_10840,N_9742,N_10490);
and U10841 (N_10841,N_9219,N_10288);
or U10842 (N_10842,N_9073,N_10277);
nor U10843 (N_10843,N_10295,N_9824);
xnor U10844 (N_10844,N_9650,N_9413);
or U10845 (N_10845,N_10021,N_9273);
nor U10846 (N_10846,N_10117,N_9224);
nor U10847 (N_10847,N_10456,N_10414);
xor U10848 (N_10848,N_9233,N_10313);
nor U10849 (N_10849,N_10041,N_10100);
nor U10850 (N_10850,N_9103,N_9398);
xor U10851 (N_10851,N_9334,N_9870);
xor U10852 (N_10852,N_10132,N_9743);
nor U10853 (N_10853,N_9881,N_9112);
and U10854 (N_10854,N_9916,N_9946);
or U10855 (N_10855,N_10068,N_9951);
nor U10856 (N_10856,N_9671,N_10489);
nor U10857 (N_10857,N_10355,N_9698);
nor U10858 (N_10858,N_9004,N_10024);
and U10859 (N_10859,N_9844,N_10438);
nor U10860 (N_10860,N_9903,N_9464);
nor U10861 (N_10861,N_9520,N_9399);
nor U10862 (N_10862,N_9302,N_10002);
xor U10863 (N_10863,N_9683,N_10123);
nor U10864 (N_10864,N_9415,N_9728);
and U10865 (N_10865,N_9531,N_9794);
and U10866 (N_10866,N_9335,N_9107);
nand U10867 (N_10867,N_9487,N_10279);
nand U10868 (N_10868,N_10380,N_9599);
xor U10869 (N_10869,N_9372,N_10494);
and U10870 (N_10870,N_9381,N_9885);
xor U10871 (N_10871,N_10244,N_10148);
or U10872 (N_10872,N_9369,N_9044);
or U10873 (N_10873,N_9504,N_9587);
or U10874 (N_10874,N_9215,N_10134);
or U10875 (N_10875,N_9736,N_9019);
nand U10876 (N_10876,N_10289,N_9350);
nand U10877 (N_10877,N_9962,N_9817);
nor U10878 (N_10878,N_9055,N_9857);
nand U10879 (N_10879,N_10066,N_9083);
or U10880 (N_10880,N_9264,N_10088);
or U10881 (N_10881,N_10212,N_10039);
nor U10882 (N_10882,N_9331,N_10201);
xor U10883 (N_10883,N_9494,N_9293);
nor U10884 (N_10884,N_9452,N_9945);
or U10885 (N_10885,N_9023,N_9947);
nor U10886 (N_10886,N_9185,N_9058);
or U10887 (N_10887,N_9028,N_10104);
nand U10888 (N_10888,N_10439,N_9757);
nor U10889 (N_10889,N_9416,N_9917);
xor U10890 (N_10890,N_9676,N_9238);
nand U10891 (N_10891,N_10118,N_9040);
xor U10892 (N_10892,N_10090,N_9426);
nor U10893 (N_10893,N_9342,N_10102);
xnor U10894 (N_10894,N_10038,N_10311);
nor U10895 (N_10895,N_10048,N_10003);
or U10896 (N_10896,N_10321,N_9699);
xor U10897 (N_10897,N_10275,N_9529);
or U10898 (N_10898,N_9637,N_10009);
and U10899 (N_10899,N_9617,N_9538);
nand U10900 (N_10900,N_9898,N_9482);
nand U10901 (N_10901,N_10294,N_9322);
nor U10902 (N_10902,N_9731,N_10013);
nand U10903 (N_10903,N_9942,N_9217);
xnor U10904 (N_10904,N_9706,N_9405);
nand U10905 (N_10905,N_9782,N_10462);
or U10906 (N_10906,N_9976,N_10401);
xor U10907 (N_10907,N_10232,N_10415);
or U10908 (N_10908,N_10446,N_10195);
nor U10909 (N_10909,N_9967,N_10179);
nor U10910 (N_10910,N_9354,N_10437);
or U10911 (N_10911,N_9866,N_9752);
nor U10912 (N_10912,N_9532,N_9229);
and U10913 (N_10913,N_10135,N_9654);
and U10914 (N_10914,N_10128,N_10231);
nor U10915 (N_10915,N_10309,N_9193);
or U10916 (N_10916,N_9805,N_9906);
and U10917 (N_10917,N_10025,N_9395);
and U10918 (N_10918,N_10325,N_9978);
or U10919 (N_10919,N_9703,N_10265);
nand U10920 (N_10920,N_9763,N_9244);
xor U10921 (N_10921,N_10274,N_9825);
nand U10922 (N_10922,N_10243,N_10022);
xor U10923 (N_10923,N_10449,N_9209);
and U10924 (N_10924,N_9804,N_10317);
nand U10925 (N_10925,N_9659,N_10182);
nor U10926 (N_10926,N_10270,N_9348);
and U10927 (N_10927,N_10249,N_10360);
xnor U10928 (N_10928,N_10378,N_9472);
or U10929 (N_10929,N_9865,N_9956);
or U10930 (N_10930,N_10391,N_9710);
nor U10931 (N_10931,N_10276,N_9828);
xnor U10932 (N_10932,N_9733,N_10203);
nor U10933 (N_10933,N_9102,N_9872);
xor U10934 (N_10934,N_10194,N_9974);
xor U10935 (N_10935,N_10040,N_10463);
nor U10936 (N_10936,N_9509,N_9454);
or U10937 (N_10937,N_9905,N_9449);
nand U10938 (N_10938,N_10044,N_9349);
and U10939 (N_10939,N_9147,N_9719);
nand U10940 (N_10940,N_9512,N_9707);
or U10941 (N_10941,N_9908,N_10033);
nand U10942 (N_10942,N_9909,N_9672);
nand U10943 (N_10943,N_9781,N_9275);
xor U10944 (N_10944,N_9640,N_9279);
nor U10945 (N_10945,N_9270,N_9611);
nand U10946 (N_10946,N_10312,N_9017);
nor U10947 (N_10947,N_10086,N_9445);
or U10948 (N_10948,N_9914,N_10023);
nand U10949 (N_10949,N_9128,N_9549);
nor U10950 (N_10950,N_9746,N_9880);
nand U10951 (N_10951,N_9404,N_9396);
nor U10952 (N_10952,N_9201,N_10097);
nand U10953 (N_10953,N_9992,N_10065);
or U10954 (N_10954,N_9152,N_10197);
or U10955 (N_10955,N_10122,N_9370);
xnor U10956 (N_10956,N_9053,N_10151);
or U10957 (N_10957,N_9535,N_9771);
and U10958 (N_10958,N_9622,N_9556);
or U10959 (N_10959,N_9851,N_10224);
nor U10960 (N_10960,N_10352,N_9567);
or U10961 (N_10961,N_9428,N_9972);
and U10962 (N_10962,N_9133,N_10284);
xnor U10963 (N_10963,N_9070,N_9808);
xor U10964 (N_10964,N_9994,N_9749);
nor U10965 (N_10965,N_10397,N_9433);
and U10966 (N_10966,N_9551,N_9121);
xor U10967 (N_10967,N_9371,N_10445);
and U10968 (N_10968,N_10011,N_10290);
nor U10969 (N_10969,N_9184,N_10441);
and U10970 (N_10970,N_9827,N_10427);
and U10971 (N_10971,N_9536,N_10162);
nand U10972 (N_10972,N_9620,N_10190);
and U10973 (N_10973,N_10130,N_9367);
or U10974 (N_10974,N_9455,N_9374);
and U10975 (N_10975,N_10477,N_10416);
nand U10976 (N_10976,N_10406,N_9377);
and U10977 (N_10977,N_10202,N_10160);
nor U10978 (N_10978,N_9980,N_9261);
and U10979 (N_10979,N_9702,N_10390);
nand U10980 (N_10980,N_10496,N_10335);
xor U10981 (N_10981,N_9421,N_9035);
and U10982 (N_10982,N_9461,N_9655);
and U10983 (N_10983,N_9584,N_9516);
or U10984 (N_10984,N_9747,N_9501);
nor U10985 (N_10985,N_9259,N_10049);
and U10986 (N_10986,N_9829,N_9309);
xnor U10987 (N_10987,N_9954,N_9196);
or U10988 (N_10988,N_9660,N_9208);
xor U10989 (N_10989,N_9492,N_10227);
nand U10990 (N_10990,N_9256,N_10341);
xnor U10991 (N_10991,N_10245,N_10127);
nor U10992 (N_10992,N_9499,N_10074);
and U10993 (N_10993,N_10306,N_10464);
or U10994 (N_10994,N_9161,N_9011);
or U10995 (N_10995,N_10266,N_9231);
and U10996 (N_10996,N_9959,N_10421);
xnor U10997 (N_10997,N_9533,N_9656);
or U10998 (N_10998,N_9059,N_10059);
nor U10999 (N_10999,N_9358,N_9493);
nor U11000 (N_11000,N_9939,N_9718);
nor U11001 (N_11001,N_10045,N_9005);
and U11002 (N_11002,N_9104,N_9351);
and U11003 (N_11003,N_10264,N_9643);
or U11004 (N_11004,N_9241,N_9397);
xnor U11005 (N_11005,N_9344,N_9981);
nor U11006 (N_11006,N_9496,N_9840);
nor U11007 (N_11007,N_9557,N_9585);
nand U11008 (N_11008,N_9262,N_9149);
or U11009 (N_11009,N_10423,N_9625);
and U11010 (N_11010,N_9127,N_9560);
nand U11011 (N_11011,N_9434,N_9202);
or U11012 (N_11012,N_10358,N_9319);
nor U11013 (N_11013,N_10087,N_9920);
or U11014 (N_11014,N_9037,N_9306);
nand U11015 (N_11015,N_9773,N_10169);
or U11016 (N_11016,N_9285,N_9807);
and U11017 (N_11017,N_9889,N_9819);
and U11018 (N_11018,N_9130,N_10302);
nand U11019 (N_11019,N_10383,N_9042);
nand U11020 (N_11020,N_9796,N_9165);
and U11021 (N_11021,N_9612,N_9597);
xnor U11022 (N_11022,N_10120,N_10222);
nand U11023 (N_11023,N_9443,N_9686);
and U11024 (N_11024,N_9143,N_10303);
xor U11025 (N_11025,N_9960,N_9519);
nand U11026 (N_11026,N_10144,N_9153);
and U11027 (N_11027,N_9661,N_10174);
and U11028 (N_11028,N_9831,N_10336);
or U11029 (N_11029,N_9281,N_10292);
xor U11030 (N_11030,N_9313,N_9867);
and U11031 (N_11031,N_10078,N_10198);
xor U11032 (N_11032,N_10476,N_9183);
and U11033 (N_11033,N_9099,N_9101);
or U11034 (N_11034,N_9545,N_9417);
and U11035 (N_11035,N_10301,N_10101);
nor U11036 (N_11036,N_10005,N_9030);
xor U11037 (N_11037,N_9518,N_10213);
nand U11038 (N_11038,N_10436,N_9713);
nand U11039 (N_11039,N_9581,N_9624);
nor U11040 (N_11040,N_10173,N_9046);
and U11041 (N_11041,N_10156,N_10050);
xor U11042 (N_11042,N_10316,N_9614);
and U11043 (N_11043,N_9478,N_9623);
nor U11044 (N_11044,N_9979,N_9029);
and U11045 (N_11045,N_10220,N_9931);
nand U11046 (N_11046,N_10035,N_10000);
nand U11047 (N_11047,N_9497,N_9726);
nand U11048 (N_11048,N_10229,N_9111);
or U11049 (N_11049,N_10376,N_10286);
nor U11050 (N_11050,N_9548,N_9072);
xnor U11051 (N_11051,N_9064,N_9592);
xnor U11052 (N_11052,N_9424,N_9668);
nand U11053 (N_11053,N_9052,N_9990);
or U11054 (N_11054,N_9223,N_9495);
xor U11055 (N_11055,N_10466,N_9353);
or U11056 (N_11056,N_9450,N_9606);
xor U11057 (N_11057,N_9838,N_9645);
xor U11058 (N_11058,N_9475,N_9968);
or U11059 (N_11059,N_9271,N_10070);
nand U11060 (N_11060,N_9155,N_9987);
nor U11061 (N_11061,N_10072,N_10096);
and U11062 (N_11062,N_10166,N_9933);
and U11063 (N_11063,N_9132,N_9218);
or U11064 (N_11064,N_9180,N_10017);
and U11065 (N_11065,N_10319,N_9436);
nor U11066 (N_11066,N_9745,N_9856);
nor U11067 (N_11067,N_9918,N_10056);
or U11068 (N_11068,N_10460,N_9524);
nor U11069 (N_11069,N_9965,N_9589);
xnor U11070 (N_11070,N_9236,N_10133);
or U11071 (N_11071,N_9272,N_10399);
nor U11072 (N_11072,N_9761,N_9570);
nor U11073 (N_11073,N_9923,N_9048);
or U11074 (N_11074,N_9311,N_9402);
or U11075 (N_11075,N_9963,N_9204);
nand U11076 (N_11076,N_9458,N_9530);
and U11077 (N_11077,N_10409,N_10146);
nor U11078 (N_11078,N_10443,N_9887);
xnor U11079 (N_11079,N_9836,N_10137);
nand U11080 (N_11080,N_9329,N_10348);
and U11081 (N_11081,N_10253,N_10235);
xnor U11082 (N_11082,N_9056,N_10465);
nor U11083 (N_11083,N_10457,N_9964);
or U11084 (N_11084,N_9168,N_10408);
and U11085 (N_11085,N_9988,N_9242);
and U11086 (N_11086,N_10124,N_9440);
nand U11087 (N_11087,N_9021,N_9891);
nand U11088 (N_11088,N_10367,N_9691);
and U11089 (N_11089,N_10467,N_9986);
or U11090 (N_11090,N_9577,N_9084);
xor U11091 (N_11091,N_9975,N_10373);
nor U11092 (N_11092,N_9425,N_10191);
nor U11093 (N_11093,N_9694,N_9338);
nand U11094 (N_11094,N_9841,N_9928);
nor U11095 (N_11095,N_9249,N_10236);
nor U11096 (N_11096,N_9163,N_9305);
or U11097 (N_11097,N_10395,N_10047);
or U11098 (N_11098,N_10145,N_10225);
nor U11099 (N_11099,N_9192,N_9929);
and U11100 (N_11100,N_10164,N_10340);
xnor U11101 (N_11101,N_10442,N_10028);
nor U11102 (N_11102,N_9758,N_9878);
xnor U11103 (N_11103,N_9288,N_10192);
nor U11104 (N_11104,N_9636,N_9687);
nand U11105 (N_11105,N_10010,N_9298);
xnor U11106 (N_11106,N_10172,N_9814);
nand U11107 (N_11107,N_9089,N_9366);
nand U11108 (N_11108,N_10482,N_9845);
and U11109 (N_11109,N_9984,N_9768);
nor U11110 (N_11110,N_9709,N_9198);
nor U11111 (N_11111,N_9506,N_9317);
or U11112 (N_11112,N_9644,N_9065);
and U11113 (N_11113,N_9762,N_9363);
or U11114 (N_11114,N_9457,N_9724);
nor U11115 (N_11115,N_9001,N_9820);
xor U11116 (N_11116,N_9157,N_10228);
nand U11117 (N_11117,N_9901,N_10085);
xnor U11118 (N_11118,N_10163,N_9809);
nor U11119 (N_11119,N_10110,N_10487);
nand U11120 (N_11120,N_9879,N_10259);
or U11121 (N_11121,N_9864,N_9002);
and U11122 (N_11122,N_10255,N_9257);
or U11123 (N_11123,N_10256,N_9086);
xnor U11124 (N_11124,N_10075,N_9131);
nor U11125 (N_11125,N_9221,N_9720);
and U11126 (N_11126,N_10402,N_9171);
and U11127 (N_11127,N_9194,N_9823);
xor U11128 (N_11128,N_9882,N_10200);
nand U11129 (N_11129,N_9590,N_10177);
xor U11130 (N_11130,N_10379,N_9092);
nor U11131 (N_11131,N_10057,N_9109);
nand U11132 (N_11132,N_9902,N_9316);
or U11133 (N_11133,N_9653,N_10109);
and U11134 (N_11134,N_9675,N_10094);
and U11135 (N_11135,N_9609,N_10327);
xor U11136 (N_11136,N_10111,N_9136);
or U11137 (N_11137,N_9697,N_9564);
nor U11138 (N_11138,N_10114,N_9113);
or U11139 (N_11139,N_9323,N_9634);
and U11140 (N_11140,N_10326,N_10432);
and U11141 (N_11141,N_10006,N_9935);
nor U11142 (N_11142,N_9813,N_10282);
or U11143 (N_11143,N_9460,N_10428);
nor U11144 (N_11144,N_9164,N_10026);
or U11145 (N_11145,N_9629,N_9320);
xor U11146 (N_11146,N_9148,N_9695);
or U11147 (N_11147,N_10019,N_10241);
xnor U11148 (N_11148,N_9409,N_9176);
xnor U11149 (N_11149,N_9038,N_9364);
nand U11150 (N_11150,N_9159,N_10268);
nor U11151 (N_11151,N_9508,N_9621);
xor U11152 (N_11152,N_9146,N_9561);
or U11153 (N_11153,N_9753,N_9362);
and U11154 (N_11154,N_9041,N_9766);
and U11155 (N_11155,N_10329,N_10300);
xor U11156 (N_11156,N_9619,N_9124);
nand U11157 (N_11157,N_10455,N_9613);
or U11158 (N_11158,N_9199,N_10374);
or U11159 (N_11159,N_10333,N_9263);
or U11160 (N_11160,N_9944,N_9020);
nand U11161 (N_11161,N_10180,N_10281);
or U11162 (N_11162,N_10119,N_10343);
and U11163 (N_11163,N_9571,N_9212);
nand U11164 (N_11164,N_10061,N_9085);
xnor U11165 (N_11165,N_10185,N_10310);
or U11166 (N_11166,N_9177,N_10493);
or U11167 (N_11167,N_10396,N_9141);
or U11168 (N_11168,N_9822,N_9583);
nand U11169 (N_11169,N_9108,N_9081);
and U11170 (N_11170,N_9759,N_9737);
nand U11171 (N_11171,N_10159,N_9013);
or U11172 (N_11172,N_10211,N_10393);
and U11173 (N_11173,N_9748,N_9705);
and U11174 (N_11174,N_9943,N_9527);
nand U11175 (N_11175,N_10431,N_10426);
nor U11176 (N_11176,N_9476,N_9511);
nor U11177 (N_11177,N_9566,N_9347);
nor U11178 (N_11178,N_10474,N_9154);
xnor U11179 (N_11179,N_10237,N_10435);
and U11180 (N_11180,N_9090,N_9784);
nand U11181 (N_11181,N_10452,N_9786);
or U11182 (N_11182,N_10483,N_9296);
or U11183 (N_11183,N_10076,N_9602);
xnor U11184 (N_11184,N_10392,N_10141);
nor U11185 (N_11185,N_9803,N_10461);
and U11186 (N_11186,N_10254,N_9540);
and U11187 (N_11187,N_9230,N_9765);
and U11188 (N_11188,N_9308,N_9488);
or U11189 (N_11189,N_9340,N_10407);
or U11190 (N_11190,N_9304,N_9129);
nand U11191 (N_11191,N_9009,N_9798);
xnor U11192 (N_11192,N_9776,N_9948);
or U11193 (N_11193,N_9294,N_10304);
nand U11194 (N_11194,N_10196,N_9075);
and U11195 (N_11195,N_9716,N_10388);
and U11196 (N_11196,N_10298,N_9373);
nor U11197 (N_11197,N_9206,N_9696);
xor U11198 (N_11198,N_10107,N_10337);
or U11199 (N_11199,N_9971,N_9775);
and U11200 (N_11200,N_9119,N_10469);
or U11201 (N_11201,N_9169,N_10305);
xor U11202 (N_11202,N_10350,N_10154);
and U11203 (N_11203,N_9934,N_9790);
nor U11204 (N_11204,N_10136,N_9444);
xor U11205 (N_11205,N_10252,N_9894);
nand U11206 (N_11206,N_10287,N_9580);
and U11207 (N_11207,N_9414,N_10205);
and U11208 (N_11208,N_9662,N_9897);
and U11209 (N_11209,N_9480,N_10342);
and U11210 (N_11210,N_9062,N_10369);
nand U11211 (N_11211,N_10209,N_10069);
xor U11212 (N_11212,N_9324,N_9039);
xnor U11213 (N_11213,N_9178,N_10280);
nand U11214 (N_11214,N_9451,N_9708);
or U11215 (N_11215,N_9628,N_9106);
nor U11216 (N_11216,N_9893,N_9435);
nand U11217 (N_11217,N_9588,N_10112);
and U11218 (N_11218,N_9669,N_10053);
or U11219 (N_11219,N_9711,N_9356);
and U11220 (N_11220,N_10356,N_10140);
xor U11221 (N_11221,N_10161,N_9252);
and U11222 (N_11222,N_9376,N_10081);
xnor U11223 (N_11223,N_9863,N_10183);
or U11224 (N_11224,N_9861,N_9498);
or U11225 (N_11225,N_9014,N_9280);
xnor U11226 (N_11226,N_10315,N_10371);
nand U11227 (N_11227,N_9074,N_9361);
nor U11228 (N_11228,N_10470,N_10272);
nor U11229 (N_11229,N_9031,N_9783);
or U11230 (N_11230,N_9642,N_10098);
nor U11231 (N_11231,N_9024,N_10147);
nor U11232 (N_11232,N_9448,N_10055);
nor U11233 (N_11233,N_10008,N_9576);
and U11234 (N_11234,N_9886,N_10031);
nand U11235 (N_11235,N_9474,N_9470);
nand U11236 (N_11236,N_9355,N_9117);
nor U11237 (N_11237,N_9463,N_9126);
and U11238 (N_11238,N_10113,N_9810);
or U11239 (N_11239,N_9858,N_9120);
nor U11240 (N_11240,N_10206,N_10171);
xnor U11241 (N_11241,N_9431,N_10479);
nand U11242 (N_11242,N_9125,N_9666);
or U11243 (N_11243,N_9063,N_9114);
xor U11244 (N_11244,N_9573,N_10175);
xor U11245 (N_11245,N_9000,N_9525);
nor U11246 (N_11246,N_9077,N_10143);
xnor U11247 (N_11247,N_10318,N_9922);
nand U11248 (N_11248,N_9207,N_9078);
nor U11249 (N_11249,N_9615,N_9684);
nand U11250 (N_11250,N_10493,N_10392);
nand U11251 (N_11251,N_9015,N_9894);
and U11252 (N_11252,N_9027,N_9306);
or U11253 (N_11253,N_9405,N_9436);
xnor U11254 (N_11254,N_10236,N_9167);
xor U11255 (N_11255,N_9595,N_9243);
nand U11256 (N_11256,N_10292,N_9278);
nand U11257 (N_11257,N_10330,N_9288);
nand U11258 (N_11258,N_10196,N_9511);
and U11259 (N_11259,N_9999,N_10345);
nand U11260 (N_11260,N_9031,N_9007);
xor U11261 (N_11261,N_9100,N_9583);
nor U11262 (N_11262,N_9380,N_9717);
or U11263 (N_11263,N_10319,N_9255);
or U11264 (N_11264,N_9359,N_10200);
xor U11265 (N_11265,N_9714,N_9311);
and U11266 (N_11266,N_9647,N_9027);
nand U11267 (N_11267,N_9726,N_10081);
or U11268 (N_11268,N_10325,N_9185);
nand U11269 (N_11269,N_9364,N_9652);
nor U11270 (N_11270,N_9032,N_9223);
nand U11271 (N_11271,N_9055,N_10149);
xor U11272 (N_11272,N_10372,N_10229);
xnor U11273 (N_11273,N_9737,N_9006);
or U11274 (N_11274,N_10329,N_9036);
and U11275 (N_11275,N_9510,N_10243);
nor U11276 (N_11276,N_10005,N_9696);
or U11277 (N_11277,N_9079,N_9046);
nor U11278 (N_11278,N_9387,N_9642);
and U11279 (N_11279,N_10149,N_9461);
and U11280 (N_11280,N_10388,N_9100);
nor U11281 (N_11281,N_10040,N_9364);
nand U11282 (N_11282,N_10426,N_10298);
nor U11283 (N_11283,N_9300,N_9354);
xnor U11284 (N_11284,N_10233,N_9902);
and U11285 (N_11285,N_10263,N_10156);
nand U11286 (N_11286,N_9834,N_10177);
and U11287 (N_11287,N_10018,N_9370);
nand U11288 (N_11288,N_9924,N_9417);
nor U11289 (N_11289,N_9734,N_9235);
and U11290 (N_11290,N_10482,N_9733);
xnor U11291 (N_11291,N_9643,N_9783);
or U11292 (N_11292,N_9370,N_9620);
or U11293 (N_11293,N_10064,N_10437);
or U11294 (N_11294,N_10144,N_9674);
nand U11295 (N_11295,N_9366,N_10361);
nor U11296 (N_11296,N_10207,N_9373);
nor U11297 (N_11297,N_10091,N_9531);
xor U11298 (N_11298,N_9249,N_9117);
nand U11299 (N_11299,N_9286,N_9371);
xnor U11300 (N_11300,N_10049,N_9088);
nor U11301 (N_11301,N_10306,N_10249);
and U11302 (N_11302,N_10218,N_10090);
nor U11303 (N_11303,N_9294,N_10213);
or U11304 (N_11304,N_10379,N_9396);
nand U11305 (N_11305,N_9584,N_9426);
nor U11306 (N_11306,N_9699,N_9176);
and U11307 (N_11307,N_10357,N_9697);
nor U11308 (N_11308,N_9247,N_10365);
nand U11309 (N_11309,N_9913,N_9193);
nand U11310 (N_11310,N_10008,N_9412);
or U11311 (N_11311,N_9860,N_10424);
nand U11312 (N_11312,N_9672,N_9577);
nor U11313 (N_11313,N_10285,N_9172);
nand U11314 (N_11314,N_10489,N_10375);
xnor U11315 (N_11315,N_9969,N_9871);
xnor U11316 (N_11316,N_10314,N_9353);
xnor U11317 (N_11317,N_10478,N_9071);
and U11318 (N_11318,N_9977,N_9835);
or U11319 (N_11319,N_10138,N_9537);
or U11320 (N_11320,N_9769,N_9062);
and U11321 (N_11321,N_9231,N_9320);
and U11322 (N_11322,N_10159,N_9668);
or U11323 (N_11323,N_10284,N_9661);
xnor U11324 (N_11324,N_9917,N_10164);
or U11325 (N_11325,N_9230,N_9775);
and U11326 (N_11326,N_10375,N_9218);
and U11327 (N_11327,N_10102,N_10154);
xnor U11328 (N_11328,N_9963,N_9566);
nor U11329 (N_11329,N_9631,N_9275);
and U11330 (N_11330,N_9558,N_9232);
or U11331 (N_11331,N_9006,N_10403);
nor U11332 (N_11332,N_9369,N_10163);
or U11333 (N_11333,N_9292,N_10221);
and U11334 (N_11334,N_10069,N_10168);
nand U11335 (N_11335,N_10011,N_9576);
nor U11336 (N_11336,N_10279,N_9599);
nand U11337 (N_11337,N_9407,N_10093);
or U11338 (N_11338,N_9584,N_10415);
xnor U11339 (N_11339,N_9643,N_9860);
nand U11340 (N_11340,N_10454,N_9306);
nor U11341 (N_11341,N_9078,N_10459);
or U11342 (N_11342,N_9682,N_10392);
xnor U11343 (N_11343,N_9044,N_10190);
nor U11344 (N_11344,N_10155,N_10144);
nand U11345 (N_11345,N_9994,N_9764);
and U11346 (N_11346,N_9978,N_9805);
nor U11347 (N_11347,N_10367,N_10090);
or U11348 (N_11348,N_10285,N_9481);
or U11349 (N_11349,N_10358,N_9870);
or U11350 (N_11350,N_9136,N_10129);
xor U11351 (N_11351,N_9112,N_10005);
and U11352 (N_11352,N_9982,N_9519);
or U11353 (N_11353,N_9362,N_9376);
nor U11354 (N_11354,N_9550,N_10256);
nand U11355 (N_11355,N_9115,N_10156);
or U11356 (N_11356,N_9547,N_9197);
and U11357 (N_11357,N_10499,N_9673);
or U11358 (N_11358,N_10454,N_10444);
nand U11359 (N_11359,N_9173,N_10286);
or U11360 (N_11360,N_9404,N_9068);
and U11361 (N_11361,N_9027,N_9633);
nand U11362 (N_11362,N_9058,N_9125);
xor U11363 (N_11363,N_9315,N_9197);
or U11364 (N_11364,N_10387,N_9158);
or U11365 (N_11365,N_10243,N_9264);
nand U11366 (N_11366,N_9754,N_10144);
or U11367 (N_11367,N_10325,N_9038);
nand U11368 (N_11368,N_9092,N_9306);
xor U11369 (N_11369,N_9538,N_10278);
and U11370 (N_11370,N_9839,N_9584);
nand U11371 (N_11371,N_9057,N_10276);
xnor U11372 (N_11372,N_9168,N_10076);
or U11373 (N_11373,N_9842,N_10231);
and U11374 (N_11374,N_9770,N_10127);
nor U11375 (N_11375,N_10069,N_9601);
nor U11376 (N_11376,N_9468,N_10454);
and U11377 (N_11377,N_10062,N_9883);
or U11378 (N_11378,N_9738,N_9621);
xor U11379 (N_11379,N_9225,N_9663);
nor U11380 (N_11380,N_10493,N_9249);
or U11381 (N_11381,N_9165,N_10341);
or U11382 (N_11382,N_9234,N_9923);
or U11383 (N_11383,N_9941,N_9248);
and U11384 (N_11384,N_10035,N_9655);
nor U11385 (N_11385,N_10313,N_9302);
nor U11386 (N_11386,N_9092,N_9039);
and U11387 (N_11387,N_10209,N_9729);
or U11388 (N_11388,N_9475,N_9837);
nor U11389 (N_11389,N_9754,N_9311);
nand U11390 (N_11390,N_9526,N_9043);
nand U11391 (N_11391,N_9895,N_9475);
xor U11392 (N_11392,N_9551,N_10439);
xor U11393 (N_11393,N_9635,N_9576);
nand U11394 (N_11394,N_9554,N_9490);
xor U11395 (N_11395,N_9571,N_9515);
or U11396 (N_11396,N_10260,N_9006);
or U11397 (N_11397,N_9825,N_10419);
or U11398 (N_11398,N_10241,N_9154);
nor U11399 (N_11399,N_10111,N_9004);
nor U11400 (N_11400,N_9093,N_10363);
xor U11401 (N_11401,N_9243,N_9788);
xnor U11402 (N_11402,N_9093,N_9075);
nand U11403 (N_11403,N_10475,N_10467);
nor U11404 (N_11404,N_9536,N_9753);
nand U11405 (N_11405,N_9920,N_9295);
and U11406 (N_11406,N_9386,N_9272);
nand U11407 (N_11407,N_9133,N_9831);
and U11408 (N_11408,N_9745,N_10273);
or U11409 (N_11409,N_10017,N_9762);
or U11410 (N_11410,N_9901,N_10301);
xnor U11411 (N_11411,N_10444,N_10493);
nor U11412 (N_11412,N_10345,N_10036);
xnor U11413 (N_11413,N_9106,N_9867);
nor U11414 (N_11414,N_9818,N_9845);
xnor U11415 (N_11415,N_9921,N_10061);
nand U11416 (N_11416,N_9626,N_9449);
nand U11417 (N_11417,N_9536,N_9409);
xnor U11418 (N_11418,N_9684,N_9993);
or U11419 (N_11419,N_10256,N_10315);
nor U11420 (N_11420,N_9633,N_9015);
or U11421 (N_11421,N_9878,N_9048);
and U11422 (N_11422,N_9926,N_9594);
nand U11423 (N_11423,N_9330,N_9643);
and U11424 (N_11424,N_10414,N_9063);
or U11425 (N_11425,N_9554,N_9684);
nand U11426 (N_11426,N_9862,N_9294);
xnor U11427 (N_11427,N_9865,N_9962);
nor U11428 (N_11428,N_10325,N_10450);
nor U11429 (N_11429,N_9379,N_9559);
or U11430 (N_11430,N_10033,N_10476);
xor U11431 (N_11431,N_10038,N_9362);
nand U11432 (N_11432,N_9444,N_9489);
and U11433 (N_11433,N_9213,N_9451);
and U11434 (N_11434,N_9717,N_10149);
or U11435 (N_11435,N_9470,N_10318);
nor U11436 (N_11436,N_10072,N_9056);
xor U11437 (N_11437,N_9306,N_10373);
nor U11438 (N_11438,N_9927,N_9211);
nand U11439 (N_11439,N_9535,N_9707);
nand U11440 (N_11440,N_9681,N_9401);
nand U11441 (N_11441,N_9279,N_10430);
nand U11442 (N_11442,N_9073,N_9814);
nor U11443 (N_11443,N_9905,N_9199);
and U11444 (N_11444,N_9356,N_10189);
nor U11445 (N_11445,N_9780,N_10142);
nand U11446 (N_11446,N_9221,N_9870);
and U11447 (N_11447,N_9891,N_9892);
or U11448 (N_11448,N_9855,N_10302);
nor U11449 (N_11449,N_9763,N_9999);
nor U11450 (N_11450,N_9910,N_9995);
and U11451 (N_11451,N_9557,N_9145);
nor U11452 (N_11452,N_9738,N_9426);
nand U11453 (N_11453,N_9897,N_10476);
nor U11454 (N_11454,N_9884,N_9625);
and U11455 (N_11455,N_9018,N_9125);
and U11456 (N_11456,N_10388,N_9305);
nor U11457 (N_11457,N_9907,N_10437);
or U11458 (N_11458,N_10382,N_9393);
nand U11459 (N_11459,N_9814,N_9167);
and U11460 (N_11460,N_9169,N_10408);
xor U11461 (N_11461,N_9756,N_10464);
and U11462 (N_11462,N_9691,N_9152);
nor U11463 (N_11463,N_10227,N_9919);
nand U11464 (N_11464,N_9205,N_9085);
and U11465 (N_11465,N_9754,N_9379);
nor U11466 (N_11466,N_9978,N_9924);
or U11467 (N_11467,N_10265,N_9928);
nand U11468 (N_11468,N_9405,N_9983);
or U11469 (N_11469,N_9188,N_9731);
nand U11470 (N_11470,N_9255,N_9366);
xor U11471 (N_11471,N_9150,N_9550);
nand U11472 (N_11472,N_10496,N_9825);
nand U11473 (N_11473,N_9434,N_9537);
nor U11474 (N_11474,N_10101,N_9875);
and U11475 (N_11475,N_9036,N_9733);
and U11476 (N_11476,N_9432,N_10102);
nand U11477 (N_11477,N_9848,N_9836);
nor U11478 (N_11478,N_9057,N_9383);
nor U11479 (N_11479,N_9877,N_10121);
nand U11480 (N_11480,N_9456,N_9913);
nor U11481 (N_11481,N_10321,N_9611);
nor U11482 (N_11482,N_9496,N_10448);
nor U11483 (N_11483,N_9912,N_9226);
or U11484 (N_11484,N_9595,N_10363);
nand U11485 (N_11485,N_9095,N_9852);
nor U11486 (N_11486,N_9938,N_9892);
nor U11487 (N_11487,N_9931,N_9522);
or U11488 (N_11488,N_10182,N_10290);
nor U11489 (N_11489,N_10169,N_9632);
nor U11490 (N_11490,N_9562,N_9483);
or U11491 (N_11491,N_9686,N_9143);
xnor U11492 (N_11492,N_10489,N_10063);
or U11493 (N_11493,N_9289,N_9343);
nor U11494 (N_11494,N_10312,N_10038);
and U11495 (N_11495,N_9345,N_9098);
xor U11496 (N_11496,N_9903,N_9775);
and U11497 (N_11497,N_9408,N_9439);
nor U11498 (N_11498,N_10034,N_10097);
or U11499 (N_11499,N_10346,N_9823);
xor U11500 (N_11500,N_10231,N_9491);
xnor U11501 (N_11501,N_9496,N_10075);
nand U11502 (N_11502,N_9143,N_9919);
nor U11503 (N_11503,N_9873,N_10249);
nor U11504 (N_11504,N_9429,N_9568);
or U11505 (N_11505,N_10214,N_10063);
or U11506 (N_11506,N_9937,N_10232);
and U11507 (N_11507,N_9693,N_9010);
nand U11508 (N_11508,N_9449,N_9836);
and U11509 (N_11509,N_9044,N_10391);
nand U11510 (N_11510,N_9468,N_9494);
nor U11511 (N_11511,N_10105,N_10497);
and U11512 (N_11512,N_9994,N_9264);
nor U11513 (N_11513,N_10340,N_9898);
or U11514 (N_11514,N_10146,N_10318);
nand U11515 (N_11515,N_10213,N_10124);
or U11516 (N_11516,N_10071,N_10073);
and U11517 (N_11517,N_9169,N_9554);
nand U11518 (N_11518,N_10464,N_9672);
and U11519 (N_11519,N_10175,N_9082);
and U11520 (N_11520,N_9965,N_9346);
or U11521 (N_11521,N_9585,N_9168);
nand U11522 (N_11522,N_9001,N_9434);
nor U11523 (N_11523,N_9008,N_9671);
nand U11524 (N_11524,N_10009,N_10354);
nand U11525 (N_11525,N_9637,N_10228);
or U11526 (N_11526,N_10496,N_9850);
xnor U11527 (N_11527,N_9728,N_9840);
nand U11528 (N_11528,N_9563,N_9642);
nand U11529 (N_11529,N_9343,N_9902);
nor U11530 (N_11530,N_9421,N_9643);
xnor U11531 (N_11531,N_9147,N_9365);
nor U11532 (N_11532,N_9449,N_9062);
or U11533 (N_11533,N_9653,N_9647);
nand U11534 (N_11534,N_10409,N_10229);
and U11535 (N_11535,N_9924,N_9501);
and U11536 (N_11536,N_9516,N_10282);
nand U11537 (N_11537,N_10295,N_9022);
nand U11538 (N_11538,N_9989,N_9596);
xnor U11539 (N_11539,N_9489,N_9689);
or U11540 (N_11540,N_9448,N_9881);
xor U11541 (N_11541,N_9790,N_9621);
or U11542 (N_11542,N_9741,N_9056);
nor U11543 (N_11543,N_9110,N_9422);
or U11544 (N_11544,N_9999,N_10384);
xnor U11545 (N_11545,N_9489,N_9132);
or U11546 (N_11546,N_9575,N_10318);
or U11547 (N_11547,N_9911,N_10116);
or U11548 (N_11548,N_10357,N_9425);
and U11549 (N_11549,N_9099,N_9356);
nand U11550 (N_11550,N_10356,N_10431);
or U11551 (N_11551,N_9322,N_10127);
or U11552 (N_11552,N_9838,N_9215);
nand U11553 (N_11553,N_10009,N_10239);
nor U11554 (N_11554,N_9149,N_9485);
xnor U11555 (N_11555,N_9069,N_9386);
xnor U11556 (N_11556,N_10172,N_9621);
nand U11557 (N_11557,N_10410,N_9093);
xor U11558 (N_11558,N_9667,N_9046);
nor U11559 (N_11559,N_9502,N_9734);
and U11560 (N_11560,N_9390,N_9096);
or U11561 (N_11561,N_10183,N_10351);
or U11562 (N_11562,N_9789,N_9591);
nor U11563 (N_11563,N_9005,N_10487);
nor U11564 (N_11564,N_9481,N_10141);
nor U11565 (N_11565,N_9554,N_9665);
nor U11566 (N_11566,N_9922,N_9401);
and U11567 (N_11567,N_10339,N_10224);
xnor U11568 (N_11568,N_9312,N_9369);
and U11569 (N_11569,N_9704,N_9770);
xor U11570 (N_11570,N_9898,N_9979);
nand U11571 (N_11571,N_10375,N_10075);
xnor U11572 (N_11572,N_9797,N_9488);
nor U11573 (N_11573,N_9750,N_10310);
nand U11574 (N_11574,N_9194,N_10287);
or U11575 (N_11575,N_9027,N_9023);
and U11576 (N_11576,N_9743,N_9127);
and U11577 (N_11577,N_10152,N_9660);
nand U11578 (N_11578,N_9479,N_10369);
xnor U11579 (N_11579,N_9115,N_9028);
xnor U11580 (N_11580,N_10186,N_9688);
nor U11581 (N_11581,N_9989,N_10159);
nor U11582 (N_11582,N_9173,N_10339);
and U11583 (N_11583,N_10360,N_9323);
and U11584 (N_11584,N_9897,N_9239);
nor U11585 (N_11585,N_10419,N_9003);
and U11586 (N_11586,N_9776,N_9548);
nor U11587 (N_11587,N_9469,N_9657);
nor U11588 (N_11588,N_9038,N_9694);
nor U11589 (N_11589,N_9852,N_9637);
and U11590 (N_11590,N_10476,N_9346);
and U11591 (N_11591,N_9068,N_10328);
xor U11592 (N_11592,N_9968,N_9622);
and U11593 (N_11593,N_9613,N_9227);
or U11594 (N_11594,N_10375,N_9132);
xor U11595 (N_11595,N_9718,N_10226);
and U11596 (N_11596,N_10493,N_9619);
or U11597 (N_11597,N_9995,N_9227);
nand U11598 (N_11598,N_9933,N_10384);
xor U11599 (N_11599,N_9412,N_9356);
and U11600 (N_11600,N_9600,N_10095);
or U11601 (N_11601,N_10029,N_9241);
and U11602 (N_11602,N_9160,N_10483);
or U11603 (N_11603,N_9021,N_10019);
nand U11604 (N_11604,N_9389,N_9600);
nor U11605 (N_11605,N_10060,N_9693);
nand U11606 (N_11606,N_9967,N_10231);
and U11607 (N_11607,N_9906,N_9780);
nand U11608 (N_11608,N_10182,N_9130);
xnor U11609 (N_11609,N_9544,N_10084);
nor U11610 (N_11610,N_10096,N_9710);
xor U11611 (N_11611,N_9229,N_9304);
nand U11612 (N_11612,N_10032,N_9462);
and U11613 (N_11613,N_10179,N_10145);
or U11614 (N_11614,N_9986,N_10410);
xor U11615 (N_11615,N_9013,N_9461);
nor U11616 (N_11616,N_9209,N_10133);
or U11617 (N_11617,N_9136,N_9700);
nor U11618 (N_11618,N_9989,N_10061);
nor U11619 (N_11619,N_9170,N_9182);
or U11620 (N_11620,N_9388,N_9451);
nand U11621 (N_11621,N_10184,N_9012);
or U11622 (N_11622,N_9421,N_10128);
xor U11623 (N_11623,N_9748,N_10031);
nand U11624 (N_11624,N_9080,N_10453);
nand U11625 (N_11625,N_10445,N_9663);
and U11626 (N_11626,N_10035,N_10409);
or U11627 (N_11627,N_9257,N_9674);
nand U11628 (N_11628,N_9591,N_10219);
xnor U11629 (N_11629,N_10170,N_10458);
nand U11630 (N_11630,N_9142,N_9702);
and U11631 (N_11631,N_9272,N_9035);
xor U11632 (N_11632,N_9864,N_10152);
xnor U11633 (N_11633,N_10378,N_9024);
or U11634 (N_11634,N_9452,N_9041);
nand U11635 (N_11635,N_10212,N_10310);
and U11636 (N_11636,N_9017,N_10093);
and U11637 (N_11637,N_9912,N_10020);
nor U11638 (N_11638,N_9748,N_9438);
nor U11639 (N_11639,N_9918,N_9696);
nor U11640 (N_11640,N_9640,N_10353);
and U11641 (N_11641,N_9047,N_10409);
or U11642 (N_11642,N_10279,N_9143);
nand U11643 (N_11643,N_9869,N_9000);
nor U11644 (N_11644,N_9113,N_10256);
or U11645 (N_11645,N_9838,N_9970);
xnor U11646 (N_11646,N_9503,N_9402);
or U11647 (N_11647,N_10277,N_10281);
nor U11648 (N_11648,N_9380,N_9108);
or U11649 (N_11649,N_9363,N_10425);
xor U11650 (N_11650,N_9374,N_9009);
nor U11651 (N_11651,N_9759,N_9584);
or U11652 (N_11652,N_9662,N_9933);
nand U11653 (N_11653,N_9113,N_9762);
or U11654 (N_11654,N_9040,N_9019);
nor U11655 (N_11655,N_9148,N_9330);
or U11656 (N_11656,N_9778,N_9222);
nand U11657 (N_11657,N_9170,N_9389);
and U11658 (N_11658,N_10360,N_10480);
xor U11659 (N_11659,N_9307,N_9618);
nand U11660 (N_11660,N_9726,N_9876);
or U11661 (N_11661,N_9955,N_9071);
and U11662 (N_11662,N_9452,N_9148);
and U11663 (N_11663,N_9445,N_9433);
nor U11664 (N_11664,N_9363,N_9230);
or U11665 (N_11665,N_9072,N_9429);
and U11666 (N_11666,N_9363,N_9375);
nor U11667 (N_11667,N_9218,N_9724);
nor U11668 (N_11668,N_9366,N_9704);
xnor U11669 (N_11669,N_9311,N_10334);
nor U11670 (N_11670,N_10069,N_10381);
xor U11671 (N_11671,N_9069,N_9936);
and U11672 (N_11672,N_10495,N_9272);
nand U11673 (N_11673,N_9384,N_10423);
nor U11674 (N_11674,N_9670,N_10383);
xor U11675 (N_11675,N_10256,N_10409);
and U11676 (N_11676,N_9585,N_10483);
or U11677 (N_11677,N_9530,N_10253);
nand U11678 (N_11678,N_10246,N_9865);
xnor U11679 (N_11679,N_9663,N_10325);
nor U11680 (N_11680,N_10182,N_10240);
nand U11681 (N_11681,N_9727,N_10189);
xor U11682 (N_11682,N_9966,N_10100);
xnor U11683 (N_11683,N_10336,N_9159);
xor U11684 (N_11684,N_9255,N_10063);
nor U11685 (N_11685,N_9759,N_9900);
nand U11686 (N_11686,N_9577,N_9487);
xnor U11687 (N_11687,N_9042,N_9600);
nor U11688 (N_11688,N_9403,N_10337);
xor U11689 (N_11689,N_9334,N_10276);
and U11690 (N_11690,N_10017,N_9974);
xnor U11691 (N_11691,N_9338,N_9492);
xnor U11692 (N_11692,N_9700,N_9652);
xnor U11693 (N_11693,N_9592,N_10005);
or U11694 (N_11694,N_9238,N_9440);
and U11695 (N_11695,N_9602,N_9589);
and U11696 (N_11696,N_9624,N_9097);
or U11697 (N_11697,N_9416,N_9517);
and U11698 (N_11698,N_9189,N_9818);
xor U11699 (N_11699,N_9566,N_10473);
and U11700 (N_11700,N_9687,N_10152);
nor U11701 (N_11701,N_10343,N_9505);
nand U11702 (N_11702,N_10193,N_9957);
and U11703 (N_11703,N_10000,N_9168);
nor U11704 (N_11704,N_9714,N_9073);
nand U11705 (N_11705,N_10375,N_9453);
xnor U11706 (N_11706,N_9802,N_10398);
or U11707 (N_11707,N_9951,N_9218);
nand U11708 (N_11708,N_10216,N_9967);
nand U11709 (N_11709,N_10206,N_9342);
or U11710 (N_11710,N_9031,N_10074);
nor U11711 (N_11711,N_10448,N_10233);
xor U11712 (N_11712,N_10145,N_9394);
nor U11713 (N_11713,N_9464,N_9881);
and U11714 (N_11714,N_9294,N_10409);
or U11715 (N_11715,N_9130,N_9938);
nand U11716 (N_11716,N_10450,N_9568);
and U11717 (N_11717,N_10131,N_9485);
nor U11718 (N_11718,N_9839,N_9070);
xnor U11719 (N_11719,N_9799,N_9557);
xnor U11720 (N_11720,N_9746,N_9691);
nand U11721 (N_11721,N_10303,N_10003);
xor U11722 (N_11722,N_9815,N_10465);
and U11723 (N_11723,N_10413,N_10201);
xor U11724 (N_11724,N_10182,N_9373);
and U11725 (N_11725,N_9628,N_9297);
nand U11726 (N_11726,N_10138,N_10033);
xor U11727 (N_11727,N_9359,N_9736);
or U11728 (N_11728,N_10254,N_10112);
nor U11729 (N_11729,N_10147,N_9180);
and U11730 (N_11730,N_10073,N_9908);
or U11731 (N_11731,N_9368,N_9829);
nand U11732 (N_11732,N_9249,N_9970);
or U11733 (N_11733,N_9586,N_9822);
nor U11734 (N_11734,N_9363,N_9575);
xor U11735 (N_11735,N_10199,N_9914);
nand U11736 (N_11736,N_9422,N_9179);
nand U11737 (N_11737,N_9251,N_10154);
nor U11738 (N_11738,N_9461,N_9797);
nand U11739 (N_11739,N_9509,N_9900);
and U11740 (N_11740,N_10192,N_9740);
and U11741 (N_11741,N_10269,N_10169);
xnor U11742 (N_11742,N_10134,N_10372);
and U11743 (N_11743,N_10196,N_9250);
xor U11744 (N_11744,N_10290,N_10137);
nor U11745 (N_11745,N_10051,N_10045);
nor U11746 (N_11746,N_9032,N_9054);
and U11747 (N_11747,N_9877,N_9516);
and U11748 (N_11748,N_9522,N_10427);
and U11749 (N_11749,N_9390,N_10235);
nand U11750 (N_11750,N_10308,N_9696);
or U11751 (N_11751,N_9410,N_10105);
nand U11752 (N_11752,N_10015,N_9959);
nand U11753 (N_11753,N_9817,N_9834);
nand U11754 (N_11754,N_9650,N_10277);
nand U11755 (N_11755,N_9405,N_10348);
nor U11756 (N_11756,N_9117,N_10260);
nand U11757 (N_11757,N_9868,N_10009);
or U11758 (N_11758,N_9642,N_9493);
nand U11759 (N_11759,N_9802,N_10217);
nand U11760 (N_11760,N_10332,N_10036);
nor U11761 (N_11761,N_9451,N_9714);
nor U11762 (N_11762,N_9072,N_9954);
xnor U11763 (N_11763,N_9830,N_9263);
xnor U11764 (N_11764,N_9804,N_10325);
nand U11765 (N_11765,N_9495,N_9898);
xnor U11766 (N_11766,N_9902,N_9142);
xnor U11767 (N_11767,N_9809,N_9657);
or U11768 (N_11768,N_9888,N_9396);
nor U11769 (N_11769,N_9110,N_9978);
nor U11770 (N_11770,N_9974,N_9296);
and U11771 (N_11771,N_10279,N_10353);
nor U11772 (N_11772,N_10409,N_9271);
xnor U11773 (N_11773,N_10218,N_9728);
or U11774 (N_11774,N_9885,N_10081);
or U11775 (N_11775,N_9784,N_9564);
xnor U11776 (N_11776,N_9422,N_9425);
or U11777 (N_11777,N_9361,N_10327);
nor U11778 (N_11778,N_9466,N_9718);
or U11779 (N_11779,N_10472,N_10497);
nand U11780 (N_11780,N_9319,N_10131);
xnor U11781 (N_11781,N_9871,N_10159);
nor U11782 (N_11782,N_9292,N_10361);
and U11783 (N_11783,N_10027,N_9354);
nor U11784 (N_11784,N_9395,N_9847);
nor U11785 (N_11785,N_10315,N_10460);
and U11786 (N_11786,N_10241,N_9465);
and U11787 (N_11787,N_10154,N_10358);
xor U11788 (N_11788,N_9827,N_9561);
nand U11789 (N_11789,N_9170,N_9107);
nand U11790 (N_11790,N_9633,N_10008);
nor U11791 (N_11791,N_9889,N_9765);
xor U11792 (N_11792,N_9827,N_9574);
xnor U11793 (N_11793,N_10468,N_9003);
nand U11794 (N_11794,N_10299,N_9712);
or U11795 (N_11795,N_9374,N_9865);
nand U11796 (N_11796,N_9973,N_10390);
nand U11797 (N_11797,N_9730,N_9280);
or U11798 (N_11798,N_9382,N_9769);
nand U11799 (N_11799,N_9701,N_9130);
nand U11800 (N_11800,N_9640,N_10110);
or U11801 (N_11801,N_9136,N_9304);
xor U11802 (N_11802,N_9464,N_9059);
or U11803 (N_11803,N_9656,N_9253);
nor U11804 (N_11804,N_9854,N_9181);
nor U11805 (N_11805,N_9551,N_10442);
xor U11806 (N_11806,N_9272,N_9332);
nor U11807 (N_11807,N_9114,N_10456);
and U11808 (N_11808,N_10371,N_9598);
and U11809 (N_11809,N_10296,N_10196);
or U11810 (N_11810,N_10062,N_10099);
nand U11811 (N_11811,N_10083,N_9422);
and U11812 (N_11812,N_9334,N_9216);
or U11813 (N_11813,N_9981,N_9909);
xor U11814 (N_11814,N_9564,N_9074);
and U11815 (N_11815,N_9983,N_9442);
and U11816 (N_11816,N_9024,N_9675);
nand U11817 (N_11817,N_10372,N_9423);
xnor U11818 (N_11818,N_9146,N_9933);
and U11819 (N_11819,N_10082,N_9309);
and U11820 (N_11820,N_9020,N_9559);
or U11821 (N_11821,N_9739,N_9125);
or U11822 (N_11822,N_9954,N_9825);
xnor U11823 (N_11823,N_10155,N_9209);
xnor U11824 (N_11824,N_9692,N_9390);
or U11825 (N_11825,N_9355,N_10329);
nor U11826 (N_11826,N_9537,N_9839);
and U11827 (N_11827,N_9778,N_9928);
or U11828 (N_11828,N_10087,N_9826);
and U11829 (N_11829,N_10217,N_9909);
xnor U11830 (N_11830,N_9320,N_9102);
xnor U11831 (N_11831,N_9843,N_10325);
xor U11832 (N_11832,N_9035,N_9889);
nor U11833 (N_11833,N_10273,N_9633);
nor U11834 (N_11834,N_9289,N_9499);
or U11835 (N_11835,N_9851,N_9746);
xor U11836 (N_11836,N_9236,N_9224);
nor U11837 (N_11837,N_10201,N_10273);
xnor U11838 (N_11838,N_9800,N_9445);
or U11839 (N_11839,N_10011,N_9507);
or U11840 (N_11840,N_10046,N_9533);
nor U11841 (N_11841,N_9182,N_10304);
nor U11842 (N_11842,N_10033,N_9903);
and U11843 (N_11843,N_9965,N_10339);
and U11844 (N_11844,N_9208,N_9158);
nor U11845 (N_11845,N_9080,N_9642);
nand U11846 (N_11846,N_9201,N_10440);
nand U11847 (N_11847,N_10483,N_9147);
and U11848 (N_11848,N_10264,N_9457);
nor U11849 (N_11849,N_9848,N_9074);
and U11850 (N_11850,N_9841,N_10106);
xor U11851 (N_11851,N_9058,N_9716);
nor U11852 (N_11852,N_10386,N_10277);
nand U11853 (N_11853,N_9671,N_9993);
nor U11854 (N_11854,N_9466,N_10409);
or U11855 (N_11855,N_9168,N_9753);
nor U11856 (N_11856,N_9642,N_9167);
xnor U11857 (N_11857,N_9793,N_9607);
xor U11858 (N_11858,N_9276,N_9355);
nand U11859 (N_11859,N_10227,N_9549);
nor U11860 (N_11860,N_10245,N_10349);
and U11861 (N_11861,N_9446,N_9676);
or U11862 (N_11862,N_10163,N_9668);
nand U11863 (N_11863,N_9092,N_10346);
xor U11864 (N_11864,N_9974,N_9053);
or U11865 (N_11865,N_9344,N_9388);
and U11866 (N_11866,N_9960,N_9782);
nand U11867 (N_11867,N_9104,N_9745);
and U11868 (N_11868,N_9612,N_10076);
or U11869 (N_11869,N_9647,N_9680);
nand U11870 (N_11870,N_10420,N_9980);
nor U11871 (N_11871,N_9603,N_9968);
and U11872 (N_11872,N_9325,N_10378);
xor U11873 (N_11873,N_10430,N_9329);
and U11874 (N_11874,N_9978,N_10013);
or U11875 (N_11875,N_10034,N_10141);
xnor U11876 (N_11876,N_9085,N_9791);
or U11877 (N_11877,N_10083,N_10099);
or U11878 (N_11878,N_9333,N_10405);
and U11879 (N_11879,N_9324,N_9538);
nand U11880 (N_11880,N_9635,N_9550);
nand U11881 (N_11881,N_9351,N_10329);
nor U11882 (N_11882,N_10193,N_9242);
nor U11883 (N_11883,N_10169,N_9515);
or U11884 (N_11884,N_9391,N_9894);
nor U11885 (N_11885,N_10161,N_10077);
nor U11886 (N_11886,N_10080,N_9878);
and U11887 (N_11887,N_9703,N_10295);
nor U11888 (N_11888,N_9712,N_9289);
and U11889 (N_11889,N_10341,N_9349);
and U11890 (N_11890,N_9994,N_10400);
xor U11891 (N_11891,N_9470,N_9218);
nor U11892 (N_11892,N_9975,N_9312);
xor U11893 (N_11893,N_10183,N_10423);
and U11894 (N_11894,N_10457,N_10216);
nor U11895 (N_11895,N_9277,N_10152);
and U11896 (N_11896,N_10202,N_10144);
nor U11897 (N_11897,N_9056,N_9368);
nor U11898 (N_11898,N_9921,N_9995);
and U11899 (N_11899,N_9831,N_10279);
xor U11900 (N_11900,N_9388,N_9216);
and U11901 (N_11901,N_9772,N_9704);
xor U11902 (N_11902,N_10026,N_9226);
nor U11903 (N_11903,N_9896,N_10393);
nand U11904 (N_11904,N_9843,N_9989);
xor U11905 (N_11905,N_9107,N_9921);
or U11906 (N_11906,N_9201,N_10016);
and U11907 (N_11907,N_10311,N_9556);
or U11908 (N_11908,N_9566,N_9477);
or U11909 (N_11909,N_9859,N_9135);
nor U11910 (N_11910,N_10353,N_9564);
and U11911 (N_11911,N_9841,N_9989);
and U11912 (N_11912,N_9502,N_9137);
nor U11913 (N_11913,N_9460,N_9201);
or U11914 (N_11914,N_9966,N_9815);
and U11915 (N_11915,N_10481,N_9018);
nor U11916 (N_11916,N_9695,N_9534);
and U11917 (N_11917,N_10206,N_10368);
xor U11918 (N_11918,N_9783,N_9091);
and U11919 (N_11919,N_9369,N_9837);
nor U11920 (N_11920,N_9448,N_9177);
xor U11921 (N_11921,N_10214,N_9614);
nor U11922 (N_11922,N_9704,N_9938);
nor U11923 (N_11923,N_10191,N_9252);
xnor U11924 (N_11924,N_9773,N_10394);
or U11925 (N_11925,N_9934,N_10164);
nand U11926 (N_11926,N_9971,N_9829);
nand U11927 (N_11927,N_10267,N_10061);
nor U11928 (N_11928,N_9979,N_9620);
or U11929 (N_11929,N_10122,N_10036);
nand U11930 (N_11930,N_9816,N_10139);
or U11931 (N_11931,N_9373,N_10090);
xnor U11932 (N_11932,N_9021,N_9448);
or U11933 (N_11933,N_10247,N_9046);
xor U11934 (N_11934,N_9415,N_9072);
nor U11935 (N_11935,N_10341,N_9534);
nand U11936 (N_11936,N_10217,N_9178);
nor U11937 (N_11937,N_9153,N_9560);
nand U11938 (N_11938,N_10036,N_9896);
or U11939 (N_11939,N_10007,N_9026);
nor U11940 (N_11940,N_9418,N_9399);
xor U11941 (N_11941,N_9429,N_10126);
and U11942 (N_11942,N_9432,N_10099);
nand U11943 (N_11943,N_9959,N_9604);
or U11944 (N_11944,N_10294,N_9765);
or U11945 (N_11945,N_9172,N_9549);
or U11946 (N_11946,N_9329,N_9787);
or U11947 (N_11947,N_10085,N_9011);
nor U11948 (N_11948,N_10367,N_10481);
and U11949 (N_11949,N_9397,N_9484);
or U11950 (N_11950,N_9015,N_10496);
nand U11951 (N_11951,N_9036,N_9649);
and U11952 (N_11952,N_9181,N_10454);
nor U11953 (N_11953,N_10377,N_10430);
nor U11954 (N_11954,N_9027,N_9358);
xor U11955 (N_11955,N_9748,N_9078);
nor U11956 (N_11956,N_10113,N_9530);
and U11957 (N_11957,N_9063,N_10490);
nand U11958 (N_11958,N_9527,N_9307);
xor U11959 (N_11959,N_9392,N_10197);
or U11960 (N_11960,N_10421,N_9671);
and U11961 (N_11961,N_9340,N_10029);
or U11962 (N_11962,N_9658,N_10313);
nand U11963 (N_11963,N_9947,N_9723);
nor U11964 (N_11964,N_9049,N_9280);
nand U11965 (N_11965,N_9866,N_9867);
or U11966 (N_11966,N_9746,N_9373);
nor U11967 (N_11967,N_9716,N_10302);
nand U11968 (N_11968,N_9860,N_10329);
xor U11969 (N_11969,N_9195,N_9348);
or U11970 (N_11970,N_10392,N_9025);
xor U11971 (N_11971,N_10323,N_10287);
nand U11972 (N_11972,N_9449,N_9047);
nand U11973 (N_11973,N_9680,N_9467);
nor U11974 (N_11974,N_9651,N_9726);
and U11975 (N_11975,N_9601,N_9070);
and U11976 (N_11976,N_9884,N_9568);
or U11977 (N_11977,N_10249,N_10073);
nor U11978 (N_11978,N_9873,N_9919);
xor U11979 (N_11979,N_9740,N_9265);
xor U11980 (N_11980,N_10277,N_9107);
xor U11981 (N_11981,N_10388,N_9817);
nand U11982 (N_11982,N_9492,N_10085);
xnor U11983 (N_11983,N_10097,N_9408);
xor U11984 (N_11984,N_10318,N_9409);
or U11985 (N_11985,N_9644,N_10104);
xor U11986 (N_11986,N_10436,N_9648);
nand U11987 (N_11987,N_9528,N_9542);
xor U11988 (N_11988,N_9280,N_10477);
nand U11989 (N_11989,N_9663,N_10255);
xnor U11990 (N_11990,N_9335,N_10124);
nor U11991 (N_11991,N_9535,N_9075);
nand U11992 (N_11992,N_9748,N_9780);
and U11993 (N_11993,N_10186,N_9513);
or U11994 (N_11994,N_9014,N_10062);
and U11995 (N_11995,N_9367,N_10441);
nand U11996 (N_11996,N_9235,N_9695);
or U11997 (N_11997,N_9209,N_9501);
xor U11998 (N_11998,N_9524,N_9363);
xnor U11999 (N_11999,N_10285,N_9085);
nor U12000 (N_12000,N_10586,N_11925);
nand U12001 (N_12001,N_11336,N_11840);
and U12002 (N_12002,N_11388,N_11694);
and U12003 (N_12003,N_11538,N_11897);
nand U12004 (N_12004,N_11273,N_11816);
or U12005 (N_12005,N_11167,N_10561);
nor U12006 (N_12006,N_11696,N_11740);
or U12007 (N_12007,N_11818,N_11408);
and U12008 (N_12008,N_11998,N_10794);
or U12009 (N_12009,N_11928,N_11211);
and U12010 (N_12010,N_11900,N_10590);
or U12011 (N_12011,N_10538,N_11459);
nor U12012 (N_12012,N_10903,N_11427);
xor U12013 (N_12013,N_10793,N_10676);
nor U12014 (N_12014,N_10762,N_11393);
nand U12015 (N_12015,N_11946,N_11610);
and U12016 (N_12016,N_11786,N_11811);
or U12017 (N_12017,N_11005,N_11402);
nor U12018 (N_12018,N_11331,N_11550);
or U12019 (N_12019,N_11062,N_11356);
nand U12020 (N_12020,N_10664,N_11440);
nand U12021 (N_12021,N_11003,N_10938);
or U12022 (N_12022,N_10691,N_10928);
or U12023 (N_12023,N_11921,N_11493);
nand U12024 (N_12024,N_10509,N_11296);
xor U12025 (N_12025,N_10521,N_11228);
and U12026 (N_12026,N_11630,N_11689);
nor U12027 (N_12027,N_11040,N_11826);
or U12028 (N_12028,N_10565,N_10967);
xnor U12029 (N_12029,N_11087,N_10599);
nor U12030 (N_12030,N_11208,N_11743);
xor U12031 (N_12031,N_11148,N_11757);
or U12032 (N_12032,N_11719,N_11654);
or U12033 (N_12033,N_11418,N_11944);
and U12034 (N_12034,N_11526,N_11589);
nor U12035 (N_12035,N_10751,N_11236);
nor U12036 (N_12036,N_11978,N_10579);
nand U12037 (N_12037,N_11241,N_11354);
or U12038 (N_12038,N_11987,N_10724);
nor U12039 (N_12039,N_11127,N_10786);
nand U12040 (N_12040,N_10936,N_10965);
or U12041 (N_12041,N_11872,N_11407);
nand U12042 (N_12042,N_10842,N_10629);
or U12043 (N_12043,N_11764,N_11159);
or U12044 (N_12044,N_10602,N_11469);
nor U12045 (N_12045,N_11319,N_11749);
or U12046 (N_12046,N_11361,N_10584);
or U12047 (N_12047,N_11633,N_10893);
and U12048 (N_12048,N_11956,N_11738);
xnor U12049 (N_12049,N_10558,N_11439);
and U12050 (N_12050,N_10706,N_11165);
xor U12051 (N_12051,N_11612,N_11118);
and U12052 (N_12052,N_11675,N_11698);
nor U12053 (N_12053,N_11929,N_11381);
nor U12054 (N_12054,N_11993,N_11559);
and U12055 (N_12055,N_11212,N_10848);
or U12056 (N_12056,N_11245,N_10686);
nor U12057 (N_12057,N_11751,N_11863);
or U12058 (N_12058,N_11170,N_11824);
nand U12059 (N_12059,N_10677,N_11379);
xor U12060 (N_12060,N_11905,N_11084);
nor U12061 (N_12061,N_11020,N_11057);
nand U12062 (N_12062,N_11515,N_11025);
nor U12063 (N_12063,N_10775,N_11155);
nor U12064 (N_12064,N_11403,N_11634);
nor U12065 (N_12065,N_11590,N_11291);
and U12066 (N_12066,N_11366,N_10866);
nor U12067 (N_12067,N_11278,N_11971);
and U12068 (N_12068,N_11500,N_11188);
and U12069 (N_12069,N_10808,N_11915);
xnor U12070 (N_12070,N_11082,N_11308);
nor U12071 (N_12071,N_11293,N_11257);
or U12072 (N_12072,N_10652,N_11669);
nor U12073 (N_12073,N_11454,N_11328);
and U12074 (N_12074,N_11373,N_11452);
and U12075 (N_12075,N_11810,N_11495);
xnor U12076 (N_12076,N_11628,N_11300);
and U12077 (N_12077,N_11244,N_10941);
or U12078 (N_12078,N_10655,N_11343);
nand U12079 (N_12079,N_11773,N_10783);
nor U12080 (N_12080,N_11924,N_10680);
and U12081 (N_12081,N_11727,N_10820);
and U12082 (N_12082,N_11842,N_11390);
nand U12083 (N_12083,N_11753,N_11825);
or U12084 (N_12084,N_11617,N_10709);
nand U12085 (N_12085,N_11594,N_11798);
and U12086 (N_12086,N_11412,N_11098);
nor U12087 (N_12087,N_10773,N_11957);
or U12088 (N_12088,N_11867,N_11329);
nor U12089 (N_12089,N_10679,N_11682);
xor U12090 (N_12090,N_11490,N_11420);
xnor U12091 (N_12091,N_10707,N_10644);
nor U12092 (N_12092,N_11939,N_11405);
and U12093 (N_12093,N_10760,N_11092);
nand U12094 (N_12094,N_11133,N_11870);
or U12095 (N_12095,N_11968,N_10733);
nand U12096 (N_12096,N_11995,N_11556);
xnor U12097 (N_12097,N_11309,N_10583);
or U12098 (N_12098,N_11176,N_10767);
xnor U12099 (N_12099,N_10744,N_10812);
xnor U12100 (N_12100,N_11504,N_10728);
and U12101 (N_12101,N_10888,N_11128);
nand U12102 (N_12102,N_10520,N_11196);
or U12103 (N_12103,N_11992,N_10777);
xor U12104 (N_12104,N_11754,N_10713);
nand U12105 (N_12105,N_11520,N_11503);
nand U12106 (N_12106,N_11985,N_11482);
or U12107 (N_12107,N_10693,N_11931);
and U12108 (N_12108,N_11829,N_11624);
nor U12109 (N_12109,N_11562,N_11117);
nand U12110 (N_12110,N_10659,N_10789);
nor U12111 (N_12111,N_11114,N_11882);
or U12112 (N_12112,N_10557,N_10572);
or U12113 (N_12113,N_11609,N_11242);
or U12114 (N_12114,N_11468,N_11576);
and U12115 (N_12115,N_11618,N_11659);
or U12116 (N_12116,N_10766,N_11352);
or U12117 (N_12117,N_11606,N_10772);
and U12118 (N_12118,N_11201,N_11638);
or U12119 (N_12119,N_10821,N_11312);
and U12120 (N_12120,N_10817,N_10543);
and U12121 (N_12121,N_10857,N_11480);
nand U12122 (N_12122,N_11431,N_11279);
nor U12123 (N_12123,N_11200,N_10588);
xor U12124 (N_12124,N_11110,N_11157);
nand U12125 (N_12125,N_10831,N_11850);
nor U12126 (N_12126,N_10625,N_11434);
xor U12127 (N_12127,N_11235,N_11737);
xnor U12128 (N_12128,N_10533,N_10883);
nand U12129 (N_12129,N_11802,N_11382);
nand U12130 (N_12130,N_10585,N_11360);
and U12131 (N_12131,N_11274,N_11717);
nor U12132 (N_12132,N_11101,N_10954);
or U12133 (N_12133,N_11316,N_11375);
and U12134 (N_12134,N_11168,N_10781);
nor U12135 (N_12135,N_11024,N_11310);
or U12136 (N_12136,N_11044,N_11093);
or U12137 (N_12137,N_10705,N_10632);
nand U12138 (N_12138,N_10610,N_11006);
and U12139 (N_12139,N_11119,N_11991);
nand U12140 (N_12140,N_11879,N_10943);
nand U12141 (N_12141,N_11856,N_11547);
or U12142 (N_12142,N_10980,N_10739);
and U12143 (N_12143,N_11951,N_10921);
or U12144 (N_12144,N_10581,N_11281);
and U12145 (N_12145,N_11714,N_11711);
xor U12146 (N_12146,N_10641,N_11999);
xnor U12147 (N_12147,N_10908,N_11037);
xnor U12148 (N_12148,N_10827,N_11641);
and U12149 (N_12149,N_11304,N_11668);
and U12150 (N_12150,N_10607,N_11019);
nor U12151 (N_12151,N_11049,N_11077);
or U12152 (N_12152,N_11184,N_10663);
nor U12153 (N_12153,N_11198,N_11901);
nor U12154 (N_12154,N_10603,N_11004);
xor U12155 (N_12155,N_11699,N_11666);
nand U12156 (N_12156,N_11016,N_11186);
nor U12157 (N_12157,N_10598,N_11301);
xor U12158 (N_12158,N_11368,N_11285);
and U12159 (N_12159,N_10665,N_11191);
or U12160 (N_12160,N_11095,N_11691);
nand U12161 (N_12161,N_11750,N_10963);
or U12162 (N_12162,N_11249,N_10506);
and U12163 (N_12163,N_11701,N_11938);
and U12164 (N_12164,N_10524,N_11142);
and U12165 (N_12165,N_11539,N_11671);
nand U12166 (N_12166,N_11483,N_10912);
nand U12167 (N_12167,N_10630,N_11709);
nor U12168 (N_12168,N_11223,N_11486);
xor U12169 (N_12169,N_11894,N_11721);
nand U12170 (N_12170,N_11359,N_11739);
and U12171 (N_12171,N_10905,N_11681);
nor U12172 (N_12172,N_11075,N_11171);
nor U12173 (N_12173,N_10896,N_11700);
and U12174 (N_12174,N_10981,N_11871);
xor U12175 (N_12175,N_10951,N_11531);
nor U12176 (N_12176,N_11017,N_11056);
nor U12177 (N_12177,N_11645,N_11510);
nor U12178 (N_12178,N_10694,N_11349);
nand U12179 (N_12179,N_10519,N_10854);
nand U12180 (N_12180,N_11649,N_11665);
nor U12181 (N_12181,N_11851,N_10648);
nor U12182 (N_12182,N_11799,N_11450);
xnor U12183 (N_12183,N_10539,N_11784);
xor U12184 (N_12184,N_11853,N_11023);
or U12185 (N_12185,N_11376,N_10720);
nor U12186 (N_12186,N_11071,N_11592);
nor U12187 (N_12187,N_11177,N_11729);
or U12188 (N_12188,N_11774,N_11578);
nand U12189 (N_12189,N_11977,N_11567);
and U12190 (N_12190,N_10993,N_10681);
and U12191 (N_12191,N_11835,N_10622);
and U12192 (N_12192,N_11085,N_10640);
nor U12193 (N_12193,N_10534,N_10688);
nand U12194 (N_12194,N_11860,N_11185);
nand U12195 (N_12195,N_11619,N_11959);
nor U12196 (N_12196,N_11306,N_11113);
nand U12197 (N_12197,N_10814,N_10745);
xor U12198 (N_12198,N_11663,N_11330);
nand U12199 (N_12199,N_10824,N_10945);
or U12200 (N_12200,N_11516,N_10708);
and U12201 (N_12201,N_10968,N_11034);
nand U12202 (N_12202,N_11580,N_10756);
or U12203 (N_12203,N_11982,N_11775);
nand U12204 (N_12204,N_10560,N_11154);
and U12205 (N_12205,N_11560,N_11371);
and U12206 (N_12206,N_10881,N_11048);
nor U12207 (N_12207,N_10889,N_11413);
or U12208 (N_12208,N_10984,N_11362);
and U12209 (N_12209,N_10568,N_10589);
xor U12210 (N_12210,N_11647,N_11730);
xor U12211 (N_12211,N_10563,N_11465);
nand U12212 (N_12212,N_10913,N_10916);
or U12213 (N_12213,N_10958,N_11785);
or U12214 (N_12214,N_11035,N_11602);
nand U12215 (N_12215,N_11636,N_10529);
nor U12216 (N_12216,N_10879,N_10942);
xnor U12217 (N_12217,N_10899,N_11920);
or U12218 (N_12218,N_11270,N_11295);
or U12219 (N_12219,N_11344,N_10931);
nor U12220 (N_12220,N_10897,N_11650);
nand U12221 (N_12221,N_11736,N_11828);
nor U12222 (N_12222,N_11126,N_10701);
or U12223 (N_12223,N_11487,N_11640);
xor U12224 (N_12224,N_10547,N_11942);
nand U12225 (N_12225,N_10878,N_10907);
nand U12226 (N_12226,N_11710,N_11426);
xor U12227 (N_12227,N_10549,N_10592);
nor U12228 (N_12228,N_10935,N_10996);
or U12229 (N_12229,N_11166,N_10782);
or U12230 (N_12230,N_10776,N_11029);
nand U12231 (N_12231,N_10518,N_11912);
nand U12232 (N_12232,N_11251,N_11069);
nor U12233 (N_12233,N_10511,N_11950);
nand U12234 (N_12234,N_10890,N_10799);
and U12235 (N_12235,N_11534,N_10505);
or U12236 (N_12236,N_10608,N_11108);
xnor U12237 (N_12237,N_11374,N_10770);
nand U12238 (N_12238,N_11706,N_10872);
or U12239 (N_12239,N_10860,N_10746);
xor U12240 (N_12240,N_10868,N_10852);
xor U12241 (N_12241,N_11178,N_11346);
and U12242 (N_12242,N_11861,N_11460);
nor U12243 (N_12243,N_11783,N_10823);
nand U12244 (N_12244,N_11975,N_10939);
nor U12245 (N_12245,N_11541,N_11410);
or U12246 (N_12246,N_11868,N_11250);
and U12247 (N_12247,N_10792,N_11845);
and U12248 (N_12248,N_11506,N_11695);
or U12249 (N_12249,N_11692,N_11657);
or U12250 (N_12250,N_11372,N_10719);
or U12251 (N_12251,N_11144,N_10887);
nor U12252 (N_12252,N_10550,N_11272);
or U12253 (N_12253,N_11181,N_10597);
and U12254 (N_12254,N_10737,N_11834);
and U12255 (N_12255,N_10825,N_11333);
or U12256 (N_12256,N_10541,N_10645);
or U12257 (N_12257,N_10643,N_11135);
nand U12258 (N_12258,N_10818,N_10934);
xnor U12259 (N_12259,N_11479,N_11151);
or U12260 (N_12260,N_11747,N_11637);
or U12261 (N_12261,N_10500,N_11656);
and U12262 (N_12262,N_10870,N_11156);
nor U12263 (N_12263,N_10712,N_10853);
nor U12264 (N_12264,N_11355,N_11684);
xor U12265 (N_12265,N_10839,N_10850);
or U12266 (N_12266,N_11297,N_10999);
nand U12267 (N_12267,N_11524,N_10873);
or U12268 (N_12268,N_11066,N_11265);
or U12269 (N_12269,N_10804,N_11790);
or U12270 (N_12270,N_11927,N_11508);
and U12271 (N_12271,N_10551,N_11341);
or U12272 (N_12272,N_11467,N_11525);
xnor U12273 (N_12273,N_11256,N_11461);
or U12274 (N_12274,N_11423,N_11216);
nand U12275 (N_12275,N_11474,N_11778);
or U12276 (N_12276,N_10956,N_11875);
nand U12277 (N_12277,N_10787,N_11464);
nand U12278 (N_12278,N_11219,N_11953);
or U12279 (N_12279,N_11591,N_10914);
and U12280 (N_12280,N_11943,N_11444);
or U12281 (N_12281,N_11478,N_11801);
and U12282 (N_12282,N_10562,N_10983);
and U12283 (N_12283,N_10990,N_11313);
nand U12284 (N_12284,N_11015,N_10695);
nand U12285 (N_12285,N_11246,N_11494);
nor U12286 (N_12286,N_10575,N_11134);
or U12287 (N_12287,N_11449,N_11396);
xor U12288 (N_12288,N_11484,N_10836);
and U12289 (N_12289,N_10944,N_11160);
nor U12290 (N_12290,N_10894,N_11908);
nand U12291 (N_12291,N_10911,N_11777);
and U12292 (N_12292,N_10721,N_11443);
nor U12293 (N_12293,N_11441,N_11583);
or U12294 (N_12294,N_11353,N_11837);
nand U12295 (N_12295,N_11597,N_11140);
xor U12296 (N_12296,N_11820,N_10710);
nor U12297 (N_12297,N_11489,N_11488);
nor U12298 (N_12298,N_10542,N_10769);
and U12299 (N_12299,N_11986,N_11760);
nor U12300 (N_12300,N_11325,N_10886);
nand U12301 (N_12301,N_10976,N_11258);
and U12302 (N_12302,N_11940,N_11453);
or U12303 (N_12303,N_10569,N_11298);
xnor U12304 (N_12304,N_11586,N_10778);
and U12305 (N_12305,N_11608,N_11103);
xnor U12306 (N_12306,N_11013,N_10633);
or U12307 (N_12307,N_11728,N_11767);
xor U12308 (N_12308,N_11261,N_10570);
nand U12309 (N_12309,N_10525,N_11970);
or U12310 (N_12310,N_11400,N_11796);
or U12311 (N_12311,N_11307,N_11880);
or U12312 (N_12312,N_11429,N_10977);
or U12313 (N_12313,N_10948,N_11145);
and U12314 (N_12314,N_11394,N_10619);
nand U12315 (N_12315,N_11415,N_11831);
and U12316 (N_12316,N_11267,N_11260);
or U12317 (N_12317,N_11146,N_11895);
nand U12318 (N_12318,N_11933,N_11169);
xor U12319 (N_12319,N_11741,N_11564);
nand U12320 (N_12320,N_10807,N_11806);
and U12321 (N_12321,N_11812,N_11389);
nand U12322 (N_12322,N_10662,N_11351);
nand U12323 (N_12323,N_11239,N_10851);
and U12324 (N_12324,N_11321,N_10650);
xnor U12325 (N_12325,N_11896,N_11161);
xnor U12326 (N_12326,N_11182,N_10763);
nand U12327 (N_12327,N_11603,N_10697);
or U12328 (N_12328,N_11137,N_11342);
and U12329 (N_12329,N_10863,N_11247);
or U12330 (N_12330,N_11776,N_11664);
nand U12331 (N_12331,N_10687,N_11887);
nand U12332 (N_12332,N_11205,N_10656);
nor U12333 (N_12333,N_10621,N_10642);
nor U12334 (N_12334,N_10832,N_11593);
nand U12335 (N_12335,N_11909,N_11147);
xor U12336 (N_12336,N_11607,N_11803);
or U12337 (N_12337,N_10513,N_10779);
and U12338 (N_12338,N_11120,N_11088);
or U12339 (N_12339,N_10544,N_10991);
xor U12340 (N_12340,N_11889,N_11187);
nand U12341 (N_12341,N_11116,N_10785);
xnor U12342 (N_12342,N_10516,N_10960);
xor U12343 (N_12343,N_11063,N_10973);
or U12344 (N_12344,N_11286,N_11522);
xor U12345 (N_12345,N_11008,N_11726);
xnor U12346 (N_12346,N_10612,N_11888);
and U12347 (N_12347,N_11220,N_10992);
nand U12348 (N_12348,N_11670,N_11746);
or U12349 (N_12349,N_11955,N_10582);
nand U12350 (N_12350,N_11948,N_10735);
or U12351 (N_12351,N_11788,N_11324);
nor U12352 (N_12352,N_11994,N_11855);
or U12353 (N_12353,N_11677,N_10540);
or U12354 (N_12354,N_11544,N_10811);
or U12355 (N_12355,N_11725,N_10546);
and U12356 (N_12356,N_10885,N_11193);
nand U12357 (N_12357,N_11012,N_11386);
nor U12358 (N_12358,N_11555,N_10578);
nand U12359 (N_12359,N_11139,N_11284);
nand U12360 (N_12360,N_11175,N_11720);
nor U12361 (N_12361,N_11916,N_11437);
xnor U12362 (N_12362,N_11667,N_11742);
nand U12363 (N_12363,N_11112,N_11813);
or U12364 (N_12364,N_11819,N_11109);
nor U12365 (N_12365,N_11363,N_10768);
or U12366 (N_12366,N_11809,N_11399);
nor U12367 (N_12367,N_11574,N_10725);
nor U12368 (N_12368,N_11124,N_11910);
nor U12369 (N_12369,N_11841,N_11862);
nand U12370 (N_12370,N_10668,N_10634);
nor U12371 (N_12371,N_11099,N_10678);
or U12372 (N_12372,N_10504,N_11289);
nand U12373 (N_12373,N_11264,N_11438);
and U12374 (N_12374,N_11129,N_10552);
nand U12375 (N_12375,N_11687,N_11262);
or U12376 (N_12376,N_11568,N_10661);
or U12377 (N_12377,N_11277,N_11724);
and U12378 (N_12378,N_11766,N_11073);
and U12379 (N_12379,N_11540,N_11715);
xor U12380 (N_12380,N_11517,N_10975);
nor U12381 (N_12381,N_10522,N_11651);
xor U12382 (N_12382,N_11064,N_11337);
nor U12383 (N_12383,N_11533,N_11772);
and U12384 (N_12384,N_11830,N_11705);
nand U12385 (N_12385,N_11045,N_10702);
nor U12386 (N_12386,N_11348,N_10805);
or U12387 (N_12387,N_11322,N_10698);
and U12388 (N_12388,N_11643,N_11655);
xor U12389 (N_12389,N_11823,N_11276);
or U12390 (N_12390,N_10624,N_11416);
xor U12391 (N_12391,N_10924,N_10959);
and U12392 (N_12392,N_11893,N_11428);
nand U12393 (N_12393,N_10537,N_11595);
nand U12394 (N_12394,N_11053,N_11713);
nor U12395 (N_12395,N_11611,N_10900);
nor U12396 (N_12396,N_10871,N_11059);
or U12397 (N_12397,N_10988,N_10726);
nand U12398 (N_12398,N_10840,N_11226);
or U12399 (N_12399,N_11552,N_11890);
xor U12400 (N_12400,N_11475,N_11635);
nor U12401 (N_12401,N_11626,N_11906);
nand U12402 (N_12402,N_11290,N_10774);
xnor U12403 (N_12403,N_10974,N_11817);
xor U12404 (N_12404,N_11021,N_11756);
or U12405 (N_12405,N_11271,N_11623);
nand U12406 (N_12406,N_11625,N_10932);
and U12407 (N_12407,N_11086,N_10876);
nand U12408 (N_12408,N_11132,N_11759);
or U12409 (N_12409,N_11180,N_10605);
nor U12410 (N_12410,N_10530,N_11962);
nand U12411 (N_12411,N_11903,N_11107);
and U12412 (N_12412,N_11807,N_11558);
xor U12413 (N_12413,N_11690,N_11163);
nand U12414 (N_12414,N_10573,N_11585);
nor U12415 (N_12415,N_11572,N_10922);
xor U12416 (N_12416,N_10711,N_11227);
nand U12417 (N_12417,N_11305,N_11865);
nor U12418 (N_12418,N_10682,N_11874);
or U12419 (N_12419,N_11821,N_10593);
nand U12420 (N_12420,N_10765,N_11314);
nand U12421 (N_12421,N_10510,N_11466);
nor U12422 (N_12422,N_10971,N_11604);
and U12423 (N_12423,N_10591,N_11061);
and U12424 (N_12424,N_11979,N_11231);
and U12425 (N_12425,N_10915,N_11843);
nor U12426 (N_12426,N_11233,N_11030);
or U12427 (N_12427,N_11569,N_10955);
xnor U12428 (N_12428,N_10898,N_10649);
nor U12429 (N_12429,N_10969,N_11718);
and U12430 (N_12430,N_11252,N_11733);
and U12431 (N_12431,N_10802,N_10574);
nand U12432 (N_12432,N_11575,N_11876);
or U12433 (N_12433,N_11573,N_10809);
nor U12434 (N_12434,N_10953,N_10566);
xnor U12435 (N_12435,N_11318,N_10651);
and U12436 (N_12436,N_10616,N_11899);
nor U12437 (N_12437,N_11642,N_10564);
nor U12438 (N_12438,N_11722,N_10535);
nor U12439 (N_12439,N_11972,N_10758);
or U12440 (N_12440,N_11089,N_11854);
nand U12441 (N_12441,N_11792,N_11846);
nor U12442 (N_12442,N_11514,N_10654);
nand U12443 (N_12443,N_10699,N_10869);
or U12444 (N_12444,N_11340,N_11028);
or U12445 (N_12445,N_11512,N_11027);
and U12446 (N_12446,N_11588,N_11424);
and U12447 (N_12447,N_10754,N_10554);
nor U12448 (N_12448,N_11702,N_10856);
and U12449 (N_12449,N_11935,N_11150);
or U12450 (N_12450,N_11989,N_10638);
nand U12451 (N_12451,N_10892,N_10784);
or U12452 (N_12452,N_11254,N_10732);
xnor U12453 (N_12453,N_10617,N_11678);
xor U12454 (N_12454,N_11036,N_11422);
and U12455 (N_12455,N_11805,N_11456);
xor U12456 (N_12456,N_11288,N_11038);
or U12457 (N_12457,N_11018,N_11997);
and U12458 (N_12458,N_10571,N_10601);
nor U12459 (N_12459,N_11229,N_10736);
nand U12460 (N_12460,N_10517,N_10595);
nand U12461 (N_12461,N_10796,N_11070);
nor U12462 (N_12462,N_10759,N_11199);
xnor U12463 (N_12463,N_11787,N_11206);
xor U12464 (N_12464,N_11904,N_11898);
nand U12465 (N_12465,N_11458,N_11519);
nand U12466 (N_12466,N_10810,N_10577);
nand U12467 (N_12467,N_10502,N_10780);
nand U12468 (N_12468,N_11050,N_11563);
xor U12469 (N_12469,N_11002,N_10507);
and U12470 (N_12470,N_11587,N_11605);
nand U12471 (N_12471,N_11417,N_11115);
nand U12472 (N_12472,N_10611,N_11232);
or U12473 (N_12473,N_11283,N_11836);
or U12474 (N_12474,N_10730,N_11936);
and U12475 (N_12475,N_11964,N_11238);
nor U12476 (N_12476,N_11311,N_11067);
or U12477 (N_12477,N_11795,N_10753);
nor U12478 (N_12478,N_11406,N_10667);
nand U12479 (N_12479,N_11958,N_10683);
nor U12480 (N_12480,N_11549,N_10910);
and U12481 (N_12481,N_11907,N_11886);
nor U12482 (N_12482,N_11395,N_10800);
nor U12483 (N_12483,N_10961,N_11268);
xor U12484 (N_12484,N_10613,N_11839);
and U12485 (N_12485,N_11620,N_11794);
nor U12486 (N_12486,N_11848,N_11162);
xnor U12487 (N_12487,N_11883,N_11755);
and U12488 (N_12488,N_11864,N_10901);
and U12489 (N_12489,N_11945,N_11462);
and U12490 (N_12490,N_11697,N_10946);
or U12491 (N_12491,N_11392,N_11869);
and U12492 (N_12492,N_10614,N_10925);
nand U12493 (N_12493,N_11481,N_11613);
and U12494 (N_12494,N_11215,N_10877);
and U12495 (N_12495,N_11513,N_10596);
nor U12496 (N_12496,N_11385,N_11364);
xor U12497 (N_12497,N_10536,N_10830);
and U12498 (N_12498,N_11102,N_11652);
or U12499 (N_12499,N_11202,N_11222);
nor U12500 (N_12500,N_10741,N_10714);
and U12501 (N_12501,N_10917,N_10615);
xnor U12502 (N_12502,N_11149,N_10828);
or U12503 (N_12503,N_10639,N_11007);
or U12504 (N_12504,N_11680,N_11892);
nand U12505 (N_12505,N_10920,N_11584);
nand U12506 (N_12506,N_11885,N_11248);
and U12507 (N_12507,N_11491,N_11078);
and U12508 (N_12508,N_10523,N_10972);
and U12509 (N_12509,N_10696,N_11631);
nor U12510 (N_12510,N_11433,N_11761);
xnor U12511 (N_12511,N_10627,N_11914);
and U12512 (N_12512,N_10722,N_11536);
nand U12513 (N_12513,N_11866,N_11365);
nand U12514 (N_12514,N_11287,N_11153);
nor U12515 (N_12515,N_11302,N_11455);
xor U12516 (N_12516,N_11096,N_11765);
nor U12517 (N_12517,N_10508,N_11369);
nand U12518 (N_12518,N_11716,N_10631);
nand U12519 (N_12519,N_11781,N_10844);
and U12520 (N_12520,N_11218,N_11535);
nand U12521 (N_12521,N_11230,N_10604);
nor U12522 (N_12522,N_10755,N_11138);
nor U12523 (N_12523,N_11988,N_11704);
or U12524 (N_12524,N_11122,N_11723);
nor U12525 (N_12525,N_10791,N_11111);
xnor U12526 (N_12526,N_10891,N_10771);
or U12527 (N_12527,N_10527,N_10609);
nand U12528 (N_12528,N_11435,N_11502);
or U12529 (N_12529,N_11926,N_10855);
xnor U12530 (N_12530,N_10673,N_11543);
nand U12531 (N_12531,N_11954,N_11414);
nand U12532 (N_12532,N_11917,N_10671);
nand U12533 (N_12533,N_10929,N_10576);
nand U12534 (N_12534,N_11204,N_11622);
nor U12535 (N_12535,N_11804,N_11280);
xnor U12536 (N_12536,N_11065,N_11745);
nand U12537 (N_12537,N_11299,N_10826);
xor U12538 (N_12538,N_11320,N_11197);
xnor U12539 (N_12539,N_11601,N_10904);
xor U12540 (N_12540,N_11090,N_11963);
or U12541 (N_12541,N_11060,N_10985);
or U12542 (N_12542,N_10528,N_11207);
xor U12543 (N_12543,N_11838,N_11380);
xor U12544 (N_12544,N_11501,N_11421);
nand U12545 (N_12545,N_11496,N_11859);
xnor U12546 (N_12546,N_11158,N_11195);
and U12547 (N_12547,N_10623,N_11367);
or U12548 (N_12548,N_11571,N_11043);
xor U12549 (N_12549,N_11703,N_11734);
nand U12550 (N_12550,N_11827,N_11712);
or U12551 (N_12551,N_11852,N_11596);
nand U12552 (N_12552,N_11315,N_10880);
xor U12553 (N_12553,N_10845,N_10822);
xor U12554 (N_12554,N_11672,N_11022);
nor U12555 (N_12555,N_11976,N_11679);
and U12556 (N_12556,N_10556,N_11387);
nor U12557 (N_12557,N_11083,N_10747);
and U12558 (N_12558,N_11599,N_11557);
nor U12559 (N_12559,N_10788,N_10672);
xor U12560 (N_12560,N_10749,N_11079);
or U12561 (N_12561,N_11259,N_10835);
or U12562 (N_12562,N_10704,N_11891);
nor U12563 (N_12563,N_10841,N_11448);
nand U12564 (N_12564,N_11532,N_11789);
nor U12565 (N_12565,N_11411,N_10675);
and U12566 (N_12566,N_11451,N_10906);
and U12567 (N_12567,N_11332,N_11996);
and U12568 (N_12568,N_11731,N_11873);
nand U12569 (N_12569,N_11253,N_11551);
nand U12570 (N_12570,N_11768,N_11674);
and U12571 (N_12571,N_10764,N_11511);
nor U12572 (N_12572,N_11173,N_10926);
and U12573 (N_12573,N_10743,N_11548);
nand U12574 (N_12574,N_10670,N_10580);
xor U12575 (N_12575,N_11779,N_10626);
nor U12576 (N_12576,N_11960,N_11068);
nor U12577 (N_12577,N_11476,N_11683);
and U12578 (N_12578,N_11984,N_11243);
nor U12579 (N_12579,N_11074,N_10966);
nand U12580 (N_12580,N_11614,N_11000);
nand U12581 (N_12581,N_11350,N_10798);
and U12582 (N_12582,N_11771,N_10989);
and U12583 (N_12583,N_11881,N_10982);
nand U12584 (N_12584,N_10986,N_11629);
xnor U12585 (N_12585,N_11172,N_11661);
nand U12586 (N_12586,N_10752,N_11922);
nand U12587 (N_12587,N_11565,N_10636);
nand U12588 (N_12588,N_11190,N_11339);
nor U12589 (N_12589,N_10803,N_11902);
and U12590 (N_12590,N_11234,N_11136);
and U12591 (N_12591,N_10937,N_10861);
nand U12592 (N_12592,N_10979,N_10618);
or U12593 (N_12593,N_10555,N_10949);
nor U12594 (N_12594,N_11763,N_10952);
nor U12595 (N_12595,N_11014,N_11797);
or U12596 (N_12596,N_10715,N_10757);
nor U12597 (N_12597,N_10867,N_10909);
or U12598 (N_12598,N_11542,N_10862);
xor U12599 (N_12599,N_10962,N_11473);
xor U12600 (N_12600,N_11391,N_10742);
xnor U12601 (N_12601,N_10950,N_10987);
and U12602 (N_12602,N_10847,N_10970);
xor U12603 (N_12603,N_11537,N_11673);
xnor U12604 (N_12604,N_11477,N_11442);
xor U12605 (N_12605,N_11676,N_11470);
xor U12606 (N_12606,N_11600,N_11770);
nand U12607 (N_12607,N_10684,N_11210);
nand U12608 (N_12608,N_10567,N_11317);
xor U12609 (N_12609,N_11378,N_10834);
nor U12610 (N_12610,N_11653,N_10995);
nand U12611 (N_12611,N_10553,N_10923);
nand U12612 (N_12612,N_10657,N_11800);
nor U12613 (N_12613,N_11639,N_10884);
nor U12614 (N_12614,N_11554,N_11054);
xnor U12615 (N_12615,N_10964,N_11052);
or U12616 (N_12616,N_11577,N_11744);
nand U12617 (N_12617,N_11347,N_11032);
nand U12618 (N_12618,N_11822,N_11923);
or U12619 (N_12619,N_10515,N_11919);
or U12620 (N_12620,N_11884,N_11457);
and U12621 (N_12621,N_11303,N_11076);
nand U12622 (N_12622,N_11528,N_11338);
nor U12623 (N_12623,N_10895,N_10882);
nand U12624 (N_12624,N_11292,N_10692);
nor U12625 (N_12625,N_11980,N_10738);
nand U12626 (N_12626,N_11833,N_11937);
or U12627 (N_12627,N_11981,N_10997);
nor U12628 (N_12628,N_11194,N_10849);
and U12629 (N_12629,N_11932,N_11189);
and U12630 (N_12630,N_11275,N_10689);
or U12631 (N_12631,N_10998,N_10858);
nor U12632 (N_12632,N_11269,N_10723);
nor U12633 (N_12633,N_11498,N_11214);
and U12634 (N_12634,N_11582,N_10919);
or U12635 (N_12635,N_11934,N_10606);
xor U12636 (N_12636,N_10658,N_11732);
and U12637 (N_12637,N_11282,N_11009);
xor U12638 (N_12638,N_11941,N_11844);
nor U12639 (N_12639,N_10635,N_11499);
nand U12640 (N_12640,N_11213,N_11814);
xor U12641 (N_12641,N_11505,N_11125);
nor U12642 (N_12642,N_10930,N_11877);
xnor U12643 (N_12643,N_11463,N_11688);
and U12644 (N_12644,N_11965,N_11961);
nor U12645 (N_12645,N_11990,N_11518);
nand U12646 (N_12646,N_11263,N_11097);
and U12647 (N_12647,N_10740,N_10748);
and U12648 (N_12648,N_10646,N_11621);
nor U12649 (N_12649,N_10703,N_10628);
xor U12650 (N_12650,N_11858,N_11419);
and U12651 (N_12651,N_10843,N_11545);
or U12652 (N_12652,N_11051,N_11693);
xnor U12653 (N_12653,N_11445,N_10902);
nor U12654 (N_12654,N_10815,N_11345);
nand U12655 (N_12655,N_11918,N_10813);
or U12656 (N_12656,N_11447,N_11529);
nand U12657 (N_12657,N_11294,N_11209);
or U12658 (N_12658,N_11685,N_10819);
nor U12659 (N_12659,N_10806,N_11255);
xnor U12660 (N_12660,N_10729,N_11141);
nor U12661 (N_12661,N_11106,N_10700);
xnor U12662 (N_12662,N_11947,N_11497);
nor U12663 (N_12663,N_11523,N_11658);
nand U12664 (N_12664,N_11644,N_10875);
nand U12665 (N_12665,N_11384,N_10801);
and U12666 (N_12666,N_10666,N_10669);
and U12667 (N_12667,N_11001,N_11010);
or U12668 (N_12668,N_11782,N_11430);
nand U12669 (N_12669,N_11383,N_11748);
nor U12670 (N_12670,N_11566,N_11047);
xnor U12671 (N_12671,N_11203,N_11598);
or U12672 (N_12672,N_11632,N_10933);
xnor U12673 (N_12673,N_11121,N_10674);
or U12674 (N_12674,N_11323,N_10978);
xor U12675 (N_12675,N_11409,N_11080);
nand U12676 (N_12676,N_11974,N_11266);
xor U12677 (N_12677,N_10503,N_11570);
nand U12678 (N_12678,N_10587,N_11398);
nor U12679 (N_12679,N_10790,N_11039);
nand U12680 (N_12680,N_11507,N_10837);
nand U12681 (N_12681,N_10761,N_11967);
xnor U12682 (N_12682,N_10685,N_11404);
or U12683 (N_12683,N_11011,N_10559);
and U12684 (N_12684,N_10514,N_11769);
nand U12685 (N_12685,N_11857,N_11832);
or U12686 (N_12686,N_11432,N_11335);
or U12687 (N_12687,N_11969,N_11058);
nand U12688 (N_12688,N_11949,N_11762);
xor U12689 (N_12689,N_10816,N_11952);
xor U12690 (N_12690,N_11815,N_10526);
nand U12691 (N_12691,N_11708,N_11174);
nand U12692 (N_12692,N_10637,N_11334);
nand U12693 (N_12693,N_11615,N_10940);
nor U12694 (N_12694,N_10838,N_11237);
nor U12695 (N_12695,N_10727,N_11026);
nor U12696 (N_12696,N_11646,N_10734);
nand U12697 (N_12697,N_11033,N_11546);
xnor U12698 (N_12698,N_11911,N_11930);
nand U12699 (N_12699,N_11041,N_10690);
xnor U12700 (N_12700,N_11081,N_11358);
nand U12701 (N_12701,N_11521,N_11471);
xor U12702 (N_12702,N_11217,N_11192);
nor U12703 (N_12703,N_11849,N_11579);
xor U12704 (N_12704,N_10718,N_10865);
and U12705 (N_12705,N_11752,N_10750);
xnor U12706 (N_12706,N_11808,N_11240);
and U12707 (N_12707,N_11370,N_10531);
or U12708 (N_12708,N_11357,N_11793);
xor U12709 (N_12709,N_11553,N_11042);
nor U12710 (N_12710,N_10647,N_10859);
nand U12711 (N_12711,N_11221,N_11094);
or U12712 (N_12712,N_11791,N_11492);
nor U12713 (N_12713,N_11179,N_11143);
nand U12714 (N_12714,N_11046,N_10653);
and U12715 (N_12715,N_10594,N_11660);
nor U12716 (N_12716,N_11446,N_11581);
and U12717 (N_12717,N_11100,N_11913);
or U12718 (N_12718,N_11131,N_11152);
or U12719 (N_12719,N_10512,N_11224);
and U12720 (N_12720,N_11401,N_11164);
xor U12721 (N_12721,N_10717,N_11072);
and U12722 (N_12722,N_10846,N_11225);
xor U12723 (N_12723,N_11397,N_10501);
nand U12724 (N_12724,N_10620,N_11472);
xnor U12725 (N_12725,N_10731,N_10548);
and U12726 (N_12726,N_11425,N_10600);
or U12727 (N_12727,N_11055,N_10957);
nand U12728 (N_12728,N_11123,N_11686);
nand U12729 (N_12729,N_11104,N_10927);
nand U12730 (N_12730,N_10660,N_11627);
xnor U12731 (N_12731,N_10864,N_10795);
xnor U12732 (N_12732,N_11509,N_11485);
nand U12733 (N_12733,N_10918,N_10874);
and U12734 (N_12734,N_11561,N_10994);
and U12735 (N_12735,N_10947,N_11735);
and U12736 (N_12736,N_11091,N_10829);
and U12737 (N_12737,N_11327,N_11847);
nor U12738 (N_12738,N_11780,N_11973);
xnor U12739 (N_12739,N_11662,N_11436);
or U12740 (N_12740,N_11648,N_11105);
nor U12741 (N_12741,N_11130,N_11707);
nor U12742 (N_12742,N_10797,N_11527);
xnor U12743 (N_12743,N_11530,N_11031);
and U12744 (N_12744,N_10532,N_10545);
nand U12745 (N_12745,N_10716,N_11377);
or U12746 (N_12746,N_11983,N_11183);
or U12747 (N_12747,N_11758,N_11966);
nor U12748 (N_12748,N_11878,N_10833);
xor U12749 (N_12749,N_11326,N_11616);
nor U12750 (N_12750,N_10522,N_11681);
xnor U12751 (N_12751,N_10680,N_10569);
or U12752 (N_12752,N_10549,N_11972);
nand U12753 (N_12753,N_10857,N_11654);
and U12754 (N_12754,N_10996,N_10527);
or U12755 (N_12755,N_10965,N_11525);
and U12756 (N_12756,N_11414,N_11206);
nand U12757 (N_12757,N_11367,N_11861);
or U12758 (N_12758,N_11263,N_11264);
nor U12759 (N_12759,N_11594,N_11174);
nand U12760 (N_12760,N_11633,N_11129);
or U12761 (N_12761,N_10942,N_10912);
nor U12762 (N_12762,N_11913,N_11715);
xor U12763 (N_12763,N_11177,N_11099);
nand U12764 (N_12764,N_10839,N_11733);
nand U12765 (N_12765,N_11716,N_11993);
or U12766 (N_12766,N_11707,N_11788);
or U12767 (N_12767,N_11493,N_11723);
xor U12768 (N_12768,N_11574,N_11673);
nand U12769 (N_12769,N_11914,N_10626);
and U12770 (N_12770,N_11174,N_10677);
nor U12771 (N_12771,N_11657,N_10687);
nor U12772 (N_12772,N_11793,N_11147);
nand U12773 (N_12773,N_11810,N_10738);
and U12774 (N_12774,N_11687,N_10662);
and U12775 (N_12775,N_10993,N_11723);
or U12776 (N_12776,N_11787,N_11724);
and U12777 (N_12777,N_11525,N_11371);
nor U12778 (N_12778,N_11957,N_11888);
xnor U12779 (N_12779,N_11045,N_11474);
nor U12780 (N_12780,N_10900,N_11415);
xor U12781 (N_12781,N_11167,N_11763);
and U12782 (N_12782,N_11446,N_10651);
nand U12783 (N_12783,N_11541,N_10595);
or U12784 (N_12784,N_11369,N_11086);
xor U12785 (N_12785,N_11841,N_10760);
nand U12786 (N_12786,N_11497,N_11892);
nand U12787 (N_12787,N_10780,N_11566);
nor U12788 (N_12788,N_10775,N_10734);
and U12789 (N_12789,N_10994,N_10678);
and U12790 (N_12790,N_11010,N_10828);
or U12791 (N_12791,N_10593,N_10503);
xnor U12792 (N_12792,N_11372,N_10513);
or U12793 (N_12793,N_11512,N_11727);
xor U12794 (N_12794,N_11994,N_11073);
nor U12795 (N_12795,N_11716,N_10536);
or U12796 (N_12796,N_11845,N_10796);
and U12797 (N_12797,N_10538,N_11901);
nand U12798 (N_12798,N_10936,N_10778);
or U12799 (N_12799,N_11708,N_11016);
or U12800 (N_12800,N_11682,N_11721);
nor U12801 (N_12801,N_11700,N_10579);
nor U12802 (N_12802,N_11757,N_10600);
nand U12803 (N_12803,N_11667,N_11923);
nand U12804 (N_12804,N_11491,N_11424);
and U12805 (N_12805,N_10579,N_11774);
or U12806 (N_12806,N_11675,N_10614);
and U12807 (N_12807,N_10622,N_11641);
xor U12808 (N_12808,N_11256,N_11020);
and U12809 (N_12809,N_11694,N_10555);
xnor U12810 (N_12810,N_11148,N_11958);
nor U12811 (N_12811,N_11776,N_10717);
xnor U12812 (N_12812,N_11687,N_10944);
or U12813 (N_12813,N_10794,N_11076);
xor U12814 (N_12814,N_11980,N_11717);
and U12815 (N_12815,N_11873,N_11176);
nor U12816 (N_12816,N_11023,N_11755);
xnor U12817 (N_12817,N_11116,N_11543);
nor U12818 (N_12818,N_10986,N_11122);
nor U12819 (N_12819,N_11818,N_10969);
nand U12820 (N_12820,N_10731,N_11164);
or U12821 (N_12821,N_11544,N_11163);
nor U12822 (N_12822,N_10765,N_10988);
and U12823 (N_12823,N_11674,N_10649);
or U12824 (N_12824,N_11766,N_10943);
nand U12825 (N_12825,N_11894,N_11522);
and U12826 (N_12826,N_11629,N_10831);
and U12827 (N_12827,N_10565,N_11796);
and U12828 (N_12828,N_10760,N_11829);
nor U12829 (N_12829,N_10970,N_11444);
nor U12830 (N_12830,N_10868,N_11907);
nand U12831 (N_12831,N_11588,N_10752);
xnor U12832 (N_12832,N_11213,N_11500);
nor U12833 (N_12833,N_11716,N_11741);
and U12834 (N_12834,N_11977,N_10753);
nor U12835 (N_12835,N_11740,N_11678);
or U12836 (N_12836,N_11058,N_11047);
nand U12837 (N_12837,N_10524,N_10780);
and U12838 (N_12838,N_11838,N_11552);
nand U12839 (N_12839,N_11406,N_11626);
and U12840 (N_12840,N_11576,N_11306);
or U12841 (N_12841,N_10756,N_10526);
nand U12842 (N_12842,N_11062,N_11637);
nand U12843 (N_12843,N_11290,N_11046);
nor U12844 (N_12844,N_11348,N_11532);
xor U12845 (N_12845,N_11130,N_11922);
nand U12846 (N_12846,N_10750,N_11193);
and U12847 (N_12847,N_10922,N_11812);
or U12848 (N_12848,N_11567,N_11168);
nand U12849 (N_12849,N_11869,N_11347);
xor U12850 (N_12850,N_10820,N_11694);
nand U12851 (N_12851,N_11091,N_11728);
xor U12852 (N_12852,N_11278,N_10746);
and U12853 (N_12853,N_10707,N_11650);
nand U12854 (N_12854,N_11737,N_10613);
and U12855 (N_12855,N_11551,N_11811);
and U12856 (N_12856,N_11881,N_10918);
nand U12857 (N_12857,N_10569,N_11393);
nor U12858 (N_12858,N_11116,N_11916);
and U12859 (N_12859,N_11597,N_10996);
nor U12860 (N_12860,N_10547,N_10877);
nand U12861 (N_12861,N_10933,N_11744);
nand U12862 (N_12862,N_11007,N_11527);
and U12863 (N_12863,N_11334,N_11986);
xor U12864 (N_12864,N_11820,N_11233);
nor U12865 (N_12865,N_11947,N_11438);
nand U12866 (N_12866,N_11365,N_11454);
or U12867 (N_12867,N_11974,N_11219);
xnor U12868 (N_12868,N_11995,N_11358);
xor U12869 (N_12869,N_11977,N_11663);
nor U12870 (N_12870,N_11478,N_10649);
nor U12871 (N_12871,N_11785,N_10893);
or U12872 (N_12872,N_11123,N_11159);
nand U12873 (N_12873,N_10909,N_11616);
nand U12874 (N_12874,N_11239,N_11800);
and U12875 (N_12875,N_11833,N_10832);
nand U12876 (N_12876,N_11622,N_11107);
or U12877 (N_12877,N_10902,N_11049);
and U12878 (N_12878,N_10587,N_10765);
xor U12879 (N_12879,N_11355,N_11268);
xor U12880 (N_12880,N_10556,N_11528);
nand U12881 (N_12881,N_11101,N_11832);
and U12882 (N_12882,N_11226,N_11512);
or U12883 (N_12883,N_10833,N_10763);
and U12884 (N_12884,N_11869,N_11664);
nor U12885 (N_12885,N_10503,N_10876);
nand U12886 (N_12886,N_10548,N_11477);
and U12887 (N_12887,N_11620,N_10950);
or U12888 (N_12888,N_11912,N_11838);
nand U12889 (N_12889,N_11296,N_11856);
and U12890 (N_12890,N_11260,N_10982);
and U12891 (N_12891,N_11025,N_11311);
nand U12892 (N_12892,N_11811,N_10858);
nand U12893 (N_12893,N_11890,N_10583);
xor U12894 (N_12894,N_11746,N_11184);
and U12895 (N_12895,N_11651,N_11905);
xnor U12896 (N_12896,N_10839,N_11721);
and U12897 (N_12897,N_11708,N_10988);
and U12898 (N_12898,N_11657,N_10503);
nand U12899 (N_12899,N_11429,N_11417);
and U12900 (N_12900,N_11168,N_10655);
nor U12901 (N_12901,N_11725,N_11839);
nor U12902 (N_12902,N_11561,N_11452);
nand U12903 (N_12903,N_11964,N_10621);
and U12904 (N_12904,N_11110,N_10933);
or U12905 (N_12905,N_10506,N_11950);
nor U12906 (N_12906,N_11993,N_11357);
xor U12907 (N_12907,N_10862,N_11467);
and U12908 (N_12908,N_11916,N_11106);
xor U12909 (N_12909,N_11936,N_10716);
or U12910 (N_12910,N_10692,N_10541);
and U12911 (N_12911,N_11088,N_11952);
or U12912 (N_12912,N_11568,N_11956);
or U12913 (N_12913,N_10729,N_11405);
and U12914 (N_12914,N_10509,N_11365);
or U12915 (N_12915,N_10925,N_10517);
nand U12916 (N_12916,N_11059,N_10559);
nand U12917 (N_12917,N_11063,N_11288);
xor U12918 (N_12918,N_11276,N_11831);
and U12919 (N_12919,N_10789,N_10956);
or U12920 (N_12920,N_10825,N_10804);
or U12921 (N_12921,N_10806,N_11745);
or U12922 (N_12922,N_11505,N_11528);
or U12923 (N_12923,N_10859,N_10932);
or U12924 (N_12924,N_11797,N_10544);
xor U12925 (N_12925,N_11828,N_11321);
and U12926 (N_12926,N_10904,N_11577);
and U12927 (N_12927,N_10729,N_11281);
nand U12928 (N_12928,N_10852,N_11582);
xor U12929 (N_12929,N_11845,N_11960);
xnor U12930 (N_12930,N_11537,N_10527);
nand U12931 (N_12931,N_11342,N_11119);
and U12932 (N_12932,N_10549,N_11048);
xnor U12933 (N_12933,N_10859,N_11395);
and U12934 (N_12934,N_10592,N_11234);
and U12935 (N_12935,N_10660,N_11332);
xnor U12936 (N_12936,N_11537,N_11298);
and U12937 (N_12937,N_11027,N_10583);
nor U12938 (N_12938,N_11414,N_10847);
xnor U12939 (N_12939,N_11081,N_10639);
nand U12940 (N_12940,N_10871,N_11763);
nand U12941 (N_12941,N_10764,N_11378);
or U12942 (N_12942,N_11065,N_10945);
nand U12943 (N_12943,N_11564,N_10567);
and U12944 (N_12944,N_11801,N_11298);
and U12945 (N_12945,N_11772,N_11302);
nand U12946 (N_12946,N_10827,N_10999);
or U12947 (N_12947,N_11618,N_11004);
xnor U12948 (N_12948,N_10957,N_11944);
xnor U12949 (N_12949,N_10624,N_11392);
xnor U12950 (N_12950,N_11211,N_11128);
nor U12951 (N_12951,N_11436,N_10610);
or U12952 (N_12952,N_11461,N_10878);
nand U12953 (N_12953,N_10618,N_11961);
xor U12954 (N_12954,N_11298,N_10912);
and U12955 (N_12955,N_11857,N_11148);
nand U12956 (N_12956,N_10841,N_11685);
and U12957 (N_12957,N_10984,N_10634);
or U12958 (N_12958,N_11149,N_11359);
nand U12959 (N_12959,N_11514,N_10870);
and U12960 (N_12960,N_10736,N_10876);
or U12961 (N_12961,N_10528,N_11507);
nor U12962 (N_12962,N_11090,N_10711);
nand U12963 (N_12963,N_11025,N_10969);
nor U12964 (N_12964,N_10740,N_10864);
nor U12965 (N_12965,N_11802,N_10610);
xnor U12966 (N_12966,N_11384,N_11895);
nor U12967 (N_12967,N_10501,N_11069);
nand U12968 (N_12968,N_10610,N_11194);
or U12969 (N_12969,N_11176,N_11336);
nor U12970 (N_12970,N_11755,N_11467);
nand U12971 (N_12971,N_11564,N_11616);
xor U12972 (N_12972,N_11274,N_11501);
nand U12973 (N_12973,N_11370,N_11150);
xor U12974 (N_12974,N_11402,N_11836);
nor U12975 (N_12975,N_11396,N_10687);
nand U12976 (N_12976,N_11132,N_11615);
and U12977 (N_12977,N_10944,N_11664);
nor U12978 (N_12978,N_10578,N_10615);
nor U12979 (N_12979,N_11317,N_11718);
xnor U12980 (N_12980,N_11824,N_10836);
xor U12981 (N_12981,N_11091,N_10962);
and U12982 (N_12982,N_10871,N_10875);
or U12983 (N_12983,N_11230,N_11024);
nand U12984 (N_12984,N_11995,N_10822);
or U12985 (N_12985,N_10933,N_11197);
or U12986 (N_12986,N_11555,N_11405);
xnor U12987 (N_12987,N_10971,N_10781);
or U12988 (N_12988,N_11091,N_10606);
xor U12989 (N_12989,N_10946,N_11294);
nand U12990 (N_12990,N_11583,N_10554);
or U12991 (N_12991,N_11621,N_11122);
nor U12992 (N_12992,N_11598,N_10975);
or U12993 (N_12993,N_10535,N_11459);
nor U12994 (N_12994,N_11571,N_11388);
xor U12995 (N_12995,N_10663,N_10804);
xor U12996 (N_12996,N_11942,N_11159);
and U12997 (N_12997,N_11792,N_11693);
nand U12998 (N_12998,N_11913,N_11388);
or U12999 (N_12999,N_10812,N_10531);
or U13000 (N_13000,N_11189,N_11744);
nor U13001 (N_13001,N_11071,N_11815);
nor U13002 (N_13002,N_11716,N_10604);
nor U13003 (N_13003,N_11436,N_11279);
nor U13004 (N_13004,N_11088,N_11126);
or U13005 (N_13005,N_11724,N_10844);
or U13006 (N_13006,N_11685,N_10690);
xnor U13007 (N_13007,N_11153,N_10847);
and U13008 (N_13008,N_11631,N_11627);
nor U13009 (N_13009,N_11367,N_11535);
or U13010 (N_13010,N_11062,N_11561);
xor U13011 (N_13011,N_11097,N_11468);
and U13012 (N_13012,N_10853,N_11229);
and U13013 (N_13013,N_11117,N_10762);
nand U13014 (N_13014,N_11218,N_11069);
nor U13015 (N_13015,N_11746,N_10979);
nand U13016 (N_13016,N_11282,N_11123);
nor U13017 (N_13017,N_10750,N_11456);
xnor U13018 (N_13018,N_11688,N_11018);
nand U13019 (N_13019,N_11026,N_11286);
nor U13020 (N_13020,N_10748,N_11627);
and U13021 (N_13021,N_11342,N_11889);
xnor U13022 (N_13022,N_11049,N_10866);
xor U13023 (N_13023,N_11549,N_10625);
xnor U13024 (N_13024,N_11886,N_10543);
xnor U13025 (N_13025,N_10993,N_10616);
xor U13026 (N_13026,N_11544,N_11915);
xor U13027 (N_13027,N_11445,N_10921);
nand U13028 (N_13028,N_10684,N_11299);
and U13029 (N_13029,N_10797,N_10864);
nor U13030 (N_13030,N_11514,N_11244);
or U13031 (N_13031,N_11996,N_10933);
nand U13032 (N_13032,N_10874,N_10710);
and U13033 (N_13033,N_10886,N_11129);
xor U13034 (N_13034,N_11326,N_10735);
and U13035 (N_13035,N_11135,N_11304);
and U13036 (N_13036,N_11333,N_11805);
nand U13037 (N_13037,N_11236,N_11771);
and U13038 (N_13038,N_10705,N_11143);
or U13039 (N_13039,N_11054,N_11981);
nand U13040 (N_13040,N_11850,N_11346);
and U13041 (N_13041,N_11292,N_11583);
and U13042 (N_13042,N_11013,N_10756);
and U13043 (N_13043,N_11029,N_11129);
nor U13044 (N_13044,N_11562,N_10824);
xor U13045 (N_13045,N_10969,N_10728);
xor U13046 (N_13046,N_10638,N_11797);
nor U13047 (N_13047,N_11298,N_11277);
nand U13048 (N_13048,N_10962,N_11366);
xor U13049 (N_13049,N_11251,N_11538);
nor U13050 (N_13050,N_10605,N_11537);
xnor U13051 (N_13051,N_11898,N_11835);
nor U13052 (N_13052,N_11462,N_11022);
nand U13053 (N_13053,N_10696,N_10581);
and U13054 (N_13054,N_11448,N_11402);
xnor U13055 (N_13055,N_11671,N_10612);
xor U13056 (N_13056,N_11630,N_11442);
or U13057 (N_13057,N_11459,N_11706);
nand U13058 (N_13058,N_10760,N_11501);
nor U13059 (N_13059,N_11577,N_10738);
or U13060 (N_13060,N_11091,N_10887);
nor U13061 (N_13061,N_11092,N_11132);
nor U13062 (N_13062,N_11651,N_10585);
or U13063 (N_13063,N_11417,N_11086);
nand U13064 (N_13064,N_10874,N_11430);
nor U13065 (N_13065,N_10945,N_11553);
nand U13066 (N_13066,N_11405,N_11306);
nand U13067 (N_13067,N_11246,N_10515);
and U13068 (N_13068,N_11776,N_11656);
nand U13069 (N_13069,N_11663,N_10951);
nor U13070 (N_13070,N_11544,N_11088);
nand U13071 (N_13071,N_11121,N_11989);
xor U13072 (N_13072,N_11998,N_11675);
and U13073 (N_13073,N_11193,N_11925);
or U13074 (N_13074,N_11636,N_10683);
xor U13075 (N_13075,N_11960,N_11738);
nor U13076 (N_13076,N_11872,N_11501);
or U13077 (N_13077,N_11507,N_11875);
nand U13078 (N_13078,N_10932,N_11800);
or U13079 (N_13079,N_11965,N_11648);
xor U13080 (N_13080,N_11735,N_11104);
or U13081 (N_13081,N_11440,N_10520);
xor U13082 (N_13082,N_11143,N_10593);
nand U13083 (N_13083,N_10585,N_11488);
and U13084 (N_13084,N_10608,N_11344);
and U13085 (N_13085,N_10821,N_10932);
nor U13086 (N_13086,N_10963,N_11252);
nor U13087 (N_13087,N_10964,N_10940);
and U13088 (N_13088,N_11234,N_11025);
nand U13089 (N_13089,N_11105,N_11486);
nor U13090 (N_13090,N_11225,N_11763);
and U13091 (N_13091,N_11813,N_11224);
xnor U13092 (N_13092,N_11790,N_10706);
and U13093 (N_13093,N_11109,N_11583);
nand U13094 (N_13094,N_11474,N_10546);
and U13095 (N_13095,N_11223,N_11439);
nor U13096 (N_13096,N_11607,N_10638);
nor U13097 (N_13097,N_10970,N_11671);
xnor U13098 (N_13098,N_11378,N_11352);
or U13099 (N_13099,N_10951,N_10801);
nand U13100 (N_13100,N_11381,N_10877);
and U13101 (N_13101,N_11598,N_10853);
nor U13102 (N_13102,N_10802,N_11718);
nor U13103 (N_13103,N_11523,N_11577);
nor U13104 (N_13104,N_11175,N_11674);
nand U13105 (N_13105,N_11201,N_10621);
and U13106 (N_13106,N_11841,N_11531);
or U13107 (N_13107,N_11274,N_11512);
and U13108 (N_13108,N_11823,N_10663);
or U13109 (N_13109,N_11277,N_11213);
xor U13110 (N_13110,N_10881,N_11333);
and U13111 (N_13111,N_11838,N_10528);
nand U13112 (N_13112,N_10890,N_10841);
nand U13113 (N_13113,N_10979,N_11894);
and U13114 (N_13114,N_11381,N_11170);
and U13115 (N_13115,N_11506,N_10689);
and U13116 (N_13116,N_11582,N_11929);
nor U13117 (N_13117,N_11911,N_10702);
nand U13118 (N_13118,N_10977,N_11743);
or U13119 (N_13119,N_11131,N_11635);
xnor U13120 (N_13120,N_10884,N_11494);
nand U13121 (N_13121,N_11851,N_11042);
and U13122 (N_13122,N_11794,N_11813);
xor U13123 (N_13123,N_11873,N_11076);
nor U13124 (N_13124,N_11164,N_11171);
nor U13125 (N_13125,N_11042,N_10697);
nor U13126 (N_13126,N_10632,N_10874);
nor U13127 (N_13127,N_11296,N_10594);
xor U13128 (N_13128,N_11055,N_11854);
xor U13129 (N_13129,N_11473,N_11426);
nand U13130 (N_13130,N_11546,N_10854);
or U13131 (N_13131,N_10908,N_11427);
xor U13132 (N_13132,N_11680,N_11905);
and U13133 (N_13133,N_11891,N_11734);
xnor U13134 (N_13134,N_11121,N_11637);
nor U13135 (N_13135,N_10773,N_11383);
and U13136 (N_13136,N_11127,N_10903);
or U13137 (N_13137,N_10963,N_11058);
or U13138 (N_13138,N_11611,N_11343);
xor U13139 (N_13139,N_10937,N_11050);
and U13140 (N_13140,N_10906,N_10755);
nand U13141 (N_13141,N_11751,N_11502);
and U13142 (N_13142,N_11231,N_11312);
and U13143 (N_13143,N_10999,N_10728);
nor U13144 (N_13144,N_10860,N_10582);
nand U13145 (N_13145,N_11601,N_11565);
or U13146 (N_13146,N_10773,N_11054);
xnor U13147 (N_13147,N_11243,N_11235);
and U13148 (N_13148,N_10867,N_11535);
xor U13149 (N_13149,N_11764,N_11856);
and U13150 (N_13150,N_11608,N_10884);
nand U13151 (N_13151,N_11732,N_11694);
xnor U13152 (N_13152,N_11971,N_10677);
xor U13153 (N_13153,N_11577,N_10889);
or U13154 (N_13154,N_11459,N_11892);
nor U13155 (N_13155,N_10736,N_11268);
xor U13156 (N_13156,N_11505,N_10973);
nor U13157 (N_13157,N_11329,N_11416);
nand U13158 (N_13158,N_11791,N_11314);
nand U13159 (N_13159,N_11727,N_11990);
or U13160 (N_13160,N_10545,N_11035);
xnor U13161 (N_13161,N_11989,N_11421);
xor U13162 (N_13162,N_11243,N_11629);
nand U13163 (N_13163,N_11789,N_11818);
or U13164 (N_13164,N_11809,N_11511);
xor U13165 (N_13165,N_11208,N_10546);
xnor U13166 (N_13166,N_11475,N_11208);
nor U13167 (N_13167,N_10697,N_11794);
nor U13168 (N_13168,N_10597,N_11548);
and U13169 (N_13169,N_11180,N_11936);
or U13170 (N_13170,N_11966,N_11231);
xor U13171 (N_13171,N_11070,N_11996);
or U13172 (N_13172,N_11500,N_11764);
xnor U13173 (N_13173,N_10688,N_11389);
nor U13174 (N_13174,N_11625,N_11733);
or U13175 (N_13175,N_10719,N_11949);
and U13176 (N_13176,N_10832,N_10708);
nand U13177 (N_13177,N_11692,N_11626);
and U13178 (N_13178,N_11167,N_11967);
xor U13179 (N_13179,N_11801,N_11085);
xnor U13180 (N_13180,N_10962,N_11879);
nor U13181 (N_13181,N_11890,N_11478);
or U13182 (N_13182,N_10994,N_11814);
nor U13183 (N_13183,N_11879,N_11910);
xor U13184 (N_13184,N_11001,N_11285);
nor U13185 (N_13185,N_11198,N_11728);
nor U13186 (N_13186,N_11355,N_11325);
and U13187 (N_13187,N_11943,N_10638);
and U13188 (N_13188,N_10860,N_10720);
or U13189 (N_13189,N_11564,N_11950);
or U13190 (N_13190,N_10870,N_11186);
xnor U13191 (N_13191,N_11671,N_11913);
and U13192 (N_13192,N_11673,N_11155);
nand U13193 (N_13193,N_11872,N_11424);
nand U13194 (N_13194,N_10509,N_11395);
nand U13195 (N_13195,N_10817,N_10831);
nand U13196 (N_13196,N_11382,N_10953);
xor U13197 (N_13197,N_10530,N_10991);
and U13198 (N_13198,N_11490,N_11224);
xnor U13199 (N_13199,N_11385,N_11594);
nand U13200 (N_13200,N_11675,N_10864);
and U13201 (N_13201,N_11234,N_11265);
nor U13202 (N_13202,N_10553,N_11704);
and U13203 (N_13203,N_11393,N_10505);
nor U13204 (N_13204,N_11817,N_10669);
or U13205 (N_13205,N_10610,N_10973);
nand U13206 (N_13206,N_10892,N_11423);
or U13207 (N_13207,N_10902,N_11518);
and U13208 (N_13208,N_10764,N_10798);
and U13209 (N_13209,N_10862,N_10526);
and U13210 (N_13210,N_10659,N_11502);
and U13211 (N_13211,N_11968,N_11706);
or U13212 (N_13212,N_11244,N_10683);
nand U13213 (N_13213,N_10728,N_11325);
nand U13214 (N_13214,N_11723,N_10780);
and U13215 (N_13215,N_11044,N_10957);
nor U13216 (N_13216,N_10840,N_11361);
and U13217 (N_13217,N_10778,N_11922);
nor U13218 (N_13218,N_10650,N_10647);
nand U13219 (N_13219,N_10939,N_11744);
xnor U13220 (N_13220,N_11416,N_11783);
nand U13221 (N_13221,N_11698,N_11586);
and U13222 (N_13222,N_11708,N_11633);
nand U13223 (N_13223,N_11674,N_11399);
xnor U13224 (N_13224,N_10567,N_10903);
xor U13225 (N_13225,N_11464,N_10781);
nor U13226 (N_13226,N_11772,N_11551);
or U13227 (N_13227,N_11561,N_11552);
or U13228 (N_13228,N_11742,N_10712);
nand U13229 (N_13229,N_10907,N_11510);
nor U13230 (N_13230,N_10836,N_10853);
and U13231 (N_13231,N_11702,N_11204);
and U13232 (N_13232,N_11035,N_11720);
or U13233 (N_13233,N_11508,N_11989);
or U13234 (N_13234,N_11552,N_10858);
and U13235 (N_13235,N_11099,N_11647);
and U13236 (N_13236,N_10976,N_10695);
or U13237 (N_13237,N_11612,N_10713);
nor U13238 (N_13238,N_10591,N_10926);
and U13239 (N_13239,N_11186,N_11988);
or U13240 (N_13240,N_11518,N_10566);
nor U13241 (N_13241,N_10849,N_11480);
or U13242 (N_13242,N_11341,N_11609);
nor U13243 (N_13243,N_11597,N_11951);
or U13244 (N_13244,N_11302,N_11320);
nand U13245 (N_13245,N_11780,N_10927);
nand U13246 (N_13246,N_11927,N_10951);
nand U13247 (N_13247,N_11582,N_11456);
xnor U13248 (N_13248,N_11161,N_11648);
and U13249 (N_13249,N_11387,N_11187);
nand U13250 (N_13250,N_10786,N_11698);
nand U13251 (N_13251,N_11876,N_10760);
and U13252 (N_13252,N_10636,N_10520);
xor U13253 (N_13253,N_10987,N_10795);
and U13254 (N_13254,N_11178,N_11760);
xor U13255 (N_13255,N_10500,N_11354);
nor U13256 (N_13256,N_11746,N_11024);
nand U13257 (N_13257,N_11766,N_11277);
xor U13258 (N_13258,N_10528,N_11098);
nor U13259 (N_13259,N_11935,N_11891);
and U13260 (N_13260,N_11132,N_11965);
and U13261 (N_13261,N_11847,N_11677);
nand U13262 (N_13262,N_11249,N_11494);
nor U13263 (N_13263,N_11002,N_10929);
and U13264 (N_13264,N_10529,N_11255);
nand U13265 (N_13265,N_11396,N_11238);
nor U13266 (N_13266,N_10635,N_10533);
nor U13267 (N_13267,N_11226,N_11037);
nand U13268 (N_13268,N_11628,N_11834);
and U13269 (N_13269,N_11275,N_11343);
or U13270 (N_13270,N_11859,N_11498);
nor U13271 (N_13271,N_11968,N_11923);
xor U13272 (N_13272,N_10975,N_11531);
nand U13273 (N_13273,N_11794,N_10516);
xnor U13274 (N_13274,N_11550,N_10855);
nand U13275 (N_13275,N_11694,N_11024);
and U13276 (N_13276,N_11316,N_11065);
xor U13277 (N_13277,N_11527,N_10603);
nor U13278 (N_13278,N_11082,N_10759);
or U13279 (N_13279,N_11310,N_11334);
and U13280 (N_13280,N_11312,N_11052);
and U13281 (N_13281,N_10995,N_10826);
xnor U13282 (N_13282,N_11652,N_10657);
or U13283 (N_13283,N_11791,N_11711);
nand U13284 (N_13284,N_10674,N_10941);
nor U13285 (N_13285,N_11166,N_11899);
or U13286 (N_13286,N_11842,N_11427);
nor U13287 (N_13287,N_11565,N_10657);
or U13288 (N_13288,N_10868,N_11540);
nand U13289 (N_13289,N_10924,N_10555);
nand U13290 (N_13290,N_11286,N_11122);
xor U13291 (N_13291,N_11593,N_10737);
and U13292 (N_13292,N_10653,N_11875);
nor U13293 (N_13293,N_11674,N_11980);
and U13294 (N_13294,N_11975,N_11510);
and U13295 (N_13295,N_11661,N_11722);
xor U13296 (N_13296,N_11547,N_11466);
or U13297 (N_13297,N_10987,N_11951);
and U13298 (N_13298,N_11487,N_11512);
or U13299 (N_13299,N_11673,N_10951);
xor U13300 (N_13300,N_11794,N_11294);
nand U13301 (N_13301,N_11482,N_11144);
xor U13302 (N_13302,N_10595,N_10895);
or U13303 (N_13303,N_11426,N_10502);
and U13304 (N_13304,N_10685,N_11323);
xnor U13305 (N_13305,N_11188,N_10715);
xnor U13306 (N_13306,N_11906,N_10801);
xnor U13307 (N_13307,N_11010,N_11978);
and U13308 (N_13308,N_11928,N_10567);
nor U13309 (N_13309,N_11308,N_10968);
and U13310 (N_13310,N_11409,N_10837);
nand U13311 (N_13311,N_11251,N_11557);
or U13312 (N_13312,N_11533,N_10749);
and U13313 (N_13313,N_10773,N_10859);
nand U13314 (N_13314,N_10869,N_11201);
nand U13315 (N_13315,N_11940,N_11974);
and U13316 (N_13316,N_10622,N_10500);
and U13317 (N_13317,N_11272,N_11986);
nand U13318 (N_13318,N_11108,N_10748);
nand U13319 (N_13319,N_11714,N_11950);
or U13320 (N_13320,N_11585,N_11285);
and U13321 (N_13321,N_10784,N_10546);
nand U13322 (N_13322,N_11294,N_11670);
nand U13323 (N_13323,N_11437,N_10634);
and U13324 (N_13324,N_10833,N_11340);
nor U13325 (N_13325,N_11679,N_11068);
or U13326 (N_13326,N_10862,N_11508);
xor U13327 (N_13327,N_10803,N_10645);
xnor U13328 (N_13328,N_11397,N_11697);
and U13329 (N_13329,N_11558,N_11539);
xor U13330 (N_13330,N_10549,N_11701);
xor U13331 (N_13331,N_11645,N_10849);
xnor U13332 (N_13332,N_11580,N_11239);
or U13333 (N_13333,N_10546,N_10839);
nor U13334 (N_13334,N_11251,N_10748);
or U13335 (N_13335,N_11948,N_10652);
nand U13336 (N_13336,N_11909,N_11195);
and U13337 (N_13337,N_11685,N_11508);
nor U13338 (N_13338,N_11356,N_11952);
xor U13339 (N_13339,N_11172,N_11283);
nand U13340 (N_13340,N_11406,N_10800);
or U13341 (N_13341,N_11697,N_11172);
and U13342 (N_13342,N_11109,N_11738);
nand U13343 (N_13343,N_11527,N_11399);
xnor U13344 (N_13344,N_11627,N_11835);
and U13345 (N_13345,N_11266,N_11259);
or U13346 (N_13346,N_10730,N_11592);
nand U13347 (N_13347,N_11724,N_11658);
and U13348 (N_13348,N_11874,N_11016);
nand U13349 (N_13349,N_10839,N_10815);
and U13350 (N_13350,N_11233,N_11019);
nor U13351 (N_13351,N_11828,N_11678);
nand U13352 (N_13352,N_11518,N_11974);
and U13353 (N_13353,N_11303,N_11058);
or U13354 (N_13354,N_10674,N_11864);
nor U13355 (N_13355,N_11881,N_11385);
or U13356 (N_13356,N_11735,N_10662);
nand U13357 (N_13357,N_10679,N_11494);
nor U13358 (N_13358,N_11397,N_10691);
nand U13359 (N_13359,N_10854,N_11389);
or U13360 (N_13360,N_10520,N_10843);
or U13361 (N_13361,N_11062,N_10621);
nor U13362 (N_13362,N_11713,N_11090);
nor U13363 (N_13363,N_10796,N_11501);
or U13364 (N_13364,N_11201,N_11231);
nand U13365 (N_13365,N_11657,N_11426);
nor U13366 (N_13366,N_11127,N_11164);
and U13367 (N_13367,N_10743,N_11226);
nor U13368 (N_13368,N_11928,N_11408);
and U13369 (N_13369,N_10955,N_11359);
nand U13370 (N_13370,N_11455,N_10766);
or U13371 (N_13371,N_11550,N_10606);
nand U13372 (N_13372,N_10931,N_10695);
or U13373 (N_13373,N_11302,N_11984);
nor U13374 (N_13374,N_11038,N_11088);
xor U13375 (N_13375,N_11178,N_10909);
xor U13376 (N_13376,N_11245,N_11359);
or U13377 (N_13377,N_11283,N_11515);
or U13378 (N_13378,N_10593,N_11741);
or U13379 (N_13379,N_11957,N_11987);
and U13380 (N_13380,N_10979,N_11413);
and U13381 (N_13381,N_10587,N_10972);
or U13382 (N_13382,N_11978,N_11677);
nor U13383 (N_13383,N_11347,N_11993);
nand U13384 (N_13384,N_10997,N_10811);
and U13385 (N_13385,N_11970,N_11232);
nor U13386 (N_13386,N_11496,N_11382);
xnor U13387 (N_13387,N_10828,N_11690);
xor U13388 (N_13388,N_11614,N_11982);
nand U13389 (N_13389,N_11591,N_11136);
or U13390 (N_13390,N_11215,N_10567);
and U13391 (N_13391,N_11887,N_11848);
xnor U13392 (N_13392,N_10544,N_10667);
and U13393 (N_13393,N_10691,N_11290);
nor U13394 (N_13394,N_11776,N_11130);
xor U13395 (N_13395,N_11427,N_11992);
and U13396 (N_13396,N_11008,N_11933);
nor U13397 (N_13397,N_10749,N_10719);
and U13398 (N_13398,N_11360,N_11884);
nor U13399 (N_13399,N_10629,N_11426);
or U13400 (N_13400,N_10680,N_10567);
or U13401 (N_13401,N_10732,N_11697);
nor U13402 (N_13402,N_10973,N_11951);
or U13403 (N_13403,N_11721,N_11544);
and U13404 (N_13404,N_11360,N_11120);
xnor U13405 (N_13405,N_10701,N_11834);
nor U13406 (N_13406,N_10576,N_11812);
and U13407 (N_13407,N_11789,N_11339);
or U13408 (N_13408,N_10802,N_11048);
xnor U13409 (N_13409,N_11432,N_10601);
nor U13410 (N_13410,N_10762,N_10900);
nand U13411 (N_13411,N_11586,N_10829);
nand U13412 (N_13412,N_11957,N_10859);
nor U13413 (N_13413,N_10782,N_10566);
nand U13414 (N_13414,N_11285,N_10772);
and U13415 (N_13415,N_10721,N_10971);
and U13416 (N_13416,N_10867,N_10903);
or U13417 (N_13417,N_11641,N_10887);
nor U13418 (N_13418,N_11243,N_11490);
or U13419 (N_13419,N_10742,N_10818);
nand U13420 (N_13420,N_10926,N_10928);
nand U13421 (N_13421,N_11993,N_10522);
xnor U13422 (N_13422,N_11007,N_10934);
nor U13423 (N_13423,N_11018,N_11498);
and U13424 (N_13424,N_11097,N_10595);
nand U13425 (N_13425,N_11470,N_11533);
nor U13426 (N_13426,N_11420,N_11940);
nor U13427 (N_13427,N_10564,N_10766);
xor U13428 (N_13428,N_11036,N_11381);
nand U13429 (N_13429,N_10616,N_11070);
nand U13430 (N_13430,N_10984,N_11621);
and U13431 (N_13431,N_11576,N_11490);
or U13432 (N_13432,N_11840,N_11648);
nand U13433 (N_13433,N_10774,N_11379);
nand U13434 (N_13434,N_11497,N_11144);
xor U13435 (N_13435,N_10850,N_10766);
and U13436 (N_13436,N_10675,N_11987);
xor U13437 (N_13437,N_11552,N_10944);
xor U13438 (N_13438,N_11029,N_11697);
nand U13439 (N_13439,N_11895,N_10922);
nor U13440 (N_13440,N_11338,N_10533);
and U13441 (N_13441,N_10687,N_11911);
nand U13442 (N_13442,N_11960,N_10781);
nand U13443 (N_13443,N_11890,N_10871);
or U13444 (N_13444,N_11506,N_11589);
and U13445 (N_13445,N_10613,N_11615);
or U13446 (N_13446,N_10839,N_11599);
nand U13447 (N_13447,N_10583,N_11772);
nand U13448 (N_13448,N_11048,N_10715);
and U13449 (N_13449,N_10972,N_11669);
or U13450 (N_13450,N_11903,N_11221);
nor U13451 (N_13451,N_10976,N_10513);
nor U13452 (N_13452,N_11109,N_10571);
and U13453 (N_13453,N_11260,N_11762);
and U13454 (N_13454,N_11897,N_10835);
nand U13455 (N_13455,N_10756,N_10937);
nand U13456 (N_13456,N_10616,N_11320);
or U13457 (N_13457,N_11169,N_11901);
nor U13458 (N_13458,N_11777,N_11420);
or U13459 (N_13459,N_10984,N_10750);
or U13460 (N_13460,N_11283,N_10540);
nand U13461 (N_13461,N_10764,N_10982);
and U13462 (N_13462,N_10954,N_11041);
xor U13463 (N_13463,N_11428,N_11381);
or U13464 (N_13464,N_10871,N_11954);
nand U13465 (N_13465,N_11386,N_10609);
nand U13466 (N_13466,N_11848,N_11436);
xnor U13467 (N_13467,N_11968,N_10529);
nor U13468 (N_13468,N_11764,N_11834);
nor U13469 (N_13469,N_10555,N_11418);
or U13470 (N_13470,N_10861,N_10774);
or U13471 (N_13471,N_10549,N_10759);
and U13472 (N_13472,N_11380,N_10749);
nand U13473 (N_13473,N_11500,N_11727);
or U13474 (N_13474,N_10759,N_11094);
or U13475 (N_13475,N_10707,N_11797);
xor U13476 (N_13476,N_11765,N_11616);
nand U13477 (N_13477,N_10658,N_10555);
nor U13478 (N_13478,N_11853,N_10716);
and U13479 (N_13479,N_10828,N_11602);
or U13480 (N_13480,N_11586,N_11905);
nand U13481 (N_13481,N_11413,N_10859);
and U13482 (N_13482,N_11774,N_11924);
xnor U13483 (N_13483,N_11192,N_10661);
xor U13484 (N_13484,N_11972,N_11948);
nand U13485 (N_13485,N_10768,N_11528);
nor U13486 (N_13486,N_10914,N_11602);
nor U13487 (N_13487,N_11080,N_11628);
xor U13488 (N_13488,N_11978,N_10745);
nor U13489 (N_13489,N_10518,N_10644);
or U13490 (N_13490,N_11424,N_11917);
xnor U13491 (N_13491,N_10820,N_10723);
xnor U13492 (N_13492,N_11971,N_11635);
nor U13493 (N_13493,N_11651,N_10777);
and U13494 (N_13494,N_11818,N_11766);
xnor U13495 (N_13495,N_11393,N_11780);
nand U13496 (N_13496,N_11965,N_11055);
nand U13497 (N_13497,N_10874,N_10669);
and U13498 (N_13498,N_11066,N_10905);
nand U13499 (N_13499,N_11939,N_10690);
nor U13500 (N_13500,N_12558,N_12000);
xnor U13501 (N_13501,N_13095,N_12909);
and U13502 (N_13502,N_13165,N_13104);
nor U13503 (N_13503,N_12842,N_13158);
nor U13504 (N_13504,N_12657,N_13319);
nor U13505 (N_13505,N_12918,N_12216);
nand U13506 (N_13506,N_12617,N_12434);
nor U13507 (N_13507,N_13237,N_12259);
nor U13508 (N_13508,N_12070,N_12645);
xor U13509 (N_13509,N_12827,N_13309);
nand U13510 (N_13510,N_13068,N_13234);
and U13511 (N_13511,N_12838,N_13103);
xor U13512 (N_13512,N_12149,N_13343);
nand U13513 (N_13513,N_12920,N_12686);
nand U13514 (N_13514,N_13163,N_12462);
and U13515 (N_13515,N_12321,N_12507);
nor U13516 (N_13516,N_13026,N_12288);
nor U13517 (N_13517,N_13116,N_12375);
and U13518 (N_13518,N_12812,N_12243);
nand U13519 (N_13519,N_12448,N_12287);
and U13520 (N_13520,N_13069,N_13266);
xnor U13521 (N_13521,N_12622,N_12214);
or U13522 (N_13522,N_13423,N_12575);
or U13523 (N_13523,N_12994,N_12658);
nand U13524 (N_13524,N_13204,N_13169);
or U13525 (N_13525,N_12353,N_13098);
nand U13526 (N_13526,N_12295,N_12407);
or U13527 (N_13527,N_13414,N_12406);
and U13528 (N_13528,N_12568,N_12146);
or U13529 (N_13529,N_12841,N_12416);
nor U13530 (N_13530,N_12897,N_12690);
and U13531 (N_13531,N_12650,N_13498);
nor U13532 (N_13532,N_12627,N_12505);
nor U13533 (N_13533,N_13185,N_13445);
or U13534 (N_13534,N_13194,N_12183);
nand U13535 (N_13535,N_13294,N_12802);
and U13536 (N_13536,N_13032,N_12563);
or U13537 (N_13537,N_13226,N_12527);
and U13538 (N_13538,N_12394,N_12364);
xnor U13539 (N_13539,N_12385,N_12002);
nor U13540 (N_13540,N_12153,N_12386);
nor U13541 (N_13541,N_12176,N_12671);
and U13542 (N_13542,N_12667,N_12262);
or U13543 (N_13543,N_12552,N_12097);
xor U13544 (N_13544,N_13182,N_12514);
and U13545 (N_13545,N_13313,N_13058);
nand U13546 (N_13546,N_12982,N_12450);
nand U13547 (N_13547,N_12119,N_12706);
xor U13548 (N_13548,N_13089,N_13245);
xnor U13549 (N_13549,N_13388,N_13004);
xnor U13550 (N_13550,N_13008,N_12720);
or U13551 (N_13551,N_12319,N_12378);
nand U13552 (N_13552,N_12754,N_12465);
nor U13553 (N_13553,N_13341,N_12009);
nand U13554 (N_13554,N_12508,N_12863);
or U13555 (N_13555,N_12976,N_13457);
xnor U13556 (N_13556,N_12785,N_13320);
or U13557 (N_13557,N_13386,N_12776);
and U13558 (N_13558,N_12299,N_12362);
xor U13559 (N_13559,N_12055,N_13330);
or U13560 (N_13560,N_12726,N_12087);
nand U13561 (N_13561,N_12439,N_12652);
nand U13562 (N_13562,N_12056,N_13249);
nor U13563 (N_13563,N_13499,N_12155);
or U13564 (N_13564,N_13323,N_12290);
and U13565 (N_13565,N_12495,N_13461);
xnor U13566 (N_13566,N_12526,N_13228);
nor U13567 (N_13567,N_13391,N_12502);
and U13568 (N_13568,N_12503,N_12731);
xnor U13569 (N_13569,N_12561,N_12583);
xor U13570 (N_13570,N_12150,N_13208);
nand U13571 (N_13571,N_12529,N_12955);
and U13572 (N_13572,N_13418,N_12922);
nand U13573 (N_13573,N_12094,N_13495);
and U13574 (N_13574,N_13028,N_12784);
or U13575 (N_13575,N_13367,N_12033);
or U13576 (N_13576,N_12964,N_13238);
xor U13577 (N_13577,N_12993,N_12557);
nand U13578 (N_13578,N_13299,N_13361);
or U13579 (N_13579,N_12478,N_12732);
xnor U13580 (N_13580,N_12068,N_13113);
xor U13581 (N_13581,N_12931,N_12887);
nand U13582 (N_13582,N_13213,N_13020);
xor U13583 (N_13583,N_12408,N_12674);
xnor U13584 (N_13584,N_13394,N_13417);
and U13585 (N_13585,N_12206,N_12882);
nor U13586 (N_13586,N_12591,N_12152);
nand U13587 (N_13587,N_12130,N_12515);
or U13588 (N_13588,N_13354,N_13203);
nor U13589 (N_13589,N_12967,N_12270);
nor U13590 (N_13590,N_12142,N_13421);
nor U13591 (N_13591,N_12469,N_12555);
or U13592 (N_13592,N_13351,N_12835);
nor U13593 (N_13593,N_13419,N_12898);
nor U13594 (N_13594,N_12626,N_12940);
and U13595 (N_13595,N_12231,N_12168);
nor U13596 (N_13596,N_13278,N_12379);
xor U13597 (N_13597,N_13007,N_12062);
nor U13598 (N_13598,N_12553,N_12770);
nand U13599 (N_13599,N_12410,N_12984);
or U13600 (N_13600,N_12343,N_12774);
or U13601 (N_13601,N_12883,N_13493);
nor U13602 (N_13602,N_12285,N_12170);
and U13603 (N_13603,N_12913,N_12317);
nor U13604 (N_13604,N_12892,N_12830);
nor U13605 (N_13605,N_12683,N_13215);
nand U13606 (N_13606,N_12934,N_12661);
xor U13607 (N_13607,N_12843,N_13356);
nand U13608 (N_13608,N_13040,N_12173);
xnor U13609 (N_13609,N_12884,N_13131);
nor U13610 (N_13610,N_13373,N_12860);
nor U13611 (N_13611,N_12966,N_12672);
or U13612 (N_13612,N_13154,N_12769);
xnor U13613 (N_13613,N_12534,N_12020);
and U13614 (N_13614,N_12151,N_13168);
and U13615 (N_13615,N_12161,N_13362);
nand U13616 (N_13616,N_12393,N_13171);
nor U13617 (N_13617,N_12189,N_13325);
xor U13618 (N_13618,N_12349,N_12877);
nor U13619 (N_13619,N_13065,N_12158);
or U13620 (N_13620,N_12419,N_12264);
nand U13621 (N_13621,N_12134,N_12044);
nand U13622 (N_13622,N_13398,N_13297);
nand U13623 (N_13623,N_12813,N_13030);
or U13624 (N_13624,N_12197,N_13409);
nand U13625 (N_13625,N_13257,N_12422);
or U13626 (N_13626,N_12054,N_12912);
nand U13627 (N_13627,N_12900,N_13440);
or U13628 (N_13628,N_12577,N_12085);
xnor U13629 (N_13629,N_12245,N_12005);
and U13630 (N_13630,N_12643,N_12950);
or U13631 (N_13631,N_12533,N_12590);
and U13632 (N_13632,N_13273,N_12923);
nor U13633 (N_13633,N_12480,N_13491);
and U13634 (N_13634,N_12392,N_12129);
and U13635 (N_13635,N_13144,N_12704);
xnor U13636 (N_13636,N_13400,N_12397);
and U13637 (N_13637,N_13081,N_13043);
and U13638 (N_13638,N_12653,N_12954);
and U13639 (N_13639,N_12609,N_12429);
nand U13640 (N_13640,N_12840,N_12099);
nand U13641 (N_13641,N_12449,N_13346);
xor U13642 (N_13642,N_12511,N_12562);
nand U13643 (N_13643,N_13025,N_12972);
nand U13644 (N_13644,N_12127,N_12023);
or U13645 (N_13645,N_13370,N_12866);
and U13646 (N_13646,N_13124,N_12438);
nand U13647 (N_13647,N_12095,N_12177);
and U13648 (N_13648,N_12342,N_12942);
and U13649 (N_13649,N_12071,N_12953);
and U13650 (N_13650,N_12907,N_12952);
nor U13651 (N_13651,N_12461,N_13413);
and U13652 (N_13652,N_12513,N_12028);
nor U13653 (N_13653,N_12398,N_12600);
xor U13654 (N_13654,N_13360,N_13059);
nand U13655 (N_13655,N_12905,N_12010);
nand U13656 (N_13656,N_12693,N_12293);
and U13657 (N_13657,N_12999,N_12181);
nor U13658 (N_13658,N_12535,N_12615);
xnor U13659 (N_13659,N_13022,N_13101);
nor U13660 (N_13660,N_13250,N_12037);
nand U13661 (N_13661,N_12484,N_12607);
or U13662 (N_13662,N_12681,N_13047);
or U13663 (N_13663,N_13239,N_13242);
xnor U13664 (N_13664,N_12579,N_13286);
nand U13665 (N_13665,N_12601,N_13014);
nand U13666 (N_13666,N_12987,N_12226);
nor U13667 (N_13667,N_12791,N_13251);
or U13668 (N_13668,N_12702,N_12137);
nor U13669 (N_13669,N_12413,N_12516);
xnor U13670 (N_13670,N_12793,N_12329);
xor U13671 (N_13671,N_12623,N_12807);
nand U13672 (N_13672,N_12052,N_12576);
nand U13673 (N_13673,N_12756,N_12805);
or U13674 (N_13674,N_12598,N_13492);
and U13675 (N_13675,N_12676,N_13038);
nand U13676 (N_13676,N_12989,N_12796);
xor U13677 (N_13677,N_13195,N_12747);
and U13678 (N_13678,N_12811,N_13324);
xnor U13679 (N_13679,N_13255,N_12716);
or U13680 (N_13680,N_13055,N_12477);
xor U13681 (N_13681,N_12744,N_12082);
or U13682 (N_13682,N_12107,N_12935);
or U13683 (N_13683,N_12207,N_12852);
nor U13684 (N_13684,N_13090,N_13267);
xor U13685 (N_13685,N_12192,N_12175);
nand U13686 (N_13686,N_12403,N_13114);
nor U13687 (N_13687,N_13329,N_12944);
xor U13688 (N_13688,N_12361,N_12330);
and U13689 (N_13689,N_12347,N_12629);
and U13690 (N_13690,N_12902,N_13379);
or U13691 (N_13691,N_13444,N_12211);
nand U13692 (N_13692,N_12673,N_12316);
nor U13693 (N_13693,N_12179,N_12586);
nor U13694 (N_13694,N_12749,N_12808);
nand U13695 (N_13695,N_12306,N_12460);
nor U13696 (N_13696,N_12133,N_12560);
nand U13697 (N_13697,N_13146,N_13312);
and U13698 (N_13698,N_12339,N_13214);
and U13699 (N_13699,N_13316,N_13156);
nand U13700 (N_13700,N_13034,N_12696);
and U13701 (N_13701,N_12008,N_12937);
and U13702 (N_13702,N_12510,N_13223);
xor U13703 (N_13703,N_12414,N_12700);
xor U13704 (N_13704,N_12881,N_12402);
xnor U13705 (N_13705,N_13383,N_13137);
or U13706 (N_13706,N_13295,N_12272);
nand U13707 (N_13707,N_13322,N_12546);
nand U13708 (N_13708,N_12286,N_12483);
xor U13709 (N_13709,N_12276,N_12388);
nor U13710 (N_13710,N_12228,N_12616);
or U13711 (N_13711,N_13128,N_12297);
xnor U13712 (N_13712,N_13450,N_12034);
nor U13713 (N_13713,N_12543,N_13363);
and U13714 (N_13714,N_12668,N_13305);
xor U13715 (N_13715,N_12701,N_12694);
nor U13716 (N_13716,N_12752,N_12518);
nor U13717 (N_13717,N_13254,N_12090);
or U13718 (N_13718,N_12167,N_12389);
nor U13719 (N_13719,N_13233,N_12337);
and U13720 (N_13720,N_13331,N_13206);
nor U13721 (N_13721,N_12431,N_13080);
and U13722 (N_13722,N_13201,N_13100);
or U13723 (N_13723,N_12823,N_12986);
nor U13724 (N_13724,N_13121,N_13129);
nor U13725 (N_13725,N_12938,N_12336);
or U13726 (N_13726,N_12219,N_12525);
nor U13727 (N_13727,N_13046,N_12267);
and U13728 (N_13728,N_13123,N_12049);
nand U13729 (N_13729,N_12740,N_12006);
and U13730 (N_13730,N_12022,N_13264);
and U13731 (N_13731,N_12331,N_12418);
xor U13732 (N_13732,N_13284,N_13212);
or U13733 (N_13733,N_12684,N_12069);
and U13734 (N_13734,N_13280,N_13377);
nand U13735 (N_13735,N_12233,N_13172);
nand U13736 (N_13736,N_12890,N_12303);
xnor U13737 (N_13737,N_12939,N_12366);
nor U13738 (N_13738,N_12359,N_12113);
xor U13739 (N_13739,N_12217,N_12766);
and U13740 (N_13740,N_13357,N_13350);
or U13741 (N_13741,N_12715,N_13380);
and U13742 (N_13742,N_13127,N_12584);
and U13743 (N_13743,N_12888,N_13184);
or U13744 (N_13744,N_12171,N_12415);
or U13745 (N_13745,N_12757,N_12642);
or U13746 (N_13746,N_12880,N_13265);
nand U13747 (N_13747,N_13192,N_12496);
xor U13748 (N_13748,N_12798,N_13452);
and U13749 (N_13749,N_12417,N_13023);
and U13750 (N_13750,N_13407,N_12481);
nor U13751 (N_13751,N_12244,N_12831);
and U13752 (N_13752,N_12550,N_12445);
xnor U13753 (N_13753,N_12611,N_12395);
or U13754 (N_13754,N_13359,N_12196);
and U13755 (N_13755,N_12220,N_13064);
nor U13756 (N_13756,N_12335,N_12426);
nand U13757 (N_13757,N_12662,N_12369);
nand U13758 (N_13758,N_12868,N_13092);
xor U13759 (N_13759,N_12501,N_13235);
xor U13760 (N_13760,N_12194,N_12135);
nor U13761 (N_13761,N_13241,N_13480);
nor U13762 (N_13762,N_13497,N_12848);
xnor U13763 (N_13763,N_12936,N_12352);
and U13764 (N_13764,N_12614,N_12261);
nand U13765 (N_13765,N_13135,N_12030);
xor U13766 (N_13766,N_13109,N_12363);
or U13767 (N_13767,N_12540,N_12790);
xnor U13768 (N_13768,N_13490,N_12806);
nor U13769 (N_13769,N_13411,N_13436);
xor U13770 (N_13770,N_13397,N_12430);
nand U13771 (N_13771,N_12844,N_12734);
or U13772 (N_13772,N_13134,N_13406);
and U13773 (N_13773,N_12644,N_12539);
xor U13774 (N_13774,N_12433,N_13384);
or U13775 (N_13775,N_12160,N_13476);
or U13776 (N_13776,N_12574,N_12132);
and U13777 (N_13777,N_13196,N_12745);
nand U13778 (N_13778,N_13066,N_12436);
or U13779 (N_13779,N_12582,N_13037);
and U13780 (N_13780,N_13220,N_12677);
or U13781 (N_13781,N_13140,N_12588);
xor U13782 (N_13782,N_12633,N_12489);
or U13783 (N_13783,N_12190,N_13456);
nand U13784 (N_13784,N_13447,N_12159);
nand U13785 (N_13785,N_13017,N_12530);
xor U13786 (N_13786,N_12669,N_12029);
xor U13787 (N_13787,N_12273,N_13118);
xnor U13788 (N_13788,N_12929,N_13344);
or U13789 (N_13789,N_12320,N_13211);
or U13790 (N_13790,N_13410,N_12919);
and U13791 (N_13791,N_13395,N_12066);
and U13792 (N_13792,N_13460,N_12504);
and U13793 (N_13793,N_13258,N_12845);
nand U13794 (N_13794,N_12487,N_12688);
and U13795 (N_13795,N_12472,N_13151);
and U13796 (N_13796,N_12140,N_13096);
and U13797 (N_13797,N_13326,N_13160);
xor U13798 (N_13798,N_12382,N_12664);
or U13799 (N_13799,N_12663,N_12506);
nand U13800 (N_13800,N_12456,N_13375);
xnor U13801 (N_13801,N_12255,N_13292);
nand U13802 (N_13802,N_13405,N_12400);
xor U13803 (N_13803,N_12679,N_13145);
nor U13804 (N_13804,N_12828,N_12188);
nand U13805 (N_13805,N_12618,N_12545);
or U13806 (N_13806,N_13321,N_13272);
xnor U13807 (N_13807,N_12794,N_13256);
and U13808 (N_13808,N_12230,N_13368);
nor U13809 (N_13809,N_12046,N_12334);
or U13810 (N_13810,N_13166,N_12763);
nand U13811 (N_13811,N_13448,N_13246);
nand U13812 (N_13812,N_12846,N_12311);
nor U13813 (N_13813,N_13304,N_12454);
or U13814 (N_13814,N_12943,N_12820);
xor U13815 (N_13815,N_12145,N_13438);
nor U13816 (N_13816,N_12968,N_13314);
xor U13817 (N_13817,N_12819,N_12391);
and U13818 (N_13818,N_12258,N_13051);
xnor U13819 (N_13819,N_12691,N_13473);
and U13820 (N_13820,N_13381,N_13177);
xor U13821 (N_13821,N_12640,N_12241);
xnor U13822 (N_13822,N_12559,N_12750);
xnor U13823 (N_13823,N_12101,N_12076);
and U13824 (N_13824,N_13427,N_13084);
nor U13825 (N_13825,N_13161,N_13050);
xor U13826 (N_13826,N_12200,N_13013);
nor U13827 (N_13827,N_13041,N_12915);
xor U13828 (N_13828,N_13307,N_12777);
nand U13829 (N_13829,N_12473,N_13333);
nand U13830 (N_13830,N_13259,N_13031);
xnor U13831 (N_13831,N_12300,N_13496);
xnor U13832 (N_13832,N_12310,N_12411);
nand U13833 (N_13833,N_13225,N_13477);
and U13834 (N_13834,N_13083,N_13401);
or U13835 (N_13835,N_12593,N_12628);
or U13836 (N_13836,N_13252,N_12594);
nand U13837 (N_13837,N_13396,N_13253);
nand U13838 (N_13838,N_12497,N_12779);
xnor U13839 (N_13839,N_12064,N_12722);
nand U13840 (N_13840,N_12136,N_12974);
nand U13841 (N_13841,N_12592,N_12581);
nor U13842 (N_13842,N_12238,N_12441);
nor U13843 (N_13843,N_13337,N_12743);
or U13844 (N_13844,N_12224,N_12098);
nand U13845 (N_13845,N_12072,N_13062);
xor U13846 (N_13846,N_12862,N_12043);
and U13847 (N_13847,N_12970,N_12960);
xnor U13848 (N_13848,N_13119,N_13334);
nand U13849 (N_13849,N_13230,N_13178);
xor U13850 (N_13850,N_13479,N_12815);
xnor U13851 (N_13851,N_12865,N_13443);
or U13852 (N_13852,N_12075,N_12492);
or U13853 (N_13853,N_13282,N_12079);
xor U13854 (N_13854,N_13317,N_13045);
or U13855 (N_13855,N_12788,N_13029);
or U13856 (N_13856,N_12965,N_12390);
or U13857 (N_13857,N_12093,N_12724);
xnor U13858 (N_13858,N_13277,N_12309);
nand U13859 (N_13859,N_12237,N_12755);
and U13860 (N_13860,N_13247,N_13489);
or U13861 (N_13861,N_12759,N_12131);
nand U13862 (N_13862,N_12872,N_12123);
or U13863 (N_13863,N_13345,N_12458);
or U13864 (N_13864,N_12067,N_12738);
nor U13865 (N_13865,N_13173,N_12187);
and U13866 (N_13866,N_12482,N_12787);
nand U13867 (N_13867,N_13152,N_12512);
nor U13868 (N_13868,N_12120,N_12758);
or U13869 (N_13869,N_13308,N_12396);
and U13870 (N_13870,N_12283,N_13229);
nand U13871 (N_13871,N_12893,N_13422);
nor U13872 (N_13872,N_13276,N_13102);
nand U13873 (N_13873,N_13200,N_12762);
nand U13874 (N_13874,N_13449,N_12257);
nand U13875 (N_13875,N_13073,N_13126);
nor U13876 (N_13876,N_13120,N_12692);
nor U13877 (N_13877,N_12695,N_12963);
nor U13878 (N_13878,N_13216,N_13382);
nor U13879 (N_13879,N_13475,N_12017);
and U13880 (N_13880,N_12589,N_13481);
and U13881 (N_13881,N_13222,N_12685);
and U13882 (N_13882,N_12003,N_13306);
and U13883 (N_13883,N_12926,N_13376);
xnor U13884 (N_13884,N_13087,N_12365);
or U13885 (N_13885,N_12274,N_12971);
or U13886 (N_13886,N_12795,N_12631);
and U13887 (N_13887,N_12878,N_12603);
xor U13888 (N_13888,N_13130,N_13459);
nor U13889 (N_13889,N_13079,N_13385);
xor U13890 (N_13890,N_12263,N_12873);
nor U13891 (N_13891,N_12199,N_12718);
nand U13892 (N_13892,N_12144,N_12240);
and U13893 (N_13893,N_12027,N_13056);
xor U13894 (N_13894,N_12169,N_13060);
and U13895 (N_13895,N_12304,N_12485);
nand U13896 (N_13896,N_13108,N_12229);
xnor U13897 (N_13897,N_12871,N_13143);
xor U13898 (N_13898,N_13402,N_13052);
nor U13899 (N_13899,N_12567,N_12855);
and U13900 (N_13900,N_12102,N_12980);
and U13901 (N_13901,N_12235,N_12057);
nand U13902 (N_13902,N_12797,N_12073);
nand U13903 (N_13903,N_13300,N_12383);
nand U13904 (N_13904,N_13487,N_12201);
nor U13905 (N_13905,N_13378,N_13164);
xor U13906 (N_13906,N_12947,N_13416);
and U13907 (N_13907,N_12111,N_13063);
and U13908 (N_13908,N_13455,N_12799);
or U13909 (N_13909,N_13112,N_13133);
nor U13910 (N_13910,N_13310,N_12531);
or U13911 (N_13911,N_12500,N_13468);
nand U13912 (N_13912,N_12876,N_12440);
xor U13913 (N_13913,N_12091,N_12610);
nand U13914 (N_13914,N_13012,N_12457);
and U13915 (N_13915,N_12193,N_13111);
nand U13916 (N_13916,N_12894,N_12867);
nor U13917 (N_13917,N_12409,N_12624);
nor U13918 (N_13918,N_13082,N_12714);
and U13919 (N_13919,N_13393,N_12746);
xor U13920 (N_13920,N_13198,N_12182);
and U13921 (N_13921,N_12348,N_12325);
and U13922 (N_13922,N_12370,N_13125);
and U13923 (N_13923,N_13467,N_12308);
xnor U13924 (N_13924,N_13430,N_12051);
xor U13925 (N_13925,N_12015,N_12910);
nor U13926 (N_13926,N_12771,N_13117);
and U13927 (N_13927,N_12801,N_12859);
and U13928 (N_13928,N_13353,N_12381);
nand U13929 (N_13929,N_13471,N_13039);
nor U13930 (N_13930,N_12452,N_13077);
and U13931 (N_13931,N_12063,N_13268);
xnor U13932 (N_13932,N_12247,N_13426);
and U13933 (N_13933,N_12857,N_12004);
xor U13934 (N_13934,N_12026,N_12421);
or U13935 (N_13935,N_12768,N_13465);
nor U13936 (N_13936,N_12985,N_12314);
nand U13937 (N_13937,N_12148,N_12162);
and U13938 (N_13938,N_12765,N_13466);
xnor U13939 (N_13939,N_13287,N_12053);
nor U13940 (N_13940,N_12707,N_12675);
xor U13941 (N_13941,N_12346,N_12602);
and U13942 (N_13942,N_12916,N_12467);
and U13943 (N_13943,N_12854,N_13006);
nand U13944 (N_13944,N_13110,N_13094);
nor U13945 (N_13945,N_12651,N_13053);
nand U13946 (N_13946,N_12753,N_13170);
xor U13947 (N_13947,N_12112,N_12014);
or U13948 (N_13948,N_12498,N_12198);
nand U13949 (N_13949,N_12108,N_12138);
or U13950 (N_13950,N_12870,N_12992);
and U13951 (N_13951,N_12141,N_12405);
nor U13952 (N_13952,N_12665,N_12242);
nand U13953 (N_13953,N_12520,N_12350);
or U13954 (N_13954,N_12646,N_12814);
nand U13955 (N_13955,N_12470,N_13269);
or U13956 (N_13956,N_13352,N_13148);
or U13957 (N_13957,N_12373,N_12251);
nor U13958 (N_13958,N_13371,N_12280);
xnor U13959 (N_13959,N_12326,N_13054);
or U13960 (N_13960,N_13451,N_12837);
xor U13961 (N_13961,N_12463,N_13186);
and U13962 (N_13962,N_12659,N_12632);
xor U13963 (N_13963,N_12647,N_12727);
xnor U13964 (N_13964,N_12537,N_13389);
xor U13965 (N_13965,N_12327,N_12065);
nand U13966 (N_13966,N_12147,N_12995);
nand U13967 (N_13967,N_13336,N_12951);
or U13968 (N_13968,N_12089,N_12708);
or U13969 (N_13969,N_13224,N_13298);
nor U13970 (N_13970,N_13019,N_12570);
nand U13971 (N_13971,N_13048,N_12983);
or U13972 (N_13972,N_13187,N_12118);
xor U13973 (N_13973,N_12446,N_12621);
nor U13974 (N_13974,N_12712,N_12804);
xnor U13975 (N_13975,N_12875,N_13458);
or U13976 (N_13976,N_13155,N_13236);
and U13977 (N_13977,N_12269,N_12522);
or U13978 (N_13978,N_12115,N_13424);
nand U13979 (N_13979,N_12164,N_12914);
xnor U13980 (N_13980,N_12444,N_13188);
or U13981 (N_13981,N_12524,N_13009);
and U13982 (N_13982,N_12977,N_12959);
or U13983 (N_13983,N_12532,N_12698);
and U13984 (N_13984,N_13097,N_13387);
xor U13985 (N_13985,N_12656,N_12019);
nor U13986 (N_13986,N_12957,N_12377);
nand U13987 (N_13987,N_12117,N_12428);
nand U13988 (N_13988,N_12184,N_13181);
and U13989 (N_13989,N_12474,N_13016);
nor U13990 (N_13990,N_12494,N_12048);
and U13991 (N_13991,N_12333,N_12466);
nand U13992 (N_13992,N_13086,N_13311);
nor U13993 (N_13993,N_12901,N_13365);
nand U13994 (N_13994,N_13035,N_12917);
nor U13995 (N_13995,N_12641,N_12001);
xnor U13996 (N_13996,N_12163,N_12945);
xnor U13997 (N_13997,N_12031,N_12988);
nor U13998 (N_13998,N_12687,N_12682);
xnor U13999 (N_13999,N_12488,N_12059);
nand U14000 (N_14000,N_12816,N_12869);
nand U14001 (N_14001,N_13167,N_13036);
or U14002 (N_14002,N_13366,N_12899);
or U14003 (N_14003,N_12822,N_12523);
or U14004 (N_14004,N_13275,N_13088);
or U14005 (N_14005,N_12847,N_12585);
xnor U14006 (N_14006,N_12105,N_12821);
or U14007 (N_14007,N_13005,N_12476);
nor U14008 (N_14008,N_12921,N_12432);
nor U14009 (N_14009,N_13243,N_13289);
or U14010 (N_14010,N_12850,N_12648);
nand U14011 (N_14011,N_12620,N_13302);
or U14012 (N_14012,N_12542,N_13027);
or U14013 (N_14013,N_12376,N_12368);
and U14014 (N_14014,N_12271,N_12824);
or U14015 (N_14015,N_12032,N_12891);
nand U14016 (N_14016,N_12709,N_13420);
nand U14017 (N_14017,N_13244,N_12074);
nor U14018 (N_14018,N_12660,N_13328);
nand U14019 (N_14019,N_13075,N_12116);
and U14020 (N_14020,N_12367,N_13176);
nor U14021 (N_14021,N_12345,N_12166);
or U14022 (N_14022,N_12246,N_12289);
or U14023 (N_14023,N_12566,N_12281);
nor U14024 (N_14024,N_13369,N_12941);
or U14025 (N_14025,N_12730,N_12284);
and U14026 (N_14026,N_13431,N_12517);
nor U14027 (N_14027,N_12975,N_12826);
nand U14028 (N_14028,N_12092,N_12719);
or U14029 (N_14029,N_12035,N_12580);
nand U14030 (N_14030,N_12997,N_12895);
xnor U14031 (N_14031,N_13227,N_13454);
nor U14032 (N_14032,N_13159,N_13342);
or U14033 (N_14033,N_12572,N_12932);
nor U14034 (N_14034,N_13141,N_12680);
or U14035 (N_14035,N_12371,N_13115);
and U14036 (N_14036,N_13147,N_12471);
nor U14037 (N_14037,N_12962,N_12829);
and U14038 (N_14038,N_13446,N_12736);
or U14039 (N_14039,N_12475,N_12832);
nand U14040 (N_14040,N_12998,N_13153);
nor U14041 (N_14041,N_12016,N_12556);
and U14042 (N_14042,N_12423,N_12751);
and U14043 (N_14043,N_12697,N_13355);
nor U14044 (N_14044,N_12227,N_13434);
xnor U14045 (N_14045,N_13070,N_13301);
nor U14046 (N_14046,N_12851,N_13248);
and U14047 (N_14047,N_12298,N_12260);
nor U14048 (N_14048,N_12927,N_12282);
nand U14049 (N_14049,N_12425,N_12312);
or U14050 (N_14050,N_12420,N_13033);
nand U14051 (N_14051,N_12165,N_13240);
and U14052 (N_14052,N_12125,N_12569);
nor U14053 (N_14053,N_12924,N_12178);
or U14054 (N_14054,N_12538,N_13000);
nand U14055 (N_14055,N_13180,N_13260);
or U14056 (N_14056,N_12705,N_13085);
and U14057 (N_14057,N_12268,N_12903);
nor U14058 (N_14058,N_12380,N_13441);
xor U14059 (N_14059,N_12979,N_13003);
and U14060 (N_14060,N_13486,N_12025);
nor U14061 (N_14061,N_13270,N_13429);
xor U14062 (N_14062,N_13474,N_12521);
and U14063 (N_14063,N_12549,N_13193);
xor U14064 (N_14064,N_12265,N_12157);
or U14065 (N_14065,N_13432,N_12077);
xor U14066 (N_14066,N_12279,N_12741);
nand U14067 (N_14067,N_12639,N_12908);
xnor U14068 (N_14068,N_12236,N_12996);
xnor U14069 (N_14069,N_13207,N_13018);
xnor U14070 (N_14070,N_12124,N_12354);
nand U14071 (N_14071,N_13439,N_12928);
nand U14072 (N_14072,N_13106,N_13078);
xnor U14073 (N_14073,N_12399,N_13099);
nand U14074 (N_14074,N_12024,N_12948);
and U14075 (N_14075,N_12404,N_12222);
nand U14076 (N_14076,N_13024,N_12764);
or U14077 (N_14077,N_12861,N_13011);
and U14078 (N_14078,N_12748,N_12041);
or U14079 (N_14079,N_12783,N_13315);
or U14080 (N_14080,N_13364,N_12038);
and U14081 (N_14081,N_12649,N_12789);
nand U14082 (N_14082,N_13162,N_13274);
xor U14083 (N_14083,N_12981,N_12013);
and U14084 (N_14084,N_12143,N_12635);
nor U14085 (N_14085,N_13189,N_13074);
xnor U14086 (N_14086,N_12990,N_13091);
xnor U14087 (N_14087,N_12464,N_13093);
nand U14088 (N_14088,N_12729,N_13290);
xnor U14089 (N_14089,N_12301,N_12060);
xnor U14090 (N_14090,N_13049,N_12864);
nand U14091 (N_14091,N_12185,N_13463);
and U14092 (N_14092,N_12904,N_12775);
nor U14093 (N_14093,N_12833,N_12086);
nand U14094 (N_14094,N_13122,N_12551);
or U14095 (N_14095,N_12356,N_12541);
and U14096 (N_14096,N_12536,N_12737);
nor U14097 (N_14097,N_12604,N_13202);
and U14098 (N_14098,N_12424,N_13469);
nor U14099 (N_14099,N_13428,N_12340);
and U14100 (N_14100,N_13175,N_13340);
nand U14101 (N_14101,N_12573,N_12933);
nand U14102 (N_14102,N_12739,N_12874);
or U14103 (N_14103,N_12374,N_12323);
or U14104 (N_14104,N_12703,N_13335);
nand U14105 (N_14105,N_13232,N_12978);
and U14106 (N_14106,N_13218,N_12858);
and U14107 (N_14107,N_12204,N_12443);
or U14108 (N_14108,N_12126,N_13339);
or U14109 (N_14109,N_12786,N_12275);
xnor U14110 (N_14110,N_12218,N_12186);
xor U14111 (N_14111,N_12961,N_12772);
nor U14112 (N_14112,N_12202,N_12442);
xor U14113 (N_14113,N_12225,N_12435);
and U14114 (N_14114,N_13288,N_12886);
nand U14115 (N_14115,N_12215,N_12427);
and U14116 (N_14116,N_12780,N_12612);
or U14117 (N_14117,N_13001,N_13425);
nand U14118 (N_14118,N_12121,N_12313);
xnor U14119 (N_14119,N_13494,N_12879);
and U14120 (N_14120,N_13072,N_13217);
and U14121 (N_14121,N_13482,N_12174);
xnor U14122 (N_14122,N_12114,N_12195);
nor U14123 (N_14123,N_12294,N_12012);
nor U14124 (N_14124,N_12717,N_12358);
nor U14125 (N_14125,N_12578,N_13199);
nand U14126 (N_14126,N_12047,N_12341);
or U14127 (N_14127,N_13279,N_12172);
nor U14128 (N_14128,N_12606,N_12554);
nand U14129 (N_14129,N_12725,N_12723);
xor U14130 (N_14130,N_12767,N_12106);
nor U14131 (N_14131,N_12110,N_12088);
nor U14132 (N_14132,N_13390,N_12372);
and U14133 (N_14133,N_13399,N_12773);
xor U14134 (N_14134,N_12084,N_12670);
or U14135 (N_14135,N_12332,N_12699);
nand U14136 (N_14136,N_13138,N_13453);
nand U14137 (N_14137,N_12666,N_12232);
xor U14138 (N_14138,N_12599,N_12351);
nor U14139 (N_14139,N_12213,N_12083);
or U14140 (N_14140,N_12810,N_13002);
xnor U14141 (N_14141,N_12782,N_12039);
nor U14142 (N_14142,N_12096,N_12991);
and U14143 (N_14143,N_13470,N_12278);
and U14144 (N_14144,N_12493,N_12315);
nor U14145 (N_14145,N_12252,N_12637);
and U14146 (N_14146,N_12803,N_12253);
nor U14147 (N_14147,N_12058,N_13107);
nor U14148 (N_14148,N_12911,N_12519);
and U14149 (N_14149,N_12239,N_12205);
and U14150 (N_14150,N_13190,N_12011);
xnor U14151 (N_14151,N_12248,N_13472);
xor U14152 (N_14152,N_12344,N_12018);
nor U14153 (N_14153,N_13136,N_12209);
nor U14154 (N_14154,N_13157,N_12412);
and U14155 (N_14155,N_12080,N_12447);
nor U14156 (N_14156,N_12036,N_12254);
xnor U14157 (N_14157,N_12930,N_12817);
nor U14158 (N_14158,N_12437,N_12654);
nor U14159 (N_14159,N_12548,N_13408);
or U14160 (N_14160,N_13057,N_13076);
or U14161 (N_14161,N_13210,N_13437);
or U14162 (N_14162,N_13293,N_13303);
nand U14163 (N_14163,N_12689,N_13231);
nand U14164 (N_14164,N_12250,N_12479);
nor U14165 (N_14165,N_13374,N_13464);
nand U14166 (N_14166,N_13435,N_13139);
nand U14167 (N_14167,N_12081,N_12613);
nor U14168 (N_14168,N_13462,N_12778);
or U14169 (N_14169,N_12809,N_13415);
nand U14170 (N_14170,N_13179,N_12360);
and U14171 (N_14171,N_13010,N_13263);
nor U14172 (N_14172,N_12834,N_12728);
and U14173 (N_14173,N_13338,N_12956);
xor U14174 (N_14174,N_13296,N_12212);
nand U14175 (N_14175,N_13433,N_13285);
and U14176 (N_14176,N_12781,N_13150);
nor U14177 (N_14177,N_12459,N_12721);
or U14178 (N_14178,N_12302,N_13358);
or U14179 (N_14179,N_12625,N_12042);
or U14180 (N_14180,N_12925,N_12596);
and U14181 (N_14181,N_12486,N_12451);
xnor U14182 (N_14182,N_12597,N_12638);
nand U14183 (N_14183,N_12849,N_12528);
nor U14184 (N_14184,N_12499,N_12792);
nor U14185 (N_14185,N_12885,N_12455);
nor U14186 (N_14186,N_12509,N_13149);
or U14187 (N_14187,N_12760,N_12007);
xnor U14188 (N_14188,N_12896,N_12711);
or U14189 (N_14189,N_12234,N_12608);
and U14190 (N_14190,N_12050,N_13291);
nand U14191 (N_14191,N_13488,N_13205);
and U14192 (N_14192,N_12122,N_12305);
nand U14193 (N_14193,N_12357,N_12742);
nand U14194 (N_14194,N_12384,N_13412);
and U14195 (N_14195,N_12818,N_13283);
and U14196 (N_14196,N_12468,N_12328);
and U14197 (N_14197,N_12210,N_13262);
nor U14198 (N_14198,N_12571,N_13392);
or U14199 (N_14199,N_12544,N_13318);
and U14200 (N_14200,N_12307,N_12836);
nand U14201 (N_14201,N_13221,N_12277);
and U14202 (N_14202,N_12969,N_12292);
or U14203 (N_14203,N_13372,N_13183);
or U14204 (N_14204,N_12839,N_13483);
nor U14205 (N_14205,N_12889,N_12949);
or U14206 (N_14206,N_12564,N_13403);
nor U14207 (N_14207,N_12853,N_12710);
and U14208 (N_14208,N_13485,N_13142);
nand U14209 (N_14209,N_13271,N_13174);
and U14210 (N_14210,N_13042,N_12203);
xnor U14211 (N_14211,N_12139,N_12355);
and U14212 (N_14212,N_13478,N_12634);
or U14213 (N_14213,N_13347,N_12338);
xor U14214 (N_14214,N_12713,N_13191);
nand U14215 (N_14215,N_12191,N_12605);
nand U14216 (N_14216,N_12973,N_13105);
xnor U14217 (N_14217,N_12040,N_12547);
nor U14218 (N_14218,N_13332,N_12128);
xor U14219 (N_14219,N_12958,N_12735);
or U14220 (N_14220,N_12636,N_12453);
or U14221 (N_14221,N_12733,N_12761);
nand U14222 (N_14222,N_12103,N_13132);
or U14223 (N_14223,N_12825,N_12221);
nor U14224 (N_14224,N_12223,N_12045);
or U14225 (N_14225,N_13071,N_12856);
or U14226 (N_14226,N_12100,N_12322);
xor U14227 (N_14227,N_12565,N_12156);
or U14228 (N_14228,N_13061,N_13349);
nor U14229 (N_14229,N_12296,N_12208);
xor U14230 (N_14230,N_13348,N_13015);
xnor U14231 (N_14231,N_12061,N_13327);
xor U14232 (N_14232,N_12387,N_12401);
and U14233 (N_14233,N_12256,N_13197);
nand U14234 (N_14234,N_12946,N_13044);
nand U14235 (N_14235,N_12109,N_12595);
nor U14236 (N_14236,N_12630,N_12318);
and U14237 (N_14237,N_13281,N_12324);
nor U14238 (N_14238,N_13404,N_12154);
or U14239 (N_14239,N_12021,N_12078);
xor U14240 (N_14240,N_12104,N_13442);
nor U14241 (N_14241,N_12266,N_12587);
or U14242 (N_14242,N_12249,N_12800);
nor U14243 (N_14243,N_12619,N_13261);
nand U14244 (N_14244,N_12490,N_13219);
xnor U14245 (N_14245,N_12655,N_13209);
nand U14246 (N_14246,N_12491,N_13484);
and U14247 (N_14247,N_13067,N_12906);
nor U14248 (N_14248,N_12678,N_13021);
nand U14249 (N_14249,N_12180,N_12291);
nand U14250 (N_14250,N_12063,N_12444);
and U14251 (N_14251,N_12738,N_12356);
nand U14252 (N_14252,N_12776,N_12850);
nor U14253 (N_14253,N_13272,N_12541);
xnor U14254 (N_14254,N_12231,N_13224);
and U14255 (N_14255,N_13470,N_13001);
nand U14256 (N_14256,N_12604,N_13168);
nand U14257 (N_14257,N_12324,N_12813);
nand U14258 (N_14258,N_13194,N_13255);
and U14259 (N_14259,N_12173,N_12827);
nor U14260 (N_14260,N_12084,N_12331);
or U14261 (N_14261,N_13173,N_12803);
nor U14262 (N_14262,N_13218,N_12229);
or U14263 (N_14263,N_12095,N_13157);
xnor U14264 (N_14264,N_12147,N_13322);
and U14265 (N_14265,N_12950,N_12490);
or U14266 (N_14266,N_13445,N_12483);
nand U14267 (N_14267,N_12636,N_12167);
or U14268 (N_14268,N_12038,N_12058);
nand U14269 (N_14269,N_12386,N_12286);
and U14270 (N_14270,N_12435,N_13065);
and U14271 (N_14271,N_12719,N_12880);
nor U14272 (N_14272,N_13446,N_13306);
nor U14273 (N_14273,N_12586,N_12443);
xnor U14274 (N_14274,N_12063,N_12883);
and U14275 (N_14275,N_12044,N_13032);
and U14276 (N_14276,N_13121,N_12491);
nor U14277 (N_14277,N_12406,N_12952);
nor U14278 (N_14278,N_12254,N_13113);
xor U14279 (N_14279,N_13232,N_12175);
and U14280 (N_14280,N_12614,N_12967);
and U14281 (N_14281,N_12725,N_12216);
and U14282 (N_14282,N_12607,N_12537);
and U14283 (N_14283,N_13266,N_12927);
nor U14284 (N_14284,N_12381,N_12449);
nor U14285 (N_14285,N_13413,N_13418);
nand U14286 (N_14286,N_13398,N_13437);
xor U14287 (N_14287,N_12442,N_12809);
or U14288 (N_14288,N_12083,N_12753);
and U14289 (N_14289,N_12719,N_12863);
nor U14290 (N_14290,N_13405,N_13057);
nand U14291 (N_14291,N_12873,N_13026);
xor U14292 (N_14292,N_13106,N_12253);
xor U14293 (N_14293,N_13352,N_12879);
and U14294 (N_14294,N_12950,N_12774);
nor U14295 (N_14295,N_13168,N_12185);
nor U14296 (N_14296,N_12640,N_13447);
or U14297 (N_14297,N_12641,N_12960);
nor U14298 (N_14298,N_12583,N_12296);
nor U14299 (N_14299,N_13184,N_12028);
nand U14300 (N_14300,N_12907,N_13402);
and U14301 (N_14301,N_13356,N_12799);
xnor U14302 (N_14302,N_12457,N_12324);
nand U14303 (N_14303,N_12726,N_12565);
or U14304 (N_14304,N_13041,N_12572);
nor U14305 (N_14305,N_12954,N_12985);
xnor U14306 (N_14306,N_13398,N_13180);
nand U14307 (N_14307,N_13154,N_12800);
or U14308 (N_14308,N_12297,N_12956);
and U14309 (N_14309,N_12259,N_13323);
xor U14310 (N_14310,N_12874,N_12894);
nor U14311 (N_14311,N_12702,N_12663);
xnor U14312 (N_14312,N_12696,N_12686);
and U14313 (N_14313,N_12257,N_12449);
nor U14314 (N_14314,N_12232,N_12935);
nor U14315 (N_14315,N_12426,N_13168);
nand U14316 (N_14316,N_12123,N_12356);
xor U14317 (N_14317,N_13401,N_12546);
nor U14318 (N_14318,N_12366,N_12359);
nor U14319 (N_14319,N_12456,N_12351);
nand U14320 (N_14320,N_13068,N_12247);
xnor U14321 (N_14321,N_12728,N_12407);
xor U14322 (N_14322,N_12383,N_13308);
xor U14323 (N_14323,N_13066,N_13153);
or U14324 (N_14324,N_12056,N_12328);
and U14325 (N_14325,N_12870,N_12880);
or U14326 (N_14326,N_12175,N_13469);
nand U14327 (N_14327,N_13418,N_12196);
nand U14328 (N_14328,N_12098,N_13117);
nor U14329 (N_14329,N_12179,N_12632);
nor U14330 (N_14330,N_12326,N_12930);
nor U14331 (N_14331,N_12899,N_12895);
nor U14332 (N_14332,N_12279,N_13017);
and U14333 (N_14333,N_13291,N_12454);
or U14334 (N_14334,N_12062,N_13159);
nor U14335 (N_14335,N_13462,N_13247);
nand U14336 (N_14336,N_12635,N_13062);
nor U14337 (N_14337,N_12199,N_12716);
or U14338 (N_14338,N_13369,N_13103);
nor U14339 (N_14339,N_12815,N_13313);
xnor U14340 (N_14340,N_13369,N_12783);
xnor U14341 (N_14341,N_13172,N_13128);
nor U14342 (N_14342,N_12613,N_12629);
xnor U14343 (N_14343,N_12324,N_12215);
xor U14344 (N_14344,N_12407,N_13183);
nand U14345 (N_14345,N_12977,N_13497);
nand U14346 (N_14346,N_13074,N_12500);
or U14347 (N_14347,N_12784,N_13161);
or U14348 (N_14348,N_13151,N_12495);
and U14349 (N_14349,N_13363,N_12922);
and U14350 (N_14350,N_12146,N_12165);
xor U14351 (N_14351,N_13190,N_12903);
xnor U14352 (N_14352,N_12024,N_12726);
nand U14353 (N_14353,N_13186,N_13335);
and U14354 (N_14354,N_12989,N_12964);
nor U14355 (N_14355,N_13228,N_13122);
nand U14356 (N_14356,N_13156,N_13045);
and U14357 (N_14357,N_12712,N_12756);
nand U14358 (N_14358,N_12706,N_12987);
nor U14359 (N_14359,N_12141,N_12057);
xnor U14360 (N_14360,N_12179,N_12207);
xor U14361 (N_14361,N_12120,N_12608);
xor U14362 (N_14362,N_12390,N_12666);
xnor U14363 (N_14363,N_13004,N_13285);
nand U14364 (N_14364,N_12994,N_12893);
and U14365 (N_14365,N_13334,N_12873);
xor U14366 (N_14366,N_13009,N_13256);
or U14367 (N_14367,N_13031,N_12699);
xnor U14368 (N_14368,N_13231,N_12888);
xor U14369 (N_14369,N_12385,N_13417);
nor U14370 (N_14370,N_12227,N_13035);
nor U14371 (N_14371,N_12835,N_12602);
nor U14372 (N_14372,N_12304,N_12482);
nor U14373 (N_14373,N_12927,N_12395);
and U14374 (N_14374,N_12604,N_12405);
and U14375 (N_14375,N_12313,N_13052);
xnor U14376 (N_14376,N_12295,N_13145);
or U14377 (N_14377,N_12698,N_13132);
xor U14378 (N_14378,N_13023,N_12381);
and U14379 (N_14379,N_13218,N_12628);
or U14380 (N_14380,N_13274,N_12273);
or U14381 (N_14381,N_13215,N_13151);
nand U14382 (N_14382,N_13161,N_12005);
xnor U14383 (N_14383,N_12847,N_12758);
or U14384 (N_14384,N_12814,N_12341);
nand U14385 (N_14385,N_12374,N_12074);
and U14386 (N_14386,N_12788,N_12210);
nand U14387 (N_14387,N_12766,N_12006);
and U14388 (N_14388,N_12575,N_13357);
or U14389 (N_14389,N_12945,N_13390);
nor U14390 (N_14390,N_12984,N_13260);
and U14391 (N_14391,N_12702,N_12346);
nand U14392 (N_14392,N_12845,N_13340);
nor U14393 (N_14393,N_12458,N_12337);
and U14394 (N_14394,N_13132,N_12209);
or U14395 (N_14395,N_12573,N_13103);
nand U14396 (N_14396,N_13221,N_12158);
xnor U14397 (N_14397,N_12516,N_12285);
and U14398 (N_14398,N_12660,N_13017);
and U14399 (N_14399,N_13027,N_12228);
or U14400 (N_14400,N_13294,N_12959);
or U14401 (N_14401,N_12650,N_12832);
nor U14402 (N_14402,N_12577,N_13208);
nor U14403 (N_14403,N_12857,N_13003);
nand U14404 (N_14404,N_12399,N_13493);
nand U14405 (N_14405,N_12125,N_13352);
or U14406 (N_14406,N_12694,N_12451);
xnor U14407 (N_14407,N_13288,N_13462);
nand U14408 (N_14408,N_12645,N_12863);
or U14409 (N_14409,N_12233,N_12699);
nor U14410 (N_14410,N_12884,N_12455);
nand U14411 (N_14411,N_12696,N_13239);
xnor U14412 (N_14412,N_13273,N_12074);
and U14413 (N_14413,N_12082,N_12855);
xor U14414 (N_14414,N_13077,N_13418);
nor U14415 (N_14415,N_12869,N_13013);
or U14416 (N_14416,N_12317,N_12331);
xor U14417 (N_14417,N_13174,N_12897);
nor U14418 (N_14418,N_13279,N_13208);
nor U14419 (N_14419,N_12262,N_12747);
or U14420 (N_14420,N_13038,N_13235);
or U14421 (N_14421,N_12361,N_12216);
nor U14422 (N_14422,N_13212,N_13013);
or U14423 (N_14423,N_12147,N_12652);
or U14424 (N_14424,N_12210,N_13335);
nor U14425 (N_14425,N_12123,N_12308);
or U14426 (N_14426,N_13174,N_12384);
xor U14427 (N_14427,N_12698,N_12697);
nor U14428 (N_14428,N_12542,N_13315);
nand U14429 (N_14429,N_12091,N_12026);
xor U14430 (N_14430,N_12381,N_13294);
and U14431 (N_14431,N_12534,N_13061);
nand U14432 (N_14432,N_12250,N_12137);
nand U14433 (N_14433,N_13288,N_13382);
nor U14434 (N_14434,N_12423,N_12765);
xor U14435 (N_14435,N_12637,N_12427);
xnor U14436 (N_14436,N_12005,N_12666);
xnor U14437 (N_14437,N_13354,N_12768);
xor U14438 (N_14438,N_12669,N_12404);
xor U14439 (N_14439,N_12064,N_12606);
xor U14440 (N_14440,N_12430,N_12733);
nand U14441 (N_14441,N_13080,N_12804);
xnor U14442 (N_14442,N_12607,N_13359);
or U14443 (N_14443,N_12191,N_12810);
and U14444 (N_14444,N_12832,N_13116);
nor U14445 (N_14445,N_13127,N_12738);
nor U14446 (N_14446,N_12650,N_12779);
and U14447 (N_14447,N_12162,N_12471);
and U14448 (N_14448,N_12375,N_13123);
xnor U14449 (N_14449,N_13410,N_12311);
and U14450 (N_14450,N_13489,N_12724);
and U14451 (N_14451,N_12076,N_13149);
and U14452 (N_14452,N_12787,N_12622);
or U14453 (N_14453,N_13310,N_12781);
xor U14454 (N_14454,N_12757,N_12048);
nor U14455 (N_14455,N_13292,N_13467);
and U14456 (N_14456,N_13363,N_13035);
nand U14457 (N_14457,N_13371,N_13017);
nand U14458 (N_14458,N_12424,N_12760);
nand U14459 (N_14459,N_12370,N_12487);
nand U14460 (N_14460,N_12686,N_13088);
nand U14461 (N_14461,N_13039,N_12044);
or U14462 (N_14462,N_12385,N_12977);
or U14463 (N_14463,N_12320,N_13435);
and U14464 (N_14464,N_12875,N_12581);
and U14465 (N_14465,N_12471,N_12590);
xor U14466 (N_14466,N_13164,N_12877);
and U14467 (N_14467,N_12215,N_12927);
or U14468 (N_14468,N_13145,N_13423);
xor U14469 (N_14469,N_12654,N_13366);
nand U14470 (N_14470,N_13483,N_12979);
or U14471 (N_14471,N_12303,N_13166);
nor U14472 (N_14472,N_12301,N_12609);
nand U14473 (N_14473,N_13445,N_12170);
or U14474 (N_14474,N_12827,N_12944);
nand U14475 (N_14475,N_12118,N_12595);
nor U14476 (N_14476,N_12718,N_12161);
xnor U14477 (N_14477,N_13349,N_12633);
and U14478 (N_14478,N_13222,N_12678);
and U14479 (N_14479,N_12665,N_12530);
nand U14480 (N_14480,N_13410,N_13352);
nor U14481 (N_14481,N_13254,N_12247);
xor U14482 (N_14482,N_12940,N_13410);
and U14483 (N_14483,N_13451,N_12471);
xnor U14484 (N_14484,N_12735,N_12767);
nand U14485 (N_14485,N_13362,N_12797);
nand U14486 (N_14486,N_12902,N_13405);
or U14487 (N_14487,N_12401,N_12369);
nand U14488 (N_14488,N_12024,N_12758);
or U14489 (N_14489,N_13218,N_13102);
or U14490 (N_14490,N_13262,N_12302);
nand U14491 (N_14491,N_13105,N_12729);
or U14492 (N_14492,N_12363,N_12670);
nor U14493 (N_14493,N_13119,N_13117);
and U14494 (N_14494,N_12425,N_12914);
nand U14495 (N_14495,N_12785,N_12893);
nor U14496 (N_14496,N_12493,N_12191);
xor U14497 (N_14497,N_12156,N_12670);
nand U14498 (N_14498,N_13044,N_12004);
or U14499 (N_14499,N_12256,N_12798);
nand U14500 (N_14500,N_12009,N_12629);
or U14501 (N_14501,N_12072,N_12611);
xor U14502 (N_14502,N_12164,N_12792);
and U14503 (N_14503,N_12338,N_12177);
or U14504 (N_14504,N_13371,N_13169);
xor U14505 (N_14505,N_12953,N_13418);
xnor U14506 (N_14506,N_13356,N_13083);
or U14507 (N_14507,N_13197,N_13280);
and U14508 (N_14508,N_12319,N_12502);
nor U14509 (N_14509,N_12136,N_12297);
nor U14510 (N_14510,N_13275,N_13204);
nand U14511 (N_14511,N_13256,N_12624);
xnor U14512 (N_14512,N_13434,N_12995);
nor U14513 (N_14513,N_12705,N_12937);
and U14514 (N_14514,N_12216,N_12902);
nor U14515 (N_14515,N_12689,N_13162);
or U14516 (N_14516,N_12770,N_12741);
or U14517 (N_14517,N_12887,N_13082);
and U14518 (N_14518,N_12726,N_13129);
nand U14519 (N_14519,N_12226,N_13284);
and U14520 (N_14520,N_12094,N_13437);
xnor U14521 (N_14521,N_12728,N_12835);
nor U14522 (N_14522,N_12034,N_12268);
xnor U14523 (N_14523,N_13022,N_13108);
nand U14524 (N_14524,N_12223,N_13244);
xor U14525 (N_14525,N_12147,N_12855);
nor U14526 (N_14526,N_12541,N_12117);
nand U14527 (N_14527,N_13400,N_12419);
and U14528 (N_14528,N_12178,N_12835);
xor U14529 (N_14529,N_12538,N_12139);
nand U14530 (N_14530,N_12172,N_12987);
nor U14531 (N_14531,N_12049,N_12955);
nand U14532 (N_14532,N_12068,N_12852);
nor U14533 (N_14533,N_13423,N_12823);
and U14534 (N_14534,N_12237,N_13204);
nand U14535 (N_14535,N_13195,N_12274);
and U14536 (N_14536,N_12334,N_12202);
or U14537 (N_14537,N_12260,N_12701);
and U14538 (N_14538,N_13362,N_12101);
or U14539 (N_14539,N_13090,N_12608);
nor U14540 (N_14540,N_12441,N_13082);
xnor U14541 (N_14541,N_12398,N_12326);
nor U14542 (N_14542,N_12751,N_12977);
xnor U14543 (N_14543,N_13347,N_12900);
nor U14544 (N_14544,N_12385,N_13197);
nand U14545 (N_14545,N_12699,N_12297);
or U14546 (N_14546,N_12055,N_13344);
or U14547 (N_14547,N_12362,N_12246);
and U14548 (N_14548,N_13421,N_12331);
nand U14549 (N_14549,N_13415,N_12006);
and U14550 (N_14550,N_12240,N_13274);
xor U14551 (N_14551,N_12529,N_13055);
xnor U14552 (N_14552,N_12438,N_12786);
and U14553 (N_14553,N_13322,N_12986);
nor U14554 (N_14554,N_13383,N_12024);
xor U14555 (N_14555,N_12854,N_12934);
or U14556 (N_14556,N_12839,N_12452);
xor U14557 (N_14557,N_12308,N_12737);
or U14558 (N_14558,N_12701,N_13119);
and U14559 (N_14559,N_13074,N_12588);
xnor U14560 (N_14560,N_13037,N_12719);
and U14561 (N_14561,N_13085,N_12364);
and U14562 (N_14562,N_12659,N_12080);
nand U14563 (N_14563,N_12107,N_12022);
nand U14564 (N_14564,N_13415,N_12865);
and U14565 (N_14565,N_12881,N_12650);
and U14566 (N_14566,N_13330,N_12257);
nor U14567 (N_14567,N_13173,N_13459);
and U14568 (N_14568,N_12492,N_13083);
and U14569 (N_14569,N_12271,N_13192);
and U14570 (N_14570,N_12099,N_13454);
and U14571 (N_14571,N_12238,N_13427);
xnor U14572 (N_14572,N_12206,N_12920);
xor U14573 (N_14573,N_12618,N_12385);
nor U14574 (N_14574,N_12076,N_13452);
nand U14575 (N_14575,N_12241,N_12833);
xnor U14576 (N_14576,N_12487,N_12586);
and U14577 (N_14577,N_12814,N_12369);
nand U14578 (N_14578,N_12742,N_12747);
and U14579 (N_14579,N_12786,N_13016);
nor U14580 (N_14580,N_12594,N_12499);
nand U14581 (N_14581,N_12309,N_13049);
nor U14582 (N_14582,N_12957,N_12052);
xor U14583 (N_14583,N_13303,N_12399);
nor U14584 (N_14584,N_12705,N_13064);
nand U14585 (N_14585,N_12380,N_13402);
and U14586 (N_14586,N_13373,N_12960);
or U14587 (N_14587,N_12190,N_12516);
or U14588 (N_14588,N_12751,N_12883);
or U14589 (N_14589,N_13078,N_12817);
and U14590 (N_14590,N_12352,N_12762);
or U14591 (N_14591,N_12755,N_12122);
and U14592 (N_14592,N_12133,N_12729);
and U14593 (N_14593,N_12865,N_12769);
nand U14594 (N_14594,N_13278,N_13070);
nor U14595 (N_14595,N_12712,N_13185);
nor U14596 (N_14596,N_13250,N_12306);
or U14597 (N_14597,N_12179,N_13194);
nor U14598 (N_14598,N_13078,N_12035);
nor U14599 (N_14599,N_13138,N_12388);
or U14600 (N_14600,N_13149,N_13314);
nor U14601 (N_14601,N_13445,N_12255);
or U14602 (N_14602,N_13120,N_13288);
xor U14603 (N_14603,N_12048,N_12684);
and U14604 (N_14604,N_13085,N_12182);
nand U14605 (N_14605,N_13342,N_12690);
nand U14606 (N_14606,N_12210,N_12389);
nor U14607 (N_14607,N_12579,N_13260);
or U14608 (N_14608,N_12065,N_12378);
nand U14609 (N_14609,N_12363,N_13382);
and U14610 (N_14610,N_12819,N_12492);
and U14611 (N_14611,N_12177,N_12942);
xor U14612 (N_14612,N_12040,N_12518);
and U14613 (N_14613,N_12286,N_13181);
and U14614 (N_14614,N_12288,N_12139);
xnor U14615 (N_14615,N_13255,N_12517);
or U14616 (N_14616,N_12437,N_12543);
nor U14617 (N_14617,N_13153,N_13291);
nor U14618 (N_14618,N_12579,N_12953);
xor U14619 (N_14619,N_13036,N_13456);
xor U14620 (N_14620,N_12489,N_12676);
xnor U14621 (N_14621,N_13030,N_12363);
xor U14622 (N_14622,N_12859,N_12604);
and U14623 (N_14623,N_13040,N_13227);
nor U14624 (N_14624,N_12998,N_12157);
or U14625 (N_14625,N_13276,N_12520);
nand U14626 (N_14626,N_12785,N_12133);
xor U14627 (N_14627,N_13326,N_12175);
nand U14628 (N_14628,N_12084,N_12284);
nand U14629 (N_14629,N_13280,N_12912);
nor U14630 (N_14630,N_13353,N_13125);
or U14631 (N_14631,N_12001,N_12676);
nor U14632 (N_14632,N_12218,N_12394);
nor U14633 (N_14633,N_12716,N_12873);
xor U14634 (N_14634,N_12195,N_12817);
and U14635 (N_14635,N_12699,N_13102);
and U14636 (N_14636,N_12166,N_12998);
nor U14637 (N_14637,N_12098,N_12067);
and U14638 (N_14638,N_12924,N_12998);
nand U14639 (N_14639,N_12619,N_12106);
or U14640 (N_14640,N_12794,N_12643);
xor U14641 (N_14641,N_13162,N_13379);
xnor U14642 (N_14642,N_12909,N_12654);
and U14643 (N_14643,N_12791,N_12704);
and U14644 (N_14644,N_12953,N_12813);
xnor U14645 (N_14645,N_12823,N_12065);
xnor U14646 (N_14646,N_12020,N_12957);
nor U14647 (N_14647,N_12514,N_12352);
xor U14648 (N_14648,N_12179,N_12133);
and U14649 (N_14649,N_12587,N_13476);
nand U14650 (N_14650,N_12441,N_12457);
xor U14651 (N_14651,N_12304,N_13012);
nor U14652 (N_14652,N_12101,N_12016);
nor U14653 (N_14653,N_12853,N_12488);
or U14654 (N_14654,N_13073,N_12264);
xnor U14655 (N_14655,N_13237,N_12101);
or U14656 (N_14656,N_12088,N_13359);
and U14657 (N_14657,N_12875,N_12489);
nand U14658 (N_14658,N_13282,N_13124);
xnor U14659 (N_14659,N_13004,N_13353);
and U14660 (N_14660,N_12586,N_12172);
nand U14661 (N_14661,N_12102,N_12553);
nor U14662 (N_14662,N_12389,N_13267);
xor U14663 (N_14663,N_12889,N_12005);
nand U14664 (N_14664,N_12628,N_12294);
or U14665 (N_14665,N_13187,N_12227);
or U14666 (N_14666,N_12988,N_12215);
and U14667 (N_14667,N_12024,N_12995);
xor U14668 (N_14668,N_13064,N_13179);
and U14669 (N_14669,N_12600,N_13294);
nand U14670 (N_14670,N_13220,N_12582);
or U14671 (N_14671,N_12204,N_12782);
nor U14672 (N_14672,N_13336,N_12551);
xor U14673 (N_14673,N_12203,N_12039);
xnor U14674 (N_14674,N_12334,N_12274);
nor U14675 (N_14675,N_12459,N_12361);
xor U14676 (N_14676,N_13429,N_12105);
xor U14677 (N_14677,N_12671,N_13410);
xnor U14678 (N_14678,N_12439,N_12955);
nand U14679 (N_14679,N_13005,N_12636);
nand U14680 (N_14680,N_12213,N_13415);
and U14681 (N_14681,N_12285,N_12688);
nand U14682 (N_14682,N_12694,N_13018);
and U14683 (N_14683,N_12362,N_12028);
nor U14684 (N_14684,N_12072,N_12599);
and U14685 (N_14685,N_13488,N_12675);
or U14686 (N_14686,N_13094,N_12764);
nand U14687 (N_14687,N_12814,N_12535);
nor U14688 (N_14688,N_12144,N_13102);
or U14689 (N_14689,N_12347,N_12206);
xor U14690 (N_14690,N_12793,N_12630);
nor U14691 (N_14691,N_12491,N_12675);
xor U14692 (N_14692,N_12448,N_13442);
xnor U14693 (N_14693,N_12267,N_12400);
xor U14694 (N_14694,N_12071,N_13172);
nor U14695 (N_14695,N_13362,N_12271);
xor U14696 (N_14696,N_12055,N_12359);
nor U14697 (N_14697,N_13141,N_12266);
and U14698 (N_14698,N_12736,N_12287);
and U14699 (N_14699,N_13356,N_12094);
nor U14700 (N_14700,N_12945,N_12069);
and U14701 (N_14701,N_13135,N_13365);
nor U14702 (N_14702,N_12941,N_12279);
or U14703 (N_14703,N_12179,N_12829);
xor U14704 (N_14704,N_12566,N_12014);
nor U14705 (N_14705,N_12278,N_12622);
xnor U14706 (N_14706,N_12516,N_13353);
nand U14707 (N_14707,N_13162,N_12587);
nor U14708 (N_14708,N_12767,N_13154);
xor U14709 (N_14709,N_12845,N_13492);
nor U14710 (N_14710,N_12582,N_13160);
xnor U14711 (N_14711,N_12190,N_12370);
nand U14712 (N_14712,N_12473,N_12060);
and U14713 (N_14713,N_13456,N_12242);
nand U14714 (N_14714,N_13254,N_13316);
nor U14715 (N_14715,N_13275,N_13126);
and U14716 (N_14716,N_13363,N_12965);
nand U14717 (N_14717,N_12304,N_12948);
and U14718 (N_14718,N_12779,N_12346);
xor U14719 (N_14719,N_12803,N_12361);
or U14720 (N_14720,N_12392,N_12267);
nand U14721 (N_14721,N_13289,N_12344);
nand U14722 (N_14722,N_12684,N_12403);
xnor U14723 (N_14723,N_12169,N_13380);
and U14724 (N_14724,N_13264,N_12818);
nor U14725 (N_14725,N_12111,N_12741);
xor U14726 (N_14726,N_12056,N_12590);
nor U14727 (N_14727,N_13421,N_12439);
nand U14728 (N_14728,N_12461,N_13195);
xor U14729 (N_14729,N_12505,N_12486);
and U14730 (N_14730,N_13115,N_13081);
nand U14731 (N_14731,N_12596,N_12654);
xnor U14732 (N_14732,N_12152,N_12694);
or U14733 (N_14733,N_13121,N_13368);
nand U14734 (N_14734,N_12481,N_12985);
nor U14735 (N_14735,N_13458,N_13066);
and U14736 (N_14736,N_13173,N_12179);
xnor U14737 (N_14737,N_12078,N_12056);
nand U14738 (N_14738,N_13432,N_13191);
nand U14739 (N_14739,N_12534,N_12543);
xor U14740 (N_14740,N_13216,N_12114);
xnor U14741 (N_14741,N_12263,N_12255);
nand U14742 (N_14742,N_13205,N_12349);
or U14743 (N_14743,N_12707,N_13078);
nand U14744 (N_14744,N_12148,N_13000);
nand U14745 (N_14745,N_13370,N_13107);
xor U14746 (N_14746,N_12111,N_12821);
nand U14747 (N_14747,N_13009,N_13493);
xnor U14748 (N_14748,N_12989,N_13055);
or U14749 (N_14749,N_12609,N_12478);
or U14750 (N_14750,N_12591,N_12341);
nand U14751 (N_14751,N_13116,N_12948);
and U14752 (N_14752,N_12042,N_12925);
nor U14753 (N_14753,N_13025,N_12729);
or U14754 (N_14754,N_13113,N_12046);
xor U14755 (N_14755,N_12980,N_13394);
and U14756 (N_14756,N_13153,N_12170);
nor U14757 (N_14757,N_12893,N_12674);
nand U14758 (N_14758,N_12570,N_12303);
and U14759 (N_14759,N_12049,N_12626);
and U14760 (N_14760,N_12298,N_13196);
nand U14761 (N_14761,N_13258,N_12147);
xnor U14762 (N_14762,N_13107,N_13258);
xor U14763 (N_14763,N_12933,N_12307);
xor U14764 (N_14764,N_12968,N_12599);
nor U14765 (N_14765,N_12858,N_12837);
or U14766 (N_14766,N_12160,N_12687);
nor U14767 (N_14767,N_13311,N_13250);
or U14768 (N_14768,N_12126,N_12178);
and U14769 (N_14769,N_13093,N_12205);
nand U14770 (N_14770,N_13284,N_12252);
xnor U14771 (N_14771,N_12934,N_12771);
or U14772 (N_14772,N_13004,N_12708);
or U14773 (N_14773,N_12753,N_13417);
or U14774 (N_14774,N_12318,N_12355);
or U14775 (N_14775,N_12706,N_13100);
nand U14776 (N_14776,N_13405,N_13314);
xnor U14777 (N_14777,N_12442,N_13330);
xnor U14778 (N_14778,N_13111,N_12629);
nand U14779 (N_14779,N_12542,N_12157);
or U14780 (N_14780,N_13486,N_12643);
nand U14781 (N_14781,N_12461,N_12342);
and U14782 (N_14782,N_12240,N_12192);
xnor U14783 (N_14783,N_13260,N_13285);
nand U14784 (N_14784,N_13492,N_12672);
nand U14785 (N_14785,N_12735,N_12498);
nor U14786 (N_14786,N_12354,N_12325);
or U14787 (N_14787,N_13312,N_12480);
xnor U14788 (N_14788,N_12415,N_12848);
xor U14789 (N_14789,N_12642,N_12801);
nand U14790 (N_14790,N_12516,N_12251);
and U14791 (N_14791,N_12171,N_12807);
nor U14792 (N_14792,N_12581,N_12890);
xor U14793 (N_14793,N_12128,N_12282);
nor U14794 (N_14794,N_13138,N_12070);
xnor U14795 (N_14795,N_12010,N_12607);
nor U14796 (N_14796,N_13146,N_13169);
and U14797 (N_14797,N_12013,N_13327);
nand U14798 (N_14798,N_13383,N_12536);
nand U14799 (N_14799,N_12757,N_12287);
nor U14800 (N_14800,N_12411,N_12233);
xnor U14801 (N_14801,N_12832,N_12860);
or U14802 (N_14802,N_12186,N_12258);
nand U14803 (N_14803,N_12107,N_12858);
or U14804 (N_14804,N_13308,N_12118);
nor U14805 (N_14805,N_12518,N_12096);
or U14806 (N_14806,N_13016,N_12056);
or U14807 (N_14807,N_12141,N_13370);
nor U14808 (N_14808,N_12706,N_12618);
nand U14809 (N_14809,N_12378,N_12441);
nor U14810 (N_14810,N_12306,N_12919);
nor U14811 (N_14811,N_12807,N_13114);
or U14812 (N_14812,N_12207,N_12056);
xor U14813 (N_14813,N_13340,N_12125);
or U14814 (N_14814,N_12915,N_13460);
or U14815 (N_14815,N_12432,N_12186);
nand U14816 (N_14816,N_12137,N_13198);
and U14817 (N_14817,N_12208,N_12979);
xor U14818 (N_14818,N_13392,N_12191);
nor U14819 (N_14819,N_12519,N_13173);
or U14820 (N_14820,N_12546,N_13150);
xor U14821 (N_14821,N_13239,N_12283);
or U14822 (N_14822,N_12043,N_13040);
nand U14823 (N_14823,N_12740,N_12410);
nor U14824 (N_14824,N_12352,N_12957);
and U14825 (N_14825,N_12391,N_13271);
nor U14826 (N_14826,N_12109,N_13403);
nor U14827 (N_14827,N_13184,N_12400);
and U14828 (N_14828,N_13016,N_12051);
nor U14829 (N_14829,N_12894,N_12984);
and U14830 (N_14830,N_12807,N_12936);
xor U14831 (N_14831,N_12940,N_12612);
and U14832 (N_14832,N_12383,N_13423);
xnor U14833 (N_14833,N_13328,N_12311);
and U14834 (N_14834,N_12479,N_12117);
nand U14835 (N_14835,N_13277,N_12050);
xor U14836 (N_14836,N_13072,N_12216);
and U14837 (N_14837,N_12289,N_13297);
or U14838 (N_14838,N_12947,N_12534);
nand U14839 (N_14839,N_13063,N_13025);
xor U14840 (N_14840,N_12776,N_12759);
nand U14841 (N_14841,N_12623,N_12217);
nor U14842 (N_14842,N_12098,N_13186);
and U14843 (N_14843,N_13055,N_12648);
and U14844 (N_14844,N_13263,N_12184);
nand U14845 (N_14845,N_13133,N_12179);
xnor U14846 (N_14846,N_12584,N_12692);
nor U14847 (N_14847,N_12304,N_13118);
nand U14848 (N_14848,N_12499,N_12416);
xor U14849 (N_14849,N_13331,N_13053);
nor U14850 (N_14850,N_12491,N_12994);
nor U14851 (N_14851,N_13122,N_13187);
nor U14852 (N_14852,N_12802,N_12682);
xor U14853 (N_14853,N_12100,N_12427);
or U14854 (N_14854,N_12345,N_13355);
nand U14855 (N_14855,N_12496,N_12825);
or U14856 (N_14856,N_12943,N_12798);
and U14857 (N_14857,N_12305,N_12201);
nand U14858 (N_14858,N_13400,N_12552);
or U14859 (N_14859,N_12478,N_12741);
and U14860 (N_14860,N_12162,N_12023);
nor U14861 (N_14861,N_13079,N_12014);
nand U14862 (N_14862,N_12101,N_12460);
nor U14863 (N_14863,N_12468,N_12951);
xor U14864 (N_14864,N_12294,N_13105);
xnor U14865 (N_14865,N_12959,N_12091);
or U14866 (N_14866,N_12423,N_12775);
or U14867 (N_14867,N_13027,N_12810);
and U14868 (N_14868,N_12564,N_12138);
xnor U14869 (N_14869,N_13432,N_12609);
nand U14870 (N_14870,N_12775,N_12366);
nor U14871 (N_14871,N_13138,N_12497);
xnor U14872 (N_14872,N_12464,N_12020);
and U14873 (N_14873,N_13465,N_12179);
nand U14874 (N_14874,N_13473,N_12388);
nor U14875 (N_14875,N_12431,N_12391);
xnor U14876 (N_14876,N_12141,N_12411);
and U14877 (N_14877,N_12424,N_12729);
xor U14878 (N_14878,N_13032,N_12038);
and U14879 (N_14879,N_12573,N_12886);
nand U14880 (N_14880,N_12020,N_12331);
or U14881 (N_14881,N_12524,N_13060);
xnor U14882 (N_14882,N_12280,N_12687);
or U14883 (N_14883,N_13441,N_12503);
nor U14884 (N_14884,N_12592,N_12756);
nor U14885 (N_14885,N_12119,N_12948);
nor U14886 (N_14886,N_13015,N_13255);
and U14887 (N_14887,N_12916,N_12514);
nand U14888 (N_14888,N_12445,N_13085);
nor U14889 (N_14889,N_13176,N_12701);
xor U14890 (N_14890,N_12709,N_12930);
xor U14891 (N_14891,N_12428,N_13157);
nor U14892 (N_14892,N_12425,N_12686);
xnor U14893 (N_14893,N_13024,N_13116);
xor U14894 (N_14894,N_12593,N_13190);
or U14895 (N_14895,N_12054,N_12561);
nor U14896 (N_14896,N_12140,N_12241);
xor U14897 (N_14897,N_13381,N_12588);
and U14898 (N_14898,N_13277,N_12094);
or U14899 (N_14899,N_13240,N_13023);
or U14900 (N_14900,N_12070,N_12993);
nor U14901 (N_14901,N_12918,N_12351);
nand U14902 (N_14902,N_12543,N_12981);
xnor U14903 (N_14903,N_12414,N_12556);
or U14904 (N_14904,N_12728,N_12068);
or U14905 (N_14905,N_13380,N_13431);
nor U14906 (N_14906,N_12677,N_12525);
nor U14907 (N_14907,N_12648,N_13036);
nand U14908 (N_14908,N_13235,N_12681);
nand U14909 (N_14909,N_13123,N_12463);
and U14910 (N_14910,N_12168,N_13325);
or U14911 (N_14911,N_12618,N_12445);
nor U14912 (N_14912,N_12163,N_12630);
nand U14913 (N_14913,N_13389,N_12133);
nand U14914 (N_14914,N_12583,N_12917);
xor U14915 (N_14915,N_12705,N_12038);
and U14916 (N_14916,N_12028,N_12293);
and U14917 (N_14917,N_12936,N_12233);
xor U14918 (N_14918,N_12549,N_12727);
xnor U14919 (N_14919,N_13332,N_12293);
nor U14920 (N_14920,N_12852,N_13084);
nand U14921 (N_14921,N_12574,N_13150);
and U14922 (N_14922,N_12032,N_13013);
nand U14923 (N_14923,N_12125,N_12941);
nand U14924 (N_14924,N_13031,N_12051);
or U14925 (N_14925,N_12378,N_12803);
or U14926 (N_14926,N_13475,N_13004);
and U14927 (N_14927,N_12164,N_13484);
xor U14928 (N_14928,N_13159,N_13034);
or U14929 (N_14929,N_12531,N_12566);
or U14930 (N_14930,N_13325,N_13370);
xnor U14931 (N_14931,N_12142,N_13373);
nand U14932 (N_14932,N_13229,N_13480);
nand U14933 (N_14933,N_12890,N_13380);
or U14934 (N_14934,N_12234,N_12277);
nor U14935 (N_14935,N_12956,N_12391);
xnor U14936 (N_14936,N_12419,N_12319);
xnor U14937 (N_14937,N_13012,N_13442);
xnor U14938 (N_14938,N_13447,N_13104);
nand U14939 (N_14939,N_13293,N_13435);
xor U14940 (N_14940,N_12864,N_12414);
nor U14941 (N_14941,N_12131,N_13256);
or U14942 (N_14942,N_12414,N_12713);
nor U14943 (N_14943,N_12587,N_13028);
or U14944 (N_14944,N_12326,N_12420);
nor U14945 (N_14945,N_12395,N_12034);
and U14946 (N_14946,N_12602,N_13276);
nor U14947 (N_14947,N_12251,N_12263);
xor U14948 (N_14948,N_13233,N_12616);
nand U14949 (N_14949,N_13011,N_13226);
or U14950 (N_14950,N_12773,N_12645);
xor U14951 (N_14951,N_12757,N_12899);
xnor U14952 (N_14952,N_12418,N_13267);
or U14953 (N_14953,N_12220,N_12199);
and U14954 (N_14954,N_12149,N_13483);
nand U14955 (N_14955,N_13065,N_13289);
nor U14956 (N_14956,N_12786,N_12848);
nand U14957 (N_14957,N_13344,N_12392);
or U14958 (N_14958,N_13425,N_13288);
nand U14959 (N_14959,N_12999,N_12524);
or U14960 (N_14960,N_12964,N_13423);
nor U14961 (N_14961,N_12114,N_12677);
or U14962 (N_14962,N_13136,N_12279);
nor U14963 (N_14963,N_13457,N_12924);
or U14964 (N_14964,N_12558,N_13264);
xor U14965 (N_14965,N_12169,N_12953);
xnor U14966 (N_14966,N_12906,N_12798);
and U14967 (N_14967,N_12774,N_12157);
xnor U14968 (N_14968,N_12757,N_12772);
and U14969 (N_14969,N_12529,N_12010);
and U14970 (N_14970,N_13017,N_12036);
and U14971 (N_14971,N_12463,N_13444);
nand U14972 (N_14972,N_12547,N_12988);
nand U14973 (N_14973,N_13484,N_13358);
or U14974 (N_14974,N_13329,N_12926);
xor U14975 (N_14975,N_12869,N_13014);
and U14976 (N_14976,N_12624,N_13463);
or U14977 (N_14977,N_12915,N_12225);
nor U14978 (N_14978,N_12470,N_13286);
xnor U14979 (N_14979,N_13209,N_13344);
or U14980 (N_14980,N_12826,N_12298);
and U14981 (N_14981,N_12550,N_13499);
xor U14982 (N_14982,N_13101,N_12417);
nand U14983 (N_14983,N_13439,N_13417);
or U14984 (N_14984,N_12934,N_12494);
xnor U14985 (N_14985,N_12289,N_12393);
nor U14986 (N_14986,N_12307,N_13158);
or U14987 (N_14987,N_12881,N_12047);
xnor U14988 (N_14988,N_12973,N_13400);
or U14989 (N_14989,N_12511,N_12748);
and U14990 (N_14990,N_12250,N_13119);
nand U14991 (N_14991,N_13070,N_12777);
xor U14992 (N_14992,N_12595,N_12900);
nand U14993 (N_14993,N_13080,N_13063);
or U14994 (N_14994,N_12907,N_12118);
xnor U14995 (N_14995,N_13461,N_13430);
or U14996 (N_14996,N_13455,N_13414);
nand U14997 (N_14997,N_12633,N_13262);
and U14998 (N_14998,N_12531,N_13083);
xnor U14999 (N_14999,N_12565,N_13476);
xor U15000 (N_15000,N_14192,N_14926);
xor U15001 (N_15001,N_13522,N_14576);
or U15002 (N_15002,N_14792,N_13643);
or U15003 (N_15003,N_13916,N_13551);
nor U15004 (N_15004,N_14168,N_14065);
or U15005 (N_15005,N_13568,N_13603);
nor U15006 (N_15006,N_14759,N_14656);
nor U15007 (N_15007,N_13515,N_14943);
nor U15008 (N_15008,N_14970,N_14379);
xnor U15009 (N_15009,N_14664,N_14446);
xnor U15010 (N_15010,N_14835,N_13820);
nor U15011 (N_15011,N_13783,N_14532);
or U15012 (N_15012,N_13656,N_14972);
and U15013 (N_15013,N_14208,N_14511);
and U15014 (N_15014,N_14851,N_14684);
or U15015 (N_15015,N_14639,N_13792);
nor U15016 (N_15016,N_14255,N_13553);
xnor U15017 (N_15017,N_14375,N_14782);
and U15018 (N_15018,N_13786,N_13833);
nor U15019 (N_15019,N_13529,N_14914);
nand U15020 (N_15020,N_13558,N_14003);
xnor U15021 (N_15021,N_14220,N_14384);
or U15022 (N_15022,N_14296,N_14070);
nand U15023 (N_15023,N_14510,N_13793);
xor U15024 (N_15024,N_13507,N_14572);
and U15025 (N_15025,N_14916,N_14424);
or U15026 (N_15026,N_13716,N_14597);
nand U15027 (N_15027,N_14527,N_13582);
nor U15028 (N_15028,N_13790,N_14534);
and U15029 (N_15029,N_13672,N_14956);
nand U15030 (N_15030,N_13858,N_14668);
nand U15031 (N_15031,N_13771,N_14740);
nand U15032 (N_15032,N_14377,N_14310);
and U15033 (N_15033,N_13687,N_13733);
or U15034 (N_15034,N_14921,N_13893);
xnor U15035 (N_15035,N_13794,N_14254);
and U15036 (N_15036,N_13729,N_13525);
or U15037 (N_15037,N_13676,N_14072);
and U15038 (N_15038,N_14177,N_14992);
and U15039 (N_15039,N_13599,N_14338);
and U15040 (N_15040,N_13514,N_14502);
or U15041 (N_15041,N_13964,N_13844);
or U15042 (N_15042,N_14867,N_14616);
and U15043 (N_15043,N_14725,N_14685);
or U15044 (N_15044,N_13500,N_14112);
or U15045 (N_15045,N_14876,N_14460);
and U15046 (N_15046,N_14928,N_13947);
nor U15047 (N_15047,N_14455,N_13696);
and U15048 (N_15048,N_13800,N_13879);
nand U15049 (N_15049,N_13978,N_13692);
nor U15050 (N_15050,N_13565,N_14425);
nor U15051 (N_15051,N_14710,N_13503);
nor U15052 (N_15052,N_14017,N_14577);
nor U15053 (N_15053,N_14433,N_14324);
and U15054 (N_15054,N_14204,N_14610);
or U15055 (N_15055,N_14404,N_14328);
nor U15056 (N_15056,N_14445,N_13691);
xnor U15057 (N_15057,N_13952,N_14189);
or U15058 (N_15058,N_14228,N_14669);
nand U15059 (N_15059,N_13695,N_13831);
nand U15060 (N_15060,N_14720,N_13632);
xnor U15061 (N_15061,N_14207,N_14562);
nor U15062 (N_15062,N_14804,N_14357);
and U15063 (N_15063,N_14183,N_14327);
xor U15064 (N_15064,N_14073,N_14233);
or U15065 (N_15065,N_14783,N_14627);
nor U15066 (N_15066,N_14487,N_14227);
xnor U15067 (N_15067,N_13910,N_14235);
nor U15068 (N_15068,N_14309,N_14631);
nor U15069 (N_15069,N_14093,N_14282);
or U15070 (N_15070,N_14146,N_13704);
and U15071 (N_15071,N_13639,N_14398);
nand U15072 (N_15072,N_13875,N_14981);
and U15073 (N_15073,N_14945,N_14621);
or U15074 (N_15074,N_13699,N_14909);
or U15075 (N_15075,N_14430,N_13864);
or U15076 (N_15076,N_13649,N_14880);
xnor U15077 (N_15077,N_14673,N_14524);
nor U15078 (N_15078,N_14801,N_13766);
nand U15079 (N_15079,N_14126,N_14193);
or U15080 (N_15080,N_13828,N_13606);
nor U15081 (N_15081,N_14142,N_14537);
nor U15082 (N_15082,N_13637,N_14078);
and U15083 (N_15083,N_14104,N_14300);
or U15084 (N_15084,N_14030,N_14137);
nand U15085 (N_15085,N_14677,N_13622);
nor U15086 (N_15086,N_14154,N_14733);
or U15087 (N_15087,N_14329,N_14251);
nand U15088 (N_15088,N_14226,N_13777);
and U15089 (N_15089,N_14635,N_14064);
or U15090 (N_15090,N_13521,N_13850);
and U15091 (N_15091,N_13872,N_14515);
xnor U15092 (N_15092,N_14658,N_13824);
and U15093 (N_15093,N_14596,N_14295);
nand U15094 (N_15094,N_14590,N_13636);
and U15095 (N_15095,N_13537,N_14859);
or U15096 (N_15096,N_14214,N_13905);
or U15097 (N_15097,N_14691,N_14431);
nor U15098 (N_15098,N_13818,N_14463);
or U15099 (N_15099,N_13907,N_14854);
nand U15100 (N_15100,N_13948,N_13690);
and U15101 (N_15101,N_14831,N_14202);
nand U15102 (N_15102,N_14195,N_13745);
nand U15103 (N_15103,N_13671,N_14369);
or U15104 (N_15104,N_13957,N_14780);
and U15105 (N_15105,N_13902,N_14151);
or U15106 (N_15106,N_14812,N_14931);
xnor U15107 (N_15107,N_14567,N_14418);
nand U15108 (N_15108,N_14018,N_13935);
xnor U15109 (N_15109,N_14185,N_14935);
and U15110 (N_15110,N_13886,N_14023);
xor U15111 (N_15111,N_13899,N_14167);
or U15112 (N_15112,N_14815,N_14860);
or U15113 (N_15113,N_13594,N_14737);
nand U15114 (N_15114,N_14279,N_13531);
or U15115 (N_15115,N_13655,N_13502);
nor U15116 (N_15116,N_13621,N_14690);
xor U15117 (N_15117,N_14541,N_14062);
xnor U15118 (N_15118,N_14654,N_14741);
xor U15119 (N_15119,N_13708,N_14407);
and U15120 (N_15120,N_14245,N_14175);
and U15121 (N_15121,N_14781,N_14444);
and U15122 (N_15122,N_13680,N_14770);
xor U15123 (N_15123,N_13659,N_14488);
xnor U15124 (N_15124,N_14092,N_14393);
and U15125 (N_15125,N_14350,N_14557);
and U15126 (N_15126,N_14963,N_14573);
or U15127 (N_15127,N_14739,N_13980);
and U15128 (N_15128,N_14139,N_14449);
nand U15129 (N_15129,N_14191,N_13511);
and U15130 (N_15130,N_14081,N_14007);
and U15131 (N_15131,N_13741,N_13926);
nand U15132 (N_15132,N_14097,N_14272);
nand U15133 (N_15133,N_14661,N_14163);
nor U15134 (N_15134,N_13719,N_13744);
xnor U15135 (N_15135,N_13617,N_13891);
or U15136 (N_15136,N_14910,N_14754);
nor U15137 (N_15137,N_14108,N_14774);
xor U15138 (N_15138,N_13545,N_14938);
nor U15139 (N_15139,N_13764,N_13732);
nor U15140 (N_15140,N_14459,N_14258);
nand U15141 (N_15141,N_14618,N_13533);
and U15142 (N_15142,N_13657,N_14147);
or U15143 (N_15143,N_14440,N_14707);
or U15144 (N_15144,N_14494,N_14231);
xnor U15145 (N_15145,N_14670,N_14060);
nand U15146 (N_15146,N_13909,N_14713);
nand U15147 (N_15147,N_13735,N_14634);
or U15148 (N_15148,N_14587,N_14964);
nor U15149 (N_15149,N_14410,N_14464);
nor U15150 (N_15150,N_13566,N_14717);
nor U15151 (N_15151,N_13703,N_13989);
nor U15152 (N_15152,N_14819,N_14046);
nor U15153 (N_15153,N_13915,N_14349);
or U15154 (N_15154,N_14390,N_13943);
xnor U15155 (N_15155,N_14057,N_14009);
or U15156 (N_15156,N_14508,N_14428);
xnor U15157 (N_15157,N_14679,N_14480);
nor U15158 (N_15158,N_14752,N_14897);
nor U15159 (N_15159,N_14313,N_14955);
or U15160 (N_15160,N_14264,N_14273);
nand U15161 (N_15161,N_14100,N_13832);
nor U15162 (N_15162,N_14458,N_13609);
nand U15163 (N_15163,N_13731,N_13738);
nand U15164 (N_15164,N_14960,N_14165);
nor U15165 (N_15165,N_14413,N_13789);
xnor U15166 (N_15166,N_14262,N_14048);
and U15167 (N_15167,N_14820,N_14021);
nor U15168 (N_15168,N_14331,N_14355);
nand U15169 (N_15169,N_14732,N_14686);
or U15170 (N_15170,N_14423,N_14514);
xnor U15171 (N_15171,N_14320,N_13560);
and U15172 (N_15172,N_13624,N_14600);
nor U15173 (N_15173,N_14968,N_14611);
xor U15174 (N_15174,N_14560,N_13647);
or U15175 (N_15175,N_14594,N_14522);
and U15176 (N_15176,N_14850,N_13702);
and U15177 (N_15177,N_14913,N_14341);
or U15178 (N_15178,N_14025,N_13711);
nor U15179 (N_15179,N_14063,N_14244);
or U15180 (N_15180,N_13852,N_14246);
and U15181 (N_15181,N_13562,N_14019);
nand U15182 (N_15182,N_14721,N_13693);
nand U15183 (N_15183,N_14497,N_13953);
nor U15184 (N_15184,N_14760,N_14376);
nand U15185 (N_15185,N_14075,N_14076);
or U15186 (N_15186,N_14363,N_13998);
nand U15187 (N_15187,N_13974,N_14116);
xnor U15188 (N_15188,N_14134,N_13936);
nand U15189 (N_15189,N_14209,N_14787);
and U15190 (N_15190,N_14866,N_13635);
nand U15191 (N_15191,N_14746,N_14419);
nor U15192 (N_15192,N_14603,N_14000);
nor U15193 (N_15193,N_14879,N_13973);
nand U15194 (N_15194,N_13922,N_13835);
nand U15195 (N_15195,N_14012,N_13889);
and U15196 (N_15196,N_14130,N_14750);
nand U15197 (N_15197,N_13767,N_14270);
nand U15198 (N_15198,N_13640,N_14588);
or U15199 (N_15199,N_14304,N_14796);
nand U15200 (N_15200,N_13765,N_13572);
nor U15201 (N_15201,N_14817,N_13940);
xnor U15202 (N_15202,N_13892,N_14676);
nand U15203 (N_15203,N_13987,N_14539);
nand U15204 (N_15204,N_14799,N_13623);
and U15205 (N_15205,N_13721,N_13933);
xnor U15206 (N_15206,N_14682,N_13966);
xor U15207 (N_15207,N_13638,N_13965);
and U15208 (N_15208,N_13904,N_13868);
and U15209 (N_15209,N_14132,N_13941);
or U15210 (N_15210,N_13642,N_14305);
and U15211 (N_15211,N_14237,N_14748);
or U15212 (N_15212,N_14793,N_13781);
or U15213 (N_15213,N_14547,N_14852);
and U15214 (N_15214,N_14096,N_14113);
nand U15215 (N_15215,N_14026,N_14899);
nor U15216 (N_15216,N_13684,N_14751);
or U15217 (N_15217,N_14267,N_13976);
nor U15218 (N_15218,N_14283,N_14486);
or U15219 (N_15219,N_13924,N_14103);
nor U15220 (N_15220,N_14633,N_14749);
or U15221 (N_15221,N_13903,N_14889);
nand U15222 (N_15222,N_13887,N_14360);
or U15223 (N_15223,N_14698,N_14215);
or U15224 (N_15224,N_13616,N_13627);
or U15225 (N_15225,N_13580,N_14589);
and U15226 (N_15226,N_14037,N_13612);
xnor U15227 (N_15227,N_14550,N_13994);
xnor U15228 (N_15228,N_13804,N_14932);
or U15229 (N_15229,N_13710,N_14439);
nand U15230 (N_15230,N_13768,N_14705);
xnor U15231 (N_15231,N_13917,N_14450);
or U15232 (N_15232,N_13871,N_14252);
nand U15233 (N_15233,N_14263,N_13720);
and U15234 (N_15234,N_13920,N_14545);
and U15235 (N_15235,N_13602,N_13688);
nand U15236 (N_15236,N_13923,N_13587);
nor U15237 (N_15237,N_14085,N_14447);
xnor U15238 (N_15238,N_13896,N_13501);
or U15239 (N_15239,N_14453,N_14632);
nand U15240 (N_15240,N_13664,N_13955);
and U15241 (N_15241,N_13588,N_14659);
and U15242 (N_15242,N_13770,N_14917);
xnor U15243 (N_15243,N_14569,N_14953);
xnor U15244 (N_15244,N_14901,N_14959);
nor U15245 (N_15245,N_14821,N_14402);
nand U15246 (N_15246,N_14500,N_13961);
nor U15247 (N_15247,N_14333,N_13563);
nand U15248 (N_15248,N_14517,N_13773);
xor U15249 (N_15249,N_13524,N_14259);
and U15250 (N_15250,N_14745,N_14672);
nand U15251 (N_15251,N_14675,N_14342);
and U15252 (N_15252,N_14947,N_13860);
nand U15253 (N_15253,N_14987,N_14150);
nor U15254 (N_15254,N_13725,N_13849);
xnor U15255 (N_15255,N_14105,N_14271);
or U15256 (N_15256,N_14161,N_13788);
and U15257 (N_15257,N_14747,N_14039);
xor U15258 (N_15258,N_14591,N_13542);
or U15259 (N_15259,N_14095,N_14394);
nor U15260 (N_15260,N_14544,N_14996);
or U15261 (N_15261,N_13779,N_13536);
xor U15262 (N_15262,N_14802,N_14087);
nand U15263 (N_15263,N_13870,N_14074);
nor U15264 (N_15264,N_14697,N_13983);
nand U15265 (N_15265,N_14624,N_13661);
or U15266 (N_15266,N_14316,N_14422);
xnor U15267 (N_15267,N_14709,N_14561);
nor U15268 (N_15268,N_13798,N_14991);
and U15269 (N_15269,N_13592,N_14335);
or U15270 (N_15270,N_14609,N_14548);
nand U15271 (N_15271,N_14767,N_13866);
nor U15272 (N_15272,N_14432,N_13705);
xnor U15273 (N_15273,N_14753,N_14640);
and U15274 (N_15274,N_14036,N_13707);
xnor U15275 (N_15275,N_13730,N_13570);
xnor U15276 (N_15276,N_14563,N_14602);
xor U15277 (N_15277,N_13811,N_14873);
nor U15278 (N_15278,N_13668,N_14274);
nor U15279 (N_15279,N_14814,N_14553);
nand U15280 (N_15280,N_14367,N_14689);
nand U15281 (N_15281,N_14182,N_14663);
nor U15282 (N_15282,N_14776,N_13857);
and U15283 (N_15283,N_14838,N_14711);
and U15284 (N_15284,N_14140,N_13982);
and U15285 (N_15285,N_14442,N_13823);
xnor U15286 (N_15286,N_14015,N_14729);
and U15287 (N_15287,N_14373,N_13593);
and U15288 (N_15288,N_14979,N_14171);
xnor U15289 (N_15289,N_13611,N_14612);
or U15290 (N_15290,N_14181,N_14371);
and U15291 (N_15291,N_14099,N_14948);
xnor U15292 (N_15292,N_13816,N_13669);
nor U15293 (N_15293,N_14114,N_13752);
and U15294 (N_15294,N_13598,N_13706);
and U15295 (N_15295,N_13520,N_14798);
and U15296 (N_15296,N_13747,N_14683);
or U15297 (N_15297,N_14178,N_14388);
or U15298 (N_15298,N_13508,N_14934);
or U15299 (N_15299,N_13977,N_14554);
and U15300 (N_15300,N_14861,N_13506);
or U15301 (N_15301,N_13934,N_14180);
xor U15302 (N_15302,N_14941,N_13797);
nand U15303 (N_15303,N_14980,N_14196);
and U15304 (N_15304,N_14915,N_14041);
xnor U15305 (N_15305,N_14348,N_13628);
or U15306 (N_15306,N_14011,N_14002);
xor U15307 (N_15307,N_13644,N_14647);
nor U15308 (N_15308,N_14863,N_14865);
or U15309 (N_15309,N_14020,N_14975);
or U15310 (N_15310,N_14605,N_14368);
or U15311 (N_15311,N_14149,N_13761);
nor U15312 (N_15312,N_14571,N_14726);
nor U15313 (N_15313,N_14230,N_13890);
nand U15314 (N_15314,N_13574,N_14253);
nand U15315 (N_15315,N_14216,N_14702);
and U15316 (N_15316,N_14894,N_14535);
nor U15317 (N_15317,N_14907,N_14013);
xnor U15318 (N_15318,N_14608,N_13846);
and U15319 (N_15319,N_14387,N_13620);
or U15320 (N_15320,N_13911,N_14905);
nand U15321 (N_15321,N_14408,N_14038);
xor U15322 (N_15322,N_14766,N_14834);
nand U15323 (N_15323,N_14623,N_14718);
or U15324 (N_15324,N_13589,N_14001);
nand U15325 (N_15325,N_14277,N_14939);
or U15326 (N_15326,N_14050,N_14556);
xnor U15327 (N_15327,N_14275,N_13999);
nand U15328 (N_15328,N_13753,N_14878);
nor U15329 (N_15329,N_14703,N_14478);
or U15330 (N_15330,N_14033,N_14667);
nand U15331 (N_15331,N_14540,N_14645);
xnor U15332 (N_15332,N_14551,N_13838);
xor U15333 (N_15333,N_13762,N_14925);
nor U15334 (N_15334,N_13746,N_13658);
or U15335 (N_15335,N_14764,N_14736);
and U15336 (N_15336,N_14565,N_14839);
xnor U15337 (N_15337,N_13854,N_14918);
xor U15338 (N_15338,N_14847,N_14825);
xor U15339 (N_15339,N_13869,N_14791);
and U15340 (N_15340,N_14778,N_13807);
xor U15341 (N_15341,N_13990,N_14681);
nand U15342 (N_15342,N_14286,N_14827);
or U15343 (N_15343,N_14503,N_14164);
or U15344 (N_15344,N_14687,N_13600);
or U15345 (N_15345,N_13806,N_14281);
xor U15346 (N_15346,N_14421,N_14531);
nor U15347 (N_15347,N_13697,N_13931);
or U15348 (N_15348,N_14117,N_14538);
nor U15349 (N_15349,N_14769,N_14261);
nor U15350 (N_15350,N_13576,N_13984);
xor U15351 (N_15351,N_13581,N_14239);
and U15352 (N_15352,N_13956,N_14330);
and U15353 (N_15353,N_13686,N_14044);
nand U15354 (N_15354,N_13660,N_14314);
xnor U15355 (N_15355,N_14416,N_14989);
and U15356 (N_15356,N_14622,N_13613);
xnor U15357 (N_15357,N_14877,N_14203);
nand U15358 (N_15358,N_14701,N_13584);
nand U15359 (N_15359,N_14971,N_14386);
nor U15360 (N_15360,N_13694,N_13713);
or U15361 (N_15361,N_13803,N_14625);
and U15362 (N_15362,N_13504,N_14582);
nor U15363 (N_15363,N_13583,N_13775);
or U15364 (N_15364,N_14080,N_14528);
and U15365 (N_15365,N_13527,N_13736);
and U15366 (N_15366,N_13897,N_14641);
and U15367 (N_15367,N_14496,N_14974);
nor U15368 (N_15368,N_14326,N_14091);
nor U15369 (N_15369,N_13618,N_14200);
xnor U15370 (N_15370,N_13512,N_14122);
nand U15371 (N_15371,N_14437,N_14518);
nor U15372 (N_15372,N_13505,N_13601);
xor U15373 (N_15373,N_13678,N_14649);
xor U15374 (N_15374,N_14643,N_14045);
or U15375 (N_15375,N_13554,N_14874);
or U15376 (N_15376,N_13969,N_14016);
nand U15377 (N_15377,N_13681,N_14358);
nor U15378 (N_15378,N_14242,N_13760);
or U15379 (N_15379,N_13754,N_14700);
nor U15380 (N_15380,N_14476,N_14443);
and U15381 (N_15381,N_14024,N_14429);
xnor U15382 (N_15382,N_14481,N_13547);
nand U15383 (N_15383,N_14699,N_13571);
and U15384 (N_15384,N_14395,N_13701);
or U15385 (N_15385,N_13573,N_14332);
nand U15386 (N_15386,N_13817,N_14483);
or U15387 (N_15387,N_14704,N_14456);
or U15388 (N_15388,N_14218,N_14806);
xnor U15389 (N_15389,N_13908,N_14241);
or U15390 (N_15390,N_14288,N_14123);
nand U15391 (N_15391,N_14303,N_14797);
nor U15392 (N_15392,N_14593,N_14465);
xnor U15393 (N_15393,N_14301,N_14498);
or U15394 (N_15394,N_14638,N_14990);
or U15395 (N_15395,N_14257,N_14680);
xnor U15396 (N_15396,N_14131,N_14035);
and U15397 (N_15397,N_14477,N_14366);
xnor U15398 (N_15398,N_13971,N_14864);
or U15399 (N_15399,N_14153,N_13959);
xnor U15400 (N_15400,N_14543,N_14484);
nor U15401 (N_15401,N_13847,N_14415);
xnor U15402 (N_15402,N_14022,N_13772);
xnor U15403 (N_15403,N_14457,N_14994);
xor U15404 (N_15404,N_13787,N_14929);
xor U15405 (N_15405,N_13546,N_13629);
nor U15406 (N_15406,N_14454,N_14856);
nand U15407 (N_15407,N_14762,N_14969);
nor U15408 (N_15408,N_13991,N_14723);
nand U15409 (N_15409,N_14006,N_14004);
or U15410 (N_15410,N_14120,N_14937);
xnor U15411 (N_15411,N_14389,N_13586);
nor U15412 (N_15412,N_13539,N_14813);
nor U15413 (N_15413,N_13825,N_14471);
nor U15414 (N_15414,N_14607,N_14743);
and U15415 (N_15415,N_14724,N_14089);
and U15416 (N_15416,N_14206,N_14922);
nor U15417 (N_15417,N_14771,N_14849);
nor U15418 (N_15418,N_14107,N_14409);
xnor U15419 (N_15419,N_13698,N_14344);
nor U15420 (N_15420,N_13535,N_13510);
nand U15421 (N_15421,N_14693,N_13986);
xor U15422 (N_15422,N_14224,N_14197);
xor U15423 (N_15423,N_13837,N_14521);
nand U15424 (N_15424,N_14052,N_13873);
nand U15425 (N_15425,N_14617,N_14930);
nor U15426 (N_15426,N_13848,N_14158);
nor U15427 (N_15427,N_13925,N_13597);
or U15428 (N_15428,N_13756,N_13791);
xnor U15429 (N_15429,N_14810,N_14405);
nor U15430 (N_15430,N_14053,N_13541);
xnor U15431 (N_15431,N_13591,N_14927);
nand U15432 (N_15432,N_13810,N_14294);
and U15433 (N_15433,N_13895,N_14805);
and U15434 (N_15434,N_14157,N_14179);
nor U15435 (N_15435,N_14490,N_14942);
nor U15436 (N_15436,N_13822,N_13932);
and U15437 (N_15437,N_14308,N_14887);
and U15438 (N_15438,N_14302,N_13673);
and U15439 (N_15439,N_14276,N_14660);
nand U15440 (N_15440,N_13718,N_14598);
xnor U15441 (N_15441,N_14055,N_14533);
xnor U15442 (N_15442,N_14297,N_14761);
or U15443 (N_15443,N_14155,N_14223);
nor U15444 (N_15444,N_14674,N_13865);
nand U15445 (N_15445,N_14256,N_14688);
nand U15446 (N_15446,N_14082,N_14614);
or U15447 (N_15447,N_13914,N_14712);
xor U15448 (N_15448,N_14650,N_14102);
nand U15449 (N_15449,N_14347,N_13526);
and U15450 (N_15450,N_14592,N_13614);
nor U15451 (N_15451,N_13958,N_14731);
nor U15452 (N_15452,N_13841,N_13727);
and U15453 (N_15453,N_14900,N_13740);
nor U15454 (N_15454,N_14757,N_14232);
and U15455 (N_15455,N_14706,N_14293);
xor U15456 (N_15456,N_14174,N_14414);
nand U15457 (N_15457,N_14946,N_13518);
nor U15458 (N_15458,N_14364,N_14268);
nor U15459 (N_15459,N_14957,N_13985);
nor U15460 (N_15460,N_14495,N_14967);
nand U15461 (N_15461,N_14311,N_14129);
and U15462 (N_15462,N_14637,N_14187);
xor U15463 (N_15463,N_14287,N_14381);
nor U15464 (N_15464,N_14896,N_14855);
xor U15465 (N_15465,N_13683,N_14162);
nand U15466 (N_15466,N_14727,N_13596);
nand U15467 (N_15467,N_14067,N_13954);
or U15468 (N_15468,N_13665,N_13607);
xor U15469 (N_15469,N_14885,N_14823);
and U15470 (N_15470,N_13928,N_14325);
xor U15471 (N_15471,N_14999,N_14708);
or U15472 (N_15472,N_14474,N_13590);
nand U15473 (N_15473,N_13859,N_14786);
and U15474 (N_15474,N_13840,N_14606);
nor U15475 (N_15475,N_13992,N_14811);
xor U15476 (N_15476,N_14118,N_14578);
nand U15477 (N_15477,N_14775,N_14128);
or U15478 (N_15478,N_14784,N_13595);
nand U15479 (N_15479,N_14613,N_13748);
or U15480 (N_15480,N_14352,N_14417);
nand U15481 (N_15481,N_14205,N_13667);
nand U15482 (N_15482,N_13814,N_14858);
nand U15483 (N_15483,N_13557,N_14221);
xor U15484 (N_15484,N_13757,N_13712);
nor U15485 (N_15485,N_14289,N_14115);
or U15486 (N_15486,N_14362,N_14125);
xor U15487 (N_15487,N_13517,N_14803);
or U15488 (N_15488,N_14652,N_14365);
xnor U15489 (N_15489,N_13567,N_14626);
nor U15490 (N_15490,N_13679,N_13821);
xnor U15491 (N_15491,N_14346,N_13845);
nor U15492 (N_15492,N_14575,N_14840);
nand U15493 (N_15493,N_14620,N_13843);
nand U15494 (N_15494,N_14436,N_14213);
nor U15495 (N_15495,N_14317,N_14936);
nand U15496 (N_15496,N_14523,N_14520);
and U15497 (N_15497,N_14692,N_14119);
and U15498 (N_15498,N_14356,N_13724);
and U15499 (N_15499,N_14435,N_14315);
nor U15500 (N_15500,N_14868,N_14247);
or U15501 (N_15501,N_13842,N_13993);
xor U15502 (N_15502,N_14875,N_14846);
nand U15503 (N_15503,N_14580,N_13970);
and U15504 (N_15504,N_14795,N_14133);
nor U15505 (N_15505,N_14034,N_14061);
and U15506 (N_15506,N_14043,N_13862);
or U15507 (N_15507,N_14260,N_13853);
nor U15508 (N_15508,N_13880,N_13942);
xor U15509 (N_15509,N_14671,N_14426);
and U15510 (N_15510,N_13608,N_13769);
xnor U15511 (N_15511,N_14694,N_14777);
or U15512 (N_15512,N_13950,N_14452);
or U15513 (N_15513,N_14266,N_14944);
nand U15514 (N_15514,N_14378,N_13929);
and U15515 (N_15515,N_14982,N_14604);
or U15516 (N_15516,N_14843,N_13856);
nand U15517 (N_15517,N_14411,N_14420);
and U15518 (N_15518,N_14353,N_14441);
xnor U15519 (N_15519,N_14298,N_14285);
nand U15520 (N_15520,N_13674,N_14728);
and U15521 (N_15521,N_14492,N_13653);
or U15522 (N_15522,N_14678,N_14291);
nor U15523 (N_15523,N_14581,N_14949);
and U15524 (N_15524,N_14501,N_13530);
or U15525 (N_15525,N_13784,N_14832);
or U15526 (N_15526,N_14985,N_14219);
and U15527 (N_15527,N_14662,N_14124);
nor U15528 (N_15528,N_13556,N_13827);
nand U15529 (N_15529,N_14568,N_14920);
and U15530 (N_15530,N_13900,N_14079);
xor U15531 (N_15531,N_14042,N_14370);
nand U15532 (N_15532,N_14127,N_14898);
nand U15533 (N_15533,N_14470,N_14343);
and U15534 (N_15534,N_14385,N_13626);
and U15535 (N_15535,N_14836,N_14822);
or U15536 (N_15536,N_14842,N_14427);
or U15537 (N_15537,N_13569,N_14049);
and U15538 (N_15538,N_14323,N_14135);
or U15539 (N_15539,N_14217,N_14351);
or U15540 (N_15540,N_14380,N_14619);
or U15541 (N_15541,N_13949,N_14715);
and U15542 (N_15542,N_13799,N_14383);
or U15543 (N_15543,N_14401,N_14837);
and U15544 (N_15544,N_13912,N_13631);
and U15545 (N_15545,N_14888,N_13855);
or U15546 (N_15546,N_13516,N_13749);
nand U15547 (N_15547,N_14983,N_13538);
or U15548 (N_15548,N_14467,N_14961);
xor U15549 (N_15549,N_14919,N_14475);
nand U15550 (N_15550,N_14029,N_14526);
nor U15551 (N_15551,N_13715,N_14564);
nor U15552 (N_15552,N_14977,N_13634);
nor U15553 (N_15553,N_14392,N_13918);
or U15554 (N_15554,N_13937,N_14841);
nand U15555 (N_15555,N_13714,N_13826);
nand U15556 (N_15556,N_13881,N_14853);
or U15557 (N_15557,N_13780,N_14199);
and U15558 (N_15558,N_13913,N_14758);
xor U15559 (N_15559,N_13564,N_13555);
nand U15560 (N_15560,N_14871,N_14318);
xor U15561 (N_15561,N_14469,N_14773);
or U15562 (N_15562,N_14644,N_14763);
or U15563 (N_15563,N_14695,N_13919);
nand U15564 (N_15564,N_14986,N_13625);
nor U15565 (N_15565,N_13774,N_14583);
nor U15566 (N_15566,N_14027,N_14278);
or U15567 (N_15567,N_14069,N_14579);
nor U15568 (N_15568,N_14339,N_14211);
or U15569 (N_15569,N_14482,N_13876);
nand U15570 (N_15570,N_14629,N_14642);
or U15571 (N_15571,N_13577,N_14194);
nand U15572 (N_15572,N_13963,N_14321);
nor U15573 (N_15573,N_13619,N_14586);
and U15574 (N_15574,N_14785,N_13975);
nand U15575 (N_15575,N_13641,N_13550);
nor U15576 (N_15576,N_13548,N_13785);
xnor U15577 (N_15577,N_13812,N_14912);
xnor U15578 (N_15578,N_14504,N_14159);
and U15579 (N_15579,N_14870,N_13945);
nor U15580 (N_15580,N_14529,N_13939);
or U15581 (N_15581,N_14978,N_13877);
nand U15582 (N_15582,N_14491,N_14238);
and U15583 (N_15583,N_14993,N_14090);
nor U15584 (N_15584,N_14552,N_13962);
or U15585 (N_15585,N_14472,N_13523);
xor U15586 (N_15586,N_14988,N_14696);
or U15587 (N_15587,N_14646,N_14319);
and U15588 (N_15588,N_13650,N_13763);
nand U15589 (N_15589,N_13700,N_13677);
or U15590 (N_15590,N_14779,N_13813);
nor U15591 (N_15591,N_14269,N_14396);
xor U15592 (N_15592,N_14152,N_14908);
and U15593 (N_15593,N_14883,N_14098);
nand U15594 (N_15594,N_13805,N_14201);
and U15595 (N_15595,N_14666,N_13559);
or U15596 (N_15596,N_14451,N_14923);
or U15597 (N_15597,N_13540,N_13878);
or U15598 (N_15598,N_14950,N_14893);
or U15599 (N_15599,N_14566,N_13979);
and U15600 (N_15600,N_14106,N_13630);
or U15601 (N_15601,N_14083,N_13561);
or U15602 (N_15602,N_14292,N_14906);
or U15603 (N_15603,N_13532,N_14924);
xnor U15604 (N_15604,N_13610,N_13662);
nor U15605 (N_15605,N_14966,N_14904);
nand U15606 (N_15606,N_14809,N_14794);
and U15607 (N_15607,N_14911,N_14824);
nor U15608 (N_15608,N_14615,N_14653);
xor U15609 (N_15609,N_14473,N_14354);
nor U15610 (N_15610,N_13645,N_14322);
nor U15611 (N_15611,N_14808,N_13682);
nor U15612 (N_15612,N_14665,N_14307);
nor U15613 (N_15613,N_13689,N_14059);
and U15614 (N_15614,N_14507,N_14397);
or U15615 (N_15615,N_13685,N_13654);
or U15616 (N_15616,N_13927,N_14058);
nand U15617 (N_15617,N_14008,N_14558);
nor U15618 (N_15618,N_14892,N_13759);
and U15619 (N_15619,N_14438,N_14555);
or U15620 (N_15620,N_13884,N_14361);
nand U15621 (N_15621,N_14337,N_13802);
nand U15622 (N_15622,N_14895,N_13863);
nand U15623 (N_15623,N_14222,N_13894);
xnor U15624 (N_15624,N_14312,N_13722);
nand U15625 (N_15625,N_14848,N_14570);
xnor U15626 (N_15626,N_13778,N_14265);
and U15627 (N_15627,N_14111,N_14462);
xnor U15628 (N_15628,N_14054,N_14005);
or U15629 (N_15629,N_13543,N_14845);
xor U15630 (N_15630,N_13819,N_14229);
xor U15631 (N_15631,N_14940,N_14014);
and U15632 (N_15632,N_14857,N_14630);
or U15633 (N_15633,N_14225,N_14031);
or U15634 (N_15634,N_14828,N_13972);
or U15635 (N_15635,N_14084,N_14768);
xnor U15636 (N_15636,N_13652,N_13967);
or U15637 (N_15637,N_14466,N_14984);
and U15638 (N_15638,N_14493,N_14789);
nor U15639 (N_15639,N_13839,N_14340);
and U15640 (N_15640,N_14170,N_14077);
nor U15641 (N_15641,N_14816,N_13544);
nand U15642 (N_15642,N_14485,N_14299);
nand U15643 (N_15643,N_14765,N_13552);
or U15644 (N_15644,N_14240,N_13758);
xor U15645 (N_15645,N_14788,N_13921);
xor U15646 (N_15646,N_14032,N_13861);
nor U15647 (N_15647,N_13944,N_14862);
nor U15648 (N_15648,N_14735,N_14585);
nand U15649 (N_15649,N_13796,N_14094);
nor U15650 (N_15650,N_13809,N_13742);
nor U15651 (N_15651,N_13885,N_13513);
nor U15652 (N_15652,N_14574,N_14280);
nor U15653 (N_15653,N_14138,N_14512);
nand U15654 (N_15654,N_14844,N_14468);
nor U15655 (N_15655,N_14198,N_14890);
xor U15656 (N_15656,N_14143,N_14998);
nand U15657 (N_15657,N_14954,N_14144);
xnor U15658 (N_15658,N_14234,N_14599);
nor U15659 (N_15659,N_14290,N_14738);
nor U15660 (N_15660,N_14086,N_14066);
and U15661 (N_15661,N_14212,N_14903);
nand U15662 (N_15662,N_14595,N_13604);
nor U15663 (N_15663,N_14169,N_14028);
xnor U15664 (N_15664,N_14040,N_13834);
xnor U15665 (N_15665,N_13675,N_14188);
nor U15666 (N_15666,N_14121,N_14755);
nand U15667 (N_15667,N_13997,N_14530);
and U15668 (N_15668,N_13734,N_14479);
nor U15669 (N_15669,N_14306,N_13519);
and U15670 (N_15670,N_13882,N_14141);
xnor U15671 (N_15671,N_13801,N_14248);
and U15672 (N_15672,N_14902,N_14790);
xnor U15673 (N_15673,N_13615,N_13874);
nand U15674 (N_15674,N_14536,N_14818);
nand U15675 (N_15675,N_14601,N_14730);
or U15676 (N_15676,N_14186,N_13648);
and U15677 (N_15677,N_14101,N_14249);
and U15678 (N_15678,N_13728,N_14412);
or U15679 (N_15679,N_14655,N_14088);
nand U15680 (N_15680,N_14160,N_14176);
and U15681 (N_15681,N_14513,N_14719);
and U15682 (N_15682,N_14406,N_14506);
and U15683 (N_15683,N_13739,N_13509);
or U15684 (N_15684,N_14399,N_13996);
and U15685 (N_15685,N_14714,N_13737);
nand U15686 (N_15686,N_13906,N_14243);
nand U15687 (N_15687,N_13575,N_14636);
and U15688 (N_15688,N_13988,N_14756);
nand U15689 (N_15689,N_13579,N_13528);
nand U15690 (N_15690,N_14047,N_13782);
nand U15691 (N_15691,N_14995,N_14716);
xor U15692 (N_15692,N_14546,N_14359);
and U15693 (N_15693,N_14236,N_13888);
nor U15694 (N_15694,N_14584,N_13968);
and U15695 (N_15695,N_13867,N_13808);
and U15696 (N_15696,N_13633,N_13815);
nand U15697 (N_15697,N_13946,N_14461);
nand U15698 (N_15698,N_14881,N_14382);
or U15699 (N_15699,N_14400,N_14372);
or U15700 (N_15700,N_14071,N_13981);
and U15701 (N_15701,N_14145,N_13666);
and U15702 (N_15702,N_14156,N_13717);
or U15703 (N_15703,N_13726,N_14345);
nand U15704 (N_15704,N_13585,N_13709);
or U15705 (N_15705,N_14109,N_14334);
or U15706 (N_15706,N_14559,N_14056);
nand U15707 (N_15707,N_13578,N_14933);
nand U15708 (N_15708,N_14952,N_14826);
nand U15709 (N_15709,N_13751,N_14973);
xnor U15710 (N_15710,N_14391,N_13534);
xor U15711 (N_15711,N_14882,N_14374);
or U15712 (N_15712,N_14010,N_13605);
xnor U15713 (N_15713,N_14829,N_13663);
and U15714 (N_15714,N_14742,N_13723);
xor U15715 (N_15715,N_14148,N_14951);
nor U15716 (N_15716,N_14833,N_14284);
xor U15717 (N_15717,N_14166,N_14434);
nor U15718 (N_15718,N_14891,N_13836);
nor U15719 (N_15719,N_13750,N_13951);
nand U15720 (N_15720,N_14184,N_13651);
xnor U15721 (N_15721,N_13776,N_14505);
or U15722 (N_15722,N_13851,N_14136);
and U15723 (N_15723,N_13646,N_14962);
or U15724 (N_15724,N_13755,N_14651);
nand U15725 (N_15725,N_14807,N_14210);
and U15726 (N_15726,N_14172,N_14872);
nor U15727 (N_15727,N_14734,N_13830);
nor U15728 (N_15728,N_13883,N_14886);
or U15729 (N_15729,N_14648,N_13960);
and U15730 (N_15730,N_14830,N_14516);
nor U15731 (N_15731,N_14800,N_14519);
nor U15732 (N_15732,N_13795,N_13938);
xnor U15733 (N_15733,N_14722,N_14489);
nor U15734 (N_15734,N_14403,N_14869);
and U15735 (N_15735,N_14965,N_13898);
nand U15736 (N_15736,N_14884,N_14958);
or U15737 (N_15737,N_14976,N_14110);
nand U15738 (N_15738,N_14549,N_13901);
and U15739 (N_15739,N_13549,N_14068);
or U15740 (N_15740,N_14525,N_14772);
and U15741 (N_15741,N_14448,N_14051);
xnor U15742 (N_15742,N_14336,N_13930);
and U15743 (N_15743,N_14997,N_13743);
nand U15744 (N_15744,N_13829,N_14250);
nor U15745 (N_15745,N_13995,N_14657);
nor U15746 (N_15746,N_14173,N_14744);
and U15747 (N_15747,N_14499,N_14542);
xnor U15748 (N_15748,N_14509,N_14628);
nand U15749 (N_15749,N_14190,N_13670);
nand U15750 (N_15750,N_14741,N_14310);
nor U15751 (N_15751,N_14082,N_13580);
and U15752 (N_15752,N_14946,N_14287);
nor U15753 (N_15753,N_14287,N_14197);
nand U15754 (N_15754,N_14000,N_14326);
and U15755 (N_15755,N_13745,N_14991);
xnor U15756 (N_15756,N_14688,N_14372);
xor U15757 (N_15757,N_14373,N_14134);
nor U15758 (N_15758,N_13511,N_14755);
nor U15759 (N_15759,N_13936,N_14017);
nand U15760 (N_15760,N_14633,N_14690);
or U15761 (N_15761,N_14433,N_14732);
or U15762 (N_15762,N_14225,N_13645);
nor U15763 (N_15763,N_13907,N_14291);
nor U15764 (N_15764,N_14642,N_13957);
or U15765 (N_15765,N_13736,N_14616);
nor U15766 (N_15766,N_14922,N_14992);
or U15767 (N_15767,N_14034,N_13753);
nand U15768 (N_15768,N_14790,N_14820);
and U15769 (N_15769,N_14271,N_14112);
nand U15770 (N_15770,N_13996,N_13627);
or U15771 (N_15771,N_14966,N_14122);
xor U15772 (N_15772,N_14937,N_14197);
xor U15773 (N_15773,N_14878,N_14110);
xor U15774 (N_15774,N_14380,N_13703);
and U15775 (N_15775,N_14878,N_14151);
xnor U15776 (N_15776,N_13833,N_14953);
and U15777 (N_15777,N_13937,N_14523);
and U15778 (N_15778,N_13729,N_14756);
nand U15779 (N_15779,N_14232,N_14611);
nand U15780 (N_15780,N_13844,N_14878);
nor U15781 (N_15781,N_13944,N_13862);
xor U15782 (N_15782,N_14667,N_13977);
and U15783 (N_15783,N_14962,N_14367);
or U15784 (N_15784,N_13505,N_13949);
nand U15785 (N_15785,N_13867,N_13951);
xor U15786 (N_15786,N_13837,N_14478);
nand U15787 (N_15787,N_14027,N_14133);
or U15788 (N_15788,N_14580,N_13689);
or U15789 (N_15789,N_13536,N_14558);
and U15790 (N_15790,N_13623,N_13909);
nand U15791 (N_15791,N_13755,N_14082);
xor U15792 (N_15792,N_14055,N_14375);
and U15793 (N_15793,N_14107,N_14057);
and U15794 (N_15794,N_14670,N_14431);
xnor U15795 (N_15795,N_14304,N_14802);
xnor U15796 (N_15796,N_14698,N_14562);
xnor U15797 (N_15797,N_13972,N_14906);
nor U15798 (N_15798,N_14515,N_14543);
xor U15799 (N_15799,N_14654,N_14635);
xnor U15800 (N_15800,N_14407,N_13541);
nor U15801 (N_15801,N_13917,N_14864);
or U15802 (N_15802,N_14261,N_13730);
xor U15803 (N_15803,N_14371,N_14446);
and U15804 (N_15804,N_14908,N_13668);
nand U15805 (N_15805,N_14567,N_14504);
or U15806 (N_15806,N_14011,N_13745);
nand U15807 (N_15807,N_13662,N_13905);
or U15808 (N_15808,N_14931,N_14659);
and U15809 (N_15809,N_14243,N_14112);
nor U15810 (N_15810,N_13760,N_14618);
nand U15811 (N_15811,N_14494,N_14751);
xnor U15812 (N_15812,N_14717,N_14314);
nand U15813 (N_15813,N_14543,N_14224);
nor U15814 (N_15814,N_13691,N_14794);
nor U15815 (N_15815,N_14525,N_14408);
or U15816 (N_15816,N_14835,N_14357);
nand U15817 (N_15817,N_13545,N_13541);
xnor U15818 (N_15818,N_14138,N_14236);
or U15819 (N_15819,N_14496,N_14426);
and U15820 (N_15820,N_14368,N_14656);
or U15821 (N_15821,N_14130,N_14731);
or U15822 (N_15822,N_14562,N_13921);
xnor U15823 (N_15823,N_14575,N_13798);
or U15824 (N_15824,N_14382,N_14742);
and U15825 (N_15825,N_14447,N_14828);
xor U15826 (N_15826,N_14698,N_13726);
or U15827 (N_15827,N_13627,N_13949);
xor U15828 (N_15828,N_14380,N_14127);
and U15829 (N_15829,N_14304,N_14878);
or U15830 (N_15830,N_14876,N_13711);
nor U15831 (N_15831,N_13888,N_14184);
or U15832 (N_15832,N_13506,N_14787);
or U15833 (N_15833,N_14874,N_13871);
or U15834 (N_15834,N_14457,N_13951);
xor U15835 (N_15835,N_14720,N_13529);
and U15836 (N_15836,N_14892,N_14227);
or U15837 (N_15837,N_14110,N_13718);
xnor U15838 (N_15838,N_13682,N_13592);
nand U15839 (N_15839,N_14774,N_13650);
and U15840 (N_15840,N_14368,N_14703);
and U15841 (N_15841,N_13586,N_13920);
nand U15842 (N_15842,N_14615,N_14924);
or U15843 (N_15843,N_13780,N_14464);
xnor U15844 (N_15844,N_14288,N_13994);
or U15845 (N_15845,N_14375,N_13571);
nand U15846 (N_15846,N_14538,N_14136);
nor U15847 (N_15847,N_13560,N_14515);
nor U15848 (N_15848,N_14111,N_14278);
nor U15849 (N_15849,N_13722,N_13647);
nor U15850 (N_15850,N_14081,N_14805);
or U15851 (N_15851,N_14504,N_14221);
nor U15852 (N_15852,N_14872,N_13909);
and U15853 (N_15853,N_13979,N_14385);
nand U15854 (N_15854,N_14788,N_13754);
xnor U15855 (N_15855,N_14826,N_13566);
or U15856 (N_15856,N_13912,N_13757);
nor U15857 (N_15857,N_14516,N_14845);
or U15858 (N_15858,N_14781,N_13648);
and U15859 (N_15859,N_14878,N_14828);
xnor U15860 (N_15860,N_14346,N_14748);
or U15861 (N_15861,N_14918,N_14678);
and U15862 (N_15862,N_14210,N_13629);
nand U15863 (N_15863,N_13738,N_14512);
nor U15864 (N_15864,N_14395,N_14224);
nand U15865 (N_15865,N_14621,N_13965);
nor U15866 (N_15866,N_14071,N_14894);
xnor U15867 (N_15867,N_13605,N_14507);
xnor U15868 (N_15868,N_14394,N_14018);
xor U15869 (N_15869,N_14466,N_13836);
xnor U15870 (N_15870,N_14306,N_14246);
nor U15871 (N_15871,N_14118,N_13691);
or U15872 (N_15872,N_13637,N_14266);
nor U15873 (N_15873,N_13519,N_14048);
or U15874 (N_15874,N_14633,N_13652);
and U15875 (N_15875,N_14719,N_13859);
and U15876 (N_15876,N_13714,N_14044);
xor U15877 (N_15877,N_14216,N_14877);
nand U15878 (N_15878,N_14298,N_14244);
or U15879 (N_15879,N_13500,N_13728);
xnor U15880 (N_15880,N_14503,N_14862);
or U15881 (N_15881,N_14166,N_13814);
and U15882 (N_15882,N_14884,N_13917);
or U15883 (N_15883,N_14155,N_14535);
or U15884 (N_15884,N_14112,N_14183);
nor U15885 (N_15885,N_14188,N_13838);
nor U15886 (N_15886,N_14076,N_13530);
nand U15887 (N_15887,N_14141,N_14301);
and U15888 (N_15888,N_13788,N_14664);
nor U15889 (N_15889,N_14333,N_14803);
xor U15890 (N_15890,N_14416,N_14295);
and U15891 (N_15891,N_13613,N_14613);
or U15892 (N_15892,N_13915,N_13576);
and U15893 (N_15893,N_14162,N_14599);
or U15894 (N_15894,N_14322,N_13795);
nor U15895 (N_15895,N_13753,N_13934);
xor U15896 (N_15896,N_13858,N_13704);
nor U15897 (N_15897,N_14554,N_13575);
nor U15898 (N_15898,N_14626,N_14422);
nor U15899 (N_15899,N_14545,N_14750);
or U15900 (N_15900,N_13827,N_14685);
nor U15901 (N_15901,N_13728,N_14923);
nor U15902 (N_15902,N_14240,N_14753);
xnor U15903 (N_15903,N_14867,N_14224);
or U15904 (N_15904,N_14991,N_13863);
nor U15905 (N_15905,N_14932,N_14576);
xnor U15906 (N_15906,N_14583,N_13601);
nand U15907 (N_15907,N_14854,N_14699);
nand U15908 (N_15908,N_14638,N_14838);
nor U15909 (N_15909,N_14208,N_14822);
or U15910 (N_15910,N_14585,N_13697);
nand U15911 (N_15911,N_14377,N_14474);
xor U15912 (N_15912,N_13869,N_13837);
nor U15913 (N_15913,N_14852,N_13526);
xor U15914 (N_15914,N_14166,N_13630);
or U15915 (N_15915,N_14610,N_14673);
or U15916 (N_15916,N_14673,N_14213);
xnor U15917 (N_15917,N_14268,N_14536);
and U15918 (N_15918,N_13701,N_14689);
xor U15919 (N_15919,N_14282,N_13566);
xor U15920 (N_15920,N_14206,N_14066);
xor U15921 (N_15921,N_14427,N_13631);
nand U15922 (N_15922,N_14558,N_14154);
nand U15923 (N_15923,N_14712,N_14518);
and U15924 (N_15924,N_14088,N_13513);
xor U15925 (N_15925,N_13930,N_14725);
nor U15926 (N_15926,N_14663,N_13802);
nand U15927 (N_15927,N_13733,N_14875);
xor U15928 (N_15928,N_13611,N_13787);
or U15929 (N_15929,N_14375,N_14827);
nand U15930 (N_15930,N_14650,N_14396);
nand U15931 (N_15931,N_14003,N_14867);
nand U15932 (N_15932,N_13591,N_14039);
nor U15933 (N_15933,N_13626,N_13971);
or U15934 (N_15934,N_13647,N_13892);
nor U15935 (N_15935,N_14612,N_14872);
nand U15936 (N_15936,N_13890,N_14519);
xnor U15937 (N_15937,N_13711,N_14205);
xnor U15938 (N_15938,N_13853,N_14485);
or U15939 (N_15939,N_13960,N_14566);
or U15940 (N_15940,N_13506,N_14469);
and U15941 (N_15941,N_14109,N_14761);
nor U15942 (N_15942,N_14400,N_13855);
and U15943 (N_15943,N_13851,N_13587);
and U15944 (N_15944,N_14484,N_14356);
nor U15945 (N_15945,N_14999,N_14409);
or U15946 (N_15946,N_14618,N_14311);
nand U15947 (N_15947,N_14151,N_14270);
nand U15948 (N_15948,N_14595,N_14150);
xor U15949 (N_15949,N_13792,N_13538);
nand U15950 (N_15950,N_14923,N_14253);
or U15951 (N_15951,N_14116,N_14078);
or U15952 (N_15952,N_14155,N_14618);
nor U15953 (N_15953,N_14160,N_14376);
xnor U15954 (N_15954,N_14453,N_14222);
nand U15955 (N_15955,N_14322,N_14667);
xor U15956 (N_15956,N_13864,N_13921);
and U15957 (N_15957,N_13832,N_14466);
nor U15958 (N_15958,N_13565,N_14011);
or U15959 (N_15959,N_14456,N_13974);
nor U15960 (N_15960,N_14951,N_14124);
nor U15961 (N_15961,N_13650,N_14028);
nand U15962 (N_15962,N_14953,N_14540);
xor U15963 (N_15963,N_14500,N_14472);
nand U15964 (N_15964,N_14518,N_13647);
nor U15965 (N_15965,N_14349,N_14047);
xnor U15966 (N_15966,N_14127,N_14110);
xor U15967 (N_15967,N_13711,N_14339);
nand U15968 (N_15968,N_14558,N_13863);
nand U15969 (N_15969,N_14780,N_13501);
nor U15970 (N_15970,N_14362,N_14314);
xnor U15971 (N_15971,N_14246,N_14774);
and U15972 (N_15972,N_14471,N_14515);
or U15973 (N_15973,N_14319,N_14752);
nor U15974 (N_15974,N_13845,N_14977);
nand U15975 (N_15975,N_13958,N_13796);
and U15976 (N_15976,N_14924,N_14089);
and U15977 (N_15977,N_13845,N_14778);
xor U15978 (N_15978,N_13910,N_14141);
or U15979 (N_15979,N_14333,N_14337);
xnor U15980 (N_15980,N_14151,N_13751);
or U15981 (N_15981,N_13803,N_14938);
nand U15982 (N_15982,N_13903,N_13879);
or U15983 (N_15983,N_14483,N_14755);
nor U15984 (N_15984,N_14344,N_14321);
nand U15985 (N_15985,N_13509,N_14281);
nand U15986 (N_15986,N_14290,N_14314);
or U15987 (N_15987,N_14990,N_14932);
or U15988 (N_15988,N_14452,N_14006);
and U15989 (N_15989,N_14681,N_14888);
xnor U15990 (N_15990,N_13707,N_13860);
or U15991 (N_15991,N_14779,N_14720);
nand U15992 (N_15992,N_14456,N_14506);
and U15993 (N_15993,N_14124,N_13810);
and U15994 (N_15994,N_14932,N_14505);
nor U15995 (N_15995,N_13973,N_14558);
and U15996 (N_15996,N_13743,N_14991);
xnor U15997 (N_15997,N_13723,N_14992);
xnor U15998 (N_15998,N_14854,N_14520);
and U15999 (N_15999,N_14032,N_13540);
or U16000 (N_16000,N_14310,N_14280);
nor U16001 (N_16001,N_14856,N_13763);
or U16002 (N_16002,N_13833,N_14479);
nor U16003 (N_16003,N_13756,N_14887);
xor U16004 (N_16004,N_13549,N_13713);
and U16005 (N_16005,N_13840,N_14565);
and U16006 (N_16006,N_14164,N_14993);
or U16007 (N_16007,N_14669,N_14015);
nor U16008 (N_16008,N_14562,N_13543);
nand U16009 (N_16009,N_13741,N_13589);
or U16010 (N_16010,N_14623,N_14802);
xnor U16011 (N_16011,N_14894,N_13798);
xor U16012 (N_16012,N_13600,N_14127);
and U16013 (N_16013,N_14562,N_14308);
nand U16014 (N_16014,N_14495,N_14522);
xnor U16015 (N_16015,N_14253,N_14863);
and U16016 (N_16016,N_14818,N_13667);
nand U16017 (N_16017,N_13766,N_14086);
xor U16018 (N_16018,N_14167,N_14363);
or U16019 (N_16019,N_14004,N_14164);
nand U16020 (N_16020,N_14801,N_13550);
or U16021 (N_16021,N_14007,N_14114);
xnor U16022 (N_16022,N_14593,N_14162);
xnor U16023 (N_16023,N_14982,N_13552);
or U16024 (N_16024,N_13580,N_14173);
nor U16025 (N_16025,N_13584,N_13589);
or U16026 (N_16026,N_14838,N_13670);
nand U16027 (N_16027,N_13611,N_13932);
nand U16028 (N_16028,N_14976,N_13801);
and U16029 (N_16029,N_13519,N_13507);
nor U16030 (N_16030,N_13822,N_14387);
nand U16031 (N_16031,N_14348,N_14106);
nand U16032 (N_16032,N_14668,N_14488);
and U16033 (N_16033,N_13720,N_13523);
nand U16034 (N_16034,N_13709,N_14428);
or U16035 (N_16035,N_14762,N_14796);
xor U16036 (N_16036,N_13549,N_13760);
and U16037 (N_16037,N_14789,N_13509);
and U16038 (N_16038,N_14239,N_14540);
nand U16039 (N_16039,N_14801,N_14911);
nor U16040 (N_16040,N_14922,N_14439);
nand U16041 (N_16041,N_14880,N_14293);
xnor U16042 (N_16042,N_14199,N_13810);
nand U16043 (N_16043,N_13804,N_14087);
nand U16044 (N_16044,N_13996,N_14375);
or U16045 (N_16045,N_14564,N_14391);
nor U16046 (N_16046,N_13853,N_14635);
nor U16047 (N_16047,N_14591,N_14732);
nand U16048 (N_16048,N_13692,N_13652);
and U16049 (N_16049,N_13523,N_14957);
and U16050 (N_16050,N_14852,N_14787);
or U16051 (N_16051,N_14481,N_13967);
or U16052 (N_16052,N_14336,N_14113);
nand U16053 (N_16053,N_13982,N_14231);
xnor U16054 (N_16054,N_13705,N_14540);
nor U16055 (N_16055,N_14351,N_14405);
and U16056 (N_16056,N_14390,N_14469);
and U16057 (N_16057,N_14400,N_13931);
nand U16058 (N_16058,N_14887,N_14080);
nand U16059 (N_16059,N_14757,N_13559);
and U16060 (N_16060,N_13993,N_13886);
xor U16061 (N_16061,N_13532,N_14541);
nand U16062 (N_16062,N_14702,N_14445);
or U16063 (N_16063,N_14068,N_14351);
and U16064 (N_16064,N_14694,N_14607);
nor U16065 (N_16065,N_14397,N_13669);
and U16066 (N_16066,N_13564,N_14755);
and U16067 (N_16067,N_14318,N_14800);
nor U16068 (N_16068,N_13645,N_13910);
xor U16069 (N_16069,N_13895,N_13556);
nor U16070 (N_16070,N_14428,N_14431);
and U16071 (N_16071,N_13663,N_14165);
or U16072 (N_16072,N_13794,N_14038);
xnor U16073 (N_16073,N_14982,N_14581);
nand U16074 (N_16074,N_14200,N_14447);
and U16075 (N_16075,N_14586,N_14603);
or U16076 (N_16076,N_13598,N_13618);
xnor U16077 (N_16077,N_14252,N_14995);
nand U16078 (N_16078,N_14876,N_14499);
and U16079 (N_16079,N_14673,N_14582);
xor U16080 (N_16080,N_14359,N_14993);
xor U16081 (N_16081,N_14248,N_14901);
and U16082 (N_16082,N_13892,N_13891);
and U16083 (N_16083,N_13503,N_13882);
and U16084 (N_16084,N_14809,N_14028);
and U16085 (N_16085,N_13735,N_14978);
nor U16086 (N_16086,N_14566,N_14116);
xnor U16087 (N_16087,N_14436,N_13748);
nor U16088 (N_16088,N_13594,N_14207);
nand U16089 (N_16089,N_13807,N_14767);
nand U16090 (N_16090,N_14003,N_14271);
nand U16091 (N_16091,N_14529,N_13956);
nor U16092 (N_16092,N_13650,N_14473);
and U16093 (N_16093,N_14298,N_14729);
xnor U16094 (N_16094,N_14339,N_14074);
xor U16095 (N_16095,N_14144,N_14538);
xor U16096 (N_16096,N_14824,N_13948);
and U16097 (N_16097,N_13579,N_14453);
nor U16098 (N_16098,N_14173,N_14724);
and U16099 (N_16099,N_13915,N_13536);
and U16100 (N_16100,N_14507,N_14918);
and U16101 (N_16101,N_14107,N_14883);
nand U16102 (N_16102,N_13677,N_13545);
and U16103 (N_16103,N_13710,N_13677);
xnor U16104 (N_16104,N_14482,N_14563);
nor U16105 (N_16105,N_14505,N_13684);
nor U16106 (N_16106,N_14187,N_13672);
nor U16107 (N_16107,N_14179,N_13831);
or U16108 (N_16108,N_14862,N_13659);
and U16109 (N_16109,N_14402,N_13799);
nand U16110 (N_16110,N_14639,N_14689);
xor U16111 (N_16111,N_13900,N_14421);
xor U16112 (N_16112,N_14977,N_13643);
or U16113 (N_16113,N_14857,N_14691);
nand U16114 (N_16114,N_13953,N_14018);
nand U16115 (N_16115,N_13758,N_13527);
xnor U16116 (N_16116,N_14514,N_14290);
nand U16117 (N_16117,N_13563,N_13698);
nand U16118 (N_16118,N_14009,N_13655);
and U16119 (N_16119,N_13758,N_14217);
or U16120 (N_16120,N_13772,N_14734);
nand U16121 (N_16121,N_13845,N_14239);
xor U16122 (N_16122,N_14789,N_14062);
and U16123 (N_16123,N_13555,N_14358);
nand U16124 (N_16124,N_13792,N_13880);
nor U16125 (N_16125,N_14536,N_14490);
nor U16126 (N_16126,N_13780,N_13779);
xnor U16127 (N_16127,N_14779,N_14337);
nand U16128 (N_16128,N_13989,N_14598);
and U16129 (N_16129,N_13691,N_13652);
or U16130 (N_16130,N_14626,N_13818);
xor U16131 (N_16131,N_13982,N_14019);
xor U16132 (N_16132,N_14495,N_14844);
xor U16133 (N_16133,N_13821,N_14881);
xor U16134 (N_16134,N_14129,N_14008);
or U16135 (N_16135,N_14182,N_14831);
and U16136 (N_16136,N_13900,N_13769);
or U16137 (N_16137,N_14033,N_14531);
or U16138 (N_16138,N_13819,N_13683);
nand U16139 (N_16139,N_14034,N_14146);
nand U16140 (N_16140,N_13553,N_14700);
and U16141 (N_16141,N_14379,N_14112);
and U16142 (N_16142,N_13666,N_13655);
nand U16143 (N_16143,N_14761,N_14689);
nor U16144 (N_16144,N_14442,N_14952);
or U16145 (N_16145,N_13729,N_13530);
and U16146 (N_16146,N_14966,N_14417);
xnor U16147 (N_16147,N_14442,N_14240);
nand U16148 (N_16148,N_14559,N_14008);
xnor U16149 (N_16149,N_14180,N_14188);
and U16150 (N_16150,N_14519,N_14832);
and U16151 (N_16151,N_13605,N_13526);
xnor U16152 (N_16152,N_13910,N_14356);
nand U16153 (N_16153,N_14456,N_13903);
xor U16154 (N_16154,N_14912,N_14450);
nor U16155 (N_16155,N_14552,N_14788);
nand U16156 (N_16156,N_14588,N_13901);
nor U16157 (N_16157,N_13536,N_14651);
nand U16158 (N_16158,N_13623,N_14817);
nand U16159 (N_16159,N_14366,N_13789);
nor U16160 (N_16160,N_14037,N_14855);
nand U16161 (N_16161,N_14108,N_14872);
nor U16162 (N_16162,N_14428,N_14532);
xnor U16163 (N_16163,N_13692,N_14770);
and U16164 (N_16164,N_14753,N_14873);
nand U16165 (N_16165,N_14254,N_13804);
and U16166 (N_16166,N_14201,N_14399);
and U16167 (N_16167,N_14559,N_14087);
xnor U16168 (N_16168,N_14002,N_13851);
and U16169 (N_16169,N_14406,N_13987);
nand U16170 (N_16170,N_13860,N_14568);
xnor U16171 (N_16171,N_14303,N_14729);
nor U16172 (N_16172,N_14893,N_14645);
nor U16173 (N_16173,N_14912,N_14567);
or U16174 (N_16174,N_14617,N_13813);
nand U16175 (N_16175,N_14129,N_13580);
nand U16176 (N_16176,N_14685,N_13944);
and U16177 (N_16177,N_14427,N_13911);
xnor U16178 (N_16178,N_13627,N_14539);
xor U16179 (N_16179,N_14956,N_13651);
nand U16180 (N_16180,N_14624,N_14572);
nand U16181 (N_16181,N_14809,N_13842);
and U16182 (N_16182,N_14591,N_14789);
xor U16183 (N_16183,N_14940,N_14785);
nand U16184 (N_16184,N_13626,N_14307);
nor U16185 (N_16185,N_14060,N_14258);
xnor U16186 (N_16186,N_13679,N_13801);
xor U16187 (N_16187,N_13624,N_14136);
and U16188 (N_16188,N_14270,N_14487);
or U16189 (N_16189,N_14257,N_14696);
nand U16190 (N_16190,N_14287,N_14578);
nand U16191 (N_16191,N_14417,N_13862);
nand U16192 (N_16192,N_13549,N_14337);
or U16193 (N_16193,N_13921,N_13709);
xnor U16194 (N_16194,N_14573,N_13834);
or U16195 (N_16195,N_13531,N_14170);
and U16196 (N_16196,N_13778,N_14372);
or U16197 (N_16197,N_13537,N_14425);
and U16198 (N_16198,N_14512,N_13881);
or U16199 (N_16199,N_14737,N_14932);
and U16200 (N_16200,N_13837,N_13960);
nor U16201 (N_16201,N_13942,N_14304);
or U16202 (N_16202,N_14895,N_14754);
nand U16203 (N_16203,N_14810,N_13951);
nor U16204 (N_16204,N_14182,N_14550);
xor U16205 (N_16205,N_14804,N_14992);
and U16206 (N_16206,N_13756,N_14922);
and U16207 (N_16207,N_14997,N_14379);
xnor U16208 (N_16208,N_14588,N_13811);
xnor U16209 (N_16209,N_14779,N_13557);
xnor U16210 (N_16210,N_13649,N_14838);
nor U16211 (N_16211,N_13869,N_13586);
nand U16212 (N_16212,N_14336,N_14368);
nand U16213 (N_16213,N_14973,N_14391);
or U16214 (N_16214,N_13559,N_14167);
xor U16215 (N_16215,N_13642,N_14314);
and U16216 (N_16216,N_14792,N_14153);
or U16217 (N_16217,N_13906,N_13676);
nand U16218 (N_16218,N_14694,N_14652);
nor U16219 (N_16219,N_14032,N_13955);
or U16220 (N_16220,N_14791,N_13649);
nor U16221 (N_16221,N_14493,N_14622);
or U16222 (N_16222,N_13676,N_13547);
and U16223 (N_16223,N_13569,N_14789);
xnor U16224 (N_16224,N_13532,N_14460);
and U16225 (N_16225,N_14640,N_14772);
and U16226 (N_16226,N_14164,N_13691);
or U16227 (N_16227,N_13576,N_14114);
or U16228 (N_16228,N_13710,N_14670);
nor U16229 (N_16229,N_14581,N_13716);
xor U16230 (N_16230,N_14068,N_13634);
nor U16231 (N_16231,N_13712,N_14583);
xor U16232 (N_16232,N_14530,N_14124);
nand U16233 (N_16233,N_13508,N_14060);
and U16234 (N_16234,N_13668,N_14334);
or U16235 (N_16235,N_13607,N_13781);
nand U16236 (N_16236,N_14010,N_14724);
nor U16237 (N_16237,N_14388,N_14511);
and U16238 (N_16238,N_14186,N_14584);
nor U16239 (N_16239,N_14733,N_14869);
nor U16240 (N_16240,N_14110,N_13991);
nor U16241 (N_16241,N_14188,N_13794);
xor U16242 (N_16242,N_14803,N_14052);
nand U16243 (N_16243,N_14432,N_14907);
xor U16244 (N_16244,N_13576,N_14031);
or U16245 (N_16245,N_14434,N_14169);
and U16246 (N_16246,N_14991,N_14383);
xnor U16247 (N_16247,N_14223,N_14613);
nand U16248 (N_16248,N_14636,N_13730);
or U16249 (N_16249,N_14418,N_14121);
and U16250 (N_16250,N_14312,N_14013);
nand U16251 (N_16251,N_14166,N_13797);
nor U16252 (N_16252,N_13982,N_14701);
nand U16253 (N_16253,N_13733,N_14898);
nand U16254 (N_16254,N_13860,N_14413);
nand U16255 (N_16255,N_14089,N_13641);
or U16256 (N_16256,N_14349,N_14082);
nand U16257 (N_16257,N_14752,N_14919);
and U16258 (N_16258,N_14159,N_14760);
and U16259 (N_16259,N_13702,N_14654);
or U16260 (N_16260,N_14803,N_14307);
or U16261 (N_16261,N_14832,N_14767);
and U16262 (N_16262,N_14564,N_13668);
and U16263 (N_16263,N_14505,N_13653);
or U16264 (N_16264,N_13670,N_14901);
or U16265 (N_16265,N_14154,N_14184);
nor U16266 (N_16266,N_14964,N_14032);
and U16267 (N_16267,N_14237,N_14722);
or U16268 (N_16268,N_13519,N_14793);
nor U16269 (N_16269,N_14330,N_14757);
nand U16270 (N_16270,N_13919,N_13820);
xnor U16271 (N_16271,N_13616,N_13577);
nor U16272 (N_16272,N_14485,N_14186);
nand U16273 (N_16273,N_14469,N_13838);
or U16274 (N_16274,N_13835,N_14325);
or U16275 (N_16275,N_13898,N_14187);
and U16276 (N_16276,N_14439,N_13845);
and U16277 (N_16277,N_13913,N_13718);
nand U16278 (N_16278,N_14901,N_14062);
or U16279 (N_16279,N_14571,N_14865);
nand U16280 (N_16280,N_14785,N_14541);
nor U16281 (N_16281,N_13598,N_14404);
xor U16282 (N_16282,N_14487,N_14800);
and U16283 (N_16283,N_13969,N_14253);
xor U16284 (N_16284,N_13678,N_13563);
or U16285 (N_16285,N_13845,N_13982);
and U16286 (N_16286,N_13959,N_14982);
nor U16287 (N_16287,N_14016,N_13812);
or U16288 (N_16288,N_14084,N_13634);
xnor U16289 (N_16289,N_13621,N_13680);
nand U16290 (N_16290,N_14362,N_13823);
nand U16291 (N_16291,N_13562,N_14299);
xnor U16292 (N_16292,N_14070,N_14045);
or U16293 (N_16293,N_14611,N_14693);
nor U16294 (N_16294,N_14454,N_14794);
or U16295 (N_16295,N_14732,N_13753);
nor U16296 (N_16296,N_14626,N_13720);
or U16297 (N_16297,N_14578,N_13658);
nor U16298 (N_16298,N_13739,N_14724);
nor U16299 (N_16299,N_14088,N_14461);
or U16300 (N_16300,N_14008,N_13965);
nand U16301 (N_16301,N_14969,N_14617);
nand U16302 (N_16302,N_14463,N_14812);
or U16303 (N_16303,N_13745,N_14735);
or U16304 (N_16304,N_14921,N_13636);
xnor U16305 (N_16305,N_13659,N_13596);
nand U16306 (N_16306,N_13863,N_14602);
xor U16307 (N_16307,N_14552,N_14183);
or U16308 (N_16308,N_14023,N_14527);
and U16309 (N_16309,N_14618,N_13781);
or U16310 (N_16310,N_14769,N_14025);
xnor U16311 (N_16311,N_13972,N_14894);
and U16312 (N_16312,N_14646,N_14062);
and U16313 (N_16313,N_13759,N_14816);
or U16314 (N_16314,N_13880,N_14513);
nor U16315 (N_16315,N_13666,N_14903);
nor U16316 (N_16316,N_13623,N_14945);
and U16317 (N_16317,N_14229,N_14029);
nor U16318 (N_16318,N_14184,N_13606);
nand U16319 (N_16319,N_13885,N_13653);
and U16320 (N_16320,N_14888,N_14852);
xnor U16321 (N_16321,N_14576,N_13517);
or U16322 (N_16322,N_14797,N_13648);
nor U16323 (N_16323,N_14585,N_14660);
nor U16324 (N_16324,N_13862,N_14290);
xnor U16325 (N_16325,N_13503,N_13877);
and U16326 (N_16326,N_14484,N_13722);
and U16327 (N_16327,N_14030,N_13723);
and U16328 (N_16328,N_13980,N_14139);
nand U16329 (N_16329,N_13582,N_14259);
nor U16330 (N_16330,N_14949,N_13676);
or U16331 (N_16331,N_14147,N_14755);
nor U16332 (N_16332,N_14988,N_13592);
xnor U16333 (N_16333,N_14344,N_14766);
and U16334 (N_16334,N_13698,N_14895);
nand U16335 (N_16335,N_13907,N_14705);
or U16336 (N_16336,N_14539,N_13693);
nand U16337 (N_16337,N_13641,N_14402);
nor U16338 (N_16338,N_14749,N_14450);
xnor U16339 (N_16339,N_14621,N_14746);
and U16340 (N_16340,N_14173,N_13587);
nor U16341 (N_16341,N_14990,N_14885);
nand U16342 (N_16342,N_14594,N_14206);
and U16343 (N_16343,N_13983,N_13681);
nor U16344 (N_16344,N_14826,N_13822);
and U16345 (N_16345,N_14670,N_14262);
nor U16346 (N_16346,N_13702,N_14653);
or U16347 (N_16347,N_13689,N_13515);
and U16348 (N_16348,N_13837,N_14001);
nand U16349 (N_16349,N_14938,N_13569);
nor U16350 (N_16350,N_14726,N_14933);
nand U16351 (N_16351,N_14934,N_13819);
and U16352 (N_16352,N_13975,N_13656);
or U16353 (N_16353,N_14006,N_14292);
nand U16354 (N_16354,N_13978,N_14883);
nand U16355 (N_16355,N_14872,N_13808);
or U16356 (N_16356,N_13563,N_13905);
or U16357 (N_16357,N_14343,N_14782);
xnor U16358 (N_16358,N_14077,N_14286);
or U16359 (N_16359,N_14390,N_14553);
or U16360 (N_16360,N_13814,N_14474);
and U16361 (N_16361,N_14399,N_13739);
or U16362 (N_16362,N_13732,N_14915);
nor U16363 (N_16363,N_13616,N_13867);
xor U16364 (N_16364,N_14608,N_14691);
and U16365 (N_16365,N_14485,N_14700);
and U16366 (N_16366,N_13799,N_13977);
or U16367 (N_16367,N_14356,N_13950);
nor U16368 (N_16368,N_14585,N_13984);
nand U16369 (N_16369,N_14327,N_14273);
or U16370 (N_16370,N_14468,N_14197);
or U16371 (N_16371,N_14985,N_13530);
and U16372 (N_16372,N_14303,N_14008);
or U16373 (N_16373,N_13892,N_14948);
nor U16374 (N_16374,N_14559,N_14707);
and U16375 (N_16375,N_14402,N_14812);
and U16376 (N_16376,N_14823,N_14495);
xnor U16377 (N_16377,N_14455,N_13967);
and U16378 (N_16378,N_13970,N_14499);
xnor U16379 (N_16379,N_13541,N_14109);
xnor U16380 (N_16380,N_13743,N_14410);
xnor U16381 (N_16381,N_14422,N_13985);
nor U16382 (N_16382,N_14678,N_13971);
or U16383 (N_16383,N_14180,N_14936);
nand U16384 (N_16384,N_13631,N_14522);
nor U16385 (N_16385,N_14520,N_14403);
xnor U16386 (N_16386,N_14113,N_13837);
and U16387 (N_16387,N_14468,N_14713);
nand U16388 (N_16388,N_14125,N_14807);
and U16389 (N_16389,N_14355,N_14116);
and U16390 (N_16390,N_14208,N_14420);
and U16391 (N_16391,N_13658,N_14045);
nor U16392 (N_16392,N_14091,N_14107);
and U16393 (N_16393,N_13870,N_14346);
nand U16394 (N_16394,N_14731,N_14315);
or U16395 (N_16395,N_13781,N_14868);
and U16396 (N_16396,N_13514,N_13534);
or U16397 (N_16397,N_14963,N_14210);
nor U16398 (N_16398,N_14499,N_14084);
nor U16399 (N_16399,N_14494,N_14105);
nor U16400 (N_16400,N_14001,N_13947);
xnor U16401 (N_16401,N_14785,N_14310);
nor U16402 (N_16402,N_13671,N_14853);
xor U16403 (N_16403,N_14321,N_14945);
and U16404 (N_16404,N_13737,N_13771);
nand U16405 (N_16405,N_14761,N_14130);
nand U16406 (N_16406,N_14956,N_14866);
nor U16407 (N_16407,N_13885,N_14097);
nand U16408 (N_16408,N_13946,N_14016);
nand U16409 (N_16409,N_14889,N_14241);
xor U16410 (N_16410,N_14820,N_14573);
or U16411 (N_16411,N_13634,N_14967);
or U16412 (N_16412,N_14643,N_13792);
and U16413 (N_16413,N_14565,N_13927);
or U16414 (N_16414,N_14098,N_13732);
or U16415 (N_16415,N_14511,N_14455);
nor U16416 (N_16416,N_14682,N_13544);
nand U16417 (N_16417,N_14353,N_13658);
or U16418 (N_16418,N_14684,N_14165);
nand U16419 (N_16419,N_14730,N_13725);
nand U16420 (N_16420,N_14538,N_13707);
xor U16421 (N_16421,N_13893,N_14292);
nor U16422 (N_16422,N_14654,N_13513);
and U16423 (N_16423,N_14699,N_13906);
and U16424 (N_16424,N_14644,N_13792);
nor U16425 (N_16425,N_14880,N_14836);
nand U16426 (N_16426,N_14972,N_14590);
or U16427 (N_16427,N_14750,N_14419);
or U16428 (N_16428,N_14231,N_14825);
xor U16429 (N_16429,N_14819,N_14930);
xor U16430 (N_16430,N_14695,N_13904);
nand U16431 (N_16431,N_14270,N_13880);
nor U16432 (N_16432,N_14733,N_14095);
or U16433 (N_16433,N_13782,N_14959);
nand U16434 (N_16434,N_14381,N_14192);
nor U16435 (N_16435,N_14706,N_14110);
or U16436 (N_16436,N_13683,N_14173);
xor U16437 (N_16437,N_14863,N_14882);
or U16438 (N_16438,N_14236,N_14589);
and U16439 (N_16439,N_13795,N_13799);
xor U16440 (N_16440,N_13882,N_13951);
nor U16441 (N_16441,N_14870,N_14926);
and U16442 (N_16442,N_13592,N_14706);
xor U16443 (N_16443,N_14612,N_14539);
xor U16444 (N_16444,N_14071,N_13834);
and U16445 (N_16445,N_14122,N_14567);
xnor U16446 (N_16446,N_14527,N_14942);
nor U16447 (N_16447,N_14997,N_14327);
xnor U16448 (N_16448,N_14314,N_14928);
xnor U16449 (N_16449,N_13796,N_14033);
xor U16450 (N_16450,N_13623,N_14078);
or U16451 (N_16451,N_14420,N_13509);
nand U16452 (N_16452,N_13621,N_13884);
xor U16453 (N_16453,N_14570,N_14185);
and U16454 (N_16454,N_13890,N_14614);
and U16455 (N_16455,N_14007,N_14681);
and U16456 (N_16456,N_14233,N_13658);
xnor U16457 (N_16457,N_13753,N_14463);
nor U16458 (N_16458,N_13757,N_13673);
xor U16459 (N_16459,N_13691,N_13533);
nor U16460 (N_16460,N_14707,N_14623);
nor U16461 (N_16461,N_14114,N_14943);
nor U16462 (N_16462,N_14153,N_14998);
or U16463 (N_16463,N_14624,N_13755);
nor U16464 (N_16464,N_14924,N_14168);
xor U16465 (N_16465,N_14862,N_14662);
xor U16466 (N_16466,N_14216,N_14582);
nand U16467 (N_16467,N_14380,N_13557);
nor U16468 (N_16468,N_13968,N_14923);
and U16469 (N_16469,N_14362,N_13970);
nand U16470 (N_16470,N_14622,N_14744);
and U16471 (N_16471,N_14817,N_13794);
nand U16472 (N_16472,N_13837,N_14514);
nor U16473 (N_16473,N_14944,N_14713);
nand U16474 (N_16474,N_13873,N_14596);
nand U16475 (N_16475,N_14677,N_13935);
or U16476 (N_16476,N_14808,N_13575);
nand U16477 (N_16477,N_13968,N_14208);
nor U16478 (N_16478,N_13934,N_14266);
xnor U16479 (N_16479,N_14815,N_14499);
and U16480 (N_16480,N_14020,N_14894);
xnor U16481 (N_16481,N_14082,N_13743);
and U16482 (N_16482,N_14715,N_14412);
nor U16483 (N_16483,N_14651,N_14082);
nand U16484 (N_16484,N_13993,N_13834);
and U16485 (N_16485,N_13552,N_13712);
nor U16486 (N_16486,N_14643,N_14588);
xnor U16487 (N_16487,N_14494,N_13610);
xnor U16488 (N_16488,N_14552,N_14752);
xor U16489 (N_16489,N_14699,N_14915);
nor U16490 (N_16490,N_14553,N_14884);
nor U16491 (N_16491,N_13548,N_14057);
nand U16492 (N_16492,N_14476,N_14350);
and U16493 (N_16493,N_14803,N_13577);
xor U16494 (N_16494,N_14467,N_13941);
and U16495 (N_16495,N_13962,N_13666);
or U16496 (N_16496,N_14030,N_13689);
nand U16497 (N_16497,N_13896,N_14392);
or U16498 (N_16498,N_14094,N_14856);
and U16499 (N_16499,N_14180,N_14870);
or U16500 (N_16500,N_15603,N_16138);
nand U16501 (N_16501,N_15076,N_16320);
or U16502 (N_16502,N_15300,N_16217);
and U16503 (N_16503,N_16075,N_16426);
nand U16504 (N_16504,N_15859,N_16039);
and U16505 (N_16505,N_15381,N_15037);
nand U16506 (N_16506,N_16049,N_15971);
and U16507 (N_16507,N_15138,N_15715);
nand U16508 (N_16508,N_15288,N_16251);
and U16509 (N_16509,N_15703,N_15332);
and U16510 (N_16510,N_15224,N_15841);
and U16511 (N_16511,N_15519,N_15633);
xor U16512 (N_16512,N_16152,N_16370);
nor U16513 (N_16513,N_15311,N_16231);
and U16514 (N_16514,N_15092,N_15154);
nor U16515 (N_16515,N_16159,N_15686);
or U16516 (N_16516,N_16469,N_16275);
xnor U16517 (N_16517,N_16022,N_15094);
nor U16518 (N_16518,N_15369,N_16279);
xor U16519 (N_16519,N_16126,N_16488);
or U16520 (N_16520,N_15872,N_16015);
nor U16521 (N_16521,N_16074,N_15909);
nor U16522 (N_16522,N_16236,N_16172);
and U16523 (N_16523,N_16157,N_15817);
nand U16524 (N_16524,N_15487,N_16215);
xor U16525 (N_16525,N_15081,N_16286);
xor U16526 (N_16526,N_16062,N_15621);
and U16527 (N_16527,N_15934,N_15446);
nor U16528 (N_16528,N_15953,N_15478);
xor U16529 (N_16529,N_16086,N_15833);
or U16530 (N_16530,N_15191,N_16077);
and U16531 (N_16531,N_16476,N_15040);
nand U16532 (N_16532,N_15305,N_16165);
or U16533 (N_16533,N_15575,N_15577);
nor U16534 (N_16534,N_16403,N_15276);
and U16535 (N_16535,N_16479,N_15712);
and U16536 (N_16536,N_15629,N_16333);
or U16537 (N_16537,N_16404,N_15054);
or U16538 (N_16538,N_16250,N_15800);
nand U16539 (N_16539,N_16164,N_15752);
nand U16540 (N_16540,N_16495,N_15461);
or U16541 (N_16541,N_16253,N_16282);
nand U16542 (N_16542,N_16451,N_16263);
nand U16543 (N_16543,N_16471,N_16298);
xnor U16544 (N_16544,N_15198,N_16130);
xor U16545 (N_16545,N_15626,N_16027);
nor U16546 (N_16546,N_15088,N_15313);
xor U16547 (N_16547,N_16043,N_16428);
or U16548 (N_16548,N_15331,N_15738);
nor U16549 (N_16549,N_15214,N_15182);
nand U16550 (N_16550,N_16063,N_16432);
xor U16551 (N_16551,N_15901,N_15539);
nor U16552 (N_16552,N_16127,N_15551);
and U16553 (N_16553,N_16220,N_15125);
xor U16554 (N_16554,N_15257,N_16387);
nand U16555 (N_16555,N_15486,N_15969);
or U16556 (N_16556,N_15220,N_15212);
nand U16557 (N_16557,N_15156,N_15126);
or U16558 (N_16558,N_15618,N_16017);
nand U16559 (N_16559,N_15274,N_16323);
nand U16560 (N_16560,N_15380,N_15111);
xnor U16561 (N_16561,N_15516,N_15046);
or U16562 (N_16562,N_15496,N_15407);
or U16563 (N_16563,N_16407,N_15162);
nor U16564 (N_16564,N_15917,N_15860);
nor U16565 (N_16565,N_15824,N_15667);
xnor U16566 (N_16566,N_15634,N_15627);
nand U16567 (N_16567,N_15526,N_16416);
and U16568 (N_16568,N_15511,N_15748);
or U16569 (N_16569,N_16028,N_16460);
nand U16570 (N_16570,N_15883,N_15813);
xnor U16571 (N_16571,N_15199,N_15957);
nor U16572 (N_16572,N_16444,N_15882);
and U16573 (N_16573,N_16142,N_15109);
or U16574 (N_16574,N_16131,N_15064);
xor U16575 (N_16575,N_15253,N_15973);
nand U16576 (N_16576,N_15096,N_15783);
and U16577 (N_16577,N_16352,N_15339);
and U16578 (N_16578,N_15875,N_16485);
xnor U16579 (N_16579,N_16340,N_16041);
and U16580 (N_16580,N_16299,N_16170);
nand U16581 (N_16581,N_15733,N_15700);
or U16582 (N_16582,N_15421,N_16242);
nor U16583 (N_16583,N_15694,N_16035);
or U16584 (N_16584,N_16128,N_15013);
or U16585 (N_16585,N_15740,N_16259);
or U16586 (N_16586,N_16477,N_15206);
xor U16587 (N_16587,N_15753,N_16110);
and U16588 (N_16588,N_15312,N_16269);
or U16589 (N_16589,N_16174,N_15522);
xor U16590 (N_16590,N_15003,N_15583);
nor U16591 (N_16591,N_16154,N_15664);
nand U16592 (N_16592,N_15058,N_15683);
nor U16593 (N_16593,N_15786,N_15216);
and U16594 (N_16594,N_15816,N_15015);
or U16595 (N_16595,N_15590,N_16399);
xnor U16596 (N_16596,N_15405,N_15561);
and U16597 (N_16597,N_16365,N_15249);
nand U16598 (N_16598,N_15576,N_16106);
or U16599 (N_16599,N_16307,N_16067);
or U16600 (N_16600,N_16301,N_15586);
xor U16601 (N_16601,N_15255,N_16466);
or U16602 (N_16602,N_15924,N_15308);
nor U16603 (N_16603,N_15361,N_16442);
or U16604 (N_16604,N_16367,N_16045);
and U16605 (N_16605,N_15533,N_15788);
nor U16606 (N_16606,N_15028,N_16037);
and U16607 (N_16607,N_15525,N_16033);
and U16608 (N_16608,N_15853,N_16278);
or U16609 (N_16609,N_16099,N_15422);
or U16610 (N_16610,N_15245,N_15069);
nand U16611 (N_16611,N_15950,N_15676);
xnor U16612 (N_16612,N_15543,N_16085);
or U16613 (N_16613,N_15822,N_15981);
and U16614 (N_16614,N_15677,N_15523);
or U16615 (N_16615,N_15277,N_15579);
xor U16616 (N_16616,N_15404,N_16261);
xnor U16617 (N_16617,N_16197,N_15892);
nand U16618 (N_16618,N_15776,N_15649);
or U16619 (N_16619,N_15134,N_15679);
xor U16620 (N_16620,N_16003,N_15080);
xnor U16621 (N_16621,N_15920,N_15630);
nor U16622 (N_16622,N_16104,N_16338);
nor U16623 (N_16623,N_15747,N_16223);
xor U16624 (N_16624,N_15565,N_16235);
nor U16625 (N_16625,N_15855,N_15742);
nor U16626 (N_16626,N_15763,N_15432);
nand U16627 (N_16627,N_15647,N_16200);
and U16628 (N_16628,N_16392,N_15019);
nor U16629 (N_16629,N_15790,N_15002);
or U16630 (N_16630,N_16265,N_15884);
nand U16631 (N_16631,N_16313,N_15400);
nand U16632 (N_16632,N_15636,N_15434);
and U16633 (N_16633,N_15090,N_15394);
xor U16634 (N_16634,N_15409,N_15616);
nand U16635 (N_16635,N_15863,N_16010);
xnor U16636 (N_16636,N_15945,N_16443);
xor U16637 (N_16637,N_16397,N_15620);
nor U16638 (N_16638,N_16098,N_15357);
and U16639 (N_16639,N_16100,N_15508);
nor U16640 (N_16640,N_15371,N_15808);
nand U16641 (N_16641,N_15186,N_15267);
or U16642 (N_16642,N_15153,N_16198);
xor U16643 (N_16643,N_15250,N_15021);
and U16644 (N_16644,N_16424,N_16494);
xor U16645 (N_16645,N_15184,N_15903);
xor U16646 (N_16646,N_15190,N_16262);
and U16647 (N_16647,N_15470,N_15500);
nor U16648 (N_16648,N_15759,N_15897);
or U16649 (N_16649,N_16393,N_15463);
or U16650 (N_16650,N_15506,N_15646);
nand U16651 (N_16651,N_16321,N_15870);
nand U16652 (N_16652,N_16115,N_15704);
xor U16653 (N_16653,N_15902,N_16061);
nand U16654 (N_16654,N_15871,N_15730);
and U16655 (N_16655,N_15454,N_16285);
nand U16656 (N_16656,N_15417,N_15809);
and U16657 (N_16657,N_15567,N_16246);
and U16658 (N_16658,N_15702,N_16461);
nand U16659 (N_16659,N_15531,N_16047);
and U16660 (N_16660,N_15047,N_15607);
nor U16661 (N_16661,N_15864,N_15393);
nand U16662 (N_16662,N_15135,N_15885);
nand U16663 (N_16663,N_15062,N_15235);
nor U16664 (N_16664,N_15236,N_16328);
and U16665 (N_16665,N_15628,N_16491);
xnor U16666 (N_16666,N_15077,N_15197);
nand U16667 (N_16667,N_16454,N_15291);
or U16668 (N_16668,N_15681,N_15105);
xnor U16669 (N_16669,N_15761,N_15641);
nand U16670 (N_16670,N_15272,N_16457);
nor U16671 (N_16671,N_15513,N_16309);
or U16672 (N_16672,N_16341,N_15129);
or U16673 (N_16673,N_15472,N_15280);
and U16674 (N_16674,N_16468,N_16482);
xnor U16675 (N_16675,N_15782,N_15798);
xor U16676 (N_16676,N_15972,N_16336);
nand U16677 (N_16677,N_15563,N_16306);
xnor U16678 (N_16678,N_15209,N_16066);
nor U16679 (N_16679,N_15294,N_15152);
nand U16680 (N_16680,N_15874,N_15119);
xnor U16681 (N_16681,N_16401,N_15128);
nor U16682 (N_16682,N_15102,N_16327);
and U16683 (N_16683,N_15985,N_15919);
or U16684 (N_16684,N_15072,N_16032);
nor U16685 (N_16685,N_16023,N_16182);
nand U16686 (N_16686,N_15296,N_15203);
nor U16687 (N_16687,N_15990,N_15437);
xnor U16688 (N_16688,N_15839,N_16417);
nand U16689 (N_16689,N_16334,N_15710);
nand U16690 (N_16690,N_15247,N_15442);
xnor U16691 (N_16691,N_15682,N_15113);
xor U16692 (N_16692,N_15986,N_15244);
nand U16693 (N_16693,N_15321,N_15414);
xor U16694 (N_16694,N_15074,N_16020);
xor U16695 (N_16695,N_15123,N_15553);
or U16696 (N_16696,N_16402,N_16438);
or U16697 (N_16697,N_16410,N_15708);
nor U16698 (N_16698,N_16331,N_15701);
and U16699 (N_16699,N_15039,N_16178);
nand U16700 (N_16700,N_15388,N_15947);
nor U16701 (N_16701,N_16470,N_15755);
nor U16702 (N_16702,N_16400,N_16339);
nand U16703 (N_16703,N_15655,N_16146);
xnor U16704 (N_16704,N_16486,N_16216);
xor U16705 (N_16705,N_15427,N_15344);
nand U16706 (N_16706,N_16359,N_15643);
nor U16707 (N_16707,N_15354,N_15270);
xnor U16708 (N_16708,N_15671,N_15520);
xor U16709 (N_16709,N_15631,N_16084);
nor U16710 (N_16710,N_16069,N_15844);
nand U16711 (N_16711,N_16136,N_15443);
xnor U16712 (N_16712,N_15391,N_15876);
nor U16713 (N_16713,N_16330,N_15743);
or U16714 (N_16714,N_15145,N_15281);
nand U16715 (N_16715,N_16446,N_16219);
nor U16716 (N_16716,N_15222,N_15079);
and U16717 (N_16717,N_16463,N_16380);
and U16718 (N_16718,N_15852,N_15410);
xnor U16719 (N_16719,N_15491,N_16237);
xnor U16720 (N_16720,N_15570,N_15426);
and U16721 (N_16721,N_16496,N_15057);
or U16722 (N_16722,N_15115,N_16158);
xnor U16723 (N_16723,N_15205,N_15771);
or U16724 (N_16724,N_15796,N_15136);
or U16725 (N_16725,N_15044,N_15906);
nor U16726 (N_16726,N_15815,N_15322);
or U16727 (N_16727,N_15379,N_16427);
nand U16728 (N_16728,N_15569,N_15714);
and U16729 (N_16729,N_16009,N_15777);
nor U16730 (N_16730,N_16076,N_16267);
or U16731 (N_16731,N_15493,N_15043);
nor U16732 (N_16732,N_15795,N_15177);
nor U16733 (N_16733,N_16445,N_16291);
or U16734 (N_16734,N_15299,N_15595);
xnor U16735 (N_16735,N_15176,N_15401);
or U16736 (N_16736,N_15555,N_15159);
and U16737 (N_16737,N_16293,N_15794);
nor U16738 (N_16738,N_16021,N_15574);
and U16739 (N_16739,N_16283,N_15416);
nor U16740 (N_16740,N_15540,N_16042);
and U16741 (N_16741,N_16135,N_15286);
nor U16742 (N_16742,N_16412,N_15886);
or U16743 (N_16743,N_15928,N_15942);
nand U16744 (N_16744,N_16190,N_16053);
xnor U16745 (N_16745,N_15155,N_16305);
xor U16746 (N_16746,N_16490,N_16101);
nor U16747 (N_16747,N_16150,N_16430);
nand U16748 (N_16748,N_15887,N_16266);
xor U16749 (N_16749,N_16065,N_15665);
or U16750 (N_16750,N_16008,N_16078);
or U16751 (N_16751,N_16125,N_16120);
xor U16752 (N_16752,N_15507,N_15211);
nand U16753 (N_16753,N_15598,N_15801);
and U16754 (N_16754,N_15262,N_15638);
nand U16755 (N_16755,N_15256,N_16016);
nor U16756 (N_16756,N_15589,N_15617);
nand U16757 (N_16757,N_15325,N_16358);
or U16758 (N_16758,N_15615,N_16357);
and U16759 (N_16759,N_15012,N_15368);
or U16760 (N_16760,N_16222,N_15592);
and U16761 (N_16761,N_15370,N_15684);
or U16762 (N_16762,N_16249,N_15987);
nor U16763 (N_16763,N_15034,N_15071);
nand U16764 (N_16764,N_15541,N_16363);
and U16765 (N_16765,N_15314,N_15178);
nor U16766 (N_16766,N_16378,N_16292);
or U16767 (N_16767,N_16132,N_15122);
or U16768 (N_16768,N_15110,N_15904);
or U16769 (N_16769,N_15196,N_16360);
nor U16770 (N_16770,N_15004,N_15020);
or U16771 (N_16771,N_16089,N_15566);
or U16772 (N_16772,N_16189,N_15975);
nand U16773 (N_16773,N_15610,N_15818);
and U16774 (N_16774,N_15365,N_15834);
xnor U16775 (N_16775,N_15766,N_15830);
or U16776 (N_16776,N_15952,N_16173);
xnor U16777 (N_16777,N_15140,N_15221);
nor U16778 (N_16778,N_15208,N_16163);
and U16779 (N_16779,N_15678,N_15739);
nand U16780 (N_16780,N_15053,N_16284);
nor U16781 (N_16781,N_15049,N_15722);
nor U16782 (N_16782,N_15095,N_15226);
xor U16783 (N_16783,N_15218,N_15232);
xnor U16784 (N_16784,N_15440,N_15623);
or U16785 (N_16785,N_15735,N_15916);
or U16786 (N_16786,N_15915,N_15979);
nand U16787 (N_16787,N_15927,N_16413);
or U16788 (N_16788,N_16192,N_16398);
nand U16789 (N_16789,N_16090,N_16122);
or U16790 (N_16790,N_15754,N_16345);
xnor U16791 (N_16791,N_15041,N_15756);
and U16792 (N_16792,N_15489,N_16145);
and U16793 (N_16793,N_15358,N_16274);
nor U16794 (N_16794,N_16257,N_15348);
or U16795 (N_16795,N_16384,N_15545);
and U16796 (N_16796,N_15836,N_15444);
and U16797 (N_16797,N_15606,N_15991);
and U16798 (N_16798,N_15784,N_15423);
nand U16799 (N_16799,N_15572,N_15195);
xor U16800 (N_16800,N_16248,N_15130);
and U16801 (N_16801,N_16489,N_15499);
and U16802 (N_16802,N_15692,N_15303);
nand U16803 (N_16803,N_16083,N_15424);
nor U16804 (N_16804,N_15078,N_15117);
or U16805 (N_16805,N_15552,N_15494);
nor U16806 (N_16806,N_15173,N_15418);
nand U16807 (N_16807,N_15802,N_15768);
or U16808 (N_16808,N_16337,N_16386);
nand U16809 (N_16809,N_15112,N_15939);
nor U16810 (N_16810,N_15749,N_15832);
and U16811 (N_16811,N_16467,N_16119);
nor U16812 (N_16812,N_16255,N_15146);
xor U16813 (N_16813,N_15335,N_15293);
or U16814 (N_16814,N_15711,N_16361);
nor U16815 (N_16815,N_16177,N_15137);
or U16816 (N_16816,N_15689,N_15512);
nor U16817 (N_16817,N_15007,N_16272);
and U16818 (N_16818,N_16474,N_15227);
and U16819 (N_16819,N_15659,N_15382);
and U16820 (N_16820,N_15468,N_15896);
xor U16821 (N_16821,N_15502,N_16107);
xnor U16822 (N_16822,N_15982,N_15843);
nand U16823 (N_16823,N_15083,N_15068);
nand U16824 (N_16824,N_15086,N_15680);
nor U16825 (N_16825,N_15035,N_15477);
and U16826 (N_16826,N_15264,N_16013);
nand U16827 (N_16827,N_15150,N_16183);
xnor U16828 (N_16828,N_16419,N_15501);
nand U16829 (N_16829,N_15524,N_16472);
nor U16830 (N_16830,N_15419,N_16133);
xor U16831 (N_16831,N_15275,N_15160);
and U16832 (N_16832,N_16289,N_15658);
and U16833 (N_16833,N_16353,N_15793);
or U16834 (N_16834,N_16218,N_15429);
nand U16835 (N_16835,N_15403,N_15898);
nand U16836 (N_16836,N_15457,N_16184);
nor U16837 (N_16837,N_15447,N_16102);
nor U16838 (N_16838,N_15338,N_15022);
and U16839 (N_16839,N_15425,N_15148);
xnor U16840 (N_16840,N_15932,N_16350);
nor U16841 (N_16841,N_15387,N_16070);
nor U16842 (N_16842,N_16240,N_15485);
xor U16843 (N_16843,N_15030,N_16391);
or U16844 (N_16844,N_15736,N_15789);
and U16845 (N_16845,N_16459,N_15814);
nand U16846 (N_16846,N_15842,N_16295);
nor U16847 (N_16847,N_15283,N_15383);
nand U16848 (N_16848,N_15347,N_15827);
nor U16849 (N_16849,N_15869,N_16205);
xor U16850 (N_16850,N_15464,N_16388);
nor U16851 (N_16851,N_16207,N_15542);
or U16852 (N_16852,N_16036,N_15373);
and U16853 (N_16853,N_15231,N_15131);
nor U16854 (N_16854,N_15282,N_15171);
or U16855 (N_16855,N_16029,N_16319);
nor U16856 (N_16856,N_15453,N_15888);
nand U16857 (N_16857,N_15854,N_15549);
or U16858 (N_16858,N_16088,N_15479);
xnor U16859 (N_16859,N_15480,N_15336);
xnor U16860 (N_16860,N_15497,N_16004);
xnor U16861 (N_16861,N_15826,N_16091);
or U16862 (N_16862,N_15016,N_15352);
xor U16863 (N_16863,N_15573,N_15894);
and U16864 (N_16864,N_15873,N_16256);
and U16865 (N_16865,N_16314,N_15905);
and U16866 (N_16866,N_15023,N_15139);
nor U16867 (N_16867,N_16385,N_15609);
nor U16868 (N_16868,N_15510,N_16310);
or U16869 (N_16869,N_15612,N_15217);
xnor U16870 (N_16870,N_15670,N_15114);
nor U16871 (N_16871,N_16448,N_15835);
nand U16872 (N_16872,N_16143,N_15052);
nand U16873 (N_16873,N_15690,N_15124);
xor U16874 (N_16874,N_15900,N_15911);
nand U16875 (N_16875,N_15433,N_16019);
nand U16876 (N_16876,N_15614,N_16153);
and U16877 (N_16877,N_16332,N_15536);
nor U16878 (N_16878,N_15943,N_15765);
and U16879 (N_16879,N_15017,N_15439);
nand U16880 (N_16880,N_15101,N_15328);
and U16881 (N_16881,N_16124,N_15687);
or U16882 (N_16882,N_16281,N_15448);
or U16883 (N_16883,N_15170,N_15287);
nand U16884 (N_16884,N_16175,N_15997);
and U16885 (N_16885,N_15923,N_15718);
nand U16886 (N_16886,N_16300,N_15757);
and U16887 (N_16887,N_15849,N_15377);
or U16888 (N_16888,N_16429,N_15980);
or U16889 (N_16889,N_16434,N_16422);
and U16890 (N_16890,N_16245,N_15751);
nand U16891 (N_16891,N_15038,N_16453);
xor U16892 (N_16892,N_15261,N_15548);
nand U16893 (N_16893,N_15121,N_16287);
or U16894 (N_16894,N_15949,N_15838);
nand U16895 (N_16895,N_16317,N_15051);
nor U16896 (N_16896,N_15334,N_15922);
and U16897 (N_16897,N_15207,N_15964);
xnor U16898 (N_16898,N_16395,N_16156);
nor U16899 (N_16899,N_15600,N_15877);
nor U16900 (N_16900,N_16382,N_16093);
nor U16901 (N_16901,N_15865,N_16040);
or U16902 (N_16902,N_16421,N_15241);
and U16903 (N_16903,N_15251,N_15758);
or U16904 (N_16904,N_15880,N_15602);
nor U16905 (N_16905,N_15668,N_15709);
nand U16906 (N_16906,N_15451,N_15343);
or U16907 (N_16907,N_15812,N_16436);
and U16908 (N_16908,N_15165,N_15465);
xnor U16909 (N_16909,N_16465,N_16326);
or U16910 (N_16910,N_15116,N_15360);
or U16911 (N_16911,N_16221,N_15104);
or U16912 (N_16912,N_15716,N_15108);
and U16913 (N_16913,N_15935,N_15717);
nor U16914 (N_16914,N_15133,N_15645);
xor U16915 (N_16915,N_16418,N_15469);
nor U16916 (N_16916,N_15557,N_16046);
nor U16917 (N_16917,N_16176,N_15306);
nor U16918 (N_16918,N_15862,N_15913);
xnor U16919 (N_16919,N_16288,N_15554);
nor U16920 (N_16920,N_15158,N_15831);
or U16921 (N_16921,N_16073,N_16194);
nand U16922 (N_16922,N_16423,N_15958);
or U16923 (N_16923,N_15662,N_15910);
or U16924 (N_16924,N_15055,N_15596);
or U16925 (N_16925,N_15639,N_15045);
nor U16926 (N_16926,N_15989,N_15385);
nor U16927 (N_16927,N_16377,N_16038);
nand U16928 (N_16928,N_15324,N_16225);
or U16929 (N_16929,N_15697,N_15201);
nand U16930 (N_16930,N_15803,N_16208);
or U16931 (N_16931,N_15430,N_16097);
and U16932 (N_16932,N_16082,N_15144);
and U16933 (N_16933,N_15652,N_16280);
and U16934 (N_16934,N_16121,N_15132);
nor U16935 (N_16935,N_15825,N_15696);
or U16936 (N_16936,N_15799,N_15406);
xnor U16937 (N_16937,N_15390,N_16057);
nand U16938 (N_16938,N_15940,N_15234);
xnor U16939 (N_16939,N_16068,N_16484);
xor U16940 (N_16940,N_15537,N_16000);
or U16941 (N_16941,N_15141,N_16396);
or U16942 (N_16942,N_15781,N_16243);
or U16943 (N_16943,N_15240,N_16195);
nor U16944 (N_16944,N_16180,N_15562);
nand U16945 (N_16945,N_16228,N_15026);
nand U16946 (N_16946,N_15315,N_15149);
nand U16947 (N_16947,N_15285,N_15867);
or U16948 (N_16948,N_15319,N_15725);
nand U16949 (N_16949,N_15413,N_16449);
and U16950 (N_16950,N_15588,N_15775);
nand U16951 (N_16951,N_15415,N_15168);
or U16952 (N_16952,N_15669,N_16343);
and U16953 (N_16953,N_16206,N_15961);
nand U16954 (N_16954,N_15329,N_15219);
nor U16955 (N_16955,N_16230,N_15558);
nor U16956 (N_16956,N_15837,N_16113);
and U16957 (N_16957,N_15091,N_15265);
xor U16958 (N_16958,N_15587,N_15359);
and U16959 (N_16959,N_15346,N_16234);
xnor U16960 (N_16960,N_16139,N_15402);
nor U16961 (N_16961,N_15918,N_15840);
nand U16962 (N_16962,N_15693,N_15938);
nor U16963 (N_16963,N_16227,N_16167);
nand U16964 (N_16964,N_16433,N_15481);
or U16965 (N_16965,N_15084,N_16059);
xor U16966 (N_16966,N_15951,N_15847);
and U16967 (N_16967,N_15921,N_15509);
nand U16968 (N_16968,N_15977,N_15597);
nor U16969 (N_16969,N_15611,N_15650);
nand U16970 (N_16970,N_15345,N_16191);
or U16971 (N_16971,N_15466,N_16425);
nand U16972 (N_16972,N_15750,N_15036);
xor U16973 (N_16973,N_15675,N_15225);
or U16974 (N_16974,N_15372,N_16498);
and U16975 (N_16975,N_15356,N_15169);
xor U16976 (N_16976,N_16092,N_15243);
nor U16977 (N_16977,N_16268,N_16052);
or U16978 (N_16978,N_16364,N_16303);
or U16979 (N_16979,N_15698,N_16487);
nand U16980 (N_16980,N_15237,N_15828);
and U16981 (N_16981,N_15778,N_15550);
or U16982 (N_16982,N_15821,N_15956);
or U16983 (N_16983,N_15157,N_16405);
or U16984 (N_16984,N_16497,N_15933);
and U16985 (N_16985,N_15948,N_15707);
or U16986 (N_16986,N_15666,N_16018);
and U16987 (N_16987,N_15899,N_16409);
xor U16988 (N_16988,N_15441,N_16050);
nor U16989 (N_16989,N_15723,N_15966);
xor U16990 (N_16990,N_15857,N_15163);
or U16991 (N_16991,N_16270,N_15632);
and U16992 (N_16992,N_16369,N_15866);
or U16993 (N_16993,N_16411,N_16224);
nor U16994 (N_16994,N_15528,N_16187);
nor U16995 (N_16995,N_15762,N_15672);
nor U16996 (N_16996,N_16315,N_15366);
xnor U16997 (N_16997,N_16229,N_16081);
nor U16998 (N_16998,N_16342,N_15396);
or U16999 (N_16999,N_16080,N_15529);
and U17000 (N_17000,N_15648,N_15353);
nand U17001 (N_17001,N_15498,N_15556);
or U17002 (N_17002,N_15992,N_15881);
nand U17003 (N_17003,N_15653,N_15151);
nor U17004 (N_17004,N_15504,N_15323);
nand U17005 (N_17005,N_15326,N_15355);
or U17006 (N_17006,N_16149,N_15926);
nor U17007 (N_17007,N_15295,N_16161);
and U17008 (N_17008,N_15238,N_15999);
nand U17009 (N_17009,N_16064,N_16406);
or U17010 (N_17010,N_15066,N_16366);
nor U17011 (N_17011,N_15823,N_15000);
and U17012 (N_17012,N_15011,N_15908);
or U17013 (N_17013,N_16114,N_15488);
nand U17014 (N_17014,N_16351,N_15029);
xor U17015 (N_17015,N_15582,N_15591);
nand U17016 (N_17016,N_15118,N_16140);
and U17017 (N_17017,N_15791,N_16455);
and U17018 (N_17018,N_16051,N_15228);
xor U17019 (N_17019,N_15067,N_15063);
nor U17020 (N_17020,N_15374,N_15517);
nand U17021 (N_17021,N_16437,N_15024);
nand U17022 (N_17022,N_16232,N_15010);
xnor U17023 (N_17023,N_15780,N_15518);
and U17024 (N_17024,N_15848,N_15578);
nand U17025 (N_17025,N_16464,N_15252);
and U17026 (N_17026,N_16002,N_15258);
nand U17027 (N_17027,N_15937,N_15931);
nand U17028 (N_17028,N_16079,N_16493);
and U17029 (N_17029,N_15087,N_15774);
or U17030 (N_17030,N_15744,N_15787);
xor U17031 (N_17031,N_15266,N_15375);
and U17032 (N_17032,N_15333,N_15161);
or U17033 (N_17033,N_16024,N_16095);
or U17034 (N_17034,N_15891,N_16129);
or U17035 (N_17035,N_16329,N_15976);
or U17036 (N_17036,N_15605,N_15890);
nand U17037 (N_17037,N_15613,N_15732);
or U17038 (N_17038,N_15560,N_15398);
nor U17039 (N_17039,N_16390,N_16296);
and U17040 (N_17040,N_16054,N_15770);
nor U17041 (N_17041,N_15340,N_15056);
or U17042 (N_17042,N_15955,N_15963);
nor U17043 (N_17043,N_15811,N_15483);
xor U17044 (N_17044,N_16211,N_16210);
nor U17045 (N_17045,N_16007,N_15005);
nand U17046 (N_17046,N_15449,N_15376);
nor U17047 (N_17047,N_15797,N_15351);
or U17048 (N_17048,N_16186,N_15785);
xnor U17049 (N_17049,N_16111,N_15025);
and U17050 (N_17050,N_15490,N_15175);
nand U17051 (N_17051,N_16462,N_15093);
or U17052 (N_17052,N_16096,N_15246);
xnor U17053 (N_17053,N_15213,N_16151);
and U17054 (N_17054,N_15445,N_15399);
or U17055 (N_17055,N_16214,N_15967);
or U17056 (N_17056,N_15279,N_16316);
and U17057 (N_17057,N_15965,N_15929);
nand U17058 (N_17058,N_15856,N_16117);
xor U17059 (N_17059,N_16318,N_15637);
and U17060 (N_17060,N_15089,N_15959);
nor U17061 (N_17061,N_16346,N_15189);
nor U17062 (N_17062,N_16264,N_15691);
nand U17063 (N_17063,N_15559,N_15484);
nor U17064 (N_17064,N_15193,N_15408);
or U17065 (N_17065,N_15893,N_15914);
and U17066 (N_17066,N_16254,N_15100);
and U17067 (N_17067,N_15996,N_15065);
or U17068 (N_17068,N_15097,N_16044);
nor U17069 (N_17069,N_15584,N_15741);
nor U17070 (N_17070,N_16260,N_16103);
nand U17071 (N_17071,N_15660,N_15458);
or U17072 (N_17072,N_15688,N_15106);
or U17073 (N_17073,N_15059,N_15450);
or U17074 (N_17074,N_15642,N_15673);
nor U17075 (N_17075,N_15179,N_15438);
or U17076 (N_17076,N_15622,N_15546);
or U17077 (N_17077,N_16308,N_15970);
xor U17078 (N_17078,N_15014,N_16277);
or U17079 (N_17079,N_15395,N_15378);
nand U17080 (N_17080,N_15930,N_15292);
nand U17081 (N_17081,N_15720,N_16233);
and U17082 (N_17082,N_15297,N_16025);
or U17083 (N_17083,N_15164,N_15107);
and U17084 (N_17084,N_16492,N_16499);
xnor U17085 (N_17085,N_15362,N_15601);
or U17086 (N_17086,N_15174,N_16420);
or U17087 (N_17087,N_16030,N_16238);
nor U17088 (N_17088,N_16108,N_16123);
and U17089 (N_17089,N_15188,N_16355);
nand U17090 (N_17090,N_15482,N_15230);
nor U17091 (N_17091,N_16302,N_15654);
or U17092 (N_17092,N_16447,N_15310);
or U17093 (N_17093,N_15731,N_16247);
and U17094 (N_17094,N_15459,N_16431);
xnor U17095 (N_17095,N_16118,N_16325);
and U17096 (N_17096,N_15263,N_15239);
xnor U17097 (N_17097,N_15316,N_16169);
xor U17098 (N_17098,N_15006,N_15127);
or U17099 (N_17099,N_16144,N_16199);
nor U17100 (N_17100,N_16375,N_15724);
or U17101 (N_17101,N_15644,N_16297);
and U17102 (N_17102,N_15183,N_15033);
xor U17103 (N_17103,N_16389,N_16112);
or U17104 (N_17104,N_16322,N_15185);
or U17105 (N_17105,N_15767,N_16204);
xor U17106 (N_17106,N_16202,N_16273);
nand U17107 (N_17107,N_15503,N_15290);
or U17108 (N_17108,N_15495,N_16356);
or U17109 (N_17109,N_16034,N_15850);
nor U17110 (N_17110,N_16155,N_16212);
or U17111 (N_17111,N_15941,N_15706);
or U17112 (N_17112,N_15846,N_15363);
or U17113 (N_17113,N_15473,N_15721);
or U17114 (N_17114,N_16087,N_15142);
nor U17115 (N_17115,N_15968,N_15544);
or U17116 (N_17116,N_16005,N_15284);
xnor U17117 (N_17117,N_15663,N_16371);
and U17118 (N_17118,N_15269,N_15745);
and U17119 (N_17119,N_15779,N_16258);
xnor U17120 (N_17120,N_15229,N_15215);
nor U17121 (N_17121,N_15187,N_16324);
or U17122 (N_17122,N_15350,N_15492);
nor U17123 (N_17123,N_16372,N_16148);
and U17124 (N_17124,N_15223,N_15307);
and U17125 (N_17125,N_15436,N_15367);
xor U17126 (N_17126,N_15851,N_16383);
and U17127 (N_17127,N_15527,N_15460);
nand U17128 (N_17128,N_16379,N_15719);
and U17129 (N_17129,N_15397,N_16012);
nor U17130 (N_17130,N_16440,N_16137);
xor U17131 (N_17131,N_16188,N_15384);
nand U17132 (N_17132,N_15534,N_15599);
nor U17133 (N_17133,N_15925,N_15298);
and U17134 (N_17134,N_15727,N_15978);
or U17135 (N_17135,N_15060,N_16160);
xor U17136 (N_17136,N_15167,N_15571);
and U17137 (N_17137,N_15661,N_16252);
nor U17138 (N_17138,N_15845,N_16026);
nor U17139 (N_17139,N_15858,N_15624);
and U17140 (N_17140,N_15505,N_15760);
or U17141 (N_17141,N_15073,N_15580);
nor U17142 (N_17142,N_16179,N_15820);
and U17143 (N_17143,N_16311,N_15764);
and U17144 (N_17144,N_15521,N_16031);
xnor U17145 (N_17145,N_16480,N_15120);
xnor U17146 (N_17146,N_15829,N_16349);
or U17147 (N_17147,N_15538,N_15705);
nor U17148 (N_17148,N_15386,N_15946);
and U17149 (N_17149,N_15085,N_16414);
nand U17150 (N_17150,N_16006,N_15805);
and U17151 (N_17151,N_16335,N_16071);
nor U17152 (N_17152,N_16381,N_16141);
nand U17153 (N_17153,N_15868,N_15268);
or U17154 (N_17154,N_15713,N_15772);
nand U17155 (N_17155,N_16415,N_15912);
nor U17156 (N_17156,N_15954,N_15050);
nand U17157 (N_17157,N_15515,N_15983);
xnor U17158 (N_17158,N_15420,N_16109);
nand U17159 (N_17159,N_15773,N_15192);
and U17160 (N_17160,N_15640,N_15181);
xnor U17161 (N_17161,N_15320,N_15301);
xor U17162 (N_17162,N_16456,N_15242);
xor U17163 (N_17163,N_15018,N_15172);
and U17164 (N_17164,N_15456,N_15027);
or U17165 (N_17165,N_15593,N_15042);
or U17166 (N_17166,N_16209,N_15233);
and U17167 (N_17167,N_15431,N_15734);
and U17168 (N_17168,N_15364,N_16394);
xnor U17169 (N_17169,N_16473,N_15810);
and U17170 (N_17170,N_16475,N_16271);
xnor U17171 (N_17171,N_15304,N_15674);
nand U17172 (N_17172,N_16304,N_15342);
nor U17173 (N_17173,N_16276,N_15260);
nand U17174 (N_17174,N_15075,N_15452);
nor U17175 (N_17175,N_15194,N_15535);
or U17176 (N_17176,N_15435,N_15210);
xnor U17177 (N_17177,N_16376,N_15962);
and U17178 (N_17178,N_16056,N_16185);
or U17179 (N_17179,N_15988,N_15082);
nand U17180 (N_17180,N_15728,N_15317);
and U17181 (N_17181,N_15455,N_15532);
or U17182 (N_17182,N_16344,N_15289);
xor U17183 (N_17183,N_16441,N_15993);
and U17184 (N_17184,N_15467,N_16168);
nand U17185 (N_17185,N_15302,N_16226);
and U17186 (N_17186,N_16181,N_15254);
xnor U17187 (N_17187,N_16203,N_15984);
nor U17188 (N_17188,N_15604,N_15608);
xor U17189 (N_17189,N_16290,N_15878);
nor U17190 (N_17190,N_16196,N_15585);
and U17191 (N_17191,N_15514,N_15994);
nor U17192 (N_17192,N_15568,N_16213);
nand U17193 (N_17193,N_15048,N_16239);
and U17194 (N_17194,N_15726,N_16134);
and U17195 (N_17195,N_16094,N_16450);
xor U17196 (N_17196,N_15807,N_15936);
and U17197 (N_17197,N_15806,N_15009);
and U17198 (N_17198,N_15737,N_16439);
nand U17199 (N_17199,N_15944,N_15031);
nand U17200 (N_17200,N_15995,N_15907);
and U17201 (N_17201,N_16348,N_15998);
or U17202 (N_17202,N_16373,N_16478);
or U17203 (N_17203,N_16193,N_15547);
nor U17204 (N_17204,N_15327,N_16312);
and U17205 (N_17205,N_15098,N_15143);
or U17206 (N_17206,N_16166,N_15769);
xnor U17207 (N_17207,N_15273,N_15389);
and U17208 (N_17208,N_16483,N_15619);
nand U17209 (N_17209,N_16171,N_15099);
nand U17210 (N_17210,N_16060,N_15960);
xnor U17211 (N_17211,N_15792,N_15476);
and U17212 (N_17212,N_16458,N_15337);
xnor U17213 (N_17213,N_16001,N_16435);
and U17214 (N_17214,N_15349,N_15103);
xor U17215 (N_17215,N_16162,N_15341);
xnor U17216 (N_17216,N_15428,N_15695);
xor U17217 (N_17217,N_15746,N_15581);
xor U17218 (N_17218,N_15974,N_15412);
xnor U17219 (N_17219,N_16105,N_16452);
xor U17220 (N_17220,N_15625,N_16116);
and U17221 (N_17221,N_15202,N_16408);
xor U17222 (N_17222,N_16481,N_15474);
nor U17223 (N_17223,N_15309,N_15657);
xnor U17224 (N_17224,N_15475,N_16072);
or U17225 (N_17225,N_15564,N_15861);
nor U17226 (N_17226,N_15392,N_15008);
or U17227 (N_17227,N_15147,N_16147);
nand U17228 (N_17228,N_16055,N_15070);
and U17229 (N_17229,N_16014,N_15530);
or U17230 (N_17230,N_15259,N_15200);
or U17231 (N_17231,N_16011,N_15204);
nand U17232 (N_17232,N_15278,N_15819);
and U17233 (N_17233,N_15271,N_16058);
and U17234 (N_17234,N_15656,N_15061);
or U17235 (N_17235,N_15879,N_16048);
xor U17236 (N_17236,N_15462,N_15594);
or U17237 (N_17237,N_16368,N_15804);
xnor U17238 (N_17238,N_16347,N_16201);
nand U17239 (N_17239,N_15685,N_15699);
xnor U17240 (N_17240,N_15001,N_16294);
nor U17241 (N_17241,N_15411,N_15651);
or U17242 (N_17242,N_16241,N_16354);
nor U17243 (N_17243,N_15895,N_15248);
or U17244 (N_17244,N_16362,N_15729);
xnor U17245 (N_17245,N_16244,N_15166);
and U17246 (N_17246,N_15318,N_15471);
nor U17247 (N_17247,N_15635,N_16374);
xor U17248 (N_17248,N_15180,N_15032);
nor U17249 (N_17249,N_15330,N_15889);
nand U17250 (N_17250,N_15467,N_16315);
nand U17251 (N_17251,N_15512,N_15842);
and U17252 (N_17252,N_15563,N_16371);
and U17253 (N_17253,N_15752,N_15264);
and U17254 (N_17254,N_15206,N_15767);
xnor U17255 (N_17255,N_15223,N_15099);
nor U17256 (N_17256,N_15308,N_15935);
xor U17257 (N_17257,N_16271,N_15962);
nor U17258 (N_17258,N_15255,N_16454);
or U17259 (N_17259,N_15999,N_16377);
and U17260 (N_17260,N_15281,N_15322);
or U17261 (N_17261,N_15968,N_16027);
nand U17262 (N_17262,N_15589,N_16191);
or U17263 (N_17263,N_16283,N_16280);
or U17264 (N_17264,N_15687,N_16388);
and U17265 (N_17265,N_15249,N_15988);
nand U17266 (N_17266,N_16365,N_15416);
nor U17267 (N_17267,N_15521,N_15879);
or U17268 (N_17268,N_15598,N_15884);
or U17269 (N_17269,N_15223,N_15438);
and U17270 (N_17270,N_15707,N_15559);
nand U17271 (N_17271,N_15391,N_15895);
nand U17272 (N_17272,N_15994,N_16085);
or U17273 (N_17273,N_15925,N_15426);
and U17274 (N_17274,N_15866,N_15153);
and U17275 (N_17275,N_16243,N_15811);
nand U17276 (N_17276,N_15562,N_15191);
xnor U17277 (N_17277,N_15097,N_16472);
nor U17278 (N_17278,N_15113,N_15367);
nor U17279 (N_17279,N_15306,N_16005);
nand U17280 (N_17280,N_15778,N_15966);
and U17281 (N_17281,N_15320,N_15434);
nand U17282 (N_17282,N_15619,N_15412);
and U17283 (N_17283,N_16484,N_15731);
nor U17284 (N_17284,N_15817,N_16215);
or U17285 (N_17285,N_15102,N_15259);
nor U17286 (N_17286,N_15999,N_16431);
xor U17287 (N_17287,N_16133,N_15266);
or U17288 (N_17288,N_15184,N_16441);
and U17289 (N_17289,N_15257,N_15204);
nor U17290 (N_17290,N_16106,N_16098);
or U17291 (N_17291,N_16180,N_15122);
and U17292 (N_17292,N_15071,N_15173);
or U17293 (N_17293,N_15173,N_16199);
or U17294 (N_17294,N_15037,N_16445);
nand U17295 (N_17295,N_15370,N_16310);
nand U17296 (N_17296,N_16297,N_15562);
xnor U17297 (N_17297,N_15071,N_16333);
and U17298 (N_17298,N_16355,N_16196);
or U17299 (N_17299,N_16114,N_15417);
or U17300 (N_17300,N_15180,N_15935);
nand U17301 (N_17301,N_16145,N_16110);
xor U17302 (N_17302,N_16467,N_15302);
nor U17303 (N_17303,N_16187,N_16232);
nor U17304 (N_17304,N_15357,N_16483);
xor U17305 (N_17305,N_15038,N_15034);
nand U17306 (N_17306,N_16217,N_15111);
nor U17307 (N_17307,N_15060,N_16483);
nand U17308 (N_17308,N_15752,N_15153);
nand U17309 (N_17309,N_15449,N_16160);
and U17310 (N_17310,N_15282,N_15312);
or U17311 (N_17311,N_15590,N_15087);
nor U17312 (N_17312,N_15271,N_15865);
xor U17313 (N_17313,N_15150,N_16242);
nor U17314 (N_17314,N_15709,N_15258);
or U17315 (N_17315,N_16349,N_15731);
xor U17316 (N_17316,N_15257,N_15621);
and U17317 (N_17317,N_16137,N_16495);
or U17318 (N_17318,N_15088,N_16298);
xor U17319 (N_17319,N_15493,N_15580);
nand U17320 (N_17320,N_15728,N_16454);
and U17321 (N_17321,N_16189,N_15158);
or U17322 (N_17322,N_15679,N_15391);
or U17323 (N_17323,N_15764,N_15793);
nor U17324 (N_17324,N_16323,N_16062);
nor U17325 (N_17325,N_15111,N_16319);
xor U17326 (N_17326,N_15047,N_16054);
nor U17327 (N_17327,N_15820,N_15431);
xor U17328 (N_17328,N_15192,N_15517);
nand U17329 (N_17329,N_16365,N_16377);
nor U17330 (N_17330,N_15177,N_15739);
xnor U17331 (N_17331,N_16297,N_15472);
and U17332 (N_17332,N_15899,N_15300);
nor U17333 (N_17333,N_16336,N_15684);
nor U17334 (N_17334,N_16102,N_16121);
or U17335 (N_17335,N_15825,N_15760);
or U17336 (N_17336,N_15448,N_16173);
and U17337 (N_17337,N_16359,N_15530);
and U17338 (N_17338,N_15564,N_15969);
nor U17339 (N_17339,N_15608,N_16158);
nand U17340 (N_17340,N_15719,N_15303);
xor U17341 (N_17341,N_15305,N_15701);
or U17342 (N_17342,N_15621,N_15781);
or U17343 (N_17343,N_16463,N_15522);
or U17344 (N_17344,N_15116,N_16407);
nand U17345 (N_17345,N_15853,N_15635);
or U17346 (N_17346,N_15638,N_16415);
and U17347 (N_17347,N_15121,N_16073);
and U17348 (N_17348,N_16038,N_15553);
xnor U17349 (N_17349,N_16278,N_16215);
nand U17350 (N_17350,N_16126,N_15151);
and U17351 (N_17351,N_15475,N_15615);
and U17352 (N_17352,N_15748,N_15889);
and U17353 (N_17353,N_16470,N_15032);
and U17354 (N_17354,N_16299,N_15391);
and U17355 (N_17355,N_15010,N_16038);
or U17356 (N_17356,N_15563,N_15676);
or U17357 (N_17357,N_15994,N_16476);
or U17358 (N_17358,N_15241,N_15353);
and U17359 (N_17359,N_15838,N_15231);
nor U17360 (N_17360,N_15599,N_16208);
and U17361 (N_17361,N_15590,N_15704);
nor U17362 (N_17362,N_16348,N_16218);
and U17363 (N_17363,N_16252,N_16006);
nand U17364 (N_17364,N_16176,N_15804);
or U17365 (N_17365,N_15695,N_15931);
xnor U17366 (N_17366,N_15493,N_15052);
or U17367 (N_17367,N_15237,N_15176);
nand U17368 (N_17368,N_15407,N_15140);
and U17369 (N_17369,N_15735,N_15922);
and U17370 (N_17370,N_16216,N_15280);
nand U17371 (N_17371,N_15996,N_15031);
nor U17372 (N_17372,N_15065,N_15157);
or U17373 (N_17373,N_15494,N_15815);
xnor U17374 (N_17374,N_15363,N_15880);
nand U17375 (N_17375,N_15701,N_15000);
and U17376 (N_17376,N_15775,N_16299);
or U17377 (N_17377,N_15167,N_15064);
nor U17378 (N_17378,N_15567,N_16309);
xnor U17379 (N_17379,N_15488,N_16108);
xor U17380 (N_17380,N_16005,N_15556);
xor U17381 (N_17381,N_16278,N_15709);
nand U17382 (N_17382,N_15072,N_15748);
and U17383 (N_17383,N_15818,N_15615);
and U17384 (N_17384,N_15630,N_15898);
nor U17385 (N_17385,N_16460,N_15539);
and U17386 (N_17386,N_16228,N_16158);
and U17387 (N_17387,N_15729,N_15480);
nor U17388 (N_17388,N_15596,N_15301);
and U17389 (N_17389,N_15902,N_15638);
nor U17390 (N_17390,N_15765,N_16263);
nand U17391 (N_17391,N_15171,N_16079);
xor U17392 (N_17392,N_15242,N_15484);
or U17393 (N_17393,N_15021,N_15508);
xor U17394 (N_17394,N_16291,N_16160);
nand U17395 (N_17395,N_15490,N_15518);
or U17396 (N_17396,N_15724,N_15694);
xnor U17397 (N_17397,N_15958,N_16102);
xor U17398 (N_17398,N_15590,N_16472);
xnor U17399 (N_17399,N_15467,N_16233);
or U17400 (N_17400,N_15770,N_16283);
xor U17401 (N_17401,N_15827,N_15181);
or U17402 (N_17402,N_15130,N_16086);
nand U17403 (N_17403,N_15811,N_15831);
nand U17404 (N_17404,N_15655,N_15146);
and U17405 (N_17405,N_15451,N_16487);
nor U17406 (N_17406,N_15478,N_15824);
or U17407 (N_17407,N_15396,N_15942);
xnor U17408 (N_17408,N_15679,N_15000);
nor U17409 (N_17409,N_15346,N_16131);
nand U17410 (N_17410,N_15885,N_16280);
nor U17411 (N_17411,N_15679,N_15480);
xnor U17412 (N_17412,N_16434,N_16243);
nand U17413 (N_17413,N_15961,N_16376);
nor U17414 (N_17414,N_16484,N_15268);
nand U17415 (N_17415,N_16202,N_15626);
nor U17416 (N_17416,N_15501,N_15608);
nor U17417 (N_17417,N_15184,N_16114);
nand U17418 (N_17418,N_15401,N_15456);
nand U17419 (N_17419,N_15108,N_15029);
and U17420 (N_17420,N_15513,N_15344);
nand U17421 (N_17421,N_16369,N_16342);
or U17422 (N_17422,N_15434,N_16202);
and U17423 (N_17423,N_15516,N_15681);
or U17424 (N_17424,N_16424,N_15291);
or U17425 (N_17425,N_15213,N_15714);
nand U17426 (N_17426,N_15906,N_15963);
nand U17427 (N_17427,N_16215,N_15404);
or U17428 (N_17428,N_16382,N_15759);
xnor U17429 (N_17429,N_15349,N_15345);
nor U17430 (N_17430,N_15754,N_16225);
nand U17431 (N_17431,N_15574,N_16118);
nor U17432 (N_17432,N_16255,N_15634);
nand U17433 (N_17433,N_15084,N_15029);
nor U17434 (N_17434,N_15908,N_16347);
nor U17435 (N_17435,N_15892,N_15252);
nor U17436 (N_17436,N_15390,N_15619);
and U17437 (N_17437,N_16049,N_15232);
or U17438 (N_17438,N_15826,N_15107);
nor U17439 (N_17439,N_16049,N_15857);
nand U17440 (N_17440,N_15924,N_15463);
or U17441 (N_17441,N_15550,N_16472);
nand U17442 (N_17442,N_15528,N_15001);
nand U17443 (N_17443,N_15040,N_15233);
or U17444 (N_17444,N_15110,N_15081);
xnor U17445 (N_17445,N_15525,N_15194);
and U17446 (N_17446,N_15550,N_15980);
and U17447 (N_17447,N_15522,N_16099);
nand U17448 (N_17448,N_15927,N_15298);
or U17449 (N_17449,N_15108,N_15457);
and U17450 (N_17450,N_15776,N_16007);
nand U17451 (N_17451,N_15991,N_15270);
or U17452 (N_17452,N_16238,N_15674);
xnor U17453 (N_17453,N_15113,N_16145);
nor U17454 (N_17454,N_15084,N_16080);
nor U17455 (N_17455,N_16208,N_15745);
nand U17456 (N_17456,N_15633,N_15770);
nor U17457 (N_17457,N_15345,N_15090);
nand U17458 (N_17458,N_15909,N_15846);
nor U17459 (N_17459,N_16477,N_15784);
xor U17460 (N_17460,N_15634,N_15885);
nor U17461 (N_17461,N_16155,N_16036);
and U17462 (N_17462,N_15078,N_15537);
or U17463 (N_17463,N_15085,N_16075);
nor U17464 (N_17464,N_15490,N_15591);
nor U17465 (N_17465,N_15686,N_15436);
nor U17466 (N_17466,N_15104,N_16232);
and U17467 (N_17467,N_15901,N_15557);
nor U17468 (N_17468,N_15745,N_16245);
nor U17469 (N_17469,N_15267,N_15376);
nor U17470 (N_17470,N_15732,N_16260);
and U17471 (N_17471,N_15693,N_16216);
nand U17472 (N_17472,N_15565,N_15288);
xor U17473 (N_17473,N_15304,N_16234);
nand U17474 (N_17474,N_15843,N_16220);
nand U17475 (N_17475,N_15952,N_15055);
xnor U17476 (N_17476,N_16353,N_16236);
nor U17477 (N_17477,N_15842,N_16456);
and U17478 (N_17478,N_16168,N_15071);
and U17479 (N_17479,N_16256,N_16404);
or U17480 (N_17480,N_15844,N_15432);
nor U17481 (N_17481,N_15154,N_15466);
xnor U17482 (N_17482,N_16098,N_15523);
nor U17483 (N_17483,N_16270,N_16064);
xnor U17484 (N_17484,N_15160,N_16012);
or U17485 (N_17485,N_15209,N_15650);
xor U17486 (N_17486,N_16147,N_16481);
nor U17487 (N_17487,N_15496,N_15356);
and U17488 (N_17488,N_15149,N_15228);
or U17489 (N_17489,N_15090,N_15574);
nand U17490 (N_17490,N_15373,N_15236);
and U17491 (N_17491,N_15907,N_15904);
xnor U17492 (N_17492,N_15781,N_15042);
and U17493 (N_17493,N_15057,N_15003);
and U17494 (N_17494,N_15565,N_15649);
nor U17495 (N_17495,N_16369,N_15608);
nand U17496 (N_17496,N_15499,N_15778);
nand U17497 (N_17497,N_15111,N_15257);
nand U17498 (N_17498,N_15069,N_16009);
or U17499 (N_17499,N_16170,N_15390);
nor U17500 (N_17500,N_16271,N_15822);
or U17501 (N_17501,N_15690,N_15220);
nor U17502 (N_17502,N_15684,N_15428);
or U17503 (N_17503,N_16233,N_15518);
or U17504 (N_17504,N_15519,N_15484);
nand U17505 (N_17505,N_15590,N_15755);
and U17506 (N_17506,N_16263,N_15768);
or U17507 (N_17507,N_16056,N_16096);
and U17508 (N_17508,N_15534,N_15383);
or U17509 (N_17509,N_16040,N_15473);
nand U17510 (N_17510,N_15040,N_16105);
nor U17511 (N_17511,N_16161,N_15978);
and U17512 (N_17512,N_16273,N_16149);
nand U17513 (N_17513,N_15519,N_16474);
or U17514 (N_17514,N_16093,N_15195);
nor U17515 (N_17515,N_16108,N_15215);
xor U17516 (N_17516,N_15230,N_15065);
nor U17517 (N_17517,N_16206,N_15275);
nor U17518 (N_17518,N_16160,N_15700);
or U17519 (N_17519,N_15237,N_15555);
nand U17520 (N_17520,N_15583,N_15926);
or U17521 (N_17521,N_16434,N_16005);
and U17522 (N_17522,N_15503,N_15412);
nand U17523 (N_17523,N_15132,N_15478);
and U17524 (N_17524,N_16407,N_15946);
and U17525 (N_17525,N_16119,N_15740);
xnor U17526 (N_17526,N_16449,N_15388);
xnor U17527 (N_17527,N_15201,N_16340);
and U17528 (N_17528,N_16159,N_15533);
xnor U17529 (N_17529,N_15407,N_15260);
nand U17530 (N_17530,N_16332,N_15796);
nor U17531 (N_17531,N_15940,N_16203);
and U17532 (N_17532,N_15357,N_15782);
xnor U17533 (N_17533,N_15131,N_16317);
nor U17534 (N_17534,N_15591,N_15546);
xor U17535 (N_17535,N_15666,N_15946);
nand U17536 (N_17536,N_15781,N_15392);
or U17537 (N_17537,N_16367,N_15250);
and U17538 (N_17538,N_15267,N_15253);
and U17539 (N_17539,N_16199,N_15302);
xor U17540 (N_17540,N_15943,N_15939);
or U17541 (N_17541,N_16404,N_15565);
nand U17542 (N_17542,N_15471,N_15132);
or U17543 (N_17543,N_16281,N_15029);
nor U17544 (N_17544,N_15274,N_15520);
or U17545 (N_17545,N_16361,N_15934);
nand U17546 (N_17546,N_15404,N_16031);
and U17547 (N_17547,N_16204,N_15528);
and U17548 (N_17548,N_16415,N_16389);
and U17549 (N_17549,N_15626,N_16059);
xnor U17550 (N_17550,N_15842,N_15322);
and U17551 (N_17551,N_16425,N_15370);
nor U17552 (N_17552,N_15785,N_16006);
xor U17553 (N_17553,N_15810,N_16165);
or U17554 (N_17554,N_15411,N_15034);
nand U17555 (N_17555,N_15614,N_15205);
nand U17556 (N_17556,N_15693,N_16210);
and U17557 (N_17557,N_15058,N_15367);
nor U17558 (N_17558,N_15514,N_16291);
nor U17559 (N_17559,N_16482,N_16200);
xor U17560 (N_17560,N_15463,N_16226);
xnor U17561 (N_17561,N_15887,N_16452);
and U17562 (N_17562,N_15561,N_16452);
nand U17563 (N_17563,N_15490,N_15106);
nor U17564 (N_17564,N_16401,N_15281);
or U17565 (N_17565,N_16175,N_16198);
nor U17566 (N_17566,N_15235,N_15871);
or U17567 (N_17567,N_15406,N_15620);
xnor U17568 (N_17568,N_16287,N_16250);
or U17569 (N_17569,N_15169,N_15721);
nand U17570 (N_17570,N_16136,N_15906);
nand U17571 (N_17571,N_15550,N_16457);
nor U17572 (N_17572,N_15880,N_15108);
and U17573 (N_17573,N_15819,N_15219);
xor U17574 (N_17574,N_16118,N_15897);
nor U17575 (N_17575,N_15930,N_15144);
or U17576 (N_17576,N_16189,N_15096);
xor U17577 (N_17577,N_15429,N_16180);
nand U17578 (N_17578,N_15705,N_15040);
and U17579 (N_17579,N_16485,N_15263);
xor U17580 (N_17580,N_15089,N_15779);
xnor U17581 (N_17581,N_15366,N_15428);
and U17582 (N_17582,N_16342,N_15857);
nor U17583 (N_17583,N_15716,N_15110);
or U17584 (N_17584,N_16374,N_16023);
nand U17585 (N_17585,N_15944,N_15729);
nor U17586 (N_17586,N_15045,N_15721);
nand U17587 (N_17587,N_16111,N_15449);
and U17588 (N_17588,N_15712,N_15923);
and U17589 (N_17589,N_16475,N_15114);
or U17590 (N_17590,N_16024,N_15759);
and U17591 (N_17591,N_16183,N_16472);
and U17592 (N_17592,N_15881,N_15134);
or U17593 (N_17593,N_15142,N_15518);
nand U17594 (N_17594,N_15431,N_16251);
nor U17595 (N_17595,N_15078,N_15209);
xnor U17596 (N_17596,N_15380,N_15884);
and U17597 (N_17597,N_16425,N_15086);
and U17598 (N_17598,N_16450,N_16018);
or U17599 (N_17599,N_15896,N_15145);
or U17600 (N_17600,N_15611,N_16416);
nor U17601 (N_17601,N_15795,N_15555);
nand U17602 (N_17602,N_16138,N_16180);
and U17603 (N_17603,N_15962,N_16284);
and U17604 (N_17604,N_15875,N_16335);
or U17605 (N_17605,N_15930,N_15726);
nor U17606 (N_17606,N_16444,N_16326);
nand U17607 (N_17607,N_15834,N_15670);
xor U17608 (N_17608,N_15811,N_15139);
or U17609 (N_17609,N_15590,N_15583);
and U17610 (N_17610,N_15038,N_15272);
and U17611 (N_17611,N_15814,N_15812);
and U17612 (N_17612,N_15516,N_15876);
and U17613 (N_17613,N_16421,N_16387);
or U17614 (N_17614,N_16377,N_16395);
nand U17615 (N_17615,N_16247,N_15889);
or U17616 (N_17616,N_15708,N_15433);
nor U17617 (N_17617,N_16237,N_16117);
and U17618 (N_17618,N_15246,N_15385);
or U17619 (N_17619,N_15229,N_15613);
or U17620 (N_17620,N_15493,N_16183);
nand U17621 (N_17621,N_15444,N_16357);
nor U17622 (N_17622,N_16215,N_15322);
nor U17623 (N_17623,N_16192,N_16230);
xor U17624 (N_17624,N_15743,N_15224);
or U17625 (N_17625,N_16235,N_16294);
xor U17626 (N_17626,N_16097,N_16206);
nor U17627 (N_17627,N_15449,N_15822);
or U17628 (N_17628,N_15790,N_15181);
xor U17629 (N_17629,N_15992,N_15755);
nand U17630 (N_17630,N_15280,N_15151);
xnor U17631 (N_17631,N_16192,N_15720);
nand U17632 (N_17632,N_15234,N_15410);
nand U17633 (N_17633,N_16116,N_15479);
or U17634 (N_17634,N_15971,N_15532);
or U17635 (N_17635,N_15500,N_15256);
nor U17636 (N_17636,N_15982,N_15367);
and U17637 (N_17637,N_15227,N_16432);
or U17638 (N_17638,N_15646,N_16409);
and U17639 (N_17639,N_15082,N_16328);
and U17640 (N_17640,N_16146,N_15180);
nor U17641 (N_17641,N_15684,N_15699);
xnor U17642 (N_17642,N_16031,N_15548);
and U17643 (N_17643,N_15991,N_16461);
nor U17644 (N_17644,N_15903,N_15805);
and U17645 (N_17645,N_15599,N_15448);
or U17646 (N_17646,N_15943,N_15341);
nand U17647 (N_17647,N_16435,N_16303);
and U17648 (N_17648,N_15967,N_15162);
and U17649 (N_17649,N_16190,N_15747);
or U17650 (N_17650,N_15361,N_15596);
or U17651 (N_17651,N_15146,N_16123);
or U17652 (N_17652,N_15824,N_15318);
nor U17653 (N_17653,N_16130,N_15924);
nand U17654 (N_17654,N_15866,N_15033);
and U17655 (N_17655,N_15447,N_15753);
nand U17656 (N_17656,N_16281,N_15399);
xor U17657 (N_17657,N_15838,N_15181);
nor U17658 (N_17658,N_15023,N_15493);
xnor U17659 (N_17659,N_15254,N_16136);
xor U17660 (N_17660,N_15527,N_15110);
nand U17661 (N_17661,N_15568,N_16013);
nand U17662 (N_17662,N_16061,N_15574);
and U17663 (N_17663,N_15884,N_15327);
or U17664 (N_17664,N_15957,N_16145);
and U17665 (N_17665,N_15943,N_16417);
or U17666 (N_17666,N_15113,N_16149);
and U17667 (N_17667,N_15437,N_15045);
nor U17668 (N_17668,N_15048,N_16069);
and U17669 (N_17669,N_16354,N_16029);
xnor U17670 (N_17670,N_15939,N_16323);
and U17671 (N_17671,N_16024,N_16248);
nor U17672 (N_17672,N_15404,N_15258);
nor U17673 (N_17673,N_15012,N_16448);
or U17674 (N_17674,N_15115,N_15849);
and U17675 (N_17675,N_15442,N_15998);
nor U17676 (N_17676,N_15030,N_16255);
nor U17677 (N_17677,N_15238,N_16296);
nand U17678 (N_17678,N_15323,N_15328);
xnor U17679 (N_17679,N_15139,N_15798);
and U17680 (N_17680,N_15734,N_15736);
and U17681 (N_17681,N_15659,N_16271);
nand U17682 (N_17682,N_16381,N_15561);
xor U17683 (N_17683,N_16176,N_15528);
and U17684 (N_17684,N_15129,N_16065);
nor U17685 (N_17685,N_16030,N_15447);
nand U17686 (N_17686,N_16321,N_15792);
nand U17687 (N_17687,N_15122,N_16434);
nand U17688 (N_17688,N_15185,N_15151);
xor U17689 (N_17689,N_15918,N_16137);
nand U17690 (N_17690,N_15765,N_15560);
and U17691 (N_17691,N_16240,N_16372);
nand U17692 (N_17692,N_16470,N_16182);
or U17693 (N_17693,N_16261,N_16452);
nor U17694 (N_17694,N_15470,N_16285);
and U17695 (N_17695,N_15444,N_15422);
nand U17696 (N_17696,N_15935,N_15047);
and U17697 (N_17697,N_15047,N_15684);
nand U17698 (N_17698,N_15950,N_16202);
and U17699 (N_17699,N_16430,N_15795);
or U17700 (N_17700,N_15265,N_15388);
nor U17701 (N_17701,N_16197,N_16375);
xor U17702 (N_17702,N_16368,N_15364);
xor U17703 (N_17703,N_16038,N_16189);
and U17704 (N_17704,N_16321,N_15235);
or U17705 (N_17705,N_16056,N_15308);
and U17706 (N_17706,N_16243,N_15600);
xnor U17707 (N_17707,N_15738,N_16387);
nor U17708 (N_17708,N_15190,N_15119);
and U17709 (N_17709,N_15448,N_15508);
or U17710 (N_17710,N_15428,N_15024);
and U17711 (N_17711,N_16228,N_15544);
or U17712 (N_17712,N_15136,N_15719);
nand U17713 (N_17713,N_15392,N_16096);
xor U17714 (N_17714,N_15307,N_16478);
nor U17715 (N_17715,N_16008,N_15291);
nand U17716 (N_17716,N_15711,N_15964);
nand U17717 (N_17717,N_15922,N_15134);
nand U17718 (N_17718,N_15144,N_16219);
nand U17719 (N_17719,N_16468,N_16151);
and U17720 (N_17720,N_15358,N_15170);
or U17721 (N_17721,N_15382,N_15185);
and U17722 (N_17722,N_16363,N_15540);
or U17723 (N_17723,N_15393,N_15527);
nand U17724 (N_17724,N_15217,N_16478);
xnor U17725 (N_17725,N_15671,N_15525);
nand U17726 (N_17726,N_16071,N_15972);
xnor U17727 (N_17727,N_15709,N_15409);
nor U17728 (N_17728,N_15138,N_16108);
or U17729 (N_17729,N_15432,N_15920);
nor U17730 (N_17730,N_15139,N_16353);
and U17731 (N_17731,N_15036,N_16253);
nand U17732 (N_17732,N_16358,N_15233);
xnor U17733 (N_17733,N_16315,N_15160);
and U17734 (N_17734,N_16121,N_15117);
or U17735 (N_17735,N_15624,N_15628);
xor U17736 (N_17736,N_16327,N_15609);
or U17737 (N_17737,N_15393,N_15267);
and U17738 (N_17738,N_15642,N_15231);
xnor U17739 (N_17739,N_15659,N_16326);
nand U17740 (N_17740,N_16039,N_15350);
and U17741 (N_17741,N_16360,N_16005);
and U17742 (N_17742,N_15268,N_15021);
nor U17743 (N_17743,N_15761,N_15254);
xnor U17744 (N_17744,N_16406,N_15296);
xor U17745 (N_17745,N_15597,N_15551);
nor U17746 (N_17746,N_15230,N_15937);
xnor U17747 (N_17747,N_16308,N_15560);
nand U17748 (N_17748,N_16000,N_16334);
nand U17749 (N_17749,N_16451,N_16255);
nand U17750 (N_17750,N_16085,N_16225);
and U17751 (N_17751,N_15814,N_16135);
nand U17752 (N_17752,N_16044,N_15812);
or U17753 (N_17753,N_16445,N_15049);
nand U17754 (N_17754,N_15851,N_15669);
xor U17755 (N_17755,N_15275,N_15191);
nand U17756 (N_17756,N_15638,N_16106);
xor U17757 (N_17757,N_15638,N_15556);
nand U17758 (N_17758,N_16092,N_15568);
xnor U17759 (N_17759,N_15795,N_15689);
xor U17760 (N_17760,N_15227,N_16252);
nor U17761 (N_17761,N_15793,N_15059);
xor U17762 (N_17762,N_15705,N_15496);
nand U17763 (N_17763,N_16021,N_15839);
or U17764 (N_17764,N_15491,N_16282);
and U17765 (N_17765,N_15228,N_16081);
nand U17766 (N_17766,N_15708,N_15873);
nand U17767 (N_17767,N_16162,N_15440);
xnor U17768 (N_17768,N_15035,N_15051);
xnor U17769 (N_17769,N_16203,N_16197);
nand U17770 (N_17770,N_15319,N_16361);
xor U17771 (N_17771,N_16122,N_16064);
nor U17772 (N_17772,N_15382,N_16116);
nand U17773 (N_17773,N_15232,N_15702);
or U17774 (N_17774,N_15583,N_15348);
or U17775 (N_17775,N_16407,N_16050);
nand U17776 (N_17776,N_15004,N_15381);
and U17777 (N_17777,N_15038,N_15786);
and U17778 (N_17778,N_15380,N_15548);
xnor U17779 (N_17779,N_16385,N_15983);
and U17780 (N_17780,N_15295,N_15904);
and U17781 (N_17781,N_15116,N_15606);
nand U17782 (N_17782,N_15520,N_15455);
or U17783 (N_17783,N_15701,N_15372);
or U17784 (N_17784,N_15750,N_15148);
xnor U17785 (N_17785,N_15652,N_16190);
and U17786 (N_17786,N_15098,N_15731);
nor U17787 (N_17787,N_15032,N_15536);
or U17788 (N_17788,N_15599,N_15132);
or U17789 (N_17789,N_16499,N_15298);
nand U17790 (N_17790,N_16041,N_16494);
or U17791 (N_17791,N_15637,N_15825);
nor U17792 (N_17792,N_16326,N_16221);
xnor U17793 (N_17793,N_15284,N_15592);
xnor U17794 (N_17794,N_15368,N_16033);
and U17795 (N_17795,N_15838,N_15699);
and U17796 (N_17796,N_16258,N_16426);
or U17797 (N_17797,N_15593,N_16496);
or U17798 (N_17798,N_15574,N_15289);
nand U17799 (N_17799,N_15174,N_15732);
nor U17800 (N_17800,N_15295,N_15676);
xnor U17801 (N_17801,N_15567,N_15211);
or U17802 (N_17802,N_15679,N_16395);
or U17803 (N_17803,N_15487,N_15784);
and U17804 (N_17804,N_15539,N_16307);
nor U17805 (N_17805,N_15060,N_16378);
nor U17806 (N_17806,N_15351,N_16444);
and U17807 (N_17807,N_15691,N_15610);
and U17808 (N_17808,N_15239,N_15943);
and U17809 (N_17809,N_16297,N_15475);
nand U17810 (N_17810,N_15390,N_15986);
nor U17811 (N_17811,N_15917,N_15198);
and U17812 (N_17812,N_16014,N_15311);
xor U17813 (N_17813,N_15008,N_15477);
or U17814 (N_17814,N_15897,N_15148);
xnor U17815 (N_17815,N_15803,N_16284);
xnor U17816 (N_17816,N_15754,N_16487);
xor U17817 (N_17817,N_15382,N_15109);
or U17818 (N_17818,N_15858,N_16139);
xor U17819 (N_17819,N_15704,N_15126);
nand U17820 (N_17820,N_16358,N_15890);
or U17821 (N_17821,N_16448,N_15696);
nor U17822 (N_17822,N_16351,N_15077);
nand U17823 (N_17823,N_15313,N_15689);
nor U17824 (N_17824,N_16062,N_15946);
nand U17825 (N_17825,N_15765,N_15304);
nor U17826 (N_17826,N_16025,N_16158);
nor U17827 (N_17827,N_15151,N_15409);
nor U17828 (N_17828,N_15015,N_16164);
nor U17829 (N_17829,N_15497,N_16407);
nand U17830 (N_17830,N_15388,N_15051);
or U17831 (N_17831,N_16424,N_15304);
nor U17832 (N_17832,N_15471,N_15365);
or U17833 (N_17833,N_15715,N_16494);
or U17834 (N_17834,N_15492,N_15849);
nand U17835 (N_17835,N_15293,N_15504);
nand U17836 (N_17836,N_15699,N_15921);
and U17837 (N_17837,N_15969,N_15768);
xor U17838 (N_17838,N_15084,N_16461);
nand U17839 (N_17839,N_15998,N_16077);
nand U17840 (N_17840,N_15254,N_15285);
xor U17841 (N_17841,N_16125,N_16141);
nand U17842 (N_17842,N_16092,N_15503);
and U17843 (N_17843,N_15062,N_15264);
xor U17844 (N_17844,N_15286,N_15661);
nand U17845 (N_17845,N_16328,N_15733);
xor U17846 (N_17846,N_16063,N_15365);
and U17847 (N_17847,N_15534,N_15574);
or U17848 (N_17848,N_15794,N_16276);
and U17849 (N_17849,N_15386,N_15057);
nand U17850 (N_17850,N_15509,N_15725);
nor U17851 (N_17851,N_16247,N_16085);
nor U17852 (N_17852,N_16191,N_15564);
nand U17853 (N_17853,N_16473,N_16179);
xnor U17854 (N_17854,N_16216,N_15556);
nand U17855 (N_17855,N_16446,N_15304);
or U17856 (N_17856,N_15058,N_15643);
xnor U17857 (N_17857,N_15613,N_15829);
and U17858 (N_17858,N_16424,N_15594);
nand U17859 (N_17859,N_16211,N_15544);
nor U17860 (N_17860,N_15951,N_16409);
nor U17861 (N_17861,N_15709,N_15869);
nor U17862 (N_17862,N_15744,N_15998);
nor U17863 (N_17863,N_16040,N_15311);
and U17864 (N_17864,N_16175,N_15396);
nor U17865 (N_17865,N_15088,N_15732);
or U17866 (N_17866,N_16117,N_16047);
nand U17867 (N_17867,N_16210,N_15137);
nor U17868 (N_17868,N_16109,N_15745);
nor U17869 (N_17869,N_16243,N_15228);
nor U17870 (N_17870,N_15125,N_15953);
nand U17871 (N_17871,N_15108,N_15458);
xnor U17872 (N_17872,N_16191,N_15654);
nor U17873 (N_17873,N_15064,N_16341);
xor U17874 (N_17874,N_16067,N_15842);
xor U17875 (N_17875,N_15046,N_15250);
and U17876 (N_17876,N_15115,N_15065);
nand U17877 (N_17877,N_15028,N_15448);
xnor U17878 (N_17878,N_15808,N_15342);
and U17879 (N_17879,N_16312,N_15711);
and U17880 (N_17880,N_15448,N_16215);
nand U17881 (N_17881,N_15199,N_16252);
nor U17882 (N_17882,N_15615,N_15154);
xnor U17883 (N_17883,N_16414,N_15388);
or U17884 (N_17884,N_15725,N_15603);
and U17885 (N_17885,N_15400,N_15837);
nand U17886 (N_17886,N_16236,N_16315);
xor U17887 (N_17887,N_16394,N_15338);
nor U17888 (N_17888,N_15162,N_15863);
or U17889 (N_17889,N_16347,N_15686);
and U17890 (N_17890,N_15697,N_16234);
or U17891 (N_17891,N_16275,N_15989);
and U17892 (N_17892,N_16169,N_15605);
xor U17893 (N_17893,N_15979,N_15885);
and U17894 (N_17894,N_15722,N_16008);
nor U17895 (N_17895,N_15258,N_15741);
and U17896 (N_17896,N_16428,N_15385);
or U17897 (N_17897,N_15787,N_15502);
nor U17898 (N_17898,N_15948,N_15796);
nor U17899 (N_17899,N_16111,N_16436);
nand U17900 (N_17900,N_15058,N_16058);
nor U17901 (N_17901,N_15723,N_16435);
xnor U17902 (N_17902,N_16088,N_15261);
or U17903 (N_17903,N_15228,N_15924);
and U17904 (N_17904,N_15965,N_16491);
nor U17905 (N_17905,N_16329,N_15522);
or U17906 (N_17906,N_15664,N_16047);
nor U17907 (N_17907,N_15996,N_15910);
and U17908 (N_17908,N_16447,N_16022);
xnor U17909 (N_17909,N_16156,N_15446);
xnor U17910 (N_17910,N_15312,N_15773);
or U17911 (N_17911,N_15798,N_15906);
nor U17912 (N_17912,N_15625,N_15034);
nand U17913 (N_17913,N_15883,N_15333);
or U17914 (N_17914,N_15244,N_16320);
nor U17915 (N_17915,N_15759,N_16355);
nor U17916 (N_17916,N_15298,N_15140);
xnor U17917 (N_17917,N_16269,N_16075);
or U17918 (N_17918,N_15317,N_15598);
nand U17919 (N_17919,N_15214,N_15871);
or U17920 (N_17920,N_16356,N_15952);
xor U17921 (N_17921,N_15286,N_16210);
xnor U17922 (N_17922,N_15448,N_15435);
xor U17923 (N_17923,N_15961,N_16239);
or U17924 (N_17924,N_15146,N_16317);
nor U17925 (N_17925,N_15511,N_15281);
or U17926 (N_17926,N_15314,N_16061);
or U17927 (N_17927,N_15938,N_16150);
nor U17928 (N_17928,N_15810,N_15694);
nand U17929 (N_17929,N_15307,N_16192);
nand U17930 (N_17930,N_15175,N_15917);
and U17931 (N_17931,N_15741,N_15923);
nor U17932 (N_17932,N_15330,N_16137);
and U17933 (N_17933,N_15110,N_15870);
and U17934 (N_17934,N_16073,N_15793);
or U17935 (N_17935,N_15746,N_15044);
and U17936 (N_17936,N_15363,N_15923);
xor U17937 (N_17937,N_15627,N_15936);
xnor U17938 (N_17938,N_16117,N_16333);
nand U17939 (N_17939,N_16192,N_16006);
or U17940 (N_17940,N_15011,N_15436);
xor U17941 (N_17941,N_16453,N_15903);
nand U17942 (N_17942,N_15652,N_15535);
nor U17943 (N_17943,N_15218,N_15647);
xnor U17944 (N_17944,N_15739,N_16329);
or U17945 (N_17945,N_15449,N_15081);
xnor U17946 (N_17946,N_16178,N_15075);
nand U17947 (N_17947,N_15539,N_15841);
or U17948 (N_17948,N_16435,N_15336);
and U17949 (N_17949,N_15725,N_16385);
or U17950 (N_17950,N_15150,N_16307);
xnor U17951 (N_17951,N_15570,N_15608);
xor U17952 (N_17952,N_15964,N_15404);
nand U17953 (N_17953,N_15445,N_15795);
or U17954 (N_17954,N_15966,N_15180);
nor U17955 (N_17955,N_15455,N_15359);
and U17956 (N_17956,N_15713,N_15324);
and U17957 (N_17957,N_15118,N_15915);
nand U17958 (N_17958,N_15279,N_16355);
and U17959 (N_17959,N_16412,N_15482);
and U17960 (N_17960,N_15170,N_15905);
xnor U17961 (N_17961,N_16460,N_15501);
nor U17962 (N_17962,N_15158,N_16025);
or U17963 (N_17963,N_15521,N_15300);
nor U17964 (N_17964,N_16356,N_16119);
nor U17965 (N_17965,N_15083,N_15570);
or U17966 (N_17966,N_16480,N_16109);
or U17967 (N_17967,N_16070,N_16221);
xnor U17968 (N_17968,N_15550,N_16244);
and U17969 (N_17969,N_16452,N_15326);
or U17970 (N_17970,N_15004,N_15794);
xnor U17971 (N_17971,N_16347,N_15406);
or U17972 (N_17972,N_16009,N_15173);
and U17973 (N_17973,N_16432,N_15831);
xor U17974 (N_17974,N_15006,N_15149);
and U17975 (N_17975,N_16098,N_16291);
or U17976 (N_17976,N_16214,N_16473);
nand U17977 (N_17977,N_15194,N_16362);
or U17978 (N_17978,N_16345,N_15159);
nand U17979 (N_17979,N_16422,N_15079);
nand U17980 (N_17980,N_15060,N_15892);
xnor U17981 (N_17981,N_15740,N_15587);
nor U17982 (N_17982,N_16099,N_16335);
nor U17983 (N_17983,N_15177,N_16029);
nand U17984 (N_17984,N_16070,N_15700);
nand U17985 (N_17985,N_15268,N_15430);
nor U17986 (N_17986,N_15838,N_15761);
nor U17987 (N_17987,N_15909,N_15162);
nor U17988 (N_17988,N_15151,N_15760);
nand U17989 (N_17989,N_16386,N_16445);
or U17990 (N_17990,N_15895,N_15374);
nor U17991 (N_17991,N_15428,N_15331);
and U17992 (N_17992,N_15315,N_15342);
xor U17993 (N_17993,N_15269,N_15913);
and U17994 (N_17994,N_15596,N_15382);
xor U17995 (N_17995,N_15149,N_16163);
or U17996 (N_17996,N_16264,N_16479);
xnor U17997 (N_17997,N_16282,N_15532);
nand U17998 (N_17998,N_15661,N_15868);
or U17999 (N_17999,N_16321,N_15316);
nor U18000 (N_18000,N_17957,N_17832);
nor U18001 (N_18001,N_16732,N_17351);
and U18002 (N_18002,N_17309,N_17479);
nor U18003 (N_18003,N_17138,N_17075);
xor U18004 (N_18004,N_17888,N_16999);
or U18005 (N_18005,N_17781,N_17488);
nand U18006 (N_18006,N_17838,N_17910);
or U18007 (N_18007,N_17719,N_17234);
nor U18008 (N_18008,N_16972,N_16872);
xor U18009 (N_18009,N_16751,N_17690);
and U18010 (N_18010,N_16736,N_17023);
nor U18011 (N_18011,N_17913,N_17988);
xor U18012 (N_18012,N_17874,N_17044);
or U18013 (N_18013,N_17821,N_17318);
nand U18014 (N_18014,N_17501,N_16748);
nor U18015 (N_18015,N_17817,N_16841);
nor U18016 (N_18016,N_17671,N_16975);
or U18017 (N_18017,N_16527,N_17028);
nor U18018 (N_18018,N_16821,N_17416);
and U18019 (N_18019,N_17646,N_16850);
nor U18020 (N_18020,N_16686,N_16608);
and U18021 (N_18021,N_16888,N_17734);
xnor U18022 (N_18022,N_17751,N_16961);
or U18023 (N_18023,N_17836,N_16662);
xnor U18024 (N_18024,N_17993,N_16645);
or U18025 (N_18025,N_16644,N_17964);
nand U18026 (N_18026,N_16853,N_16650);
xor U18027 (N_18027,N_17928,N_17718);
nand U18028 (N_18028,N_16601,N_17389);
nor U18029 (N_18029,N_17731,N_17546);
nor U18030 (N_18030,N_17859,N_17872);
or U18031 (N_18031,N_17325,N_16965);
and U18032 (N_18032,N_16604,N_16772);
xor U18033 (N_18033,N_17217,N_16825);
and U18034 (N_18034,N_17580,N_16523);
nand U18035 (N_18035,N_16613,N_16976);
nor U18036 (N_18036,N_17653,N_17732);
nand U18037 (N_18037,N_17446,N_16913);
and U18038 (N_18038,N_17692,N_17035);
xor U18039 (N_18039,N_17634,N_17638);
nor U18040 (N_18040,N_16820,N_17729);
xnor U18041 (N_18041,N_17244,N_16747);
xor U18042 (N_18042,N_17271,N_17721);
or U18043 (N_18043,N_17557,N_17857);
or U18044 (N_18044,N_17236,N_17068);
and U18045 (N_18045,N_17034,N_17815);
or U18046 (N_18046,N_17001,N_17121);
and U18047 (N_18047,N_17795,N_17551);
or U18048 (N_18048,N_16918,N_17039);
or U18049 (N_18049,N_17435,N_16842);
and U18050 (N_18050,N_17677,N_16861);
or U18051 (N_18051,N_17590,N_16970);
and U18052 (N_18052,N_17357,N_17515);
xor U18053 (N_18053,N_17730,N_17208);
nand U18054 (N_18054,N_17024,N_17885);
or U18055 (N_18055,N_17008,N_17126);
or U18056 (N_18056,N_17490,N_17599);
xor U18057 (N_18057,N_17432,N_17554);
nor U18058 (N_18058,N_17958,N_17015);
nor U18059 (N_18059,N_17969,N_17549);
nor U18060 (N_18060,N_16630,N_17502);
nor U18061 (N_18061,N_17960,N_17425);
and U18062 (N_18062,N_16863,N_17756);
xnor U18063 (N_18063,N_16755,N_17245);
nand U18064 (N_18064,N_17996,N_17214);
or U18065 (N_18065,N_16845,N_16809);
nor U18066 (N_18066,N_17649,N_17179);
or U18067 (N_18067,N_17555,N_17867);
xor U18068 (N_18068,N_17655,N_17892);
and U18069 (N_18069,N_17049,N_16948);
xnor U18070 (N_18070,N_16723,N_16596);
or U18071 (N_18071,N_16540,N_17575);
xor U18072 (N_18072,N_16835,N_17430);
nor U18073 (N_18073,N_17529,N_16974);
and U18074 (N_18074,N_16661,N_16980);
or U18075 (N_18075,N_17429,N_16562);
and U18076 (N_18076,N_16549,N_17084);
or U18077 (N_18077,N_16561,N_17368);
or U18078 (N_18078,N_17322,N_17173);
xor U18079 (N_18079,N_17114,N_17990);
nand U18080 (N_18080,N_17887,N_17582);
and U18081 (N_18081,N_17989,N_17311);
and U18082 (N_18082,N_17469,N_17806);
nand U18083 (N_18083,N_17376,N_16854);
xor U18084 (N_18084,N_17539,N_16810);
nor U18085 (N_18085,N_17705,N_17308);
and U18086 (N_18086,N_16646,N_16683);
and U18087 (N_18087,N_17123,N_16602);
nand U18088 (N_18088,N_17824,N_16622);
and U18089 (N_18089,N_17141,N_16628);
xnor U18090 (N_18090,N_16934,N_17863);
xnor U18091 (N_18091,N_17641,N_17998);
nand U18092 (N_18092,N_17113,N_16735);
and U18093 (N_18093,N_17890,N_17150);
or U18094 (N_18094,N_17019,N_17133);
xnor U18095 (N_18095,N_17940,N_16771);
and U18096 (N_18096,N_16876,N_17080);
nand U18097 (N_18097,N_17424,N_17831);
nand U18098 (N_18098,N_17936,N_16884);
and U18099 (N_18099,N_17697,N_17074);
or U18100 (N_18100,N_16515,N_17828);
nor U18101 (N_18101,N_16826,N_17540);
xnor U18102 (N_18102,N_17603,N_16846);
or U18103 (N_18103,N_17514,N_17346);
xnor U18104 (N_18104,N_16541,N_17253);
nand U18105 (N_18105,N_17541,N_17714);
xnor U18106 (N_18106,N_16758,N_17755);
nor U18107 (N_18107,N_16942,N_17413);
nor U18108 (N_18108,N_17012,N_17746);
nand U18109 (N_18109,N_17449,N_16658);
nor U18110 (N_18110,N_17796,N_17047);
and U18111 (N_18111,N_17902,N_17330);
nor U18112 (N_18112,N_17421,N_17401);
or U18113 (N_18113,N_17427,N_16651);
and U18114 (N_18114,N_16564,N_17343);
and U18115 (N_18115,N_17240,N_17182);
nand U18116 (N_18116,N_17526,N_17196);
or U18117 (N_18117,N_16746,N_17807);
nand U18118 (N_18118,N_16875,N_16859);
nand U18119 (N_18119,N_17199,N_17313);
and U18120 (N_18120,N_17433,N_16839);
or U18121 (N_18121,N_17959,N_17232);
nand U18122 (N_18122,N_16691,N_16706);
and U18123 (N_18123,N_17904,N_17760);
nand U18124 (N_18124,N_17334,N_16804);
and U18125 (N_18125,N_17187,N_17818);
or U18126 (N_18126,N_17263,N_17802);
nand U18127 (N_18127,N_16937,N_17443);
xnor U18128 (N_18128,N_17628,N_17737);
and U18129 (N_18129,N_17862,N_17131);
or U18130 (N_18130,N_17680,N_17278);
nand U18131 (N_18131,N_16763,N_16827);
or U18132 (N_18132,N_17260,N_17743);
xor U18133 (N_18133,N_17060,N_17669);
nor U18134 (N_18134,N_17591,N_17144);
and U18135 (N_18135,N_16895,N_17915);
and U18136 (N_18136,N_17648,N_16855);
nand U18137 (N_18137,N_16538,N_17595);
or U18138 (N_18138,N_17175,N_17406);
nor U18139 (N_18139,N_16674,N_17605);
nor U18140 (N_18140,N_17399,N_17745);
and U18141 (N_18141,N_16881,N_17917);
nor U18142 (N_18142,N_17383,N_16631);
xor U18143 (N_18143,N_16618,N_17508);
nor U18144 (N_18144,N_17335,N_17316);
or U18145 (N_18145,N_17820,N_17953);
xnor U18146 (N_18146,N_16572,N_17883);
nand U18147 (N_18147,N_17209,N_17579);
and U18148 (N_18148,N_17375,N_17854);
or U18149 (N_18149,N_17947,N_16958);
nor U18150 (N_18150,N_16693,N_17945);
nor U18151 (N_18151,N_17477,N_16817);
nand U18152 (N_18152,N_17265,N_16525);
nand U18153 (N_18153,N_16621,N_17623);
xnor U18154 (N_18154,N_16762,N_17492);
or U18155 (N_18155,N_17987,N_17137);
nand U18156 (N_18156,N_16521,N_17762);
nor U18157 (N_18157,N_16998,N_17676);
nand U18158 (N_18158,N_16689,N_16616);
nand U18159 (N_18159,N_17227,N_16950);
xnor U18160 (N_18160,N_16698,N_16520);
or U18161 (N_18161,N_16929,N_17468);
nor U18162 (N_18162,N_17124,N_17530);
and U18163 (N_18163,N_17592,N_16624);
nand U18164 (N_18164,N_17345,N_17444);
nand U18165 (N_18165,N_17774,N_17152);
nor U18166 (N_18166,N_16892,N_16798);
xnor U18167 (N_18167,N_17951,N_17129);
nor U18168 (N_18168,N_16802,N_17307);
xnor U18169 (N_18169,N_17331,N_16848);
nor U18170 (N_18170,N_17544,N_16529);
xnor U18171 (N_18171,N_17125,N_16886);
and U18172 (N_18172,N_16620,N_17533);
xor U18173 (N_18173,N_16641,N_16860);
nand U18174 (N_18174,N_17261,N_17107);
xor U18175 (N_18175,N_17552,N_17564);
xor U18176 (N_18176,N_17610,N_16593);
nand U18177 (N_18177,N_17397,N_17486);
nor U18178 (N_18178,N_17127,N_17464);
xor U18179 (N_18179,N_17087,N_16806);
and U18180 (N_18180,N_17929,N_16777);
and U18181 (N_18181,N_17914,N_17221);
nand U18182 (N_18182,N_16916,N_17574);
nor U18183 (N_18183,N_17809,N_17000);
or U18184 (N_18184,N_17098,N_16738);
or U18185 (N_18185,N_17378,N_17534);
nor U18186 (N_18186,N_17747,N_16780);
or U18187 (N_18187,N_17689,N_16653);
and U18188 (N_18188,N_16774,N_17104);
or U18189 (N_18189,N_17342,N_17411);
and U18190 (N_18190,N_17513,N_17727);
nor U18191 (N_18191,N_17447,N_17556);
nand U18192 (N_18192,N_17215,N_17819);
and U18193 (N_18193,N_17100,N_17506);
and U18194 (N_18194,N_17639,N_17115);
nand U18195 (N_18195,N_17827,N_16941);
and U18196 (N_18196,N_17059,N_16807);
xnor U18197 (N_18197,N_17329,N_17441);
nor U18198 (N_18198,N_17426,N_16752);
nand U18199 (N_18199,N_17640,N_16740);
nor U18200 (N_18200,N_17673,N_17157);
and U18201 (N_18201,N_16640,N_16659);
nand U18202 (N_18202,N_16677,N_17893);
and U18203 (N_18203,N_16627,N_16514);
nand U18204 (N_18204,N_17407,N_17973);
nand U18205 (N_18205,N_16639,N_17725);
nor U18206 (N_18206,N_16589,N_17153);
and U18207 (N_18207,N_16894,N_16784);
xnor U18208 (N_18208,N_17586,N_17102);
nand U18209 (N_18209,N_16675,N_16778);
nor U18210 (N_18210,N_16503,N_17600);
and U18211 (N_18211,N_16742,N_17735);
nor U18212 (N_18212,N_17791,N_16508);
nor U18213 (N_18213,N_17076,N_16957);
and U18214 (N_18214,N_17630,N_17282);
nor U18215 (N_18215,N_16764,N_16552);
and U18216 (N_18216,N_17758,N_17200);
nand U18217 (N_18217,N_16586,N_17460);
or U18218 (N_18218,N_17078,N_17779);
xnor U18219 (N_18219,N_17291,N_17931);
xnor U18220 (N_18220,N_16971,N_17233);
xor U18221 (N_18221,N_16545,N_17195);
nor U18222 (N_18222,N_17920,N_16576);
nand U18223 (N_18223,N_17687,N_17272);
and U18224 (N_18224,N_17298,N_16829);
or U18225 (N_18225,N_17935,N_17470);
or U18226 (N_18226,N_16800,N_17310);
nor U18227 (N_18227,N_16874,N_16714);
and U18228 (N_18228,N_17471,N_17204);
and U18229 (N_18229,N_16547,N_16933);
or U18230 (N_18230,N_17889,N_17674);
nand U18231 (N_18231,N_17986,N_16502);
or U18232 (N_18232,N_16898,N_17884);
or U18233 (N_18233,N_16730,N_16966);
nor U18234 (N_18234,N_17037,N_16963);
xnor U18235 (N_18235,N_17905,N_17877);
nor U18236 (N_18236,N_17520,N_16991);
xnor U18237 (N_18237,N_17467,N_17394);
and U18238 (N_18238,N_16930,N_16687);
or U18239 (N_18239,N_17652,N_17361);
and U18240 (N_18240,N_17328,N_17950);
and U18241 (N_18241,N_17771,N_17417);
and U18242 (N_18242,N_17249,N_17768);
nor U18243 (N_18243,N_17009,N_16907);
and U18244 (N_18244,N_16647,N_17594);
nor U18245 (N_18245,N_17593,N_17943);
nand U18246 (N_18246,N_16581,N_17999);
and U18247 (N_18247,N_16799,N_17786);
or U18248 (N_18248,N_17352,N_17572);
nand U18249 (N_18249,N_17581,N_17903);
nand U18250 (N_18250,N_17116,N_16956);
nand U18251 (N_18251,N_17082,N_17238);
nand U18252 (N_18252,N_17911,N_16781);
xnor U18253 (N_18253,N_16951,N_17493);
xnor U18254 (N_18254,N_17942,N_16978);
and U18255 (N_18255,N_16877,N_17081);
nand U18256 (N_18256,N_17511,N_17901);
or U18257 (N_18257,N_17979,N_17724);
and U18258 (N_18258,N_17487,N_16943);
or U18259 (N_18259,N_17038,N_17485);
nand U18260 (N_18260,N_17553,N_17491);
and U18261 (N_18261,N_17839,N_17625);
nand U18262 (N_18262,N_16773,N_17624);
and U18263 (N_18263,N_17522,N_17212);
and U18264 (N_18264,N_16559,N_16731);
xnor U18265 (N_18265,N_17712,N_16793);
nor U18266 (N_18266,N_17360,N_17171);
nand U18267 (N_18267,N_16532,N_17315);
or U18268 (N_18268,N_17972,N_17358);
nor U18269 (N_18269,N_16588,N_17284);
and U18270 (N_18270,N_16605,N_16657);
nand U18271 (N_18271,N_16759,N_17856);
nand U18272 (N_18272,N_17650,N_17803);
nor U18273 (N_18273,N_17757,N_17454);
or U18274 (N_18274,N_17861,N_17483);
xnor U18275 (N_18275,N_17198,N_17504);
nand U18276 (N_18276,N_17143,N_17845);
and U18277 (N_18277,N_17881,N_17955);
or U18278 (N_18278,N_17275,N_17169);
and U18279 (N_18279,N_17631,N_16928);
and U18280 (N_18280,N_17823,N_17843);
or U18281 (N_18281,N_17805,N_17984);
and U18282 (N_18282,N_17256,N_17231);
and U18283 (N_18283,N_16813,N_17645);
xor U18284 (N_18284,N_16887,N_17063);
and U18285 (N_18285,N_17866,N_17708);
xnor U18286 (N_18286,N_17808,N_17090);
or U18287 (N_18287,N_16896,N_16721);
nand U18288 (N_18288,N_16664,N_17897);
xnor U18289 (N_18289,N_16590,N_17042);
and U18290 (N_18290,N_17543,N_17402);
and U18291 (N_18291,N_17388,N_17926);
nor U18292 (N_18292,N_17612,N_17665);
or U18293 (N_18293,N_17029,N_17036);
nor U18294 (N_18294,N_17395,N_16921);
xnor U18295 (N_18295,N_16739,N_17804);
xor U18296 (N_18296,N_17442,N_17415);
or U18297 (N_18297,N_17844,N_17642);
nand U18298 (N_18298,N_17093,N_17379);
nand U18299 (N_18299,N_17007,N_16932);
nand U18300 (N_18300,N_16680,N_16979);
and U18301 (N_18301,N_17776,N_17602);
nand U18302 (N_18302,N_17025,N_17667);
or U18303 (N_18303,N_17122,N_16917);
nor U18304 (N_18304,N_17053,N_16560);
and U18305 (N_18305,N_17128,N_16579);
nand U18306 (N_18306,N_16858,N_17033);
nand U18307 (N_18307,N_16592,N_16708);
or U18308 (N_18308,N_17283,N_17451);
nand U18309 (N_18309,N_17202,N_17014);
nor U18310 (N_18310,N_16968,N_16612);
xor U18311 (N_18311,N_17419,N_17158);
or U18312 (N_18312,N_17392,N_16695);
or U18313 (N_18313,N_16993,N_17020);
and U18314 (N_18314,N_17868,N_17041);
nand U18315 (N_18315,N_16707,N_17437);
or U18316 (N_18316,N_17583,N_17482);
xor U18317 (N_18317,N_17742,N_17154);
or U18318 (N_18318,N_16871,N_17478);
nand U18319 (N_18319,N_17072,N_17722);
or U18320 (N_18320,N_16851,N_16788);
nand U18321 (N_18321,N_17643,N_16823);
and U18322 (N_18322,N_17016,N_17299);
and U18323 (N_18323,N_17438,N_17149);
and U18324 (N_18324,N_16787,N_16879);
nand U18325 (N_18325,N_17961,N_17302);
or U18326 (N_18326,N_16870,N_16583);
nand U18327 (N_18327,N_16598,N_17934);
nand U18328 (N_18328,N_17830,N_17966);
xor U18329 (N_18329,N_17288,N_16517);
xor U18330 (N_18330,N_17787,N_17405);
nor U18331 (N_18331,N_17627,N_17775);
nor U18332 (N_18332,N_16789,N_17668);
and U18333 (N_18333,N_17633,N_16988);
nor U18334 (N_18334,N_17085,N_16949);
nand U18335 (N_18335,N_17609,N_17290);
and U18336 (N_18336,N_16669,N_16997);
nor U18337 (N_18337,N_17191,N_16803);
nand U18338 (N_18338,N_17258,N_17670);
nor U18339 (N_18339,N_17531,N_17364);
xor U18340 (N_18340,N_17374,N_17925);
nand U18341 (N_18341,N_17851,N_17850);
or U18342 (N_18342,N_17664,N_16811);
nor U18343 (N_18343,N_17369,N_17661);
or U18344 (N_18344,N_17494,N_16619);
xnor U18345 (N_18345,N_17778,N_17281);
or U18346 (N_18346,N_16632,N_17753);
nor U18347 (N_18347,N_17542,N_16544);
xor U18348 (N_18348,N_17414,N_17252);
xnor U18349 (N_18349,N_16911,N_17338);
or U18350 (N_18350,N_17323,N_17382);
nor U18351 (N_18351,N_17611,N_17254);
nor U18352 (N_18352,N_17206,N_16847);
nand U18353 (N_18353,N_17792,N_17472);
xnor U18354 (N_18354,N_17390,N_16500);
and U18355 (N_18355,N_17408,N_16765);
or U18356 (N_18356,N_16571,N_17228);
nand U18357 (N_18357,N_17637,N_17162);
xnor U18358 (N_18358,N_16805,N_17057);
and U18359 (N_18359,N_16709,N_17651);
nor U18360 (N_18360,N_17907,N_17339);
and U18361 (N_18361,N_17597,N_17095);
xor U18362 (N_18362,N_17013,N_16533);
and U18363 (N_18363,N_17880,N_17246);
or U18364 (N_18364,N_16690,N_16548);
or U18365 (N_18365,N_17666,N_17788);
nor U18366 (N_18366,N_16741,N_17793);
nand U18367 (N_18367,N_16724,N_17396);
and U18368 (N_18368,N_17176,N_17816);
nor U18369 (N_18369,N_17678,N_16885);
xor U18370 (N_18370,N_17834,N_17201);
or U18371 (N_18371,N_17073,N_17213);
xnor U18372 (N_18372,N_17837,N_17975);
nand U18373 (N_18373,N_17733,N_17043);
nor U18374 (N_18374,N_17525,N_16554);
xor U18375 (N_18375,N_17944,N_16946);
xor U18376 (N_18376,N_17703,N_17569);
nand U18377 (N_18377,N_17615,N_17250);
nor U18378 (N_18378,N_17151,N_16969);
xnor U18379 (N_18379,N_17174,N_17237);
and U18380 (N_18380,N_17096,N_16745);
and U18381 (N_18381,N_17326,N_17156);
and U18382 (N_18382,N_16577,N_16761);
and U18383 (N_18383,N_17693,N_17381);
nor U18384 (N_18384,N_17045,N_16655);
nor U18385 (N_18385,N_17918,N_16652);
or U18386 (N_18386,N_17848,N_16678);
xor U18387 (N_18387,N_16831,N_17241);
nand U18388 (N_18388,N_17377,N_16582);
nor U18389 (N_18389,N_17118,N_16530);
nand U18390 (N_18390,N_17420,N_16959);
xor U18391 (N_18391,N_17785,N_16866);
nand U18392 (N_18392,N_16909,N_17120);
nand U18393 (N_18393,N_17711,N_17922);
nand U18394 (N_18394,N_17709,N_17462);
xnor U18395 (N_18395,N_17584,N_17279);
xor U18396 (N_18396,N_17371,N_17900);
nor U18397 (N_18397,N_17192,N_17303);
xnor U18398 (N_18398,N_16703,N_17606);
nand U18399 (N_18399,N_17409,N_17235);
nand U18400 (N_18400,N_16716,N_17230);
and U18401 (N_18401,N_17713,N_16717);
nor U18402 (N_18402,N_17939,N_17380);
or U18403 (N_18403,N_17461,N_17225);
xnor U18404 (N_18404,N_17662,N_16995);
and U18405 (N_18405,N_17203,N_17521);
nand U18406 (N_18406,N_17186,N_17262);
and U18407 (N_18407,N_17932,N_16812);
nand U18408 (N_18408,N_17387,N_17882);
and U18409 (N_18409,N_17341,N_17985);
xnor U18410 (N_18410,N_16537,N_16786);
and U18411 (N_18411,N_16656,N_17632);
or U18412 (N_18412,N_17548,N_16947);
xor U18413 (N_18413,N_17287,N_17306);
xnor U18414 (N_18414,N_16603,N_16637);
nand U18415 (N_18415,N_17864,N_16543);
xnor U18416 (N_18416,N_17489,N_17205);
xor U18417 (N_18417,N_16938,N_17536);
or U18418 (N_18418,N_17337,N_17923);
nand U18419 (N_18419,N_16986,N_17780);
and U18420 (N_18420,N_17616,N_17423);
and U18421 (N_18421,N_17978,N_16511);
nor U18422 (N_18422,N_17140,N_17145);
nor U18423 (N_18423,N_17285,N_16828);
or U18424 (N_18424,N_17782,N_16510);
nand U18425 (N_18425,N_17344,N_17749);
nor U18426 (N_18426,N_16779,N_17223);
or U18427 (N_18427,N_17040,N_17058);
and U18428 (N_18428,N_16926,N_17517);
or U18429 (N_18429,N_16939,N_17453);
xnor U18430 (N_18430,N_17190,N_16534);
nor U18431 (N_18431,N_17276,N_17507);
xor U18432 (N_18432,N_16699,N_17992);
nor U18433 (N_18433,N_16996,N_16819);
and U18434 (N_18434,N_16519,N_16833);
nor U18435 (N_18435,N_17112,N_17359);
or U18436 (N_18436,N_16908,N_17974);
xnor U18437 (N_18437,N_16719,N_17794);
or U18438 (N_18438,N_17560,N_16873);
and U18439 (N_18439,N_17067,N_17702);
xnor U18440 (N_18440,N_17784,N_16915);
and U18441 (N_18441,N_17495,N_17142);
xor U18442 (N_18442,N_17117,N_17908);
xnor U18443 (N_18443,N_16862,N_17728);
xor U18444 (N_18444,N_16531,N_16808);
and U18445 (N_18445,N_16750,N_16575);
and U18446 (N_18446,N_17391,N_17064);
or U18447 (N_18447,N_17163,N_16557);
nand U18448 (N_18448,N_17229,N_16518);
xnor U18449 (N_18449,N_17155,N_17826);
and U18450 (N_18450,N_17754,N_16776);
and U18451 (N_18451,N_17320,N_17841);
nand U18452 (N_18452,N_17933,N_16945);
xnor U18453 (N_18453,N_17952,N_17002);
or U18454 (N_18454,N_17962,N_17193);
xnor U18455 (N_18455,N_16610,N_16796);
nor U18456 (N_18456,N_17134,N_17010);
xnor U18457 (N_18457,N_17672,N_17321);
nand U18458 (N_18458,N_17614,N_17340);
xor U18459 (N_18459,N_17032,N_16625);
or U18460 (N_18460,N_17132,N_17535);
or U18461 (N_18461,N_16900,N_17255);
xor U18462 (N_18462,N_17954,N_16615);
and U18463 (N_18463,N_17077,N_17736);
xor U18464 (N_18464,N_16556,N_16600);
nand U18465 (N_18465,N_17436,N_17005);
or U18466 (N_18466,N_16749,N_17403);
xnor U18467 (N_18467,N_17647,N_17739);
nor U18468 (N_18468,N_16766,N_16700);
and U18469 (N_18469,N_17484,N_17620);
and U18470 (N_18470,N_16940,N_16584);
and U18471 (N_18471,N_16922,N_17448);
nor U18472 (N_18472,N_16783,N_17207);
xor U18473 (N_18473,N_17797,N_17617);
xor U18474 (N_18474,N_17519,N_17658);
xor U18475 (N_18475,N_17715,N_17527);
nand U18476 (N_18476,N_17801,N_17108);
nor U18477 (N_18477,N_16635,N_17891);
nor U18478 (N_18478,N_16756,N_16891);
xor U18479 (N_18479,N_17537,N_17938);
and U18480 (N_18480,N_16790,N_17130);
xnor U18481 (N_18481,N_16864,N_17400);
or U18482 (N_18482,N_17937,N_17251);
xor U18483 (N_18483,N_17264,N_17773);
nor U18484 (N_18484,N_16815,N_17219);
or U18485 (N_18485,N_17577,N_17626);
or U18486 (N_18486,N_17516,N_17790);
nand U18487 (N_18487,N_17510,N_17312);
or U18488 (N_18488,N_17066,N_17347);
or U18489 (N_18489,N_16585,N_17300);
or U18490 (N_18490,N_17991,N_16754);
and U18491 (N_18491,N_17295,N_17497);
or U18492 (N_18492,N_17750,N_17598);
or U18493 (N_18493,N_17571,N_17393);
nand U18494 (N_18494,N_17941,N_16672);
or U18495 (N_18495,N_17977,N_16953);
xor U18496 (N_18496,N_16648,N_17286);
nand U18497 (N_18497,N_16818,N_17684);
or U18498 (N_18498,N_17243,N_16878);
and U18499 (N_18499,N_17906,N_17355);
or U18500 (N_18500,N_16507,N_17688);
and U18501 (N_18501,N_17948,N_17601);
xnor U18502 (N_18502,N_17070,N_16501);
xnor U18503 (N_18503,N_17629,N_17685);
nand U18504 (N_18504,N_17356,N_17224);
xnor U18505 (N_18505,N_17052,N_17829);
xor U18506 (N_18506,N_17168,N_17319);
or U18507 (N_18507,N_16516,N_17026);
and U18508 (N_18508,N_16535,N_16743);
nor U18509 (N_18509,N_16775,N_17798);
xnor U18510 (N_18510,N_16967,N_16566);
nand U18511 (N_18511,N_16580,N_17105);
or U18512 (N_18512,N_16712,N_17147);
or U18513 (N_18513,N_17896,N_16768);
nand U18514 (N_18514,N_17588,N_17017);
xnor U18515 (N_18515,N_16713,N_17457);
and U18516 (N_18516,N_16512,N_17842);
nor U18517 (N_18517,N_16832,N_17873);
nand U18518 (N_18518,N_17965,N_17194);
nor U18519 (N_18519,N_17197,N_17744);
or U18520 (N_18520,N_17410,N_17853);
nand U18521 (N_18521,N_16667,N_17607);
nand U18522 (N_18522,N_17297,N_17875);
and U18523 (N_18523,N_16617,N_17135);
nor U18524 (N_18524,N_17148,N_16711);
and U18525 (N_18525,N_16679,N_17267);
or U18526 (N_18526,N_17825,N_17006);
or U18527 (N_18527,N_17568,N_16505);
nand U18528 (N_18528,N_17505,N_17619);
or U18529 (N_18529,N_17898,N_16567);
nor U18530 (N_18530,N_17869,N_16867);
and U18531 (N_18531,N_16983,N_17110);
nand U18532 (N_18532,N_17474,N_17720);
and U18533 (N_18533,N_17604,N_17317);
nand U18534 (N_18534,N_17211,N_17088);
nor U18535 (N_18535,N_17178,N_16914);
nor U18536 (N_18536,N_17563,N_17846);
nand U18537 (N_18537,N_16573,N_17970);
nand U18538 (N_18538,N_17811,N_17459);
nor U18539 (N_18539,N_16654,N_17949);
xor U18540 (N_18540,N_17686,N_16550);
and U18541 (N_18541,N_17277,N_17894);
and U18542 (N_18542,N_17878,N_17289);
nand U18543 (N_18543,N_17398,N_16663);
or U18544 (N_18544,N_16694,N_17086);
nor U18545 (N_18545,N_17353,N_17269);
nand U18546 (N_18546,N_17418,N_16836);
nor U18547 (N_18547,N_17723,N_16705);
nand U18548 (N_18548,N_16982,N_17741);
nand U18549 (N_18549,N_17763,N_17170);
or U18550 (N_18550,N_17119,N_16889);
xnor U18551 (N_18551,N_17681,N_17273);
or U18552 (N_18552,N_16607,N_16558);
nand U18553 (N_18553,N_17550,N_17899);
and U18554 (N_18554,N_16606,N_16944);
nor U18555 (N_18555,N_17912,N_16923);
nor U18556 (N_18556,N_17248,N_16595);
and U18557 (N_18557,N_16671,N_17466);
nand U18558 (N_18558,N_17094,N_17799);
nand U18559 (N_18559,N_17558,N_16767);
nand U18560 (N_18560,N_17473,N_17363);
or U18561 (N_18561,N_17764,N_17847);
nand U18562 (N_18562,N_16513,N_17465);
or U18563 (N_18563,N_17699,N_17635);
or U18564 (N_18564,N_16642,N_16676);
nor U18565 (N_18565,N_17840,N_17759);
xor U18566 (N_18566,N_17567,N_17046);
nand U18567 (N_18567,N_16962,N_16989);
or U18568 (N_18568,N_17663,N_16797);
xor U18569 (N_18569,N_16984,N_16729);
or U18570 (N_18570,N_17404,N_17752);
nor U18571 (N_18571,N_17349,N_16760);
or U18572 (N_18572,N_17089,N_16890);
and U18573 (N_18573,N_17139,N_17852);
nor U18574 (N_18574,N_17305,N_17092);
xnor U18575 (N_18575,N_17679,N_17091);
and U18576 (N_18576,N_17812,N_16955);
or U18577 (N_18577,N_16536,N_17576);
and U18578 (N_18578,N_16734,N_17748);
nand U18579 (N_18579,N_17886,N_16737);
or U18580 (N_18580,N_16629,N_17675);
xor U18581 (N_18581,N_16919,N_17636);
xnor U18582 (N_18582,N_17698,N_17021);
nand U18583 (N_18583,N_17879,N_17570);
nand U18584 (N_18584,N_17716,N_16733);
nand U18585 (N_18585,N_16728,N_16553);
nor U18586 (N_18586,N_17216,N_16726);
and U18587 (N_18587,N_17445,N_17218);
nor U18588 (N_18588,N_17103,N_17280);
or U18589 (N_18589,N_17097,N_17810);
nand U18590 (N_18590,N_17370,N_16634);
nand U18591 (N_18591,N_16936,N_17324);
xnor U18592 (N_18592,N_16574,N_17366);
or U18593 (N_18593,N_16569,N_16504);
and U18594 (N_18594,N_17161,N_17919);
nand U18595 (N_18595,N_16704,N_16960);
nor U18596 (N_18596,N_17769,N_16685);
and U18597 (N_18597,N_17384,N_17858);
or U18598 (N_18598,N_17696,N_16824);
or U18599 (N_18599,N_16869,N_16725);
nor U18600 (N_18600,N_17833,N_17835);
and U18601 (N_18601,N_17498,N_17644);
xor U18602 (N_18602,N_17022,N_17870);
and U18603 (N_18603,N_16843,N_17700);
and U18604 (N_18604,N_17691,N_16792);
and U18605 (N_18605,N_17164,N_16856);
nand U18606 (N_18606,N_17332,N_17695);
nand U18607 (N_18607,N_17587,N_17373);
nand U18608 (N_18608,N_16785,N_16791);
and U18609 (N_18609,N_17585,N_17386);
nand U18610 (N_18610,N_16973,N_16905);
nor U18611 (N_18611,N_17983,N_17440);
nand U18612 (N_18612,N_16865,N_16688);
nand U18613 (N_18613,N_16565,N_16506);
nand U18614 (N_18614,N_17767,N_16660);
nor U18615 (N_18615,N_17220,N_17738);
xor U18616 (N_18616,N_17456,N_16883);
nand U18617 (N_18617,N_17956,N_17971);
nand U18618 (N_18618,N_16684,N_16816);
nand U18619 (N_18619,N_16852,N_17004);
nor U18620 (N_18620,N_16901,N_17524);
nand U18621 (N_18621,N_17480,N_17946);
or U18622 (N_18622,N_17481,N_16857);
nor U18623 (N_18623,N_16643,N_16594);
xor U18624 (N_18624,N_16801,N_16844);
xnor U18625 (N_18625,N_17876,N_16757);
or U18626 (N_18626,N_17622,N_16599);
xnor U18627 (N_18627,N_16591,N_17654);
or U18628 (N_18628,N_16849,N_17659);
or U18629 (N_18629,N_16681,N_16665);
xor U18630 (N_18630,N_17968,N_17512);
xnor U18631 (N_18631,N_16782,N_16990);
or U18632 (N_18632,N_17354,N_16899);
nor U18633 (N_18633,N_17247,N_17963);
and U18634 (N_18634,N_17761,N_17242);
nor U18635 (N_18635,N_17458,N_17509);
and U18636 (N_18636,N_17431,N_16838);
xor U18637 (N_18637,N_17777,N_17270);
nand U18638 (N_18638,N_17657,N_17726);
xor U18639 (N_18639,N_16570,N_17336);
nand U18640 (N_18640,N_17800,N_16673);
xnor U18641 (N_18641,N_17921,N_16985);
nor U18642 (N_18642,N_16954,N_17292);
and U18643 (N_18643,N_17031,N_16904);
and U18644 (N_18644,N_17849,N_16528);
or U18645 (N_18645,N_17916,N_16977);
nand U18646 (N_18646,N_17545,N_16597);
and U18647 (N_18647,N_16701,N_17995);
nor U18648 (N_18648,N_17180,N_17562);
nand U18649 (N_18649,N_17146,N_17997);
nor U18650 (N_18650,N_17189,N_16638);
nor U18651 (N_18651,N_17367,N_17701);
or U18652 (N_18652,N_17565,N_17304);
or U18653 (N_18653,N_17450,N_16546);
nand U18654 (N_18654,N_17532,N_16649);
and U18655 (N_18655,N_17050,N_17766);
or U18656 (N_18656,N_17618,N_17710);
and U18657 (N_18657,N_17365,N_16633);
and U18658 (N_18658,N_17184,N_17621);
nor U18659 (N_18659,N_17268,N_17385);
xor U18660 (N_18660,N_16578,N_17274);
or U18661 (N_18661,N_17559,N_17596);
or U18662 (N_18662,N_17704,N_16668);
and U18663 (N_18663,N_17188,N_17500);
nand U18664 (N_18664,N_16710,N_17578);
xor U18665 (N_18665,N_16834,N_17860);
and U18666 (N_18666,N_17056,N_17071);
and U18667 (N_18667,N_16682,N_16814);
or U18668 (N_18668,N_17109,N_17982);
and U18669 (N_18669,N_17222,N_17160);
nor U18670 (N_18670,N_17296,N_17523);
nor U18671 (N_18671,N_17683,N_17561);
nor U18672 (N_18672,N_17707,N_17475);
nand U18673 (N_18673,N_17257,N_17981);
nor U18674 (N_18674,N_16509,N_16555);
or U18675 (N_18675,N_16840,N_16994);
xor U18676 (N_18676,N_17930,N_17813);
or U18677 (N_18677,N_17476,N_17333);
or U18678 (N_18678,N_16702,N_17172);
or U18679 (N_18679,N_16542,N_17210);
and U18680 (N_18680,N_16964,N_17372);
nor U18681 (N_18681,N_17717,N_17538);
or U18682 (N_18682,N_17682,N_17927);
nor U18683 (N_18683,N_17159,N_17226);
nor U18684 (N_18684,N_17924,N_16539);
or U18685 (N_18685,N_16696,N_16551);
xnor U18686 (N_18686,N_16903,N_16981);
and U18687 (N_18687,N_17967,N_16868);
and U18688 (N_18688,N_16902,N_17499);
nand U18689 (N_18689,N_16626,N_16910);
xor U18690 (N_18690,N_16609,N_16522);
nor U18691 (N_18691,N_17166,N_16636);
or U18692 (N_18692,N_17770,N_17694);
nand U18693 (N_18693,N_16753,N_17177);
or U18694 (N_18694,N_17062,N_16524);
nor U18695 (N_18695,N_16697,N_16666);
xnor U18696 (N_18696,N_17412,N_17167);
nor U18697 (N_18697,N_17239,N_17865);
nand U18698 (N_18698,N_17099,N_17789);
and U18699 (N_18699,N_16722,N_17871);
nand U18700 (N_18700,N_16830,N_17055);
nor U18701 (N_18701,N_16611,N_17706);
nor U18702 (N_18702,N_17660,N_17083);
or U18703 (N_18703,N_17822,N_17065);
nor U18704 (N_18704,N_17327,N_17566);
xnor U18705 (N_18705,N_16920,N_16670);
and U18706 (N_18706,N_17814,N_17185);
or U18707 (N_18707,N_16893,N_16952);
or U18708 (N_18708,N_17428,N_17293);
or U18709 (N_18709,N_16718,N_16720);
nand U18710 (N_18710,N_17048,N_17895);
and U18711 (N_18711,N_16882,N_17314);
and U18712 (N_18712,N_17452,N_17350);
xnor U18713 (N_18713,N_17496,N_17613);
or U18714 (N_18714,N_16924,N_17463);
nor U18715 (N_18715,N_17294,N_16931);
nand U18716 (N_18716,N_17765,N_17054);
nor U18717 (N_18717,N_17079,N_17994);
nor U18718 (N_18718,N_16727,N_16568);
xor U18719 (N_18719,N_16795,N_17980);
nand U18720 (N_18720,N_16992,N_17547);
nor U18721 (N_18721,N_17030,N_16744);
xnor U18722 (N_18722,N_17783,N_17003);
xnor U18723 (N_18723,N_17434,N_17503);
or U18724 (N_18724,N_17051,N_16715);
xnor U18725 (N_18725,N_17181,N_17528);
nand U18726 (N_18726,N_17573,N_17018);
and U18727 (N_18727,N_16925,N_16769);
or U18728 (N_18728,N_17259,N_17165);
or U18729 (N_18729,N_17111,N_17136);
nand U18730 (N_18730,N_17106,N_17909);
nand U18731 (N_18731,N_16770,N_16880);
xnor U18732 (N_18732,N_17362,N_16897);
and U18733 (N_18733,N_16912,N_17740);
and U18734 (N_18734,N_16935,N_17183);
xnor U18735 (N_18735,N_17422,N_17301);
xor U18736 (N_18736,N_17608,N_17266);
xor U18737 (N_18737,N_16794,N_16526);
or U18738 (N_18738,N_17061,N_17772);
xnor U18739 (N_18739,N_17589,N_17011);
and U18740 (N_18740,N_16822,N_17101);
nand U18741 (N_18741,N_16987,N_16927);
and U18742 (N_18742,N_17855,N_17976);
and U18743 (N_18743,N_16906,N_16623);
xnor U18744 (N_18744,N_16563,N_17348);
or U18745 (N_18745,N_16837,N_17069);
or U18746 (N_18746,N_16614,N_17518);
nor U18747 (N_18747,N_17455,N_16587);
nor U18748 (N_18748,N_17439,N_17027);
xor U18749 (N_18749,N_17656,N_16692);
xor U18750 (N_18750,N_17737,N_16961);
or U18751 (N_18751,N_17239,N_16777);
nor U18752 (N_18752,N_17055,N_17050);
nand U18753 (N_18753,N_16605,N_17059);
and U18754 (N_18754,N_17596,N_16991);
and U18755 (N_18755,N_16567,N_17061);
xnor U18756 (N_18756,N_17047,N_17401);
nand U18757 (N_18757,N_16733,N_17534);
nor U18758 (N_18758,N_17817,N_17500);
xor U18759 (N_18759,N_17903,N_17363);
nand U18760 (N_18760,N_17014,N_16552);
and U18761 (N_18761,N_16979,N_17651);
xnor U18762 (N_18762,N_17489,N_17664);
or U18763 (N_18763,N_17233,N_16603);
xnor U18764 (N_18764,N_17563,N_17517);
nand U18765 (N_18765,N_17090,N_16619);
or U18766 (N_18766,N_17651,N_17655);
and U18767 (N_18767,N_17399,N_17588);
or U18768 (N_18768,N_16844,N_17482);
nand U18769 (N_18769,N_17070,N_17119);
and U18770 (N_18770,N_17418,N_17961);
xnor U18771 (N_18771,N_17813,N_17163);
and U18772 (N_18772,N_16841,N_17658);
or U18773 (N_18773,N_17412,N_17710);
or U18774 (N_18774,N_16953,N_17282);
or U18775 (N_18775,N_17056,N_17433);
xnor U18776 (N_18776,N_16521,N_17766);
nand U18777 (N_18777,N_17364,N_16962);
xnor U18778 (N_18778,N_17384,N_17705);
and U18779 (N_18779,N_17288,N_17737);
xnor U18780 (N_18780,N_17275,N_17839);
and U18781 (N_18781,N_16893,N_16848);
xnor U18782 (N_18782,N_17584,N_17727);
or U18783 (N_18783,N_16731,N_17685);
nand U18784 (N_18784,N_17311,N_17979);
or U18785 (N_18785,N_16856,N_17005);
nor U18786 (N_18786,N_17140,N_17734);
nand U18787 (N_18787,N_16692,N_17518);
or U18788 (N_18788,N_17985,N_17698);
xnor U18789 (N_18789,N_17684,N_17539);
xnor U18790 (N_18790,N_16864,N_17014);
or U18791 (N_18791,N_17292,N_17338);
nand U18792 (N_18792,N_17299,N_17178);
or U18793 (N_18793,N_17653,N_17763);
nor U18794 (N_18794,N_17971,N_17751);
and U18795 (N_18795,N_17591,N_16778);
xnor U18796 (N_18796,N_16803,N_17565);
and U18797 (N_18797,N_17915,N_17113);
or U18798 (N_18798,N_16920,N_16694);
and U18799 (N_18799,N_16826,N_17343);
xor U18800 (N_18800,N_17747,N_17999);
xor U18801 (N_18801,N_17182,N_17078);
and U18802 (N_18802,N_17070,N_17010);
or U18803 (N_18803,N_16970,N_17571);
and U18804 (N_18804,N_17738,N_16524);
xnor U18805 (N_18805,N_16784,N_17739);
xnor U18806 (N_18806,N_17688,N_16649);
nand U18807 (N_18807,N_16869,N_16852);
or U18808 (N_18808,N_16634,N_16508);
nand U18809 (N_18809,N_17537,N_16680);
nand U18810 (N_18810,N_16752,N_17396);
nor U18811 (N_18811,N_16814,N_17723);
or U18812 (N_18812,N_17476,N_17854);
nor U18813 (N_18813,N_17424,N_17093);
and U18814 (N_18814,N_16610,N_17780);
xor U18815 (N_18815,N_17116,N_16751);
nor U18816 (N_18816,N_16831,N_17575);
nor U18817 (N_18817,N_17681,N_17859);
and U18818 (N_18818,N_16808,N_17710);
nand U18819 (N_18819,N_17484,N_17603);
and U18820 (N_18820,N_16902,N_17185);
and U18821 (N_18821,N_17215,N_16781);
and U18822 (N_18822,N_17220,N_16949);
nor U18823 (N_18823,N_16597,N_16914);
nor U18824 (N_18824,N_17065,N_17184);
xor U18825 (N_18825,N_17327,N_17545);
nor U18826 (N_18826,N_16588,N_17823);
nor U18827 (N_18827,N_17855,N_17171);
nor U18828 (N_18828,N_16699,N_17750);
and U18829 (N_18829,N_17495,N_17344);
or U18830 (N_18830,N_17244,N_17177);
or U18831 (N_18831,N_16770,N_17605);
xor U18832 (N_18832,N_16738,N_17452);
xnor U18833 (N_18833,N_17099,N_16691);
xnor U18834 (N_18834,N_17625,N_17290);
and U18835 (N_18835,N_17837,N_16557);
nand U18836 (N_18836,N_16911,N_17051);
xnor U18837 (N_18837,N_17973,N_16874);
xor U18838 (N_18838,N_16923,N_17277);
nor U18839 (N_18839,N_17642,N_17914);
nand U18840 (N_18840,N_16573,N_17196);
nor U18841 (N_18841,N_16971,N_17095);
xnor U18842 (N_18842,N_17468,N_17534);
or U18843 (N_18843,N_17796,N_16629);
nand U18844 (N_18844,N_16661,N_17632);
or U18845 (N_18845,N_16884,N_17456);
xor U18846 (N_18846,N_17968,N_17875);
or U18847 (N_18847,N_17391,N_17228);
or U18848 (N_18848,N_17327,N_16895);
xnor U18849 (N_18849,N_17277,N_16582);
nor U18850 (N_18850,N_17608,N_16640);
nor U18851 (N_18851,N_17348,N_17877);
and U18852 (N_18852,N_16745,N_17179);
nor U18853 (N_18853,N_16788,N_16648);
nand U18854 (N_18854,N_17259,N_17322);
or U18855 (N_18855,N_17258,N_16825);
nor U18856 (N_18856,N_16743,N_17581);
nor U18857 (N_18857,N_17839,N_17259);
and U18858 (N_18858,N_16684,N_17676);
nand U18859 (N_18859,N_17278,N_17773);
nor U18860 (N_18860,N_17314,N_16538);
nand U18861 (N_18861,N_16860,N_16624);
xor U18862 (N_18862,N_16845,N_16709);
nand U18863 (N_18863,N_17560,N_16865);
or U18864 (N_18864,N_17181,N_16985);
or U18865 (N_18865,N_16613,N_16769);
xnor U18866 (N_18866,N_17635,N_16707);
and U18867 (N_18867,N_17985,N_17038);
nand U18868 (N_18868,N_17514,N_17767);
xor U18869 (N_18869,N_17523,N_17222);
or U18870 (N_18870,N_17534,N_17441);
and U18871 (N_18871,N_17193,N_17919);
xor U18872 (N_18872,N_17450,N_17211);
nor U18873 (N_18873,N_17783,N_16727);
and U18874 (N_18874,N_17551,N_16832);
nand U18875 (N_18875,N_16704,N_17115);
and U18876 (N_18876,N_16872,N_16965);
nor U18877 (N_18877,N_17440,N_16807);
and U18878 (N_18878,N_17284,N_16890);
and U18879 (N_18879,N_17904,N_17628);
or U18880 (N_18880,N_17082,N_17444);
nor U18881 (N_18881,N_16880,N_17427);
and U18882 (N_18882,N_16723,N_16714);
and U18883 (N_18883,N_16790,N_17258);
nor U18884 (N_18884,N_16902,N_17389);
xor U18885 (N_18885,N_16768,N_17438);
nand U18886 (N_18886,N_17158,N_16578);
nand U18887 (N_18887,N_17969,N_17343);
or U18888 (N_18888,N_16646,N_17326);
and U18889 (N_18889,N_16771,N_17050);
or U18890 (N_18890,N_17258,N_17625);
nand U18891 (N_18891,N_16770,N_17754);
and U18892 (N_18892,N_17375,N_17657);
nand U18893 (N_18893,N_17019,N_16817);
nand U18894 (N_18894,N_16985,N_16671);
and U18895 (N_18895,N_17201,N_16966);
nand U18896 (N_18896,N_17512,N_16852);
and U18897 (N_18897,N_16686,N_16916);
xor U18898 (N_18898,N_16918,N_16839);
nand U18899 (N_18899,N_17185,N_16881);
and U18900 (N_18900,N_16664,N_17041);
nand U18901 (N_18901,N_17056,N_17285);
and U18902 (N_18902,N_16906,N_17784);
and U18903 (N_18903,N_16766,N_17400);
and U18904 (N_18904,N_17136,N_17244);
xor U18905 (N_18905,N_17825,N_17574);
or U18906 (N_18906,N_17843,N_17190);
and U18907 (N_18907,N_17334,N_16543);
xnor U18908 (N_18908,N_17457,N_17223);
nor U18909 (N_18909,N_16767,N_17017);
or U18910 (N_18910,N_16816,N_17300);
nor U18911 (N_18911,N_17411,N_17430);
and U18912 (N_18912,N_17150,N_17576);
and U18913 (N_18913,N_16927,N_16744);
nor U18914 (N_18914,N_16669,N_17722);
or U18915 (N_18915,N_17336,N_17134);
and U18916 (N_18916,N_16901,N_16938);
nor U18917 (N_18917,N_17914,N_16773);
nor U18918 (N_18918,N_16696,N_16704);
xnor U18919 (N_18919,N_16508,N_16613);
xnor U18920 (N_18920,N_16767,N_17247);
nor U18921 (N_18921,N_17819,N_16689);
and U18922 (N_18922,N_16952,N_17376);
or U18923 (N_18923,N_17150,N_17312);
or U18924 (N_18924,N_17041,N_16936);
xor U18925 (N_18925,N_17957,N_17598);
and U18926 (N_18926,N_17893,N_17557);
nand U18927 (N_18927,N_16973,N_17687);
nor U18928 (N_18928,N_16850,N_17993);
or U18929 (N_18929,N_17921,N_17895);
xnor U18930 (N_18930,N_17674,N_16861);
xnor U18931 (N_18931,N_17993,N_17018);
xor U18932 (N_18932,N_17994,N_17000);
xor U18933 (N_18933,N_17093,N_16913);
and U18934 (N_18934,N_17289,N_17049);
or U18935 (N_18935,N_17100,N_16893);
xor U18936 (N_18936,N_16853,N_17309);
nand U18937 (N_18937,N_16996,N_17682);
nor U18938 (N_18938,N_17813,N_17206);
nor U18939 (N_18939,N_16974,N_16763);
nor U18940 (N_18940,N_16641,N_16694);
nor U18941 (N_18941,N_17016,N_17108);
xor U18942 (N_18942,N_17532,N_17153);
and U18943 (N_18943,N_17941,N_17122);
nand U18944 (N_18944,N_16800,N_17220);
nand U18945 (N_18945,N_16539,N_17144);
xor U18946 (N_18946,N_17754,N_17724);
or U18947 (N_18947,N_16804,N_16910);
xnor U18948 (N_18948,N_16696,N_17140);
xnor U18949 (N_18949,N_17788,N_16910);
xor U18950 (N_18950,N_17374,N_17426);
nand U18951 (N_18951,N_17870,N_16708);
nor U18952 (N_18952,N_17071,N_17022);
nand U18953 (N_18953,N_17157,N_16681);
and U18954 (N_18954,N_17047,N_16718);
nand U18955 (N_18955,N_16662,N_16789);
nand U18956 (N_18956,N_17789,N_17162);
xnor U18957 (N_18957,N_17012,N_17061);
or U18958 (N_18958,N_16725,N_16971);
nor U18959 (N_18959,N_16794,N_17236);
nor U18960 (N_18960,N_17876,N_16958);
nor U18961 (N_18961,N_17037,N_16624);
or U18962 (N_18962,N_17429,N_17745);
nand U18963 (N_18963,N_17782,N_17017);
and U18964 (N_18964,N_16948,N_17237);
xor U18965 (N_18965,N_17720,N_17801);
xnor U18966 (N_18966,N_17400,N_17312);
or U18967 (N_18967,N_17755,N_16526);
nand U18968 (N_18968,N_17777,N_17302);
nand U18969 (N_18969,N_16554,N_17536);
nand U18970 (N_18970,N_17697,N_17813);
nand U18971 (N_18971,N_16519,N_17394);
nor U18972 (N_18972,N_17529,N_17822);
nand U18973 (N_18973,N_17945,N_17985);
nor U18974 (N_18974,N_17614,N_17693);
and U18975 (N_18975,N_16667,N_17921);
nand U18976 (N_18976,N_17791,N_16671);
nor U18977 (N_18977,N_17621,N_17173);
nor U18978 (N_18978,N_17703,N_17114);
and U18979 (N_18979,N_17808,N_17924);
and U18980 (N_18980,N_17440,N_17051);
or U18981 (N_18981,N_17764,N_17801);
or U18982 (N_18982,N_16807,N_16540);
nand U18983 (N_18983,N_17098,N_17224);
nand U18984 (N_18984,N_16754,N_17257);
and U18985 (N_18985,N_17918,N_17347);
xor U18986 (N_18986,N_17462,N_16699);
nor U18987 (N_18987,N_17745,N_17772);
xnor U18988 (N_18988,N_16838,N_17477);
nand U18989 (N_18989,N_16794,N_17398);
nor U18990 (N_18990,N_17667,N_16622);
and U18991 (N_18991,N_16679,N_17084);
nand U18992 (N_18992,N_17584,N_17902);
or U18993 (N_18993,N_17379,N_17301);
and U18994 (N_18994,N_16590,N_17064);
xnor U18995 (N_18995,N_16915,N_16835);
nor U18996 (N_18996,N_17189,N_16791);
or U18997 (N_18997,N_17892,N_16637);
xor U18998 (N_18998,N_17181,N_17491);
and U18999 (N_18999,N_17565,N_17231);
nand U19000 (N_19000,N_17513,N_17050);
nor U19001 (N_19001,N_17713,N_17153);
nor U19002 (N_19002,N_17912,N_16570);
nor U19003 (N_19003,N_17969,N_16673);
nor U19004 (N_19004,N_17169,N_17707);
xnor U19005 (N_19005,N_17254,N_17564);
or U19006 (N_19006,N_17632,N_17217);
nor U19007 (N_19007,N_17152,N_17530);
and U19008 (N_19008,N_17477,N_17840);
nor U19009 (N_19009,N_16987,N_16513);
xor U19010 (N_19010,N_16853,N_17916);
or U19011 (N_19011,N_17470,N_17608);
nor U19012 (N_19012,N_17318,N_17942);
xnor U19013 (N_19013,N_17836,N_16934);
or U19014 (N_19014,N_17429,N_16814);
nand U19015 (N_19015,N_17667,N_17547);
xor U19016 (N_19016,N_17159,N_17844);
xor U19017 (N_19017,N_17049,N_17113);
xor U19018 (N_19018,N_17555,N_17110);
xor U19019 (N_19019,N_17207,N_16665);
or U19020 (N_19020,N_17771,N_17327);
xor U19021 (N_19021,N_17422,N_16864);
nor U19022 (N_19022,N_16551,N_17075);
and U19023 (N_19023,N_17495,N_17989);
xor U19024 (N_19024,N_16852,N_17717);
and U19025 (N_19025,N_16507,N_17570);
nand U19026 (N_19026,N_17298,N_17285);
and U19027 (N_19027,N_17638,N_17360);
and U19028 (N_19028,N_17270,N_17778);
nor U19029 (N_19029,N_17369,N_17343);
nor U19030 (N_19030,N_17250,N_16545);
nand U19031 (N_19031,N_16915,N_16712);
and U19032 (N_19032,N_16845,N_16521);
nor U19033 (N_19033,N_17703,N_17676);
nor U19034 (N_19034,N_17460,N_17058);
and U19035 (N_19035,N_17890,N_17397);
nand U19036 (N_19036,N_17959,N_17836);
or U19037 (N_19037,N_17245,N_17754);
or U19038 (N_19038,N_17182,N_17405);
and U19039 (N_19039,N_16858,N_16823);
nor U19040 (N_19040,N_17419,N_17130);
nand U19041 (N_19041,N_17422,N_16724);
xor U19042 (N_19042,N_16839,N_17909);
or U19043 (N_19043,N_17814,N_16557);
xor U19044 (N_19044,N_16890,N_16501);
or U19045 (N_19045,N_16864,N_17649);
nor U19046 (N_19046,N_16552,N_16821);
nand U19047 (N_19047,N_17021,N_17287);
and U19048 (N_19048,N_16713,N_17739);
nand U19049 (N_19049,N_17638,N_16948);
and U19050 (N_19050,N_17044,N_17459);
or U19051 (N_19051,N_17006,N_17958);
or U19052 (N_19052,N_17767,N_16640);
and U19053 (N_19053,N_17242,N_17215);
nand U19054 (N_19054,N_17662,N_17987);
xnor U19055 (N_19055,N_16750,N_17721);
nor U19056 (N_19056,N_16867,N_16684);
xnor U19057 (N_19057,N_17800,N_17790);
xor U19058 (N_19058,N_17650,N_17822);
or U19059 (N_19059,N_17543,N_16938);
xor U19060 (N_19060,N_17413,N_17033);
and U19061 (N_19061,N_17690,N_16645);
and U19062 (N_19062,N_17798,N_17036);
and U19063 (N_19063,N_17341,N_16791);
xnor U19064 (N_19064,N_17410,N_17782);
xor U19065 (N_19065,N_17520,N_16865);
nand U19066 (N_19066,N_17623,N_17978);
nor U19067 (N_19067,N_16604,N_17053);
or U19068 (N_19068,N_17919,N_16780);
or U19069 (N_19069,N_17893,N_16623);
xnor U19070 (N_19070,N_17153,N_16897);
nand U19071 (N_19071,N_16794,N_16599);
or U19072 (N_19072,N_17659,N_17637);
and U19073 (N_19073,N_16601,N_16649);
or U19074 (N_19074,N_16724,N_17441);
nor U19075 (N_19075,N_16698,N_16979);
xor U19076 (N_19076,N_17909,N_16891);
and U19077 (N_19077,N_17261,N_16856);
nor U19078 (N_19078,N_17927,N_17475);
nor U19079 (N_19079,N_17657,N_16751);
nand U19080 (N_19080,N_16831,N_16997);
nor U19081 (N_19081,N_17091,N_17913);
xnor U19082 (N_19082,N_17740,N_17898);
and U19083 (N_19083,N_17868,N_17226);
nand U19084 (N_19084,N_17521,N_17107);
and U19085 (N_19085,N_17065,N_17438);
and U19086 (N_19086,N_17599,N_17538);
xor U19087 (N_19087,N_17716,N_16994);
nand U19088 (N_19088,N_17269,N_17542);
xnor U19089 (N_19089,N_17670,N_17402);
nor U19090 (N_19090,N_17576,N_17204);
xnor U19091 (N_19091,N_17753,N_17972);
or U19092 (N_19092,N_17833,N_17700);
nand U19093 (N_19093,N_17737,N_17257);
nand U19094 (N_19094,N_17086,N_16903);
nand U19095 (N_19095,N_17502,N_17997);
and U19096 (N_19096,N_16711,N_17474);
nand U19097 (N_19097,N_17871,N_17237);
nand U19098 (N_19098,N_16818,N_17598);
and U19099 (N_19099,N_16868,N_17962);
and U19100 (N_19100,N_16843,N_16520);
or U19101 (N_19101,N_16873,N_17013);
or U19102 (N_19102,N_17085,N_17667);
nor U19103 (N_19103,N_16693,N_17870);
xnor U19104 (N_19104,N_16554,N_17992);
xnor U19105 (N_19105,N_17688,N_17286);
or U19106 (N_19106,N_17161,N_16795);
and U19107 (N_19107,N_16771,N_17844);
or U19108 (N_19108,N_17820,N_16855);
and U19109 (N_19109,N_17049,N_17349);
or U19110 (N_19110,N_17925,N_16755);
nand U19111 (N_19111,N_16853,N_17186);
nand U19112 (N_19112,N_16580,N_16768);
xor U19113 (N_19113,N_16511,N_16798);
or U19114 (N_19114,N_17409,N_17604);
nor U19115 (N_19115,N_17100,N_17001);
nand U19116 (N_19116,N_16646,N_17117);
nand U19117 (N_19117,N_16667,N_16661);
and U19118 (N_19118,N_17218,N_16901);
or U19119 (N_19119,N_17979,N_17629);
nand U19120 (N_19120,N_17580,N_16540);
xor U19121 (N_19121,N_17474,N_16512);
nand U19122 (N_19122,N_17035,N_16698);
xor U19123 (N_19123,N_17872,N_17807);
and U19124 (N_19124,N_16993,N_17861);
xnor U19125 (N_19125,N_17142,N_17120);
or U19126 (N_19126,N_16933,N_16749);
nand U19127 (N_19127,N_17986,N_16895);
xor U19128 (N_19128,N_16895,N_17391);
and U19129 (N_19129,N_17263,N_17514);
and U19130 (N_19130,N_17492,N_17003);
nand U19131 (N_19131,N_16779,N_16735);
or U19132 (N_19132,N_17763,N_17299);
or U19133 (N_19133,N_17312,N_16931);
and U19134 (N_19134,N_17808,N_17869);
or U19135 (N_19135,N_17912,N_16926);
and U19136 (N_19136,N_16627,N_17042);
nor U19137 (N_19137,N_17277,N_17646);
nor U19138 (N_19138,N_16826,N_17172);
and U19139 (N_19139,N_17105,N_16715);
nor U19140 (N_19140,N_17087,N_16964);
or U19141 (N_19141,N_16577,N_17394);
nand U19142 (N_19142,N_16603,N_16975);
and U19143 (N_19143,N_17603,N_16909);
nor U19144 (N_19144,N_16694,N_17953);
and U19145 (N_19145,N_16676,N_17257);
nand U19146 (N_19146,N_17436,N_16685);
or U19147 (N_19147,N_17169,N_17769);
and U19148 (N_19148,N_17274,N_16913);
or U19149 (N_19149,N_16785,N_17285);
xnor U19150 (N_19150,N_17757,N_16578);
nor U19151 (N_19151,N_17687,N_17351);
or U19152 (N_19152,N_17332,N_17194);
nor U19153 (N_19153,N_17520,N_16810);
and U19154 (N_19154,N_17876,N_17224);
and U19155 (N_19155,N_17734,N_17655);
and U19156 (N_19156,N_17303,N_16547);
and U19157 (N_19157,N_17548,N_17781);
nand U19158 (N_19158,N_16583,N_17912);
and U19159 (N_19159,N_17146,N_17138);
nor U19160 (N_19160,N_16779,N_17506);
and U19161 (N_19161,N_17760,N_16880);
or U19162 (N_19162,N_16713,N_17598);
nor U19163 (N_19163,N_16698,N_16906);
nor U19164 (N_19164,N_17141,N_17526);
nor U19165 (N_19165,N_17561,N_17485);
and U19166 (N_19166,N_17499,N_17915);
nand U19167 (N_19167,N_17419,N_17241);
or U19168 (N_19168,N_16866,N_17510);
nor U19169 (N_19169,N_17604,N_16650);
and U19170 (N_19170,N_16871,N_17611);
and U19171 (N_19171,N_16881,N_16656);
xnor U19172 (N_19172,N_17090,N_17593);
nand U19173 (N_19173,N_17069,N_17861);
xnor U19174 (N_19174,N_16579,N_17347);
xor U19175 (N_19175,N_17031,N_16727);
or U19176 (N_19176,N_16950,N_16602);
nor U19177 (N_19177,N_17495,N_17406);
and U19178 (N_19178,N_17679,N_16687);
or U19179 (N_19179,N_17141,N_17917);
nor U19180 (N_19180,N_17345,N_16926);
and U19181 (N_19181,N_16845,N_17448);
or U19182 (N_19182,N_16572,N_17016);
nand U19183 (N_19183,N_17737,N_16857);
nor U19184 (N_19184,N_17509,N_17786);
xnor U19185 (N_19185,N_17437,N_17393);
xor U19186 (N_19186,N_17225,N_16786);
and U19187 (N_19187,N_17077,N_16643);
nand U19188 (N_19188,N_17295,N_17270);
nor U19189 (N_19189,N_17517,N_17742);
xor U19190 (N_19190,N_17043,N_16767);
nor U19191 (N_19191,N_17923,N_17987);
and U19192 (N_19192,N_17075,N_17469);
xnor U19193 (N_19193,N_17725,N_17030);
and U19194 (N_19194,N_17533,N_16783);
xor U19195 (N_19195,N_17952,N_17644);
or U19196 (N_19196,N_17492,N_17277);
or U19197 (N_19197,N_17210,N_17265);
nand U19198 (N_19198,N_16595,N_16899);
nand U19199 (N_19199,N_17031,N_17332);
xnor U19200 (N_19200,N_16784,N_17774);
nand U19201 (N_19201,N_17851,N_16694);
nor U19202 (N_19202,N_17561,N_17729);
xnor U19203 (N_19203,N_17971,N_17472);
nand U19204 (N_19204,N_16888,N_16784);
or U19205 (N_19205,N_17072,N_16999);
and U19206 (N_19206,N_17535,N_17954);
nand U19207 (N_19207,N_16578,N_16603);
or U19208 (N_19208,N_17171,N_16599);
or U19209 (N_19209,N_16779,N_16865);
nor U19210 (N_19210,N_17992,N_17847);
nor U19211 (N_19211,N_17068,N_17237);
xor U19212 (N_19212,N_16680,N_16936);
nand U19213 (N_19213,N_16939,N_17846);
nor U19214 (N_19214,N_17389,N_16874);
nor U19215 (N_19215,N_17994,N_17680);
and U19216 (N_19216,N_17721,N_17647);
nor U19217 (N_19217,N_17352,N_16762);
or U19218 (N_19218,N_17842,N_17600);
or U19219 (N_19219,N_17842,N_17712);
or U19220 (N_19220,N_17926,N_16666);
nor U19221 (N_19221,N_16568,N_16596);
or U19222 (N_19222,N_17448,N_17394);
nor U19223 (N_19223,N_17933,N_17838);
and U19224 (N_19224,N_16562,N_17654);
nor U19225 (N_19225,N_17685,N_17588);
xor U19226 (N_19226,N_16851,N_16930);
nor U19227 (N_19227,N_16743,N_16610);
xor U19228 (N_19228,N_17862,N_17948);
and U19229 (N_19229,N_17417,N_16989);
xnor U19230 (N_19230,N_17468,N_16743);
nor U19231 (N_19231,N_17841,N_17243);
nor U19232 (N_19232,N_17522,N_17217);
and U19233 (N_19233,N_17900,N_16991);
and U19234 (N_19234,N_17715,N_16548);
nand U19235 (N_19235,N_16658,N_16586);
nand U19236 (N_19236,N_17848,N_17716);
and U19237 (N_19237,N_17394,N_16822);
or U19238 (N_19238,N_16535,N_17017);
and U19239 (N_19239,N_16847,N_17430);
nor U19240 (N_19240,N_17693,N_17364);
and U19241 (N_19241,N_17138,N_17148);
nand U19242 (N_19242,N_16586,N_16635);
and U19243 (N_19243,N_17991,N_16777);
nor U19244 (N_19244,N_17507,N_17469);
or U19245 (N_19245,N_16723,N_17841);
or U19246 (N_19246,N_16627,N_17682);
or U19247 (N_19247,N_17351,N_17101);
nor U19248 (N_19248,N_16893,N_17933);
or U19249 (N_19249,N_17498,N_16546);
xor U19250 (N_19250,N_17141,N_17597);
or U19251 (N_19251,N_17586,N_17573);
nor U19252 (N_19252,N_17743,N_17483);
nand U19253 (N_19253,N_17293,N_16996);
xor U19254 (N_19254,N_17335,N_16641);
nor U19255 (N_19255,N_17028,N_16568);
or U19256 (N_19256,N_17944,N_16954);
xor U19257 (N_19257,N_17720,N_16514);
xnor U19258 (N_19258,N_17235,N_17280);
and U19259 (N_19259,N_16591,N_16918);
and U19260 (N_19260,N_17021,N_17609);
nor U19261 (N_19261,N_17840,N_17829);
or U19262 (N_19262,N_17055,N_17339);
nand U19263 (N_19263,N_17858,N_16805);
nor U19264 (N_19264,N_17202,N_16820);
or U19265 (N_19265,N_17074,N_17189);
and U19266 (N_19266,N_17452,N_16839);
nand U19267 (N_19267,N_17838,N_16777);
and U19268 (N_19268,N_16853,N_17957);
or U19269 (N_19269,N_17921,N_17164);
and U19270 (N_19270,N_16522,N_17415);
nor U19271 (N_19271,N_16879,N_17528);
and U19272 (N_19272,N_16620,N_17625);
xnor U19273 (N_19273,N_17044,N_16594);
and U19274 (N_19274,N_16937,N_16543);
and U19275 (N_19275,N_17196,N_17868);
or U19276 (N_19276,N_17111,N_17613);
and U19277 (N_19277,N_17687,N_16878);
nor U19278 (N_19278,N_17118,N_16916);
or U19279 (N_19279,N_16867,N_17492);
nor U19280 (N_19280,N_17632,N_16967);
and U19281 (N_19281,N_16962,N_17148);
nor U19282 (N_19282,N_16541,N_17344);
nor U19283 (N_19283,N_16985,N_17186);
nor U19284 (N_19284,N_17072,N_16678);
and U19285 (N_19285,N_17964,N_17091);
or U19286 (N_19286,N_17454,N_16771);
xor U19287 (N_19287,N_17501,N_17632);
and U19288 (N_19288,N_17736,N_16523);
xnor U19289 (N_19289,N_16503,N_17569);
nor U19290 (N_19290,N_17181,N_17539);
xnor U19291 (N_19291,N_17401,N_17221);
xnor U19292 (N_19292,N_17363,N_17072);
and U19293 (N_19293,N_17832,N_17005);
xnor U19294 (N_19294,N_16929,N_17093);
and U19295 (N_19295,N_16761,N_16671);
xor U19296 (N_19296,N_17339,N_17815);
xor U19297 (N_19297,N_17634,N_17156);
xor U19298 (N_19298,N_17756,N_17740);
or U19299 (N_19299,N_17245,N_16607);
and U19300 (N_19300,N_17176,N_17350);
or U19301 (N_19301,N_17567,N_16685);
and U19302 (N_19302,N_16661,N_17822);
and U19303 (N_19303,N_17935,N_17898);
nor U19304 (N_19304,N_16607,N_17309);
and U19305 (N_19305,N_16890,N_17942);
nor U19306 (N_19306,N_16626,N_17244);
nor U19307 (N_19307,N_17726,N_16626);
or U19308 (N_19308,N_17030,N_16818);
xor U19309 (N_19309,N_17645,N_17768);
nand U19310 (N_19310,N_16973,N_17292);
xnor U19311 (N_19311,N_17189,N_17323);
nor U19312 (N_19312,N_16599,N_17850);
nor U19313 (N_19313,N_17460,N_17503);
or U19314 (N_19314,N_17994,N_17653);
and U19315 (N_19315,N_17097,N_17656);
nor U19316 (N_19316,N_17712,N_17674);
nand U19317 (N_19317,N_17090,N_17963);
and U19318 (N_19318,N_16815,N_17059);
nand U19319 (N_19319,N_17345,N_17600);
and U19320 (N_19320,N_17475,N_17885);
nand U19321 (N_19321,N_17129,N_17376);
and U19322 (N_19322,N_17903,N_17897);
xor U19323 (N_19323,N_17937,N_16540);
or U19324 (N_19324,N_16582,N_16626);
or U19325 (N_19325,N_17292,N_17369);
and U19326 (N_19326,N_16665,N_17171);
or U19327 (N_19327,N_17958,N_16663);
or U19328 (N_19328,N_17742,N_17222);
xnor U19329 (N_19329,N_17964,N_17026);
xor U19330 (N_19330,N_17023,N_17185);
and U19331 (N_19331,N_17082,N_16725);
nor U19332 (N_19332,N_17699,N_17488);
xor U19333 (N_19333,N_16745,N_16765);
nor U19334 (N_19334,N_17770,N_16808);
or U19335 (N_19335,N_17264,N_16731);
nand U19336 (N_19336,N_17778,N_16968);
or U19337 (N_19337,N_17887,N_17850);
or U19338 (N_19338,N_16831,N_16658);
and U19339 (N_19339,N_17863,N_16512);
or U19340 (N_19340,N_16514,N_17159);
xnor U19341 (N_19341,N_16944,N_16776);
nand U19342 (N_19342,N_16914,N_17997);
nand U19343 (N_19343,N_16835,N_17814);
or U19344 (N_19344,N_17071,N_17656);
nand U19345 (N_19345,N_16544,N_17675);
xnor U19346 (N_19346,N_17878,N_17972);
xnor U19347 (N_19347,N_16694,N_17615);
xnor U19348 (N_19348,N_17923,N_16779);
nand U19349 (N_19349,N_17723,N_16917);
nand U19350 (N_19350,N_17652,N_17440);
xor U19351 (N_19351,N_16636,N_16789);
or U19352 (N_19352,N_17717,N_17381);
or U19353 (N_19353,N_17284,N_17402);
xnor U19354 (N_19354,N_16674,N_17604);
and U19355 (N_19355,N_17314,N_17431);
nor U19356 (N_19356,N_17626,N_17970);
xnor U19357 (N_19357,N_17938,N_17035);
and U19358 (N_19358,N_17229,N_17729);
or U19359 (N_19359,N_17367,N_17713);
nor U19360 (N_19360,N_17783,N_17593);
and U19361 (N_19361,N_16766,N_17353);
or U19362 (N_19362,N_17162,N_17198);
xor U19363 (N_19363,N_17721,N_17523);
nor U19364 (N_19364,N_17521,N_17767);
and U19365 (N_19365,N_17581,N_17123);
xnor U19366 (N_19366,N_17218,N_17487);
or U19367 (N_19367,N_17184,N_17677);
nor U19368 (N_19368,N_17597,N_16912);
and U19369 (N_19369,N_17631,N_17179);
and U19370 (N_19370,N_17982,N_17009);
xor U19371 (N_19371,N_16692,N_16673);
and U19372 (N_19372,N_16624,N_16877);
nand U19373 (N_19373,N_17137,N_17067);
and U19374 (N_19374,N_16634,N_17170);
nand U19375 (N_19375,N_17782,N_17992);
or U19376 (N_19376,N_16833,N_16944);
or U19377 (N_19377,N_17755,N_16842);
nand U19378 (N_19378,N_16881,N_17407);
and U19379 (N_19379,N_17420,N_17201);
xnor U19380 (N_19380,N_17860,N_17796);
nor U19381 (N_19381,N_16911,N_17663);
xor U19382 (N_19382,N_16973,N_17503);
or U19383 (N_19383,N_16640,N_17993);
nor U19384 (N_19384,N_16551,N_17842);
nand U19385 (N_19385,N_16769,N_17387);
nand U19386 (N_19386,N_17192,N_16655);
nand U19387 (N_19387,N_17904,N_17590);
nand U19388 (N_19388,N_17893,N_17039);
nand U19389 (N_19389,N_17617,N_16792);
or U19390 (N_19390,N_16956,N_17891);
xnor U19391 (N_19391,N_17712,N_16706);
or U19392 (N_19392,N_16878,N_16660);
xnor U19393 (N_19393,N_17105,N_17773);
nand U19394 (N_19394,N_17628,N_17874);
and U19395 (N_19395,N_16634,N_17735);
and U19396 (N_19396,N_17711,N_16877);
or U19397 (N_19397,N_16514,N_17005);
and U19398 (N_19398,N_17265,N_17394);
nand U19399 (N_19399,N_17483,N_16639);
nand U19400 (N_19400,N_17349,N_16879);
nor U19401 (N_19401,N_17616,N_16869);
xnor U19402 (N_19402,N_17086,N_17080);
nor U19403 (N_19403,N_16739,N_17014);
and U19404 (N_19404,N_16997,N_16828);
xor U19405 (N_19405,N_17202,N_17669);
xor U19406 (N_19406,N_17727,N_17593);
xnor U19407 (N_19407,N_16886,N_17305);
nor U19408 (N_19408,N_16684,N_17819);
xnor U19409 (N_19409,N_17758,N_17372);
or U19410 (N_19410,N_17593,N_17105);
or U19411 (N_19411,N_16603,N_16687);
nor U19412 (N_19412,N_17175,N_17311);
xnor U19413 (N_19413,N_17287,N_17046);
or U19414 (N_19414,N_16554,N_17991);
and U19415 (N_19415,N_17105,N_17024);
or U19416 (N_19416,N_16712,N_16957);
nor U19417 (N_19417,N_17381,N_17149);
and U19418 (N_19418,N_17006,N_16941);
and U19419 (N_19419,N_16903,N_17277);
or U19420 (N_19420,N_17194,N_17588);
nor U19421 (N_19421,N_17621,N_17806);
nor U19422 (N_19422,N_17578,N_16744);
nand U19423 (N_19423,N_16852,N_17767);
or U19424 (N_19424,N_17232,N_16944);
and U19425 (N_19425,N_16688,N_16698);
and U19426 (N_19426,N_17481,N_17189);
nand U19427 (N_19427,N_16926,N_16801);
nor U19428 (N_19428,N_17092,N_17012);
nand U19429 (N_19429,N_17784,N_17822);
and U19430 (N_19430,N_17982,N_16551);
nor U19431 (N_19431,N_17478,N_17991);
nand U19432 (N_19432,N_17304,N_17470);
or U19433 (N_19433,N_17402,N_16910);
and U19434 (N_19434,N_16805,N_17954);
nand U19435 (N_19435,N_17224,N_17039);
or U19436 (N_19436,N_17249,N_17181);
or U19437 (N_19437,N_16878,N_16998);
and U19438 (N_19438,N_17167,N_16788);
nand U19439 (N_19439,N_16975,N_16973);
nor U19440 (N_19440,N_17237,N_17950);
xnor U19441 (N_19441,N_17144,N_17024);
or U19442 (N_19442,N_17264,N_17045);
nand U19443 (N_19443,N_16888,N_16577);
nor U19444 (N_19444,N_16569,N_17776);
or U19445 (N_19445,N_16591,N_17933);
and U19446 (N_19446,N_16665,N_17699);
and U19447 (N_19447,N_16852,N_17206);
or U19448 (N_19448,N_16919,N_16570);
xnor U19449 (N_19449,N_16885,N_17329);
nor U19450 (N_19450,N_17717,N_17337);
and U19451 (N_19451,N_17080,N_17962);
and U19452 (N_19452,N_16957,N_16803);
xnor U19453 (N_19453,N_17159,N_16583);
nor U19454 (N_19454,N_17388,N_17396);
or U19455 (N_19455,N_17479,N_17695);
xor U19456 (N_19456,N_17506,N_16593);
nand U19457 (N_19457,N_17921,N_16626);
and U19458 (N_19458,N_17725,N_16697);
and U19459 (N_19459,N_16882,N_17207);
or U19460 (N_19460,N_17573,N_16945);
nand U19461 (N_19461,N_16797,N_17625);
nor U19462 (N_19462,N_17649,N_17264);
nand U19463 (N_19463,N_16742,N_17047);
xnor U19464 (N_19464,N_17293,N_17623);
or U19465 (N_19465,N_16573,N_17840);
nor U19466 (N_19466,N_17959,N_16878);
nor U19467 (N_19467,N_17167,N_16882);
xor U19468 (N_19468,N_17943,N_17296);
and U19469 (N_19469,N_17603,N_16966);
or U19470 (N_19470,N_17790,N_17826);
xnor U19471 (N_19471,N_17514,N_17670);
or U19472 (N_19472,N_17346,N_17772);
xor U19473 (N_19473,N_17136,N_17127);
or U19474 (N_19474,N_17111,N_17560);
xor U19475 (N_19475,N_17090,N_17096);
and U19476 (N_19476,N_17086,N_16723);
nand U19477 (N_19477,N_17551,N_17399);
xor U19478 (N_19478,N_17978,N_16527);
nand U19479 (N_19479,N_16699,N_17740);
or U19480 (N_19480,N_16727,N_17982);
and U19481 (N_19481,N_17460,N_17475);
and U19482 (N_19482,N_17697,N_17909);
or U19483 (N_19483,N_17766,N_17368);
or U19484 (N_19484,N_16928,N_17182);
and U19485 (N_19485,N_17609,N_16630);
nor U19486 (N_19486,N_17178,N_17398);
nand U19487 (N_19487,N_17704,N_17792);
or U19488 (N_19488,N_17454,N_16608);
nor U19489 (N_19489,N_17941,N_17343);
nand U19490 (N_19490,N_17116,N_17219);
or U19491 (N_19491,N_16737,N_16702);
xor U19492 (N_19492,N_16592,N_17955);
xnor U19493 (N_19493,N_17250,N_17277);
nor U19494 (N_19494,N_17180,N_17565);
or U19495 (N_19495,N_16995,N_17750);
nor U19496 (N_19496,N_17689,N_16991);
or U19497 (N_19497,N_17080,N_16602);
nor U19498 (N_19498,N_16703,N_16574);
and U19499 (N_19499,N_16674,N_17865);
or U19500 (N_19500,N_18269,N_18307);
and U19501 (N_19501,N_18022,N_18171);
nor U19502 (N_19502,N_18557,N_18305);
nand U19503 (N_19503,N_18961,N_19341);
and U19504 (N_19504,N_18430,N_18152);
or U19505 (N_19505,N_18830,N_19101);
nand U19506 (N_19506,N_19215,N_18038);
xnor U19507 (N_19507,N_18742,N_18591);
and U19508 (N_19508,N_18309,N_18739);
and U19509 (N_19509,N_19053,N_18151);
and U19510 (N_19510,N_18319,N_19096);
nor U19511 (N_19511,N_18174,N_19130);
xnor U19512 (N_19512,N_19041,N_18988);
and U19513 (N_19513,N_18561,N_19131);
xnor U19514 (N_19514,N_18857,N_18869);
xnor U19515 (N_19515,N_18413,N_19342);
nor U19516 (N_19516,N_18956,N_19435);
and U19517 (N_19517,N_19234,N_18111);
nor U19518 (N_19518,N_18280,N_18959);
and U19519 (N_19519,N_18429,N_18075);
and U19520 (N_19520,N_18207,N_18998);
xor U19521 (N_19521,N_19492,N_18406);
xnor U19522 (N_19522,N_19357,N_19111);
xor U19523 (N_19523,N_19316,N_18975);
or U19524 (N_19524,N_18662,N_18006);
xnor U19525 (N_19525,N_19244,N_18925);
xor U19526 (N_19526,N_18908,N_18845);
xor U19527 (N_19527,N_18437,N_18537);
nor U19528 (N_19528,N_19441,N_18829);
or U19529 (N_19529,N_18923,N_18387);
nor U19530 (N_19530,N_19179,N_18167);
or U19531 (N_19531,N_18905,N_18405);
nor U19532 (N_19532,N_18364,N_18861);
and U19533 (N_19533,N_18211,N_19248);
nand U19534 (N_19534,N_18454,N_18196);
xnor U19535 (N_19535,N_18618,N_18545);
xnor U19536 (N_19536,N_19344,N_18617);
or U19537 (N_19537,N_18994,N_18805);
nand U19538 (N_19538,N_19254,N_19010);
or U19539 (N_19539,N_18021,N_18627);
and U19540 (N_19540,N_19323,N_18051);
xor U19541 (N_19541,N_18997,N_18121);
and U19542 (N_19542,N_19263,N_18137);
or U19543 (N_19543,N_18297,N_18717);
or U19544 (N_19544,N_18189,N_18225);
or U19545 (N_19545,N_18809,N_19166);
and U19546 (N_19546,N_18817,N_18026);
and U19547 (N_19547,N_18448,N_18042);
or U19548 (N_19548,N_18694,N_18090);
or U19549 (N_19549,N_18820,N_19337);
nor U19550 (N_19550,N_18741,N_18419);
xnor U19551 (N_19551,N_18782,N_18621);
or U19552 (N_19552,N_18835,N_19436);
and U19553 (N_19553,N_18578,N_18093);
nand U19554 (N_19554,N_19196,N_19207);
xor U19555 (N_19555,N_19392,N_18025);
nor U19556 (N_19556,N_18163,N_18446);
and U19557 (N_19557,N_19233,N_18145);
or U19558 (N_19558,N_18815,N_19093);
and U19559 (N_19559,N_19307,N_18254);
xor U19560 (N_19560,N_19035,N_18453);
or U19561 (N_19561,N_19083,N_19349);
nand U19562 (N_19562,N_19330,N_18227);
xnor U19563 (N_19563,N_18023,N_19170);
and U19564 (N_19564,N_18910,N_18142);
nand U19565 (N_19565,N_19328,N_18015);
nor U19566 (N_19566,N_18941,N_18543);
nand U19567 (N_19567,N_18053,N_18938);
nand U19568 (N_19568,N_18549,N_18973);
and U19569 (N_19569,N_18004,N_19048);
xnor U19570 (N_19570,N_19407,N_19222);
nand U19571 (N_19571,N_18314,N_18032);
nor U19572 (N_19572,N_19438,N_19168);
nor U19573 (N_19573,N_19102,N_19421);
xnor U19574 (N_19574,N_19277,N_19326);
and U19575 (N_19575,N_19183,N_19311);
and U19576 (N_19576,N_18170,N_19125);
nor U19577 (N_19577,N_18426,N_18002);
xnor U19578 (N_19578,N_19430,N_18718);
nor U19579 (N_19579,N_18271,N_19391);
nand U19580 (N_19580,N_18791,N_18298);
xor U19581 (N_19581,N_18416,N_19081);
nand U19582 (N_19582,N_18386,N_19003);
or U19583 (N_19583,N_19494,N_19006);
nand U19584 (N_19584,N_19481,N_18186);
nor U19585 (N_19585,N_18489,N_18045);
xor U19586 (N_19586,N_18204,N_19106);
or U19587 (N_19587,N_18728,N_19230);
and U19588 (N_19588,N_18456,N_19008);
nor U19589 (N_19589,N_19015,N_18408);
nor U19590 (N_19590,N_18572,N_18885);
xor U19591 (N_19591,N_18834,N_19406);
nor U19592 (N_19592,N_18256,N_19158);
nor U19593 (N_19593,N_19178,N_19180);
xor U19594 (N_19594,N_18631,N_18864);
or U19595 (N_19595,N_19389,N_18881);
and U19596 (N_19596,N_18306,N_18899);
or U19597 (N_19597,N_19442,N_18643);
or U19598 (N_19598,N_18232,N_18176);
or U19599 (N_19599,N_18380,N_19173);
and U19600 (N_19600,N_18206,N_19029);
and U19601 (N_19601,N_19383,N_19470);
nand U19602 (N_19602,N_19126,N_19068);
xor U19603 (N_19603,N_18262,N_18969);
nor U19604 (N_19604,N_19428,N_18982);
nor U19605 (N_19605,N_18190,N_18548);
xor U19606 (N_19606,N_19270,N_19043);
and U19607 (N_19607,N_18073,N_18619);
and U19608 (N_19608,N_18625,N_18596);
and U19609 (N_19609,N_18526,N_19051);
nor U19610 (N_19610,N_18913,N_19187);
nor U19611 (N_19611,N_18036,N_18381);
or U19612 (N_19612,N_19107,N_18503);
xor U19613 (N_19613,N_18699,N_18246);
xnor U19614 (N_19614,N_18274,N_18930);
nand U19615 (N_19615,N_19221,N_19459);
nand U19616 (N_19616,N_18601,N_18346);
and U19617 (N_19617,N_18390,N_19191);
or U19618 (N_19618,N_18629,N_18005);
nor U19619 (N_19619,N_18392,N_18642);
and U19620 (N_19620,N_18275,N_19242);
or U19621 (N_19621,N_18035,N_18593);
and U19622 (N_19622,N_18100,N_19335);
and U19623 (N_19623,N_19352,N_18794);
nand U19624 (N_19624,N_18674,N_19315);
xor U19625 (N_19625,N_19231,N_18415);
xnor U19626 (N_19626,N_19240,N_18808);
and U19627 (N_19627,N_18219,N_18579);
or U19628 (N_19628,N_19305,N_18746);
and U19629 (N_19629,N_19480,N_18872);
and U19630 (N_19630,N_18963,N_18332);
nand U19631 (N_19631,N_18356,N_18081);
or U19632 (N_19632,N_18821,N_18716);
or U19633 (N_19633,N_19278,N_19448);
nor U19634 (N_19634,N_18584,N_18187);
and U19635 (N_19635,N_18486,N_18544);
and U19636 (N_19636,N_19265,N_19299);
nor U19637 (N_19637,N_18721,N_18528);
nand U19638 (N_19638,N_18607,N_18551);
nor U19639 (N_19639,N_18731,N_18926);
xor U19640 (N_19640,N_18842,N_18072);
and U19641 (N_19641,N_19033,N_18276);
or U19642 (N_19642,N_18412,N_18838);
nor U19643 (N_19643,N_18865,N_18304);
xor U19644 (N_19644,N_19232,N_19202);
or U19645 (N_19645,N_19446,N_18825);
and U19646 (N_19646,N_19151,N_18116);
or U19647 (N_19647,N_19425,N_19289);
nand U19648 (N_19648,N_18921,N_18811);
nand U19649 (N_19649,N_18554,N_18962);
and U19650 (N_19650,N_18637,N_18542);
or U19651 (N_19651,N_18311,N_19269);
or U19652 (N_19652,N_19264,N_19274);
or U19653 (N_19653,N_18494,N_18535);
and U19654 (N_19654,N_18786,N_18466);
or U19655 (N_19655,N_18303,N_18009);
or U19656 (N_19656,N_19312,N_18434);
or U19657 (N_19657,N_19325,N_19137);
nor U19658 (N_19658,N_19149,N_19487);
or U19659 (N_19659,N_19467,N_18553);
nor U19660 (N_19660,N_18239,N_18340);
nand U19661 (N_19661,N_18198,N_19171);
or U19662 (N_19662,N_18576,N_18059);
and U19663 (N_19663,N_18652,N_18933);
or U19664 (N_19664,N_19078,N_18368);
xnor U19665 (N_19665,N_18457,N_19287);
or U19666 (N_19666,N_18952,N_18730);
xnor U19667 (N_19667,N_18855,N_18449);
nor U19668 (N_19668,N_18780,N_18282);
or U19669 (N_19669,N_18079,N_18411);
nand U19670 (N_19670,N_18039,N_18148);
nor U19671 (N_19671,N_18562,N_19123);
and U19672 (N_19672,N_18240,N_19057);
or U19673 (N_19673,N_18495,N_18477);
or U19674 (N_19674,N_19229,N_19482);
xor U19675 (N_19675,N_18020,N_19455);
and U19676 (N_19676,N_18164,N_18610);
nand U19677 (N_19677,N_18669,N_19141);
or U19678 (N_19678,N_18402,N_18445);
xor U19679 (N_19679,N_19145,N_19022);
xor U19680 (N_19680,N_19030,N_19476);
nor U19681 (N_19681,N_19372,N_19243);
nor U19682 (N_19682,N_19351,N_19063);
and U19683 (N_19683,N_18673,N_18900);
nand U19684 (N_19684,N_19212,N_18441);
and U19685 (N_19685,N_18894,N_18365);
nor U19686 (N_19686,N_18832,N_18192);
nand U19687 (N_19687,N_18439,N_18612);
or U19688 (N_19688,N_18658,N_18342);
xor U19689 (N_19689,N_18224,N_18614);
xnor U19690 (N_19690,N_18824,N_18028);
or U19691 (N_19691,N_18278,N_19012);
nand U19692 (N_19692,N_19408,N_18783);
and U19693 (N_19693,N_18985,N_19009);
nand U19694 (N_19694,N_19100,N_19115);
nor U19695 (N_19695,N_19380,N_18810);
or U19696 (N_19696,N_18770,N_18713);
xor U19697 (N_19697,N_18889,N_18491);
and U19698 (N_19698,N_18436,N_18632);
xnor U19699 (N_19699,N_19154,N_19127);
or U19700 (N_19700,N_18143,N_18487);
or U19701 (N_19701,N_19143,N_18054);
and U19702 (N_19702,N_18481,N_18972);
and U19703 (N_19703,N_19318,N_18818);
xor U19704 (N_19704,N_19452,N_18118);
and U19705 (N_19705,N_18657,N_19339);
nand U19706 (N_19706,N_18907,N_18775);
or U19707 (N_19707,N_18223,N_18539);
xnor U19708 (N_19708,N_18604,N_18213);
or U19709 (N_19709,N_19049,N_18928);
and U19710 (N_19710,N_18740,N_18571);
xor U19711 (N_19711,N_19276,N_18338);
and U19712 (N_19712,N_18299,N_18797);
and U19713 (N_19713,N_19086,N_18476);
or U19714 (N_19714,N_19472,N_19427);
or U19715 (N_19715,N_19150,N_19386);
nor U19716 (N_19716,N_19350,N_19366);
nor U19717 (N_19717,N_19493,N_18635);
nor U19718 (N_19718,N_19024,N_19275);
nor U19719 (N_19719,N_18606,N_18114);
or U19720 (N_19720,N_19479,N_18709);
and U19721 (N_19721,N_18049,N_18144);
xnor U19722 (N_19722,N_18229,N_19090);
and U19723 (N_19723,N_18464,N_19114);
or U19724 (N_19724,N_18147,N_18315);
or U19725 (N_19725,N_19046,N_18279);
nand U19726 (N_19726,N_18991,N_18744);
nand U19727 (N_19727,N_18678,N_19411);
nor U19728 (N_19728,N_18257,N_18689);
nor U19729 (N_19729,N_18550,N_18083);
nor U19730 (N_19730,N_18914,N_18541);
xnor U19731 (N_19731,N_19238,N_18388);
nor U19732 (N_19732,N_19272,N_19044);
nor U19733 (N_19733,N_18410,N_18609);
xor U19734 (N_19734,N_19110,N_18583);
nand U19735 (N_19735,N_19412,N_19120);
nand U19736 (N_19736,N_19450,N_18498);
xnor U19737 (N_19737,N_19443,N_18769);
and U19738 (N_19738,N_18839,N_18261);
and U19739 (N_19739,N_19290,N_19208);
or U19740 (N_19740,N_19317,N_18670);
xnor U19741 (N_19741,N_18676,N_19279);
and U19742 (N_19742,N_18724,N_18605);
or U19743 (N_19743,N_18097,N_18953);
and U19744 (N_19744,N_19061,N_19437);
or U19745 (N_19745,N_18816,N_18955);
nor U19746 (N_19746,N_18360,N_19060);
nor U19747 (N_19747,N_19065,N_19292);
or U19748 (N_19748,N_19136,N_18029);
nor U19749 (N_19749,N_18250,N_19266);
and U19750 (N_19750,N_18628,N_19175);
nor U19751 (N_19751,N_18706,N_19226);
or U19752 (N_19752,N_18397,N_18667);
nor U19753 (N_19753,N_18697,N_18455);
nand U19754 (N_19754,N_18329,N_18870);
nand U19755 (N_19755,N_19302,N_18231);
and U19756 (N_19756,N_19416,N_19458);
xor U19757 (N_19757,N_18895,N_19117);
or U19758 (N_19758,N_18420,N_19034);
or U19759 (N_19759,N_18107,N_19308);
or U19760 (N_19760,N_18650,N_18203);
xnor U19761 (N_19761,N_19332,N_18715);
or U19762 (N_19762,N_18520,N_18277);
or U19763 (N_19763,N_19002,N_18241);
nand U19764 (N_19764,N_18559,N_18761);
and U19765 (N_19765,N_19192,N_18385);
or U19766 (N_19766,N_19082,N_18695);
nand U19767 (N_19767,N_19108,N_19201);
nor U19768 (N_19768,N_18105,N_19354);
nor U19769 (N_19769,N_19236,N_18680);
xor U19770 (N_19770,N_18751,N_19210);
nor U19771 (N_19771,N_18874,N_18892);
or U19772 (N_19772,N_19485,N_18488);
nor U19773 (N_19773,N_18949,N_18126);
and U19774 (N_19774,N_18611,N_18139);
and U19775 (N_19775,N_18951,N_18055);
and U19776 (N_19776,N_18210,N_18932);
nand U19777 (N_19777,N_18555,N_18787);
xnor U19778 (N_19778,N_18316,N_18513);
or U19779 (N_19779,N_19146,N_19403);
nor U19780 (N_19780,N_18616,N_18188);
or U19781 (N_19781,N_19404,N_18837);
nand U19782 (N_19782,N_18301,N_19422);
and U19783 (N_19783,N_18504,N_18878);
nand U19784 (N_19784,N_18506,N_18518);
or U19785 (N_19785,N_18654,N_19410);
nor U19786 (N_19786,N_18812,N_18165);
nor U19787 (N_19787,N_18876,N_18463);
nand U19788 (N_19788,N_18313,N_19356);
nand U19789 (N_19789,N_18123,N_19050);
xor U19790 (N_19790,N_19249,N_18157);
xnor U19791 (N_19791,N_18376,N_18472);
nor U19792 (N_19792,N_18078,N_19301);
xor U19793 (N_19793,N_18714,N_18964);
or U19794 (N_19794,N_18336,N_18600);
nor U19795 (N_19795,N_19075,N_18681);
and U19796 (N_19796,N_18031,N_19495);
xor U19797 (N_19797,N_18580,N_18971);
or U19798 (N_19798,N_18101,N_18597);
and U19799 (N_19799,N_19205,N_18841);
xor U19800 (N_19800,N_18321,N_18266);
xor U19801 (N_19801,N_19097,N_19016);
xor U19802 (N_19802,N_18379,N_18359);
or U19803 (N_19803,N_18208,N_18814);
xor U19804 (N_19804,N_18685,N_18369);
xnor U19805 (N_19805,N_19295,N_18218);
xnor U19806 (N_19806,N_18427,N_18019);
or U19807 (N_19807,N_18756,N_18570);
nor U19808 (N_19808,N_18175,N_18996);
or U19809 (N_19809,N_19280,N_19135);
nand U19810 (N_19810,N_18801,N_18008);
nand U19811 (N_19811,N_18462,N_18317);
xnor U19812 (N_19812,N_19214,N_18088);
nand U19813 (N_19813,N_18183,N_18840);
xnor U19814 (N_19814,N_19071,N_18538);
nor U19815 (N_19815,N_18660,N_18484);
and U19816 (N_19816,N_19098,N_19070);
xnor U19817 (N_19817,N_18155,N_18358);
nand U19818 (N_19818,N_18470,N_18394);
nand U19819 (N_19819,N_18409,N_18194);
nand U19820 (N_19820,N_18981,N_18846);
xnor U19821 (N_19821,N_18113,N_18773);
or U19822 (N_19822,N_18659,N_19461);
and U19823 (N_19823,N_18747,N_18977);
and U19824 (N_19824,N_18060,N_18902);
nand U19825 (N_19825,N_18771,N_18065);
or U19826 (N_19826,N_18950,N_18260);
and U19827 (N_19827,N_18140,N_18592);
xor U19828 (N_19828,N_18112,N_18016);
or U19829 (N_19829,N_19094,N_18636);
and U19830 (N_19830,N_19257,N_19095);
nand U19831 (N_19831,N_18851,N_19076);
and U19832 (N_19832,N_19159,N_18873);
or U19833 (N_19833,N_18182,N_19285);
nor U19834 (N_19834,N_18912,N_19304);
nor U19835 (N_19835,N_18327,N_19157);
nor U19836 (N_19836,N_18033,N_18896);
xor U19837 (N_19837,N_18201,N_19224);
xnor U19838 (N_19838,N_19400,N_18736);
nand U19839 (N_19839,N_18626,N_18337);
and U19840 (N_19840,N_19011,N_19398);
nand U19841 (N_19841,N_18354,N_19186);
nand U19842 (N_19842,N_19155,N_19142);
and U19843 (N_19843,N_18258,N_19334);
or U19844 (N_19844,N_18440,N_18124);
or U19845 (N_19845,N_19319,N_19447);
or U19846 (N_19846,N_19054,N_18334);
and U19847 (N_19847,N_18987,N_18682);
and U19848 (N_19848,N_19468,N_19119);
nor U19849 (N_19849,N_18954,N_18252);
and U19850 (N_19850,N_18759,N_19080);
xor U19851 (N_19851,N_18451,N_18483);
nor U19852 (N_19852,N_18687,N_18285);
nand U19853 (N_19853,N_19194,N_19466);
nor U19854 (N_19854,N_19160,N_18178);
or U19855 (N_19855,N_19184,N_18357);
nand U19856 (N_19856,N_18712,N_18935);
nand U19857 (N_19857,N_18490,N_18986);
nor U19858 (N_19858,N_18173,N_18345);
nand U19859 (N_19859,N_18141,N_19105);
or U19860 (N_19860,N_19377,N_19206);
nor U19861 (N_19861,N_18447,N_18668);
xor U19862 (N_19862,N_18048,N_18244);
xor U19863 (N_19863,N_18853,N_18395);
or U19864 (N_19864,N_18980,N_18711);
nand U19865 (N_19865,N_18265,N_18983);
xor U19866 (N_19866,N_18161,N_19491);
or U19867 (N_19867,N_18150,N_18527);
nand U19868 (N_19868,N_18819,N_19027);
nand U19869 (N_19869,N_19069,N_19116);
nand U19870 (N_19870,N_19169,N_19134);
nand U19871 (N_19871,N_19031,N_18071);
nor U19872 (N_19872,N_18799,N_18286);
and U19873 (N_19873,N_18887,N_18943);
nor U19874 (N_19874,N_18577,N_18245);
and U19875 (N_19875,N_19219,N_19445);
and U19876 (N_19876,N_18735,N_18478);
and U19877 (N_19877,N_18407,N_18209);
nor U19878 (N_19878,N_18960,N_18401);
and U19879 (N_19879,N_18293,N_18339);
nor U19880 (N_19880,N_19132,N_19394);
xnor U19881 (N_19881,N_18967,N_18757);
nand U19882 (N_19882,N_18166,N_19393);
nor U19883 (N_19883,N_18560,N_18723);
and U19884 (N_19884,N_18129,N_18804);
nand U19885 (N_19885,N_18001,N_18509);
nor U19886 (N_19886,N_18867,N_18133);
nor U19887 (N_19887,N_19294,N_19381);
and U19888 (N_19888,N_18061,N_18017);
nand U19889 (N_19889,N_18848,N_18574);
and U19890 (N_19890,N_18566,N_18130);
nand U19891 (N_19891,N_19129,N_18034);
and U19892 (N_19892,N_18993,N_18267);
and U19893 (N_19893,N_19293,N_18177);
xnor U19894 (N_19894,N_18469,N_18523);
xnor U19895 (N_19895,N_18431,N_18911);
nor U19896 (N_19896,N_18037,N_18595);
nor U19897 (N_19897,N_19471,N_18929);
nand U19898 (N_19898,N_18940,N_19163);
and U19899 (N_19899,N_19037,N_18511);
nor U19900 (N_19900,N_19498,N_18886);
nor U19901 (N_19901,N_18904,N_18665);
nor U19902 (N_19902,N_19322,N_18671);
or U19903 (N_19903,N_18202,N_18630);
nor U19904 (N_19904,N_18435,N_19310);
nand U19905 (N_19905,N_19478,N_18355);
and U19906 (N_19906,N_18199,N_19434);
and U19907 (N_19907,N_18027,N_19036);
nor U19908 (N_19908,N_18375,N_18086);
and U19909 (N_19909,N_19193,N_18418);
nand U19910 (N_19910,N_18999,N_19052);
or U19911 (N_19911,N_18110,N_19138);
xnor U19912 (N_19912,N_18168,N_18888);
or U19913 (N_19913,N_18132,N_18362);
nand U19914 (N_19914,N_19042,N_18529);
and U19915 (N_19915,N_19088,N_19039);
nor U19916 (N_19916,N_18030,N_18270);
or U19917 (N_19917,N_18608,N_19217);
nor U19918 (N_19918,N_18014,N_18692);
and U19919 (N_19919,N_19079,N_19162);
nand U19920 (N_19920,N_18496,N_19488);
xnor U19921 (N_19921,N_18575,N_19040);
and U19922 (N_19922,N_19113,N_19415);
or U19923 (N_19923,N_19001,N_18403);
xnor U19924 (N_19924,N_18095,N_18531);
xnor U19925 (N_19925,N_19432,N_19139);
and U19926 (N_19926,N_19195,N_18802);
or U19927 (N_19927,N_18957,N_18517);
nor U19928 (N_19928,N_18581,N_18222);
xnor U19929 (N_19929,N_19228,N_18745);
nand U19930 (N_19930,N_18871,N_18701);
and U19931 (N_19931,N_18565,N_18798);
nand U19932 (N_19932,N_18589,N_18762);
and U19933 (N_19933,N_18158,N_18564);
or U19934 (N_19934,N_19329,N_18655);
or U19935 (N_19935,N_18916,N_18844);
or U19936 (N_19936,N_19396,N_18287);
and U19937 (N_19937,N_19260,N_18727);
xnor U19938 (N_19938,N_18281,N_18686);
and U19939 (N_19939,N_18530,N_19144);
nor U19940 (N_19940,N_19298,N_18363);
nor U19941 (N_19941,N_18263,N_19176);
or U19942 (N_19942,N_18793,N_18558);
nand U19943 (N_19943,N_18302,N_19190);
or U19944 (N_19944,N_18942,N_18080);
xnor U19945 (N_19945,N_18289,N_19204);
nand U19946 (N_19946,N_18349,N_19062);
nor U19947 (N_19947,N_18897,N_18467);
or U19948 (N_19948,N_18640,N_18353);
nand U19949 (N_19949,N_18138,N_18044);
xor U19950 (N_19950,N_18854,N_18777);
xnor U19951 (N_19951,N_18508,N_19433);
xor U19952 (N_19952,N_19172,N_18587);
xor U19953 (N_19953,N_19247,N_18465);
nand U19954 (N_19954,N_18880,N_18594);
nor U19955 (N_19955,N_18312,N_18989);
nor U19956 (N_19956,N_18965,N_18522);
or U19957 (N_19957,N_19387,N_19359);
or U19958 (N_19958,N_18092,N_18047);
or U19959 (N_19959,N_18296,N_18428);
nand U19960 (N_19960,N_18656,N_18396);
or U19961 (N_19961,N_19005,N_18862);
and U19962 (N_19962,N_19309,N_18146);
xor U19963 (N_19963,N_18990,N_19336);
and U19964 (N_19964,N_18253,N_18471);
or U19965 (N_19965,N_18290,N_19087);
nor U19966 (N_19966,N_18233,N_18195);
or U19967 (N_19967,N_19331,N_19104);
or U19968 (N_19968,N_18502,N_18666);
or U19969 (N_19969,N_18404,N_18807);
or U19970 (N_19970,N_18242,N_18131);
and U19971 (N_19971,N_19368,N_18255);
nand U19972 (N_19972,N_18691,N_18300);
xor U19973 (N_19973,N_19072,N_18806);
nand U19974 (N_19974,N_18688,N_18729);
or U19975 (N_19975,N_19378,N_18333);
or U19976 (N_19976,N_18647,N_18292);
nor U19977 (N_19977,N_18639,N_18507);
and U19978 (N_19978,N_18458,N_18373);
and U19979 (N_19979,N_19121,N_18310);
nand U19980 (N_19980,N_19283,N_19321);
and U19981 (N_19981,N_18970,N_18512);
and U19982 (N_19982,N_19382,N_19475);
and U19983 (N_19983,N_18623,N_19379);
nand U19984 (N_19984,N_18228,N_18939);
or U19985 (N_19985,N_18737,N_18398);
nor U19986 (N_19986,N_18251,N_18119);
nor U19987 (N_19987,N_18370,N_18534);
nor U19988 (N_19988,N_19313,N_18108);
nor U19989 (N_19989,N_18700,N_18624);
xor U19990 (N_19990,N_18103,N_19007);
and U19991 (N_19991,N_19147,N_19397);
nand U19992 (N_19992,N_19038,N_18444);
nor U19993 (N_19993,N_18516,N_19182);
nor U19994 (N_19994,N_18524,N_18785);
or U19995 (N_19995,N_19419,N_19128);
and U19996 (N_19996,N_19164,N_18567);
and U19997 (N_19997,N_19227,N_19089);
nand U19998 (N_19998,N_18879,N_19250);
and U19999 (N_19999,N_18084,N_18831);
xor U20000 (N_20000,N_18226,N_19401);
xnor U20001 (N_20001,N_19338,N_19497);
nand U20002 (N_20002,N_18180,N_18294);
and U20003 (N_20003,N_18000,N_18361);
xor U20004 (N_20004,N_18236,N_18698);
or U20005 (N_20005,N_18937,N_18089);
nand U20006 (N_20006,N_19241,N_19066);
or U20007 (N_20007,N_18500,N_19140);
or U20008 (N_20008,N_19369,N_19281);
nand U20009 (N_20009,N_19374,N_18927);
nor U20010 (N_20010,N_18085,N_18077);
or U20011 (N_20011,N_18115,N_18181);
nor U20012 (N_20012,N_18767,N_19025);
and U20013 (N_20013,N_18012,N_18796);
and U20014 (N_20014,N_19109,N_18273);
xor U20015 (N_20015,N_18536,N_18040);
or U20016 (N_20016,N_18109,N_18324);
nor U20017 (N_20017,N_18371,N_18391);
nor U20018 (N_20018,N_18399,N_18764);
xor U20019 (N_20019,N_18283,N_18013);
or U20020 (N_20020,N_18850,N_19363);
xnor U20021 (N_20021,N_18521,N_19439);
and U20022 (N_20022,N_19343,N_19177);
or U20023 (N_20023,N_18732,N_19477);
nor U20024 (N_20024,N_18320,N_18979);
nand U20025 (N_20025,N_18160,N_19073);
and U20026 (N_20026,N_19327,N_19246);
or U20027 (N_20027,N_19203,N_19286);
and U20028 (N_20028,N_19440,N_18863);
or U20029 (N_20029,N_18169,N_19490);
nand U20030 (N_20030,N_18615,N_18884);
or U20031 (N_20031,N_19463,N_18215);
and U20032 (N_20032,N_19340,N_19303);
or U20033 (N_20033,N_18127,N_18351);
nor U20034 (N_20034,N_18122,N_19362);
or U20035 (N_20035,N_19103,N_18172);
and U20036 (N_20036,N_18421,N_18069);
nor U20037 (N_20037,N_18046,N_19099);
and U20038 (N_20038,N_18052,N_18098);
nor U20039 (N_20039,N_19324,N_18460);
or U20040 (N_20040,N_18847,N_18284);
nand U20041 (N_20041,N_18193,N_19499);
or U20042 (N_20042,N_18585,N_18719);
nand U20043 (N_20043,N_19085,N_18752);
nor U20044 (N_20044,N_18883,N_18331);
or U20045 (N_20045,N_19174,N_19414);
nand U20046 (N_20046,N_19355,N_18212);
or U20047 (N_20047,N_19489,N_18622);
nand U20048 (N_20048,N_18992,N_19431);
and U20049 (N_20049,N_19261,N_18828);
nor U20050 (N_20050,N_18947,N_18099);
xor U20051 (N_20051,N_18546,N_18672);
nor U20052 (N_20052,N_18134,N_18344);
xnor U20053 (N_20053,N_19161,N_19032);
and U20054 (N_20054,N_18318,N_19465);
xnor U20055 (N_20055,N_18779,N_18859);
xor U20056 (N_20056,N_18238,N_18058);
nor U20057 (N_20057,N_18753,N_19273);
nor U20058 (N_20058,N_18322,N_18492);
nor U20059 (N_20059,N_18803,N_18683);
or U20060 (N_20060,N_18573,N_18649);
nand U20061 (N_20061,N_18149,N_18868);
nand U20062 (N_20062,N_19019,N_19454);
or U20063 (N_20063,N_18734,N_19122);
nand U20064 (N_20064,N_18645,N_18915);
or U20065 (N_20065,N_19297,N_18184);
or U20066 (N_20066,N_18249,N_18563);
xnor U20067 (N_20067,N_19358,N_18547);
and U20068 (N_20068,N_18159,N_18323);
or U20069 (N_20069,N_18860,N_18205);
nor U20070 (N_20070,N_18350,N_19112);
xnor U20071 (N_20071,N_18795,N_18919);
nand U20072 (N_20072,N_18823,N_18056);
or U20073 (N_20073,N_18532,N_18106);
or U20074 (N_20074,N_18651,N_18893);
nand U20075 (N_20075,N_18063,N_18974);
nor U20076 (N_20076,N_18480,N_19402);
xnor U20077 (N_20077,N_18720,N_19199);
and U20078 (N_20078,N_18772,N_19423);
and U20079 (N_20079,N_18755,N_18646);
or U20080 (N_20080,N_19255,N_18722);
nor U20081 (N_20081,N_18128,N_18903);
nand U20082 (N_20082,N_19405,N_18826);
nor U20083 (N_20083,N_18917,N_18482);
and U20084 (N_20084,N_19424,N_18707);
nand U20085 (N_20085,N_18781,N_18918);
nand U20086 (N_20086,N_18291,N_18091);
nor U20087 (N_20087,N_18041,N_18220);
or U20088 (N_20088,N_18393,N_18613);
nor U20089 (N_20089,N_18922,N_18474);
or U20090 (N_20090,N_19474,N_18423);
nor U20091 (N_20091,N_18978,N_18776);
or U20092 (N_20092,N_19074,N_18976);
nand U20093 (N_20093,N_18308,N_18268);
nor U20094 (N_20094,N_18104,N_19084);
or U20095 (N_20095,N_18382,N_18708);
nor U20096 (N_20096,N_18179,N_18050);
and U20097 (N_20097,N_18010,N_18726);
nor U20098 (N_20098,N_19152,N_18367);
nand U20099 (N_20099,N_18094,N_18383);
nand U20100 (N_20100,N_19252,N_18154);
nand U20101 (N_20101,N_19417,N_19197);
nand U20102 (N_20102,N_19388,N_18066);
nor U20103 (N_20103,N_18217,N_18946);
nor U20104 (N_20104,N_18068,N_19347);
nand U20105 (N_20105,N_19268,N_18493);
or U20106 (N_20106,N_18259,N_18120);
xnor U20107 (N_20107,N_19409,N_19216);
and U20108 (N_20108,N_18944,N_18366);
nand U20109 (N_20109,N_19284,N_18326);
nor U20110 (N_20110,N_18653,N_19256);
xor U20111 (N_20111,N_18750,N_19218);
xnor U20112 (N_20112,N_18501,N_19267);
or U20113 (N_20113,N_18384,N_18214);
xnor U20114 (N_20114,N_18710,N_18018);
xor U20115 (N_20115,N_19373,N_18191);
nor U20116 (N_20116,N_18485,N_18822);
nor U20117 (N_20117,N_18648,N_18414);
and U20118 (N_20118,N_19385,N_19413);
nand U20119 (N_20119,N_19018,N_18754);
nor U20120 (N_20120,N_19156,N_19348);
xnor U20121 (N_20121,N_19365,N_18638);
or U20122 (N_20122,N_18082,N_19185);
nor U20123 (N_20123,N_19188,N_19282);
or U20124 (N_20124,N_19077,N_18664);
or U20125 (N_20125,N_18468,N_19059);
xnor U20126 (N_20126,N_18076,N_18552);
nand U20127 (N_20127,N_19296,N_18264);
nand U20128 (N_20128,N_18136,N_18288);
or U20129 (N_20129,N_18774,N_18684);
or U20130 (N_20130,N_19181,N_19056);
and U20131 (N_20131,N_19047,N_18519);
nor U20132 (N_20132,N_19211,N_19306);
xor U20133 (N_20133,N_19288,N_18906);
and U20134 (N_20134,N_18505,N_18766);
nand U20135 (N_20135,N_19067,N_18760);
nor U20136 (N_20136,N_18514,N_18067);
xor U20137 (N_20137,N_18378,N_18620);
or U20138 (N_20138,N_18661,N_18433);
nor U20139 (N_20139,N_19486,N_18738);
and U20140 (N_20140,N_18556,N_19320);
or U20141 (N_20141,N_19253,N_18230);
and U20142 (N_20142,N_18003,N_18425);
nand U20143 (N_20143,N_18945,N_19395);
nor U20144 (N_20144,N_18598,N_18966);
and U20145 (N_20145,N_19420,N_18096);
nand U20146 (N_20146,N_19209,N_18330);
xor U20147 (N_20147,N_19225,N_19004);
xor U20148 (N_20148,N_18377,N_18705);
xnor U20149 (N_20149,N_19462,N_18335);
xor U20150 (N_20150,N_18586,N_19258);
nand U20151 (N_20151,N_18763,N_19045);
nand U20152 (N_20152,N_18920,N_19367);
and U20153 (N_20153,N_18235,N_18043);
nand U20154 (N_20154,N_19064,N_19376);
or U20155 (N_20155,N_18590,N_18702);
nand U20156 (N_20156,N_19239,N_18784);
or U20157 (N_20157,N_19399,N_19092);
xor U20158 (N_20158,N_18934,N_18891);
or U20159 (N_20159,N_18968,N_19021);
xor U20160 (N_20160,N_18582,N_19484);
nor U20161 (N_20161,N_18568,N_19223);
xnor U20162 (N_20162,N_18877,N_18634);
xor U20163 (N_20163,N_18858,N_19473);
nor U20164 (N_20164,N_18792,N_19483);
xnor U20165 (N_20165,N_18422,N_18703);
nand U20166 (N_20166,N_18995,N_19091);
or U20167 (N_20167,N_19456,N_18102);
nor U20168 (N_20168,N_19444,N_18064);
xor U20169 (N_20169,N_18087,N_19055);
nor U20170 (N_20170,N_18898,N_18325);
xnor U20171 (N_20171,N_18372,N_19449);
xor U20172 (N_20172,N_18931,N_18461);
and U20173 (N_20173,N_19235,N_19345);
or U20174 (N_20174,N_19020,N_18389);
or U20175 (N_20175,N_18641,N_18602);
or U20176 (N_20176,N_18352,N_18343);
or U20177 (N_20177,N_18984,N_18758);
nor U20178 (N_20178,N_18866,N_19371);
xnor U20179 (N_20179,N_18499,N_18475);
or U20180 (N_20180,N_19361,N_19013);
nand U20181 (N_20181,N_18243,N_18827);
or U20182 (N_20182,N_18024,N_18765);
or U20183 (N_20183,N_19390,N_19189);
nor U20184 (N_20184,N_18341,N_18533);
or U20185 (N_20185,N_19496,N_19133);
nor U20186 (N_20186,N_18443,N_18833);
nand U20187 (N_20187,N_18479,N_18473);
nand U20188 (N_20188,N_19353,N_19346);
nor U20189 (N_20189,N_18836,N_18497);
nand U20190 (N_20190,N_18843,N_19300);
xor U20191 (N_20191,N_19451,N_18856);
nand U20192 (N_20192,N_18540,N_18442);
or U20193 (N_20193,N_18234,N_18599);
nor U20194 (N_20194,N_18725,N_19457);
nor U20195 (N_20195,N_19153,N_18374);
xnor U20196 (N_20196,N_19453,N_18948);
nor U20197 (N_20197,N_18074,N_18459);
xor U20198 (N_20198,N_18958,N_19237);
nand U20199 (N_20199,N_18813,N_18675);
nand U20200 (N_20200,N_19220,N_19426);
nand U20201 (N_20201,N_18295,N_19167);
and U20202 (N_20202,N_18588,N_18890);
or U20203 (N_20203,N_18882,N_19058);
or U20204 (N_20204,N_18603,N_19271);
nor U20205 (N_20205,N_19464,N_18677);
xor U20206 (N_20206,N_18247,N_18852);
or U20207 (N_20207,N_18875,N_19360);
and U20208 (N_20208,N_18901,N_18788);
xnor U20209 (N_20209,N_19262,N_18197);
or U20210 (N_20210,N_18135,N_19259);
xnor U20211 (N_20211,N_18185,N_18452);
and U20212 (N_20212,N_19148,N_19000);
or U20213 (N_20213,N_19333,N_18070);
or U20214 (N_20214,N_18924,N_19200);
and U20215 (N_20215,N_18733,N_19314);
and U20216 (N_20216,N_18156,N_18849);
xor U20217 (N_20217,N_18237,N_19429);
or U20218 (N_20218,N_18569,N_18153);
and U20219 (N_20219,N_18162,N_19124);
xor U20220 (N_20220,N_18748,N_18400);
nand U20221 (N_20221,N_18663,N_18800);
nor U20222 (N_20222,N_18432,N_18696);
nand U20223 (N_20223,N_18057,N_18216);
and U20224 (N_20224,N_18510,N_18424);
nand U20225 (N_20225,N_18272,N_19026);
nand U20226 (N_20226,N_19028,N_18011);
xor U20227 (N_20227,N_18743,N_19375);
nand U20228 (N_20228,N_18525,N_19469);
nand U20229 (N_20229,N_19023,N_18248);
or U20230 (N_20230,N_18749,N_18515);
nor U20231 (N_20231,N_18768,N_18417);
xor U20232 (N_20232,N_18007,N_18117);
nor U20233 (N_20233,N_19418,N_18789);
nand U20234 (N_20234,N_18062,N_19291);
and U20235 (N_20235,N_18704,N_19017);
nor U20236 (N_20236,N_18693,N_19370);
or U20237 (N_20237,N_19014,N_18690);
nor U20238 (N_20238,N_19364,N_19460);
nor U20239 (N_20239,N_18936,N_18679);
nor U20240 (N_20240,N_19118,N_19245);
and U20241 (N_20241,N_18221,N_18125);
xnor U20242 (N_20242,N_19251,N_19198);
nand U20243 (N_20243,N_18438,N_18328);
xor U20244 (N_20244,N_19213,N_18909);
xnor U20245 (N_20245,N_19165,N_18790);
and U20246 (N_20246,N_18633,N_18348);
nand U20247 (N_20247,N_18450,N_18644);
nor U20248 (N_20248,N_19384,N_18778);
or U20249 (N_20249,N_18347,N_18200);
and U20250 (N_20250,N_18839,N_18991);
or U20251 (N_20251,N_18747,N_18766);
xor U20252 (N_20252,N_19066,N_18193);
nand U20253 (N_20253,N_19207,N_19497);
nor U20254 (N_20254,N_18873,N_18674);
nor U20255 (N_20255,N_18446,N_19067);
and U20256 (N_20256,N_18505,N_18926);
nor U20257 (N_20257,N_19463,N_18023);
or U20258 (N_20258,N_19225,N_18870);
xor U20259 (N_20259,N_18660,N_18843);
and U20260 (N_20260,N_19489,N_19112);
nor U20261 (N_20261,N_18052,N_18210);
and U20262 (N_20262,N_19362,N_18679);
xnor U20263 (N_20263,N_18551,N_18894);
nand U20264 (N_20264,N_19271,N_19287);
and U20265 (N_20265,N_18186,N_18033);
xor U20266 (N_20266,N_19085,N_18899);
or U20267 (N_20267,N_19236,N_18936);
and U20268 (N_20268,N_18766,N_18057);
xor U20269 (N_20269,N_19462,N_19196);
and U20270 (N_20270,N_19330,N_18684);
nand U20271 (N_20271,N_19079,N_19088);
and U20272 (N_20272,N_19303,N_18234);
and U20273 (N_20273,N_19073,N_18135);
xor U20274 (N_20274,N_19145,N_18387);
and U20275 (N_20275,N_18598,N_18520);
xnor U20276 (N_20276,N_19450,N_18860);
and U20277 (N_20277,N_19405,N_18325);
or U20278 (N_20278,N_19401,N_18631);
and U20279 (N_20279,N_18279,N_18767);
nand U20280 (N_20280,N_18001,N_18546);
or U20281 (N_20281,N_19225,N_19076);
nor U20282 (N_20282,N_18316,N_18451);
xor U20283 (N_20283,N_19073,N_18329);
nand U20284 (N_20284,N_18671,N_19329);
xor U20285 (N_20285,N_19124,N_18133);
or U20286 (N_20286,N_18083,N_19119);
nand U20287 (N_20287,N_18088,N_18167);
nand U20288 (N_20288,N_19037,N_18666);
xor U20289 (N_20289,N_18922,N_19463);
xor U20290 (N_20290,N_18340,N_18287);
xnor U20291 (N_20291,N_19028,N_18275);
nand U20292 (N_20292,N_18014,N_19268);
nor U20293 (N_20293,N_18112,N_18656);
xor U20294 (N_20294,N_18118,N_19450);
nor U20295 (N_20295,N_18485,N_18573);
nor U20296 (N_20296,N_19429,N_18309);
or U20297 (N_20297,N_18113,N_18557);
or U20298 (N_20298,N_19449,N_19133);
or U20299 (N_20299,N_18800,N_18967);
nand U20300 (N_20300,N_18365,N_19215);
or U20301 (N_20301,N_18185,N_19254);
nor U20302 (N_20302,N_18057,N_19331);
nor U20303 (N_20303,N_19274,N_18461);
xor U20304 (N_20304,N_18229,N_18596);
nor U20305 (N_20305,N_19042,N_19127);
nand U20306 (N_20306,N_19358,N_19203);
and U20307 (N_20307,N_18214,N_18861);
xnor U20308 (N_20308,N_18348,N_19241);
and U20309 (N_20309,N_19195,N_18554);
nand U20310 (N_20310,N_18775,N_19028);
and U20311 (N_20311,N_18853,N_18381);
nor U20312 (N_20312,N_18038,N_18930);
or U20313 (N_20313,N_18994,N_19058);
xor U20314 (N_20314,N_19428,N_19017);
nand U20315 (N_20315,N_18009,N_18342);
and U20316 (N_20316,N_18600,N_19348);
nand U20317 (N_20317,N_18960,N_19104);
xor U20318 (N_20318,N_18448,N_18636);
nand U20319 (N_20319,N_18359,N_18805);
nand U20320 (N_20320,N_18111,N_18211);
or U20321 (N_20321,N_18089,N_18669);
and U20322 (N_20322,N_18506,N_18960);
xor U20323 (N_20323,N_18181,N_19490);
nand U20324 (N_20324,N_18339,N_18280);
or U20325 (N_20325,N_19347,N_18770);
xnor U20326 (N_20326,N_19062,N_18220);
or U20327 (N_20327,N_18820,N_18895);
xnor U20328 (N_20328,N_18441,N_19060);
xor U20329 (N_20329,N_18546,N_19059);
or U20330 (N_20330,N_18374,N_19182);
nand U20331 (N_20331,N_18943,N_19223);
xnor U20332 (N_20332,N_19448,N_18504);
nor U20333 (N_20333,N_19371,N_18715);
or U20334 (N_20334,N_18555,N_18671);
nor U20335 (N_20335,N_18044,N_18102);
nor U20336 (N_20336,N_18075,N_19240);
xnor U20337 (N_20337,N_19455,N_19230);
nand U20338 (N_20338,N_18892,N_18870);
nand U20339 (N_20339,N_19492,N_19162);
nand U20340 (N_20340,N_18765,N_18720);
xor U20341 (N_20341,N_18594,N_19294);
xnor U20342 (N_20342,N_18714,N_19431);
nand U20343 (N_20343,N_19472,N_19360);
nand U20344 (N_20344,N_18695,N_18580);
nor U20345 (N_20345,N_18765,N_19010);
and U20346 (N_20346,N_18694,N_19110);
nor U20347 (N_20347,N_19426,N_18073);
xnor U20348 (N_20348,N_19331,N_18046);
and U20349 (N_20349,N_19342,N_18717);
xor U20350 (N_20350,N_18156,N_18283);
or U20351 (N_20351,N_18249,N_18578);
or U20352 (N_20352,N_18781,N_18709);
xor U20353 (N_20353,N_19436,N_19021);
xor U20354 (N_20354,N_18021,N_18828);
and U20355 (N_20355,N_18647,N_18575);
or U20356 (N_20356,N_19346,N_18055);
nor U20357 (N_20357,N_18947,N_18047);
nand U20358 (N_20358,N_19420,N_18860);
nand U20359 (N_20359,N_18780,N_19422);
xor U20360 (N_20360,N_18515,N_19469);
nor U20361 (N_20361,N_18680,N_19499);
and U20362 (N_20362,N_18121,N_18902);
nor U20363 (N_20363,N_18115,N_18651);
nor U20364 (N_20364,N_18190,N_18305);
nand U20365 (N_20365,N_18235,N_19108);
nand U20366 (N_20366,N_19101,N_18299);
nor U20367 (N_20367,N_18226,N_18543);
nand U20368 (N_20368,N_18895,N_18932);
nand U20369 (N_20369,N_18402,N_19388);
or U20370 (N_20370,N_18749,N_19441);
and U20371 (N_20371,N_18214,N_18569);
and U20372 (N_20372,N_18817,N_18398);
and U20373 (N_20373,N_18153,N_19160);
xor U20374 (N_20374,N_18909,N_18854);
xor U20375 (N_20375,N_19055,N_18372);
xor U20376 (N_20376,N_18530,N_18407);
nor U20377 (N_20377,N_18288,N_19114);
xnor U20378 (N_20378,N_18785,N_18870);
nor U20379 (N_20379,N_18329,N_18812);
nor U20380 (N_20380,N_19268,N_18851);
or U20381 (N_20381,N_18451,N_18894);
xor U20382 (N_20382,N_18174,N_19026);
or U20383 (N_20383,N_18628,N_18654);
nand U20384 (N_20384,N_18202,N_19497);
xnor U20385 (N_20385,N_18913,N_19312);
nor U20386 (N_20386,N_19479,N_18415);
or U20387 (N_20387,N_18103,N_18407);
or U20388 (N_20388,N_18115,N_18844);
nand U20389 (N_20389,N_19184,N_19232);
xnor U20390 (N_20390,N_19401,N_19423);
nor U20391 (N_20391,N_18416,N_18060);
nand U20392 (N_20392,N_18393,N_18856);
xor U20393 (N_20393,N_18347,N_18836);
nor U20394 (N_20394,N_18652,N_18387);
nor U20395 (N_20395,N_19273,N_19350);
xnor U20396 (N_20396,N_18286,N_18424);
and U20397 (N_20397,N_19389,N_18661);
xor U20398 (N_20398,N_19476,N_18846);
xor U20399 (N_20399,N_19030,N_18744);
and U20400 (N_20400,N_18524,N_18001);
nand U20401 (N_20401,N_18578,N_18473);
nand U20402 (N_20402,N_18304,N_18042);
and U20403 (N_20403,N_19368,N_18776);
xor U20404 (N_20404,N_19105,N_18845);
xor U20405 (N_20405,N_19107,N_19104);
nand U20406 (N_20406,N_18532,N_19120);
and U20407 (N_20407,N_18876,N_18961);
nor U20408 (N_20408,N_18521,N_18980);
or U20409 (N_20409,N_19453,N_19174);
xnor U20410 (N_20410,N_19100,N_19246);
and U20411 (N_20411,N_19143,N_18396);
or U20412 (N_20412,N_18933,N_18604);
and U20413 (N_20413,N_18898,N_18660);
nand U20414 (N_20414,N_18036,N_18348);
or U20415 (N_20415,N_19475,N_19171);
and U20416 (N_20416,N_18101,N_18523);
or U20417 (N_20417,N_18912,N_18891);
xor U20418 (N_20418,N_19129,N_18129);
nand U20419 (N_20419,N_19368,N_18114);
or U20420 (N_20420,N_18565,N_19122);
or U20421 (N_20421,N_19363,N_18081);
or U20422 (N_20422,N_18691,N_18258);
or U20423 (N_20423,N_18974,N_19146);
nand U20424 (N_20424,N_19185,N_18755);
nand U20425 (N_20425,N_18467,N_18250);
nor U20426 (N_20426,N_18521,N_19161);
xnor U20427 (N_20427,N_18325,N_18614);
or U20428 (N_20428,N_18642,N_18400);
nor U20429 (N_20429,N_18490,N_18400);
nand U20430 (N_20430,N_18924,N_18431);
nand U20431 (N_20431,N_18392,N_18721);
nand U20432 (N_20432,N_19491,N_18415);
nand U20433 (N_20433,N_18630,N_18247);
xnor U20434 (N_20434,N_19173,N_18389);
or U20435 (N_20435,N_18689,N_18835);
nand U20436 (N_20436,N_19183,N_19061);
nor U20437 (N_20437,N_18517,N_19384);
or U20438 (N_20438,N_18941,N_19350);
nor U20439 (N_20439,N_19027,N_18075);
xor U20440 (N_20440,N_18193,N_18012);
nand U20441 (N_20441,N_19188,N_18465);
nand U20442 (N_20442,N_19047,N_19032);
and U20443 (N_20443,N_18901,N_19050);
or U20444 (N_20444,N_18359,N_18856);
nor U20445 (N_20445,N_18761,N_19151);
nand U20446 (N_20446,N_18756,N_18358);
nand U20447 (N_20447,N_18958,N_18369);
xnor U20448 (N_20448,N_18384,N_18285);
or U20449 (N_20449,N_18985,N_19323);
or U20450 (N_20450,N_19398,N_18217);
and U20451 (N_20451,N_18219,N_18390);
nor U20452 (N_20452,N_18729,N_18722);
nor U20453 (N_20453,N_18284,N_18426);
and U20454 (N_20454,N_18925,N_18412);
nand U20455 (N_20455,N_19372,N_18249);
xor U20456 (N_20456,N_18377,N_18928);
or U20457 (N_20457,N_18561,N_18538);
or U20458 (N_20458,N_18369,N_18642);
and U20459 (N_20459,N_18651,N_18926);
nand U20460 (N_20460,N_19114,N_18132);
or U20461 (N_20461,N_18746,N_19134);
or U20462 (N_20462,N_18712,N_19314);
xor U20463 (N_20463,N_19254,N_19448);
and U20464 (N_20464,N_19041,N_18633);
nor U20465 (N_20465,N_19308,N_18095);
or U20466 (N_20466,N_18550,N_18531);
nand U20467 (N_20467,N_18846,N_18120);
nand U20468 (N_20468,N_18383,N_18365);
and U20469 (N_20469,N_19008,N_19050);
xnor U20470 (N_20470,N_18552,N_18569);
or U20471 (N_20471,N_18918,N_18175);
or U20472 (N_20472,N_18606,N_18163);
xnor U20473 (N_20473,N_19395,N_18442);
or U20474 (N_20474,N_18042,N_19064);
nand U20475 (N_20475,N_18690,N_18645);
and U20476 (N_20476,N_18051,N_19103);
nor U20477 (N_20477,N_18556,N_19265);
or U20478 (N_20478,N_18954,N_18270);
nand U20479 (N_20479,N_19230,N_19361);
nor U20480 (N_20480,N_18211,N_19088);
nand U20481 (N_20481,N_18198,N_18411);
nor U20482 (N_20482,N_18463,N_18540);
nand U20483 (N_20483,N_18184,N_18002);
nand U20484 (N_20484,N_19308,N_19146);
nor U20485 (N_20485,N_18642,N_18247);
and U20486 (N_20486,N_18900,N_19347);
or U20487 (N_20487,N_19390,N_19114);
nor U20488 (N_20488,N_19045,N_19419);
nor U20489 (N_20489,N_19370,N_18439);
or U20490 (N_20490,N_19220,N_18772);
or U20491 (N_20491,N_19499,N_18643);
or U20492 (N_20492,N_19299,N_18394);
nand U20493 (N_20493,N_19112,N_18756);
or U20494 (N_20494,N_19408,N_18374);
and U20495 (N_20495,N_18215,N_18975);
or U20496 (N_20496,N_18580,N_19134);
nor U20497 (N_20497,N_18051,N_19002);
and U20498 (N_20498,N_18528,N_18967);
xnor U20499 (N_20499,N_18588,N_19068);
nand U20500 (N_20500,N_18336,N_18952);
or U20501 (N_20501,N_18418,N_18561);
and U20502 (N_20502,N_18206,N_19222);
or U20503 (N_20503,N_19482,N_18135);
and U20504 (N_20504,N_18248,N_19128);
and U20505 (N_20505,N_18506,N_18799);
nor U20506 (N_20506,N_18040,N_19231);
nand U20507 (N_20507,N_18905,N_18524);
nor U20508 (N_20508,N_18621,N_18063);
or U20509 (N_20509,N_18902,N_18414);
nor U20510 (N_20510,N_18824,N_18606);
nand U20511 (N_20511,N_18992,N_18573);
xnor U20512 (N_20512,N_18912,N_18764);
nor U20513 (N_20513,N_18286,N_18105);
nor U20514 (N_20514,N_18165,N_19062);
and U20515 (N_20515,N_18685,N_19325);
xor U20516 (N_20516,N_18501,N_19318);
or U20517 (N_20517,N_18629,N_19247);
or U20518 (N_20518,N_18733,N_18184);
nand U20519 (N_20519,N_18358,N_19202);
nand U20520 (N_20520,N_19028,N_18808);
nand U20521 (N_20521,N_19446,N_19081);
nand U20522 (N_20522,N_19318,N_18245);
or U20523 (N_20523,N_18541,N_18173);
nor U20524 (N_20524,N_18502,N_19163);
and U20525 (N_20525,N_18296,N_18822);
nand U20526 (N_20526,N_19391,N_18062);
xor U20527 (N_20527,N_18437,N_19312);
nor U20528 (N_20528,N_19291,N_18296);
nand U20529 (N_20529,N_19274,N_18004);
and U20530 (N_20530,N_18965,N_18586);
and U20531 (N_20531,N_18881,N_18180);
nor U20532 (N_20532,N_18417,N_18956);
and U20533 (N_20533,N_19446,N_18036);
and U20534 (N_20534,N_19147,N_19226);
xor U20535 (N_20535,N_19402,N_18049);
and U20536 (N_20536,N_18217,N_18382);
nand U20537 (N_20537,N_18997,N_18996);
or U20538 (N_20538,N_18019,N_18008);
nand U20539 (N_20539,N_19016,N_19296);
xnor U20540 (N_20540,N_18238,N_18201);
nor U20541 (N_20541,N_18330,N_18559);
nand U20542 (N_20542,N_19432,N_18397);
nor U20543 (N_20543,N_18482,N_18373);
nor U20544 (N_20544,N_18972,N_18828);
xnor U20545 (N_20545,N_18243,N_18432);
nor U20546 (N_20546,N_19289,N_18886);
and U20547 (N_20547,N_18456,N_18137);
nor U20548 (N_20548,N_18740,N_18072);
xnor U20549 (N_20549,N_18530,N_18739);
nand U20550 (N_20550,N_18756,N_18320);
or U20551 (N_20551,N_18654,N_19404);
and U20552 (N_20552,N_19210,N_18589);
xor U20553 (N_20553,N_18506,N_18089);
xnor U20554 (N_20554,N_18583,N_18470);
and U20555 (N_20555,N_19434,N_19076);
and U20556 (N_20556,N_19364,N_18157);
xor U20557 (N_20557,N_19191,N_18578);
xnor U20558 (N_20558,N_18710,N_18253);
nand U20559 (N_20559,N_19331,N_18846);
nand U20560 (N_20560,N_18715,N_19203);
nor U20561 (N_20561,N_18174,N_18817);
or U20562 (N_20562,N_18570,N_19479);
nand U20563 (N_20563,N_18028,N_19213);
or U20564 (N_20564,N_18395,N_18006);
nand U20565 (N_20565,N_18491,N_19206);
xor U20566 (N_20566,N_18274,N_19071);
xor U20567 (N_20567,N_19465,N_19191);
or U20568 (N_20568,N_18706,N_18749);
and U20569 (N_20569,N_18760,N_18022);
nand U20570 (N_20570,N_18337,N_18843);
or U20571 (N_20571,N_18511,N_18726);
xor U20572 (N_20572,N_18307,N_18893);
nand U20573 (N_20573,N_19379,N_18181);
nor U20574 (N_20574,N_18469,N_18237);
or U20575 (N_20575,N_19236,N_18071);
and U20576 (N_20576,N_19431,N_18332);
xor U20577 (N_20577,N_18154,N_19093);
nand U20578 (N_20578,N_19148,N_19247);
and U20579 (N_20579,N_19281,N_18609);
and U20580 (N_20580,N_19112,N_18497);
nor U20581 (N_20581,N_18705,N_19345);
nand U20582 (N_20582,N_18198,N_18306);
or U20583 (N_20583,N_18264,N_18131);
nor U20584 (N_20584,N_18711,N_18079);
nor U20585 (N_20585,N_18486,N_19447);
and U20586 (N_20586,N_18942,N_18047);
and U20587 (N_20587,N_18915,N_18359);
nand U20588 (N_20588,N_19455,N_18427);
nor U20589 (N_20589,N_18404,N_18289);
and U20590 (N_20590,N_19458,N_18989);
xor U20591 (N_20591,N_18100,N_19422);
and U20592 (N_20592,N_18772,N_18538);
xnor U20593 (N_20593,N_18022,N_18667);
xor U20594 (N_20594,N_18855,N_18081);
nand U20595 (N_20595,N_19457,N_19290);
xor U20596 (N_20596,N_18185,N_18966);
nand U20597 (N_20597,N_18985,N_19014);
and U20598 (N_20598,N_18017,N_18765);
xor U20599 (N_20599,N_19031,N_18475);
xor U20600 (N_20600,N_18417,N_18127);
nand U20601 (N_20601,N_19115,N_19288);
nor U20602 (N_20602,N_19146,N_19407);
nand U20603 (N_20603,N_18549,N_19234);
and U20604 (N_20604,N_19347,N_19376);
and U20605 (N_20605,N_18786,N_18192);
or U20606 (N_20606,N_19373,N_19210);
nand U20607 (N_20607,N_18984,N_18460);
nand U20608 (N_20608,N_18249,N_19083);
and U20609 (N_20609,N_18878,N_19204);
xnor U20610 (N_20610,N_18009,N_18679);
and U20611 (N_20611,N_18188,N_18342);
nor U20612 (N_20612,N_18564,N_19266);
nor U20613 (N_20613,N_19125,N_19322);
nand U20614 (N_20614,N_18785,N_18720);
or U20615 (N_20615,N_18595,N_18124);
and U20616 (N_20616,N_18569,N_19191);
nand U20617 (N_20617,N_18342,N_18960);
and U20618 (N_20618,N_18881,N_18525);
nor U20619 (N_20619,N_18095,N_19169);
xor U20620 (N_20620,N_18820,N_18028);
xor U20621 (N_20621,N_18343,N_18444);
and U20622 (N_20622,N_18397,N_19134);
nand U20623 (N_20623,N_19017,N_19278);
nor U20624 (N_20624,N_19092,N_18653);
xnor U20625 (N_20625,N_18294,N_18281);
xor U20626 (N_20626,N_18624,N_19223);
or U20627 (N_20627,N_18980,N_19025);
or U20628 (N_20628,N_18619,N_18064);
nand U20629 (N_20629,N_19048,N_18501);
or U20630 (N_20630,N_19032,N_18833);
xor U20631 (N_20631,N_18253,N_18794);
xor U20632 (N_20632,N_18553,N_19238);
and U20633 (N_20633,N_18939,N_19400);
xor U20634 (N_20634,N_18664,N_18361);
nand U20635 (N_20635,N_18300,N_19442);
and U20636 (N_20636,N_18778,N_18434);
or U20637 (N_20637,N_18597,N_18955);
xor U20638 (N_20638,N_18893,N_19476);
and U20639 (N_20639,N_18522,N_19034);
nor U20640 (N_20640,N_19373,N_18117);
nor U20641 (N_20641,N_18526,N_18431);
nor U20642 (N_20642,N_19404,N_18572);
xor U20643 (N_20643,N_19167,N_19428);
or U20644 (N_20644,N_18130,N_18474);
or U20645 (N_20645,N_18048,N_18447);
nor U20646 (N_20646,N_18453,N_19128);
xor U20647 (N_20647,N_18064,N_18232);
or U20648 (N_20648,N_18954,N_18828);
or U20649 (N_20649,N_18774,N_18245);
or U20650 (N_20650,N_19104,N_19014);
nand U20651 (N_20651,N_18635,N_18266);
xor U20652 (N_20652,N_18685,N_18355);
or U20653 (N_20653,N_19263,N_19031);
or U20654 (N_20654,N_18927,N_18233);
nand U20655 (N_20655,N_18417,N_19431);
and U20656 (N_20656,N_19070,N_19167);
xor U20657 (N_20657,N_19310,N_18207);
or U20658 (N_20658,N_19222,N_18041);
or U20659 (N_20659,N_18897,N_19390);
nand U20660 (N_20660,N_18536,N_19499);
xnor U20661 (N_20661,N_19248,N_19181);
or U20662 (N_20662,N_18504,N_19026);
xnor U20663 (N_20663,N_18617,N_18653);
xnor U20664 (N_20664,N_19145,N_18167);
and U20665 (N_20665,N_18703,N_19407);
nor U20666 (N_20666,N_18177,N_19176);
and U20667 (N_20667,N_18059,N_19359);
nand U20668 (N_20668,N_18656,N_18618);
and U20669 (N_20669,N_19406,N_19025);
and U20670 (N_20670,N_19498,N_19079);
nand U20671 (N_20671,N_18906,N_18486);
nand U20672 (N_20672,N_18709,N_18396);
nor U20673 (N_20673,N_19061,N_18577);
and U20674 (N_20674,N_18463,N_18390);
and U20675 (N_20675,N_18574,N_18522);
nand U20676 (N_20676,N_18421,N_18991);
and U20677 (N_20677,N_18734,N_18449);
or U20678 (N_20678,N_19408,N_18401);
and U20679 (N_20679,N_18892,N_18385);
xnor U20680 (N_20680,N_19436,N_18707);
and U20681 (N_20681,N_18362,N_19363);
xnor U20682 (N_20682,N_18398,N_19018);
nor U20683 (N_20683,N_18767,N_18478);
nor U20684 (N_20684,N_18841,N_18646);
nand U20685 (N_20685,N_18519,N_18995);
or U20686 (N_20686,N_18436,N_19009);
nand U20687 (N_20687,N_18176,N_18963);
and U20688 (N_20688,N_18081,N_18984);
xor U20689 (N_20689,N_19298,N_19302);
nor U20690 (N_20690,N_18119,N_18713);
and U20691 (N_20691,N_18546,N_18715);
or U20692 (N_20692,N_18260,N_19248);
nand U20693 (N_20693,N_19021,N_19168);
nor U20694 (N_20694,N_18483,N_19410);
nor U20695 (N_20695,N_18320,N_18789);
xor U20696 (N_20696,N_18836,N_19361);
nor U20697 (N_20697,N_18536,N_18061);
nand U20698 (N_20698,N_18697,N_19269);
and U20699 (N_20699,N_19385,N_18523);
or U20700 (N_20700,N_18080,N_18177);
nand U20701 (N_20701,N_19133,N_19293);
nand U20702 (N_20702,N_19366,N_18389);
nand U20703 (N_20703,N_19104,N_19362);
and U20704 (N_20704,N_19014,N_18756);
xnor U20705 (N_20705,N_19184,N_19299);
or U20706 (N_20706,N_18808,N_18362);
or U20707 (N_20707,N_18643,N_19010);
xor U20708 (N_20708,N_18485,N_18889);
or U20709 (N_20709,N_19228,N_18546);
or U20710 (N_20710,N_18754,N_18421);
xnor U20711 (N_20711,N_18609,N_19269);
and U20712 (N_20712,N_19301,N_18871);
xnor U20713 (N_20713,N_19207,N_19369);
nand U20714 (N_20714,N_18974,N_19219);
nor U20715 (N_20715,N_18932,N_19038);
nand U20716 (N_20716,N_18316,N_18197);
nor U20717 (N_20717,N_19480,N_18135);
nand U20718 (N_20718,N_18249,N_19425);
and U20719 (N_20719,N_18307,N_18202);
nor U20720 (N_20720,N_18214,N_19017);
and U20721 (N_20721,N_19118,N_19234);
xor U20722 (N_20722,N_19073,N_18602);
or U20723 (N_20723,N_19266,N_18150);
nand U20724 (N_20724,N_18551,N_18816);
nor U20725 (N_20725,N_18391,N_19064);
or U20726 (N_20726,N_18327,N_18788);
nor U20727 (N_20727,N_18596,N_19159);
or U20728 (N_20728,N_18042,N_19186);
xor U20729 (N_20729,N_18764,N_19136);
xnor U20730 (N_20730,N_18818,N_18213);
nor U20731 (N_20731,N_19322,N_18274);
nand U20732 (N_20732,N_18581,N_19080);
nor U20733 (N_20733,N_18607,N_19006);
or U20734 (N_20734,N_18526,N_18995);
and U20735 (N_20735,N_18278,N_18329);
nand U20736 (N_20736,N_18751,N_18463);
or U20737 (N_20737,N_18724,N_18863);
nand U20738 (N_20738,N_18979,N_18576);
xnor U20739 (N_20739,N_18926,N_18023);
and U20740 (N_20740,N_18331,N_18304);
or U20741 (N_20741,N_18309,N_18051);
nor U20742 (N_20742,N_18219,N_18506);
nand U20743 (N_20743,N_18528,N_19175);
or U20744 (N_20744,N_19209,N_18596);
xnor U20745 (N_20745,N_19114,N_18751);
or U20746 (N_20746,N_18410,N_18771);
and U20747 (N_20747,N_18458,N_18969);
xnor U20748 (N_20748,N_19347,N_18961);
nor U20749 (N_20749,N_18484,N_19206);
nand U20750 (N_20750,N_18283,N_18963);
or U20751 (N_20751,N_19268,N_18049);
or U20752 (N_20752,N_18744,N_18688);
nand U20753 (N_20753,N_19347,N_18189);
and U20754 (N_20754,N_18576,N_19042);
or U20755 (N_20755,N_18797,N_19251);
xor U20756 (N_20756,N_19036,N_18352);
or U20757 (N_20757,N_18107,N_18260);
and U20758 (N_20758,N_18228,N_19372);
or U20759 (N_20759,N_19013,N_18772);
or U20760 (N_20760,N_19393,N_18083);
and U20761 (N_20761,N_19462,N_18163);
nand U20762 (N_20762,N_19362,N_18883);
or U20763 (N_20763,N_18643,N_19412);
or U20764 (N_20764,N_18384,N_19058);
or U20765 (N_20765,N_18924,N_19262);
and U20766 (N_20766,N_18110,N_19488);
xor U20767 (N_20767,N_19153,N_18471);
xor U20768 (N_20768,N_18016,N_18138);
xor U20769 (N_20769,N_19387,N_18254);
or U20770 (N_20770,N_18028,N_18585);
or U20771 (N_20771,N_18200,N_18841);
xor U20772 (N_20772,N_19304,N_18419);
and U20773 (N_20773,N_19306,N_19115);
and U20774 (N_20774,N_19284,N_18636);
nor U20775 (N_20775,N_18329,N_19316);
and U20776 (N_20776,N_18437,N_18895);
xor U20777 (N_20777,N_18346,N_19193);
nand U20778 (N_20778,N_18881,N_19249);
xor U20779 (N_20779,N_19000,N_18495);
nand U20780 (N_20780,N_19135,N_18308);
nor U20781 (N_20781,N_18184,N_19007);
or U20782 (N_20782,N_19221,N_19425);
nand U20783 (N_20783,N_18054,N_18797);
nor U20784 (N_20784,N_18336,N_19448);
xor U20785 (N_20785,N_18084,N_18586);
and U20786 (N_20786,N_19433,N_18461);
nor U20787 (N_20787,N_19062,N_18396);
nand U20788 (N_20788,N_18860,N_18917);
nand U20789 (N_20789,N_18958,N_18890);
nand U20790 (N_20790,N_18660,N_18047);
nand U20791 (N_20791,N_18156,N_18052);
nand U20792 (N_20792,N_18975,N_18145);
xor U20793 (N_20793,N_18085,N_19420);
and U20794 (N_20794,N_18288,N_19336);
nand U20795 (N_20795,N_18444,N_18130);
and U20796 (N_20796,N_18022,N_19152);
nor U20797 (N_20797,N_18169,N_19007);
nand U20798 (N_20798,N_18273,N_18116);
and U20799 (N_20799,N_18977,N_18415);
nor U20800 (N_20800,N_18117,N_19153);
and U20801 (N_20801,N_18795,N_18316);
and U20802 (N_20802,N_18492,N_18124);
nand U20803 (N_20803,N_18242,N_18374);
nor U20804 (N_20804,N_18459,N_19470);
nand U20805 (N_20805,N_18712,N_19123);
nand U20806 (N_20806,N_18693,N_19176);
and U20807 (N_20807,N_19266,N_19305);
and U20808 (N_20808,N_19480,N_18493);
or U20809 (N_20809,N_19284,N_19274);
xor U20810 (N_20810,N_18147,N_18030);
or U20811 (N_20811,N_18637,N_18841);
and U20812 (N_20812,N_18075,N_18693);
nand U20813 (N_20813,N_19107,N_18606);
or U20814 (N_20814,N_18155,N_19404);
nand U20815 (N_20815,N_19092,N_19327);
and U20816 (N_20816,N_19242,N_18515);
and U20817 (N_20817,N_18245,N_18318);
or U20818 (N_20818,N_18023,N_18570);
or U20819 (N_20819,N_18451,N_18876);
nor U20820 (N_20820,N_18323,N_19317);
xor U20821 (N_20821,N_18318,N_18098);
or U20822 (N_20822,N_18269,N_19344);
nand U20823 (N_20823,N_18970,N_18727);
xor U20824 (N_20824,N_18314,N_19372);
and U20825 (N_20825,N_18807,N_18511);
nand U20826 (N_20826,N_19468,N_19034);
and U20827 (N_20827,N_19103,N_19202);
or U20828 (N_20828,N_18649,N_18334);
xor U20829 (N_20829,N_18010,N_19200);
and U20830 (N_20830,N_19485,N_19182);
xnor U20831 (N_20831,N_18158,N_18239);
nand U20832 (N_20832,N_18668,N_18645);
xor U20833 (N_20833,N_18850,N_18621);
xnor U20834 (N_20834,N_18216,N_19087);
nand U20835 (N_20835,N_19173,N_18758);
or U20836 (N_20836,N_19416,N_18959);
xnor U20837 (N_20837,N_18645,N_19243);
and U20838 (N_20838,N_19080,N_19125);
nor U20839 (N_20839,N_18139,N_18189);
or U20840 (N_20840,N_19484,N_19411);
and U20841 (N_20841,N_18447,N_18983);
and U20842 (N_20842,N_18910,N_19265);
and U20843 (N_20843,N_18656,N_18267);
nor U20844 (N_20844,N_18082,N_19467);
xnor U20845 (N_20845,N_18254,N_18227);
and U20846 (N_20846,N_18467,N_18120);
xnor U20847 (N_20847,N_18083,N_18371);
and U20848 (N_20848,N_18109,N_19210);
or U20849 (N_20849,N_19068,N_18701);
or U20850 (N_20850,N_19048,N_19133);
nor U20851 (N_20851,N_18487,N_18380);
nand U20852 (N_20852,N_19129,N_18830);
nand U20853 (N_20853,N_18271,N_19025);
xor U20854 (N_20854,N_19158,N_18280);
and U20855 (N_20855,N_18796,N_18248);
and U20856 (N_20856,N_18077,N_18430);
and U20857 (N_20857,N_18808,N_19316);
and U20858 (N_20858,N_18874,N_18957);
and U20859 (N_20859,N_18026,N_19450);
or U20860 (N_20860,N_18184,N_19103);
or U20861 (N_20861,N_18208,N_18166);
xor U20862 (N_20862,N_18086,N_18711);
and U20863 (N_20863,N_18226,N_18382);
nor U20864 (N_20864,N_18153,N_19320);
or U20865 (N_20865,N_18528,N_18094);
and U20866 (N_20866,N_19206,N_18010);
or U20867 (N_20867,N_19388,N_19335);
or U20868 (N_20868,N_18137,N_18738);
nor U20869 (N_20869,N_19034,N_18563);
nor U20870 (N_20870,N_18607,N_19327);
nand U20871 (N_20871,N_18506,N_18329);
xor U20872 (N_20872,N_18921,N_18055);
nand U20873 (N_20873,N_19233,N_18383);
xnor U20874 (N_20874,N_18456,N_18808);
nor U20875 (N_20875,N_19015,N_19402);
and U20876 (N_20876,N_18405,N_18500);
nor U20877 (N_20877,N_19264,N_18745);
or U20878 (N_20878,N_18454,N_18299);
nor U20879 (N_20879,N_18783,N_19177);
and U20880 (N_20880,N_18155,N_18242);
nand U20881 (N_20881,N_18307,N_18642);
xor U20882 (N_20882,N_18837,N_18146);
xnor U20883 (N_20883,N_18638,N_19220);
and U20884 (N_20884,N_18140,N_18922);
nor U20885 (N_20885,N_19369,N_18308);
or U20886 (N_20886,N_18866,N_18151);
xnor U20887 (N_20887,N_18066,N_18304);
nand U20888 (N_20888,N_18091,N_19013);
and U20889 (N_20889,N_19356,N_19137);
nor U20890 (N_20890,N_18674,N_18378);
and U20891 (N_20891,N_19033,N_18686);
xor U20892 (N_20892,N_19420,N_18438);
and U20893 (N_20893,N_18358,N_19420);
nor U20894 (N_20894,N_18954,N_19052);
xor U20895 (N_20895,N_18120,N_18743);
or U20896 (N_20896,N_18041,N_18805);
or U20897 (N_20897,N_19128,N_19076);
nor U20898 (N_20898,N_18590,N_18573);
nor U20899 (N_20899,N_18852,N_19413);
and U20900 (N_20900,N_19112,N_18242);
or U20901 (N_20901,N_18431,N_18140);
and U20902 (N_20902,N_18805,N_18242);
or U20903 (N_20903,N_18759,N_18198);
or U20904 (N_20904,N_19236,N_18432);
xnor U20905 (N_20905,N_18297,N_19273);
nor U20906 (N_20906,N_19001,N_18926);
and U20907 (N_20907,N_18995,N_18708);
or U20908 (N_20908,N_18006,N_18909);
nand U20909 (N_20909,N_18470,N_19079);
nor U20910 (N_20910,N_18055,N_19471);
nand U20911 (N_20911,N_18647,N_18992);
xnor U20912 (N_20912,N_18142,N_19339);
xnor U20913 (N_20913,N_18252,N_18180);
or U20914 (N_20914,N_18639,N_18562);
and U20915 (N_20915,N_19295,N_18627);
and U20916 (N_20916,N_18676,N_18495);
nor U20917 (N_20917,N_18444,N_18622);
and U20918 (N_20918,N_18226,N_18090);
nor U20919 (N_20919,N_18094,N_19093);
xor U20920 (N_20920,N_18488,N_18018);
xor U20921 (N_20921,N_18339,N_19392);
or U20922 (N_20922,N_18916,N_18557);
xnor U20923 (N_20923,N_19255,N_19041);
nand U20924 (N_20924,N_19456,N_18113);
nand U20925 (N_20925,N_19332,N_18882);
and U20926 (N_20926,N_18746,N_18769);
and U20927 (N_20927,N_18231,N_19272);
nand U20928 (N_20928,N_19099,N_18919);
nor U20929 (N_20929,N_18841,N_18466);
nor U20930 (N_20930,N_19271,N_18915);
nand U20931 (N_20931,N_19256,N_19354);
nand U20932 (N_20932,N_18213,N_18833);
and U20933 (N_20933,N_19128,N_18671);
nand U20934 (N_20934,N_18149,N_18611);
or U20935 (N_20935,N_18768,N_18538);
and U20936 (N_20936,N_19388,N_19030);
nand U20937 (N_20937,N_18408,N_19137);
nand U20938 (N_20938,N_19479,N_18311);
nor U20939 (N_20939,N_18624,N_19092);
nor U20940 (N_20940,N_19227,N_18713);
nor U20941 (N_20941,N_18170,N_19320);
nand U20942 (N_20942,N_18952,N_18258);
nor U20943 (N_20943,N_18465,N_18579);
or U20944 (N_20944,N_18070,N_18111);
nor U20945 (N_20945,N_18409,N_18105);
xnor U20946 (N_20946,N_18325,N_18290);
nor U20947 (N_20947,N_19382,N_19097);
or U20948 (N_20948,N_18137,N_19333);
or U20949 (N_20949,N_18961,N_19141);
xor U20950 (N_20950,N_18576,N_18729);
xnor U20951 (N_20951,N_18172,N_19031);
nor U20952 (N_20952,N_18069,N_18370);
nand U20953 (N_20953,N_19350,N_19102);
or U20954 (N_20954,N_18668,N_19328);
nor U20955 (N_20955,N_18493,N_18476);
xor U20956 (N_20956,N_18520,N_18330);
nor U20957 (N_20957,N_18924,N_19263);
and U20958 (N_20958,N_19381,N_18101);
and U20959 (N_20959,N_19219,N_18943);
and U20960 (N_20960,N_18131,N_19461);
nand U20961 (N_20961,N_18923,N_19225);
nor U20962 (N_20962,N_18214,N_19027);
nor U20963 (N_20963,N_18709,N_18601);
nor U20964 (N_20964,N_18278,N_19343);
or U20965 (N_20965,N_18103,N_18547);
xnor U20966 (N_20966,N_18506,N_19272);
nand U20967 (N_20967,N_18511,N_19055);
and U20968 (N_20968,N_18775,N_18443);
nor U20969 (N_20969,N_18182,N_18904);
and U20970 (N_20970,N_18844,N_18587);
xnor U20971 (N_20971,N_18336,N_18722);
nand U20972 (N_20972,N_19155,N_18066);
nor U20973 (N_20973,N_18332,N_18324);
nor U20974 (N_20974,N_18291,N_18606);
nor U20975 (N_20975,N_18069,N_19256);
nand U20976 (N_20976,N_18527,N_19063);
nand U20977 (N_20977,N_18994,N_18982);
nand U20978 (N_20978,N_18001,N_18280);
nand U20979 (N_20979,N_19353,N_18214);
xor U20980 (N_20980,N_19003,N_18467);
nor U20981 (N_20981,N_19473,N_19406);
and U20982 (N_20982,N_18666,N_18187);
and U20983 (N_20983,N_18609,N_19205);
and U20984 (N_20984,N_18853,N_19423);
and U20985 (N_20985,N_18822,N_19283);
and U20986 (N_20986,N_18239,N_18052);
or U20987 (N_20987,N_18751,N_18191);
nor U20988 (N_20988,N_18234,N_19368);
or U20989 (N_20989,N_19386,N_19277);
nor U20990 (N_20990,N_19122,N_18303);
and U20991 (N_20991,N_19117,N_18998);
xor U20992 (N_20992,N_19474,N_18501);
nor U20993 (N_20993,N_18357,N_19266);
xor U20994 (N_20994,N_18854,N_18449);
nand U20995 (N_20995,N_19084,N_18415);
nand U20996 (N_20996,N_19027,N_18370);
xnor U20997 (N_20997,N_18569,N_19239);
or U20998 (N_20998,N_18225,N_19156);
nand U20999 (N_20999,N_18988,N_18276);
or U21000 (N_21000,N_19966,N_19909);
and U21001 (N_21001,N_20219,N_20551);
nand U21002 (N_21002,N_19818,N_20559);
nand U21003 (N_21003,N_20063,N_20158);
nand U21004 (N_21004,N_19795,N_19689);
nor U21005 (N_21005,N_20879,N_20554);
and U21006 (N_21006,N_20250,N_20782);
and U21007 (N_21007,N_20701,N_20286);
nand U21008 (N_21008,N_20562,N_19581);
and U21009 (N_21009,N_20951,N_20118);
nor U21010 (N_21010,N_19666,N_20657);
and U21011 (N_21011,N_20536,N_20043);
and U21012 (N_21012,N_20626,N_19964);
xnor U21013 (N_21013,N_20045,N_20520);
or U21014 (N_21014,N_20647,N_20290);
nor U21015 (N_21015,N_19644,N_20304);
or U21016 (N_21016,N_20269,N_20732);
and U21017 (N_21017,N_19612,N_20104);
xor U21018 (N_21018,N_19529,N_19675);
nand U21019 (N_21019,N_19796,N_19955);
nand U21020 (N_21020,N_19989,N_20513);
nand U21021 (N_21021,N_19752,N_20548);
nor U21022 (N_21022,N_19789,N_20639);
xor U21023 (N_21023,N_20855,N_20524);
xnor U21024 (N_21024,N_20825,N_20744);
xor U21025 (N_21025,N_20653,N_20727);
or U21026 (N_21026,N_19533,N_20152);
xnor U21027 (N_21027,N_19972,N_20968);
xnor U21028 (N_21028,N_20083,N_20799);
and U21029 (N_21029,N_20365,N_20185);
nand U21030 (N_21030,N_20109,N_20485);
and U21031 (N_21031,N_20486,N_20511);
or U21032 (N_21032,N_20500,N_20635);
or U21033 (N_21033,N_20337,N_19862);
nand U21034 (N_21034,N_20489,N_19942);
nand U21035 (N_21035,N_20060,N_20357);
or U21036 (N_21036,N_20009,N_19518);
or U21037 (N_21037,N_20203,N_19803);
nand U21038 (N_21038,N_20106,N_19651);
xnor U21039 (N_21039,N_20863,N_19530);
xnor U21040 (N_21040,N_20595,N_20627);
or U21041 (N_21041,N_20521,N_20138);
nor U21042 (N_21042,N_20332,N_20920);
nand U21043 (N_21043,N_19608,N_20382);
xnor U21044 (N_21044,N_20765,N_20556);
or U21045 (N_21045,N_20044,N_20409);
xnor U21046 (N_21046,N_20102,N_20617);
and U21047 (N_21047,N_20945,N_20658);
and U21048 (N_21048,N_19591,N_20291);
nor U21049 (N_21049,N_20004,N_19606);
nor U21050 (N_21050,N_19549,N_19903);
or U21051 (N_21051,N_19978,N_20175);
or U21052 (N_21052,N_20070,N_19735);
nand U21053 (N_21053,N_20275,N_20887);
or U21054 (N_21054,N_20734,N_20006);
xnor U21055 (N_21055,N_20037,N_20475);
nand U21056 (N_21056,N_19917,N_20568);
or U21057 (N_21057,N_19805,N_19676);
or U21058 (N_21058,N_20469,N_19846);
nor U21059 (N_21059,N_20849,N_20592);
xnor U21060 (N_21060,N_20046,N_20088);
xor U21061 (N_21061,N_20430,N_19649);
or U21062 (N_21062,N_20114,N_20522);
or U21063 (N_21063,N_20764,N_20552);
nand U21064 (N_21064,N_20650,N_20867);
nand U21065 (N_21065,N_20735,N_19714);
xnor U21066 (N_21066,N_20420,N_19564);
or U21067 (N_21067,N_19703,N_20916);
xnor U21068 (N_21068,N_20501,N_19881);
xor U21069 (N_21069,N_19828,N_20610);
and U21070 (N_21070,N_19993,N_19965);
nand U21071 (N_21071,N_20050,N_20167);
or U21072 (N_21072,N_20053,N_19835);
nand U21073 (N_21073,N_19585,N_20597);
nor U21074 (N_21074,N_20515,N_19988);
or U21075 (N_21075,N_20832,N_19894);
xor U21076 (N_21076,N_19886,N_19624);
and U21077 (N_21077,N_20176,N_20582);
or U21078 (N_21078,N_20302,N_20202);
nand U21079 (N_21079,N_19815,N_19563);
nand U21080 (N_21080,N_20633,N_20504);
nor U21081 (N_21081,N_19844,N_20300);
or U21082 (N_21082,N_19641,N_19732);
nand U21083 (N_21083,N_20209,N_20233);
xor U21084 (N_21084,N_19670,N_20164);
xor U21085 (N_21085,N_20977,N_19901);
nor U21086 (N_21086,N_20819,N_20499);
nand U21087 (N_21087,N_20533,N_19587);
or U21088 (N_21088,N_20098,N_19938);
or U21089 (N_21089,N_19876,N_20605);
or U21090 (N_21090,N_20638,N_20681);
nand U21091 (N_21091,N_19939,N_20007);
nand U21092 (N_21092,N_20682,N_20367);
or U21093 (N_21093,N_20873,N_20204);
nor U21094 (N_21094,N_20231,N_20813);
and U21095 (N_21095,N_19838,N_20897);
xor U21096 (N_21096,N_20995,N_20343);
nand U21097 (N_21097,N_19990,N_20465);
or U21098 (N_21098,N_19584,N_19637);
nor U21099 (N_21099,N_19638,N_19706);
or U21100 (N_21100,N_19619,N_20924);
and U21101 (N_21101,N_20677,N_20205);
or U21102 (N_21102,N_20718,N_20604);
xnor U21103 (N_21103,N_20086,N_20576);
xor U21104 (N_21104,N_19571,N_20492);
or U21105 (N_21105,N_19793,N_20856);
xnor U21106 (N_21106,N_20493,N_20603);
nor U21107 (N_21107,N_19621,N_19946);
nor U21108 (N_21108,N_20170,N_20428);
and U21109 (N_21109,N_20122,N_20768);
and U21110 (N_21110,N_19614,N_20839);
or U21111 (N_21111,N_19761,N_20889);
and U21112 (N_21112,N_20966,N_19708);
or U21113 (N_21113,N_19842,N_20463);
nand U21114 (N_21114,N_19544,N_20229);
nand U21115 (N_21115,N_20666,N_20906);
nor U21116 (N_21116,N_19680,N_20422);
xnor U21117 (N_21117,N_20763,N_20611);
xor U21118 (N_21118,N_19896,N_19520);
xnor U21119 (N_21119,N_20704,N_20488);
and U21120 (N_21120,N_20079,N_20096);
nor U21121 (N_21121,N_19729,N_20184);
nor U21122 (N_21122,N_19888,N_19570);
or U21123 (N_21123,N_19932,N_20312);
nor U21124 (N_21124,N_20862,N_20441);
nor U21125 (N_21125,N_20890,N_20155);
nor U21126 (N_21126,N_19745,N_19987);
nand U21127 (N_21127,N_19500,N_20566);
nor U21128 (N_21128,N_19810,N_19702);
xor U21129 (N_21129,N_20431,N_20348);
nand U21130 (N_21130,N_20778,N_19884);
nor U21131 (N_21131,N_19879,N_19869);
and U21132 (N_21132,N_19904,N_20599);
or U21133 (N_21133,N_20539,N_19726);
xnor U21134 (N_21134,N_20543,N_19741);
and U21135 (N_21135,N_20243,N_20808);
nor U21136 (N_21136,N_20921,N_19860);
nand U21137 (N_21137,N_20035,N_20974);
or U21138 (N_21138,N_20391,N_19502);
and U21139 (N_21139,N_20115,N_20038);
xnor U21140 (N_21140,N_20609,N_20029);
xnor U21141 (N_21141,N_20905,N_20900);
and U21142 (N_21142,N_20917,N_20642);
nor U21143 (N_21143,N_20412,N_20178);
and U21144 (N_21144,N_20976,N_20589);
and U21145 (N_21145,N_20410,N_20301);
xor U21146 (N_21146,N_19858,N_19751);
and U21147 (N_21147,N_20885,N_19652);
or U21148 (N_21148,N_20117,N_20833);
or U21149 (N_21149,N_20777,N_20121);
xnor U21150 (N_21150,N_20452,N_20810);
xor U21151 (N_21151,N_20986,N_19687);
and U21152 (N_21152,N_20023,N_20816);
xor U21153 (N_21153,N_19753,N_20941);
xnor U21154 (N_21154,N_20895,N_20829);
xor U21155 (N_21155,N_20462,N_20450);
and U21156 (N_21156,N_20632,N_19770);
or U21157 (N_21157,N_20123,N_19690);
and U21158 (N_21158,N_20415,N_19885);
xnor U21159 (N_21159,N_20722,N_19738);
nand U21160 (N_21160,N_19593,N_19892);
and U21161 (N_21161,N_19731,N_20298);
nor U21162 (N_21162,N_20919,N_20600);
xnor U21163 (N_21163,N_20743,N_20996);
nand U21164 (N_21164,N_20481,N_20745);
xor U21165 (N_21165,N_19683,N_19850);
nor U21166 (N_21166,N_19613,N_20788);
and U21167 (N_21167,N_19669,N_19890);
and U21168 (N_21168,N_20324,N_20807);
nand U21169 (N_21169,N_20091,N_19820);
or U21170 (N_21170,N_20991,N_19656);
nor U21171 (N_21171,N_20378,N_20192);
xnor U21172 (N_21172,N_20623,N_19546);
or U21173 (N_21173,N_20072,N_20852);
xnor U21174 (N_21174,N_20326,N_19873);
or U21175 (N_21175,N_20308,N_20295);
xnor U21176 (N_21176,N_19566,N_19826);
xor U21177 (N_21177,N_20069,N_19711);
or U21178 (N_21178,N_20001,N_20094);
and U21179 (N_21179,N_20198,N_20311);
or U21180 (N_21180,N_20020,N_20442);
nand U21181 (N_21181,N_20015,N_20546);
nor U21182 (N_21182,N_20847,N_19762);
nor U21183 (N_21183,N_20396,N_19897);
nand U21184 (N_21184,N_19663,N_19986);
nor U21185 (N_21185,N_20097,N_19961);
xnor U21186 (N_21186,N_20055,N_19799);
or U21187 (N_21187,N_20937,N_19739);
and U21188 (N_21188,N_19562,N_20257);
nor U21189 (N_21189,N_20661,N_20160);
xnor U21190 (N_21190,N_20540,N_20956);
nand U21191 (N_21191,N_20297,N_20443);
nand U21192 (N_21192,N_20439,N_20436);
nor U21193 (N_21193,N_20981,N_19557);
xnor U21194 (N_21194,N_19539,N_20142);
and U21195 (N_21195,N_19664,N_20588);
or U21196 (N_21196,N_20421,N_20861);
or U21197 (N_21197,N_19999,N_20684);
xor U21198 (N_21198,N_19588,N_20509);
or U21199 (N_21199,N_20717,N_20387);
nor U21200 (N_21200,N_20621,N_20831);
or U21201 (N_21201,N_19697,N_20624);
and U21202 (N_21202,N_20418,N_20051);
xor U21203 (N_21203,N_20779,N_20282);
nor U21204 (N_21204,N_20584,N_20569);
or U21205 (N_21205,N_20914,N_20187);
nand U21206 (N_21206,N_20542,N_20695);
nor U21207 (N_21207,N_19535,N_20003);
nor U21208 (N_21208,N_19742,N_19540);
and U21209 (N_21209,N_20135,N_20911);
and U21210 (N_21210,N_19740,N_19945);
or U21211 (N_21211,N_20320,N_20190);
nand U21212 (N_21212,N_20802,N_20375);
xnor U21213 (N_21213,N_20416,N_19684);
nand U21214 (N_21214,N_19537,N_19692);
xor U21215 (N_21215,N_20640,N_20608);
and U21216 (N_21216,N_19596,N_20830);
and U21217 (N_21217,N_19808,N_20712);
nand U21218 (N_21218,N_19715,N_20634);
nand U21219 (N_21219,N_20822,N_19699);
and U21220 (N_21220,N_19506,N_19766);
or U21221 (N_21221,N_20517,N_20703);
and U21222 (N_21222,N_19620,N_20793);
or U21223 (N_21223,N_20893,N_20739);
xnor U21224 (N_21224,N_20494,N_20074);
nor U21225 (N_21225,N_19893,N_19594);
nand U21226 (N_21226,N_19730,N_19548);
xor U21227 (N_21227,N_20179,N_20093);
or U21228 (N_21228,N_19630,N_20618);
nand U21229 (N_21229,N_19908,N_19545);
nor U21230 (N_21230,N_20721,N_20913);
nand U21231 (N_21231,N_19686,N_20265);
nor U21232 (N_21232,N_19800,N_20244);
nor U21233 (N_21233,N_19734,N_20750);
and U21234 (N_21234,N_20273,N_20838);
or U21235 (N_21235,N_20468,N_20678);
or U21236 (N_21236,N_20570,N_20528);
and U21237 (N_21237,N_19700,N_20221);
xnor U21238 (N_21238,N_20947,N_20978);
nor U21239 (N_21239,N_19722,N_19604);
nand U21240 (N_21240,N_19723,N_19754);
nor U21241 (N_21241,N_20859,N_20218);
nand U21242 (N_21242,N_19555,N_19509);
xnor U21243 (N_21243,N_19511,N_20261);
or U21244 (N_21244,N_20456,N_20054);
or U21245 (N_21245,N_19919,N_20958);
nand U21246 (N_21246,N_19528,N_19671);
nor U21247 (N_21247,N_20168,N_20449);
nand U21248 (N_21248,N_19611,N_20502);
nor U21249 (N_21249,N_19995,N_19553);
or U21250 (N_21250,N_20362,N_20025);
xnor U21251 (N_21251,N_20159,N_20200);
nand U21252 (N_21252,N_20547,N_20724);
nand U21253 (N_21253,N_20406,N_20903);
and U21254 (N_21254,N_19954,N_20398);
nand U21255 (N_21255,N_19646,N_20136);
nor U21256 (N_21256,N_19554,N_19940);
or U21257 (N_21257,N_19532,N_20073);
xor U21258 (N_21258,N_20674,N_19821);
nand U21259 (N_21259,N_19824,N_19625);
nand U21260 (N_21260,N_20791,N_19543);
nand U21261 (N_21261,N_20157,N_20034);
nor U21262 (N_21262,N_20596,N_19707);
xor U21263 (N_21263,N_20153,N_19759);
xor U21264 (N_21264,N_20130,N_20815);
nand U21265 (N_21265,N_19633,N_20289);
nand U21266 (N_21266,N_19960,N_19781);
xor U21267 (N_21267,N_20383,N_20884);
xor U21268 (N_21268,N_20390,N_20961);
nand U21269 (N_21269,N_20898,N_20834);
xnor U21270 (N_21270,N_20821,N_19602);
nand U21271 (N_21271,N_20933,N_20005);
and U21272 (N_21272,N_19765,N_20564);
nand U21273 (N_21273,N_20993,N_20189);
nand U21274 (N_21274,N_19631,N_19550);
xor U21275 (N_21275,N_20555,N_20835);
xnor U21276 (N_21276,N_19950,N_19639);
and U21277 (N_21277,N_19867,N_20534);
nand U21278 (N_21278,N_20369,N_20665);
xnor U21279 (N_21279,N_20953,N_20236);
xnor U21280 (N_21280,N_20655,N_19949);
nand U21281 (N_21281,N_20644,N_20801);
and U21282 (N_21282,N_20535,N_19769);
xnor U21283 (N_21283,N_20972,N_20028);
or U21284 (N_21284,N_19512,N_20201);
xor U21285 (N_21285,N_19616,N_20707);
and U21286 (N_21286,N_19837,N_19601);
nor U21287 (N_21287,N_20258,N_20846);
xnor U21288 (N_21288,N_19527,N_20111);
nand U21289 (N_21289,N_19674,N_20886);
nand U21290 (N_21290,N_20419,N_20907);
nor U21291 (N_21291,N_20141,N_20030);
and U21292 (N_21292,N_19609,N_20561);
nor U21293 (N_21293,N_20692,N_20228);
or U21294 (N_21294,N_20918,N_19979);
xnor U21295 (N_21295,N_19748,N_20466);
and U21296 (N_21296,N_19851,N_19777);
or U21297 (N_21297,N_20973,N_19970);
nor U21298 (N_21298,N_19763,N_20246);
nand U21299 (N_21299,N_19559,N_20950);
nor U21300 (N_21300,N_20663,N_20997);
nand U21301 (N_21301,N_20759,N_20414);
or U21302 (N_21302,N_19561,N_20042);
xor U21303 (N_21303,N_20370,N_20685);
xor U21304 (N_21304,N_20649,N_19819);
nor U21305 (N_21305,N_19757,N_20374);
xnor U21306 (N_21306,N_20110,N_19785);
and U21307 (N_21307,N_20773,N_19573);
nand U21308 (N_21308,N_20532,N_20222);
xnor U21309 (N_21309,N_19900,N_20591);
nand U21310 (N_21310,N_20057,N_20150);
and U21311 (N_21311,N_19934,N_20388);
or U21312 (N_21312,N_20938,N_20350);
and U21313 (N_21313,N_19576,N_20758);
nor U21314 (N_21314,N_19541,N_20713);
nand U21315 (N_21315,N_19503,N_20964);
or U21316 (N_21316,N_20751,N_19967);
nor U21317 (N_21317,N_20319,N_19716);
xnor U21318 (N_21318,N_19538,N_19635);
nand U21319 (N_21319,N_20689,N_20746);
xnor U21320 (N_21320,N_20901,N_20676);
nor U21321 (N_21321,N_20059,N_19992);
nand U21322 (N_21322,N_20241,N_20989);
nor U21323 (N_21323,N_20785,N_20165);
nor U21324 (N_21324,N_19957,N_20174);
nand U21325 (N_21325,N_20162,N_19727);
or U21326 (N_21326,N_19848,N_19774);
nor U21327 (N_21327,N_19705,N_20602);
nor U21328 (N_21328,N_20939,N_20352);
xor U21329 (N_21329,N_20823,N_19840);
nand U21330 (N_21330,N_20393,N_20427);
and U21331 (N_21331,N_20770,N_19918);
and U21332 (N_21332,N_20929,N_20593);
xor U21333 (N_21333,N_20127,N_20954);
and U21334 (N_21334,N_19660,N_20081);
xnor U21335 (N_21335,N_20256,N_19627);
or U21336 (N_21336,N_20235,N_20446);
or U21337 (N_21337,N_20423,N_20748);
and U21338 (N_21338,N_20180,N_20811);
nand U21339 (N_21339,N_20963,N_20537);
and U21340 (N_21340,N_20875,N_19760);
xor U21341 (N_21341,N_20659,N_20310);
nand U21342 (N_21342,N_20720,N_20182);
or U21343 (N_21343,N_19650,N_19586);
nor U21344 (N_21344,N_20287,N_19750);
nand U21345 (N_21345,N_19605,N_20840);
nand U21346 (N_21346,N_19784,N_19704);
nor U21347 (N_21347,N_19944,N_20022);
nand U21348 (N_21348,N_20143,N_20550);
xnor U21349 (N_21349,N_19994,N_20095);
and U21350 (N_21350,N_19685,N_20698);
and U21351 (N_21351,N_19975,N_19825);
nor U21352 (N_21352,N_20379,N_19985);
nor U21353 (N_21353,N_20648,N_20844);
and U21354 (N_21354,N_19984,N_20480);
or U21355 (N_21355,N_20353,N_20670);
nand U21356 (N_21356,N_20266,N_20132);
and U21357 (N_21357,N_20014,N_20786);
nor U21358 (N_21358,N_20908,N_20740);
nand U21359 (N_21359,N_20498,N_20538);
and U21360 (N_21360,N_20899,N_20339);
and U21361 (N_21361,N_20281,N_20223);
xor U21362 (N_21362,N_20573,N_20694);
nand U21363 (N_21363,N_20460,N_20395);
xnor U21364 (N_21364,N_20103,N_19952);
or U21365 (N_21365,N_19556,N_19854);
and U21366 (N_21366,N_20870,N_19929);
nor U21367 (N_21367,N_20242,N_19580);
and U21368 (N_21368,N_20679,N_19839);
nand U21369 (N_21369,N_19578,N_20195);
xor U21370 (N_21370,N_20868,N_19899);
nand U21371 (N_21371,N_20651,N_20331);
nand U21372 (N_21372,N_20299,N_20140);
or U21373 (N_21373,N_19636,N_19673);
nor U21374 (N_21374,N_20757,N_20214);
or U21375 (N_21375,N_20686,N_20262);
nand U21376 (N_21376,N_19875,N_20514);
or U21377 (N_21377,N_19654,N_20667);
xor U21378 (N_21378,N_19859,N_20448);
nand U21379 (N_21379,N_19951,N_20212);
and U21380 (N_21380,N_20809,N_19747);
or U21381 (N_21381,N_19688,N_20148);
nand U21382 (N_21382,N_20172,N_20307);
or U21383 (N_21383,N_20078,N_20615);
nand U21384 (N_21384,N_20668,N_20904);
or U21385 (N_21385,N_19780,N_20248);
xnor U21386 (N_21386,N_20737,N_20417);
xor U21387 (N_21387,N_20245,N_20373);
xor U21388 (N_21388,N_20206,N_19640);
and U21389 (N_21389,N_20936,N_20794);
xnor U21390 (N_21390,N_20392,N_20891);
nand U21391 (N_21391,N_20032,N_19790);
nand U21392 (N_21392,N_20129,N_20725);
nor U21393 (N_21393,N_19720,N_20193);
xor U21394 (N_21394,N_20285,N_19870);
and U21395 (N_21395,N_20268,N_20560);
or U21396 (N_21396,N_20173,N_20454);
nor U21397 (N_21397,N_20013,N_19693);
xnor U21398 (N_21398,N_20702,N_20518);
nand U21399 (N_21399,N_19921,N_20935);
xnor U21400 (N_21400,N_20896,N_20333);
and U21401 (N_21401,N_19567,N_19816);
nand U21402 (N_21402,N_19982,N_20487);
and U21403 (N_21403,N_19749,N_19515);
and U21404 (N_21404,N_20804,N_19665);
or U21405 (N_21405,N_20781,N_20280);
and U21406 (N_21406,N_20544,N_19926);
or U21407 (N_21407,N_20836,N_20571);
xnor U21408 (N_21408,N_20614,N_20878);
and U21409 (N_21409,N_20747,N_20065);
xnor U21410 (N_21410,N_20181,N_19632);
or U21411 (N_21411,N_20578,N_20161);
xnor U21412 (N_21412,N_20402,N_19628);
and U21413 (N_21413,N_19600,N_19871);
or U21414 (N_21414,N_19504,N_20426);
xor U21415 (N_21415,N_20824,N_20076);
or U21416 (N_21416,N_20048,N_20928);
xnor U21417 (N_21417,N_20820,N_20075);
xor U21418 (N_21418,N_20817,N_20372);
or U21419 (N_21419,N_20199,N_19983);
and U21420 (N_21420,N_19958,N_19746);
xor U21421 (N_21421,N_20220,N_19874);
or U21422 (N_21422,N_19798,N_19809);
and U21423 (N_21423,N_19768,N_20283);
or U21424 (N_21424,N_19657,N_20344);
or U21425 (N_21425,N_20771,N_20309);
and U21426 (N_21426,N_19531,N_19930);
nand U21427 (N_21427,N_20407,N_19889);
nand U21428 (N_21428,N_20645,N_19920);
and U21429 (N_21429,N_20687,N_20024);
nand U21430 (N_21430,N_20858,N_19510);
or U21431 (N_21431,N_20590,N_20349);
or U21432 (N_21432,N_20188,N_20960);
and U21433 (N_21433,N_20252,N_19565);
and U21434 (N_21434,N_20041,N_20116);
and U21435 (N_21435,N_20026,N_20361);
xnor U21436 (N_21436,N_20139,N_20982);
nand U21437 (N_21437,N_19887,N_20505);
xnor U21438 (N_21438,N_20728,N_19925);
nand U21439 (N_21439,N_20691,N_20545);
or U21440 (N_21440,N_19667,N_20549);
xnor U21441 (N_21441,N_20031,N_20798);
or U21442 (N_21442,N_19823,N_20381);
nor U21443 (N_21443,N_19943,N_19607);
nor U21444 (N_21444,N_19836,N_20039);
xnor U21445 (N_21445,N_20384,N_19857);
nand U21446 (N_21446,N_20107,N_19847);
and U21447 (N_21447,N_20479,N_20985);
xnor U21448 (N_21448,N_20292,N_20008);
nor U21449 (N_21449,N_20894,N_19880);
or U21450 (N_21450,N_20806,N_20965);
and U21451 (N_21451,N_20437,N_20455);
or U21452 (N_21452,N_20249,N_20071);
and U21453 (N_21453,N_19572,N_20323);
or U21454 (N_21454,N_19797,N_19634);
nor U21455 (N_21455,N_20359,N_19976);
or U21456 (N_21456,N_20775,N_19791);
and U21457 (N_21457,N_20021,N_20967);
nand U21458 (N_21458,N_20092,N_20510);
nor U21459 (N_21459,N_19782,N_20880);
nand U21460 (N_21460,N_20338,N_19691);
nand U21461 (N_21461,N_20058,N_20210);
xnor U21462 (N_21462,N_19913,N_19744);
and U21463 (N_21463,N_20983,N_20272);
and U21464 (N_21464,N_19813,N_19931);
and U21465 (N_21465,N_19872,N_20910);
xor U21466 (N_21466,N_20277,N_20567);
or U21467 (N_21467,N_19804,N_19682);
or U21468 (N_21468,N_19902,N_20738);
nand U21469 (N_21469,N_19807,N_20099);
nor U21470 (N_21470,N_20151,N_20408);
and U21471 (N_21471,N_19802,N_19598);
nand U21472 (N_21472,N_20087,N_19536);
nand U21473 (N_21473,N_20010,N_20656);
nand U21474 (N_21474,N_19912,N_20563);
nor U21475 (N_21475,N_20274,N_19615);
and U21476 (N_21476,N_19696,N_20607);
xnor U21477 (N_21477,N_20356,N_20169);
nor U21478 (N_21478,N_20998,N_19721);
xor U21479 (N_21479,N_20660,N_20496);
and U21480 (N_21480,N_20413,N_20680);
and U21481 (N_21481,N_20512,N_20346);
and U21482 (N_21482,N_20263,N_19834);
xnor U21483 (N_21483,N_19679,N_20753);
xnor U21484 (N_21484,N_20011,N_19560);
xnor U21485 (N_21485,N_20191,N_19855);
and U21486 (N_21486,N_19891,N_20119);
nand U21487 (N_21487,N_20226,N_20690);
xor U21488 (N_21488,N_20137,N_20363);
or U21489 (N_21489,N_19589,N_19622);
and U21490 (N_21490,N_19776,N_19668);
or U21491 (N_21491,N_20865,N_20495);
nor U21492 (N_21492,N_20519,N_20368);
xor U21493 (N_21493,N_20224,N_19883);
nand U21494 (N_21494,N_19724,N_20012);
nand U21495 (N_21495,N_19928,N_20787);
nor U21496 (N_21496,N_19778,N_19662);
nor U21497 (N_21497,N_20577,N_20800);
and U21498 (N_21498,N_20927,N_20587);
or U21499 (N_21499,N_20636,N_20047);
xnor U21500 (N_21500,N_20756,N_19787);
and U21501 (N_21501,N_19599,N_20783);
xor U21502 (N_21502,N_20328,N_19980);
or U21503 (N_21503,N_19517,N_19969);
nand U21504 (N_21504,N_20061,N_20451);
and U21505 (N_21505,N_20062,N_19534);
or U21506 (N_21506,N_20579,N_20124);
nor U21507 (N_21507,N_20818,N_19956);
xor U21508 (N_21508,N_20774,N_20795);
nand U21509 (N_21509,N_19648,N_20016);
nor U21510 (N_21510,N_19907,N_20149);
nor U21511 (N_21511,N_20325,N_20729);
and U21512 (N_21512,N_20260,N_19806);
xor U21513 (N_21513,N_20002,N_19525);
or U21514 (N_21514,N_20944,N_20719);
nand U21515 (N_21515,N_20380,N_19779);
or U21516 (N_21516,N_20888,N_20902);
nor U21517 (N_21517,N_20276,N_19658);
xnor U21518 (N_21518,N_19756,N_20789);
xnor U21519 (N_21519,N_19953,N_20217);
and U21520 (N_21520,N_19629,N_20464);
nand U21521 (N_21521,N_20503,N_19856);
nor U21522 (N_21522,N_20733,N_20238);
nor U21523 (N_21523,N_20476,N_20754);
or U21524 (N_21524,N_20612,N_20812);
and U21525 (N_21525,N_20447,N_20864);
or U21526 (N_21526,N_20558,N_20459);
nand U21527 (N_21527,N_19643,N_20952);
nand U21528 (N_21528,N_20270,N_20970);
xor U21529 (N_21529,N_20523,N_20874);
nor U21530 (N_21530,N_20438,N_19569);
xor U21531 (N_21531,N_20697,N_19597);
nor U21532 (N_21532,N_20208,N_20303);
nor U21533 (N_21533,N_20869,N_20400);
and U21534 (N_21534,N_19941,N_19733);
nor U21535 (N_21535,N_20761,N_20925);
nand U21536 (N_21536,N_19814,N_20036);
and U21537 (N_21537,N_20581,N_20156);
and U21538 (N_21538,N_20336,N_20335);
or U21539 (N_21539,N_19962,N_19959);
and U21540 (N_21540,N_20876,N_20403);
xor U21541 (N_21541,N_19677,N_20067);
nand U21542 (N_21542,N_20033,N_20313);
and U21543 (N_21543,N_19653,N_20749);
nor U21544 (N_21544,N_19737,N_20445);
and U21545 (N_21545,N_20622,N_20483);
nor U21546 (N_21546,N_19701,N_19817);
or U21547 (N_21547,N_20068,N_19542);
or U21548 (N_21548,N_19717,N_20527);
or U21549 (N_21549,N_20969,N_19725);
or U21550 (N_21550,N_20457,N_20017);
nand U21551 (N_21551,N_19575,N_19694);
or U21552 (N_21552,N_19830,N_20284);
nor U21553 (N_21553,N_19878,N_20959);
or U21554 (N_21554,N_20988,N_20772);
or U21555 (N_21555,N_20146,N_20850);
or U21556 (N_21556,N_20101,N_20955);
and U21557 (N_21557,N_20018,N_20296);
or U21558 (N_21558,N_20125,N_20341);
xor U21559 (N_21559,N_20715,N_20731);
or U21560 (N_21560,N_20848,N_19968);
nand U21561 (N_21561,N_20696,N_19853);
xor U21562 (N_21562,N_20987,N_20842);
or U21563 (N_21563,N_20672,N_19516);
xnor U21564 (N_21564,N_20113,N_19501);
xor U21565 (N_21565,N_19863,N_20726);
xor U21566 (N_21566,N_20979,N_20232);
or U21567 (N_21567,N_20932,N_19914);
nor U21568 (N_21568,N_19743,N_20253);
or U21569 (N_21569,N_20797,N_20664);
xor U21570 (N_21570,N_20723,N_19645);
and U21571 (N_21571,N_20131,N_20377);
and U21572 (N_21572,N_20760,N_19882);
and U21573 (N_21573,N_20112,N_19568);
nor U21574 (N_21574,N_20145,N_20949);
nand U21575 (N_21575,N_20405,N_20315);
xnor U21576 (N_21576,N_19864,N_20183);
and U21577 (N_21577,N_20683,N_19558);
xor U21578 (N_21578,N_20946,N_19861);
nand U21579 (N_21579,N_20334,N_19574);
and U21580 (N_21580,N_20166,N_20688);
nand U21581 (N_21581,N_19603,N_20355);
or U21582 (N_21582,N_19521,N_19583);
and U21583 (N_21583,N_20803,N_20052);
xnor U21584 (N_21584,N_20490,N_20147);
and U21585 (N_21585,N_19811,N_19905);
and U21586 (N_21586,N_20586,N_20999);
and U21587 (N_21587,N_19911,N_19590);
and U21588 (N_21588,N_19552,N_20752);
xor U21589 (N_21589,N_19832,N_20837);
and U21590 (N_21590,N_20598,N_20931);
nand U21591 (N_21591,N_20128,N_20766);
nand U21592 (N_21592,N_20019,N_20557);
nand U21593 (N_21593,N_20671,N_19996);
and U21594 (N_21594,N_19868,N_20213);
and U21595 (N_21595,N_19719,N_20971);
xnor U21596 (N_21596,N_19822,N_20484);
or U21597 (N_21597,N_20251,N_20706);
nor U21598 (N_21598,N_20458,N_20574);
nor U21599 (N_21599,N_20240,N_19963);
xnor U21600 (N_21600,N_20705,N_19998);
nand U21601 (N_21601,N_20444,N_19915);
and U21602 (N_21602,N_19523,N_20585);
or U21603 (N_21603,N_20980,N_20089);
nor U21604 (N_21604,N_20389,N_20892);
and U21605 (N_21605,N_20975,N_20401);
nor U21606 (N_21606,N_19801,N_19712);
or U21607 (N_21607,N_20144,N_20227);
nand U21608 (N_21608,N_19519,N_20371);
nand U21609 (N_21609,N_19623,N_19845);
and U21610 (N_21610,N_20853,N_20435);
xor U21611 (N_21611,N_19526,N_19618);
xnor U21612 (N_21612,N_20606,N_20990);
nor U21613 (N_21613,N_20366,N_19947);
nor U21614 (N_21614,N_20860,N_20317);
nor U21615 (N_21615,N_20472,N_19661);
nand U21616 (N_21616,N_20133,N_20742);
nor U21617 (N_21617,N_19514,N_20186);
nor U21618 (N_21618,N_20620,N_20628);
and U21619 (N_21619,N_20805,N_20049);
or U21620 (N_21620,N_20425,N_19937);
and U21621 (N_21621,N_20082,N_20957);
nor U21622 (N_21622,N_19865,N_19595);
and U21623 (N_21623,N_20216,N_20424);
nor U21624 (N_21624,N_20327,N_20108);
nand U21625 (N_21625,N_20040,N_20854);
or U21626 (N_21626,N_20883,N_20525);
or U21627 (N_21627,N_19659,N_19710);
nor U21628 (N_21628,N_19933,N_19786);
and U21629 (N_21629,N_20594,N_20473);
nor U21630 (N_21630,N_19577,N_20741);
and U21631 (N_21631,N_20294,N_19977);
and U21632 (N_21632,N_19916,N_20234);
and U21633 (N_21633,N_19681,N_20776);
nand U21634 (N_21634,N_20826,N_20432);
xnor U21635 (N_21635,N_19898,N_20619);
and U21636 (N_21636,N_20279,N_20736);
nand U21637 (N_21637,N_19642,N_19507);
xnor U21638 (N_21638,N_20293,N_20474);
nor U21639 (N_21639,N_19758,N_20580);
or U21640 (N_21640,N_20271,N_19579);
xor U21641 (N_21641,N_20278,N_20508);
or U21642 (N_21642,N_20767,N_20881);
nor U21643 (N_21643,N_19866,N_20364);
xnor U21644 (N_21644,N_20434,N_20716);
nand U21645 (N_21645,N_20654,N_20652);
nor U21646 (N_21646,N_20411,N_20267);
and U21647 (N_21647,N_20247,N_20877);
nor U21648 (N_21648,N_20616,N_20530);
nor U21649 (N_21649,N_20948,N_20064);
xnor U21650 (N_21650,N_20675,N_19672);
nand U21651 (N_21651,N_19626,N_19764);
nand U21652 (N_21652,N_20828,N_19841);
or U21653 (N_21653,N_19678,N_20711);
nand U21654 (N_21654,N_20843,N_20814);
or U21655 (N_21655,N_20796,N_20673);
and U21656 (N_21656,N_19713,N_19829);
nor U21657 (N_21657,N_20077,N_20909);
nand U21658 (N_21658,N_20497,N_19792);
nand U21659 (N_21659,N_20306,N_19906);
or U21660 (N_21660,N_20386,N_20940);
or U21661 (N_21661,N_20662,N_19582);
and U21662 (N_21662,N_19877,N_19610);
nor U21663 (N_21663,N_20066,N_20641);
xor U21664 (N_21664,N_20329,N_20871);
nand U21665 (N_21665,N_20553,N_20316);
nand U21666 (N_21666,N_19522,N_19849);
or U21667 (N_21667,N_20330,N_20942);
and U21668 (N_21668,N_19997,N_19647);
xor U21669 (N_21669,N_20376,N_19772);
nor U21670 (N_21670,N_20482,N_20347);
xnor U21671 (N_21671,N_20477,N_20340);
nor U21672 (N_21672,N_20507,N_20399);
and U21673 (N_21673,N_19794,N_19617);
or U21674 (N_21674,N_20934,N_19736);
or U21675 (N_21675,N_20453,N_20994);
xnor U21676 (N_21676,N_20429,N_20467);
nor U21677 (N_21677,N_20478,N_20237);
nor U21678 (N_21678,N_20780,N_19973);
and U21679 (N_21679,N_20882,N_20541);
nor U21680 (N_21680,N_20404,N_20926);
xnor U21681 (N_21681,N_20572,N_19695);
nand U21682 (N_21682,N_19788,N_20631);
and U21683 (N_21683,N_19910,N_20930);
nand U21684 (N_21684,N_20625,N_20962);
or U21685 (N_21685,N_20714,N_20239);
xor U21686 (N_21686,N_19827,N_20710);
and U21687 (N_21687,N_20084,N_20196);
and U21688 (N_21688,N_20085,N_19923);
and U21689 (N_21689,N_20915,N_20526);
nand U21690 (N_21690,N_20090,N_20851);
or U21691 (N_21691,N_20360,N_19655);
or U21692 (N_21692,N_20197,N_19895);
nand U21693 (N_21693,N_20637,N_19547);
or U21694 (N_21694,N_19936,N_19922);
xor U21695 (N_21695,N_19843,N_20461);
nand U21696 (N_21696,N_20984,N_20943);
nor U21697 (N_21697,N_20358,N_20565);
or U21698 (N_21698,N_20194,N_20120);
xor U21699 (N_21699,N_20385,N_19551);
and U21700 (N_21700,N_20769,N_20255);
or U21701 (N_21701,N_20215,N_20629);
nor U21702 (N_21702,N_19831,N_20321);
nor U21703 (N_21703,N_19924,N_20700);
xnor U21704 (N_21704,N_19833,N_19783);
or U21705 (N_21705,N_20531,N_20643);
and U21706 (N_21706,N_19991,N_19771);
nor U21707 (N_21707,N_20646,N_20992);
or U21708 (N_21708,N_19773,N_19508);
nor U21709 (N_21709,N_19718,N_20506);
or U21710 (N_21710,N_20105,N_20730);
xor U21711 (N_21711,N_20230,N_19948);
and U21712 (N_21712,N_19505,N_20207);
nor U21713 (N_21713,N_20351,N_20693);
nor U21714 (N_21714,N_20314,N_20318);
and U21715 (N_21715,N_19935,N_20669);
nand U21716 (N_21716,N_20211,N_19852);
nor U21717 (N_21717,N_20177,N_20923);
and U21718 (N_21718,N_19927,N_20471);
or U21719 (N_21719,N_20254,N_20583);
xnor U21720 (N_21720,N_20171,N_20784);
or U21721 (N_21721,N_19698,N_20912);
and U21722 (N_21722,N_20305,N_20529);
xnor U21723 (N_21723,N_20790,N_20699);
nand U21724 (N_21724,N_20288,N_20100);
xnor U21725 (N_21725,N_20433,N_20259);
nor U21726 (N_21726,N_19755,N_19524);
or U21727 (N_21727,N_20575,N_19709);
xnor U21728 (N_21728,N_19971,N_20709);
xnor U21729 (N_21729,N_20345,N_19592);
xnor U21730 (N_21730,N_20516,N_19767);
nand U21731 (N_21731,N_20225,N_20708);
and U21732 (N_21732,N_20755,N_20000);
xnor U21733 (N_21733,N_20354,N_20126);
nor U21734 (N_21734,N_19513,N_19728);
xnor U21735 (N_21735,N_19981,N_20027);
xor U21736 (N_21736,N_20163,N_20827);
nand U21737 (N_21737,N_20922,N_20056);
xor U21738 (N_21738,N_20841,N_20080);
nand U21739 (N_21739,N_20872,N_20792);
or U21740 (N_21740,N_19974,N_20762);
nand U21741 (N_21741,N_20845,N_20866);
xnor U21742 (N_21742,N_20134,N_20397);
nor U21743 (N_21743,N_20440,N_20154);
xor U21744 (N_21744,N_20491,N_20322);
xnor U21745 (N_21745,N_20630,N_19812);
nor U21746 (N_21746,N_20613,N_20394);
nor U21747 (N_21747,N_19775,N_20264);
xor U21748 (N_21748,N_20601,N_20857);
nor U21749 (N_21749,N_20470,N_20342);
xor U21750 (N_21750,N_20249,N_19723);
and U21751 (N_21751,N_20155,N_20827);
nand U21752 (N_21752,N_20695,N_19579);
and U21753 (N_21753,N_19902,N_20327);
xor U21754 (N_21754,N_19863,N_19589);
nand U21755 (N_21755,N_20840,N_20269);
nor U21756 (N_21756,N_20574,N_20644);
nor U21757 (N_21757,N_20067,N_20704);
xor U21758 (N_21758,N_19705,N_20392);
nor U21759 (N_21759,N_19757,N_20686);
xor U21760 (N_21760,N_20474,N_19910);
nor U21761 (N_21761,N_20711,N_20053);
or U21762 (N_21762,N_19919,N_19762);
or U21763 (N_21763,N_20537,N_20150);
nor U21764 (N_21764,N_20301,N_20920);
nand U21765 (N_21765,N_20790,N_20752);
nand U21766 (N_21766,N_19891,N_20552);
and U21767 (N_21767,N_20355,N_20554);
or U21768 (N_21768,N_20263,N_19919);
nand U21769 (N_21769,N_20608,N_20994);
and U21770 (N_21770,N_20710,N_20086);
nor U21771 (N_21771,N_19988,N_20301);
nor U21772 (N_21772,N_20922,N_20036);
nand U21773 (N_21773,N_20380,N_19872);
nand U21774 (N_21774,N_20962,N_20585);
nor U21775 (N_21775,N_19918,N_20329);
or U21776 (N_21776,N_20344,N_19993);
xnor U21777 (N_21777,N_20312,N_19727);
nand U21778 (N_21778,N_20015,N_20792);
nor U21779 (N_21779,N_19996,N_20749);
nand U21780 (N_21780,N_20826,N_19790);
xnor U21781 (N_21781,N_20271,N_19680);
nand U21782 (N_21782,N_20885,N_19771);
or U21783 (N_21783,N_20034,N_19871);
or U21784 (N_21784,N_20542,N_19825);
and U21785 (N_21785,N_19628,N_20450);
xor U21786 (N_21786,N_20998,N_20073);
nand U21787 (N_21787,N_19578,N_20093);
and U21788 (N_21788,N_20701,N_20614);
nor U21789 (N_21789,N_20499,N_19999);
and U21790 (N_21790,N_19915,N_19627);
nor U21791 (N_21791,N_20974,N_20378);
nand U21792 (N_21792,N_19877,N_20971);
nand U21793 (N_21793,N_20897,N_20214);
nand U21794 (N_21794,N_20720,N_20866);
nand U21795 (N_21795,N_20268,N_20871);
xnor U21796 (N_21796,N_19772,N_20411);
nor U21797 (N_21797,N_20025,N_20737);
nor U21798 (N_21798,N_20543,N_19579);
or U21799 (N_21799,N_19773,N_19671);
xnor U21800 (N_21800,N_19801,N_19825);
and U21801 (N_21801,N_19996,N_20318);
and U21802 (N_21802,N_20764,N_20054);
and U21803 (N_21803,N_20977,N_19519);
xor U21804 (N_21804,N_20637,N_20476);
or U21805 (N_21805,N_20245,N_20344);
nand U21806 (N_21806,N_20800,N_20771);
or U21807 (N_21807,N_19597,N_20712);
nor U21808 (N_21808,N_20353,N_20916);
and U21809 (N_21809,N_19882,N_20982);
nor U21810 (N_21810,N_20834,N_19981);
and U21811 (N_21811,N_19597,N_20045);
nand U21812 (N_21812,N_19743,N_19990);
nor U21813 (N_21813,N_19691,N_19897);
and U21814 (N_21814,N_19754,N_20623);
xnor U21815 (N_21815,N_20509,N_20082);
nor U21816 (N_21816,N_20696,N_20326);
or U21817 (N_21817,N_19966,N_20753);
nand U21818 (N_21818,N_19719,N_20724);
xnor U21819 (N_21819,N_19983,N_19820);
nand U21820 (N_21820,N_19971,N_20433);
and U21821 (N_21821,N_19890,N_19856);
and U21822 (N_21822,N_19898,N_20810);
xor U21823 (N_21823,N_19998,N_20850);
nor U21824 (N_21824,N_19944,N_19739);
nor U21825 (N_21825,N_20577,N_19595);
nand U21826 (N_21826,N_20394,N_20452);
nand U21827 (N_21827,N_20558,N_19641);
and U21828 (N_21828,N_20698,N_19589);
and U21829 (N_21829,N_20727,N_20235);
and U21830 (N_21830,N_20431,N_20805);
nor U21831 (N_21831,N_20534,N_20583);
nor U21832 (N_21832,N_20327,N_20763);
nor U21833 (N_21833,N_20854,N_20152);
or U21834 (N_21834,N_20179,N_20990);
nand U21835 (N_21835,N_20361,N_20908);
xnor U21836 (N_21836,N_20086,N_20784);
xor U21837 (N_21837,N_20767,N_19758);
or U21838 (N_21838,N_19933,N_20224);
nor U21839 (N_21839,N_20974,N_20781);
and U21840 (N_21840,N_19855,N_20418);
nand U21841 (N_21841,N_19944,N_19748);
nand U21842 (N_21842,N_19982,N_20338);
nor U21843 (N_21843,N_20373,N_20763);
or U21844 (N_21844,N_20752,N_20649);
nor U21845 (N_21845,N_20397,N_20075);
nor U21846 (N_21846,N_20446,N_20290);
nand U21847 (N_21847,N_19976,N_19842);
and U21848 (N_21848,N_20932,N_19506);
nand U21849 (N_21849,N_20294,N_19545);
or U21850 (N_21850,N_19989,N_20274);
or U21851 (N_21851,N_19785,N_20686);
xor U21852 (N_21852,N_20935,N_20553);
xor U21853 (N_21853,N_20108,N_20716);
or U21854 (N_21854,N_19591,N_19601);
xor U21855 (N_21855,N_19733,N_20852);
nor U21856 (N_21856,N_19789,N_19572);
or U21857 (N_21857,N_19592,N_19935);
and U21858 (N_21858,N_19598,N_19764);
nor U21859 (N_21859,N_20618,N_20498);
xor U21860 (N_21860,N_19563,N_20897);
nor U21861 (N_21861,N_20428,N_19696);
xnor U21862 (N_21862,N_20077,N_20239);
and U21863 (N_21863,N_20600,N_20746);
or U21864 (N_21864,N_19752,N_20614);
nand U21865 (N_21865,N_19736,N_19915);
nand U21866 (N_21866,N_20730,N_20122);
xnor U21867 (N_21867,N_19634,N_19829);
xnor U21868 (N_21868,N_19921,N_20984);
and U21869 (N_21869,N_20853,N_20498);
nor U21870 (N_21870,N_20117,N_19767);
nand U21871 (N_21871,N_20830,N_19985);
nor U21872 (N_21872,N_19525,N_20895);
xor U21873 (N_21873,N_19815,N_20541);
or U21874 (N_21874,N_20319,N_20318);
or U21875 (N_21875,N_19591,N_20799);
xor U21876 (N_21876,N_19603,N_20584);
xor U21877 (N_21877,N_19512,N_20054);
nand U21878 (N_21878,N_20312,N_20705);
or U21879 (N_21879,N_19721,N_20850);
xnor U21880 (N_21880,N_20307,N_20261);
and U21881 (N_21881,N_20035,N_20965);
or U21882 (N_21882,N_20551,N_20741);
and U21883 (N_21883,N_20764,N_19790);
xnor U21884 (N_21884,N_20852,N_20302);
nor U21885 (N_21885,N_19749,N_19625);
nand U21886 (N_21886,N_20216,N_20105);
and U21887 (N_21887,N_19927,N_19866);
nor U21888 (N_21888,N_20886,N_20724);
and U21889 (N_21889,N_20000,N_20629);
nand U21890 (N_21890,N_20596,N_19946);
xor U21891 (N_21891,N_20793,N_20260);
xnor U21892 (N_21892,N_19980,N_19783);
nand U21893 (N_21893,N_19808,N_20496);
and U21894 (N_21894,N_20756,N_20282);
or U21895 (N_21895,N_20505,N_20230);
or U21896 (N_21896,N_19771,N_20049);
or U21897 (N_21897,N_20364,N_20445);
and U21898 (N_21898,N_19697,N_20691);
nand U21899 (N_21899,N_19532,N_20876);
xor U21900 (N_21900,N_19992,N_20562);
xor U21901 (N_21901,N_20643,N_20662);
nor U21902 (N_21902,N_20148,N_20334);
and U21903 (N_21903,N_20151,N_20506);
and U21904 (N_21904,N_19576,N_19807);
xnor U21905 (N_21905,N_20745,N_20872);
nor U21906 (N_21906,N_20002,N_20232);
or U21907 (N_21907,N_19681,N_20326);
xnor U21908 (N_21908,N_19892,N_20485);
xor U21909 (N_21909,N_20366,N_19754);
and U21910 (N_21910,N_19679,N_20421);
nand U21911 (N_21911,N_20212,N_20828);
or U21912 (N_21912,N_19771,N_20590);
nand U21913 (N_21913,N_20738,N_19872);
xnor U21914 (N_21914,N_20359,N_20713);
nand U21915 (N_21915,N_20796,N_19563);
xnor U21916 (N_21916,N_19755,N_20651);
and U21917 (N_21917,N_20734,N_20294);
xor U21918 (N_21918,N_19922,N_20574);
or U21919 (N_21919,N_20879,N_19888);
and U21920 (N_21920,N_20741,N_20213);
nor U21921 (N_21921,N_20745,N_20225);
or U21922 (N_21922,N_20138,N_20740);
or U21923 (N_21923,N_20007,N_20577);
or U21924 (N_21924,N_20404,N_20875);
or U21925 (N_21925,N_20347,N_20480);
nor U21926 (N_21926,N_20584,N_19559);
nand U21927 (N_21927,N_20791,N_20113);
xnor U21928 (N_21928,N_20067,N_20309);
or U21929 (N_21929,N_20096,N_19968);
nor U21930 (N_21930,N_20753,N_20823);
and U21931 (N_21931,N_20865,N_20626);
and U21932 (N_21932,N_19775,N_20326);
nor U21933 (N_21933,N_20966,N_19544);
nor U21934 (N_21934,N_20548,N_20180);
nor U21935 (N_21935,N_20087,N_20855);
and U21936 (N_21936,N_19787,N_20691);
xor U21937 (N_21937,N_20052,N_20805);
xnor U21938 (N_21938,N_20630,N_19525);
and U21939 (N_21939,N_19974,N_20282);
or U21940 (N_21940,N_20229,N_19691);
and U21941 (N_21941,N_19795,N_19869);
xor U21942 (N_21942,N_19690,N_20430);
and U21943 (N_21943,N_20796,N_20773);
nor U21944 (N_21944,N_20890,N_20979);
and U21945 (N_21945,N_19948,N_20942);
nor U21946 (N_21946,N_20475,N_19588);
or U21947 (N_21947,N_19655,N_19569);
or U21948 (N_21948,N_20366,N_20712);
nand U21949 (N_21949,N_20480,N_20941);
and U21950 (N_21950,N_20543,N_19720);
nor U21951 (N_21951,N_20336,N_19755);
nand U21952 (N_21952,N_20967,N_20681);
and U21953 (N_21953,N_20692,N_19952);
xor U21954 (N_21954,N_19665,N_20298);
nand U21955 (N_21955,N_19648,N_20123);
nor U21956 (N_21956,N_20578,N_20575);
and U21957 (N_21957,N_20662,N_20788);
and U21958 (N_21958,N_20264,N_20721);
nand U21959 (N_21959,N_19839,N_20676);
nor U21960 (N_21960,N_19988,N_20917);
nand U21961 (N_21961,N_19947,N_20888);
or U21962 (N_21962,N_19611,N_19719);
nand U21963 (N_21963,N_20374,N_20032);
and U21964 (N_21964,N_20334,N_20737);
nand U21965 (N_21965,N_20250,N_20692);
or U21966 (N_21966,N_19677,N_20646);
nand U21967 (N_21967,N_20830,N_20701);
and U21968 (N_21968,N_20645,N_19677);
nor U21969 (N_21969,N_20884,N_19508);
nand U21970 (N_21970,N_20473,N_20954);
nand U21971 (N_21971,N_19976,N_20402);
nor U21972 (N_21972,N_19578,N_20718);
xor U21973 (N_21973,N_20478,N_20927);
and U21974 (N_21974,N_20628,N_20417);
nand U21975 (N_21975,N_20027,N_20032);
nor U21976 (N_21976,N_19645,N_20443);
xor U21977 (N_21977,N_20198,N_20238);
and U21978 (N_21978,N_20924,N_19890);
nand U21979 (N_21979,N_19910,N_20426);
or U21980 (N_21980,N_19994,N_20849);
xor U21981 (N_21981,N_20247,N_20325);
or U21982 (N_21982,N_19804,N_20862);
xnor U21983 (N_21983,N_19659,N_19561);
nand U21984 (N_21984,N_20828,N_20410);
or U21985 (N_21985,N_20520,N_20217);
nor U21986 (N_21986,N_20572,N_20178);
or U21987 (N_21987,N_19779,N_19989);
nand U21988 (N_21988,N_20969,N_20399);
nor U21989 (N_21989,N_20539,N_19623);
and U21990 (N_21990,N_20306,N_19815);
xnor U21991 (N_21991,N_20690,N_20588);
and U21992 (N_21992,N_20981,N_19925);
nor U21993 (N_21993,N_20123,N_20103);
nand U21994 (N_21994,N_20693,N_20169);
or U21995 (N_21995,N_20939,N_20682);
nand U21996 (N_21996,N_19925,N_20107);
and U21997 (N_21997,N_20233,N_19547);
and U21998 (N_21998,N_19930,N_20507);
nor U21999 (N_21999,N_20207,N_20191);
xor U22000 (N_22000,N_20427,N_19689);
xnor U22001 (N_22001,N_19631,N_20127);
nand U22002 (N_22002,N_20108,N_19994);
nor U22003 (N_22003,N_20704,N_19971);
xor U22004 (N_22004,N_20533,N_19832);
nor U22005 (N_22005,N_19835,N_20538);
xor U22006 (N_22006,N_19732,N_20206);
or U22007 (N_22007,N_19532,N_20605);
xnor U22008 (N_22008,N_20784,N_20391);
and U22009 (N_22009,N_20800,N_20429);
nand U22010 (N_22010,N_19929,N_19737);
xnor U22011 (N_22011,N_19649,N_20633);
nand U22012 (N_22012,N_20885,N_20628);
xor U22013 (N_22013,N_20226,N_20420);
nand U22014 (N_22014,N_20553,N_20407);
nand U22015 (N_22015,N_20788,N_20335);
nand U22016 (N_22016,N_20534,N_19639);
nand U22017 (N_22017,N_19610,N_20623);
nor U22018 (N_22018,N_19791,N_19523);
and U22019 (N_22019,N_20395,N_20037);
and U22020 (N_22020,N_20644,N_20748);
and U22021 (N_22021,N_20426,N_20308);
and U22022 (N_22022,N_19741,N_19969);
nor U22023 (N_22023,N_20453,N_20302);
and U22024 (N_22024,N_20650,N_19800);
or U22025 (N_22025,N_20118,N_20283);
and U22026 (N_22026,N_20930,N_20069);
or U22027 (N_22027,N_20821,N_20982);
nor U22028 (N_22028,N_20137,N_19912);
or U22029 (N_22029,N_20677,N_20931);
nand U22030 (N_22030,N_19863,N_20349);
nand U22031 (N_22031,N_20232,N_19519);
xnor U22032 (N_22032,N_20270,N_20692);
and U22033 (N_22033,N_19669,N_19626);
or U22034 (N_22034,N_20071,N_20463);
nand U22035 (N_22035,N_20634,N_20641);
or U22036 (N_22036,N_20696,N_20187);
nor U22037 (N_22037,N_19550,N_20786);
xor U22038 (N_22038,N_20663,N_20033);
nor U22039 (N_22039,N_20680,N_20753);
and U22040 (N_22040,N_20124,N_20275);
nor U22041 (N_22041,N_19757,N_20945);
xor U22042 (N_22042,N_20202,N_19863);
or U22043 (N_22043,N_20797,N_19897);
xnor U22044 (N_22044,N_20214,N_20914);
and U22045 (N_22045,N_20939,N_20832);
and U22046 (N_22046,N_20094,N_20627);
xor U22047 (N_22047,N_19689,N_20154);
nor U22048 (N_22048,N_19642,N_19580);
nand U22049 (N_22049,N_20032,N_19973);
nor U22050 (N_22050,N_20757,N_20706);
xnor U22051 (N_22051,N_20588,N_19957);
xor U22052 (N_22052,N_20273,N_19882);
nor U22053 (N_22053,N_20030,N_20905);
nand U22054 (N_22054,N_20004,N_20746);
or U22055 (N_22055,N_19915,N_20973);
nand U22056 (N_22056,N_20517,N_20548);
xnor U22057 (N_22057,N_20512,N_20356);
or U22058 (N_22058,N_19505,N_20587);
and U22059 (N_22059,N_19622,N_20592);
xor U22060 (N_22060,N_20249,N_20232);
or U22061 (N_22061,N_19921,N_19598);
or U22062 (N_22062,N_19802,N_20855);
nand U22063 (N_22063,N_19801,N_20650);
nor U22064 (N_22064,N_19889,N_20523);
nand U22065 (N_22065,N_20609,N_20023);
nand U22066 (N_22066,N_20414,N_20816);
nand U22067 (N_22067,N_20088,N_19786);
and U22068 (N_22068,N_20775,N_19662);
nor U22069 (N_22069,N_19671,N_20499);
or U22070 (N_22070,N_20226,N_20862);
and U22071 (N_22071,N_20427,N_20774);
and U22072 (N_22072,N_19649,N_20135);
or U22073 (N_22073,N_20368,N_20153);
nand U22074 (N_22074,N_19547,N_20278);
nor U22075 (N_22075,N_19824,N_20653);
and U22076 (N_22076,N_19649,N_19854);
nor U22077 (N_22077,N_20737,N_20148);
nand U22078 (N_22078,N_20988,N_19725);
xnor U22079 (N_22079,N_20781,N_20400);
and U22080 (N_22080,N_19633,N_20753);
nand U22081 (N_22081,N_20604,N_20048);
nand U22082 (N_22082,N_19588,N_20547);
and U22083 (N_22083,N_20890,N_20359);
nor U22084 (N_22084,N_20408,N_20509);
and U22085 (N_22085,N_19753,N_19684);
nor U22086 (N_22086,N_20687,N_20928);
or U22087 (N_22087,N_19914,N_20809);
or U22088 (N_22088,N_20922,N_20101);
nand U22089 (N_22089,N_19892,N_20316);
xor U22090 (N_22090,N_20660,N_20125);
or U22091 (N_22091,N_20716,N_20706);
nand U22092 (N_22092,N_20864,N_20225);
nand U22093 (N_22093,N_19900,N_20557);
xor U22094 (N_22094,N_19510,N_19949);
or U22095 (N_22095,N_20007,N_19746);
nand U22096 (N_22096,N_20931,N_20705);
and U22097 (N_22097,N_20398,N_19666);
xor U22098 (N_22098,N_20398,N_20637);
or U22099 (N_22099,N_19786,N_20416);
xor U22100 (N_22100,N_19785,N_20210);
and U22101 (N_22101,N_20719,N_19744);
nor U22102 (N_22102,N_20642,N_20366);
xor U22103 (N_22103,N_20077,N_20055);
nor U22104 (N_22104,N_20345,N_19841);
xnor U22105 (N_22105,N_20797,N_20380);
xor U22106 (N_22106,N_19581,N_20968);
xor U22107 (N_22107,N_20661,N_20767);
and U22108 (N_22108,N_19547,N_19960);
nand U22109 (N_22109,N_19776,N_19822);
or U22110 (N_22110,N_20436,N_19883);
xnor U22111 (N_22111,N_20720,N_20817);
nand U22112 (N_22112,N_20476,N_19592);
and U22113 (N_22113,N_20047,N_20694);
nand U22114 (N_22114,N_20154,N_19691);
nand U22115 (N_22115,N_20892,N_20383);
nand U22116 (N_22116,N_19893,N_20845);
nor U22117 (N_22117,N_20390,N_20748);
nand U22118 (N_22118,N_19690,N_20013);
xor U22119 (N_22119,N_20088,N_20540);
and U22120 (N_22120,N_20508,N_20790);
nor U22121 (N_22121,N_20214,N_20001);
nand U22122 (N_22122,N_20412,N_19815);
nand U22123 (N_22123,N_20023,N_20615);
nand U22124 (N_22124,N_20966,N_19841);
nor U22125 (N_22125,N_20191,N_20482);
or U22126 (N_22126,N_19683,N_20119);
xor U22127 (N_22127,N_20623,N_20093);
and U22128 (N_22128,N_20917,N_19905);
or U22129 (N_22129,N_19597,N_20085);
xor U22130 (N_22130,N_19954,N_20189);
or U22131 (N_22131,N_20092,N_20013);
and U22132 (N_22132,N_19979,N_20770);
nor U22133 (N_22133,N_19606,N_20217);
nand U22134 (N_22134,N_20652,N_20869);
nor U22135 (N_22135,N_20481,N_20796);
nor U22136 (N_22136,N_19904,N_20241);
xnor U22137 (N_22137,N_20845,N_20398);
nor U22138 (N_22138,N_20223,N_20486);
and U22139 (N_22139,N_19668,N_20641);
xnor U22140 (N_22140,N_20204,N_20969);
nand U22141 (N_22141,N_20604,N_20927);
xnor U22142 (N_22142,N_20186,N_19542);
nand U22143 (N_22143,N_20136,N_20180);
and U22144 (N_22144,N_20409,N_20331);
xnor U22145 (N_22145,N_20822,N_19539);
and U22146 (N_22146,N_20183,N_19986);
and U22147 (N_22147,N_19713,N_19566);
and U22148 (N_22148,N_20580,N_19810);
xor U22149 (N_22149,N_20715,N_19961);
or U22150 (N_22150,N_20671,N_20504);
nor U22151 (N_22151,N_20043,N_20352);
and U22152 (N_22152,N_20146,N_20081);
and U22153 (N_22153,N_19893,N_20822);
nor U22154 (N_22154,N_20529,N_19713);
and U22155 (N_22155,N_19902,N_20811);
nor U22156 (N_22156,N_20857,N_20669);
xnor U22157 (N_22157,N_20837,N_20251);
and U22158 (N_22158,N_19774,N_20328);
nor U22159 (N_22159,N_20529,N_20918);
nor U22160 (N_22160,N_19990,N_20200);
and U22161 (N_22161,N_20089,N_20599);
and U22162 (N_22162,N_19595,N_20057);
nor U22163 (N_22163,N_20925,N_19709);
xor U22164 (N_22164,N_20256,N_20666);
xnor U22165 (N_22165,N_19531,N_20346);
and U22166 (N_22166,N_20755,N_20756);
xor U22167 (N_22167,N_20941,N_20385);
nand U22168 (N_22168,N_20492,N_19955);
nor U22169 (N_22169,N_20195,N_20733);
nor U22170 (N_22170,N_20108,N_20630);
and U22171 (N_22171,N_20927,N_19985);
nor U22172 (N_22172,N_20557,N_19529);
xor U22173 (N_22173,N_20925,N_19735);
xor U22174 (N_22174,N_20591,N_19872);
or U22175 (N_22175,N_19645,N_20224);
or U22176 (N_22176,N_19842,N_20682);
xnor U22177 (N_22177,N_20261,N_20104);
and U22178 (N_22178,N_20732,N_20705);
and U22179 (N_22179,N_20053,N_20407);
nand U22180 (N_22180,N_20321,N_20744);
nor U22181 (N_22181,N_20270,N_19870);
or U22182 (N_22182,N_20847,N_19991);
or U22183 (N_22183,N_20926,N_20857);
and U22184 (N_22184,N_20004,N_19637);
or U22185 (N_22185,N_20205,N_19986);
xnor U22186 (N_22186,N_20627,N_19511);
or U22187 (N_22187,N_20125,N_20614);
and U22188 (N_22188,N_20971,N_19735);
or U22189 (N_22189,N_20061,N_19886);
or U22190 (N_22190,N_20660,N_20518);
nand U22191 (N_22191,N_20269,N_20654);
nand U22192 (N_22192,N_20429,N_20361);
and U22193 (N_22193,N_20035,N_20426);
nand U22194 (N_22194,N_19756,N_19500);
or U22195 (N_22195,N_20151,N_19700);
nand U22196 (N_22196,N_19775,N_19525);
or U22197 (N_22197,N_20001,N_20777);
or U22198 (N_22198,N_20100,N_20832);
nand U22199 (N_22199,N_19703,N_20150);
or U22200 (N_22200,N_20600,N_20559);
nand U22201 (N_22201,N_19950,N_20413);
nor U22202 (N_22202,N_19618,N_20209);
or U22203 (N_22203,N_20282,N_19528);
xor U22204 (N_22204,N_20501,N_20711);
xor U22205 (N_22205,N_19906,N_20384);
or U22206 (N_22206,N_20226,N_20161);
and U22207 (N_22207,N_20100,N_20465);
or U22208 (N_22208,N_20275,N_20425);
xnor U22209 (N_22209,N_19728,N_19854);
or U22210 (N_22210,N_19577,N_20350);
or U22211 (N_22211,N_20563,N_20480);
or U22212 (N_22212,N_20097,N_19842);
nand U22213 (N_22213,N_20659,N_20782);
xor U22214 (N_22214,N_20657,N_19919);
nor U22215 (N_22215,N_20371,N_20571);
nand U22216 (N_22216,N_20094,N_19823);
xor U22217 (N_22217,N_19550,N_20034);
xnor U22218 (N_22218,N_20389,N_19716);
and U22219 (N_22219,N_19582,N_20737);
nand U22220 (N_22220,N_20764,N_19782);
and U22221 (N_22221,N_19648,N_20618);
xnor U22222 (N_22222,N_20094,N_20668);
xor U22223 (N_22223,N_20909,N_20129);
or U22224 (N_22224,N_20640,N_20337);
nand U22225 (N_22225,N_19882,N_20099);
and U22226 (N_22226,N_20104,N_20777);
or U22227 (N_22227,N_19983,N_20689);
and U22228 (N_22228,N_20578,N_20943);
and U22229 (N_22229,N_20411,N_20976);
nor U22230 (N_22230,N_19996,N_20940);
or U22231 (N_22231,N_20632,N_19970);
or U22232 (N_22232,N_19591,N_20588);
and U22233 (N_22233,N_20822,N_20389);
nand U22234 (N_22234,N_20035,N_20683);
or U22235 (N_22235,N_19752,N_19782);
nor U22236 (N_22236,N_20812,N_19709);
nor U22237 (N_22237,N_20205,N_20559);
and U22238 (N_22238,N_19595,N_20055);
xnor U22239 (N_22239,N_19743,N_19723);
xnor U22240 (N_22240,N_20311,N_20471);
nand U22241 (N_22241,N_19988,N_20283);
xnor U22242 (N_22242,N_20015,N_19825);
nand U22243 (N_22243,N_20745,N_20521);
nand U22244 (N_22244,N_20165,N_20577);
or U22245 (N_22245,N_19706,N_20875);
or U22246 (N_22246,N_19695,N_20954);
nand U22247 (N_22247,N_20607,N_19975);
nand U22248 (N_22248,N_19608,N_19757);
and U22249 (N_22249,N_19549,N_20232);
xnor U22250 (N_22250,N_20225,N_20073);
xor U22251 (N_22251,N_19862,N_20186);
nand U22252 (N_22252,N_19595,N_19502);
nand U22253 (N_22253,N_20812,N_20038);
nor U22254 (N_22254,N_20845,N_20587);
xnor U22255 (N_22255,N_20527,N_20604);
xor U22256 (N_22256,N_20937,N_20673);
nor U22257 (N_22257,N_19563,N_20475);
or U22258 (N_22258,N_19528,N_20354);
nor U22259 (N_22259,N_20483,N_20440);
nand U22260 (N_22260,N_20212,N_19934);
or U22261 (N_22261,N_20513,N_20897);
xor U22262 (N_22262,N_20565,N_19508);
xor U22263 (N_22263,N_20581,N_19966);
xor U22264 (N_22264,N_20285,N_20658);
and U22265 (N_22265,N_20016,N_19607);
xor U22266 (N_22266,N_20913,N_19543);
nor U22267 (N_22267,N_20939,N_20899);
or U22268 (N_22268,N_19876,N_20249);
nand U22269 (N_22269,N_20015,N_20005);
nand U22270 (N_22270,N_20192,N_20317);
xnor U22271 (N_22271,N_20988,N_20177);
and U22272 (N_22272,N_20872,N_20388);
nand U22273 (N_22273,N_20685,N_19815);
or U22274 (N_22274,N_19775,N_20152);
xnor U22275 (N_22275,N_20117,N_20343);
xor U22276 (N_22276,N_19939,N_19708);
or U22277 (N_22277,N_20463,N_20462);
or U22278 (N_22278,N_20780,N_19716);
or U22279 (N_22279,N_19967,N_20934);
nor U22280 (N_22280,N_19846,N_19906);
nor U22281 (N_22281,N_20457,N_20067);
nand U22282 (N_22282,N_20580,N_20162);
or U22283 (N_22283,N_20690,N_19713);
and U22284 (N_22284,N_19954,N_20858);
or U22285 (N_22285,N_20736,N_20397);
nor U22286 (N_22286,N_20960,N_20088);
xor U22287 (N_22287,N_20185,N_20230);
and U22288 (N_22288,N_20105,N_20872);
nor U22289 (N_22289,N_20521,N_19513);
xor U22290 (N_22290,N_20072,N_20928);
nand U22291 (N_22291,N_19675,N_20375);
nand U22292 (N_22292,N_19530,N_20877);
or U22293 (N_22293,N_19865,N_20616);
nand U22294 (N_22294,N_20489,N_20526);
and U22295 (N_22295,N_19660,N_20660);
xor U22296 (N_22296,N_19639,N_20696);
nand U22297 (N_22297,N_20938,N_20550);
xnor U22298 (N_22298,N_20831,N_20285);
nand U22299 (N_22299,N_20116,N_20861);
and U22300 (N_22300,N_19875,N_20981);
and U22301 (N_22301,N_20439,N_19556);
xnor U22302 (N_22302,N_19627,N_19838);
and U22303 (N_22303,N_20659,N_20780);
nor U22304 (N_22304,N_19828,N_20398);
nor U22305 (N_22305,N_20815,N_20295);
and U22306 (N_22306,N_19952,N_20123);
nor U22307 (N_22307,N_20131,N_20836);
nand U22308 (N_22308,N_19844,N_20086);
nor U22309 (N_22309,N_20042,N_20948);
and U22310 (N_22310,N_19682,N_19526);
or U22311 (N_22311,N_19829,N_20003);
nor U22312 (N_22312,N_20025,N_20023);
xor U22313 (N_22313,N_20577,N_20752);
or U22314 (N_22314,N_20683,N_20330);
or U22315 (N_22315,N_19616,N_20201);
nand U22316 (N_22316,N_19630,N_19850);
nor U22317 (N_22317,N_20562,N_20601);
and U22318 (N_22318,N_20166,N_20475);
xor U22319 (N_22319,N_20425,N_20515);
nor U22320 (N_22320,N_19995,N_20120);
nor U22321 (N_22321,N_20038,N_19695);
xnor U22322 (N_22322,N_20376,N_20126);
nand U22323 (N_22323,N_20910,N_20943);
xnor U22324 (N_22324,N_19943,N_20213);
and U22325 (N_22325,N_20651,N_20660);
nand U22326 (N_22326,N_20368,N_19694);
and U22327 (N_22327,N_20403,N_20851);
and U22328 (N_22328,N_20142,N_19880);
nor U22329 (N_22329,N_20358,N_20836);
or U22330 (N_22330,N_20831,N_20778);
xnor U22331 (N_22331,N_20406,N_20576);
and U22332 (N_22332,N_19726,N_19541);
or U22333 (N_22333,N_19956,N_19931);
xnor U22334 (N_22334,N_20117,N_19779);
or U22335 (N_22335,N_19595,N_20821);
nor U22336 (N_22336,N_19907,N_20119);
or U22337 (N_22337,N_19951,N_20927);
nand U22338 (N_22338,N_20733,N_20987);
xor U22339 (N_22339,N_19690,N_20325);
nand U22340 (N_22340,N_20189,N_19503);
and U22341 (N_22341,N_20802,N_20889);
and U22342 (N_22342,N_20632,N_20178);
nand U22343 (N_22343,N_20573,N_20331);
nand U22344 (N_22344,N_20447,N_20405);
and U22345 (N_22345,N_19530,N_19788);
nand U22346 (N_22346,N_20768,N_20371);
and U22347 (N_22347,N_19541,N_20135);
and U22348 (N_22348,N_20856,N_19625);
and U22349 (N_22349,N_20836,N_19543);
or U22350 (N_22350,N_19542,N_19504);
nor U22351 (N_22351,N_19930,N_20985);
or U22352 (N_22352,N_20152,N_20737);
xnor U22353 (N_22353,N_20354,N_19770);
nor U22354 (N_22354,N_19828,N_19712);
or U22355 (N_22355,N_19988,N_19518);
or U22356 (N_22356,N_20314,N_19501);
or U22357 (N_22357,N_19868,N_19808);
nor U22358 (N_22358,N_19875,N_19505);
and U22359 (N_22359,N_19891,N_19833);
nor U22360 (N_22360,N_20412,N_19810);
and U22361 (N_22361,N_20546,N_19924);
nand U22362 (N_22362,N_20980,N_20144);
nor U22363 (N_22363,N_20024,N_20128);
or U22364 (N_22364,N_20410,N_19711);
and U22365 (N_22365,N_20242,N_20732);
and U22366 (N_22366,N_20874,N_20648);
nor U22367 (N_22367,N_19513,N_20207);
nor U22368 (N_22368,N_20224,N_20991);
nand U22369 (N_22369,N_19597,N_20523);
nand U22370 (N_22370,N_19838,N_20996);
and U22371 (N_22371,N_20408,N_19853);
and U22372 (N_22372,N_19805,N_20329);
and U22373 (N_22373,N_20239,N_20589);
xor U22374 (N_22374,N_20483,N_20236);
xor U22375 (N_22375,N_19938,N_20892);
xor U22376 (N_22376,N_20358,N_19992);
xor U22377 (N_22377,N_20024,N_20686);
nand U22378 (N_22378,N_20879,N_20926);
nor U22379 (N_22379,N_20581,N_20084);
nand U22380 (N_22380,N_20199,N_19935);
nor U22381 (N_22381,N_20181,N_19613);
xnor U22382 (N_22382,N_20222,N_20908);
and U22383 (N_22383,N_20299,N_19845);
and U22384 (N_22384,N_20140,N_19714);
nor U22385 (N_22385,N_20549,N_19811);
and U22386 (N_22386,N_20728,N_20175);
and U22387 (N_22387,N_20969,N_20789);
nand U22388 (N_22388,N_19581,N_19821);
and U22389 (N_22389,N_20135,N_19692);
or U22390 (N_22390,N_20152,N_20587);
and U22391 (N_22391,N_20461,N_19659);
and U22392 (N_22392,N_19707,N_20751);
nand U22393 (N_22393,N_20198,N_20592);
nor U22394 (N_22394,N_19902,N_20892);
and U22395 (N_22395,N_19523,N_20189);
xnor U22396 (N_22396,N_20498,N_20682);
nor U22397 (N_22397,N_20738,N_20923);
nand U22398 (N_22398,N_20620,N_20075);
and U22399 (N_22399,N_19833,N_20300);
and U22400 (N_22400,N_19510,N_20088);
nand U22401 (N_22401,N_20966,N_19898);
nand U22402 (N_22402,N_19557,N_20908);
or U22403 (N_22403,N_19899,N_19632);
nor U22404 (N_22404,N_20132,N_20546);
or U22405 (N_22405,N_19543,N_20228);
xnor U22406 (N_22406,N_20155,N_20053);
and U22407 (N_22407,N_20363,N_20033);
and U22408 (N_22408,N_20685,N_20474);
nand U22409 (N_22409,N_20390,N_20361);
nand U22410 (N_22410,N_19630,N_20277);
or U22411 (N_22411,N_20828,N_20832);
nor U22412 (N_22412,N_19864,N_20366);
and U22413 (N_22413,N_19608,N_20170);
nor U22414 (N_22414,N_20119,N_20288);
nor U22415 (N_22415,N_20156,N_19549);
or U22416 (N_22416,N_20617,N_19900);
nand U22417 (N_22417,N_20510,N_19752);
xor U22418 (N_22418,N_20212,N_20409);
and U22419 (N_22419,N_20245,N_20688);
or U22420 (N_22420,N_20542,N_19864);
xnor U22421 (N_22421,N_20236,N_19948);
and U22422 (N_22422,N_19549,N_20813);
nand U22423 (N_22423,N_19801,N_19894);
xnor U22424 (N_22424,N_19640,N_20341);
and U22425 (N_22425,N_20818,N_20641);
nand U22426 (N_22426,N_19651,N_20636);
xor U22427 (N_22427,N_19766,N_19953);
xor U22428 (N_22428,N_20345,N_19804);
or U22429 (N_22429,N_19817,N_20707);
xor U22430 (N_22430,N_20588,N_20983);
or U22431 (N_22431,N_20057,N_20649);
nand U22432 (N_22432,N_20217,N_20781);
and U22433 (N_22433,N_19527,N_20995);
nand U22434 (N_22434,N_19571,N_19596);
and U22435 (N_22435,N_20966,N_20663);
xor U22436 (N_22436,N_20990,N_20001);
xnor U22437 (N_22437,N_20809,N_19622);
and U22438 (N_22438,N_19883,N_20270);
or U22439 (N_22439,N_19512,N_20832);
xor U22440 (N_22440,N_20206,N_19759);
and U22441 (N_22441,N_20247,N_20386);
or U22442 (N_22442,N_20385,N_20176);
nand U22443 (N_22443,N_20328,N_19605);
nand U22444 (N_22444,N_20739,N_20702);
nand U22445 (N_22445,N_20698,N_19879);
nand U22446 (N_22446,N_19594,N_19995);
nand U22447 (N_22447,N_20333,N_19863);
nor U22448 (N_22448,N_19586,N_20508);
and U22449 (N_22449,N_20178,N_20916);
xnor U22450 (N_22450,N_20787,N_20061);
nor U22451 (N_22451,N_20654,N_19723);
nand U22452 (N_22452,N_19503,N_19579);
nor U22453 (N_22453,N_20519,N_20486);
and U22454 (N_22454,N_20889,N_20810);
or U22455 (N_22455,N_20578,N_20753);
and U22456 (N_22456,N_20841,N_19958);
nor U22457 (N_22457,N_20633,N_19500);
nand U22458 (N_22458,N_19712,N_20824);
nor U22459 (N_22459,N_20748,N_20241);
nor U22460 (N_22460,N_20323,N_20165);
and U22461 (N_22461,N_20138,N_20531);
or U22462 (N_22462,N_20777,N_20014);
xnor U22463 (N_22463,N_20393,N_20628);
and U22464 (N_22464,N_20579,N_20174);
and U22465 (N_22465,N_20241,N_20853);
nand U22466 (N_22466,N_20640,N_20156);
nor U22467 (N_22467,N_20379,N_20829);
or U22468 (N_22468,N_19584,N_19968);
nand U22469 (N_22469,N_20719,N_19631);
nor U22470 (N_22470,N_20528,N_20905);
nand U22471 (N_22471,N_20973,N_19811);
xnor U22472 (N_22472,N_20802,N_20300);
or U22473 (N_22473,N_19791,N_20227);
or U22474 (N_22474,N_20409,N_20192);
or U22475 (N_22475,N_20499,N_20951);
xnor U22476 (N_22476,N_19952,N_20125);
xnor U22477 (N_22477,N_19762,N_20818);
and U22478 (N_22478,N_19921,N_20895);
xor U22479 (N_22479,N_19617,N_19737);
nand U22480 (N_22480,N_20388,N_20401);
xor U22481 (N_22481,N_20134,N_20378);
nor U22482 (N_22482,N_20447,N_20199);
and U22483 (N_22483,N_20047,N_20246);
xor U22484 (N_22484,N_20172,N_19887);
nor U22485 (N_22485,N_20335,N_20624);
and U22486 (N_22486,N_19937,N_20129);
nand U22487 (N_22487,N_19522,N_20054);
nor U22488 (N_22488,N_20495,N_19809);
nor U22489 (N_22489,N_20720,N_20084);
xor U22490 (N_22490,N_19890,N_20705);
nor U22491 (N_22491,N_20729,N_20825);
nor U22492 (N_22492,N_20852,N_20564);
or U22493 (N_22493,N_20918,N_20551);
and U22494 (N_22494,N_19685,N_20145);
nor U22495 (N_22495,N_20324,N_20182);
xor U22496 (N_22496,N_20187,N_20634);
and U22497 (N_22497,N_19760,N_19549);
nand U22498 (N_22498,N_20157,N_19724);
nor U22499 (N_22499,N_20599,N_20566);
nor U22500 (N_22500,N_21675,N_22448);
or U22501 (N_22501,N_21254,N_21657);
nand U22502 (N_22502,N_21865,N_22404);
xnor U22503 (N_22503,N_21289,N_21364);
xor U22504 (N_22504,N_22096,N_22063);
nor U22505 (N_22505,N_21767,N_21804);
or U22506 (N_22506,N_21144,N_22323);
or U22507 (N_22507,N_21568,N_21445);
nor U22508 (N_22508,N_21511,N_21719);
xor U22509 (N_22509,N_21407,N_22278);
and U22510 (N_22510,N_21149,N_21901);
nor U22511 (N_22511,N_21346,N_21942);
xnor U22512 (N_22512,N_21746,N_21319);
xor U22513 (N_22513,N_22035,N_21612);
nand U22514 (N_22514,N_21832,N_21374);
nand U22515 (N_22515,N_21361,N_22335);
nor U22516 (N_22516,N_21064,N_21480);
and U22517 (N_22517,N_22496,N_21936);
and U22518 (N_22518,N_21070,N_21978);
or U22519 (N_22519,N_21425,N_22131);
or U22520 (N_22520,N_21862,N_21922);
or U22521 (N_22521,N_22019,N_21234);
nor U22522 (N_22522,N_22055,N_21146);
xor U22523 (N_22523,N_22119,N_21123);
nand U22524 (N_22524,N_21822,N_21178);
xor U22525 (N_22525,N_22249,N_22324);
and U22526 (N_22526,N_22393,N_21111);
and U22527 (N_22527,N_22214,N_22481);
nand U22528 (N_22528,N_21646,N_21184);
or U22529 (N_22529,N_21388,N_22356);
and U22530 (N_22530,N_22498,N_22106);
and U22531 (N_22531,N_21148,N_21994);
or U22532 (N_22532,N_22417,N_21837);
nor U22533 (N_22533,N_22385,N_21641);
xnor U22534 (N_22534,N_22003,N_21637);
nor U22535 (N_22535,N_21773,N_21105);
nand U22536 (N_22536,N_21427,N_22144);
nand U22537 (N_22537,N_21573,N_21975);
and U22538 (N_22538,N_21513,N_21626);
nand U22539 (N_22539,N_21439,N_21341);
or U22540 (N_22540,N_21337,N_22142);
nor U22541 (N_22541,N_22007,N_21741);
xor U22542 (N_22542,N_22499,N_21658);
or U22543 (N_22543,N_21372,N_22107);
and U22544 (N_22544,N_21733,N_22363);
and U22545 (N_22545,N_21005,N_22384);
and U22546 (N_22546,N_22456,N_21463);
and U22547 (N_22547,N_21759,N_21898);
or U22548 (N_22548,N_21801,N_22057);
nand U22549 (N_22549,N_21928,N_21417);
or U22550 (N_22550,N_21321,N_21494);
xnor U22551 (N_22551,N_22155,N_21878);
nor U22552 (N_22552,N_22315,N_21690);
nand U22553 (N_22553,N_22258,N_22039);
or U22554 (N_22554,N_21840,N_21044);
or U22555 (N_22555,N_22082,N_22112);
or U22556 (N_22556,N_21309,N_21958);
nor U22557 (N_22557,N_22203,N_21891);
nand U22558 (N_22558,N_22424,N_21405);
nor U22559 (N_22559,N_21583,N_22072);
or U22560 (N_22560,N_21279,N_21079);
xnor U22561 (N_22561,N_21382,N_21082);
or U22562 (N_22562,N_21864,N_21955);
xnor U22563 (N_22563,N_21487,N_21585);
xnor U22564 (N_22564,N_22068,N_22414);
and U22565 (N_22565,N_21877,N_21858);
and U22566 (N_22566,N_22455,N_22083);
or U22567 (N_22567,N_22040,N_21889);
xor U22568 (N_22568,N_21159,N_21045);
and U22569 (N_22569,N_22212,N_22188);
nor U22570 (N_22570,N_22291,N_22339);
nand U22571 (N_22571,N_21017,N_21711);
nor U22572 (N_22572,N_22489,N_21320);
or U22573 (N_22573,N_22129,N_22353);
nand U22574 (N_22574,N_21245,N_21007);
nor U22575 (N_22575,N_21314,N_21133);
nand U22576 (N_22576,N_21720,N_22141);
xor U22577 (N_22577,N_21293,N_22332);
and U22578 (N_22578,N_21169,N_21524);
and U22579 (N_22579,N_22017,N_21533);
or U22580 (N_22580,N_21555,N_21705);
or U22581 (N_22581,N_22317,N_21459);
and U22582 (N_22582,N_21117,N_22425);
nor U22583 (N_22583,N_22288,N_22478);
and U22584 (N_22584,N_22397,N_22190);
or U22585 (N_22585,N_22174,N_21038);
or U22586 (N_22586,N_22237,N_22463);
xor U22587 (N_22587,N_21292,N_21308);
nand U22588 (N_22588,N_21744,N_21881);
xor U22589 (N_22589,N_21244,N_22430);
xor U22590 (N_22590,N_21915,N_21677);
nand U22591 (N_22591,N_22494,N_21643);
nor U22592 (N_22592,N_22334,N_21298);
and U22593 (N_22593,N_21754,N_21941);
nor U22594 (N_22594,N_21887,N_21324);
xor U22595 (N_22595,N_21482,N_22394);
xnor U22596 (N_22596,N_21062,N_22216);
nand U22597 (N_22597,N_21917,N_22084);
xor U22598 (N_22598,N_22090,N_21563);
nor U22599 (N_22599,N_21313,N_21286);
xor U22600 (N_22600,N_22473,N_21999);
nand U22601 (N_22601,N_22330,N_21990);
and U22602 (N_22602,N_21181,N_22049);
and U22603 (N_22603,N_21725,N_21634);
nor U22604 (N_22604,N_21772,N_22041);
nor U22605 (N_22605,N_21399,N_21375);
nor U22606 (N_22606,N_22194,N_21135);
nor U22607 (N_22607,N_21454,N_22046);
and U22608 (N_22608,N_21285,N_22102);
nor U22609 (N_22609,N_21820,N_21479);
nand U22610 (N_22610,N_22105,N_21859);
or U22611 (N_22611,N_21106,N_21774);
or U22612 (N_22612,N_22423,N_21179);
and U22613 (N_22613,N_21885,N_22495);
xnor U22614 (N_22614,N_21544,N_22386);
xor U22615 (N_22615,N_21157,N_21297);
and U22616 (N_22616,N_21259,N_21014);
and U22617 (N_22617,N_22381,N_22474);
nand U22618 (N_22618,N_21226,N_21850);
xnor U22619 (N_22619,N_21795,N_21000);
nand U22620 (N_22620,N_21578,N_22239);
xor U22621 (N_22621,N_21347,N_22395);
and U22622 (N_22622,N_21470,N_22116);
nand U22623 (N_22623,N_21448,N_21561);
nand U22624 (N_22624,N_21827,N_21828);
and U22625 (N_22625,N_21271,N_21001);
nand U22626 (N_22626,N_21704,N_21531);
nand U22627 (N_22627,N_22004,N_21060);
or U22628 (N_22628,N_22198,N_21132);
xor U22629 (N_22629,N_21491,N_21108);
xnor U22630 (N_22630,N_21393,N_22338);
and U22631 (N_22631,N_22031,N_21874);
nand U22632 (N_22632,N_21876,N_22191);
and U22633 (N_22633,N_22293,N_21042);
or U22634 (N_22634,N_22059,N_22379);
and U22635 (N_22635,N_21776,N_21081);
or U22636 (N_22636,N_21593,N_22022);
nor U22637 (N_22637,N_22048,N_21846);
and U22638 (N_22638,N_22349,N_22285);
nand U22639 (N_22639,N_21302,N_21848);
nand U22640 (N_22640,N_21391,N_22151);
nand U22641 (N_22641,N_21868,N_21446);
and U22642 (N_22642,N_22294,N_21048);
xor U22643 (N_22643,N_21167,N_21002);
nand U22644 (N_22644,N_21597,N_21201);
nor U22645 (N_22645,N_22015,N_21196);
nor U22646 (N_22646,N_21666,N_22436);
and U22647 (N_22647,N_22421,N_21779);
or U22648 (N_22648,N_22118,N_21897);
nand U22649 (N_22649,N_22081,N_21582);
xor U22650 (N_22650,N_22325,N_22342);
and U22651 (N_22651,N_21629,N_21562);
or U22652 (N_22652,N_22201,N_21202);
nand U22653 (N_22653,N_21961,N_21543);
or U22654 (N_22654,N_21041,N_22305);
nand U22655 (N_22655,N_21429,N_21194);
and U22656 (N_22656,N_21537,N_22269);
nor U22657 (N_22657,N_22099,N_22235);
nor U22658 (N_22658,N_21342,N_21376);
and U22659 (N_22659,N_21488,N_22160);
xnor U22660 (N_22660,N_21006,N_22482);
nor U22661 (N_22661,N_21318,N_21571);
xor U22662 (N_22662,N_21465,N_22462);
or U22663 (N_22663,N_21198,N_21696);
nor U22664 (N_22664,N_21930,N_21932);
nand U22665 (N_22665,N_21241,N_21951);
and U22666 (N_22666,N_21505,N_21577);
or U22667 (N_22667,N_21046,N_22075);
nand U22668 (N_22668,N_21782,N_21174);
or U22669 (N_22669,N_21039,N_22266);
or U22670 (N_22670,N_22488,N_22132);
or U22671 (N_22671,N_22245,N_21836);
xor U22672 (N_22672,N_21397,N_21683);
nand U22673 (N_22673,N_22290,N_21592);
xor U22674 (N_22674,N_22023,N_21518);
or U22675 (N_22675,N_22202,N_21581);
and U22676 (N_22676,N_21963,N_22357);
and U22677 (N_22677,N_21183,N_21402);
nor U22678 (N_22678,N_22110,N_22274);
or U22679 (N_22679,N_22217,N_21525);
and U22680 (N_22680,N_21466,N_21158);
nand U22681 (N_22681,N_21145,N_21410);
nand U22682 (N_22682,N_21065,N_21778);
nor U22683 (N_22683,N_22070,N_21988);
xor U22684 (N_22684,N_21240,N_21053);
nor U22685 (N_22685,N_21280,N_21238);
nor U22686 (N_22686,N_21693,N_21945);
and U22687 (N_22687,N_21902,N_21816);
and U22688 (N_22688,N_22368,N_21606);
xor U22689 (N_22689,N_21449,N_22219);
and U22690 (N_22690,N_22163,N_21012);
or U22691 (N_22691,N_21270,N_21644);
xor U22692 (N_22692,N_21956,N_21576);
nand U22693 (N_22693,N_21926,N_22360);
and U22694 (N_22694,N_21225,N_21362);
nand U22695 (N_22695,N_21684,N_22279);
or U22696 (N_22696,N_21219,N_22336);
nand U22697 (N_22697,N_21824,N_21009);
nor U22698 (N_22698,N_22387,N_21232);
and U22699 (N_22699,N_22128,N_21110);
or U22700 (N_22700,N_22168,N_21973);
and U22701 (N_22701,N_21390,N_21189);
and U22702 (N_22702,N_21147,N_21565);
xor U22703 (N_22703,N_21129,N_21352);
xor U22704 (N_22704,N_21919,N_22087);
xnor U22705 (N_22705,N_22408,N_21025);
nand U22706 (N_22706,N_21825,N_21283);
and U22707 (N_22707,N_22350,N_21688);
xnor U22708 (N_22708,N_21246,N_22447);
nand U22709 (N_22709,N_21331,N_22162);
nor U22710 (N_22710,N_22058,N_22497);
nor U22711 (N_22711,N_21717,N_21303);
and U22712 (N_22712,N_21163,N_21277);
nor U22713 (N_22713,N_21142,N_21030);
nor U22714 (N_22714,N_22309,N_21076);
xor U22715 (N_22715,N_21713,N_22113);
nor U22716 (N_22716,N_22479,N_21895);
or U22717 (N_22717,N_21831,N_22125);
and U22718 (N_22718,N_21998,N_22001);
nand U22719 (N_22719,N_21799,N_21514);
and U22720 (N_22720,N_22009,N_21687);
and U22721 (N_22721,N_21500,N_21594);
nand U22722 (N_22722,N_21854,N_22080);
and U22723 (N_22723,N_21156,N_21103);
nor U22724 (N_22724,N_21755,N_22164);
nor U22725 (N_22725,N_21495,N_22008);
or U22726 (N_22726,N_21981,N_22139);
xnor U22727 (N_22727,N_21781,N_21984);
nand U22728 (N_22728,N_22165,N_22422);
and U22729 (N_22729,N_21236,N_21003);
or U22730 (N_22730,N_21154,N_22171);
and U22731 (N_22731,N_21193,N_22077);
and U22732 (N_22732,N_21243,N_21507);
nor U22733 (N_22733,N_22183,N_21155);
nor U22734 (N_22734,N_21310,N_22262);
and U22735 (N_22735,N_22167,N_22147);
and U22736 (N_22736,N_21510,N_21451);
and U22737 (N_22737,N_21851,N_21114);
nand U22738 (N_22738,N_21921,N_22468);
nor U22739 (N_22739,N_21925,N_21467);
or U22740 (N_22740,N_21369,N_22480);
nor U22741 (N_22741,N_21589,N_22161);
or U22742 (N_22742,N_21879,N_22490);
nand U22743 (N_22743,N_21264,N_22265);
and U22744 (N_22744,N_22218,N_21587);
nor U22745 (N_22745,N_21473,N_21966);
xor U22746 (N_22746,N_21989,N_21492);
and U22747 (N_22747,N_21140,N_21871);
nand U22748 (N_22748,N_21517,N_22121);
or U22749 (N_22749,N_21430,N_21223);
nor U22750 (N_22750,N_21419,N_21940);
and U22751 (N_22751,N_21345,N_21086);
or U22752 (N_22752,N_21261,N_21913);
nand U22753 (N_22753,N_22034,N_21783);
xor U22754 (N_22754,N_21747,N_21924);
or U22755 (N_22755,N_21287,N_21251);
and U22756 (N_22756,N_22377,N_21315);
xnor U22757 (N_22757,N_22244,N_21983);
nand U22758 (N_22758,N_21627,N_21911);
xnor U22759 (N_22759,N_21475,N_22260);
nor U22760 (N_22760,N_21164,N_21021);
nor U22761 (N_22761,N_21821,N_22086);
nand U22762 (N_22762,N_21845,N_21674);
nor U22763 (N_22763,N_21443,N_21457);
nand U22764 (N_22764,N_21377,N_21977);
nor U22765 (N_22765,N_22460,N_22108);
nor U22766 (N_22766,N_21227,N_21976);
nor U22767 (N_22767,N_21288,N_21916);
and U22768 (N_22768,N_21266,N_21695);
and U22769 (N_22769,N_21468,N_21528);
nand U22770 (N_22770,N_22427,N_22069);
nand U22771 (N_22771,N_21914,N_22405);
xor U22772 (N_22772,N_21306,N_21762);
nand U22773 (N_22773,N_21008,N_22348);
nor U22774 (N_22774,N_22442,N_21541);
and U22775 (N_22775,N_21073,N_21823);
xor U22776 (N_22776,N_21934,N_22143);
nand U22777 (N_22777,N_21617,N_22486);
and U22778 (N_22778,N_22018,N_21997);
or U22779 (N_22779,N_21431,N_21250);
or U22780 (N_22780,N_21075,N_22210);
nand U22781 (N_22781,N_21182,N_22440);
nor U22782 (N_22782,N_22391,N_21549);
or U22783 (N_22783,N_22060,N_22370);
nor U22784 (N_22784,N_21952,N_21722);
nor U22785 (N_22785,N_21483,N_22374);
xor U22786 (N_22786,N_21204,N_22383);
or U22787 (N_22787,N_22373,N_21662);
xnor U22788 (N_22788,N_22185,N_22465);
nand U22789 (N_22789,N_22432,N_22011);
or U22790 (N_22790,N_22002,N_21753);
or U22791 (N_22791,N_21899,N_22200);
nand U22792 (N_22792,N_21253,N_21367);
nor U22793 (N_22793,N_21161,N_22382);
nand U22794 (N_22794,N_22104,N_21900);
or U22795 (N_22795,N_21353,N_22122);
nand U22796 (N_22796,N_21462,N_21501);
and U22797 (N_22797,N_22375,N_21233);
nor U22798 (N_22798,N_21789,N_22493);
or U22799 (N_22799,N_21024,N_21819);
nand U22800 (N_22800,N_21098,N_21569);
nand U22801 (N_22801,N_22458,N_21249);
nor U22802 (N_22802,N_22042,N_21853);
or U22803 (N_22803,N_21530,N_21972);
nor U22804 (N_22804,N_21217,N_21216);
xnor U22805 (N_22805,N_22230,N_21170);
xnor U22806 (N_22806,N_22340,N_21604);
xnor U22807 (N_22807,N_21995,N_21428);
nand U22808 (N_22808,N_21113,N_22439);
and U22809 (N_22809,N_21115,N_21094);
xnor U22810 (N_22810,N_21923,N_22180);
nand U22811 (N_22811,N_21214,N_21168);
xor U22812 (N_22812,N_21265,N_22123);
or U22813 (N_22813,N_22354,N_21716);
or U22814 (N_22814,N_22076,N_22101);
and U22815 (N_22815,N_21213,N_21931);
or U22816 (N_22816,N_21171,N_21413);
nand U22817 (N_22817,N_22492,N_21317);
nor U22818 (N_22818,N_22403,N_21378);
and U22819 (N_22819,N_22233,N_21867);
xnor U22820 (N_22820,N_21992,N_22038);
nand U22821 (N_22821,N_21496,N_21740);
and U22822 (N_22822,N_21508,N_22364);
nor U22823 (N_22823,N_21034,N_21190);
nor U22824 (N_22824,N_22091,N_22308);
or U22825 (N_22825,N_22261,N_21392);
nand U22826 (N_22826,N_21020,N_22206);
nor U22827 (N_22827,N_21752,N_21013);
nand U22828 (N_22828,N_22114,N_21077);
nor U22829 (N_22829,N_21209,N_21400);
and U22830 (N_22830,N_21126,N_21329);
and U22831 (N_22831,N_21539,N_21043);
and U22832 (N_22832,N_22322,N_22032);
or U22833 (N_22833,N_22173,N_21939);
nand U22834 (N_22834,N_22156,N_22170);
nor U22835 (N_22835,N_21295,N_22193);
xor U22836 (N_22836,N_22396,N_21101);
nand U22837 (N_22837,N_21150,N_22028);
and U22838 (N_22838,N_22369,N_22213);
or U22839 (N_22839,N_21905,N_21485);
nand U22840 (N_22840,N_22254,N_21080);
xor U22841 (N_22841,N_21927,N_21621);
nor U22842 (N_22842,N_21120,N_22454);
xnor U22843 (N_22843,N_21212,N_22412);
xnor U22844 (N_22844,N_21422,N_21545);
and U22845 (N_22845,N_21838,N_21671);
or U22846 (N_22846,N_21609,N_21456);
and U22847 (N_22847,N_21833,N_21971);
nand U22848 (N_22848,N_21016,N_22136);
or U22849 (N_22849,N_21200,N_22115);
xor U22850 (N_22850,N_22301,N_22263);
and U22851 (N_22851,N_22150,N_22074);
nor U22852 (N_22852,N_21097,N_21745);
nand U22853 (N_22853,N_22148,N_21893);
nand U22854 (N_22854,N_21022,N_21398);
nor U22855 (N_22855,N_22410,N_21489);
nor U22856 (N_22856,N_22199,N_21461);
nand U22857 (N_22857,N_21197,N_21055);
or U22858 (N_22858,N_21360,N_21102);
nor U22859 (N_22859,N_21680,N_21050);
nor U22860 (N_22860,N_22461,N_21807);
nand U22861 (N_22861,N_22146,N_21188);
nand U22862 (N_22862,N_22178,N_22420);
nand U22863 (N_22863,N_21438,N_22208);
or U22864 (N_22864,N_21385,N_21712);
and U22865 (N_22865,N_22043,N_21738);
or U22866 (N_22866,N_21694,N_21262);
xnor U22867 (N_22867,N_21109,N_21718);
xor U22868 (N_22868,N_21714,N_22021);
or U22869 (N_22869,N_21811,N_21386);
xnor U22870 (N_22870,N_21325,N_21567);
or U22871 (N_22871,N_21300,N_21506);
nand U22872 (N_22872,N_22225,N_22389);
xor U22873 (N_22873,N_21996,N_22345);
nand U22874 (N_22874,N_21529,N_21379);
or U22875 (N_22875,N_21775,N_21061);
and U22876 (N_22876,N_21723,N_21328);
or U22877 (N_22877,N_21185,N_21019);
and U22878 (N_22878,N_22388,N_21269);
and U22879 (N_22879,N_21970,N_21797);
nor U22880 (N_22880,N_22270,N_22220);
and U22881 (N_22881,N_22371,N_22402);
and U22882 (N_22882,N_21894,N_21826);
or U22883 (N_22883,N_21964,N_22277);
or U22884 (N_22884,N_22145,N_22172);
or U22885 (N_22885,N_22097,N_21596);
and U22886 (N_22886,N_22413,N_21127);
nand U22887 (N_22887,N_21909,N_21869);
or U22888 (N_22888,N_22333,N_21406);
xnor U22889 (N_22889,N_22416,N_22268);
xnor U22890 (N_22890,N_22453,N_21960);
xor U22891 (N_22891,N_21408,N_21435);
nand U22892 (N_22892,N_22272,N_21031);
nor U22893 (N_22893,N_21160,N_22056);
nor U22894 (N_22894,N_22310,N_21206);
nand U22895 (N_22895,N_21558,N_21165);
and U22896 (N_22896,N_21880,N_21910);
nand U22897 (N_22897,N_22292,N_21373);
nand U22898 (N_22898,N_21237,N_21935);
nor U22899 (N_22899,N_21538,N_22399);
nor U22900 (N_22900,N_22435,N_22341);
nand U22901 (N_22901,N_21835,N_21761);
nor U22902 (N_22902,N_22337,N_21619);
and U22903 (N_22903,N_21614,N_22100);
xnor U22904 (N_22904,N_22477,N_22376);
and U22905 (N_22905,N_22429,N_22103);
or U22906 (N_22906,N_21843,N_21628);
xor U22907 (N_22907,N_21540,N_21137);
nand U22908 (N_22908,N_21040,N_22281);
xor U22909 (N_22909,N_21802,N_21095);
xor U22910 (N_22910,N_21534,N_22437);
nor U22911 (N_22911,N_22321,N_21499);
nor U22912 (N_22912,N_21312,N_21566);
xnor U22913 (N_22913,N_21847,N_21409);
or U22914 (N_22914,N_21526,N_22130);
nand U22915 (N_22915,N_22367,N_21715);
xnor U22916 (N_22916,N_22027,N_22013);
nor U22917 (N_22917,N_21504,N_21639);
nand U22918 (N_22918,N_21866,N_21728);
nand U22919 (N_22919,N_21980,N_21344);
or U22920 (N_22920,N_22483,N_21830);
and U22921 (N_22921,N_21890,N_21333);
nor U22922 (N_22922,N_21010,N_21519);
or U22923 (N_22923,N_22024,N_21950);
xnor U22924 (N_22924,N_21100,N_21231);
xnor U22925 (N_22925,N_22359,N_21959);
xnor U22926 (N_22926,N_22187,N_22111);
and U22927 (N_22927,N_21575,N_22238);
and U22928 (N_22928,N_21686,N_21230);
xor U22929 (N_22929,N_21748,N_21138);
and U22930 (N_22930,N_21294,N_21702);
xnor U22931 (N_22931,N_21588,N_21542);
and U22932 (N_22932,N_21882,N_21709);
nand U22933 (N_22933,N_21260,N_21818);
nand U22934 (N_22934,N_21692,N_21757);
xnor U22935 (N_22935,N_22316,N_21645);
and U22936 (N_22936,N_22295,N_21291);
or U22937 (N_22937,N_22476,N_22303);
nand U22938 (N_22938,N_21724,N_21829);
xor U22939 (N_22939,N_21857,N_22062);
and U22940 (N_22940,N_21296,N_22431);
or U22941 (N_22941,N_22406,N_21469);
nor U22942 (N_22942,N_21727,N_21560);
and U22943 (N_22943,N_21777,N_21788);
nand U22944 (N_22944,N_21841,N_21340);
or U22945 (N_22945,N_22409,N_21057);
nand U22946 (N_22946,N_21436,N_21125);
nand U22947 (N_22947,N_21943,N_21796);
xnor U22948 (N_22948,N_22469,N_21598);
nor U22949 (N_22949,N_22275,N_21268);
or U22950 (N_22950,N_21450,N_21503);
xor U22951 (N_22951,N_21613,N_21872);
nor U22952 (N_22952,N_22253,N_21672);
and U22953 (N_22953,N_22451,N_21652);
or U22954 (N_22954,N_22236,N_21701);
and U22955 (N_22955,N_21281,N_22014);
and U22956 (N_22956,N_21359,N_21187);
or U22957 (N_22957,N_21258,N_21486);
or U22958 (N_22958,N_22443,N_21363);
nor U22959 (N_22959,N_21944,N_21474);
and U22960 (N_22960,N_21356,N_21242);
and U22961 (N_22961,N_22065,N_21497);
nor U22962 (N_22962,N_21424,N_21625);
nor U22963 (N_22963,N_21305,N_22006);
or U22964 (N_22964,N_21371,N_22390);
xor U22965 (N_22965,N_21069,N_21912);
or U22966 (N_22966,N_21074,N_22152);
or U22967 (N_22967,N_21636,N_21834);
nand U22968 (N_22968,N_22358,N_21176);
xnor U22969 (N_22969,N_21166,N_22153);
nor U22970 (N_22970,N_21222,N_22312);
xnor U22971 (N_22971,N_21965,N_21273);
nor U22972 (N_22972,N_21967,N_21557);
or U22973 (N_22973,N_21121,N_21350);
nand U22974 (N_22974,N_21685,N_22037);
xnor U22975 (N_22975,N_21962,N_21739);
xor U22976 (N_22976,N_22380,N_21066);
nor U22977 (N_22977,N_21354,N_21812);
nor U22978 (N_22978,N_21803,N_21177);
nand U22979 (N_22979,N_21205,N_21173);
or U22980 (N_22980,N_21153,N_21937);
nand U22981 (N_22981,N_21805,N_22098);
and U22982 (N_22982,N_21118,N_21681);
xnor U22983 (N_22983,N_21343,N_22355);
and U22984 (N_22984,N_22299,N_21256);
or U22985 (N_22985,N_22211,N_22030);
nand U22986 (N_22986,N_21335,N_22186);
nand U22987 (N_22987,N_21886,N_21721);
nand U22988 (N_22988,N_22050,N_22071);
or U22989 (N_22989,N_22149,N_21063);
and U22990 (N_22990,N_21765,N_21472);
or U22991 (N_22991,N_22445,N_22307);
nand U22992 (N_22992,N_21067,N_21656);
or U22993 (N_22993,N_21968,N_22250);
and U22994 (N_22994,N_21027,N_21660);
nand U22995 (N_22995,N_21396,N_22415);
nor U22996 (N_22996,N_22246,N_22135);
nor U22997 (N_22997,N_21648,N_22433);
nor U22998 (N_22998,N_22446,N_21798);
or U22999 (N_22999,N_21018,N_22184);
nand U23000 (N_23000,N_21059,N_22079);
nor U23001 (N_23001,N_21790,N_21987);
nor U23002 (N_23002,N_22182,N_22209);
and U23003 (N_23003,N_21404,N_22227);
and U23004 (N_23004,N_21623,N_21092);
and U23005 (N_23005,N_22352,N_22255);
nand U23006 (N_23006,N_21768,N_21141);
or U23007 (N_23007,N_21366,N_21235);
and U23008 (N_23008,N_22089,N_21276);
xor U23009 (N_23009,N_22280,N_22426);
and U23010 (N_23010,N_21743,N_22464);
and U23011 (N_23011,N_21601,N_22085);
nand U23012 (N_23012,N_21647,N_22326);
nor U23013 (N_23013,N_21855,N_21883);
nand U23014 (N_23014,N_22195,N_21957);
xnor U23015 (N_23015,N_21638,N_22248);
or U23016 (N_23016,N_21348,N_22066);
and U23017 (N_23017,N_21085,N_21116);
and U23018 (N_23018,N_21764,N_22078);
nor U23019 (N_23019,N_21370,N_21599);
or U23020 (N_23020,N_21550,N_21839);
or U23021 (N_23021,N_21632,N_21661);
or U23022 (N_23022,N_22319,N_21083);
and U23023 (N_23023,N_22438,N_21982);
and U23024 (N_23024,N_21275,N_21175);
nor U23025 (N_23025,N_22092,N_22061);
nor U23026 (N_23026,N_21052,N_21809);
and U23027 (N_23027,N_21432,N_22378);
nand U23028 (N_23028,N_21920,N_21192);
or U23029 (N_23029,N_21139,N_21215);
and U23030 (N_23030,N_21654,N_22306);
and U23031 (N_23031,N_21104,N_22457);
xor U23032 (N_23032,N_21051,N_21595);
xnor U23033 (N_23033,N_21278,N_22444);
and U23034 (N_23034,N_21252,N_21616);
or U23035 (N_23035,N_22000,N_22257);
nor U23036 (N_23036,N_21056,N_22215);
nand U23037 (N_23037,N_21985,N_21698);
xor U23038 (N_23038,N_22273,N_21420);
or U23039 (N_23039,N_21036,N_21172);
nor U23040 (N_23040,N_21653,N_21954);
and U23041 (N_23041,N_21351,N_21136);
nand U23042 (N_23042,N_21515,N_21131);
nand U23043 (N_23043,N_22407,N_21130);
xor U23044 (N_23044,N_21433,N_22287);
and U23045 (N_23045,N_22095,N_21316);
xnor U23046 (N_23046,N_21929,N_22401);
nor U23047 (N_23047,N_22328,N_21330);
or U23048 (N_23048,N_22045,N_21602);
or U23049 (N_23049,N_22452,N_21143);
xnor U23050 (N_23050,N_22343,N_21304);
or U23051 (N_23051,N_21401,N_21327);
nand U23052 (N_23052,N_21049,N_21640);
nor U23053 (N_23053,N_22298,N_21707);
or U23054 (N_23054,N_21054,N_21668);
nor U23055 (N_23055,N_21785,N_22346);
xor U23056 (N_23056,N_21071,N_21806);
nand U23057 (N_23057,N_22313,N_21600);
or U23058 (N_23058,N_21394,N_21650);
xor U23059 (N_23059,N_22176,N_21607);
nand U23060 (N_23060,N_22450,N_21706);
xor U23061 (N_23061,N_22205,N_21800);
nor U23062 (N_23062,N_21415,N_22252);
and U23063 (N_23063,N_22224,N_21028);
or U23064 (N_23064,N_21863,N_21603);
xnor U23065 (N_23065,N_22033,N_22140);
and U23066 (N_23066,N_21947,N_21559);
nor U23067 (N_23067,N_21742,N_21888);
and U23068 (N_23068,N_21124,N_21763);
or U23069 (N_23069,N_21708,N_21817);
nand U23070 (N_23070,N_22197,N_21453);
nor U23071 (N_23071,N_21093,N_22177);
nand U23072 (N_23072,N_21769,N_21162);
and U23073 (N_23073,N_22311,N_21907);
xor U23074 (N_23074,N_22470,N_21186);
or U23075 (N_23075,N_22053,N_21991);
and U23076 (N_23076,N_21336,N_21758);
xor U23077 (N_23077,N_21090,N_22247);
or U23078 (N_23078,N_21437,N_21383);
and U23079 (N_23079,N_21199,N_21861);
xnor U23080 (N_23080,N_21750,N_21323);
nand U23081 (N_23081,N_22296,N_21949);
nor U23082 (N_23082,N_21896,N_22181);
nor U23083 (N_23083,N_22459,N_21068);
or U23084 (N_23084,N_22361,N_21673);
xor U23085 (N_23085,N_21792,N_22472);
and U23086 (N_23086,N_21455,N_22192);
and U23087 (N_23087,N_21730,N_21418);
nand U23088 (N_23088,N_21221,N_22372);
and U23089 (N_23089,N_21703,N_22138);
xor U23090 (N_23090,N_21191,N_21756);
nor U23091 (N_23091,N_21334,N_22175);
and U23092 (N_23092,N_21842,N_21731);
xnor U23093 (N_23093,N_21274,N_22094);
nand U23094 (N_23094,N_21938,N_21536);
and U23095 (N_23095,N_21903,N_22466);
and U23096 (N_23096,N_21047,N_21493);
or U23097 (N_23097,N_21736,N_21272);
nand U23098 (N_23098,N_21969,N_22159);
nor U23099 (N_23099,N_21023,N_21091);
and U23100 (N_23100,N_22327,N_22051);
or U23101 (N_23101,N_22264,N_22134);
xnor U23102 (N_23102,N_21387,N_21444);
and U23103 (N_23103,N_21332,N_22228);
xor U23104 (N_23104,N_21365,N_21478);
nor U23105 (N_23105,N_21326,N_22221);
xor U23106 (N_23106,N_21771,N_21037);
nor U23107 (N_23107,N_22016,N_22133);
nor U23108 (N_23108,N_21622,N_22109);
xor U23109 (N_23109,N_22047,N_22320);
nor U23110 (N_23110,N_21122,N_21460);
and U23111 (N_23111,N_22243,N_21087);
nor U23112 (N_23112,N_21512,N_21849);
nand U23113 (N_23113,N_21211,N_21072);
xnor U23114 (N_23114,N_21403,N_21808);
nand U23115 (N_23115,N_21697,N_21710);
and U23116 (N_23116,N_21322,N_22471);
or U23117 (N_23117,N_22282,N_21035);
nor U23118 (N_23118,N_21993,N_22189);
nand U23119 (N_23119,N_22126,N_21099);
nor U23120 (N_23120,N_21787,N_21282);
and U23121 (N_23121,N_21498,N_21089);
or U23122 (N_23122,N_21516,N_21311);
xnor U23123 (N_23123,N_21635,N_22428);
or U23124 (N_23124,N_21476,N_21766);
xor U23125 (N_23125,N_22231,N_21477);
nor U23126 (N_23126,N_21608,N_21033);
nor U23127 (N_23127,N_21770,N_21247);
or U23128 (N_23128,N_22067,N_22010);
or U23129 (N_23129,N_22271,N_22196);
or U23130 (N_23130,N_21535,N_21810);
and U23131 (N_23131,N_21572,N_21112);
or U23132 (N_23132,N_21659,N_21421);
nor U23133 (N_23133,N_21642,N_21452);
nor U23134 (N_23134,N_22251,N_22044);
xnor U23135 (N_23135,N_21284,N_22300);
nor U23136 (N_23136,N_21078,N_21248);
nor U23137 (N_23137,N_21464,N_22491);
nand U23138 (N_23138,N_21553,N_22229);
nor U23139 (N_23139,N_22259,N_21586);
nand U23140 (N_23140,N_22289,N_21218);
nand U23141 (N_23141,N_21546,N_21844);
nand U23142 (N_23142,N_22234,N_22240);
xnor U23143 (N_23143,N_21481,N_21203);
nand U23144 (N_23144,N_21669,N_21471);
nor U23145 (N_23145,N_21381,N_21986);
nand U23146 (N_23146,N_21933,N_21948);
nand U23147 (N_23147,N_21339,N_21906);
nand U23148 (N_23148,N_21551,N_21618);
xnor U23149 (N_23149,N_22314,N_21084);
xor U23150 (N_23150,N_21815,N_21547);
or U23151 (N_23151,N_21875,N_21860);
and U23152 (N_23152,N_22158,N_21509);
and U23153 (N_23153,N_21134,N_22127);
nor U23154 (N_23154,N_21128,N_21207);
or U23155 (N_23155,N_21229,N_21255);
or U23156 (N_23156,N_21522,N_21442);
xor U23157 (N_23157,N_21682,N_22179);
nand U23158 (N_23158,N_21918,N_22276);
nand U23159 (N_23159,N_22137,N_21210);
nand U23160 (N_23160,N_21096,N_21384);
or U23161 (N_23161,N_21904,N_21676);
and U23162 (N_23162,N_21856,N_21412);
nor U23163 (N_23163,N_21729,N_21651);
nor U23164 (N_23164,N_22222,N_21735);
or U23165 (N_23165,N_21760,N_21267);
nor U23166 (N_23166,N_22036,N_22418);
nand U23167 (N_23167,N_21107,N_21447);
xnor U23168 (N_23168,N_21590,N_21520);
xor U23169 (N_23169,N_22166,N_21458);
or U23170 (N_23170,N_21649,N_21678);
nor U23171 (N_23171,N_22073,N_21665);
xnor U23172 (N_23172,N_21521,N_21620);
or U23173 (N_23173,N_21441,N_21004);
xor U23174 (N_23174,N_21029,N_21670);
nand U23175 (N_23175,N_21523,N_21852);
xnor U23176 (N_23176,N_21564,N_22005);
nand U23177 (N_23177,N_22088,N_21426);
or U23178 (N_23178,N_21591,N_22467);
and U23179 (N_23179,N_21548,N_22362);
nor U23180 (N_23180,N_22329,N_21338);
xnor U23181 (N_23181,N_22256,N_21552);
or U23182 (N_23182,N_21734,N_21580);
nand U23183 (N_23183,N_21691,N_22054);
or U23184 (N_23184,N_21794,N_21873);
and U23185 (N_23185,N_21195,N_21679);
or U23186 (N_23186,N_21355,N_21208);
or U23187 (N_23187,N_21380,N_21793);
nand U23188 (N_23188,N_22411,N_22117);
nand U23189 (N_23189,N_21749,N_21979);
or U23190 (N_23190,N_22242,N_22204);
or U23191 (N_23191,N_21892,N_22286);
xnor U23192 (N_23192,N_22400,N_22475);
nand U23193 (N_23193,N_21088,N_22025);
nor U23194 (N_23194,N_21624,N_21434);
or U23195 (N_23195,N_21290,N_21301);
or U23196 (N_23196,N_21689,N_21349);
nand U23197 (N_23197,N_21953,N_21015);
or U23198 (N_23198,N_22318,N_21664);
xnor U23199 (N_23199,N_21751,N_21884);
nor U23200 (N_23200,N_21554,N_22398);
nand U23201 (N_23201,N_21151,N_21032);
and U23202 (N_23202,N_22093,N_21610);
xnor U23203 (N_23203,N_21667,N_21357);
xnor U23204 (N_23204,N_21224,N_21058);
and U23205 (N_23205,N_22441,N_22026);
nand U23206 (N_23206,N_22351,N_21490);
nand U23207 (N_23207,N_22419,N_21870);
or U23208 (N_23208,N_21615,N_21414);
nand U23209 (N_23209,N_21389,N_21605);
or U23210 (N_23210,N_22154,N_21484);
and U23211 (N_23211,N_22365,N_22029);
or U23212 (N_23212,N_21630,N_21780);
and U23213 (N_23213,N_21423,N_22331);
nand U23214 (N_23214,N_21726,N_22207);
nand U23215 (N_23215,N_22064,N_21611);
and U23216 (N_23216,N_21633,N_21584);
xnor U23217 (N_23217,N_22347,N_22449);
and U23218 (N_23218,N_21411,N_21663);
nor U23219 (N_23219,N_21784,N_21813);
and U23220 (N_23220,N_22485,N_21228);
nor U23221 (N_23221,N_21220,N_21786);
nor U23222 (N_23222,N_21307,N_22344);
nand U23223 (N_23223,N_22120,N_21180);
nor U23224 (N_23224,N_22283,N_21699);
nor U23225 (N_23225,N_21556,N_21440);
xnor U23226 (N_23226,N_22052,N_21368);
xnor U23227 (N_23227,N_22392,N_21791);
nor U23228 (N_23228,N_22232,N_22284);
nand U23229 (N_23229,N_22297,N_21263);
nand U23230 (N_23230,N_21152,N_22169);
or U23231 (N_23231,N_22223,N_22366);
and U23232 (N_23232,N_21631,N_22487);
and U23233 (N_23233,N_22241,N_22484);
xor U23234 (N_23234,N_22157,N_21358);
or U23235 (N_23235,N_21011,N_21239);
xnor U23236 (N_23236,N_21416,N_21579);
xor U23237 (N_23237,N_21908,N_21570);
or U23238 (N_23238,N_21299,N_21974);
or U23239 (N_23239,N_21026,N_22020);
xor U23240 (N_23240,N_22226,N_21502);
nand U23241 (N_23241,N_21732,N_22302);
nand U23242 (N_23242,N_21946,N_21257);
and U23243 (N_23243,N_21395,N_21527);
or U23244 (N_23244,N_21737,N_21814);
nand U23245 (N_23245,N_22012,N_22267);
or U23246 (N_23246,N_21655,N_21119);
or U23247 (N_23247,N_21574,N_21532);
and U23248 (N_23248,N_22434,N_21700);
xor U23249 (N_23249,N_22304,N_22124);
xnor U23250 (N_23250,N_21813,N_22081);
nand U23251 (N_23251,N_22032,N_21742);
xnor U23252 (N_23252,N_21776,N_22132);
xnor U23253 (N_23253,N_21110,N_21809);
or U23254 (N_23254,N_21355,N_21247);
nand U23255 (N_23255,N_22296,N_21775);
nand U23256 (N_23256,N_22446,N_21766);
nor U23257 (N_23257,N_21292,N_21316);
xnor U23258 (N_23258,N_21654,N_21938);
or U23259 (N_23259,N_21674,N_21539);
or U23260 (N_23260,N_21230,N_21926);
xor U23261 (N_23261,N_21981,N_22232);
or U23262 (N_23262,N_21222,N_21119);
nor U23263 (N_23263,N_22286,N_21154);
xnor U23264 (N_23264,N_22426,N_21963);
nand U23265 (N_23265,N_22487,N_22475);
and U23266 (N_23266,N_21395,N_21581);
or U23267 (N_23267,N_21564,N_22421);
and U23268 (N_23268,N_22497,N_21616);
nand U23269 (N_23269,N_21225,N_21211);
nor U23270 (N_23270,N_22470,N_21292);
xnor U23271 (N_23271,N_21949,N_21634);
or U23272 (N_23272,N_21147,N_22447);
or U23273 (N_23273,N_21082,N_21493);
and U23274 (N_23274,N_22209,N_22348);
xnor U23275 (N_23275,N_22238,N_22376);
nand U23276 (N_23276,N_22443,N_21343);
or U23277 (N_23277,N_21270,N_21919);
or U23278 (N_23278,N_21383,N_21187);
nor U23279 (N_23279,N_21643,N_21138);
and U23280 (N_23280,N_21618,N_22386);
xor U23281 (N_23281,N_21373,N_21958);
nand U23282 (N_23282,N_21521,N_22422);
or U23283 (N_23283,N_21937,N_21162);
or U23284 (N_23284,N_21933,N_21197);
xnor U23285 (N_23285,N_21712,N_22335);
nor U23286 (N_23286,N_21140,N_22489);
xor U23287 (N_23287,N_21095,N_22280);
nor U23288 (N_23288,N_21618,N_21662);
nand U23289 (N_23289,N_22212,N_21571);
xnor U23290 (N_23290,N_21584,N_22387);
or U23291 (N_23291,N_22026,N_21249);
and U23292 (N_23292,N_21846,N_22241);
nor U23293 (N_23293,N_22158,N_21647);
or U23294 (N_23294,N_21724,N_21789);
and U23295 (N_23295,N_22347,N_21514);
nor U23296 (N_23296,N_22109,N_22371);
and U23297 (N_23297,N_21721,N_22478);
and U23298 (N_23298,N_21565,N_22487);
and U23299 (N_23299,N_22082,N_22050);
xnor U23300 (N_23300,N_22331,N_21681);
nand U23301 (N_23301,N_22243,N_21569);
and U23302 (N_23302,N_22358,N_21209);
xor U23303 (N_23303,N_21349,N_21337);
xor U23304 (N_23304,N_21694,N_21814);
nand U23305 (N_23305,N_22081,N_21351);
xnor U23306 (N_23306,N_21097,N_21924);
xor U23307 (N_23307,N_21090,N_22417);
and U23308 (N_23308,N_21603,N_22188);
nand U23309 (N_23309,N_22210,N_21019);
xnor U23310 (N_23310,N_22285,N_21975);
nor U23311 (N_23311,N_21736,N_22042);
or U23312 (N_23312,N_21262,N_21958);
nand U23313 (N_23313,N_22324,N_21931);
xnor U23314 (N_23314,N_22472,N_21513);
nand U23315 (N_23315,N_21382,N_21208);
or U23316 (N_23316,N_21633,N_21599);
nor U23317 (N_23317,N_21299,N_21808);
nor U23318 (N_23318,N_22150,N_21370);
and U23319 (N_23319,N_21272,N_22439);
and U23320 (N_23320,N_22149,N_21603);
and U23321 (N_23321,N_22096,N_21085);
or U23322 (N_23322,N_22297,N_21256);
or U23323 (N_23323,N_21505,N_21247);
nand U23324 (N_23324,N_22033,N_21959);
or U23325 (N_23325,N_21627,N_21287);
xnor U23326 (N_23326,N_22271,N_21444);
or U23327 (N_23327,N_21468,N_22469);
nor U23328 (N_23328,N_21516,N_22369);
nand U23329 (N_23329,N_21833,N_21468);
and U23330 (N_23330,N_22235,N_22465);
nor U23331 (N_23331,N_21085,N_21249);
and U23332 (N_23332,N_22333,N_21992);
and U23333 (N_23333,N_22090,N_21993);
nand U23334 (N_23334,N_21102,N_21002);
and U23335 (N_23335,N_21463,N_22295);
nor U23336 (N_23336,N_21740,N_22381);
xor U23337 (N_23337,N_21263,N_21190);
xnor U23338 (N_23338,N_21199,N_21929);
xnor U23339 (N_23339,N_22118,N_22364);
xor U23340 (N_23340,N_21239,N_21873);
xor U23341 (N_23341,N_21897,N_21388);
nor U23342 (N_23342,N_21824,N_21939);
and U23343 (N_23343,N_21832,N_21133);
or U23344 (N_23344,N_22135,N_22475);
nor U23345 (N_23345,N_21266,N_21152);
xor U23346 (N_23346,N_21763,N_21732);
nand U23347 (N_23347,N_22451,N_22286);
nor U23348 (N_23348,N_22431,N_21919);
xnor U23349 (N_23349,N_21086,N_21389);
and U23350 (N_23350,N_21826,N_21410);
xnor U23351 (N_23351,N_21401,N_21346);
and U23352 (N_23352,N_21988,N_21697);
nand U23353 (N_23353,N_22157,N_22282);
nand U23354 (N_23354,N_21095,N_22289);
or U23355 (N_23355,N_21430,N_21805);
or U23356 (N_23356,N_21940,N_21563);
xor U23357 (N_23357,N_21671,N_21819);
or U23358 (N_23358,N_22387,N_22166);
nor U23359 (N_23359,N_21486,N_21720);
nor U23360 (N_23360,N_21474,N_21482);
nor U23361 (N_23361,N_21153,N_22316);
nand U23362 (N_23362,N_21342,N_22369);
nand U23363 (N_23363,N_22138,N_21637);
and U23364 (N_23364,N_22042,N_22210);
nand U23365 (N_23365,N_21083,N_21381);
nor U23366 (N_23366,N_22118,N_22312);
and U23367 (N_23367,N_22093,N_21213);
or U23368 (N_23368,N_21965,N_21615);
or U23369 (N_23369,N_21323,N_21306);
xnor U23370 (N_23370,N_21268,N_21838);
nor U23371 (N_23371,N_22067,N_21469);
nor U23372 (N_23372,N_21850,N_21856);
or U23373 (N_23373,N_21538,N_21065);
or U23374 (N_23374,N_21937,N_22046);
and U23375 (N_23375,N_21960,N_21430);
nand U23376 (N_23376,N_21722,N_21851);
and U23377 (N_23377,N_21588,N_22134);
nor U23378 (N_23378,N_21330,N_22457);
nand U23379 (N_23379,N_22105,N_21392);
xor U23380 (N_23380,N_22349,N_21194);
or U23381 (N_23381,N_21068,N_21532);
nand U23382 (N_23382,N_21451,N_22332);
or U23383 (N_23383,N_21571,N_21365);
or U23384 (N_23384,N_22095,N_21020);
and U23385 (N_23385,N_21221,N_22430);
xnor U23386 (N_23386,N_22331,N_21848);
xor U23387 (N_23387,N_21258,N_22132);
and U23388 (N_23388,N_21032,N_21599);
and U23389 (N_23389,N_22085,N_21460);
nor U23390 (N_23390,N_22123,N_21884);
and U23391 (N_23391,N_21773,N_21245);
xnor U23392 (N_23392,N_21351,N_22147);
or U23393 (N_23393,N_21174,N_22466);
nand U23394 (N_23394,N_21715,N_21375);
or U23395 (N_23395,N_21907,N_22072);
xor U23396 (N_23396,N_21276,N_21979);
nand U23397 (N_23397,N_21452,N_21193);
nand U23398 (N_23398,N_22124,N_21625);
and U23399 (N_23399,N_21038,N_21537);
nand U23400 (N_23400,N_21225,N_21195);
and U23401 (N_23401,N_21352,N_21787);
nand U23402 (N_23402,N_22220,N_22414);
nand U23403 (N_23403,N_21248,N_21502);
nor U23404 (N_23404,N_21755,N_21601);
nor U23405 (N_23405,N_21184,N_21430);
xnor U23406 (N_23406,N_21477,N_22242);
xor U23407 (N_23407,N_21432,N_21785);
and U23408 (N_23408,N_22323,N_21685);
nand U23409 (N_23409,N_22417,N_22495);
nand U23410 (N_23410,N_21879,N_21725);
xnor U23411 (N_23411,N_22224,N_21364);
nand U23412 (N_23412,N_21056,N_21747);
nand U23413 (N_23413,N_21247,N_21062);
and U23414 (N_23414,N_21147,N_22163);
nand U23415 (N_23415,N_21316,N_22465);
or U23416 (N_23416,N_22060,N_21186);
or U23417 (N_23417,N_21205,N_21633);
or U23418 (N_23418,N_22010,N_21830);
and U23419 (N_23419,N_21676,N_22096);
nand U23420 (N_23420,N_21387,N_21339);
nand U23421 (N_23421,N_21027,N_21315);
nor U23422 (N_23422,N_22119,N_21533);
xor U23423 (N_23423,N_22080,N_22486);
nand U23424 (N_23424,N_21348,N_21120);
nand U23425 (N_23425,N_21383,N_21342);
and U23426 (N_23426,N_22046,N_21045);
and U23427 (N_23427,N_22427,N_22178);
or U23428 (N_23428,N_21386,N_22369);
nand U23429 (N_23429,N_21895,N_21111);
nand U23430 (N_23430,N_21009,N_21527);
nand U23431 (N_23431,N_21700,N_21746);
or U23432 (N_23432,N_21157,N_22495);
xnor U23433 (N_23433,N_22004,N_22255);
or U23434 (N_23434,N_22317,N_21564);
xor U23435 (N_23435,N_21825,N_21959);
nand U23436 (N_23436,N_22407,N_21376);
or U23437 (N_23437,N_21308,N_21332);
nor U23438 (N_23438,N_22489,N_22195);
and U23439 (N_23439,N_21292,N_21417);
and U23440 (N_23440,N_22034,N_21415);
nand U23441 (N_23441,N_21597,N_21668);
nor U23442 (N_23442,N_22048,N_22178);
or U23443 (N_23443,N_21706,N_21032);
nor U23444 (N_23444,N_21050,N_21697);
and U23445 (N_23445,N_21733,N_21415);
xor U23446 (N_23446,N_22121,N_22329);
xor U23447 (N_23447,N_21765,N_21270);
and U23448 (N_23448,N_22110,N_22097);
and U23449 (N_23449,N_21059,N_21735);
nor U23450 (N_23450,N_21514,N_22207);
xor U23451 (N_23451,N_22084,N_21512);
and U23452 (N_23452,N_21147,N_21001);
and U23453 (N_23453,N_22167,N_22403);
or U23454 (N_23454,N_22418,N_21127);
and U23455 (N_23455,N_21216,N_21239);
or U23456 (N_23456,N_21235,N_21304);
nor U23457 (N_23457,N_21128,N_21536);
or U23458 (N_23458,N_21864,N_22095);
xor U23459 (N_23459,N_21278,N_21673);
xnor U23460 (N_23460,N_21045,N_21060);
or U23461 (N_23461,N_21581,N_21537);
nor U23462 (N_23462,N_21946,N_21663);
xor U23463 (N_23463,N_21315,N_21128);
and U23464 (N_23464,N_22105,N_22151);
xnor U23465 (N_23465,N_22002,N_21179);
nor U23466 (N_23466,N_22338,N_22248);
xnor U23467 (N_23467,N_21552,N_22335);
or U23468 (N_23468,N_22151,N_22450);
nand U23469 (N_23469,N_22200,N_21712);
nand U23470 (N_23470,N_21214,N_22139);
or U23471 (N_23471,N_22447,N_21087);
xnor U23472 (N_23472,N_21043,N_21493);
or U23473 (N_23473,N_21502,N_22456);
nor U23474 (N_23474,N_21432,N_21415);
and U23475 (N_23475,N_21251,N_21297);
nand U23476 (N_23476,N_21355,N_21338);
xnor U23477 (N_23477,N_22191,N_21653);
and U23478 (N_23478,N_22116,N_21303);
nand U23479 (N_23479,N_21024,N_22488);
nand U23480 (N_23480,N_21464,N_21185);
nor U23481 (N_23481,N_21769,N_22002);
nand U23482 (N_23482,N_21634,N_21268);
nand U23483 (N_23483,N_22250,N_21419);
nand U23484 (N_23484,N_21086,N_22150);
or U23485 (N_23485,N_22375,N_22281);
and U23486 (N_23486,N_21203,N_22294);
or U23487 (N_23487,N_21321,N_22258);
xor U23488 (N_23488,N_21614,N_22278);
or U23489 (N_23489,N_21005,N_22461);
and U23490 (N_23490,N_21559,N_21353);
or U23491 (N_23491,N_22106,N_21571);
or U23492 (N_23492,N_21244,N_22473);
xnor U23493 (N_23493,N_22456,N_21791);
nand U23494 (N_23494,N_22393,N_21781);
nor U23495 (N_23495,N_22333,N_21011);
xor U23496 (N_23496,N_22172,N_21255);
nand U23497 (N_23497,N_21037,N_22443);
xnor U23498 (N_23498,N_21612,N_21239);
nor U23499 (N_23499,N_22390,N_22131);
nor U23500 (N_23500,N_22302,N_21938);
nor U23501 (N_23501,N_22042,N_21379);
nor U23502 (N_23502,N_21007,N_21938);
and U23503 (N_23503,N_21372,N_22467);
xor U23504 (N_23504,N_21858,N_21975);
and U23505 (N_23505,N_21184,N_21001);
xnor U23506 (N_23506,N_21633,N_22128);
and U23507 (N_23507,N_22347,N_22119);
and U23508 (N_23508,N_21056,N_22423);
nand U23509 (N_23509,N_22499,N_22260);
nor U23510 (N_23510,N_22132,N_21619);
xnor U23511 (N_23511,N_21357,N_21745);
nor U23512 (N_23512,N_21833,N_21995);
nand U23513 (N_23513,N_21911,N_22301);
or U23514 (N_23514,N_21790,N_21661);
nor U23515 (N_23515,N_21501,N_21730);
xor U23516 (N_23516,N_22415,N_21003);
nand U23517 (N_23517,N_22380,N_21363);
and U23518 (N_23518,N_21338,N_21444);
or U23519 (N_23519,N_21889,N_21370);
nand U23520 (N_23520,N_21760,N_21789);
or U23521 (N_23521,N_21061,N_21967);
nand U23522 (N_23522,N_22177,N_21815);
nor U23523 (N_23523,N_21389,N_21730);
nor U23524 (N_23524,N_22280,N_21728);
nor U23525 (N_23525,N_22083,N_21895);
or U23526 (N_23526,N_21501,N_21391);
xor U23527 (N_23527,N_22437,N_22393);
or U23528 (N_23528,N_22085,N_22269);
or U23529 (N_23529,N_21435,N_21912);
and U23530 (N_23530,N_21136,N_21367);
and U23531 (N_23531,N_21388,N_22439);
xnor U23532 (N_23532,N_22023,N_21569);
nor U23533 (N_23533,N_21476,N_21504);
or U23534 (N_23534,N_22013,N_21907);
or U23535 (N_23535,N_21465,N_22216);
nor U23536 (N_23536,N_21637,N_22008);
and U23537 (N_23537,N_21746,N_22414);
nand U23538 (N_23538,N_21745,N_22163);
xnor U23539 (N_23539,N_21102,N_21562);
nand U23540 (N_23540,N_21665,N_21624);
or U23541 (N_23541,N_21730,N_22256);
xnor U23542 (N_23542,N_21290,N_21155);
nor U23543 (N_23543,N_22074,N_21285);
or U23544 (N_23544,N_22492,N_21091);
or U23545 (N_23545,N_21679,N_21528);
or U23546 (N_23546,N_21548,N_21387);
nand U23547 (N_23547,N_22388,N_21058);
and U23548 (N_23548,N_21030,N_22061);
nor U23549 (N_23549,N_21179,N_21449);
xnor U23550 (N_23550,N_21920,N_21826);
nand U23551 (N_23551,N_21764,N_21492);
or U23552 (N_23552,N_21529,N_22043);
or U23553 (N_23553,N_21262,N_21419);
or U23554 (N_23554,N_21996,N_21257);
or U23555 (N_23555,N_22305,N_21564);
nand U23556 (N_23556,N_22440,N_21229);
and U23557 (N_23557,N_21617,N_21068);
or U23558 (N_23558,N_21148,N_22104);
or U23559 (N_23559,N_21964,N_22035);
nand U23560 (N_23560,N_21550,N_22118);
nor U23561 (N_23561,N_22183,N_21456);
xor U23562 (N_23562,N_21997,N_21636);
nor U23563 (N_23563,N_21756,N_21435);
nand U23564 (N_23564,N_21534,N_21825);
and U23565 (N_23565,N_21716,N_21102);
nor U23566 (N_23566,N_21307,N_22214);
xnor U23567 (N_23567,N_22329,N_21671);
nor U23568 (N_23568,N_22123,N_21284);
xor U23569 (N_23569,N_22440,N_21251);
nand U23570 (N_23570,N_21230,N_21078);
xnor U23571 (N_23571,N_21105,N_22157);
nand U23572 (N_23572,N_22319,N_22382);
or U23573 (N_23573,N_21318,N_22035);
or U23574 (N_23574,N_21045,N_21085);
xnor U23575 (N_23575,N_21844,N_21026);
xor U23576 (N_23576,N_21353,N_21321);
and U23577 (N_23577,N_22054,N_22142);
and U23578 (N_23578,N_21425,N_21928);
or U23579 (N_23579,N_22316,N_21638);
and U23580 (N_23580,N_21665,N_21536);
xor U23581 (N_23581,N_21960,N_22176);
xor U23582 (N_23582,N_21426,N_21125);
nand U23583 (N_23583,N_21837,N_21136);
nand U23584 (N_23584,N_22008,N_21988);
or U23585 (N_23585,N_22074,N_21089);
xnor U23586 (N_23586,N_21712,N_22220);
xnor U23587 (N_23587,N_21525,N_21722);
and U23588 (N_23588,N_22322,N_21108);
xnor U23589 (N_23589,N_21683,N_22042);
xor U23590 (N_23590,N_21584,N_21250);
nor U23591 (N_23591,N_21873,N_21961);
nand U23592 (N_23592,N_21035,N_21321);
or U23593 (N_23593,N_22493,N_21567);
nor U23594 (N_23594,N_21355,N_21889);
and U23595 (N_23595,N_21524,N_22059);
nand U23596 (N_23596,N_21896,N_21538);
nand U23597 (N_23597,N_21786,N_22371);
and U23598 (N_23598,N_21869,N_21629);
or U23599 (N_23599,N_21160,N_22007);
or U23600 (N_23600,N_21973,N_22285);
or U23601 (N_23601,N_22227,N_22000);
nand U23602 (N_23602,N_21459,N_21424);
nor U23603 (N_23603,N_22470,N_21562);
nand U23604 (N_23604,N_21551,N_21233);
or U23605 (N_23605,N_21802,N_22070);
nor U23606 (N_23606,N_22022,N_21540);
or U23607 (N_23607,N_21453,N_21360);
nand U23608 (N_23608,N_22049,N_21955);
nor U23609 (N_23609,N_22245,N_22355);
nand U23610 (N_23610,N_21365,N_22449);
and U23611 (N_23611,N_21792,N_21669);
xor U23612 (N_23612,N_21073,N_21790);
and U23613 (N_23613,N_21836,N_21556);
nand U23614 (N_23614,N_21231,N_21243);
xor U23615 (N_23615,N_21786,N_21569);
and U23616 (N_23616,N_22259,N_21668);
and U23617 (N_23617,N_21626,N_21889);
nand U23618 (N_23618,N_22350,N_22465);
xnor U23619 (N_23619,N_21408,N_21676);
or U23620 (N_23620,N_21849,N_22173);
and U23621 (N_23621,N_21728,N_22309);
or U23622 (N_23622,N_21490,N_22155);
nand U23623 (N_23623,N_21370,N_22379);
or U23624 (N_23624,N_21475,N_22181);
xor U23625 (N_23625,N_21092,N_21394);
nand U23626 (N_23626,N_21059,N_21240);
or U23627 (N_23627,N_21413,N_22433);
xnor U23628 (N_23628,N_21091,N_22138);
and U23629 (N_23629,N_21686,N_21643);
nand U23630 (N_23630,N_22388,N_21674);
xor U23631 (N_23631,N_21035,N_21393);
nor U23632 (N_23632,N_21025,N_21303);
xnor U23633 (N_23633,N_21657,N_21708);
or U23634 (N_23634,N_21650,N_22209);
and U23635 (N_23635,N_21503,N_22131);
nor U23636 (N_23636,N_21776,N_21750);
and U23637 (N_23637,N_22040,N_22348);
or U23638 (N_23638,N_21299,N_21446);
xnor U23639 (N_23639,N_22126,N_21231);
or U23640 (N_23640,N_22025,N_21981);
and U23641 (N_23641,N_21305,N_22031);
and U23642 (N_23642,N_21098,N_22257);
nor U23643 (N_23643,N_21015,N_22434);
or U23644 (N_23644,N_22327,N_22216);
xnor U23645 (N_23645,N_21662,N_21564);
nor U23646 (N_23646,N_21805,N_21057);
nand U23647 (N_23647,N_22333,N_21370);
and U23648 (N_23648,N_21232,N_22132);
xnor U23649 (N_23649,N_21962,N_21882);
nand U23650 (N_23650,N_21745,N_21039);
nand U23651 (N_23651,N_22173,N_21810);
and U23652 (N_23652,N_22439,N_22254);
xnor U23653 (N_23653,N_21627,N_22482);
nor U23654 (N_23654,N_21458,N_21023);
nor U23655 (N_23655,N_21691,N_22239);
and U23656 (N_23656,N_21250,N_21972);
nor U23657 (N_23657,N_22171,N_21732);
or U23658 (N_23658,N_21823,N_22364);
xor U23659 (N_23659,N_22344,N_22271);
nor U23660 (N_23660,N_21888,N_21595);
xnor U23661 (N_23661,N_21644,N_21442);
nor U23662 (N_23662,N_21391,N_21659);
nand U23663 (N_23663,N_21911,N_21869);
xor U23664 (N_23664,N_22168,N_21125);
xor U23665 (N_23665,N_22274,N_21148);
xnor U23666 (N_23666,N_21165,N_22207);
and U23667 (N_23667,N_21076,N_22307);
xor U23668 (N_23668,N_22022,N_22375);
xnor U23669 (N_23669,N_22218,N_21088);
nand U23670 (N_23670,N_21538,N_22047);
and U23671 (N_23671,N_21974,N_22277);
nor U23672 (N_23672,N_22369,N_21185);
and U23673 (N_23673,N_21530,N_21952);
nor U23674 (N_23674,N_21467,N_21296);
or U23675 (N_23675,N_22091,N_21226);
xor U23676 (N_23676,N_21384,N_21544);
nand U23677 (N_23677,N_21544,N_21317);
and U23678 (N_23678,N_21891,N_21754);
nor U23679 (N_23679,N_21149,N_22352);
or U23680 (N_23680,N_21700,N_21379);
nor U23681 (N_23681,N_21555,N_22051);
or U23682 (N_23682,N_22049,N_22087);
and U23683 (N_23683,N_21815,N_22200);
xnor U23684 (N_23684,N_21579,N_22385);
xor U23685 (N_23685,N_22126,N_21375);
xor U23686 (N_23686,N_21323,N_21954);
or U23687 (N_23687,N_22082,N_21996);
nor U23688 (N_23688,N_21404,N_22172);
nand U23689 (N_23689,N_22259,N_21473);
nor U23690 (N_23690,N_21546,N_21767);
nor U23691 (N_23691,N_22491,N_21822);
nor U23692 (N_23692,N_21655,N_21970);
or U23693 (N_23693,N_21845,N_22372);
or U23694 (N_23694,N_22310,N_21815);
nor U23695 (N_23695,N_22308,N_21119);
and U23696 (N_23696,N_22281,N_22185);
nor U23697 (N_23697,N_21134,N_21390);
xnor U23698 (N_23698,N_21095,N_21295);
nor U23699 (N_23699,N_22471,N_21282);
or U23700 (N_23700,N_21592,N_22301);
or U23701 (N_23701,N_21948,N_21461);
and U23702 (N_23702,N_22076,N_21359);
xor U23703 (N_23703,N_21025,N_22001);
nor U23704 (N_23704,N_22435,N_21938);
nor U23705 (N_23705,N_21825,N_22377);
nand U23706 (N_23706,N_21775,N_21553);
or U23707 (N_23707,N_22451,N_21922);
or U23708 (N_23708,N_22299,N_22273);
or U23709 (N_23709,N_21247,N_21099);
and U23710 (N_23710,N_22285,N_22116);
xor U23711 (N_23711,N_21731,N_21609);
and U23712 (N_23712,N_21297,N_21726);
xor U23713 (N_23713,N_21361,N_21352);
nor U23714 (N_23714,N_21469,N_21245);
xor U23715 (N_23715,N_21732,N_21541);
nand U23716 (N_23716,N_22330,N_22078);
xnor U23717 (N_23717,N_21157,N_22007);
xor U23718 (N_23718,N_22287,N_21328);
xor U23719 (N_23719,N_21011,N_21350);
or U23720 (N_23720,N_21534,N_21752);
or U23721 (N_23721,N_21030,N_22175);
nor U23722 (N_23722,N_21915,N_21352);
and U23723 (N_23723,N_21957,N_21410);
and U23724 (N_23724,N_21762,N_21715);
xnor U23725 (N_23725,N_21084,N_22498);
nand U23726 (N_23726,N_21450,N_21114);
or U23727 (N_23727,N_21261,N_21431);
nand U23728 (N_23728,N_22263,N_22184);
and U23729 (N_23729,N_22396,N_21051);
or U23730 (N_23730,N_22307,N_21544);
and U23731 (N_23731,N_21354,N_21945);
and U23732 (N_23732,N_22152,N_21570);
or U23733 (N_23733,N_21693,N_21987);
or U23734 (N_23734,N_21364,N_21043);
nand U23735 (N_23735,N_21139,N_21497);
and U23736 (N_23736,N_22035,N_21111);
or U23737 (N_23737,N_21319,N_21076);
nor U23738 (N_23738,N_21149,N_22394);
or U23739 (N_23739,N_21525,N_21102);
nor U23740 (N_23740,N_21376,N_21139);
xor U23741 (N_23741,N_21218,N_21304);
xor U23742 (N_23742,N_21495,N_22432);
and U23743 (N_23743,N_22377,N_21612);
nor U23744 (N_23744,N_22059,N_22168);
nand U23745 (N_23745,N_21640,N_21704);
or U23746 (N_23746,N_21904,N_21354);
nand U23747 (N_23747,N_22130,N_21732);
nand U23748 (N_23748,N_21350,N_21927);
xor U23749 (N_23749,N_21426,N_21855);
or U23750 (N_23750,N_21065,N_21947);
or U23751 (N_23751,N_21726,N_21698);
xor U23752 (N_23752,N_21470,N_21965);
xnor U23753 (N_23753,N_22426,N_21786);
xnor U23754 (N_23754,N_21624,N_21832);
nor U23755 (N_23755,N_22198,N_21848);
and U23756 (N_23756,N_21851,N_21341);
xnor U23757 (N_23757,N_21556,N_22318);
or U23758 (N_23758,N_22425,N_21829);
nand U23759 (N_23759,N_21354,N_22075);
nor U23760 (N_23760,N_21291,N_21186);
or U23761 (N_23761,N_22017,N_21760);
nand U23762 (N_23762,N_21070,N_21898);
nor U23763 (N_23763,N_21302,N_22352);
or U23764 (N_23764,N_21195,N_21932);
or U23765 (N_23765,N_22137,N_21981);
or U23766 (N_23766,N_22184,N_22103);
or U23767 (N_23767,N_22282,N_21743);
xnor U23768 (N_23768,N_21232,N_21943);
nor U23769 (N_23769,N_21790,N_21181);
nor U23770 (N_23770,N_21061,N_21203);
or U23771 (N_23771,N_21915,N_21295);
and U23772 (N_23772,N_21230,N_22198);
xor U23773 (N_23773,N_21557,N_22212);
or U23774 (N_23774,N_22323,N_21842);
xor U23775 (N_23775,N_22434,N_22098);
nor U23776 (N_23776,N_22444,N_21486);
xor U23777 (N_23777,N_21744,N_21136);
nand U23778 (N_23778,N_22015,N_21036);
or U23779 (N_23779,N_22112,N_21423);
and U23780 (N_23780,N_21312,N_21521);
nand U23781 (N_23781,N_22109,N_21632);
or U23782 (N_23782,N_22402,N_22494);
nor U23783 (N_23783,N_21824,N_21222);
or U23784 (N_23784,N_22236,N_22393);
and U23785 (N_23785,N_21772,N_22295);
xor U23786 (N_23786,N_21589,N_21576);
or U23787 (N_23787,N_21484,N_22124);
nor U23788 (N_23788,N_21618,N_21515);
and U23789 (N_23789,N_21458,N_21455);
and U23790 (N_23790,N_21770,N_22403);
nor U23791 (N_23791,N_21030,N_21495);
nand U23792 (N_23792,N_21197,N_22041);
nor U23793 (N_23793,N_21138,N_21481);
xnor U23794 (N_23794,N_21084,N_22289);
xor U23795 (N_23795,N_21832,N_22131);
nand U23796 (N_23796,N_21639,N_21484);
xnor U23797 (N_23797,N_21111,N_22234);
nor U23798 (N_23798,N_21188,N_22237);
xor U23799 (N_23799,N_21932,N_21378);
and U23800 (N_23800,N_21914,N_21332);
xor U23801 (N_23801,N_21782,N_21520);
xnor U23802 (N_23802,N_21709,N_22087);
nand U23803 (N_23803,N_21379,N_21866);
nand U23804 (N_23804,N_21476,N_21512);
and U23805 (N_23805,N_21173,N_22422);
nor U23806 (N_23806,N_21698,N_22217);
or U23807 (N_23807,N_21468,N_22237);
and U23808 (N_23808,N_21429,N_21513);
nor U23809 (N_23809,N_21388,N_21164);
xor U23810 (N_23810,N_21085,N_21707);
or U23811 (N_23811,N_21029,N_21000);
and U23812 (N_23812,N_21209,N_22224);
xnor U23813 (N_23813,N_21241,N_22395);
or U23814 (N_23814,N_21381,N_21618);
or U23815 (N_23815,N_21896,N_21229);
xor U23816 (N_23816,N_21707,N_22380);
or U23817 (N_23817,N_21039,N_21238);
nand U23818 (N_23818,N_22479,N_21114);
xnor U23819 (N_23819,N_22140,N_21429);
xnor U23820 (N_23820,N_21960,N_21418);
or U23821 (N_23821,N_21022,N_21650);
nor U23822 (N_23822,N_21340,N_21824);
or U23823 (N_23823,N_22024,N_21908);
and U23824 (N_23824,N_21637,N_22381);
nor U23825 (N_23825,N_22441,N_21923);
nand U23826 (N_23826,N_22448,N_21457);
nor U23827 (N_23827,N_21172,N_21210);
xnor U23828 (N_23828,N_21526,N_22010);
or U23829 (N_23829,N_21962,N_21679);
and U23830 (N_23830,N_21277,N_22301);
nand U23831 (N_23831,N_21626,N_21888);
xnor U23832 (N_23832,N_22498,N_21913);
nor U23833 (N_23833,N_22084,N_21370);
nor U23834 (N_23834,N_22211,N_21518);
nand U23835 (N_23835,N_21435,N_22048);
nand U23836 (N_23836,N_21305,N_21299);
nand U23837 (N_23837,N_21641,N_22343);
or U23838 (N_23838,N_21171,N_21528);
xnor U23839 (N_23839,N_22291,N_22351);
nor U23840 (N_23840,N_21921,N_21006);
or U23841 (N_23841,N_21880,N_22370);
xor U23842 (N_23842,N_22165,N_21649);
xor U23843 (N_23843,N_21603,N_21927);
xnor U23844 (N_23844,N_21959,N_22023);
nand U23845 (N_23845,N_21394,N_22306);
nand U23846 (N_23846,N_21069,N_21005);
and U23847 (N_23847,N_21702,N_21015);
xnor U23848 (N_23848,N_21644,N_22326);
nand U23849 (N_23849,N_21568,N_22067);
and U23850 (N_23850,N_22443,N_21320);
or U23851 (N_23851,N_21576,N_21197);
nand U23852 (N_23852,N_21042,N_22156);
and U23853 (N_23853,N_22493,N_21783);
nor U23854 (N_23854,N_21114,N_22118);
or U23855 (N_23855,N_21297,N_22278);
nand U23856 (N_23856,N_21657,N_22263);
nand U23857 (N_23857,N_21576,N_21008);
nor U23858 (N_23858,N_22440,N_22420);
or U23859 (N_23859,N_21519,N_21729);
nor U23860 (N_23860,N_21312,N_21367);
xor U23861 (N_23861,N_21639,N_21647);
or U23862 (N_23862,N_21969,N_21384);
nor U23863 (N_23863,N_21432,N_21632);
and U23864 (N_23864,N_22477,N_21550);
xnor U23865 (N_23865,N_22386,N_22181);
xnor U23866 (N_23866,N_22478,N_21560);
and U23867 (N_23867,N_21176,N_21029);
xor U23868 (N_23868,N_21698,N_22198);
nand U23869 (N_23869,N_22412,N_21466);
xor U23870 (N_23870,N_21047,N_22440);
nand U23871 (N_23871,N_21404,N_21701);
or U23872 (N_23872,N_22269,N_22485);
and U23873 (N_23873,N_21014,N_21714);
and U23874 (N_23874,N_21919,N_21096);
xnor U23875 (N_23875,N_21082,N_22163);
nor U23876 (N_23876,N_21302,N_22393);
and U23877 (N_23877,N_21725,N_21410);
and U23878 (N_23878,N_21449,N_21694);
xnor U23879 (N_23879,N_21737,N_21057);
and U23880 (N_23880,N_22302,N_21643);
or U23881 (N_23881,N_22464,N_21324);
nand U23882 (N_23882,N_21863,N_21556);
nand U23883 (N_23883,N_21169,N_22467);
nand U23884 (N_23884,N_22142,N_21459);
and U23885 (N_23885,N_21735,N_22266);
nor U23886 (N_23886,N_22355,N_21356);
nand U23887 (N_23887,N_21504,N_22319);
nand U23888 (N_23888,N_21322,N_21963);
or U23889 (N_23889,N_22214,N_21214);
and U23890 (N_23890,N_21191,N_22151);
nor U23891 (N_23891,N_22372,N_21313);
nand U23892 (N_23892,N_22101,N_22453);
and U23893 (N_23893,N_21339,N_22309);
nor U23894 (N_23894,N_21602,N_21730);
nand U23895 (N_23895,N_22206,N_22078);
nor U23896 (N_23896,N_21224,N_21078);
or U23897 (N_23897,N_21835,N_22335);
nor U23898 (N_23898,N_22432,N_22163);
and U23899 (N_23899,N_22323,N_21834);
and U23900 (N_23900,N_21085,N_21029);
xor U23901 (N_23901,N_21521,N_21801);
xnor U23902 (N_23902,N_22181,N_22312);
or U23903 (N_23903,N_21861,N_22404);
nand U23904 (N_23904,N_21222,N_21098);
nor U23905 (N_23905,N_22222,N_22148);
or U23906 (N_23906,N_21239,N_21408);
and U23907 (N_23907,N_21982,N_21243);
or U23908 (N_23908,N_21773,N_22312);
nor U23909 (N_23909,N_21546,N_21519);
nor U23910 (N_23910,N_21129,N_21672);
and U23911 (N_23911,N_21773,N_21514);
nor U23912 (N_23912,N_22424,N_21096);
nor U23913 (N_23913,N_21594,N_21212);
xnor U23914 (N_23914,N_21577,N_21136);
and U23915 (N_23915,N_21544,N_21859);
nor U23916 (N_23916,N_21991,N_22315);
or U23917 (N_23917,N_21218,N_21688);
or U23918 (N_23918,N_21502,N_21591);
or U23919 (N_23919,N_21804,N_21485);
nor U23920 (N_23920,N_21481,N_21273);
xor U23921 (N_23921,N_21509,N_21056);
nand U23922 (N_23922,N_21389,N_21278);
or U23923 (N_23923,N_21369,N_21128);
nor U23924 (N_23924,N_22353,N_21270);
and U23925 (N_23925,N_21022,N_21750);
xnor U23926 (N_23926,N_21190,N_22029);
xnor U23927 (N_23927,N_21481,N_21031);
xor U23928 (N_23928,N_21665,N_22056);
nand U23929 (N_23929,N_22228,N_22481);
or U23930 (N_23930,N_21606,N_21917);
or U23931 (N_23931,N_21775,N_21549);
nor U23932 (N_23932,N_21140,N_22432);
xnor U23933 (N_23933,N_21169,N_21714);
or U23934 (N_23934,N_21532,N_21835);
and U23935 (N_23935,N_22140,N_22379);
nor U23936 (N_23936,N_21171,N_21889);
or U23937 (N_23937,N_22442,N_21522);
xor U23938 (N_23938,N_21900,N_21975);
or U23939 (N_23939,N_21924,N_22482);
or U23940 (N_23940,N_22324,N_21354);
nand U23941 (N_23941,N_21147,N_21188);
and U23942 (N_23942,N_21939,N_21003);
or U23943 (N_23943,N_21218,N_21995);
and U23944 (N_23944,N_21663,N_22425);
or U23945 (N_23945,N_21696,N_21901);
xor U23946 (N_23946,N_21814,N_21862);
and U23947 (N_23947,N_22051,N_21192);
nand U23948 (N_23948,N_21952,N_21914);
nor U23949 (N_23949,N_21517,N_21093);
nor U23950 (N_23950,N_21410,N_21239);
nand U23951 (N_23951,N_22474,N_21515);
and U23952 (N_23952,N_21460,N_21922);
nor U23953 (N_23953,N_22382,N_21526);
nor U23954 (N_23954,N_21899,N_21949);
nand U23955 (N_23955,N_21420,N_21426);
xnor U23956 (N_23956,N_22037,N_21218);
and U23957 (N_23957,N_21111,N_22382);
xor U23958 (N_23958,N_21449,N_21921);
nand U23959 (N_23959,N_22316,N_21277);
and U23960 (N_23960,N_22153,N_21340);
and U23961 (N_23961,N_21523,N_22075);
or U23962 (N_23962,N_22078,N_21869);
or U23963 (N_23963,N_21591,N_22128);
and U23964 (N_23964,N_22320,N_22166);
or U23965 (N_23965,N_22027,N_21540);
nand U23966 (N_23966,N_21392,N_22364);
nand U23967 (N_23967,N_21396,N_21177);
or U23968 (N_23968,N_21730,N_21195);
or U23969 (N_23969,N_21130,N_22044);
nand U23970 (N_23970,N_21882,N_22427);
nand U23971 (N_23971,N_22386,N_21800);
nor U23972 (N_23972,N_21396,N_22210);
xnor U23973 (N_23973,N_21204,N_22460);
nand U23974 (N_23974,N_22491,N_21152);
and U23975 (N_23975,N_21234,N_21018);
and U23976 (N_23976,N_21458,N_21048);
or U23977 (N_23977,N_21846,N_22336);
or U23978 (N_23978,N_22322,N_21998);
or U23979 (N_23979,N_21361,N_21215);
nor U23980 (N_23980,N_21227,N_21703);
nand U23981 (N_23981,N_21597,N_21500);
or U23982 (N_23982,N_22471,N_21668);
xor U23983 (N_23983,N_21096,N_21000);
nor U23984 (N_23984,N_21329,N_21539);
xor U23985 (N_23985,N_22118,N_21624);
nor U23986 (N_23986,N_21519,N_21098);
and U23987 (N_23987,N_22127,N_21532);
nand U23988 (N_23988,N_21148,N_21794);
and U23989 (N_23989,N_22177,N_22063);
and U23990 (N_23990,N_21354,N_22102);
and U23991 (N_23991,N_22352,N_22041);
nor U23992 (N_23992,N_21361,N_21874);
nor U23993 (N_23993,N_21263,N_21623);
xnor U23994 (N_23994,N_21147,N_21213);
nand U23995 (N_23995,N_21581,N_22006);
and U23996 (N_23996,N_22106,N_21420);
nor U23997 (N_23997,N_21621,N_21753);
xor U23998 (N_23998,N_21632,N_21199);
or U23999 (N_23999,N_21084,N_21237);
xor U24000 (N_24000,N_23093,N_23678);
nor U24001 (N_24001,N_23484,N_23392);
xor U24002 (N_24002,N_23574,N_23178);
nor U24003 (N_24003,N_23265,N_23009);
and U24004 (N_24004,N_23291,N_23783);
nand U24005 (N_24005,N_23903,N_23726);
xor U24006 (N_24006,N_22653,N_22737);
nor U24007 (N_24007,N_23494,N_23233);
nor U24008 (N_24008,N_23363,N_22953);
xor U24009 (N_24009,N_23218,N_23064);
xor U24010 (N_24010,N_23303,N_22860);
nor U24011 (N_24011,N_23342,N_23148);
xor U24012 (N_24012,N_22764,N_23229);
and U24013 (N_24013,N_23880,N_23956);
nand U24014 (N_24014,N_23656,N_23564);
nor U24015 (N_24015,N_23677,N_23247);
or U24016 (N_24016,N_23873,N_22888);
nand U24017 (N_24017,N_23081,N_23769);
nand U24018 (N_24018,N_22950,N_22952);
or U24019 (N_24019,N_23384,N_23642);
nor U24020 (N_24020,N_23274,N_23219);
nor U24021 (N_24021,N_23414,N_22602);
and U24022 (N_24022,N_22813,N_23216);
nor U24023 (N_24023,N_23536,N_23876);
nor U24024 (N_24024,N_23991,N_22980);
nor U24025 (N_24025,N_23804,N_23917);
and U24026 (N_24026,N_22578,N_23046);
or U24027 (N_24027,N_22740,N_23482);
or U24028 (N_24028,N_23417,N_22900);
and U24029 (N_24029,N_23153,N_23039);
or U24030 (N_24030,N_22798,N_22611);
or U24031 (N_24031,N_23278,N_23849);
and U24032 (N_24032,N_23404,N_22969);
nand U24033 (N_24033,N_23251,N_22864);
xor U24034 (N_24034,N_23751,N_23753);
and U24035 (N_24035,N_23271,N_22658);
nand U24036 (N_24036,N_22549,N_23292);
and U24037 (N_24037,N_22748,N_23937);
or U24038 (N_24038,N_23572,N_23275);
nor U24039 (N_24039,N_23738,N_23760);
nand U24040 (N_24040,N_23322,N_22509);
nor U24041 (N_24041,N_22745,N_23792);
nor U24042 (N_24042,N_23790,N_23050);
xnor U24043 (N_24043,N_23280,N_22782);
nor U24044 (N_24044,N_23776,N_23314);
xor U24045 (N_24045,N_23149,N_22598);
or U24046 (N_24046,N_23629,N_22552);
or U24047 (N_24047,N_23735,N_22609);
nor U24048 (N_24048,N_23758,N_23300);
nand U24049 (N_24049,N_23706,N_22743);
or U24050 (N_24050,N_22837,N_22755);
xnor U24051 (N_24051,N_23528,N_23584);
xor U24052 (N_24052,N_23550,N_23302);
and U24053 (N_24053,N_22779,N_22838);
or U24054 (N_24054,N_23512,N_23750);
xnor U24055 (N_24055,N_22536,N_23413);
xor U24056 (N_24056,N_23939,N_23968);
or U24057 (N_24057,N_23320,N_22587);
or U24058 (N_24058,N_23775,N_23490);
xor U24059 (N_24059,N_23555,N_23946);
nand U24060 (N_24060,N_23955,N_23854);
xnor U24061 (N_24061,N_22507,N_23231);
nand U24062 (N_24062,N_22982,N_23513);
and U24063 (N_24063,N_23266,N_22688);
and U24064 (N_24064,N_22849,N_23539);
and U24065 (N_24065,N_22651,N_22822);
xnor U24066 (N_24066,N_23076,N_23906);
and U24067 (N_24067,N_23249,N_22833);
nor U24068 (N_24068,N_23205,N_22853);
or U24069 (N_24069,N_23382,N_23984);
nor U24070 (N_24070,N_22520,N_23640);
and U24071 (N_24071,N_22992,N_23372);
and U24072 (N_24072,N_23001,N_23655);
nor U24073 (N_24073,N_22948,N_23426);
or U24074 (N_24074,N_22866,N_22919);
xnor U24075 (N_24075,N_22912,N_23026);
xor U24076 (N_24076,N_22519,N_23552);
or U24077 (N_24077,N_23455,N_23394);
nor U24078 (N_24078,N_23763,N_22895);
and U24079 (N_24079,N_23732,N_22683);
xor U24080 (N_24080,N_23713,N_23893);
nand U24081 (N_24081,N_23331,N_22872);
or U24082 (N_24082,N_23590,N_23953);
nand U24083 (N_24083,N_23554,N_22918);
and U24084 (N_24084,N_23096,N_23252);
nand U24085 (N_24085,N_23988,N_23442);
nand U24086 (N_24086,N_23246,N_23355);
or U24087 (N_24087,N_23890,N_23003);
nor U24088 (N_24088,N_23774,N_23729);
nor U24089 (N_24089,N_23131,N_22867);
nor U24090 (N_24090,N_23930,N_22840);
nor U24091 (N_24091,N_23217,N_23618);
nand U24092 (N_24092,N_23406,N_23118);
or U24093 (N_24093,N_23616,N_23015);
and U24094 (N_24094,N_22733,N_22712);
nor U24095 (N_24095,N_22882,N_23747);
nand U24096 (N_24096,N_23110,N_23522);
nor U24097 (N_24097,N_23307,N_23987);
or U24098 (N_24098,N_22809,N_23435);
xnor U24099 (N_24099,N_23826,N_22890);
xor U24100 (N_24100,N_22599,N_23960);
nor U24101 (N_24101,N_22789,N_23861);
and U24102 (N_24102,N_23884,N_23023);
xor U24103 (N_24103,N_23922,N_23209);
xor U24104 (N_24104,N_23843,N_22704);
or U24105 (N_24105,N_23200,N_22633);
and U24106 (N_24106,N_23881,N_23220);
nor U24107 (N_24107,N_23874,N_23600);
nor U24108 (N_24108,N_23126,N_23888);
and U24109 (N_24109,N_23586,N_23851);
or U24110 (N_24110,N_23082,N_22988);
nor U24111 (N_24111,N_22739,N_22576);
nand U24112 (N_24112,N_22521,N_23299);
and U24113 (N_24113,N_23672,N_23581);
and U24114 (N_24114,N_22725,N_23440);
xor U24115 (N_24115,N_23635,N_23954);
or U24116 (N_24116,N_22843,N_22985);
nor U24117 (N_24117,N_22772,N_23092);
and U24118 (N_24118,N_23033,N_22635);
and U24119 (N_24119,N_23277,N_22696);
xnor U24120 (N_24120,N_23059,N_22591);
xnor U24121 (N_24121,N_22652,N_22506);
xor U24122 (N_24122,N_22999,N_23571);
and U24123 (N_24123,N_23370,N_23828);
nand U24124 (N_24124,N_23969,N_23168);
nand U24125 (N_24125,N_23256,N_23237);
nor U24126 (N_24126,N_23373,N_22553);
xor U24127 (N_24127,N_23981,N_22944);
and U24128 (N_24128,N_23661,N_23514);
and U24129 (N_24129,N_23736,N_23643);
and U24130 (N_24130,N_23193,N_23585);
nor U24131 (N_24131,N_23324,N_23815);
nor U24132 (N_24132,N_23145,N_22628);
xnor U24133 (N_24133,N_23894,N_22703);
and U24134 (N_24134,N_23791,N_23399);
xnor U24135 (N_24135,N_22596,N_23974);
and U24136 (N_24136,N_22650,N_23798);
nor U24137 (N_24137,N_22961,N_23390);
or U24138 (N_24138,N_23936,N_23768);
and U24139 (N_24139,N_23606,N_23337);
or U24140 (N_24140,N_22746,N_23461);
or U24141 (N_24141,N_23632,N_23142);
or U24142 (N_24142,N_23408,N_23745);
nand U24143 (N_24143,N_22959,N_22619);
or U24144 (N_24144,N_23971,N_23340);
or U24145 (N_24145,N_23478,N_23577);
nor U24146 (N_24146,N_23483,N_23028);
or U24147 (N_24147,N_23623,N_23685);
or U24148 (N_24148,N_23005,N_23973);
nor U24149 (N_24149,N_22573,N_23961);
nor U24150 (N_24150,N_22994,N_23281);
and U24151 (N_24151,N_23610,N_23002);
or U24152 (N_24152,N_23613,N_22754);
xor U24153 (N_24153,N_23665,N_22510);
or U24154 (N_24154,N_22937,N_23710);
and U24155 (N_24155,N_23128,N_23607);
nor U24156 (N_24156,N_22747,N_22684);
xnor U24157 (N_24157,N_22511,N_23883);
or U24158 (N_24158,N_22861,N_23821);
or U24159 (N_24159,N_23165,N_22542);
nand U24160 (N_24160,N_23914,N_23493);
nor U24161 (N_24161,N_23038,N_23248);
or U24162 (N_24162,N_23063,N_22829);
nand U24163 (N_24163,N_23687,N_23173);
xor U24164 (N_24164,N_22645,N_23502);
nor U24165 (N_24165,N_23369,N_23171);
xnor U24166 (N_24166,N_22807,N_23925);
or U24167 (N_24167,N_23657,N_23544);
nor U24168 (N_24168,N_22610,N_22667);
or U24169 (N_24169,N_22532,N_22717);
xor U24170 (N_24170,N_23376,N_22824);
xnor U24171 (N_24171,N_23464,N_23226);
nand U24172 (N_24172,N_23362,N_22977);
nor U24173 (N_24173,N_23867,N_23232);
nand U24174 (N_24174,N_23570,N_22987);
and U24175 (N_24175,N_23445,N_22927);
or U24176 (N_24176,N_22941,N_23976);
xnor U24177 (N_24177,N_23159,N_23746);
or U24178 (N_24178,N_23839,N_23140);
nand U24179 (N_24179,N_22791,N_23651);
xor U24180 (N_24180,N_22891,N_22559);
or U24181 (N_24181,N_22991,N_22657);
nand U24182 (N_24182,N_23712,N_22761);
and U24183 (N_24183,N_23460,N_23386);
nor U24184 (N_24184,N_23127,N_23272);
nor U24185 (N_24185,N_22711,N_22535);
and U24186 (N_24186,N_23000,N_22562);
nand U24187 (N_24187,N_23022,N_23598);
nand U24188 (N_24188,N_22801,N_23080);
nor U24189 (N_24189,N_23594,N_22525);
xnor U24190 (N_24190,N_22719,N_23345);
nand U24191 (N_24191,N_23517,N_23695);
xnor U24192 (N_24192,N_22936,N_23488);
or U24193 (N_24193,N_22753,N_23479);
and U24194 (N_24194,N_23509,N_23170);
or U24195 (N_24195,N_22975,N_23176);
nand U24196 (N_24196,N_23359,N_23859);
xnor U24197 (N_24197,N_23680,N_22620);
nor U24198 (N_24198,N_22797,N_23241);
or U24199 (N_24199,N_22616,N_22640);
nor U24200 (N_24200,N_22502,N_22736);
xor U24201 (N_24201,N_23820,N_23945);
nor U24202 (N_24202,N_22855,N_23866);
xor U24203 (N_24203,N_23562,N_23078);
and U24204 (N_24204,N_23761,N_23367);
and U24205 (N_24205,N_23349,N_23208);
nand U24206 (N_24206,N_23994,N_23803);
and U24207 (N_24207,N_23895,N_22656);
nor U24208 (N_24208,N_22503,N_23019);
nand U24209 (N_24209,N_23767,N_23662);
xnor U24210 (N_24210,N_23926,N_23430);
nor U24211 (N_24211,N_23700,N_23155);
xor U24212 (N_24212,N_23389,N_22716);
nand U24213 (N_24213,N_23630,N_23177);
nand U24214 (N_24214,N_22618,N_22685);
and U24215 (N_24215,N_23371,N_22911);
xor U24216 (N_24216,N_23343,N_23701);
xor U24217 (N_24217,N_22744,N_23161);
and U24218 (N_24218,N_23912,N_23567);
xnor U24219 (N_24219,N_23497,N_23759);
nand U24220 (N_24220,N_22899,N_22751);
xor U24221 (N_24221,N_22957,N_23978);
or U24222 (N_24222,N_22925,N_23403);
nand U24223 (N_24223,N_22665,N_22672);
and U24224 (N_24224,N_23213,N_23310);
and U24225 (N_24225,N_22921,N_23591);
nor U24226 (N_24226,N_22881,N_23141);
or U24227 (N_24227,N_22714,N_22540);
or U24228 (N_24228,N_23206,N_23966);
or U24229 (N_24229,N_23682,N_23838);
nor U24230 (N_24230,N_23915,N_23174);
or U24231 (N_24231,N_23805,N_23060);
nand U24232 (N_24232,N_23857,N_23287);
nand U24233 (N_24233,N_23456,N_22713);
or U24234 (N_24234,N_23366,N_23401);
nor U24235 (N_24235,N_23416,N_23947);
or U24236 (N_24236,N_22623,N_23733);
xor U24237 (N_24237,N_23877,N_23381);
or U24238 (N_24238,N_23061,N_22907);
or U24239 (N_24239,N_22956,N_23253);
or U24240 (N_24240,N_23869,N_23789);
or U24241 (N_24241,N_23566,N_23079);
xor U24242 (N_24242,N_23834,N_23535);
xor U24243 (N_24243,N_23719,N_23801);
or U24244 (N_24244,N_23734,N_23311);
nor U24245 (N_24245,N_22947,N_23197);
or U24246 (N_24246,N_23658,N_23533);
nand U24247 (N_24247,N_23344,N_23722);
nand U24248 (N_24248,N_23108,N_23853);
nand U24249 (N_24249,N_23457,N_23244);
xnor U24250 (N_24250,N_22997,N_23419);
nand U24251 (N_24251,N_22889,N_23199);
nand U24252 (N_24252,N_22637,N_23167);
or U24253 (N_24253,N_23405,N_23336);
nor U24254 (N_24254,N_23365,N_22790);
xnor U24255 (N_24255,N_23619,N_22673);
nor U24256 (N_24256,N_23011,N_23236);
nand U24257 (N_24257,N_23186,N_23264);
and U24258 (N_24258,N_23516,N_23179);
or U24259 (N_24259,N_23998,N_22817);
and U24260 (N_24260,N_22862,N_23025);
and U24261 (N_24261,N_23480,N_23031);
nand U24262 (N_24262,N_22655,N_23016);
or U24263 (N_24263,N_23103,N_23901);
or U24264 (N_24264,N_23222,N_23811);
nand U24265 (N_24265,N_23130,N_22729);
nand U24266 (N_24266,N_23358,N_22939);
nand U24267 (N_24267,N_23162,N_23556);
and U24268 (N_24268,N_23975,N_23073);
and U24269 (N_24269,N_23921,N_23465);
nor U24270 (N_24270,N_23447,N_22583);
or U24271 (N_24271,N_23716,N_23786);
or U24272 (N_24272,N_23150,N_22970);
or U24273 (N_24273,N_23296,N_23989);
xnor U24274 (N_24274,N_22776,N_22989);
nor U24275 (N_24275,N_22680,N_23286);
nor U24276 (N_24276,N_22949,N_23636);
or U24277 (N_24277,N_22728,N_23752);
or U24278 (N_24278,N_23737,N_23660);
nor U24279 (N_24279,N_22879,N_23526);
xnor U24280 (N_24280,N_23052,N_22581);
nor U24281 (N_24281,N_23900,N_23357);
xnor U24282 (N_24282,N_23184,N_23950);
nand U24283 (N_24283,N_23066,N_23327);
and U24284 (N_24284,N_22516,N_22590);
xnor U24285 (N_24285,N_23317,N_23474);
xnor U24286 (N_24286,N_23608,N_23891);
nor U24287 (N_24287,N_22920,N_23850);
and U24288 (N_24288,N_23538,N_23087);
nand U24289 (N_24289,N_23439,N_23330);
nand U24290 (N_24290,N_23102,N_23885);
and U24291 (N_24291,N_23121,N_22625);
nand U24292 (N_24292,N_23112,N_23182);
nand U24293 (N_24293,N_23611,N_23565);
nor U24294 (N_24294,N_22870,N_23048);
nand U24295 (N_24295,N_22905,N_22694);
xor U24296 (N_24296,N_22508,N_23652);
nor U24297 (N_24297,N_22821,N_22836);
or U24298 (N_24298,N_23263,N_23492);
and U24299 (N_24299,N_23505,N_23578);
nor U24300 (N_24300,N_22705,N_23720);
and U24301 (N_24301,N_23012,N_23152);
or U24302 (N_24302,N_23541,N_22768);
or U24303 (N_24303,N_22514,N_23638);
xor U24304 (N_24304,N_23757,N_22677);
and U24305 (N_24305,N_23443,N_23032);
xnor U24306 (N_24306,N_23452,N_23659);
nor U24307 (N_24307,N_22819,N_22990);
and U24308 (N_24308,N_23728,N_23215);
xor U24309 (N_24309,N_23529,N_22631);
xnor U24310 (N_24310,N_22643,N_23388);
nor U24311 (N_24311,N_23739,N_23273);
or U24312 (N_24312,N_22641,N_23049);
and U24313 (N_24313,N_23020,N_23856);
and U24314 (N_24314,N_22526,N_23181);
and U24315 (N_24315,N_23870,N_23137);
nor U24316 (N_24316,N_23228,N_23276);
nor U24317 (N_24317,N_23312,N_22720);
nor U24318 (N_24318,N_22723,N_23605);
or U24319 (N_24319,N_23602,N_23519);
nand U24320 (N_24320,N_22923,N_22878);
xnor U24321 (N_24321,N_23353,N_23230);
and U24322 (N_24322,N_23862,N_22766);
and U24323 (N_24323,N_22595,N_23294);
nand U24324 (N_24324,N_22831,N_23288);
and U24325 (N_24325,N_23428,N_22557);
xor U24326 (N_24326,N_22886,N_22597);
nand U24327 (N_24327,N_22897,N_22960);
xor U24328 (N_24328,N_23972,N_22593);
or U24329 (N_24329,N_22851,N_23592);
nor U24330 (N_24330,N_23772,N_23617);
and U24331 (N_24331,N_22916,N_22796);
and U24332 (N_24332,N_23647,N_22710);
or U24333 (N_24333,N_23597,N_23301);
or U24334 (N_24334,N_23313,N_22555);
or U24335 (N_24335,N_23727,N_22522);
nand U24336 (N_24336,N_22757,N_23547);
xor U24337 (N_24337,N_22504,N_23117);
or U24338 (N_24338,N_22606,N_22906);
nor U24339 (N_24339,N_22852,N_23583);
nor U24340 (N_24340,N_23653,N_23697);
xor U24341 (N_24341,N_22662,N_23085);
and U24342 (N_24342,N_22681,N_23691);
and U24343 (N_24343,N_23589,N_22527);
and U24344 (N_24344,N_22523,N_23559);
nor U24345 (N_24345,N_23245,N_23214);
nand U24346 (N_24346,N_23420,N_23227);
or U24347 (N_24347,N_22505,N_23596);
nand U24348 (N_24348,N_23510,N_22675);
nand U24349 (N_24349,N_23021,N_23558);
nand U24350 (N_24350,N_22876,N_23957);
or U24351 (N_24351,N_22933,N_22995);
nand U24352 (N_24352,N_23160,N_23268);
and U24353 (N_24353,N_23711,N_23051);
and U24354 (N_24354,N_23633,N_23243);
nor U24355 (N_24355,N_22571,N_23489);
xnor U24356 (N_24356,N_23469,N_22986);
or U24357 (N_24357,N_22938,N_22500);
and U24358 (N_24358,N_23094,N_22541);
xor U24359 (N_24359,N_23542,N_23621);
and U24360 (N_24360,N_23681,N_23886);
xor U24361 (N_24361,N_23819,N_22967);
xnor U24362 (N_24362,N_22560,N_23400);
nor U24363 (N_24363,N_23267,N_22934);
nor U24364 (N_24364,N_22741,N_23506);
xor U24365 (N_24365,N_23283,N_22946);
or U24366 (N_24366,N_22605,N_23315);
or U24367 (N_24367,N_22615,N_23380);
xor U24368 (N_24368,N_23409,N_23996);
xnor U24369 (N_24369,N_23030,N_23507);
nor U24370 (N_24370,N_23847,N_22586);
or U24371 (N_24371,N_22730,N_22786);
and U24372 (N_24372,N_22913,N_23799);
nand U24373 (N_24373,N_23361,N_23604);
xor U24374 (N_24374,N_23860,N_23848);
xor U24375 (N_24375,N_22617,N_23599);
xor U24376 (N_24376,N_22760,N_22648);
nand U24377 (N_24377,N_23441,N_22577);
or U24378 (N_24378,N_22850,N_23568);
nor U24379 (N_24379,N_23034,N_23224);
xor U24380 (N_24380,N_22915,N_22904);
or U24381 (N_24381,N_23007,N_23808);
xnor U24382 (N_24382,N_22835,N_23622);
nand U24383 (N_24383,N_22847,N_23354);
and U24384 (N_24384,N_23203,N_23962);
nand U24385 (N_24385,N_22756,N_22863);
nor U24386 (N_24386,N_22763,N_23433);
or U24387 (N_24387,N_23645,N_22945);
and U24388 (N_24388,N_23959,N_23113);
nand U24389 (N_24389,N_23690,N_23451);
xnor U24390 (N_24390,N_23837,N_23825);
xnor U24391 (N_24391,N_23298,N_23496);
and U24392 (N_24392,N_23062,N_23100);
and U24393 (N_24393,N_22556,N_23074);
xnor U24394 (N_24394,N_22626,N_22629);
or U24395 (N_24395,N_22530,N_23135);
and U24396 (N_24396,N_23724,N_23472);
nor U24397 (N_24397,N_23258,N_22784);
or U24398 (N_24398,N_23899,N_22812);
and U24399 (N_24399,N_22512,N_23043);
nor U24400 (N_24400,N_22932,N_23679);
or U24401 (N_24401,N_23693,N_22529);
and U24402 (N_24402,N_23255,N_23377);
xor U24403 (N_24403,N_22575,N_22706);
and U24404 (N_24404,N_23316,N_22515);
nand U24405 (N_24405,N_23067,N_23902);
nor U24406 (N_24406,N_22826,N_22668);
nor U24407 (N_24407,N_23694,N_23931);
nand U24408 (N_24408,N_22868,N_23393);
nand U24409 (N_24409,N_23004,N_23044);
nand U24410 (N_24410,N_22978,N_23540);
or U24411 (N_24411,N_23924,N_22844);
nor U24412 (N_24412,N_23582,N_23527);
nor U24413 (N_24413,N_22752,N_22901);
nand U24414 (N_24414,N_23055,N_22554);
and U24415 (N_24415,N_22972,N_22954);
nand U24416 (N_24416,N_23449,N_23065);
nand U24417 (N_24417,N_22674,N_23421);
or U24418 (N_24418,N_23637,N_23948);
and U24419 (N_24419,N_23250,N_23018);
nand U24420 (N_24420,N_22871,N_22699);
nand U24421 (N_24421,N_23010,N_23411);
and U24422 (N_24422,N_23634,N_23169);
nor U24423 (N_24423,N_23183,N_22942);
or U24424 (N_24424,N_22926,N_22660);
and U24425 (N_24425,N_23158,N_22811);
and U24426 (N_24426,N_23129,N_23800);
xor U24427 (N_24427,N_23503,N_22765);
xor U24428 (N_24428,N_22546,N_23762);
or U24429 (N_24429,N_23949,N_23784);
and U24430 (N_24430,N_22827,N_23919);
xnor U24431 (N_24431,N_23952,N_22604);
and U24432 (N_24432,N_23305,N_22517);
and U24433 (N_24433,N_22544,N_23699);
nor U24434 (N_24434,N_23983,N_22708);
and U24435 (N_24435,N_23667,N_22770);
xnor U24436 (N_24436,N_23744,N_23190);
nor U24437 (N_24437,N_23887,N_23463);
xnor U24438 (N_24438,N_22721,N_23101);
and U24439 (N_24439,N_23708,N_23940);
or U24440 (N_24440,N_22898,N_23832);
xor U24441 (N_24441,N_22803,N_23098);
xor U24442 (N_24442,N_23603,N_23646);
nand U24443 (N_24443,N_23625,N_23398);
or U24444 (N_24444,N_23057,N_23326);
nor U24445 (N_24445,N_23898,N_23951);
and U24446 (N_24446,N_23378,N_23929);
and U24447 (N_24447,N_22533,N_23418);
or U24448 (N_24448,N_23201,N_22695);
and U24449 (N_24449,N_22848,N_23928);
and U24450 (N_24450,N_23341,N_23508);
nand U24451 (N_24451,N_22767,N_23427);
xor U24452 (N_24452,N_22964,N_23918);
xor U24453 (N_24453,N_22592,N_23965);
nand U24454 (N_24454,N_22566,N_23813);
and U24455 (N_24455,N_23620,N_23262);
xor U24456 (N_24456,N_23530,N_22996);
or U24457 (N_24457,N_22788,N_23029);
xnor U24458 (N_24458,N_22909,N_22682);
nand U24459 (N_24459,N_23933,N_23992);
and U24460 (N_24460,N_22664,N_23095);
xor U24461 (N_24461,N_23717,N_23072);
nor U24462 (N_24462,N_23569,N_23683);
xnor U24463 (N_24463,N_23334,N_23714);
or U24464 (N_24464,N_22731,N_22630);
xor U24465 (N_24465,N_22981,N_23054);
and U24466 (N_24466,N_23068,N_23882);
or U24467 (N_24467,N_22893,N_23781);
xnor U24468 (N_24468,N_23202,N_23718);
nand U24469 (N_24469,N_22601,N_23730);
and U24470 (N_24470,N_22671,N_22669);
or U24471 (N_24471,N_23725,N_22734);
nand U24472 (N_24472,N_23911,N_23125);
or U24473 (N_24473,N_23641,N_23122);
and U24474 (N_24474,N_23935,N_23561);
nor U24475 (N_24475,N_23089,N_23916);
xor U24476 (N_24476,N_22914,N_22579);
nand U24477 (N_24477,N_23075,N_22883);
or U24478 (N_24478,N_23740,N_23560);
xnor U24479 (N_24479,N_23579,N_23835);
nor U24480 (N_24480,N_23765,N_22565);
nand U24481 (N_24481,N_23785,N_23257);
or U24482 (N_24482,N_23858,N_22841);
xor U24483 (N_24483,N_23576,N_22715);
and U24484 (N_24484,N_23537,N_22903);
nand U24485 (N_24485,N_23115,N_22608);
xor U24486 (N_24486,N_23006,N_23356);
xnor U24487 (N_24487,N_23360,N_23396);
or U24488 (N_24488,N_22687,N_23553);
and U24489 (N_24489,N_22974,N_22777);
nor U24490 (N_24490,N_23139,N_23454);
or U24491 (N_24491,N_23521,N_23491);
nor U24492 (N_24492,N_22732,N_22922);
nor U24493 (N_24493,N_23580,N_22572);
xor U24494 (N_24494,N_23612,N_23383);
or U24495 (N_24495,N_22924,N_23707);
nor U24496 (N_24496,N_23523,N_22642);
or U24497 (N_24497,N_22561,N_23818);
and U24498 (N_24498,N_23980,N_23212);
nor U24499 (N_24499,N_23352,N_23017);
nor U24500 (N_24500,N_22799,N_23339);
nor U24501 (N_24501,N_23543,N_22892);
xnor U24502 (N_24502,N_22644,N_22589);
nand U24503 (N_24503,N_22958,N_23846);
nor U24504 (N_24504,N_23164,N_22830);
and U24505 (N_24505,N_23979,N_23470);
or U24506 (N_24506,N_23705,N_23993);
nand U24507 (N_24507,N_22774,N_23709);
nor U24508 (N_24508,N_22569,N_23041);
nor U24509 (N_24509,N_23412,N_23351);
xnor U24510 (N_24510,N_23013,N_22820);
or U24511 (N_24511,N_23787,N_23995);
and U24512 (N_24512,N_22955,N_23696);
nor U24513 (N_24513,N_22528,N_23563);
nand U24514 (N_24514,N_23982,N_23627);
or U24515 (N_24515,N_23986,N_23824);
or U24516 (N_24516,N_23347,N_23788);
and U24517 (N_24517,N_22676,N_23686);
xnor U24518 (N_24518,N_23504,N_23648);
xor U24519 (N_24519,N_23368,N_23335);
or U24520 (N_24520,N_23323,N_23188);
xor U24521 (N_24521,N_23180,N_23692);
nor U24522 (N_24522,N_23297,N_22659);
or U24523 (N_24523,N_22828,N_22607);
and U24524 (N_24524,N_22877,N_23036);
or U24525 (N_24525,N_23448,N_23106);
xor U24526 (N_24526,N_22563,N_22929);
or U24527 (N_24527,N_23109,N_23084);
xnor U24528 (N_24528,N_22908,N_22513);
and U24529 (N_24529,N_23844,N_22804);
xor U24530 (N_24530,N_23822,N_23779);
nor U24531 (N_24531,N_23318,N_23045);
and U24532 (N_24532,N_23284,N_22759);
or U24533 (N_24533,N_22951,N_23166);
nand U24534 (N_24534,N_23666,N_22588);
nand U24535 (N_24535,N_23107,N_23144);
xnor U24536 (N_24536,N_23743,N_23407);
nand U24537 (N_24537,N_23486,N_23810);
or U24538 (N_24538,N_22670,N_23111);
or U24539 (N_24539,N_23557,N_22697);
nor U24540 (N_24540,N_23802,N_22795);
xor U24541 (N_24541,N_23628,N_23796);
and U24542 (N_24542,N_23402,N_22518);
or U24543 (N_24543,N_23069,N_22701);
nor U24544 (N_24544,N_23120,N_23154);
and U24545 (N_24545,N_23868,N_22794);
and U24546 (N_24546,N_22781,N_23053);
nand U24547 (N_24547,N_22808,N_23097);
or U24548 (N_24548,N_22910,N_22663);
nand U24549 (N_24549,N_23423,N_23575);
or U24550 (N_24550,N_23524,N_23468);
and U24551 (N_24551,N_22622,N_23487);
nor U24552 (N_24552,N_23999,N_23254);
and U24553 (N_24553,N_22691,N_23501);
nand U24554 (N_24554,N_23688,N_23615);
and U24555 (N_24555,N_23221,N_23040);
nor U24556 (N_24556,N_23119,N_22501);
and U24557 (N_24557,N_23192,N_23374);
nand U24558 (N_24558,N_23664,N_22649);
nor U24559 (N_24559,N_22698,N_23941);
or U24560 (N_24560,N_23511,N_23143);
xnor U24561 (N_24561,N_23211,N_23814);
nand U24562 (N_24562,N_22634,N_23782);
and U24563 (N_24563,N_23654,N_23410);
nor U24564 (N_24564,N_22928,N_22896);
and U24565 (N_24565,N_22543,N_23806);
nand U24566 (N_24566,N_23269,N_23147);
nand U24567 (N_24567,N_22858,N_22550);
xor U24568 (N_24568,N_23963,N_23133);
and U24569 (N_24569,N_23609,N_23749);
xnor U24570 (N_24570,N_22582,N_23104);
or U24571 (N_24571,N_23473,N_23855);
and U24572 (N_24572,N_22873,N_23715);
and U24573 (N_24573,N_22638,N_23905);
nand U24574 (N_24574,N_23771,N_23191);
or U24575 (N_24575,N_22880,N_23518);
nand U24576 (N_24576,N_23573,N_23748);
xnor U24577 (N_24577,N_22545,N_22859);
xor U24578 (N_24578,N_23650,N_23425);
nor U24579 (N_24579,N_22832,N_23778);
nor U24580 (N_24580,N_23481,N_23833);
xnor U24581 (N_24581,N_23721,N_23499);
or U24582 (N_24582,N_22846,N_23437);
and U24583 (N_24583,N_23467,N_23293);
nand U24584 (N_24584,N_23593,N_22930);
nand U24585 (N_24585,N_23136,N_22823);
nor U24586 (N_24586,N_23172,N_23397);
xnor U24587 (N_24587,N_23889,N_23764);
and U24588 (N_24588,N_23500,N_22749);
xnor U24589 (N_24589,N_23282,N_23459);
nor U24590 (N_24590,N_23932,N_22702);
xor U24591 (N_24591,N_23270,N_23534);
and U24592 (N_24592,N_23138,N_23114);
and U24593 (N_24593,N_23964,N_23704);
nor U24594 (N_24594,N_23967,N_23875);
nand U24595 (N_24595,N_22940,N_23827);
and U24596 (N_24596,N_22816,N_23907);
nand U24597 (N_24597,N_23896,N_23829);
nor U24598 (N_24598,N_23466,N_23871);
nand U24599 (N_24599,N_23840,N_23495);
or U24600 (N_24600,N_22773,N_22869);
nor U24601 (N_24601,N_22722,N_23083);
xnor U24602 (N_24602,N_23675,N_23328);
nand U24603 (N_24603,N_23189,N_22584);
nand U24604 (N_24604,N_22887,N_22718);
xor U24605 (N_24605,N_22935,N_23458);
nor U24606 (N_24606,N_23639,N_23385);
nand U24607 (N_24607,N_23239,N_23422);
and U24608 (N_24608,N_23146,N_22742);
and U24609 (N_24609,N_23196,N_23731);
nor U24610 (N_24610,N_23741,N_23549);
nand U24611 (N_24611,N_23942,N_23123);
xnor U24612 (N_24612,N_22537,N_23207);
and U24613 (N_24613,N_23151,N_22614);
or U24614 (N_24614,N_23424,N_22647);
xnor U24615 (N_24615,N_22971,N_22724);
xor U24616 (N_24616,N_23668,N_22594);
nor U24617 (N_24617,N_22547,N_22931);
xnor U24618 (N_24618,N_23515,N_23124);
xor U24619 (N_24619,N_23669,N_23295);
or U24620 (N_24620,N_22839,N_22800);
xor U24621 (N_24621,N_23684,N_23644);
xor U24622 (N_24622,N_23649,N_22585);
nand U24623 (N_24623,N_23024,N_23807);
nor U24624 (N_24624,N_22806,N_22738);
or U24625 (N_24625,N_23531,N_23329);
nor U24626 (N_24626,N_23702,N_22689);
nor U24627 (N_24627,N_22885,N_22621);
and U24628 (N_24628,N_23210,N_22707);
xnor U24629 (N_24629,N_23485,N_22979);
or U24630 (N_24630,N_22787,N_22857);
and U24631 (N_24631,N_22639,N_22679);
nand U24632 (N_24632,N_23134,N_22654);
or U24633 (N_24633,N_22963,N_23816);
nor U24634 (N_24634,N_23309,N_22775);
xor U24635 (N_24635,N_23864,N_23498);
or U24636 (N_24636,N_22865,N_23525);
xor U24637 (N_24637,N_22666,N_22998);
or U24638 (N_24638,N_23204,N_23676);
nand U24639 (N_24639,N_22570,N_23588);
or U24640 (N_24640,N_22558,N_22785);
or U24641 (N_24641,N_23977,N_23185);
nand U24642 (N_24642,N_23070,N_22845);
and U24643 (N_24643,N_22943,N_22531);
nand U24644 (N_24644,N_23823,N_23350);
xor U24645 (N_24645,N_23432,N_22750);
xor U24646 (N_24646,N_23689,N_23766);
nand U24647 (N_24647,N_23897,N_22693);
xnor U24648 (N_24648,N_22983,N_23794);
and U24649 (N_24649,N_22966,N_23471);
nand U24650 (N_24650,N_23830,N_23187);
nand U24651 (N_24651,N_23663,N_23934);
xnor U24652 (N_24652,N_23997,N_23546);
nand U24653 (N_24653,N_23944,N_23863);
nand U24654 (N_24654,N_23773,N_22538);
or U24655 (N_24655,N_23754,N_23809);
nor U24656 (N_24656,N_23304,N_23225);
or U24657 (N_24657,N_23091,N_23027);
and U24658 (N_24658,N_22539,N_22875);
or U24659 (N_24659,N_23595,N_23841);
or U24660 (N_24660,N_22917,N_22690);
and U24661 (N_24661,N_23259,N_23434);
and U24662 (N_24662,N_23436,N_23910);
nor U24663 (N_24663,N_22632,N_23090);
and U24664 (N_24664,N_23476,N_22700);
nor U24665 (N_24665,N_23943,N_23742);
or U24666 (N_24666,N_23852,N_23624);
nand U24667 (N_24667,N_22600,N_23391);
nor U24668 (N_24668,N_22962,N_22814);
or U24669 (N_24669,N_22802,N_23308);
nand U24670 (N_24670,N_23797,N_22965);
xnor U24671 (N_24671,N_23387,N_22856);
nor U24672 (N_24672,N_23938,N_23545);
or U24673 (N_24673,N_22574,N_23777);
and U24674 (N_24674,N_23836,N_23132);
nand U24675 (N_24675,N_23845,N_23240);
nor U24676 (N_24676,N_23035,N_22636);
and U24677 (N_24677,N_22976,N_22792);
or U24678 (N_24678,N_23077,N_23551);
or U24679 (N_24679,N_22692,N_23319);
nand U24680 (N_24680,N_23058,N_22854);
and U24681 (N_24681,N_23755,N_23375);
nor U24682 (N_24682,N_22993,N_23842);
and U24683 (N_24683,N_23614,N_23056);
nand U24684 (N_24684,N_23198,N_23631);
nand U24685 (N_24685,N_23175,N_22624);
or U24686 (N_24686,N_23446,N_23163);
nor U24687 (N_24687,N_23793,N_23223);
xor U24688 (N_24688,N_22524,N_22783);
xor U24689 (N_24689,N_22984,N_23306);
xor U24690 (N_24690,N_23333,N_23970);
and U24691 (N_24691,N_22834,N_22567);
nor U24692 (N_24692,N_23242,N_22735);
or U24693 (N_24693,N_23321,N_23332);
xnor U24694 (N_24694,N_22548,N_22613);
or U24695 (N_24695,N_23348,N_23453);
nor U24696 (N_24696,N_23042,N_23723);
and U24697 (N_24697,N_22874,N_23325);
xnor U24698 (N_24698,N_23812,N_23438);
nor U24699 (N_24699,N_23920,N_23099);
nand U24700 (N_24700,N_22534,N_23279);
nand U24701 (N_24701,N_22769,N_23157);
and U24702 (N_24702,N_23756,N_22661);
or U24703 (N_24703,N_23260,N_23195);
or U24704 (N_24704,N_23008,N_22726);
or U24705 (N_24705,N_22842,N_23674);
xnor U24706 (N_24706,N_23338,N_23985);
nand U24707 (N_24707,N_22580,N_23395);
nor U24708 (N_24708,N_23346,N_22780);
nor U24709 (N_24709,N_23892,N_22793);
or U24710 (N_24710,N_22894,N_22884);
or U24711 (N_24711,N_23770,N_23450);
nor U24712 (N_24712,N_23795,N_22771);
nor U24713 (N_24713,N_22603,N_23462);
and U24714 (N_24714,N_23532,N_23913);
and U24715 (N_24715,N_23234,N_23990);
xor U24716 (N_24716,N_23261,N_23444);
nand U24717 (N_24717,N_22551,N_23520);
xor U24718 (N_24718,N_23927,N_22646);
nor U24719 (N_24719,N_23958,N_23703);
nor U24720 (N_24720,N_23289,N_23878);
nor U24721 (N_24721,N_22727,N_23156);
nand U24722 (N_24722,N_23872,N_22810);
xor U24723 (N_24723,N_23477,N_23909);
or U24724 (N_24724,N_23626,N_23908);
or U24725 (N_24725,N_23673,N_23548);
nor U24726 (N_24726,N_23671,N_22825);
nor U24727 (N_24727,N_22686,N_23235);
and U24728 (N_24728,N_23698,N_23285);
xor U24729 (N_24729,N_23379,N_23879);
and U24730 (N_24730,N_23088,N_22778);
and U24731 (N_24731,N_23601,N_23105);
nand U24732 (N_24732,N_22968,N_23037);
and U24733 (N_24733,N_23587,N_23817);
xor U24734 (N_24734,N_23415,N_23014);
or U24735 (N_24735,N_22762,N_22902);
xnor U24736 (N_24736,N_23071,N_23194);
and U24737 (N_24737,N_23831,N_23780);
and U24738 (N_24738,N_23429,N_22709);
or U24739 (N_24739,N_23923,N_22805);
nor U24740 (N_24740,N_23238,N_23086);
or U24741 (N_24741,N_23047,N_22627);
xor U24742 (N_24742,N_23670,N_22758);
or U24743 (N_24743,N_22612,N_23290);
xnor U24744 (N_24744,N_23364,N_22568);
and U24745 (N_24745,N_22815,N_23904);
nor U24746 (N_24746,N_23431,N_22564);
or U24747 (N_24747,N_23865,N_23116);
xor U24748 (N_24748,N_22818,N_22973);
and U24749 (N_24749,N_23475,N_22678);
and U24750 (N_24750,N_22618,N_22815);
nor U24751 (N_24751,N_23060,N_23679);
or U24752 (N_24752,N_23104,N_23775);
nor U24753 (N_24753,N_23815,N_23572);
or U24754 (N_24754,N_22622,N_22822);
xor U24755 (N_24755,N_23360,N_22683);
xor U24756 (N_24756,N_23985,N_23483);
or U24757 (N_24757,N_23410,N_22722);
nor U24758 (N_24758,N_23928,N_22766);
or U24759 (N_24759,N_23580,N_23566);
and U24760 (N_24760,N_23084,N_22964);
nor U24761 (N_24761,N_22667,N_22536);
xor U24762 (N_24762,N_23877,N_23305);
nand U24763 (N_24763,N_22735,N_23607);
nor U24764 (N_24764,N_23763,N_23031);
nand U24765 (N_24765,N_22525,N_22775);
and U24766 (N_24766,N_23228,N_23034);
nand U24767 (N_24767,N_22701,N_23659);
or U24768 (N_24768,N_23929,N_23697);
and U24769 (N_24769,N_23042,N_23111);
and U24770 (N_24770,N_23725,N_23875);
nand U24771 (N_24771,N_22726,N_22782);
or U24772 (N_24772,N_23411,N_23353);
or U24773 (N_24773,N_23648,N_23622);
xnor U24774 (N_24774,N_23418,N_22930);
and U24775 (N_24775,N_23403,N_23999);
and U24776 (N_24776,N_23794,N_22623);
or U24777 (N_24777,N_23328,N_23059);
xnor U24778 (N_24778,N_23903,N_22617);
and U24779 (N_24779,N_22687,N_23556);
xnor U24780 (N_24780,N_23580,N_22762);
and U24781 (N_24781,N_23754,N_23235);
and U24782 (N_24782,N_23576,N_23883);
xnor U24783 (N_24783,N_23052,N_22927);
and U24784 (N_24784,N_22717,N_23618);
nand U24785 (N_24785,N_23485,N_23653);
xnor U24786 (N_24786,N_23996,N_23833);
nor U24787 (N_24787,N_22740,N_22811);
nand U24788 (N_24788,N_23383,N_22811);
or U24789 (N_24789,N_22975,N_23063);
nor U24790 (N_24790,N_23504,N_23543);
or U24791 (N_24791,N_22965,N_22756);
nor U24792 (N_24792,N_22560,N_23223);
nand U24793 (N_24793,N_22501,N_22699);
nor U24794 (N_24794,N_23392,N_22849);
or U24795 (N_24795,N_23676,N_22844);
xor U24796 (N_24796,N_23329,N_23261);
and U24797 (N_24797,N_23113,N_23365);
nand U24798 (N_24798,N_23933,N_22673);
nand U24799 (N_24799,N_23987,N_23895);
or U24800 (N_24800,N_23866,N_23265);
and U24801 (N_24801,N_23939,N_23801);
xnor U24802 (N_24802,N_22709,N_23949);
xor U24803 (N_24803,N_23009,N_23574);
nand U24804 (N_24804,N_22638,N_23074);
and U24805 (N_24805,N_23811,N_23480);
xnor U24806 (N_24806,N_23642,N_23651);
nor U24807 (N_24807,N_23322,N_23928);
nand U24808 (N_24808,N_22790,N_22502);
nand U24809 (N_24809,N_23130,N_23079);
xnor U24810 (N_24810,N_23604,N_23011);
nor U24811 (N_24811,N_23924,N_22772);
or U24812 (N_24812,N_23033,N_22815);
nor U24813 (N_24813,N_22508,N_23275);
nor U24814 (N_24814,N_22659,N_23053);
xor U24815 (N_24815,N_23119,N_23041);
or U24816 (N_24816,N_23192,N_23734);
and U24817 (N_24817,N_23472,N_23952);
or U24818 (N_24818,N_23357,N_23283);
and U24819 (N_24819,N_22959,N_22963);
or U24820 (N_24820,N_22807,N_22917);
xnor U24821 (N_24821,N_23026,N_23635);
nand U24822 (N_24822,N_23961,N_23910);
nor U24823 (N_24823,N_23762,N_23527);
nand U24824 (N_24824,N_23844,N_23909);
xor U24825 (N_24825,N_23583,N_22590);
and U24826 (N_24826,N_23119,N_23174);
xor U24827 (N_24827,N_23756,N_23896);
and U24828 (N_24828,N_23016,N_22923);
nand U24829 (N_24829,N_23823,N_22644);
and U24830 (N_24830,N_23591,N_22820);
nand U24831 (N_24831,N_22651,N_23642);
or U24832 (N_24832,N_23269,N_22527);
nand U24833 (N_24833,N_22522,N_23773);
nand U24834 (N_24834,N_22562,N_23661);
nand U24835 (N_24835,N_22717,N_23772);
nand U24836 (N_24836,N_22699,N_22695);
xnor U24837 (N_24837,N_23810,N_23140);
or U24838 (N_24838,N_22618,N_22609);
and U24839 (N_24839,N_23673,N_23353);
and U24840 (N_24840,N_23462,N_22668);
or U24841 (N_24841,N_23123,N_23440);
nand U24842 (N_24842,N_23472,N_23599);
and U24843 (N_24843,N_23525,N_22731);
or U24844 (N_24844,N_23702,N_23210);
and U24845 (N_24845,N_23934,N_23646);
nor U24846 (N_24846,N_23163,N_22686);
nand U24847 (N_24847,N_23392,N_23933);
or U24848 (N_24848,N_23597,N_22526);
xor U24849 (N_24849,N_22749,N_22645);
nor U24850 (N_24850,N_23006,N_22568);
or U24851 (N_24851,N_23284,N_23048);
and U24852 (N_24852,N_22966,N_23658);
nor U24853 (N_24853,N_23186,N_23348);
or U24854 (N_24854,N_23364,N_22610);
or U24855 (N_24855,N_22510,N_22787);
nor U24856 (N_24856,N_23637,N_23891);
and U24857 (N_24857,N_22824,N_23925);
or U24858 (N_24858,N_23386,N_23537);
or U24859 (N_24859,N_23698,N_23782);
or U24860 (N_24860,N_23192,N_22640);
nor U24861 (N_24861,N_22928,N_23039);
or U24862 (N_24862,N_23396,N_23615);
nor U24863 (N_24863,N_23164,N_22688);
and U24864 (N_24864,N_23063,N_23672);
nand U24865 (N_24865,N_23338,N_22828);
nand U24866 (N_24866,N_23646,N_23092);
xor U24867 (N_24867,N_23715,N_22593);
nor U24868 (N_24868,N_22924,N_22985);
or U24869 (N_24869,N_23625,N_23862);
and U24870 (N_24870,N_22607,N_23367);
nand U24871 (N_24871,N_22953,N_23705);
nand U24872 (N_24872,N_22618,N_22514);
nand U24873 (N_24873,N_23954,N_22806);
nor U24874 (N_24874,N_22923,N_23225);
and U24875 (N_24875,N_23747,N_23797);
xnor U24876 (N_24876,N_22703,N_22969);
nor U24877 (N_24877,N_23584,N_23237);
xnor U24878 (N_24878,N_22881,N_23841);
xor U24879 (N_24879,N_22551,N_22709);
nand U24880 (N_24880,N_22617,N_23915);
nand U24881 (N_24881,N_23018,N_23705);
nor U24882 (N_24882,N_23232,N_23597);
nand U24883 (N_24883,N_22816,N_23209);
nand U24884 (N_24884,N_23112,N_23319);
xor U24885 (N_24885,N_23657,N_23134);
nand U24886 (N_24886,N_23167,N_22600);
or U24887 (N_24887,N_23957,N_22940);
and U24888 (N_24888,N_23383,N_22620);
and U24889 (N_24889,N_23162,N_22620);
and U24890 (N_24890,N_23648,N_23404);
or U24891 (N_24891,N_23103,N_23574);
nor U24892 (N_24892,N_23592,N_23577);
or U24893 (N_24893,N_23414,N_23463);
xnor U24894 (N_24894,N_22727,N_23474);
or U24895 (N_24895,N_23439,N_23928);
nand U24896 (N_24896,N_22601,N_22781);
nand U24897 (N_24897,N_23431,N_22662);
nand U24898 (N_24898,N_23604,N_22649);
or U24899 (N_24899,N_23703,N_23427);
and U24900 (N_24900,N_22801,N_22760);
nand U24901 (N_24901,N_22567,N_23132);
xnor U24902 (N_24902,N_22695,N_23442);
nand U24903 (N_24903,N_23881,N_23056);
xor U24904 (N_24904,N_23630,N_23661);
xnor U24905 (N_24905,N_23053,N_22859);
nand U24906 (N_24906,N_23238,N_22967);
nor U24907 (N_24907,N_23913,N_22882);
nand U24908 (N_24908,N_23329,N_22641);
xor U24909 (N_24909,N_23059,N_22963);
nor U24910 (N_24910,N_23061,N_22824);
nor U24911 (N_24911,N_23934,N_23836);
nand U24912 (N_24912,N_23442,N_22710);
nand U24913 (N_24913,N_23801,N_22784);
nand U24914 (N_24914,N_23946,N_22917);
xnor U24915 (N_24915,N_23343,N_23454);
nor U24916 (N_24916,N_23936,N_23171);
nand U24917 (N_24917,N_23953,N_22983);
xor U24918 (N_24918,N_23514,N_23491);
nand U24919 (N_24919,N_23740,N_23169);
or U24920 (N_24920,N_23027,N_23485);
nor U24921 (N_24921,N_23572,N_23904);
and U24922 (N_24922,N_23573,N_23605);
nor U24923 (N_24923,N_23467,N_23440);
and U24924 (N_24924,N_22972,N_23219);
and U24925 (N_24925,N_22560,N_22904);
nor U24926 (N_24926,N_22757,N_22667);
nand U24927 (N_24927,N_23440,N_23375);
nor U24928 (N_24928,N_23334,N_22606);
or U24929 (N_24929,N_23502,N_23472);
nor U24930 (N_24930,N_23523,N_23644);
xor U24931 (N_24931,N_23208,N_23407);
nand U24932 (N_24932,N_23658,N_22766);
and U24933 (N_24933,N_23383,N_23127);
and U24934 (N_24934,N_23631,N_22573);
and U24935 (N_24935,N_23364,N_22875);
or U24936 (N_24936,N_23378,N_23015);
nor U24937 (N_24937,N_23769,N_23164);
xnor U24938 (N_24938,N_23650,N_23273);
nand U24939 (N_24939,N_22973,N_22823);
nor U24940 (N_24940,N_23169,N_22898);
xnor U24941 (N_24941,N_22958,N_23247);
nor U24942 (N_24942,N_23992,N_23090);
or U24943 (N_24943,N_22685,N_22672);
xor U24944 (N_24944,N_23216,N_23208);
or U24945 (N_24945,N_22950,N_22819);
xor U24946 (N_24946,N_23201,N_23839);
or U24947 (N_24947,N_23458,N_22508);
nor U24948 (N_24948,N_23912,N_22669);
nand U24949 (N_24949,N_22982,N_23575);
xnor U24950 (N_24950,N_23097,N_23259);
nand U24951 (N_24951,N_22904,N_22672);
nor U24952 (N_24952,N_22726,N_23263);
nand U24953 (N_24953,N_22957,N_23663);
or U24954 (N_24954,N_23382,N_22579);
xor U24955 (N_24955,N_23941,N_23268);
nor U24956 (N_24956,N_22778,N_23775);
and U24957 (N_24957,N_22537,N_23590);
nand U24958 (N_24958,N_22580,N_23549);
and U24959 (N_24959,N_23146,N_23268);
nor U24960 (N_24960,N_23989,N_23288);
xnor U24961 (N_24961,N_22871,N_22756);
nand U24962 (N_24962,N_23077,N_22924);
nand U24963 (N_24963,N_22973,N_23076);
and U24964 (N_24964,N_22938,N_22777);
nand U24965 (N_24965,N_23385,N_22800);
nand U24966 (N_24966,N_23285,N_23531);
or U24967 (N_24967,N_22958,N_22661);
or U24968 (N_24968,N_23725,N_23969);
nand U24969 (N_24969,N_22500,N_23071);
nor U24970 (N_24970,N_22856,N_22681);
and U24971 (N_24971,N_23202,N_22711);
and U24972 (N_24972,N_22687,N_23736);
nand U24973 (N_24973,N_23641,N_23698);
nand U24974 (N_24974,N_22936,N_23000);
nand U24975 (N_24975,N_23149,N_22781);
nand U24976 (N_24976,N_23555,N_22915);
or U24977 (N_24977,N_23315,N_23069);
nor U24978 (N_24978,N_22953,N_23335);
xor U24979 (N_24979,N_23396,N_22519);
xor U24980 (N_24980,N_23456,N_23004);
and U24981 (N_24981,N_23200,N_23514);
and U24982 (N_24982,N_23282,N_22675);
or U24983 (N_24983,N_22734,N_22688);
nand U24984 (N_24984,N_23461,N_23401);
or U24985 (N_24985,N_23530,N_23301);
or U24986 (N_24986,N_23993,N_23278);
and U24987 (N_24987,N_23753,N_22866);
nor U24988 (N_24988,N_22658,N_23990);
xnor U24989 (N_24989,N_22658,N_23860);
or U24990 (N_24990,N_22771,N_23578);
xor U24991 (N_24991,N_22609,N_22873);
nor U24992 (N_24992,N_22647,N_23968);
and U24993 (N_24993,N_22803,N_23992);
or U24994 (N_24994,N_22528,N_23493);
or U24995 (N_24995,N_23132,N_23872);
xnor U24996 (N_24996,N_23973,N_23027);
and U24997 (N_24997,N_23659,N_23415);
nor U24998 (N_24998,N_23569,N_23663);
nor U24999 (N_24999,N_22780,N_23609);
and U25000 (N_25000,N_23436,N_23536);
nor U25001 (N_25001,N_23564,N_23100);
or U25002 (N_25002,N_23603,N_23015);
and U25003 (N_25003,N_23118,N_23462);
or U25004 (N_25004,N_23751,N_22791);
nand U25005 (N_25005,N_22633,N_22972);
or U25006 (N_25006,N_23809,N_23524);
nor U25007 (N_25007,N_23674,N_23247);
xnor U25008 (N_25008,N_23634,N_22895);
and U25009 (N_25009,N_22829,N_23821);
or U25010 (N_25010,N_22601,N_23885);
nand U25011 (N_25011,N_22981,N_22944);
nor U25012 (N_25012,N_23952,N_23610);
nand U25013 (N_25013,N_22551,N_22817);
nor U25014 (N_25014,N_23532,N_22804);
or U25015 (N_25015,N_23616,N_23911);
and U25016 (N_25016,N_23482,N_23326);
nand U25017 (N_25017,N_23675,N_22898);
or U25018 (N_25018,N_23617,N_23442);
nand U25019 (N_25019,N_23220,N_22885);
and U25020 (N_25020,N_23169,N_23396);
or U25021 (N_25021,N_23294,N_23044);
xor U25022 (N_25022,N_23054,N_23850);
or U25023 (N_25023,N_23994,N_22894);
nor U25024 (N_25024,N_23934,N_22874);
nor U25025 (N_25025,N_23762,N_23480);
nand U25026 (N_25026,N_22846,N_23170);
nor U25027 (N_25027,N_22577,N_22631);
and U25028 (N_25028,N_23253,N_22510);
and U25029 (N_25029,N_23487,N_22783);
and U25030 (N_25030,N_22921,N_23809);
xnor U25031 (N_25031,N_22739,N_22999);
or U25032 (N_25032,N_22573,N_22785);
nor U25033 (N_25033,N_23995,N_23969);
or U25034 (N_25034,N_23844,N_23900);
nand U25035 (N_25035,N_22877,N_23947);
xnor U25036 (N_25036,N_23174,N_22622);
nor U25037 (N_25037,N_23657,N_22918);
nor U25038 (N_25038,N_23846,N_23394);
or U25039 (N_25039,N_23654,N_23938);
nor U25040 (N_25040,N_23694,N_23277);
xor U25041 (N_25041,N_23061,N_23345);
and U25042 (N_25042,N_23751,N_23042);
xor U25043 (N_25043,N_22852,N_23767);
or U25044 (N_25044,N_23651,N_23240);
nor U25045 (N_25045,N_22984,N_22718);
nand U25046 (N_25046,N_23051,N_23963);
and U25047 (N_25047,N_23812,N_23498);
or U25048 (N_25048,N_23528,N_23396);
and U25049 (N_25049,N_23179,N_23808);
nor U25050 (N_25050,N_23967,N_23269);
and U25051 (N_25051,N_23218,N_22634);
or U25052 (N_25052,N_23983,N_23484);
and U25053 (N_25053,N_23159,N_22693);
nor U25054 (N_25054,N_23481,N_23782);
xor U25055 (N_25055,N_23657,N_23120);
nor U25056 (N_25056,N_23053,N_22972);
nand U25057 (N_25057,N_22980,N_22564);
or U25058 (N_25058,N_23172,N_23379);
or U25059 (N_25059,N_22872,N_23620);
and U25060 (N_25060,N_23066,N_23920);
nand U25061 (N_25061,N_22616,N_22574);
and U25062 (N_25062,N_23627,N_23266);
nand U25063 (N_25063,N_23075,N_22887);
or U25064 (N_25064,N_23979,N_23412);
and U25065 (N_25065,N_23755,N_23988);
nand U25066 (N_25066,N_23687,N_23352);
and U25067 (N_25067,N_23060,N_22561);
xor U25068 (N_25068,N_22797,N_22609);
xor U25069 (N_25069,N_22581,N_23530);
and U25070 (N_25070,N_23850,N_22786);
nand U25071 (N_25071,N_23710,N_23467);
xor U25072 (N_25072,N_23433,N_22546);
xor U25073 (N_25073,N_23116,N_23093);
nor U25074 (N_25074,N_23654,N_23796);
nand U25075 (N_25075,N_23678,N_23958);
or U25076 (N_25076,N_23272,N_23083);
and U25077 (N_25077,N_22851,N_22821);
xnor U25078 (N_25078,N_23622,N_23186);
xor U25079 (N_25079,N_22707,N_22982);
and U25080 (N_25080,N_23362,N_23889);
xor U25081 (N_25081,N_23037,N_22657);
nand U25082 (N_25082,N_23517,N_22725);
xor U25083 (N_25083,N_22649,N_23064);
or U25084 (N_25084,N_23954,N_22582);
or U25085 (N_25085,N_23123,N_23215);
or U25086 (N_25086,N_23959,N_23938);
and U25087 (N_25087,N_23448,N_23293);
xor U25088 (N_25088,N_23210,N_23806);
or U25089 (N_25089,N_22830,N_22589);
nor U25090 (N_25090,N_23097,N_23688);
nor U25091 (N_25091,N_23486,N_23313);
nor U25092 (N_25092,N_23829,N_23370);
nand U25093 (N_25093,N_23732,N_23618);
nand U25094 (N_25094,N_23759,N_23788);
nand U25095 (N_25095,N_23705,N_23073);
or U25096 (N_25096,N_23985,N_23173);
or U25097 (N_25097,N_23106,N_22652);
and U25098 (N_25098,N_23562,N_23995);
nor U25099 (N_25099,N_23988,N_23157);
nand U25100 (N_25100,N_23753,N_22841);
nand U25101 (N_25101,N_23686,N_23181);
xor U25102 (N_25102,N_23724,N_22865);
nand U25103 (N_25103,N_23497,N_23333);
and U25104 (N_25104,N_22818,N_23380);
nand U25105 (N_25105,N_23293,N_23536);
nand U25106 (N_25106,N_23044,N_23281);
or U25107 (N_25107,N_23716,N_22978);
xnor U25108 (N_25108,N_23062,N_22905);
nor U25109 (N_25109,N_22776,N_22540);
nor U25110 (N_25110,N_22866,N_22634);
nor U25111 (N_25111,N_22564,N_23183);
nor U25112 (N_25112,N_23724,N_23757);
nor U25113 (N_25113,N_23839,N_23854);
nor U25114 (N_25114,N_22524,N_23381);
nor U25115 (N_25115,N_22577,N_22693);
and U25116 (N_25116,N_23696,N_23153);
xnor U25117 (N_25117,N_23525,N_22709);
xor U25118 (N_25118,N_23608,N_22971);
or U25119 (N_25119,N_22680,N_23486);
nand U25120 (N_25120,N_23664,N_23626);
or U25121 (N_25121,N_23546,N_22588);
and U25122 (N_25122,N_23835,N_23504);
xor U25123 (N_25123,N_23843,N_22723);
nand U25124 (N_25124,N_23114,N_23071);
and U25125 (N_25125,N_23208,N_23595);
xor U25126 (N_25126,N_23008,N_23661);
xnor U25127 (N_25127,N_23523,N_22942);
xnor U25128 (N_25128,N_23666,N_22799);
nor U25129 (N_25129,N_22723,N_23428);
xnor U25130 (N_25130,N_23647,N_22600);
and U25131 (N_25131,N_23752,N_23500);
nor U25132 (N_25132,N_23701,N_23265);
nor U25133 (N_25133,N_23823,N_23899);
and U25134 (N_25134,N_23202,N_23254);
xnor U25135 (N_25135,N_23967,N_23729);
and U25136 (N_25136,N_23318,N_23122);
xnor U25137 (N_25137,N_23529,N_23816);
xnor U25138 (N_25138,N_22554,N_22995);
nor U25139 (N_25139,N_23411,N_22576);
nand U25140 (N_25140,N_23989,N_23214);
nand U25141 (N_25141,N_23814,N_23013);
nor U25142 (N_25142,N_23763,N_23019);
or U25143 (N_25143,N_23779,N_23192);
nand U25144 (N_25144,N_22828,N_22887);
nor U25145 (N_25145,N_22789,N_23316);
or U25146 (N_25146,N_23909,N_23796);
nand U25147 (N_25147,N_23403,N_23489);
nor U25148 (N_25148,N_23529,N_23116);
xor U25149 (N_25149,N_22720,N_22598);
and U25150 (N_25150,N_23851,N_23010);
and U25151 (N_25151,N_23684,N_23577);
xnor U25152 (N_25152,N_22758,N_22819);
or U25153 (N_25153,N_23328,N_22567);
nor U25154 (N_25154,N_23804,N_22544);
nand U25155 (N_25155,N_23339,N_23950);
nor U25156 (N_25156,N_22838,N_22913);
xor U25157 (N_25157,N_22652,N_22992);
xnor U25158 (N_25158,N_22742,N_23738);
xor U25159 (N_25159,N_22838,N_23948);
nand U25160 (N_25160,N_22792,N_22807);
nor U25161 (N_25161,N_23058,N_23688);
xnor U25162 (N_25162,N_23044,N_22876);
or U25163 (N_25163,N_22816,N_23600);
nor U25164 (N_25164,N_23899,N_22893);
and U25165 (N_25165,N_22732,N_23329);
and U25166 (N_25166,N_23939,N_23267);
nor U25167 (N_25167,N_22987,N_23443);
and U25168 (N_25168,N_23617,N_23976);
xor U25169 (N_25169,N_23962,N_23056);
xnor U25170 (N_25170,N_23921,N_23225);
xnor U25171 (N_25171,N_22866,N_23800);
nand U25172 (N_25172,N_22689,N_22765);
nand U25173 (N_25173,N_23490,N_22576);
nor U25174 (N_25174,N_22697,N_23553);
or U25175 (N_25175,N_22980,N_23847);
xnor U25176 (N_25176,N_23624,N_23703);
nor U25177 (N_25177,N_23506,N_22919);
or U25178 (N_25178,N_22550,N_23535);
nor U25179 (N_25179,N_23574,N_23091);
and U25180 (N_25180,N_23238,N_23287);
nand U25181 (N_25181,N_23188,N_23202);
nor U25182 (N_25182,N_23834,N_23051);
nor U25183 (N_25183,N_23691,N_23334);
nor U25184 (N_25184,N_22820,N_23920);
nand U25185 (N_25185,N_22967,N_22729);
nand U25186 (N_25186,N_23645,N_23664);
nand U25187 (N_25187,N_23639,N_22975);
xor U25188 (N_25188,N_23833,N_23156);
nor U25189 (N_25189,N_22916,N_22625);
nand U25190 (N_25190,N_23810,N_22845);
or U25191 (N_25191,N_22691,N_23744);
or U25192 (N_25192,N_23523,N_23020);
nor U25193 (N_25193,N_22991,N_23741);
nand U25194 (N_25194,N_22956,N_23316);
or U25195 (N_25195,N_23978,N_23097);
and U25196 (N_25196,N_22589,N_23351);
and U25197 (N_25197,N_23104,N_23479);
nor U25198 (N_25198,N_23852,N_23783);
nor U25199 (N_25199,N_22640,N_22634);
nor U25200 (N_25200,N_22676,N_23621);
and U25201 (N_25201,N_23532,N_23348);
xnor U25202 (N_25202,N_22526,N_23858);
or U25203 (N_25203,N_22778,N_22635);
or U25204 (N_25204,N_23643,N_22917);
or U25205 (N_25205,N_22643,N_22706);
or U25206 (N_25206,N_23264,N_22733);
xor U25207 (N_25207,N_23895,N_22840);
nand U25208 (N_25208,N_23398,N_22690);
xor U25209 (N_25209,N_22975,N_23187);
and U25210 (N_25210,N_22860,N_23967);
xnor U25211 (N_25211,N_23632,N_23798);
or U25212 (N_25212,N_23743,N_22903);
and U25213 (N_25213,N_23957,N_22868);
nand U25214 (N_25214,N_23762,N_22558);
or U25215 (N_25215,N_22597,N_23844);
nor U25216 (N_25216,N_23167,N_23524);
nand U25217 (N_25217,N_23268,N_23476);
nand U25218 (N_25218,N_23931,N_22783);
nor U25219 (N_25219,N_22590,N_23707);
or U25220 (N_25220,N_22854,N_23706);
xor U25221 (N_25221,N_22683,N_22793);
nand U25222 (N_25222,N_23078,N_23213);
nor U25223 (N_25223,N_23091,N_22578);
xnor U25224 (N_25224,N_22988,N_23030);
xnor U25225 (N_25225,N_22641,N_23711);
xor U25226 (N_25226,N_22551,N_23233);
or U25227 (N_25227,N_23947,N_23428);
or U25228 (N_25228,N_22538,N_23879);
and U25229 (N_25229,N_23849,N_23181);
or U25230 (N_25230,N_23813,N_22549);
or U25231 (N_25231,N_22680,N_23294);
xor U25232 (N_25232,N_23342,N_22809);
and U25233 (N_25233,N_23154,N_23889);
nand U25234 (N_25234,N_22812,N_23817);
or U25235 (N_25235,N_23046,N_23838);
nand U25236 (N_25236,N_22982,N_23529);
nor U25237 (N_25237,N_23551,N_23671);
xnor U25238 (N_25238,N_22676,N_22747);
or U25239 (N_25239,N_23484,N_23972);
nand U25240 (N_25240,N_23590,N_23834);
xor U25241 (N_25241,N_23573,N_23221);
xnor U25242 (N_25242,N_22514,N_23365);
or U25243 (N_25243,N_23242,N_23539);
or U25244 (N_25244,N_23024,N_22722);
nand U25245 (N_25245,N_23034,N_22980);
or U25246 (N_25246,N_23060,N_22653);
nand U25247 (N_25247,N_22845,N_23444);
nand U25248 (N_25248,N_23701,N_22955);
or U25249 (N_25249,N_23419,N_23928);
nor U25250 (N_25250,N_23130,N_23308);
and U25251 (N_25251,N_22635,N_22682);
or U25252 (N_25252,N_22864,N_23141);
or U25253 (N_25253,N_23597,N_23525);
nor U25254 (N_25254,N_23029,N_23913);
xor U25255 (N_25255,N_22749,N_23300);
xnor U25256 (N_25256,N_23033,N_23200);
and U25257 (N_25257,N_22778,N_22961);
and U25258 (N_25258,N_23405,N_23359);
nor U25259 (N_25259,N_23006,N_22991);
or U25260 (N_25260,N_22505,N_23455);
and U25261 (N_25261,N_23182,N_23119);
or U25262 (N_25262,N_23738,N_22679);
xnor U25263 (N_25263,N_23286,N_22851);
or U25264 (N_25264,N_23315,N_23236);
and U25265 (N_25265,N_22855,N_23696);
xnor U25266 (N_25266,N_23559,N_23826);
nand U25267 (N_25267,N_23389,N_23267);
nor U25268 (N_25268,N_22642,N_23137);
nor U25269 (N_25269,N_23741,N_23465);
nand U25270 (N_25270,N_23841,N_23504);
and U25271 (N_25271,N_23476,N_23839);
and U25272 (N_25272,N_23229,N_23606);
or U25273 (N_25273,N_23122,N_22751);
or U25274 (N_25274,N_23802,N_22698);
nor U25275 (N_25275,N_22756,N_23946);
nor U25276 (N_25276,N_22988,N_22737);
xor U25277 (N_25277,N_23731,N_23958);
nand U25278 (N_25278,N_22778,N_23916);
xnor U25279 (N_25279,N_23181,N_22914);
nand U25280 (N_25280,N_23686,N_23374);
nor U25281 (N_25281,N_23064,N_22974);
xnor U25282 (N_25282,N_23323,N_23723);
and U25283 (N_25283,N_23751,N_22979);
nor U25284 (N_25284,N_23722,N_23371);
or U25285 (N_25285,N_23287,N_22901);
nor U25286 (N_25286,N_23108,N_22944);
nand U25287 (N_25287,N_22735,N_22844);
and U25288 (N_25288,N_23949,N_23567);
and U25289 (N_25289,N_22710,N_23745);
nand U25290 (N_25290,N_22575,N_22675);
and U25291 (N_25291,N_23194,N_23749);
nand U25292 (N_25292,N_22782,N_23566);
or U25293 (N_25293,N_23865,N_23848);
and U25294 (N_25294,N_23144,N_22623);
or U25295 (N_25295,N_23438,N_22590);
or U25296 (N_25296,N_23889,N_23723);
xnor U25297 (N_25297,N_22578,N_22707);
and U25298 (N_25298,N_23992,N_23456);
xnor U25299 (N_25299,N_22898,N_23614);
nor U25300 (N_25300,N_22887,N_23036);
and U25301 (N_25301,N_23950,N_23071);
and U25302 (N_25302,N_23286,N_23242);
xnor U25303 (N_25303,N_22696,N_22618);
nor U25304 (N_25304,N_23460,N_23674);
and U25305 (N_25305,N_23954,N_23645);
nand U25306 (N_25306,N_23219,N_22798);
xnor U25307 (N_25307,N_23719,N_23749);
or U25308 (N_25308,N_23596,N_23219);
xor U25309 (N_25309,N_22562,N_22534);
nand U25310 (N_25310,N_23541,N_22656);
nand U25311 (N_25311,N_22918,N_22880);
xnor U25312 (N_25312,N_23598,N_22773);
nand U25313 (N_25313,N_22950,N_23880);
xnor U25314 (N_25314,N_22765,N_23451);
nand U25315 (N_25315,N_23271,N_22930);
or U25316 (N_25316,N_22718,N_23929);
or U25317 (N_25317,N_23236,N_23857);
xor U25318 (N_25318,N_23678,N_22996);
nand U25319 (N_25319,N_22919,N_22760);
xnor U25320 (N_25320,N_23676,N_23426);
xnor U25321 (N_25321,N_22738,N_23254);
or U25322 (N_25322,N_23988,N_23227);
or U25323 (N_25323,N_23406,N_23420);
nor U25324 (N_25324,N_23781,N_22730);
xnor U25325 (N_25325,N_23352,N_23094);
xnor U25326 (N_25326,N_23573,N_22763);
xnor U25327 (N_25327,N_22994,N_23508);
nand U25328 (N_25328,N_22937,N_22898);
nand U25329 (N_25329,N_23973,N_23028);
or U25330 (N_25330,N_23444,N_22809);
nor U25331 (N_25331,N_22899,N_23840);
xor U25332 (N_25332,N_23205,N_23893);
nand U25333 (N_25333,N_23367,N_23249);
nand U25334 (N_25334,N_23677,N_23683);
nand U25335 (N_25335,N_23227,N_23708);
or U25336 (N_25336,N_22614,N_23244);
or U25337 (N_25337,N_22728,N_23813);
or U25338 (N_25338,N_23201,N_23773);
or U25339 (N_25339,N_23859,N_23281);
or U25340 (N_25340,N_23174,N_23814);
nand U25341 (N_25341,N_23798,N_22992);
nand U25342 (N_25342,N_22652,N_23510);
xor U25343 (N_25343,N_23162,N_23613);
nor U25344 (N_25344,N_22835,N_23011);
xor U25345 (N_25345,N_23277,N_22787);
xor U25346 (N_25346,N_23505,N_23256);
and U25347 (N_25347,N_23358,N_23789);
nor U25348 (N_25348,N_23670,N_23729);
or U25349 (N_25349,N_23669,N_23095);
nand U25350 (N_25350,N_22727,N_22750);
or U25351 (N_25351,N_23782,N_23200);
xnor U25352 (N_25352,N_22817,N_23548);
xnor U25353 (N_25353,N_23878,N_23271);
nor U25354 (N_25354,N_23371,N_23354);
nand U25355 (N_25355,N_23062,N_22647);
or U25356 (N_25356,N_22697,N_23627);
and U25357 (N_25357,N_23519,N_23208);
or U25358 (N_25358,N_23510,N_23491);
xnor U25359 (N_25359,N_23917,N_23615);
or U25360 (N_25360,N_23586,N_23612);
nor U25361 (N_25361,N_22872,N_22809);
xnor U25362 (N_25362,N_23622,N_23574);
and U25363 (N_25363,N_22966,N_22594);
nor U25364 (N_25364,N_23388,N_22519);
and U25365 (N_25365,N_23655,N_23131);
xnor U25366 (N_25366,N_22572,N_22837);
xnor U25367 (N_25367,N_23592,N_22856);
and U25368 (N_25368,N_23556,N_23060);
nor U25369 (N_25369,N_22727,N_23347);
or U25370 (N_25370,N_23780,N_23117);
xnor U25371 (N_25371,N_22858,N_23848);
nor U25372 (N_25372,N_22994,N_23311);
and U25373 (N_25373,N_23265,N_23969);
and U25374 (N_25374,N_22586,N_23993);
and U25375 (N_25375,N_23348,N_23646);
or U25376 (N_25376,N_22749,N_23316);
nor U25377 (N_25377,N_23418,N_22563);
or U25378 (N_25378,N_23310,N_23677);
nand U25379 (N_25379,N_23207,N_23201);
nor U25380 (N_25380,N_23584,N_22901);
nor U25381 (N_25381,N_22675,N_23864);
nand U25382 (N_25382,N_23209,N_22919);
nand U25383 (N_25383,N_23628,N_23752);
nor U25384 (N_25384,N_23091,N_22732);
nand U25385 (N_25385,N_22716,N_23603);
xnor U25386 (N_25386,N_23844,N_23974);
and U25387 (N_25387,N_22700,N_23564);
nor U25388 (N_25388,N_23223,N_22822);
nand U25389 (N_25389,N_23641,N_23683);
nor U25390 (N_25390,N_22957,N_23161);
xnor U25391 (N_25391,N_23747,N_23368);
nand U25392 (N_25392,N_23003,N_23122);
nor U25393 (N_25393,N_23532,N_23454);
nor U25394 (N_25394,N_23834,N_23374);
xor U25395 (N_25395,N_23051,N_22676);
xnor U25396 (N_25396,N_22534,N_23177);
or U25397 (N_25397,N_22948,N_23350);
nand U25398 (N_25398,N_22796,N_23817);
or U25399 (N_25399,N_22689,N_23653);
and U25400 (N_25400,N_23231,N_22593);
xor U25401 (N_25401,N_23730,N_22994);
or U25402 (N_25402,N_23077,N_23878);
or U25403 (N_25403,N_23287,N_22643);
xnor U25404 (N_25404,N_23193,N_23574);
and U25405 (N_25405,N_23386,N_23008);
nand U25406 (N_25406,N_23636,N_23409);
and U25407 (N_25407,N_22887,N_23296);
or U25408 (N_25408,N_23527,N_23503);
nand U25409 (N_25409,N_23746,N_22675);
or U25410 (N_25410,N_22962,N_23226);
nor U25411 (N_25411,N_23315,N_23031);
nand U25412 (N_25412,N_23861,N_23381);
nand U25413 (N_25413,N_23721,N_22605);
and U25414 (N_25414,N_23379,N_22573);
and U25415 (N_25415,N_22639,N_23438);
xor U25416 (N_25416,N_23215,N_22743);
xnor U25417 (N_25417,N_22791,N_23974);
or U25418 (N_25418,N_23596,N_23633);
xor U25419 (N_25419,N_22665,N_23710);
nor U25420 (N_25420,N_23751,N_23604);
or U25421 (N_25421,N_23555,N_22528);
xor U25422 (N_25422,N_23464,N_22708);
nand U25423 (N_25423,N_22914,N_23340);
and U25424 (N_25424,N_23907,N_22917);
xnor U25425 (N_25425,N_23611,N_23761);
nand U25426 (N_25426,N_23174,N_22968);
and U25427 (N_25427,N_23547,N_23615);
xnor U25428 (N_25428,N_23814,N_23167);
and U25429 (N_25429,N_23708,N_23329);
nor U25430 (N_25430,N_23467,N_23673);
nor U25431 (N_25431,N_23951,N_23714);
or U25432 (N_25432,N_22724,N_23429);
xnor U25433 (N_25433,N_23706,N_23411);
xor U25434 (N_25434,N_23277,N_22833);
nor U25435 (N_25435,N_22681,N_23767);
nand U25436 (N_25436,N_23076,N_23825);
and U25437 (N_25437,N_22783,N_22670);
nor U25438 (N_25438,N_23980,N_22867);
xnor U25439 (N_25439,N_23189,N_23952);
or U25440 (N_25440,N_22943,N_23821);
nor U25441 (N_25441,N_22905,N_23882);
and U25442 (N_25442,N_22612,N_23690);
nand U25443 (N_25443,N_22601,N_23540);
nand U25444 (N_25444,N_22570,N_23737);
and U25445 (N_25445,N_22612,N_22575);
or U25446 (N_25446,N_22828,N_23876);
and U25447 (N_25447,N_22788,N_22785);
and U25448 (N_25448,N_22890,N_23986);
nand U25449 (N_25449,N_23865,N_22537);
or U25450 (N_25450,N_22963,N_23210);
or U25451 (N_25451,N_23201,N_23161);
xor U25452 (N_25452,N_23449,N_22603);
nor U25453 (N_25453,N_22508,N_23001);
nor U25454 (N_25454,N_23958,N_22844);
xor U25455 (N_25455,N_22679,N_23653);
nor U25456 (N_25456,N_23896,N_22835);
nor U25457 (N_25457,N_22596,N_23959);
nor U25458 (N_25458,N_22778,N_22810);
or U25459 (N_25459,N_22835,N_23601);
xnor U25460 (N_25460,N_23664,N_23094);
and U25461 (N_25461,N_23271,N_23744);
nand U25462 (N_25462,N_23813,N_22984);
nor U25463 (N_25463,N_23495,N_23527);
or U25464 (N_25464,N_23992,N_23552);
and U25465 (N_25465,N_23978,N_22518);
nor U25466 (N_25466,N_23239,N_22724);
nor U25467 (N_25467,N_23900,N_23487);
nand U25468 (N_25468,N_22928,N_22718);
and U25469 (N_25469,N_22938,N_23842);
nor U25470 (N_25470,N_23996,N_23209);
xnor U25471 (N_25471,N_22678,N_23270);
nand U25472 (N_25472,N_23703,N_22717);
xnor U25473 (N_25473,N_23175,N_23689);
and U25474 (N_25474,N_23224,N_22933);
nand U25475 (N_25475,N_22611,N_23335);
or U25476 (N_25476,N_22855,N_23490);
and U25477 (N_25477,N_23035,N_22961);
xor U25478 (N_25478,N_23080,N_23350);
nand U25479 (N_25479,N_23529,N_22538);
nor U25480 (N_25480,N_22846,N_23930);
and U25481 (N_25481,N_22771,N_23829);
nand U25482 (N_25482,N_23383,N_23837);
or U25483 (N_25483,N_23300,N_23013);
and U25484 (N_25484,N_23316,N_22775);
or U25485 (N_25485,N_23034,N_23564);
or U25486 (N_25486,N_23538,N_23569);
and U25487 (N_25487,N_23505,N_23837);
nand U25488 (N_25488,N_22812,N_22948);
nor U25489 (N_25489,N_23804,N_23026);
nor U25490 (N_25490,N_23309,N_23637);
nand U25491 (N_25491,N_23502,N_23414);
nor U25492 (N_25492,N_22974,N_22517);
or U25493 (N_25493,N_22963,N_23189);
nor U25494 (N_25494,N_23052,N_23348);
or U25495 (N_25495,N_22932,N_23771);
nand U25496 (N_25496,N_22610,N_23537);
xor U25497 (N_25497,N_23088,N_23344);
and U25498 (N_25498,N_23566,N_22843);
or U25499 (N_25499,N_22602,N_23967);
nand U25500 (N_25500,N_25160,N_24287);
nand U25501 (N_25501,N_24028,N_24981);
xor U25502 (N_25502,N_24175,N_24870);
nor U25503 (N_25503,N_24563,N_24033);
and U25504 (N_25504,N_25194,N_24574);
nand U25505 (N_25505,N_24910,N_24898);
nor U25506 (N_25506,N_25089,N_25246);
xnor U25507 (N_25507,N_24513,N_25058);
xor U25508 (N_25508,N_25049,N_24707);
nor U25509 (N_25509,N_24820,N_24129);
nand U25510 (N_25510,N_24905,N_24190);
nand U25511 (N_25511,N_25038,N_24749);
nor U25512 (N_25512,N_24562,N_24647);
or U25513 (N_25513,N_24788,N_24181);
nor U25514 (N_25514,N_24236,N_25168);
nand U25515 (N_25515,N_24426,N_24775);
xnor U25516 (N_25516,N_25105,N_24161);
nor U25517 (N_25517,N_25346,N_24169);
nor U25518 (N_25518,N_24079,N_24078);
nand U25519 (N_25519,N_24572,N_24178);
and U25520 (N_25520,N_24812,N_24565);
nand U25521 (N_25521,N_24208,N_24609);
nor U25522 (N_25522,N_25399,N_24684);
nand U25523 (N_25523,N_24350,N_25141);
xnor U25524 (N_25524,N_24477,N_24994);
or U25525 (N_25525,N_24310,N_25006);
nand U25526 (N_25526,N_24652,N_25376);
xor U25527 (N_25527,N_24029,N_24501);
nand U25528 (N_25528,N_25473,N_24725);
nand U25529 (N_25529,N_25499,N_24457);
nand U25530 (N_25530,N_25215,N_24286);
nand U25531 (N_25531,N_24795,N_24309);
nor U25532 (N_25532,N_24663,N_24656);
nand U25533 (N_25533,N_24458,N_25358);
nor U25534 (N_25534,N_24638,N_25057);
nand U25535 (N_25535,N_24098,N_25437);
nor U25536 (N_25536,N_25101,N_24228);
nand U25537 (N_25537,N_25349,N_24952);
nor U25538 (N_25538,N_24438,N_24015);
and U25539 (N_25539,N_24533,N_25113);
xnor U25540 (N_25540,N_24382,N_25013);
nand U25541 (N_25541,N_24058,N_24641);
nor U25542 (N_25542,N_25324,N_25288);
nor U25543 (N_25543,N_24838,N_25207);
xnor U25544 (N_25544,N_24548,N_25118);
xnor U25545 (N_25545,N_25429,N_25279);
or U25546 (N_25546,N_25483,N_25237);
nor U25547 (N_25547,N_24315,N_24727);
xnor U25548 (N_25548,N_24846,N_25003);
and U25549 (N_25549,N_25181,N_24507);
xor U25550 (N_25550,N_25129,N_24949);
and U25551 (N_25551,N_24613,N_24209);
and U25552 (N_25552,N_25425,N_24882);
and U25553 (N_25553,N_24412,N_25334);
or U25554 (N_25554,N_25068,N_24833);
and U25555 (N_25555,N_25380,N_24489);
nor U25556 (N_25556,N_24871,N_24074);
or U25557 (N_25557,N_24000,N_24582);
nand U25558 (N_25558,N_25348,N_25083);
nand U25559 (N_25559,N_25387,N_25498);
nand U25560 (N_25560,N_24690,N_25480);
or U25561 (N_25561,N_24365,N_25420);
xnor U25562 (N_25562,N_25114,N_24366);
nand U25563 (N_25563,N_24005,N_25294);
nand U25564 (N_25564,N_24325,N_24878);
or U25565 (N_25565,N_25099,N_25412);
xor U25566 (N_25566,N_24134,N_25048);
nand U25567 (N_25567,N_24774,N_24768);
xnor U25568 (N_25568,N_25484,N_25209);
and U25569 (N_25569,N_25177,N_24577);
or U25570 (N_25570,N_24844,N_24759);
nor U25571 (N_25571,N_24353,N_25024);
xnor U25572 (N_25572,N_24492,N_24635);
nand U25573 (N_25573,N_24172,N_25463);
or U25574 (N_25574,N_25262,N_24256);
xnor U25575 (N_25575,N_24369,N_24423);
and U25576 (N_25576,N_24206,N_24218);
nand U25577 (N_25577,N_24012,N_24616);
nand U25578 (N_25578,N_25169,N_24446);
nand U25579 (N_25579,N_24255,N_24372);
nand U25580 (N_25580,N_24362,N_24050);
nand U25581 (N_25581,N_24816,N_24305);
and U25582 (N_25582,N_25197,N_24311);
nor U25583 (N_25583,N_25147,N_25328);
and U25584 (N_25584,N_24606,N_24648);
xnor U25585 (N_25585,N_24540,N_25450);
xor U25586 (N_25586,N_25243,N_24530);
or U25587 (N_25587,N_25180,N_24340);
and U25588 (N_25588,N_24063,N_24946);
nor U25589 (N_25589,N_25444,N_24850);
nor U25590 (N_25590,N_25000,N_24532);
nor U25591 (N_25591,N_24519,N_25043);
or U25592 (N_25592,N_24222,N_25224);
xor U25593 (N_25593,N_24117,N_24602);
xnor U25594 (N_25594,N_24116,N_24830);
and U25595 (N_25595,N_24784,N_24667);
nand U25596 (N_25596,N_24693,N_24048);
xnor U25597 (N_25597,N_24996,N_25347);
or U25598 (N_25598,N_24723,N_25316);
and U25599 (N_25599,N_24605,N_24284);
nor U25600 (N_25600,N_24894,N_24464);
xor U25601 (N_25601,N_24569,N_25015);
or U25602 (N_25602,N_24942,N_25385);
xor U25603 (N_25603,N_25223,N_24627);
and U25604 (N_25604,N_24734,N_24941);
or U25605 (N_25605,N_24651,N_24022);
xor U25606 (N_25606,N_24025,N_24418);
nand U25607 (N_25607,N_25152,N_24586);
xnor U25608 (N_25608,N_24358,N_24702);
and U25609 (N_25609,N_25367,N_24829);
nor U25610 (N_25610,N_25255,N_25302);
xor U25611 (N_25611,N_25023,N_24230);
or U25612 (N_25612,N_24819,N_25289);
and U25613 (N_25613,N_24568,N_24499);
nor U25614 (N_25614,N_24985,N_24804);
nor U25615 (N_25615,N_24375,N_24643);
nand U25616 (N_25616,N_24642,N_25005);
and U25617 (N_25617,N_24887,N_24626);
xor U25618 (N_25618,N_24096,N_24420);
nand U25619 (N_25619,N_24755,N_25475);
nor U25620 (N_25620,N_25104,N_24732);
or U25621 (N_25621,N_25047,N_24556);
and U25622 (N_25622,N_24120,N_24242);
nor U25623 (N_25623,N_24488,N_24696);
and U25624 (N_25624,N_25256,N_24460);
xnor U25625 (N_25625,N_25155,N_25326);
xnor U25626 (N_25626,N_24908,N_24197);
xor U25627 (N_25627,N_25016,N_25350);
and U25628 (N_25628,N_24594,N_24007);
or U25629 (N_25629,N_24925,N_25336);
nand U25630 (N_25630,N_24671,N_24566);
nand U25631 (N_25631,N_25474,N_25035);
or U25632 (N_25632,N_24840,N_24171);
xor U25633 (N_25633,N_24813,N_24858);
nor U25634 (N_25634,N_24302,N_24828);
xnor U25635 (N_25635,N_25364,N_25492);
xor U25636 (N_25636,N_24183,N_24611);
nor U25637 (N_25637,N_25053,N_25183);
or U25638 (N_25638,N_24738,N_24392);
nor U25639 (N_25639,N_25112,N_24097);
and U25640 (N_25640,N_25198,N_24947);
xnor U25641 (N_25641,N_24416,N_24006);
xor U25642 (N_25642,N_24924,N_24409);
or U25643 (N_25643,N_24188,N_24436);
or U25644 (N_25644,N_24351,N_25490);
nor U25645 (N_25645,N_24285,N_24735);
and U25646 (N_25646,N_25185,N_25186);
nand U25647 (N_25647,N_24966,N_24902);
xnor U25648 (N_25648,N_24590,N_25396);
and U25649 (N_25649,N_25471,N_24751);
nand U25650 (N_25650,N_24921,N_25199);
or U25651 (N_25651,N_24388,N_24090);
and U25652 (N_25652,N_25264,N_25402);
and U25653 (N_25653,N_25284,N_24034);
and U25654 (N_25654,N_24786,N_24071);
or U25655 (N_25655,N_25460,N_25027);
or U25656 (N_25656,N_24655,N_25007);
nand U25657 (N_25657,N_25071,N_24010);
nand U25658 (N_25658,N_25355,N_24543);
nand U25659 (N_25659,N_24137,N_24212);
xor U25660 (N_25660,N_24695,N_25494);
nor U25661 (N_25661,N_25405,N_25190);
nand U25662 (N_25662,N_24639,N_24537);
nor U25663 (N_25663,N_24632,N_24658);
nand U25664 (N_25664,N_25029,N_24155);
xor U25665 (N_25665,N_24739,N_25455);
nand U25666 (N_25666,N_24988,N_24849);
nand U25667 (N_25667,N_24066,N_24177);
nand U25668 (N_25668,N_25375,N_24296);
nor U25669 (N_25669,N_25332,N_25046);
and U25670 (N_25670,N_25457,N_24918);
and U25671 (N_25671,N_24754,N_24356);
and U25672 (N_25672,N_25366,N_24879);
xor U25673 (N_25673,N_24794,N_24328);
and U25674 (N_25674,N_25384,N_25272);
xor U25675 (N_25675,N_24893,N_25028);
nand U25676 (N_25676,N_24598,N_24538);
and U25677 (N_25677,N_24054,N_25157);
nand U25678 (N_25678,N_25461,N_25259);
nor U25679 (N_25679,N_24043,N_25218);
nor U25680 (N_25680,N_24146,N_24791);
or U25681 (N_25681,N_24553,N_24825);
or U25682 (N_25682,N_25395,N_24984);
nor U25683 (N_25683,N_24099,N_24928);
nand U25684 (N_25684,N_24486,N_24313);
xnor U25685 (N_25685,N_24341,N_24835);
xnor U25686 (N_25686,N_24152,N_25430);
xor U25687 (N_25687,N_25022,N_25496);
nand U25688 (N_25688,N_24250,N_24468);
nor U25689 (N_25689,N_24432,N_24571);
and U25690 (N_25690,N_24500,N_24783);
xor U25691 (N_25691,N_24083,N_25001);
nand U25692 (N_25692,N_25351,N_24159);
nor U25693 (N_25693,N_25454,N_24357);
and U25694 (N_25694,N_24861,N_24240);
xor U25695 (N_25695,N_24772,N_24459);
nor U25696 (N_25696,N_24604,N_24980);
nor U25697 (N_25697,N_24856,N_24619);
nor U25698 (N_25698,N_25196,N_24480);
or U25699 (N_25699,N_24132,N_24195);
xnor U25700 (N_25700,N_25100,N_24895);
nand U25701 (N_25701,N_24281,N_25251);
nor U25702 (N_25702,N_24251,N_24168);
and U25703 (N_25703,N_24558,N_25136);
or U25704 (N_25704,N_25070,N_24024);
nor U25705 (N_25705,N_24913,N_25314);
xor U25706 (N_25706,N_24650,N_24347);
or U25707 (N_25707,N_24121,N_25214);
and U25708 (N_25708,N_24207,N_24922);
nand U25709 (N_25709,N_24312,N_24860);
or U25710 (N_25710,N_24086,N_24017);
nor U25711 (N_25711,N_24964,N_24403);
or U25712 (N_25712,N_24761,N_25369);
nor U25713 (N_25713,N_24634,N_24731);
nor U25714 (N_25714,N_24127,N_24442);
nand U25715 (N_25715,N_25370,N_24705);
xnor U25716 (N_25716,N_24189,N_24425);
nand U25717 (N_25717,N_24750,N_24308);
or U25718 (N_25718,N_24244,N_25149);
and U25719 (N_25719,N_24187,N_24135);
and U25720 (N_25720,N_24515,N_24093);
or U25721 (N_25721,N_24441,N_25159);
nand U25722 (N_25722,N_24371,N_24184);
and U25723 (N_25723,N_24520,N_25365);
and U25724 (N_25724,N_25133,N_24956);
nand U25725 (N_25725,N_24623,N_25495);
and U25726 (N_25726,N_25291,N_25252);
nand U25727 (N_25727,N_24151,N_24379);
xnor U25728 (N_25728,N_25254,N_24797);
and U25729 (N_25729,N_24317,N_24258);
nor U25730 (N_25730,N_24672,N_24247);
nand U25731 (N_25731,N_25482,N_24527);
xnor U25732 (N_25732,N_24587,N_24395);
xnor U25733 (N_25733,N_25121,N_24766);
nand U25734 (N_25734,N_24322,N_24386);
or U25735 (N_25735,N_25139,N_25145);
nand U25736 (N_25736,N_25312,N_24581);
nand U25737 (N_25737,N_24953,N_25012);
and U25738 (N_25738,N_25311,N_24790);
and U25739 (N_25739,N_24975,N_24331);
nand U25740 (N_25740,N_24496,N_24473);
and U25741 (N_25741,N_25257,N_25459);
and U25742 (N_25742,N_24937,N_24927);
or U25743 (N_25743,N_24254,N_24199);
nand U25744 (N_25744,N_24465,N_25076);
nor U25745 (N_25745,N_24186,N_25322);
and U25746 (N_25746,N_24675,N_25127);
or U25747 (N_25747,N_25195,N_25344);
nor U25748 (N_25748,N_24481,N_24274);
nor U25749 (N_25749,N_24900,N_24660);
nor U25750 (N_25750,N_24698,N_24510);
or U25751 (N_25751,N_25435,N_25452);
nor U25752 (N_25752,N_25270,N_25416);
or U25753 (N_25753,N_24402,N_24710);
xnor U25754 (N_25754,N_25325,N_24711);
or U25755 (N_25755,N_24881,N_24567);
nand U25756 (N_25756,N_24373,N_24760);
and U25757 (N_25757,N_24689,N_25067);
xnor U25758 (N_25758,N_24487,N_25230);
and U25759 (N_25759,N_24545,N_24780);
or U25760 (N_25760,N_24077,N_24039);
xor U25761 (N_25761,N_24396,N_25032);
and U25762 (N_25762,N_24677,N_24073);
and U25763 (N_25763,N_24799,N_24536);
nand U25764 (N_25764,N_24055,N_24541);
or U25765 (N_25765,N_24076,N_24728);
xnor U25766 (N_25766,N_24943,N_24534);
nor U25767 (N_25767,N_24235,N_25407);
nor U25768 (N_25768,N_25134,N_24597);
xnor U25769 (N_25769,N_24843,N_24821);
and U25770 (N_25770,N_24471,N_24469);
and U25771 (N_25771,N_24360,N_25439);
and U25772 (N_25772,N_25078,N_24801);
and U25773 (N_25773,N_25318,N_25410);
nor U25774 (N_25774,N_24747,N_24721);
nor U25775 (N_25775,N_24709,N_24032);
and U25776 (N_25776,N_25392,N_24729);
nor U25777 (N_25777,N_25161,N_24903);
xnor U25778 (N_25778,N_25073,N_25271);
nor U25779 (N_25779,N_24278,N_25080);
xnor U25780 (N_25780,N_24165,N_24384);
xnor U25781 (N_25781,N_24557,N_24770);
and U25782 (N_25782,N_24084,N_24339);
and U25783 (N_25783,N_24268,N_24345);
nand U25784 (N_25784,N_24726,N_24649);
and U25785 (N_25785,N_24706,N_24899);
nor U25786 (N_25786,N_24115,N_24931);
nor U25787 (N_25787,N_24653,N_24008);
xor U25788 (N_25788,N_25247,N_24466);
nor U25789 (N_25789,N_24904,N_24257);
or U25790 (N_25790,N_24011,N_24020);
nor U25791 (N_25791,N_25382,N_25119);
nand U25792 (N_25792,N_24319,N_25300);
or U25793 (N_25793,N_24912,N_24888);
nand U25794 (N_25794,N_24915,N_24971);
xnor U25795 (N_25795,N_25431,N_25229);
nor U25796 (N_25796,N_24511,N_25278);
nor U25797 (N_25797,N_24260,N_25356);
or U25798 (N_25798,N_25036,N_24238);
or U25799 (N_25799,N_24685,N_25010);
and U25800 (N_25800,N_24779,N_24225);
or U25801 (N_25801,N_24827,N_24991);
or U25802 (N_25802,N_24264,N_24892);
nor U25803 (N_25803,N_24699,N_24810);
xnor U25804 (N_25804,N_24045,N_24781);
nor U25805 (N_25805,N_25135,N_24676);
or U25806 (N_25806,N_24529,N_24013);
and U25807 (N_25807,N_25438,N_24917);
xnor U25808 (N_25808,N_24853,N_25319);
nand U25809 (N_25809,N_24620,N_24524);
nor U25810 (N_25810,N_24320,N_25309);
nor U25811 (N_25811,N_24243,N_24363);
or U25812 (N_25812,N_24452,N_25335);
nor U25813 (N_25813,N_24348,N_24631);
or U25814 (N_25814,N_24205,N_24216);
and U25815 (N_25815,N_25060,N_24472);
nand U25816 (N_25816,N_25493,N_25017);
and U25817 (N_25817,N_25333,N_24805);
and U25818 (N_25818,N_24976,N_25260);
or U25819 (N_25819,N_24769,N_24118);
or U25820 (N_25820,N_25087,N_24753);
nand U25821 (N_25821,N_24934,N_24992);
nor U25822 (N_25822,N_25175,N_24682);
nor U25823 (N_25823,N_24431,N_24686);
nor U25824 (N_25824,N_25025,N_25063);
nand U25825 (N_25825,N_24989,N_24393);
and U25826 (N_25826,N_25434,N_25306);
nand U25827 (N_25827,N_24164,N_25166);
xnor U25828 (N_25828,N_25059,N_24595);
nand U25829 (N_25829,N_24221,N_25329);
nand U25830 (N_25830,N_24578,N_24792);
and U25831 (N_25831,N_24683,N_24108);
and U25832 (N_25832,N_24326,N_24292);
and U25833 (N_25833,N_24198,N_25307);
or U25834 (N_25834,N_24051,N_24318);
or U25835 (N_25835,N_24831,N_24807);
xor U25836 (N_25836,N_24234,N_24521);
or U25837 (N_25837,N_25283,N_24239);
nor U25838 (N_25838,N_24368,N_25212);
or U25839 (N_25839,N_24282,N_24119);
xnor U25840 (N_25840,N_25249,N_25258);
xnor U25841 (N_25841,N_24935,N_24483);
and U25842 (N_25842,N_24035,N_24219);
nor U25843 (N_25843,N_24607,N_25045);
or U25844 (N_25844,N_24525,N_24376);
xnor U25845 (N_25845,N_24950,N_24301);
and U25846 (N_25846,N_25228,N_24454);
or U25847 (N_25847,N_24461,N_25189);
nor U25848 (N_25848,N_24026,N_25363);
nand U25849 (N_25849,N_24518,N_24998);
nand U25850 (N_25850,N_25021,N_24246);
and U25851 (N_25851,N_25019,N_24665);
nor U25852 (N_25852,N_25377,N_24911);
xnor U25853 (N_25853,N_24802,N_24990);
or U25854 (N_25854,N_24584,N_25220);
and U25855 (N_25855,N_24273,N_25303);
xnor U25856 (N_25856,N_24703,N_24479);
and U25857 (N_25857,N_24113,N_25341);
nand U25858 (N_25858,N_25128,N_25476);
nor U25859 (N_25859,N_25154,N_24704);
nor U25860 (N_25860,N_24453,N_24491);
nand U25861 (N_25861,N_24736,N_24385);
nand U25862 (N_25862,N_24060,N_25478);
xor U25863 (N_25863,N_24232,N_24352);
xnor U25864 (N_25864,N_24842,N_24618);
xnor U25865 (N_25865,N_24776,N_24270);
or U25866 (N_25866,N_24107,N_24072);
and U25867 (N_25867,N_24874,N_24640);
xor U25868 (N_25868,N_24406,N_24062);
xnor U25869 (N_25869,N_25123,N_25193);
nor U25870 (N_25870,N_25342,N_24397);
nor U25871 (N_25871,N_25170,N_25188);
xor U25872 (N_25872,N_24700,N_25360);
xnor U25873 (N_25873,N_24275,N_25041);
nor U25874 (N_25874,N_25276,N_24245);
and U25875 (N_25875,N_24068,N_25372);
and U25876 (N_25876,N_24601,N_24789);
nor U25877 (N_25877,N_24758,N_24104);
xor U25878 (N_25878,N_25359,N_25440);
nand U25879 (N_25879,N_24049,N_24016);
nand U25880 (N_25880,N_25225,N_25208);
xor U25881 (N_25881,N_24087,N_24939);
nor U25882 (N_25882,N_24229,N_24973);
xor U25883 (N_25883,N_24873,N_25020);
xor U25884 (N_25884,N_24413,N_25443);
or U25885 (N_25885,N_25253,N_25432);
and U25886 (N_25886,N_24977,N_25200);
xor U25887 (N_25887,N_25040,N_25448);
nand U25888 (N_25888,N_24958,N_25394);
nor U25889 (N_25889,N_24252,N_25315);
or U25890 (N_25890,N_25422,N_25442);
or U25891 (N_25891,N_24191,N_24440);
or U25892 (N_25892,N_24869,N_25092);
nor U25893 (N_25893,N_24724,N_24213);
nor U25894 (N_25894,N_24001,N_24859);
nand U25895 (N_25895,N_24681,N_24031);
nand U25896 (N_25896,N_24865,N_24451);
or U25897 (N_25897,N_24476,N_24414);
xnor U25898 (N_25898,N_24144,N_25222);
nor U25899 (N_25899,N_24929,N_24153);
nand U25900 (N_25900,N_24387,N_24624);
nor U25901 (N_25901,N_24231,N_24933);
and U25902 (N_25902,N_25340,N_24692);
nand U25903 (N_25903,N_24475,N_24854);
xor U25904 (N_25904,N_25406,N_24503);
xnor U25905 (N_25905,N_25339,N_24847);
nand U25906 (N_25906,N_24333,N_25240);
or U25907 (N_25907,N_25345,N_24439);
nand U25908 (N_25908,N_24517,N_24944);
and U25909 (N_25909,N_24421,N_25096);
nand U25910 (N_25910,N_24085,N_24972);
nand U25911 (N_25911,N_24336,N_25102);
xnor U25912 (N_25912,N_25491,N_25162);
nand U25913 (N_25913,N_24433,N_24614);
nor U25914 (N_25914,N_25091,N_24617);
nand U25915 (N_25915,N_24160,N_24139);
or U25916 (N_25916,N_24818,N_24349);
or U25917 (N_25917,N_24528,N_24550);
and U25918 (N_25918,N_24004,N_25378);
nand U25919 (N_25919,N_25368,N_25227);
xnor U25920 (N_25920,N_24809,N_24437);
nor U25921 (N_25921,N_24030,N_24694);
nor U25922 (N_25922,N_24561,N_24484);
and U25923 (N_25923,N_24448,N_25107);
nor U25924 (N_25924,N_25153,N_24424);
nor U25925 (N_25925,N_25117,N_24997);
and U25926 (N_25926,N_24002,N_25462);
xnor U25927 (N_25927,N_24542,N_24067);
nand U25928 (N_25928,N_25427,N_24193);
and U25929 (N_25929,N_24599,N_24771);
or U25930 (N_25930,N_24133,N_25282);
nand U25931 (N_25931,N_25115,N_25146);
xor U25932 (N_25932,N_25409,N_24657);
or U25933 (N_25933,N_25374,N_24088);
xnor U25934 (N_25934,N_24344,N_25267);
nor U25935 (N_25935,N_24263,N_24400);
xnor U25936 (N_25936,N_25174,N_24410);
or U25937 (N_25937,N_25469,N_25415);
and U25938 (N_25938,N_24678,N_24822);
or U25939 (N_25939,N_24192,N_24056);
or U25940 (N_25940,N_24109,N_24294);
xnor U25941 (N_25941,N_24215,N_24936);
or U25942 (N_25942,N_25379,N_25011);
nor U25943 (N_25943,N_24535,N_24307);
nand U25944 (N_25944,N_24334,N_24555);
nor U25945 (N_25945,N_25479,N_25280);
nor U25946 (N_25946,N_24450,N_25217);
nand U25947 (N_25947,N_24401,N_24354);
nand U25948 (N_25948,N_24951,N_24265);
and U25949 (N_25949,N_25082,N_24730);
and U25950 (N_25950,N_24637,N_24271);
nand U25951 (N_25951,N_24196,N_24482);
xnor U25952 (N_25952,N_24708,N_24891);
xnor U25953 (N_25953,N_24575,N_25304);
or U25954 (N_25954,N_24938,N_24886);
nand U25955 (N_25955,N_24744,N_24130);
nor U25956 (N_25956,N_25125,N_24211);
and U25957 (N_25957,N_25298,N_24262);
or U25958 (N_25958,N_24064,N_24162);
and U25959 (N_25959,N_24343,N_25213);
and U25960 (N_25960,N_24335,N_24907);
xor U25961 (N_25961,N_25414,N_24210);
xor U25962 (N_25962,N_24081,N_25261);
and U25963 (N_25963,N_24963,N_24687);
nand U25964 (N_25964,N_24154,N_24680);
and U25965 (N_25965,N_24298,N_25293);
nand U25966 (N_25966,N_24095,N_25287);
nand U25967 (N_25967,N_24866,N_24737);
nand U25968 (N_25968,N_24633,N_24701);
and U25969 (N_25969,N_25037,N_24291);
xnor U25970 (N_25970,N_24662,N_24559);
xor U25971 (N_25971,N_25064,N_24897);
nand U25972 (N_25972,N_25468,N_24009);
nor U25973 (N_25973,N_24815,N_24447);
nand U25974 (N_25974,N_25203,N_24143);
or U25975 (N_25975,N_24102,N_24122);
xnor U25976 (N_25976,N_24583,N_25362);
xnor U25977 (N_25977,N_25488,N_24014);
xor U25978 (N_25978,N_24201,N_24733);
xnor U25979 (N_25979,N_24740,N_25090);
and U25980 (N_25980,N_24712,N_25292);
or U25981 (N_25981,N_24722,N_25381);
nor U25982 (N_25982,N_24128,N_24743);
or U25983 (N_25983,N_25487,N_24621);
nand U25984 (N_25984,N_24969,N_24800);
and U25985 (N_25985,N_25056,N_25026);
xor U25986 (N_25986,N_24070,N_24855);
nand U25987 (N_25987,N_24919,N_24636);
xor U25988 (N_25988,N_25352,N_24679);
and U25989 (N_25989,N_24509,N_25130);
nand U25990 (N_25990,N_24837,N_24493);
xnor U25991 (N_25991,N_24316,N_24608);
nand U25992 (N_25992,N_24463,N_24306);
nor U25993 (N_25993,N_24741,N_24174);
or U25994 (N_25994,N_24126,N_24715);
nor U25995 (N_25995,N_25239,N_25120);
nand U25996 (N_25996,N_24042,N_24166);
and U25997 (N_25997,N_24044,N_24124);
nand U25998 (N_25998,N_24848,N_24147);
xor U25999 (N_25999,N_25338,N_25248);
nand U26000 (N_26000,N_25132,N_24596);
or U26001 (N_26001,N_25299,N_24038);
nor U26002 (N_26002,N_25131,N_25393);
nand U26003 (N_26003,N_25167,N_24478);
xor U26004 (N_26004,N_24445,N_24047);
xnor U26005 (N_26005,N_24082,N_25313);
nand U26006 (N_26006,N_25211,N_24717);
and U26007 (N_26007,N_24506,N_24645);
nand U26008 (N_26008,N_25173,N_24415);
nor U26009 (N_26009,N_25150,N_25466);
nor U26010 (N_26010,N_24092,N_24422);
nand U26011 (N_26011,N_25226,N_24808);
nand U26012 (N_26012,N_24714,N_25004);
nand U26013 (N_26013,N_25373,N_25337);
or U26014 (N_26014,N_25386,N_24052);
and U26015 (N_26015,N_24374,N_25093);
and U26016 (N_26016,N_24877,N_24290);
nand U26017 (N_26017,N_25171,N_25327);
and U26018 (N_26018,N_24021,N_25232);
or U26019 (N_26019,N_24765,N_24389);
and U26020 (N_26020,N_24430,N_25202);
nand U26021 (N_26021,N_25424,N_24823);
nor U26022 (N_26022,N_25441,N_25108);
and U26023 (N_26023,N_25447,N_25054);
xor U26024 (N_26024,N_25330,N_24142);
xnor U26025 (N_26025,N_25317,N_25467);
nor U26026 (N_26026,N_24670,N_24955);
nand U26027 (N_26027,N_24691,N_25285);
and U26028 (N_26028,N_25266,N_24644);
nor U26029 (N_26029,N_24628,N_24945);
nand U26030 (N_26030,N_25297,N_24993);
or U26031 (N_26031,N_25400,N_25403);
xor U26032 (N_26032,N_24355,N_25163);
or U26033 (N_26033,N_24136,N_24688);
xor U26034 (N_26034,N_24961,N_24592);
or U26035 (N_26035,N_25310,N_24960);
xor U26036 (N_26036,N_24674,N_24516);
nor U26037 (N_26037,N_24327,N_24867);
or U26038 (N_26038,N_24585,N_25397);
and U26039 (N_26039,N_24381,N_24610);
or U26040 (N_26040,N_24249,N_25343);
or U26041 (N_26041,N_24075,N_24417);
or U26042 (N_26042,N_24456,N_24974);
and U26043 (N_26043,N_24125,N_24223);
xor U26044 (N_26044,N_25497,N_24544);
nor U26045 (N_26045,N_25050,N_25428);
xor U26046 (N_26046,N_24580,N_24277);
nor U26047 (N_26047,N_25137,N_24539);
nand U26048 (N_26048,N_24470,N_24982);
xnor U26049 (N_26049,N_25235,N_24342);
or U26050 (N_26050,N_25086,N_24906);
xor U26051 (N_26051,N_24826,N_24300);
xnor U26052 (N_26052,N_24986,N_24752);
and U26053 (N_26053,N_25201,N_25275);
nor U26054 (N_26054,N_25323,N_25072);
or U26055 (N_26055,N_24018,N_25353);
or U26056 (N_26056,N_24720,N_24046);
xnor U26057 (N_26057,N_25419,N_24338);
xor U26058 (N_26058,N_25398,N_24554);
xnor U26059 (N_26059,N_25204,N_24814);
or U26060 (N_26060,N_25408,N_24367);
and U26061 (N_26061,N_25030,N_24272);
or U26062 (N_26062,N_25453,N_25061);
and U26063 (N_26063,N_24156,N_24449);
nor U26064 (N_26064,N_24764,N_24289);
or U26065 (N_26065,N_24773,N_24612);
and U26066 (N_26066,N_24303,N_25178);
nor U26067 (N_26067,N_25305,N_24757);
and U26068 (N_26068,N_25095,N_24176);
or U26069 (N_26069,N_24023,N_24547);
nand U26070 (N_26070,N_24661,N_25233);
nor U26071 (N_26071,N_24748,N_25269);
or U26072 (N_26072,N_24576,N_24100);
nor U26073 (N_26073,N_24940,N_24965);
and U26074 (N_26074,N_24839,N_24782);
xnor U26075 (N_26075,N_24817,N_24803);
nand U26076 (N_26076,N_25485,N_25172);
xor U26077 (N_26077,N_24896,N_24123);
and U26078 (N_26078,N_24883,N_24408);
or U26079 (N_26079,N_24824,N_24180);
or U26080 (N_26080,N_24279,N_24920);
or U26081 (N_26081,N_25320,N_25151);
nor U26082 (N_26082,N_24505,N_25401);
and U26083 (N_26083,N_24630,N_25308);
or U26084 (N_26084,N_24405,N_25124);
nand U26085 (N_26085,N_24485,N_25144);
xor U26086 (N_26086,N_24170,N_24293);
nor U26087 (N_26087,N_24194,N_24314);
nor U26088 (N_26088,N_25489,N_24872);
or U26089 (N_26089,N_25081,N_25074);
or U26090 (N_26090,N_25051,N_24202);
nand U26091 (N_26091,N_24259,N_25423);
nor U26092 (N_26092,N_24615,N_24182);
nor U26093 (N_26093,N_24467,N_24659);
or U26094 (N_26094,N_24299,N_24959);
and U26095 (N_26095,N_24057,N_25458);
nor U26096 (N_26096,N_25085,N_24359);
nand U26097 (N_26097,N_25109,N_24570);
nand U26098 (N_26098,N_25357,N_24149);
nor U26099 (N_26099,N_24462,N_24037);
and U26100 (N_26100,N_24157,N_25417);
nand U26101 (N_26101,N_24220,N_25002);
or U26102 (N_26102,N_24173,N_24253);
and U26103 (N_26103,N_24167,N_24889);
xnor U26104 (N_26104,N_25273,N_24114);
nand U26105 (N_26105,N_24080,N_24217);
xnor U26106 (N_26106,N_24065,N_24718);
and U26107 (N_26107,N_24150,N_24280);
xnor U26108 (N_26108,N_25103,N_25242);
and U26109 (N_26109,N_25097,N_25206);
or U26110 (N_26110,N_25079,N_25277);
nand U26111 (N_26111,N_25238,N_25296);
xnor U26112 (N_26112,N_24323,N_24836);
xnor U26113 (N_26113,N_25371,N_24968);
and U26114 (N_26114,N_24995,N_24185);
nand U26115 (N_26115,N_24668,N_25052);
nand U26116 (N_26116,N_24664,N_24796);
xnor U26117 (N_26117,N_24832,N_25014);
or U26118 (N_26118,N_24746,N_24512);
or U26119 (N_26119,N_25165,N_24398);
or U26120 (N_26120,N_24145,N_25456);
nor U26121 (N_26121,N_24233,N_25433);
xor U26122 (N_26122,N_25472,N_24380);
and U26123 (N_26123,N_25158,N_25390);
xor U26124 (N_26124,N_24564,N_24967);
nand U26125 (N_26125,N_24622,N_25009);
xnor U26126 (N_26126,N_25033,N_25250);
or U26127 (N_26127,N_24868,N_25421);
nor U26128 (N_26128,N_25470,N_24444);
or U26129 (N_26129,N_25236,N_24110);
nor U26130 (N_26130,N_24200,N_24502);
xnor U26131 (N_26131,N_25031,N_24923);
or U26132 (N_26132,N_25274,N_24138);
nand U26133 (N_26133,N_24103,N_25465);
or U26134 (N_26134,N_24391,N_25116);
or U26135 (N_26135,N_25404,N_24697);
or U26136 (N_26136,N_25066,N_24716);
or U26137 (N_26137,N_25069,N_24742);
nor U26138 (N_26138,N_25055,N_24756);
nor U26139 (N_26139,N_25034,N_24111);
and U26140 (N_26140,N_25383,N_24589);
or U26141 (N_26141,N_24916,N_25219);
or U26142 (N_26142,N_24112,N_24666);
xor U26143 (N_26143,N_24498,N_24494);
and U26144 (N_26144,N_25263,N_24105);
or U26145 (N_26145,N_24158,N_25187);
nand U26146 (N_26146,N_24793,N_24531);
or U26147 (N_26147,N_25354,N_24983);
nor U26148 (N_26148,N_24834,N_24591);
nand U26149 (N_26149,N_25391,N_25077);
xnor U26150 (N_26150,N_25140,N_24909);
or U26151 (N_26151,N_25301,N_24094);
xnor U26152 (N_26152,N_25042,N_24852);
nor U26153 (N_26153,N_24745,N_25182);
nor U26154 (N_26154,N_24875,N_24266);
and U26155 (N_26155,N_25221,N_24261);
and U26156 (N_26156,N_24719,N_25205);
nand U26157 (N_26157,N_24926,N_24394);
and U26158 (N_26158,N_24061,N_24880);
xnor U26159 (N_26159,N_24876,N_25290);
and U26160 (N_26160,N_24329,N_24862);
nand U26161 (N_26161,N_25106,N_24845);
nor U26162 (N_26162,N_24851,N_24003);
nand U26163 (N_26163,N_24864,N_25184);
or U26164 (N_26164,N_24593,N_24713);
nor U26165 (N_26165,N_25436,N_24522);
nand U26166 (N_26166,N_24954,N_24579);
nand U26167 (N_26167,N_25268,N_24321);
or U26168 (N_26168,N_25142,N_24979);
nand U26169 (N_26169,N_24419,N_24407);
or U26170 (N_26170,N_24885,N_24283);
xor U26171 (N_26171,N_24669,N_24490);
or U26172 (N_26172,N_24361,N_24495);
or U26173 (N_26173,N_24163,N_24364);
nand U26174 (N_26174,N_24434,N_24370);
nand U26175 (N_26175,N_24549,N_24552);
nand U26176 (N_26176,N_25110,N_24377);
nand U26177 (N_26177,N_24089,N_24806);
nor U26178 (N_26178,N_24588,N_24514);
xnor U26179 (N_26179,N_24767,N_25111);
or U26180 (N_26180,N_25445,N_24654);
nor U26181 (N_26181,N_24560,N_24332);
nand U26182 (N_26182,N_25481,N_24019);
or U26183 (N_26183,N_25138,N_24508);
nor U26184 (N_26184,N_24600,N_24646);
or U26185 (N_26185,N_25244,N_25065);
xnor U26186 (N_26186,N_25331,N_24890);
nor U26187 (N_26187,N_24404,N_25192);
xnor U26188 (N_26188,N_24248,N_25084);
xor U26189 (N_26189,N_24497,N_24504);
xnor U26190 (N_26190,N_25148,N_25241);
nand U26191 (N_26191,N_25075,N_24932);
nor U26192 (N_26192,N_24383,N_25426);
or U26193 (N_26193,N_24987,N_24276);
nand U26194 (N_26194,N_25179,N_25449);
and U26195 (N_26195,N_24295,N_24041);
nand U26196 (N_26196,N_24036,N_25210);
nand U26197 (N_26197,N_24297,N_24241);
nand U26198 (N_26198,N_24179,N_24857);
nor U26199 (N_26199,N_24390,N_25286);
and U26200 (N_26200,N_25464,N_24978);
nor U26201 (N_26201,N_24267,N_24140);
or U26202 (N_26202,N_24428,N_25098);
nand U26203 (N_26203,N_25156,N_25122);
or U26204 (N_26204,N_24040,N_24551);
nor U26205 (N_26205,N_24901,N_24573);
xnor U26206 (N_26206,N_24673,N_24059);
nand U26207 (N_26207,N_24999,N_25295);
or U26208 (N_26208,N_25321,N_24841);
nor U26209 (N_26209,N_25088,N_24798);
and U26210 (N_26210,N_24204,N_24762);
xor U26211 (N_26211,N_24930,N_25191);
or U26212 (N_26212,N_25451,N_25018);
and U26213 (N_26213,N_24884,N_25281);
nor U26214 (N_26214,N_24224,N_24227);
nand U26215 (N_26215,N_25477,N_24330);
nand U26216 (N_26216,N_24948,N_24427);
and U26217 (N_26217,N_24324,N_24269);
nand U26218 (N_26218,N_24763,N_25411);
nand U26219 (N_26219,N_25486,N_24777);
xnor U26220 (N_26220,N_25176,N_24091);
or U26221 (N_26221,N_25008,N_24787);
or U26222 (N_26222,N_24785,N_24288);
or U26223 (N_26223,N_25094,N_24962);
xor U26224 (N_26224,N_24346,N_24526);
and U26225 (N_26225,N_24148,N_25389);
nor U26226 (N_26226,N_25143,N_24811);
nor U26227 (N_26227,N_24429,N_24337);
xor U26228 (N_26228,N_24435,N_24474);
nor U26229 (N_26229,N_24629,N_24443);
xnor U26230 (N_26230,N_25418,N_24411);
nand U26231 (N_26231,N_24141,N_24027);
xnor U26232 (N_26232,N_25446,N_25413);
xnor U26233 (N_26233,N_25039,N_24203);
nand U26234 (N_26234,N_24131,N_25062);
and U26235 (N_26235,N_24778,N_24101);
or U26236 (N_26236,N_24603,N_24237);
xnor U26237 (N_26237,N_24863,N_25234);
xnor U26238 (N_26238,N_24625,N_24546);
nand U26239 (N_26239,N_24226,N_25216);
nor U26240 (N_26240,N_24957,N_25265);
nand U26241 (N_26241,N_25126,N_25388);
nor U26242 (N_26242,N_25231,N_24455);
xor U26243 (N_26243,N_24970,N_24914);
xor U26244 (N_26244,N_25044,N_25361);
nand U26245 (N_26245,N_24214,N_24053);
nor U26246 (N_26246,N_24069,N_24106);
xor U26247 (N_26247,N_24523,N_25245);
or U26248 (N_26248,N_25164,N_24378);
xor U26249 (N_26249,N_24304,N_24399);
and U26250 (N_26250,N_24074,N_24680);
nor U26251 (N_26251,N_24714,N_24851);
nand U26252 (N_26252,N_24971,N_24726);
nand U26253 (N_26253,N_24360,N_24307);
and U26254 (N_26254,N_25360,N_24908);
nor U26255 (N_26255,N_24123,N_24810);
nor U26256 (N_26256,N_25341,N_24120);
nor U26257 (N_26257,N_24444,N_25206);
or U26258 (N_26258,N_25429,N_25125);
nor U26259 (N_26259,N_24361,N_24452);
nand U26260 (N_26260,N_24718,N_24136);
nor U26261 (N_26261,N_24155,N_25448);
and U26262 (N_26262,N_24361,N_24394);
or U26263 (N_26263,N_24121,N_24667);
nor U26264 (N_26264,N_25001,N_24286);
nor U26265 (N_26265,N_24714,N_24584);
or U26266 (N_26266,N_24070,N_25186);
xor U26267 (N_26267,N_24161,N_24334);
nand U26268 (N_26268,N_25090,N_25303);
nor U26269 (N_26269,N_24072,N_25279);
and U26270 (N_26270,N_24542,N_24329);
nand U26271 (N_26271,N_25192,N_24085);
xor U26272 (N_26272,N_24020,N_24054);
and U26273 (N_26273,N_25116,N_25470);
xor U26274 (N_26274,N_25494,N_25265);
and U26275 (N_26275,N_24772,N_25144);
and U26276 (N_26276,N_24265,N_25248);
and U26277 (N_26277,N_24981,N_25304);
nand U26278 (N_26278,N_24868,N_24671);
nand U26279 (N_26279,N_25010,N_24874);
xnor U26280 (N_26280,N_25165,N_25458);
nor U26281 (N_26281,N_24902,N_24827);
and U26282 (N_26282,N_25350,N_24660);
or U26283 (N_26283,N_24249,N_24947);
nand U26284 (N_26284,N_24218,N_25445);
nand U26285 (N_26285,N_24662,N_24597);
xnor U26286 (N_26286,N_24618,N_25202);
nor U26287 (N_26287,N_24344,N_24800);
nor U26288 (N_26288,N_25300,N_25464);
or U26289 (N_26289,N_25031,N_24178);
nand U26290 (N_26290,N_24120,N_24993);
xnor U26291 (N_26291,N_24364,N_25383);
xor U26292 (N_26292,N_25303,N_24882);
nand U26293 (N_26293,N_24394,N_25359);
xnor U26294 (N_26294,N_24206,N_24822);
nand U26295 (N_26295,N_24171,N_25482);
nand U26296 (N_26296,N_25080,N_25147);
xor U26297 (N_26297,N_24955,N_25113);
xnor U26298 (N_26298,N_24588,N_24426);
nand U26299 (N_26299,N_25098,N_24839);
xor U26300 (N_26300,N_24390,N_25193);
nor U26301 (N_26301,N_24627,N_24361);
or U26302 (N_26302,N_24924,N_24291);
xnor U26303 (N_26303,N_24364,N_24956);
xor U26304 (N_26304,N_24113,N_24859);
nand U26305 (N_26305,N_24759,N_25447);
and U26306 (N_26306,N_24737,N_25166);
nand U26307 (N_26307,N_25098,N_25326);
nor U26308 (N_26308,N_25181,N_25220);
nand U26309 (N_26309,N_24854,N_24077);
or U26310 (N_26310,N_24138,N_24337);
xnor U26311 (N_26311,N_24630,N_24108);
and U26312 (N_26312,N_24637,N_24949);
nor U26313 (N_26313,N_24890,N_25112);
nand U26314 (N_26314,N_24787,N_24159);
xnor U26315 (N_26315,N_25218,N_24365);
nand U26316 (N_26316,N_24617,N_24978);
xnor U26317 (N_26317,N_24480,N_24589);
nand U26318 (N_26318,N_24274,N_24947);
xnor U26319 (N_26319,N_24927,N_25265);
or U26320 (N_26320,N_24591,N_24024);
nor U26321 (N_26321,N_24060,N_24579);
xnor U26322 (N_26322,N_24812,N_24116);
nand U26323 (N_26323,N_25268,N_24718);
and U26324 (N_26324,N_24382,N_24474);
nor U26325 (N_26325,N_24460,N_24651);
or U26326 (N_26326,N_24373,N_24666);
nor U26327 (N_26327,N_24356,N_24764);
nor U26328 (N_26328,N_24360,N_24127);
or U26329 (N_26329,N_24813,N_25246);
xnor U26330 (N_26330,N_25307,N_24911);
xnor U26331 (N_26331,N_24478,N_25496);
nand U26332 (N_26332,N_24680,N_24000);
nand U26333 (N_26333,N_25164,N_24297);
xnor U26334 (N_26334,N_25277,N_25364);
nor U26335 (N_26335,N_24827,N_24636);
nor U26336 (N_26336,N_25305,N_24004);
nor U26337 (N_26337,N_25050,N_24041);
xor U26338 (N_26338,N_24888,N_24047);
or U26339 (N_26339,N_24105,N_24605);
nand U26340 (N_26340,N_24020,N_24355);
nand U26341 (N_26341,N_24642,N_25465);
xor U26342 (N_26342,N_24883,N_24597);
xnor U26343 (N_26343,N_24538,N_24249);
or U26344 (N_26344,N_24128,N_25410);
and U26345 (N_26345,N_25458,N_24713);
xnor U26346 (N_26346,N_24647,N_24675);
nor U26347 (N_26347,N_25181,N_24030);
nand U26348 (N_26348,N_25092,N_24129);
xor U26349 (N_26349,N_24066,N_24727);
nand U26350 (N_26350,N_25185,N_25368);
and U26351 (N_26351,N_24555,N_25462);
or U26352 (N_26352,N_25350,N_24838);
or U26353 (N_26353,N_24595,N_24740);
nor U26354 (N_26354,N_24481,N_24519);
nand U26355 (N_26355,N_24438,N_24462);
or U26356 (N_26356,N_24248,N_24934);
nor U26357 (N_26357,N_25006,N_24192);
or U26358 (N_26358,N_24820,N_24639);
nor U26359 (N_26359,N_24581,N_24940);
xor U26360 (N_26360,N_24562,N_25205);
nor U26361 (N_26361,N_25416,N_25492);
nand U26362 (N_26362,N_24107,N_24293);
or U26363 (N_26363,N_24496,N_24640);
nand U26364 (N_26364,N_25426,N_24304);
or U26365 (N_26365,N_24389,N_25446);
xor U26366 (N_26366,N_24912,N_24462);
or U26367 (N_26367,N_25039,N_24081);
and U26368 (N_26368,N_24899,N_25077);
xnor U26369 (N_26369,N_24557,N_24279);
nand U26370 (N_26370,N_24139,N_24056);
nor U26371 (N_26371,N_24855,N_24965);
xnor U26372 (N_26372,N_24844,N_24576);
xor U26373 (N_26373,N_25067,N_25215);
xnor U26374 (N_26374,N_24513,N_24631);
xor U26375 (N_26375,N_24865,N_24757);
nand U26376 (N_26376,N_24441,N_25303);
nor U26377 (N_26377,N_25364,N_24662);
xor U26378 (N_26378,N_24492,N_24847);
or U26379 (N_26379,N_24413,N_24397);
and U26380 (N_26380,N_25281,N_24573);
xor U26381 (N_26381,N_24680,N_24028);
xnor U26382 (N_26382,N_24739,N_24960);
nor U26383 (N_26383,N_25169,N_25445);
and U26384 (N_26384,N_24533,N_25347);
or U26385 (N_26385,N_24689,N_24103);
or U26386 (N_26386,N_25064,N_24931);
nor U26387 (N_26387,N_24433,N_25476);
nor U26388 (N_26388,N_25195,N_24019);
and U26389 (N_26389,N_24006,N_25250);
nor U26390 (N_26390,N_25063,N_25381);
and U26391 (N_26391,N_25244,N_24057);
and U26392 (N_26392,N_24556,N_24631);
nand U26393 (N_26393,N_24530,N_24849);
or U26394 (N_26394,N_25166,N_25173);
or U26395 (N_26395,N_24770,N_24461);
nand U26396 (N_26396,N_25381,N_24055);
and U26397 (N_26397,N_24029,N_24520);
nand U26398 (N_26398,N_24969,N_24737);
or U26399 (N_26399,N_25275,N_25088);
and U26400 (N_26400,N_24039,N_24080);
nand U26401 (N_26401,N_25254,N_24995);
nand U26402 (N_26402,N_24368,N_24580);
nand U26403 (N_26403,N_24577,N_24057);
nor U26404 (N_26404,N_24040,N_24793);
or U26405 (N_26405,N_24912,N_24875);
or U26406 (N_26406,N_24410,N_24678);
nor U26407 (N_26407,N_24874,N_25229);
and U26408 (N_26408,N_25039,N_25404);
and U26409 (N_26409,N_24845,N_24303);
or U26410 (N_26410,N_24510,N_25050);
nand U26411 (N_26411,N_25343,N_24620);
and U26412 (N_26412,N_24483,N_24521);
nor U26413 (N_26413,N_24356,N_24823);
xnor U26414 (N_26414,N_24082,N_24169);
nand U26415 (N_26415,N_24719,N_24578);
and U26416 (N_26416,N_24045,N_25026);
or U26417 (N_26417,N_25002,N_24547);
nor U26418 (N_26418,N_25002,N_24327);
and U26419 (N_26419,N_24425,N_25209);
nor U26420 (N_26420,N_25406,N_25002);
xnor U26421 (N_26421,N_24509,N_24531);
and U26422 (N_26422,N_24678,N_24805);
or U26423 (N_26423,N_25047,N_25464);
nand U26424 (N_26424,N_24242,N_24816);
xor U26425 (N_26425,N_25263,N_25276);
nand U26426 (N_26426,N_24013,N_24422);
xor U26427 (N_26427,N_24753,N_25043);
and U26428 (N_26428,N_24583,N_24131);
nor U26429 (N_26429,N_24115,N_24543);
xor U26430 (N_26430,N_25286,N_25283);
xor U26431 (N_26431,N_25271,N_24382);
and U26432 (N_26432,N_24682,N_24822);
and U26433 (N_26433,N_25319,N_24967);
or U26434 (N_26434,N_25483,N_24695);
xnor U26435 (N_26435,N_24557,N_24237);
and U26436 (N_26436,N_24117,N_24782);
and U26437 (N_26437,N_24188,N_24549);
nand U26438 (N_26438,N_25147,N_24926);
nor U26439 (N_26439,N_25321,N_25393);
and U26440 (N_26440,N_24151,N_25085);
nand U26441 (N_26441,N_24789,N_24740);
and U26442 (N_26442,N_24435,N_25421);
nor U26443 (N_26443,N_24146,N_24018);
and U26444 (N_26444,N_25382,N_25248);
nor U26445 (N_26445,N_25235,N_24628);
xor U26446 (N_26446,N_24532,N_25173);
nand U26447 (N_26447,N_24623,N_24029);
or U26448 (N_26448,N_24438,N_25414);
and U26449 (N_26449,N_25384,N_24797);
and U26450 (N_26450,N_24650,N_24275);
nand U26451 (N_26451,N_24768,N_25337);
or U26452 (N_26452,N_25053,N_25007);
and U26453 (N_26453,N_24841,N_24790);
or U26454 (N_26454,N_24644,N_25337);
xor U26455 (N_26455,N_24953,N_25176);
nor U26456 (N_26456,N_24831,N_24329);
nand U26457 (N_26457,N_25246,N_25266);
and U26458 (N_26458,N_24277,N_24040);
xnor U26459 (N_26459,N_24497,N_24197);
xor U26460 (N_26460,N_24465,N_25057);
xor U26461 (N_26461,N_24100,N_24591);
xnor U26462 (N_26462,N_25147,N_25307);
or U26463 (N_26463,N_24273,N_25176);
xnor U26464 (N_26464,N_24932,N_24985);
and U26465 (N_26465,N_25249,N_25430);
nand U26466 (N_26466,N_24377,N_24180);
and U26467 (N_26467,N_24105,N_25364);
or U26468 (N_26468,N_24374,N_24663);
nor U26469 (N_26469,N_24583,N_25370);
nand U26470 (N_26470,N_25474,N_24014);
xor U26471 (N_26471,N_24381,N_24192);
xnor U26472 (N_26472,N_24910,N_25176);
nor U26473 (N_26473,N_25179,N_24859);
or U26474 (N_26474,N_25137,N_24433);
or U26475 (N_26475,N_24720,N_25283);
and U26476 (N_26476,N_24596,N_24061);
nand U26477 (N_26477,N_24409,N_24790);
nor U26478 (N_26478,N_24190,N_24203);
xor U26479 (N_26479,N_25312,N_24696);
nand U26480 (N_26480,N_24784,N_25194);
nand U26481 (N_26481,N_25414,N_24303);
nand U26482 (N_26482,N_24267,N_24929);
nand U26483 (N_26483,N_24012,N_25042);
xor U26484 (N_26484,N_24476,N_25059);
xnor U26485 (N_26485,N_24708,N_25005);
nand U26486 (N_26486,N_24795,N_24126);
nor U26487 (N_26487,N_24374,N_25137);
nand U26488 (N_26488,N_24164,N_24475);
and U26489 (N_26489,N_24776,N_24659);
nor U26490 (N_26490,N_25130,N_24684);
xor U26491 (N_26491,N_24515,N_25015);
xor U26492 (N_26492,N_25342,N_24468);
nand U26493 (N_26493,N_24094,N_24011);
nand U26494 (N_26494,N_24573,N_24272);
nand U26495 (N_26495,N_24486,N_24219);
nor U26496 (N_26496,N_24562,N_24278);
or U26497 (N_26497,N_24226,N_24239);
nand U26498 (N_26498,N_24174,N_25427);
nand U26499 (N_26499,N_24218,N_25004);
xnor U26500 (N_26500,N_24502,N_24725);
xnor U26501 (N_26501,N_24570,N_24464);
or U26502 (N_26502,N_24624,N_24606);
or U26503 (N_26503,N_24904,N_24055);
nand U26504 (N_26504,N_24807,N_24710);
xnor U26505 (N_26505,N_24914,N_25191);
and U26506 (N_26506,N_24205,N_24879);
nor U26507 (N_26507,N_25439,N_24767);
and U26508 (N_26508,N_24672,N_24449);
nand U26509 (N_26509,N_24860,N_24601);
nor U26510 (N_26510,N_24550,N_24079);
nor U26511 (N_26511,N_24874,N_25459);
or U26512 (N_26512,N_25461,N_24433);
nor U26513 (N_26513,N_24027,N_24877);
nor U26514 (N_26514,N_24466,N_24193);
xnor U26515 (N_26515,N_25091,N_25444);
nor U26516 (N_26516,N_25309,N_24349);
nand U26517 (N_26517,N_24637,N_24734);
xor U26518 (N_26518,N_25357,N_24229);
or U26519 (N_26519,N_24188,N_24739);
or U26520 (N_26520,N_25335,N_24175);
nor U26521 (N_26521,N_24803,N_25357);
xor U26522 (N_26522,N_25408,N_24294);
and U26523 (N_26523,N_24479,N_24996);
nor U26524 (N_26524,N_24287,N_25090);
xnor U26525 (N_26525,N_24551,N_25169);
nor U26526 (N_26526,N_25176,N_24235);
and U26527 (N_26527,N_24655,N_24776);
xnor U26528 (N_26528,N_24696,N_25327);
and U26529 (N_26529,N_25244,N_25004);
nor U26530 (N_26530,N_24724,N_24185);
and U26531 (N_26531,N_24676,N_24542);
or U26532 (N_26532,N_25262,N_24054);
xor U26533 (N_26533,N_25243,N_24241);
nand U26534 (N_26534,N_24196,N_24923);
nor U26535 (N_26535,N_24260,N_25318);
nand U26536 (N_26536,N_24721,N_24193);
and U26537 (N_26537,N_24144,N_25439);
nor U26538 (N_26538,N_24541,N_24051);
nor U26539 (N_26539,N_25048,N_24790);
nand U26540 (N_26540,N_24957,N_24091);
or U26541 (N_26541,N_25169,N_24165);
nor U26542 (N_26542,N_24958,N_25439);
or U26543 (N_26543,N_24146,N_25135);
and U26544 (N_26544,N_24545,N_24353);
nand U26545 (N_26545,N_25393,N_24798);
nor U26546 (N_26546,N_25493,N_24997);
and U26547 (N_26547,N_25447,N_24547);
xnor U26548 (N_26548,N_25411,N_24260);
and U26549 (N_26549,N_24226,N_25375);
nor U26550 (N_26550,N_25226,N_24398);
nor U26551 (N_26551,N_24142,N_24974);
and U26552 (N_26552,N_24064,N_25402);
and U26553 (N_26553,N_24695,N_24617);
and U26554 (N_26554,N_25482,N_24228);
nand U26555 (N_26555,N_24736,N_24530);
nand U26556 (N_26556,N_25143,N_25066);
nand U26557 (N_26557,N_25379,N_24003);
and U26558 (N_26558,N_24322,N_25174);
nand U26559 (N_26559,N_24364,N_25223);
nor U26560 (N_26560,N_24523,N_25272);
nor U26561 (N_26561,N_24657,N_25167);
and U26562 (N_26562,N_24448,N_24038);
and U26563 (N_26563,N_24419,N_24371);
and U26564 (N_26564,N_24608,N_24098);
or U26565 (N_26565,N_24035,N_24521);
nand U26566 (N_26566,N_24811,N_25070);
and U26567 (N_26567,N_25290,N_25171);
xor U26568 (N_26568,N_24077,N_24832);
nor U26569 (N_26569,N_24576,N_24649);
or U26570 (N_26570,N_25319,N_24266);
and U26571 (N_26571,N_25197,N_24845);
nand U26572 (N_26572,N_24652,N_25336);
nand U26573 (N_26573,N_24067,N_24015);
and U26574 (N_26574,N_24841,N_24274);
or U26575 (N_26575,N_24503,N_25069);
and U26576 (N_26576,N_25146,N_25219);
nand U26577 (N_26577,N_25399,N_24736);
xor U26578 (N_26578,N_24180,N_24001);
xnor U26579 (N_26579,N_25348,N_25175);
and U26580 (N_26580,N_24175,N_25088);
nor U26581 (N_26581,N_24380,N_24229);
nand U26582 (N_26582,N_24989,N_25376);
and U26583 (N_26583,N_24022,N_24060);
or U26584 (N_26584,N_25441,N_24132);
xnor U26585 (N_26585,N_24174,N_24084);
or U26586 (N_26586,N_25373,N_24762);
nor U26587 (N_26587,N_24128,N_24603);
nand U26588 (N_26588,N_24119,N_24297);
or U26589 (N_26589,N_25078,N_24382);
and U26590 (N_26590,N_24711,N_25165);
and U26591 (N_26591,N_25059,N_24507);
or U26592 (N_26592,N_25332,N_25403);
nor U26593 (N_26593,N_24321,N_24539);
or U26594 (N_26594,N_25469,N_25046);
and U26595 (N_26595,N_24541,N_25056);
or U26596 (N_26596,N_25211,N_24500);
and U26597 (N_26597,N_25443,N_24788);
or U26598 (N_26598,N_24070,N_25324);
and U26599 (N_26599,N_24295,N_25154);
or U26600 (N_26600,N_24641,N_24137);
and U26601 (N_26601,N_25170,N_24001);
xor U26602 (N_26602,N_24400,N_24169);
nor U26603 (N_26603,N_24854,N_25157);
nor U26604 (N_26604,N_25206,N_25027);
nand U26605 (N_26605,N_25195,N_24868);
and U26606 (N_26606,N_25445,N_24786);
xnor U26607 (N_26607,N_24709,N_24129);
xor U26608 (N_26608,N_24167,N_24849);
nand U26609 (N_26609,N_25092,N_25432);
and U26610 (N_26610,N_24331,N_25087);
nor U26611 (N_26611,N_24051,N_25151);
nand U26612 (N_26612,N_25163,N_25482);
nand U26613 (N_26613,N_24258,N_25337);
nor U26614 (N_26614,N_24933,N_24046);
and U26615 (N_26615,N_24759,N_25464);
and U26616 (N_26616,N_24214,N_25405);
or U26617 (N_26617,N_24630,N_25310);
nor U26618 (N_26618,N_25000,N_24616);
or U26619 (N_26619,N_24985,N_24023);
or U26620 (N_26620,N_24875,N_24788);
or U26621 (N_26621,N_24686,N_25098);
or U26622 (N_26622,N_25196,N_24025);
or U26623 (N_26623,N_24887,N_24355);
and U26624 (N_26624,N_24320,N_24684);
xnor U26625 (N_26625,N_24732,N_25308);
nor U26626 (N_26626,N_25001,N_25315);
nand U26627 (N_26627,N_24373,N_24838);
xnor U26628 (N_26628,N_25484,N_24947);
nand U26629 (N_26629,N_25374,N_24380);
xor U26630 (N_26630,N_24134,N_25467);
or U26631 (N_26631,N_24596,N_24716);
nand U26632 (N_26632,N_24467,N_25273);
nand U26633 (N_26633,N_24061,N_24565);
nor U26634 (N_26634,N_25093,N_25209);
xor U26635 (N_26635,N_24594,N_24644);
and U26636 (N_26636,N_25055,N_24964);
xor U26637 (N_26637,N_24109,N_24734);
nor U26638 (N_26638,N_25494,N_24744);
or U26639 (N_26639,N_24455,N_25097);
or U26640 (N_26640,N_24239,N_24290);
nand U26641 (N_26641,N_24258,N_25441);
and U26642 (N_26642,N_24482,N_24844);
nor U26643 (N_26643,N_24215,N_25121);
xor U26644 (N_26644,N_24847,N_25044);
nor U26645 (N_26645,N_24599,N_25289);
or U26646 (N_26646,N_24038,N_24720);
or U26647 (N_26647,N_24288,N_24205);
nand U26648 (N_26648,N_24151,N_24341);
nand U26649 (N_26649,N_24921,N_24664);
and U26650 (N_26650,N_25347,N_24863);
or U26651 (N_26651,N_25321,N_24072);
nor U26652 (N_26652,N_25073,N_24791);
xnor U26653 (N_26653,N_24852,N_25190);
nand U26654 (N_26654,N_25185,N_24396);
xor U26655 (N_26655,N_24099,N_25116);
nor U26656 (N_26656,N_24453,N_24965);
and U26657 (N_26657,N_25000,N_24357);
or U26658 (N_26658,N_24697,N_24751);
and U26659 (N_26659,N_24868,N_25277);
xnor U26660 (N_26660,N_24612,N_24091);
and U26661 (N_26661,N_24682,N_24920);
xor U26662 (N_26662,N_24228,N_25270);
and U26663 (N_26663,N_24861,N_24993);
nor U26664 (N_26664,N_25018,N_24352);
nor U26665 (N_26665,N_24976,N_24486);
xor U26666 (N_26666,N_25438,N_24045);
or U26667 (N_26667,N_25222,N_24977);
xor U26668 (N_26668,N_25316,N_25383);
nor U26669 (N_26669,N_25454,N_25319);
nor U26670 (N_26670,N_24794,N_24414);
xor U26671 (N_26671,N_25219,N_24219);
and U26672 (N_26672,N_25380,N_25038);
nor U26673 (N_26673,N_24137,N_24823);
nor U26674 (N_26674,N_24682,N_25484);
xor U26675 (N_26675,N_24315,N_24098);
and U26676 (N_26676,N_25327,N_24270);
nor U26677 (N_26677,N_24911,N_24765);
xnor U26678 (N_26678,N_24606,N_25072);
xnor U26679 (N_26679,N_24718,N_24234);
xnor U26680 (N_26680,N_24598,N_24634);
xnor U26681 (N_26681,N_24277,N_25285);
or U26682 (N_26682,N_24011,N_24996);
nor U26683 (N_26683,N_24392,N_24047);
nor U26684 (N_26684,N_24093,N_25377);
or U26685 (N_26685,N_25455,N_25314);
xor U26686 (N_26686,N_25266,N_25279);
nand U26687 (N_26687,N_24463,N_24800);
or U26688 (N_26688,N_24298,N_25075);
or U26689 (N_26689,N_25415,N_24748);
nor U26690 (N_26690,N_24775,N_25177);
nor U26691 (N_26691,N_24406,N_24531);
nand U26692 (N_26692,N_25264,N_25300);
xor U26693 (N_26693,N_25357,N_25120);
and U26694 (N_26694,N_25250,N_25404);
nor U26695 (N_26695,N_24353,N_24631);
nand U26696 (N_26696,N_24716,N_24498);
or U26697 (N_26697,N_24083,N_24837);
nor U26698 (N_26698,N_24123,N_24346);
nand U26699 (N_26699,N_25305,N_24416);
nand U26700 (N_26700,N_24267,N_24854);
nand U26701 (N_26701,N_24942,N_24248);
xor U26702 (N_26702,N_24004,N_24569);
xnor U26703 (N_26703,N_24626,N_25160);
or U26704 (N_26704,N_25202,N_25119);
nand U26705 (N_26705,N_24319,N_24159);
or U26706 (N_26706,N_24893,N_25354);
xnor U26707 (N_26707,N_25202,N_25126);
nor U26708 (N_26708,N_25141,N_24126);
nor U26709 (N_26709,N_25161,N_25095);
and U26710 (N_26710,N_24558,N_24100);
or U26711 (N_26711,N_25402,N_24809);
or U26712 (N_26712,N_24333,N_24157);
nand U26713 (N_26713,N_25440,N_24704);
nor U26714 (N_26714,N_25114,N_24159);
or U26715 (N_26715,N_24410,N_25167);
nand U26716 (N_26716,N_24460,N_24814);
xor U26717 (N_26717,N_25291,N_25468);
nor U26718 (N_26718,N_25435,N_25009);
and U26719 (N_26719,N_25248,N_24701);
nor U26720 (N_26720,N_25169,N_25172);
and U26721 (N_26721,N_24661,N_24368);
nand U26722 (N_26722,N_25055,N_24180);
xnor U26723 (N_26723,N_24143,N_24377);
nor U26724 (N_26724,N_24159,N_24120);
nor U26725 (N_26725,N_25132,N_24303);
or U26726 (N_26726,N_25323,N_24397);
or U26727 (N_26727,N_24022,N_24574);
or U26728 (N_26728,N_24766,N_24400);
xor U26729 (N_26729,N_25081,N_24131);
nor U26730 (N_26730,N_24689,N_24918);
nand U26731 (N_26731,N_24134,N_24706);
xnor U26732 (N_26732,N_24966,N_25078);
nand U26733 (N_26733,N_25282,N_24777);
or U26734 (N_26734,N_24381,N_25048);
xor U26735 (N_26735,N_25004,N_24325);
or U26736 (N_26736,N_24619,N_24376);
and U26737 (N_26737,N_24781,N_25432);
xor U26738 (N_26738,N_24240,N_25372);
and U26739 (N_26739,N_24020,N_24914);
xnor U26740 (N_26740,N_24341,N_25407);
nand U26741 (N_26741,N_25329,N_24459);
nor U26742 (N_26742,N_24797,N_24499);
and U26743 (N_26743,N_25250,N_25082);
nor U26744 (N_26744,N_25213,N_24419);
or U26745 (N_26745,N_24017,N_24795);
nor U26746 (N_26746,N_24330,N_25411);
or U26747 (N_26747,N_24198,N_25116);
or U26748 (N_26748,N_24684,N_24561);
and U26749 (N_26749,N_25201,N_24072);
and U26750 (N_26750,N_24596,N_24989);
xor U26751 (N_26751,N_25269,N_24925);
nor U26752 (N_26752,N_24586,N_24563);
nor U26753 (N_26753,N_25279,N_24470);
or U26754 (N_26754,N_24722,N_24412);
or U26755 (N_26755,N_24492,N_25288);
nand U26756 (N_26756,N_25047,N_24724);
or U26757 (N_26757,N_24727,N_25189);
nor U26758 (N_26758,N_25312,N_24961);
nor U26759 (N_26759,N_24049,N_24746);
nor U26760 (N_26760,N_24934,N_25156);
xor U26761 (N_26761,N_25117,N_25336);
xnor U26762 (N_26762,N_25278,N_24653);
or U26763 (N_26763,N_25178,N_25154);
nand U26764 (N_26764,N_24672,N_24065);
xnor U26765 (N_26765,N_24433,N_24711);
or U26766 (N_26766,N_24537,N_25404);
xnor U26767 (N_26767,N_25270,N_25137);
xor U26768 (N_26768,N_24101,N_24845);
or U26769 (N_26769,N_24807,N_25249);
nor U26770 (N_26770,N_24921,N_24822);
nand U26771 (N_26771,N_24498,N_24740);
xor U26772 (N_26772,N_24674,N_25460);
or U26773 (N_26773,N_25166,N_24482);
nor U26774 (N_26774,N_25359,N_25398);
nor U26775 (N_26775,N_25455,N_24784);
nand U26776 (N_26776,N_24863,N_25281);
and U26777 (N_26777,N_25462,N_24646);
xor U26778 (N_26778,N_25046,N_25128);
and U26779 (N_26779,N_25298,N_24326);
xor U26780 (N_26780,N_25006,N_24473);
xor U26781 (N_26781,N_24101,N_25419);
nand U26782 (N_26782,N_24325,N_25474);
nand U26783 (N_26783,N_24954,N_24600);
and U26784 (N_26784,N_24947,N_24397);
nand U26785 (N_26785,N_25184,N_25253);
nor U26786 (N_26786,N_24252,N_24659);
or U26787 (N_26787,N_24900,N_24517);
nand U26788 (N_26788,N_25044,N_25169);
or U26789 (N_26789,N_25089,N_24626);
or U26790 (N_26790,N_25192,N_24880);
and U26791 (N_26791,N_24339,N_24678);
xor U26792 (N_26792,N_24182,N_24144);
and U26793 (N_26793,N_24133,N_24759);
and U26794 (N_26794,N_24191,N_25450);
or U26795 (N_26795,N_25429,N_24292);
or U26796 (N_26796,N_25489,N_24724);
xor U26797 (N_26797,N_24278,N_25343);
xor U26798 (N_26798,N_25004,N_24389);
and U26799 (N_26799,N_25348,N_25079);
nor U26800 (N_26800,N_24583,N_25438);
or U26801 (N_26801,N_24196,N_24142);
or U26802 (N_26802,N_24418,N_24077);
and U26803 (N_26803,N_25263,N_25227);
or U26804 (N_26804,N_24877,N_24769);
nand U26805 (N_26805,N_24383,N_24164);
nor U26806 (N_26806,N_24685,N_24187);
nor U26807 (N_26807,N_25010,N_24845);
nor U26808 (N_26808,N_24269,N_24415);
nor U26809 (N_26809,N_24635,N_25477);
nor U26810 (N_26810,N_24486,N_25248);
xor U26811 (N_26811,N_24287,N_25445);
nor U26812 (N_26812,N_24751,N_24441);
and U26813 (N_26813,N_24451,N_24587);
or U26814 (N_26814,N_24857,N_24146);
and U26815 (N_26815,N_24309,N_25321);
xor U26816 (N_26816,N_24702,N_25070);
xor U26817 (N_26817,N_25154,N_24963);
or U26818 (N_26818,N_25207,N_25456);
xor U26819 (N_26819,N_24540,N_24230);
nand U26820 (N_26820,N_24882,N_24930);
and U26821 (N_26821,N_24469,N_24969);
and U26822 (N_26822,N_25136,N_24318);
nor U26823 (N_26823,N_25167,N_25099);
or U26824 (N_26824,N_24307,N_24772);
xnor U26825 (N_26825,N_24505,N_24393);
nor U26826 (N_26826,N_25098,N_24068);
nor U26827 (N_26827,N_24882,N_24380);
nor U26828 (N_26828,N_24197,N_24955);
nand U26829 (N_26829,N_25262,N_25331);
nor U26830 (N_26830,N_24200,N_24672);
xnor U26831 (N_26831,N_25345,N_24431);
xnor U26832 (N_26832,N_25093,N_24913);
or U26833 (N_26833,N_24477,N_25194);
nor U26834 (N_26834,N_24243,N_25389);
xor U26835 (N_26835,N_24344,N_25416);
nor U26836 (N_26836,N_24886,N_25425);
or U26837 (N_26837,N_24567,N_25188);
nand U26838 (N_26838,N_25231,N_24090);
xnor U26839 (N_26839,N_25026,N_24566);
or U26840 (N_26840,N_24285,N_24797);
xor U26841 (N_26841,N_25054,N_24577);
and U26842 (N_26842,N_25103,N_24138);
nand U26843 (N_26843,N_25113,N_24675);
xor U26844 (N_26844,N_25467,N_25139);
nor U26845 (N_26845,N_24134,N_25034);
xnor U26846 (N_26846,N_25185,N_24852);
nand U26847 (N_26847,N_25139,N_24592);
xnor U26848 (N_26848,N_24026,N_24577);
or U26849 (N_26849,N_25001,N_24020);
or U26850 (N_26850,N_25179,N_25167);
or U26851 (N_26851,N_24370,N_24638);
or U26852 (N_26852,N_25088,N_24743);
and U26853 (N_26853,N_24647,N_25281);
xor U26854 (N_26854,N_24100,N_25357);
and U26855 (N_26855,N_25167,N_24016);
nand U26856 (N_26856,N_24375,N_24077);
xnor U26857 (N_26857,N_24001,N_24323);
xnor U26858 (N_26858,N_24903,N_24151);
nand U26859 (N_26859,N_25232,N_25380);
nor U26860 (N_26860,N_24560,N_24940);
and U26861 (N_26861,N_24424,N_25356);
xnor U26862 (N_26862,N_25111,N_24848);
and U26863 (N_26863,N_24050,N_25493);
xnor U26864 (N_26864,N_25176,N_24745);
nand U26865 (N_26865,N_24893,N_25002);
and U26866 (N_26866,N_24131,N_24446);
nand U26867 (N_26867,N_24787,N_25403);
nor U26868 (N_26868,N_24560,N_25427);
or U26869 (N_26869,N_25175,N_24503);
or U26870 (N_26870,N_24072,N_24772);
or U26871 (N_26871,N_25360,N_24858);
or U26872 (N_26872,N_25182,N_24770);
and U26873 (N_26873,N_24984,N_24271);
nor U26874 (N_26874,N_24004,N_24010);
nand U26875 (N_26875,N_25456,N_24058);
and U26876 (N_26876,N_24546,N_24345);
xnor U26877 (N_26877,N_24891,N_25234);
nor U26878 (N_26878,N_25323,N_25132);
and U26879 (N_26879,N_25325,N_24952);
or U26880 (N_26880,N_24586,N_24374);
nand U26881 (N_26881,N_25311,N_25416);
and U26882 (N_26882,N_25442,N_24114);
and U26883 (N_26883,N_24766,N_25340);
and U26884 (N_26884,N_24618,N_24046);
or U26885 (N_26885,N_24866,N_24838);
or U26886 (N_26886,N_24576,N_25102);
and U26887 (N_26887,N_24937,N_24383);
or U26888 (N_26888,N_24489,N_24794);
and U26889 (N_26889,N_25007,N_24155);
or U26890 (N_26890,N_25299,N_24326);
and U26891 (N_26891,N_25104,N_24874);
and U26892 (N_26892,N_24274,N_25438);
nor U26893 (N_26893,N_25380,N_24446);
and U26894 (N_26894,N_25280,N_24118);
xor U26895 (N_26895,N_24491,N_24786);
nand U26896 (N_26896,N_25432,N_25221);
and U26897 (N_26897,N_24824,N_25188);
xnor U26898 (N_26898,N_25048,N_24931);
or U26899 (N_26899,N_24529,N_24249);
nor U26900 (N_26900,N_24983,N_24170);
and U26901 (N_26901,N_24138,N_24542);
or U26902 (N_26902,N_25051,N_24365);
and U26903 (N_26903,N_24096,N_24333);
and U26904 (N_26904,N_24416,N_24770);
nand U26905 (N_26905,N_24337,N_25495);
xor U26906 (N_26906,N_24394,N_25027);
nor U26907 (N_26907,N_25385,N_24470);
nor U26908 (N_26908,N_25016,N_24605);
nor U26909 (N_26909,N_24183,N_24368);
or U26910 (N_26910,N_24489,N_25029);
and U26911 (N_26911,N_25401,N_24106);
xnor U26912 (N_26912,N_24290,N_24722);
nor U26913 (N_26913,N_24095,N_24892);
nand U26914 (N_26914,N_24582,N_25110);
nand U26915 (N_26915,N_24219,N_24628);
xor U26916 (N_26916,N_24350,N_24866);
or U26917 (N_26917,N_25027,N_24037);
xor U26918 (N_26918,N_24845,N_24087);
nor U26919 (N_26919,N_25040,N_24632);
or U26920 (N_26920,N_24778,N_25025);
nor U26921 (N_26921,N_24082,N_24113);
and U26922 (N_26922,N_24454,N_25387);
or U26923 (N_26923,N_24163,N_24464);
or U26924 (N_26924,N_24169,N_24368);
xor U26925 (N_26925,N_25006,N_24404);
nand U26926 (N_26926,N_24499,N_24176);
nor U26927 (N_26927,N_24181,N_25477);
xor U26928 (N_26928,N_24577,N_24673);
or U26929 (N_26929,N_25453,N_24631);
xnor U26930 (N_26930,N_24702,N_24647);
xnor U26931 (N_26931,N_24753,N_24088);
nor U26932 (N_26932,N_24912,N_24771);
or U26933 (N_26933,N_25164,N_24283);
nor U26934 (N_26934,N_25178,N_24575);
nand U26935 (N_26935,N_24207,N_24830);
xor U26936 (N_26936,N_25214,N_24129);
nand U26937 (N_26937,N_24220,N_25196);
nand U26938 (N_26938,N_25149,N_25292);
nand U26939 (N_26939,N_25001,N_24501);
or U26940 (N_26940,N_25304,N_24237);
nor U26941 (N_26941,N_24371,N_25038);
or U26942 (N_26942,N_24481,N_24730);
and U26943 (N_26943,N_25143,N_25044);
or U26944 (N_26944,N_24082,N_24816);
xnor U26945 (N_26945,N_24496,N_24139);
or U26946 (N_26946,N_24104,N_24614);
nand U26947 (N_26947,N_24169,N_24921);
or U26948 (N_26948,N_24312,N_25300);
nand U26949 (N_26949,N_24025,N_24860);
and U26950 (N_26950,N_24603,N_24989);
nand U26951 (N_26951,N_24353,N_24997);
or U26952 (N_26952,N_24018,N_24594);
and U26953 (N_26953,N_24188,N_24324);
nor U26954 (N_26954,N_24013,N_24898);
nor U26955 (N_26955,N_24231,N_25068);
or U26956 (N_26956,N_25388,N_24740);
nand U26957 (N_26957,N_24170,N_25120);
nand U26958 (N_26958,N_25206,N_24612);
or U26959 (N_26959,N_24513,N_24560);
or U26960 (N_26960,N_24579,N_24979);
nor U26961 (N_26961,N_24098,N_24543);
and U26962 (N_26962,N_24055,N_24255);
and U26963 (N_26963,N_24140,N_25206);
or U26964 (N_26964,N_25043,N_25432);
or U26965 (N_26965,N_24771,N_24901);
xnor U26966 (N_26966,N_25366,N_25367);
xor U26967 (N_26967,N_24929,N_25038);
or U26968 (N_26968,N_24334,N_25132);
nor U26969 (N_26969,N_24786,N_24372);
nand U26970 (N_26970,N_24057,N_24234);
xnor U26971 (N_26971,N_24222,N_24429);
nor U26972 (N_26972,N_24242,N_24891);
xor U26973 (N_26973,N_24747,N_24641);
xor U26974 (N_26974,N_24645,N_24914);
or U26975 (N_26975,N_25458,N_25208);
nor U26976 (N_26976,N_24055,N_25496);
and U26977 (N_26977,N_25322,N_24970);
and U26978 (N_26978,N_24782,N_24648);
and U26979 (N_26979,N_24227,N_25210);
nand U26980 (N_26980,N_24999,N_24475);
or U26981 (N_26981,N_24715,N_24673);
and U26982 (N_26982,N_24472,N_24662);
nor U26983 (N_26983,N_25279,N_25074);
xnor U26984 (N_26984,N_24416,N_24226);
nand U26985 (N_26985,N_25151,N_24152);
or U26986 (N_26986,N_24200,N_24289);
or U26987 (N_26987,N_24180,N_24720);
nor U26988 (N_26988,N_24530,N_24154);
xnor U26989 (N_26989,N_24292,N_25162);
nand U26990 (N_26990,N_24486,N_25463);
nand U26991 (N_26991,N_24522,N_24576);
xor U26992 (N_26992,N_25381,N_24904);
nand U26993 (N_26993,N_25194,N_24599);
or U26994 (N_26994,N_24018,N_24575);
nor U26995 (N_26995,N_24805,N_25344);
xnor U26996 (N_26996,N_24957,N_24445);
and U26997 (N_26997,N_25231,N_24752);
and U26998 (N_26998,N_24858,N_24469);
xor U26999 (N_26999,N_25168,N_24715);
or U27000 (N_27000,N_26963,N_26100);
xnor U27001 (N_27001,N_25925,N_25544);
nand U27002 (N_27002,N_25876,N_26610);
and U27003 (N_27003,N_25611,N_26482);
nor U27004 (N_27004,N_25549,N_26242);
or U27005 (N_27005,N_26052,N_26089);
nand U27006 (N_27006,N_25923,N_25635);
nor U27007 (N_27007,N_25542,N_26976);
nand U27008 (N_27008,N_26200,N_26399);
xnor U27009 (N_27009,N_26601,N_25566);
nand U27010 (N_27010,N_26166,N_25939);
and U27011 (N_27011,N_26552,N_26984);
xnor U27012 (N_27012,N_26004,N_26165);
nor U27013 (N_27013,N_26347,N_25832);
and U27014 (N_27014,N_25772,N_26544);
or U27015 (N_27015,N_26603,N_25856);
and U27016 (N_27016,N_26338,N_25732);
xor U27017 (N_27017,N_25979,N_26343);
nor U27018 (N_27018,N_26651,N_26401);
nor U27019 (N_27019,N_26434,N_26251);
and U27020 (N_27020,N_26782,N_25752);
xnor U27021 (N_27021,N_26537,N_25580);
and U27022 (N_27022,N_26138,N_26076);
and U27023 (N_27023,N_26890,N_25516);
and U27024 (N_27024,N_26915,N_26659);
nor U27025 (N_27025,N_26028,N_26216);
and U27026 (N_27026,N_26406,N_26459);
and U27027 (N_27027,N_26771,N_26940);
and U27028 (N_27028,N_25731,N_26201);
or U27029 (N_27029,N_26314,N_25588);
or U27030 (N_27030,N_26041,N_25656);
xnor U27031 (N_27031,N_25593,N_25933);
and U27032 (N_27032,N_26921,N_26602);
nand U27033 (N_27033,N_26996,N_25884);
xor U27034 (N_27034,N_26789,N_26077);
nand U27035 (N_27035,N_25543,N_25576);
xnor U27036 (N_27036,N_26545,N_26755);
xnor U27037 (N_27037,N_25907,N_26954);
xor U27038 (N_27038,N_26566,N_26647);
nand U27039 (N_27039,N_26672,N_25946);
and U27040 (N_27040,N_26907,N_26247);
or U27041 (N_27041,N_25625,N_26970);
nor U27042 (N_27042,N_25938,N_26860);
or U27043 (N_27043,N_25717,N_25538);
or U27044 (N_27044,N_26148,N_25640);
or U27045 (N_27045,N_26222,N_26763);
xor U27046 (N_27046,N_26390,N_26037);
xor U27047 (N_27047,N_26155,N_25880);
or U27048 (N_27048,N_26597,N_26709);
or U27049 (N_27049,N_26561,N_26742);
xor U27050 (N_27050,N_26820,N_26839);
nand U27051 (N_27051,N_26126,N_26885);
nand U27052 (N_27052,N_26371,N_25613);
or U27053 (N_27053,N_26520,N_25646);
nor U27054 (N_27054,N_26420,N_25626);
nand U27055 (N_27055,N_25535,N_25776);
xnor U27056 (N_27056,N_25614,N_26008);
and U27057 (N_27057,N_25711,N_26623);
or U27058 (N_27058,N_26931,N_26236);
nor U27059 (N_27059,N_26365,N_25788);
or U27060 (N_27060,N_25879,N_25537);
nor U27061 (N_27061,N_25757,N_26481);
nand U27062 (N_27062,N_26643,N_26728);
or U27063 (N_27063,N_26701,N_26558);
xor U27064 (N_27064,N_26240,N_26262);
or U27065 (N_27065,N_25749,N_26075);
xor U27066 (N_27066,N_25651,N_26319);
xor U27067 (N_27067,N_25826,N_26124);
nand U27068 (N_27068,N_26211,N_26475);
nor U27069 (N_27069,N_26436,N_26140);
and U27070 (N_27070,N_26440,N_25913);
nand U27071 (N_27071,N_25501,N_26744);
nor U27072 (N_27072,N_25784,N_25709);
or U27073 (N_27073,N_25951,N_25663);
nor U27074 (N_27074,N_26062,N_26683);
nand U27075 (N_27075,N_26161,N_26500);
or U27076 (N_27076,N_25999,N_26111);
nor U27077 (N_27077,N_26467,N_26916);
nand U27078 (N_27078,N_25968,N_26613);
nor U27079 (N_27079,N_25994,N_26769);
nor U27080 (N_27080,N_25674,N_26451);
nor U27081 (N_27081,N_26241,N_26776);
nand U27082 (N_27082,N_26082,N_26445);
xnor U27083 (N_27083,N_26619,N_26836);
or U27084 (N_27084,N_26108,N_26293);
or U27085 (N_27085,N_26288,N_26644);
nand U27086 (N_27086,N_26780,N_26405);
nand U27087 (N_27087,N_26282,N_26430);
and U27088 (N_27088,N_25688,N_25834);
and U27089 (N_27089,N_25668,N_25860);
and U27090 (N_27090,N_26562,N_26478);
nor U27091 (N_27091,N_26362,N_25980);
nand U27092 (N_27092,N_26435,N_26305);
and U27093 (N_27093,N_25893,N_26326);
nor U27094 (N_27094,N_25713,N_26524);
and U27095 (N_27095,N_25703,N_26749);
nand U27096 (N_27096,N_26766,N_25574);
and U27097 (N_27097,N_26998,N_26083);
and U27098 (N_27098,N_26779,N_26381);
nand U27099 (N_27099,N_26874,N_25734);
nand U27100 (N_27100,N_26715,N_26638);
and U27101 (N_27101,N_26005,N_26385);
and U27102 (N_27102,N_26533,N_26384);
or U27103 (N_27103,N_26181,N_26360);
nor U27104 (N_27104,N_26980,N_26630);
xnor U27105 (N_27105,N_26534,N_25728);
nor U27106 (N_27106,N_25707,N_25741);
nand U27107 (N_27107,N_25724,N_26375);
or U27108 (N_27108,N_26723,N_26580);
nand U27109 (N_27109,N_26631,N_26180);
and U27110 (N_27110,N_26859,N_26007);
or U27111 (N_27111,N_25624,N_26272);
and U27112 (N_27112,N_25871,N_26967);
or U27113 (N_27113,N_25889,N_25875);
and U27114 (N_27114,N_25557,N_26993);
or U27115 (N_27115,N_26814,N_26276);
and U27116 (N_27116,N_26712,N_25921);
or U27117 (N_27117,N_25899,N_25563);
and U27118 (N_27118,N_26882,N_26622);
xnor U27119 (N_27119,N_25807,N_26373);
and U27120 (N_27120,N_25781,N_26509);
nand U27121 (N_27121,N_26513,N_26256);
nor U27122 (N_27122,N_25903,N_25519);
xor U27123 (N_27123,N_25866,N_26285);
and U27124 (N_27124,N_25607,N_26495);
or U27125 (N_27125,N_26527,N_26308);
or U27126 (N_27126,N_25528,N_26210);
and U27127 (N_27127,N_26324,N_26258);
or U27128 (N_27128,N_25701,N_26017);
and U27129 (N_27129,N_26514,N_26551);
nand U27130 (N_27130,N_26183,N_25722);
or U27131 (N_27131,N_25521,N_26118);
nor U27132 (N_27132,N_25920,N_25919);
xor U27133 (N_27133,N_26668,N_26189);
xnor U27134 (N_27134,N_26426,N_25988);
and U27135 (N_27135,N_26686,N_26521);
and U27136 (N_27136,N_26639,N_25673);
nand U27137 (N_27137,N_26920,N_26398);
nand U27138 (N_27138,N_25689,N_26454);
and U27139 (N_27139,N_25966,N_26307);
and U27140 (N_27140,N_26173,N_26429);
nand U27141 (N_27141,N_26304,N_26303);
or U27142 (N_27142,N_26460,N_25993);
xor U27143 (N_27143,N_26112,N_26031);
nor U27144 (N_27144,N_25808,N_26227);
nor U27145 (N_27145,N_25755,N_26059);
nor U27146 (N_27146,N_25585,N_26508);
nor U27147 (N_27147,N_25801,N_26707);
and U27148 (N_27148,N_26156,N_26595);
nand U27149 (N_27149,N_26797,N_26986);
or U27150 (N_27150,N_26832,N_26673);
or U27151 (N_27151,N_26355,N_25839);
nand U27152 (N_27152,N_25975,N_26556);
and U27153 (N_27153,N_26829,N_26841);
nand U27154 (N_27154,N_26669,N_25770);
nand U27155 (N_27155,N_26854,N_25702);
and U27156 (N_27156,N_25733,N_25705);
or U27157 (N_27157,N_26144,N_25685);
and U27158 (N_27158,N_26670,N_26067);
xnor U27159 (N_27159,N_25971,N_26234);
xnor U27160 (N_27160,N_26648,N_25594);
nor U27161 (N_27161,N_26952,N_25981);
nor U27162 (N_27162,N_25553,N_25854);
and U27163 (N_27163,N_26748,N_25989);
nand U27164 (N_27164,N_26574,N_25756);
and U27165 (N_27165,N_25865,N_26588);
nand U27166 (N_27166,N_26042,N_25642);
and U27167 (N_27167,N_25987,N_26237);
nand U27168 (N_27168,N_26080,N_26584);
or U27169 (N_27169,N_26257,N_26851);
and U27170 (N_27170,N_25887,N_26006);
or U27171 (N_27171,N_26152,N_26128);
nor U27172 (N_27172,N_26239,N_25530);
xnor U27173 (N_27173,N_25502,N_25882);
nand U27174 (N_27174,N_26248,N_25630);
xnor U27175 (N_27175,N_26097,N_25991);
nand U27176 (N_27176,N_26411,N_26160);
xor U27177 (N_27177,N_26287,N_26871);
or U27178 (N_27178,N_26805,N_25976);
nand U27179 (N_27179,N_26759,N_26127);
xnor U27180 (N_27180,N_26264,N_26895);
xor U27181 (N_27181,N_26966,N_26423);
xnor U27182 (N_27182,N_26999,N_25745);
xnor U27183 (N_27183,N_25598,N_26466);
xor U27184 (N_27184,N_26046,N_26635);
and U27185 (N_27185,N_26792,N_26054);
and U27186 (N_27186,N_25679,N_26091);
xnor U27187 (N_27187,N_26182,N_26765);
xnor U27188 (N_27188,N_26988,N_26229);
nand U27189 (N_27189,N_26117,N_26113);
nand U27190 (N_27190,N_25682,N_25600);
nand U27191 (N_27191,N_26098,N_26750);
nand U27192 (N_27192,N_26536,N_26599);
nor U27193 (N_27193,N_25568,N_26354);
nor U27194 (N_27194,N_25599,N_26717);
nor U27195 (N_27195,N_26051,N_25983);
and U27196 (N_27196,N_25896,N_25507);
xor U27197 (N_27197,N_26014,N_25890);
or U27198 (N_27198,N_26710,N_25931);
and U27199 (N_27199,N_25997,N_26863);
nand U27200 (N_27200,N_25855,N_25943);
nand U27201 (N_27201,N_26679,N_25824);
xor U27202 (N_27202,N_25918,N_26681);
nand U27203 (N_27203,N_25727,N_26965);
or U27204 (N_27204,N_25645,N_26719);
and U27205 (N_27205,N_26539,N_26106);
nor U27206 (N_27206,N_25506,N_26827);
nor U27207 (N_27207,N_26190,N_25671);
or U27208 (N_27208,N_25935,N_25877);
nor U27209 (N_27209,N_26981,N_26185);
and U27210 (N_27210,N_26045,N_26278);
nand U27211 (N_27211,N_25763,N_26884);
nor U27212 (N_27212,N_26188,N_26410);
or U27213 (N_27213,N_25909,N_26713);
or U27214 (N_27214,N_25730,N_26818);
or U27215 (N_27215,N_25691,N_25849);
and U27216 (N_27216,N_26629,N_26625);
nor U27217 (N_27217,N_25901,N_26852);
nand U27218 (N_27218,N_25708,N_25504);
xnor U27219 (N_27219,N_26228,N_26009);
and U27220 (N_27220,N_26102,N_26730);
xor U27221 (N_27221,N_25828,N_26957);
nor U27222 (N_27222,N_26893,N_25978);
nor U27223 (N_27223,N_26408,N_26615);
nor U27224 (N_27224,N_26081,N_25641);
nand U27225 (N_27225,N_26016,N_26912);
nand U27226 (N_27226,N_26186,N_25555);
nor U27227 (N_27227,N_26948,N_26243);
nor U27228 (N_27228,N_25868,N_26813);
and U27229 (N_27229,N_25500,N_26700);
and U27230 (N_27230,N_26026,N_25819);
or U27231 (N_27231,N_26364,N_26122);
or U27232 (N_27232,N_26589,N_25578);
xnor U27233 (N_27233,N_26132,N_26937);
nor U27234 (N_27234,N_26002,N_26058);
and U27235 (N_27235,N_25794,N_25934);
xor U27236 (N_27236,N_25726,N_25817);
xor U27237 (N_27237,N_25534,N_25508);
nor U27238 (N_27238,N_25517,N_25767);
nor U27239 (N_27239,N_25806,N_26995);
or U27240 (N_27240,N_26455,N_26951);
xor U27241 (N_27241,N_26933,N_25815);
or U27242 (N_27242,N_25622,N_25631);
xor U27243 (N_27243,N_26905,N_26409);
nor U27244 (N_27244,N_25798,N_26000);
and U27245 (N_27245,N_26032,N_25844);
or U27246 (N_27246,N_25541,N_25629);
nand U27247 (N_27247,N_26762,N_25869);
nor U27248 (N_27248,N_25522,N_26048);
or U27249 (N_27249,N_26259,N_26487);
xor U27250 (N_27250,N_26724,N_26400);
and U27251 (N_27251,N_26515,N_26439);
xor U27252 (N_27252,N_26845,N_25823);
xnor U27253 (N_27253,N_25571,N_25765);
nand U27254 (N_27254,N_26866,N_26528);
nand U27255 (N_27255,N_26560,N_26361);
nor U27256 (N_27256,N_26547,N_25782);
and U27257 (N_27257,N_26929,N_26801);
nand U27258 (N_27258,N_25954,N_25915);
nand U27259 (N_27259,N_26828,N_26575);
nor U27260 (N_27260,N_26943,N_26238);
or U27261 (N_27261,N_26857,N_26664);
xnor U27262 (N_27262,N_25892,N_25601);
and U27263 (N_27263,N_26891,N_25964);
xnor U27264 (N_27264,N_25766,N_25694);
nor U27265 (N_27265,N_26452,N_26538);
xnor U27266 (N_27266,N_25795,N_26346);
and U27267 (N_27267,N_26492,N_25654);
and U27268 (N_27268,N_26107,N_26889);
nor U27269 (N_27269,N_26203,N_25858);
xnor U27270 (N_27270,N_26213,N_26232);
or U27271 (N_27271,N_26868,N_26318);
nand U27272 (N_27272,N_26690,N_26583);
or U27273 (N_27273,N_26279,N_26947);
and U27274 (N_27274,N_25950,N_26894);
or U27275 (N_27275,N_26611,N_26987);
and U27276 (N_27276,N_25676,N_25917);
nor U27277 (N_27277,N_26869,N_26770);
xnor U27278 (N_27278,N_26019,N_25942);
nand U27279 (N_27279,N_26695,N_25972);
nor U27280 (N_27280,N_26888,N_26685);
nor U27281 (N_27281,N_26909,N_26516);
nand U27282 (N_27282,N_25829,N_26198);
nor U27283 (N_27283,N_25602,N_25783);
nor U27284 (N_27284,N_26865,N_26323);
or U27285 (N_27285,N_26864,N_25937);
nor U27286 (N_27286,N_25758,N_26675);
or U27287 (N_27287,N_25575,N_25720);
or U27288 (N_27288,N_26628,N_26233);
nor U27289 (N_27289,N_26437,N_26143);
xnor U27290 (N_27290,N_25998,N_26403);
xnor U27291 (N_27291,N_26153,N_26992);
nand U27292 (N_27292,N_26910,N_26254);
nand U27293 (N_27293,N_26585,N_26898);
or U27294 (N_27294,N_26975,N_26777);
or U27295 (N_27295,N_26641,N_26469);
xnor U27296 (N_27296,N_25761,N_25977);
nor U27297 (N_27297,N_25670,N_26844);
and U27298 (N_27298,N_26268,N_26853);
and U27299 (N_27299,N_26798,N_25905);
or U27300 (N_27300,N_26886,N_26908);
nand U27301 (N_27301,N_25827,N_26214);
nor U27302 (N_27302,N_26598,N_25505);
nand U27303 (N_27303,N_25878,N_26705);
or U27304 (N_27304,N_26919,N_26784);
or U27305 (N_27305,N_26812,N_26484);
xnor U27306 (N_27306,N_26079,N_26147);
or U27307 (N_27307,N_26191,N_26600);
nor U27308 (N_27308,N_25840,N_25650);
and U27309 (N_27309,N_25659,N_26465);
nor U27310 (N_27310,N_25963,N_26096);
or U27311 (N_27311,N_26689,N_26474);
nand U27312 (N_27312,N_26518,N_26427);
xnor U27313 (N_27313,N_25558,N_26997);
nor U27314 (N_27314,N_25714,N_25510);
nand U27315 (N_27315,N_26577,N_26275);
or U27316 (N_27316,N_26168,N_25531);
or U27317 (N_27317,N_26339,N_26468);
and U27318 (N_27318,N_26834,N_25984);
or U27319 (N_27319,N_25725,N_26476);
nand U27320 (N_27320,N_26969,N_25848);
xnor U27321 (N_27321,N_26274,N_25792);
nor U27322 (N_27322,N_26151,N_26830);
or U27323 (N_27323,N_26120,N_25872);
nor U27324 (N_27324,N_26542,N_26729);
nand U27325 (N_27325,N_26494,N_26105);
and U27326 (N_27326,N_26800,N_26913);
xor U27327 (N_27327,N_25657,N_26103);
xnor U27328 (N_27328,N_26815,N_26447);
or U27329 (N_27329,N_26959,N_26368);
nand U27330 (N_27330,N_26312,N_26511);
xnor U27331 (N_27331,N_26897,N_25660);
or U27332 (N_27332,N_26872,N_25723);
and U27333 (N_27333,N_26387,N_26367);
nor U27334 (N_27334,N_26345,N_25771);
xnor U27335 (N_27335,N_26855,N_26325);
xnor U27336 (N_27336,N_26650,N_25664);
nand U27337 (N_27337,N_26657,N_25697);
nand U27338 (N_27338,N_26530,N_26711);
and U27339 (N_27339,N_26444,N_26283);
xor U27340 (N_27340,N_25655,N_26676);
and U27341 (N_27341,N_26123,N_25825);
or U27342 (N_27342,N_26350,N_26892);
or U27343 (N_27343,N_26193,N_26896);
nor U27344 (N_27344,N_25560,N_25683);
nor U27345 (N_27345,N_26022,N_26703);
nand U27346 (N_27346,N_26737,N_26687);
and U27347 (N_27347,N_26280,N_26039);
nor U27348 (N_27348,N_26902,N_26768);
and U27349 (N_27349,N_26417,N_26121);
nor U27350 (N_27350,N_25739,N_25562);
xor U27351 (N_27351,N_25748,N_26066);
and U27352 (N_27352,N_26490,N_26374);
and U27353 (N_27353,N_25898,N_25852);
or U27354 (N_27354,N_25649,N_25559);
nand U27355 (N_27355,N_26734,N_26134);
or U27356 (N_27356,N_26671,N_26219);
nand U27357 (N_27357,N_26225,N_25718);
or U27358 (N_27358,N_26740,N_25527);
xor U27359 (N_27359,N_26491,N_26418);
nand U27360 (N_27360,N_25857,N_26245);
and U27361 (N_27361,N_26738,N_26088);
and U27362 (N_27362,N_26714,N_26942);
or U27363 (N_27363,N_26732,N_26104);
xor U27364 (N_27364,N_25678,N_26479);
xnor U27365 (N_27365,N_26821,N_26197);
or U27366 (N_27366,N_26950,N_26473);
nand U27367 (N_27367,N_25681,N_26694);
and U27368 (N_27368,N_26754,N_25965);
nor U27369 (N_27369,N_26056,N_26573);
or U27370 (N_27370,N_25513,N_25803);
nor U27371 (N_27371,N_26962,N_25514);
nor U27372 (N_27372,N_26785,N_25961);
nand U27373 (N_27373,N_26172,N_25751);
nand U27374 (N_27374,N_26392,N_26773);
and U27375 (N_27375,N_25584,N_26271);
and U27376 (N_27376,N_26502,N_26835);
and U27377 (N_27377,N_26043,N_26377);
or U27378 (N_27378,N_25744,N_26290);
nand U27379 (N_27379,N_26110,N_25740);
and U27380 (N_27380,N_25610,N_26716);
or U27381 (N_27381,N_26162,N_25836);
or U27382 (N_27382,N_26559,N_26837);
or U27383 (N_27383,N_25864,N_26425);
nand U27384 (N_27384,N_26372,N_25692);
nor U27385 (N_27385,N_26555,N_26125);
and U27386 (N_27386,N_26337,N_25632);
xnor U27387 (N_27387,N_26572,N_26115);
xor U27388 (N_27388,N_26204,N_26208);
and U27389 (N_27389,N_26317,N_26464);
or U27390 (N_27390,N_25552,N_26072);
or U27391 (N_27391,N_26010,N_25786);
nand U27392 (N_27392,N_25570,N_26071);
or U27393 (N_27393,N_25551,N_25719);
xor U27394 (N_27394,N_26861,N_26003);
and U27395 (N_27395,N_25797,N_25567);
xnor U27396 (N_27396,N_25672,N_26012);
nor U27397 (N_27397,N_25617,N_25911);
or U27398 (N_27398,N_26217,N_26667);
nand U27399 (N_27399,N_25830,N_26911);
and U27400 (N_27400,N_25843,N_26994);
nand U27401 (N_27401,N_25842,N_26205);
xor U27402 (N_27402,N_26590,N_26366);
and U27403 (N_27403,N_25737,N_26548);
xnor U27404 (N_27404,N_25564,N_26549);
nor U27405 (N_27405,N_26068,N_25870);
xor U27406 (N_27406,N_26973,N_25986);
nor U27407 (N_27407,N_26634,N_26564);
nor U27408 (N_27408,N_26906,N_26541);
nand U27409 (N_27409,N_26457,N_26531);
and U27410 (N_27410,N_26523,N_26421);
and U27411 (N_27411,N_26215,N_26141);
xnor U27412 (N_27412,N_25738,N_26774);
and U27413 (N_27413,N_26621,N_25813);
nand U27414 (N_27414,N_26579,N_26655);
nor U27415 (N_27415,N_26055,N_26231);
nand U27416 (N_27416,N_26876,N_25837);
or U27417 (N_27417,N_25603,N_25810);
xor U27418 (N_27418,N_26824,N_26982);
or U27419 (N_27419,N_25928,N_25637);
xor U27420 (N_27420,N_26535,N_26431);
and U27421 (N_27421,N_26945,N_26593);
nand U27422 (N_27422,N_26114,N_26939);
or U27423 (N_27423,N_26396,N_25586);
xnor U27424 (N_27424,N_26620,N_26788);
nand U27425 (N_27425,N_26529,N_26718);
nand U27426 (N_27426,N_26727,N_25773);
nand U27427 (N_27427,N_26154,N_25990);
nand U27428 (N_27428,N_25944,N_26674);
and U27429 (N_27429,N_26692,N_26253);
nor U27430 (N_27430,N_26171,N_26934);
or U27431 (N_27431,N_26024,N_26653);
nor U27432 (N_27432,N_26809,N_26316);
and U27433 (N_27433,N_26781,N_25960);
and U27434 (N_27434,N_25785,N_25680);
nor U27435 (N_27435,N_26512,N_25509);
nand U27436 (N_27436,N_25675,N_25862);
xor U27437 (N_27437,N_25729,N_25569);
nand U27438 (N_27438,N_25596,N_25577);
or U27439 (N_27439,N_25644,N_25546);
or U27440 (N_27440,N_25759,N_26199);
nor U27441 (N_27441,N_26532,N_26310);
nor U27442 (N_27442,N_25891,N_25547);
nand U27443 (N_27443,N_25846,N_25885);
or U27444 (N_27444,N_26764,N_26488);
nor U27445 (N_27445,N_25554,N_25859);
xnor U27446 (N_27446,N_26023,N_26637);
nand U27447 (N_27447,N_26791,N_26030);
xnor U27448 (N_27448,N_26443,N_26918);
xor U27449 (N_27449,N_25912,N_26783);
or U27450 (N_27450,N_26311,N_26879);
nor U27451 (N_27451,N_25606,N_26823);
nor U27452 (N_27452,N_26044,N_26313);
nand U27453 (N_27453,N_26831,N_25929);
or U27454 (N_27454,N_26930,N_26594);
or U27455 (N_27455,N_26989,N_26745);
xnor U27456 (N_27456,N_25589,N_25687);
and U27457 (N_27457,N_26470,N_26221);
nor U27458 (N_27458,N_26230,N_26158);
or U27459 (N_27459,N_26665,N_26568);
nor U27460 (N_27460,N_26099,N_26049);
and U27461 (N_27461,N_25747,N_26794);
or U27462 (N_27462,N_26116,N_26862);
nor U27463 (N_27463,N_26289,N_26654);
nand U27464 (N_27464,N_25618,N_26553);
nand U27465 (N_27465,N_25900,N_26069);
nor U27466 (N_27466,N_26270,N_26402);
xnor U27467 (N_27467,N_26142,N_25550);
nand U27468 (N_27468,N_25814,N_26101);
and U27469 (N_27469,N_25746,N_26087);
or U27470 (N_27470,N_26772,N_26811);
xor U27471 (N_27471,N_26169,N_26543);
nand U27472 (N_27472,N_26129,N_26775);
and U27473 (N_27473,N_25721,N_25853);
xor U27474 (N_27474,N_26050,N_26358);
or U27475 (N_27475,N_26084,N_26136);
xnor U27476 (N_27476,N_26847,N_26618);
and U27477 (N_27477,N_26725,N_26015);
or U27478 (N_27478,N_26557,N_25924);
xor U27479 (N_27479,N_26904,N_26284);
xor U27480 (N_27480,N_26846,N_26684);
nand U27481 (N_27481,N_26922,N_26333);
nand U27482 (N_27482,N_26159,N_25973);
and U27483 (N_27483,N_26064,N_26187);
nor U27484 (N_27484,N_26582,N_25936);
or U27485 (N_27485,N_25503,N_26842);
nor U27486 (N_27486,N_25953,N_26642);
nor U27487 (N_27487,N_25804,N_26021);
xnor U27488 (N_27488,N_26025,N_25619);
and U27489 (N_27489,N_25662,N_25690);
nand U27490 (N_27490,N_26501,N_26720);
or U27491 (N_27491,N_26395,N_25962);
nand U27492 (N_27492,N_25916,N_25666);
or U27493 (N_27493,N_26799,N_25532);
nor U27494 (N_27494,N_26320,N_25536);
and U27495 (N_27495,N_26721,N_26013);
or U27496 (N_27496,N_25886,N_26449);
xor U27497 (N_27497,N_25582,N_26504);
or U27498 (N_27498,N_26806,N_26540);
and U27499 (N_27499,N_26985,N_25902);
nand U27500 (N_27500,N_26422,N_25595);
or U27501 (N_27501,N_25874,N_26065);
and U27502 (N_27502,N_26804,N_26438);
or U27503 (N_27503,N_26696,N_25573);
xor U27504 (N_27504,N_25956,N_26038);
xor U27505 (N_27505,N_26751,N_26070);
xor U27506 (N_27506,N_26269,N_26493);
xnor U27507 (N_27507,N_26903,N_25699);
xor U27508 (N_27508,N_26899,N_26586);
or U27509 (N_27509,N_26736,N_26708);
nand U27510 (N_27510,N_26753,N_26605);
xnor U27511 (N_27511,N_26472,N_26757);
xnor U27512 (N_27512,N_26875,N_25684);
and U27513 (N_27513,N_26961,N_25750);
and U27514 (N_27514,N_26164,N_25957);
or U27515 (N_27515,N_26291,N_26587);
or U27516 (N_27516,N_26932,N_26607);
nand U27517 (N_27517,N_26453,N_25812);
xor U27518 (N_27518,N_26526,N_26137);
nor U27519 (N_27519,N_25805,N_26483);
and U27520 (N_27520,N_25789,N_25958);
or U27521 (N_27521,N_25914,N_26131);
xnor U27522 (N_27522,N_26645,N_26149);
nor U27523 (N_27523,N_25940,N_26565);
nand U27524 (N_27524,N_26739,N_25906);
nand U27525 (N_27525,N_26498,N_25948);
nand U27526 (N_27526,N_26887,N_25620);
and U27527 (N_27527,N_26063,N_26295);
and U27528 (N_27528,N_26609,N_26353);
nand U27529 (N_27529,N_26315,N_26485);
nand U27530 (N_27530,N_25974,N_25816);
xor U27531 (N_27531,N_26878,N_26499);
or U27532 (N_27532,N_26649,N_25910);
nand U27533 (N_27533,N_26192,N_26133);
or U27534 (N_27534,N_26036,N_25677);
nand U27535 (N_27535,N_26095,N_26196);
or U27536 (N_27536,N_26505,N_25811);
nand U27537 (N_27537,N_25628,N_26035);
nand U27538 (N_27538,N_26458,N_26414);
or U27539 (N_27539,N_26581,N_25658);
nand U27540 (N_27540,N_26462,N_25565);
nand U27541 (N_27541,N_26935,N_26020);
or U27542 (N_27542,N_25818,N_25820);
xnor U27543 (N_27543,N_26344,N_26522);
xor U27544 (N_27544,N_26486,N_25791);
or U27545 (N_27545,N_26255,N_26202);
and U27546 (N_27546,N_25511,N_26329);
nand U27547 (N_27547,N_26011,N_25590);
nor U27548 (N_27548,N_26349,N_26135);
and U27549 (N_27549,N_25932,N_26636);
and U27550 (N_27550,N_26456,N_25592);
or U27551 (N_27551,N_25608,N_26682);
or U27552 (N_27552,N_26061,N_26680);
nor U27553 (N_27553,N_26428,N_26612);
nand U27554 (N_27554,N_26880,N_25686);
or U27555 (N_27555,N_25512,N_26571);
and U27556 (N_27556,N_26407,N_26576);
or U27557 (N_27557,N_26001,N_25959);
xnor U27558 (N_27558,N_26244,N_26376);
xor U27559 (N_27559,N_26292,N_26273);
nand U27560 (N_27560,N_26808,N_26294);
xor U27561 (N_27561,N_26817,N_25985);
and U27562 (N_27562,N_26778,N_25612);
and U27563 (N_27563,N_26900,N_26109);
or U27564 (N_27564,N_26596,N_26209);
nor U27565 (N_27565,N_26163,N_26383);
xor U27566 (N_27566,N_25665,N_26397);
and U27567 (N_27567,N_26698,N_25735);
xor U27568 (N_27568,N_26393,N_25753);
xor U27569 (N_27569,N_26971,N_26761);
nand U27570 (N_27570,N_26503,N_26335);
nand U27571 (N_27571,N_26351,N_26870);
nor U27572 (N_27572,N_26260,N_26826);
nand U27573 (N_27573,N_26507,N_26220);
nor U27574 (N_27574,N_26309,N_26419);
and U27575 (N_27575,N_26092,N_26928);
or U27576 (N_27576,N_26433,N_26790);
nor U27577 (N_27577,N_26331,N_26359);
and U27578 (N_27578,N_25778,N_26979);
xnor U27579 (N_27579,N_26497,N_26741);
and U27580 (N_27580,N_26073,N_26150);
and U27581 (N_27581,N_26510,N_26266);
and U27582 (N_27582,N_26787,N_26348);
nor U27583 (N_27583,N_25894,N_26678);
xnor U27584 (N_27584,N_26550,N_26170);
xor U27585 (N_27585,N_26956,N_26146);
or U27586 (N_27586,N_25945,N_25652);
xnor U27587 (N_27587,N_26184,N_26944);
xor U27588 (N_27588,N_25861,N_26356);
and U27589 (N_27589,N_26662,N_26130);
nor U27590 (N_27590,N_26825,N_25821);
and U27591 (N_27591,N_26034,N_26179);
xnor U27592 (N_27592,N_25529,N_26819);
nand U27593 (N_27593,N_26060,N_25949);
nand U27594 (N_27594,N_26218,N_26953);
and U27595 (N_27595,N_26706,N_26570);
and U27596 (N_27596,N_26699,N_25621);
xor U27597 (N_27597,N_26843,N_26328);
or U27598 (N_27598,N_26506,N_26926);
xor U27599 (N_27599,N_26480,N_25793);
or U27600 (N_27600,N_25764,N_25704);
nor U27601 (N_27601,N_25995,N_26389);
xor U27602 (N_27602,N_25775,N_26760);
and U27603 (N_27603,N_26938,N_26990);
xor U27604 (N_27604,N_26033,N_26336);
or U27605 (N_27605,N_26614,N_26145);
and U27606 (N_27606,N_25579,N_26093);
nand U27607 (N_27607,N_26658,N_25769);
nand U27608 (N_27608,N_26833,N_25780);
nand U27609 (N_27609,N_26300,N_25967);
nor U27610 (N_27610,N_26252,N_26955);
nor U27611 (N_27611,N_26960,N_26090);
xnor U27612 (N_27612,N_26477,N_26616);
xnor U27613 (N_27613,N_26388,N_25787);
and U27614 (N_27614,N_26415,N_26416);
xnor U27615 (N_27615,N_26157,N_25800);
and U27616 (N_27616,N_26877,N_26302);
and U27617 (N_27617,N_26296,N_26578);
nor U27618 (N_27618,N_25591,N_26627);
or U27619 (N_27619,N_25867,N_26267);
and U27620 (N_27620,N_26177,N_26850);
nor U27621 (N_27621,N_25847,N_26085);
nand U27622 (N_27622,N_26299,N_26297);
xnor U27623 (N_27623,N_25881,N_26412);
and U27624 (N_27624,N_26936,N_25802);
nor U27625 (N_27625,N_26632,N_26027);
nand U27626 (N_27626,N_25833,N_26803);
nand U27627 (N_27627,N_25715,N_25895);
and U27628 (N_27628,N_26404,N_25693);
or U27629 (N_27629,N_25779,N_25653);
nand U27630 (N_27630,N_26369,N_25796);
xor U27631 (N_27631,N_26018,N_26666);
or U27632 (N_27632,N_26301,N_26281);
nor U27633 (N_27633,N_25526,N_26758);
xor U27634 (N_27634,N_25661,N_25710);
and U27635 (N_27635,N_26174,N_26786);
xnor U27636 (N_27636,N_26223,N_26917);
or U27637 (N_27637,N_26656,N_26626);
nand U27638 (N_27638,N_25520,N_26246);
or U27639 (N_27639,N_26432,N_25638);
or U27640 (N_27640,N_26357,N_26496);
or U27641 (N_27641,N_25581,N_26592);
and U27642 (N_27642,N_25604,N_26807);
nor U27643 (N_27643,N_25952,N_25831);
xor U27644 (N_27644,N_26265,N_25518);
nor U27645 (N_27645,N_26489,N_26941);
xnor U27646 (N_27646,N_26946,N_25548);
or U27647 (N_27647,N_26746,N_26250);
nor U27648 (N_27648,N_25743,N_26074);
or U27649 (N_27649,N_26040,N_26743);
and U27650 (N_27650,N_26341,N_26752);
or U27651 (N_27651,N_26604,N_26810);
nor U27652 (N_27652,N_26726,N_26261);
xnor U27653 (N_27653,N_26867,N_26591);
and U27654 (N_27654,N_26661,N_26617);
and U27655 (N_27655,N_26608,N_26178);
nor U27656 (N_27656,N_26838,N_25863);
xnor U27657 (N_27657,N_26663,N_25587);
nor U27658 (N_27658,N_26983,N_26883);
and U27659 (N_27659,N_26391,N_25524);
xor U27660 (N_27660,N_25969,N_25768);
xor U27661 (N_27661,N_25777,N_26094);
or U27662 (N_27662,N_26277,N_26342);
and U27663 (N_27663,N_25643,N_25873);
or U27664 (N_27664,N_26378,N_26461);
or U27665 (N_27665,N_26226,N_26901);
xor U27666 (N_27666,N_26958,N_25851);
xor U27667 (N_27667,N_25941,N_26795);
or U27668 (N_27668,N_26057,N_25523);
and U27669 (N_27669,N_25841,N_25633);
nor U27670 (N_27670,N_26235,N_26914);
xnor U27671 (N_27671,N_26175,N_25609);
nor U27672 (N_27672,N_25515,N_25996);
xor U27673 (N_27673,N_26519,N_25736);
xor U27674 (N_27674,N_26330,N_25790);
nand U27675 (N_27675,N_25947,N_26224);
nand U27676 (N_27676,N_25955,N_26767);
nand U27677 (N_27677,N_26394,N_26660);
or U27678 (N_27678,N_25700,N_26652);
and U27679 (N_27679,N_25742,N_26849);
xor U27680 (N_27680,N_25698,N_25838);
nor U27681 (N_27681,N_26195,N_25639);
nor U27682 (N_27682,N_26086,N_26735);
xor U27683 (N_27683,N_25712,N_26925);
and U27684 (N_27684,N_26640,N_25760);
nor U27685 (N_27685,N_26334,N_26731);
nor U27686 (N_27686,N_25623,N_26139);
or U27687 (N_27687,N_26441,N_26321);
nand U27688 (N_27688,N_26306,N_26972);
or U27689 (N_27689,N_26298,N_26978);
or U27690 (N_27690,N_25696,N_25883);
nor U27691 (N_27691,N_26167,N_26848);
or U27692 (N_27692,N_25648,N_26212);
xor U27693 (N_27693,N_26816,N_26517);
and U27694 (N_27694,N_26370,N_26340);
or U27695 (N_27695,N_25922,N_25539);
xnor U27696 (N_27696,N_25605,N_26563);
nand U27697 (N_27697,N_26691,N_26733);
and U27698 (N_27698,N_26525,N_26756);
or U27699 (N_27699,N_26119,N_26927);
or U27700 (N_27700,N_25561,N_26924);
or U27701 (N_27701,N_25897,N_26053);
nor U27702 (N_27702,N_25525,N_26352);
or U27703 (N_27703,N_25888,N_25706);
xnor U27704 (N_27704,N_26332,N_26688);
or U27705 (N_27705,N_26840,N_25583);
or U27706 (N_27706,N_26747,N_26697);
nor U27707 (N_27707,N_26991,N_25762);
xor U27708 (N_27708,N_26450,N_25545);
nand U27709 (N_27709,N_26624,N_25667);
nor U27710 (N_27710,N_26856,N_26704);
or U27711 (N_27711,N_25634,N_25845);
or U27712 (N_27712,N_25556,N_26968);
nor U27713 (N_27713,N_26327,N_26207);
nand U27714 (N_27714,N_26413,N_26448);
or U27715 (N_27715,N_25597,N_25926);
or U27716 (N_27716,N_26974,N_25835);
nor U27717 (N_27717,N_25908,N_26380);
or U27718 (N_27718,N_26554,N_26322);
xnor U27719 (N_27719,N_25927,N_25615);
xnor U27720 (N_27720,N_26633,N_26176);
or U27721 (N_27721,N_25695,N_26047);
nand U27722 (N_27722,N_26471,N_26029);
xor U27723 (N_27723,N_26646,N_26923);
nor U27724 (N_27724,N_26722,N_26881);
nor U27725 (N_27725,N_26858,N_25647);
and U27726 (N_27726,N_26606,N_26379);
nor U27727 (N_27727,N_25774,N_26446);
or U27728 (N_27728,N_25992,N_25616);
and U27729 (N_27729,N_26949,N_25970);
nor U27730 (N_27730,N_26569,N_25627);
or U27731 (N_27731,N_25754,N_25799);
nand U27732 (N_27732,N_25636,N_26386);
and U27733 (N_27733,N_26873,N_25904);
xnor U27734 (N_27734,N_26546,N_26802);
nand U27735 (N_27735,N_26567,N_26194);
xnor U27736 (N_27736,N_26286,N_26702);
nor U27737 (N_27737,N_26964,N_25930);
nand U27738 (N_27738,N_26424,N_26249);
nor U27739 (N_27739,N_26363,N_26382);
nand U27740 (N_27740,N_26463,N_25850);
nand U27741 (N_27741,N_26206,N_26078);
xor U27742 (N_27742,N_25533,N_25809);
nand U27743 (N_27743,N_26793,N_26977);
nor U27744 (N_27744,N_25669,N_25822);
nor U27745 (N_27745,N_26693,N_25982);
nor U27746 (N_27746,N_26263,N_25540);
nand U27747 (N_27747,N_26822,N_25716);
or U27748 (N_27748,N_26796,N_26677);
xor U27749 (N_27749,N_26442,N_25572);
nor U27750 (N_27750,N_26893,N_26563);
or U27751 (N_27751,N_25517,N_26604);
xor U27752 (N_27752,N_26385,N_25755);
or U27753 (N_27753,N_26772,N_26665);
xnor U27754 (N_27754,N_26222,N_26237);
or U27755 (N_27755,N_25877,N_26028);
nand U27756 (N_27756,N_25820,N_26127);
xor U27757 (N_27757,N_26576,N_25843);
nand U27758 (N_27758,N_26106,N_26801);
or U27759 (N_27759,N_25512,N_26145);
xor U27760 (N_27760,N_26306,N_26237);
or U27761 (N_27761,N_26507,N_26418);
nand U27762 (N_27762,N_26914,N_25678);
nor U27763 (N_27763,N_25972,N_26929);
xnor U27764 (N_27764,N_25737,N_25715);
nand U27765 (N_27765,N_25540,N_25708);
nand U27766 (N_27766,N_26538,N_26177);
and U27767 (N_27767,N_26467,N_26501);
and U27768 (N_27768,N_25558,N_26226);
or U27769 (N_27769,N_25752,N_25764);
or U27770 (N_27770,N_25629,N_26925);
and U27771 (N_27771,N_26030,N_25686);
or U27772 (N_27772,N_26225,N_26653);
xor U27773 (N_27773,N_26933,N_26687);
xor U27774 (N_27774,N_26296,N_26345);
or U27775 (N_27775,N_26185,N_26326);
nor U27776 (N_27776,N_26699,N_26363);
or U27777 (N_27777,N_26173,N_25733);
nor U27778 (N_27778,N_26566,N_26138);
nor U27779 (N_27779,N_26773,N_25611);
xnor U27780 (N_27780,N_26774,N_26860);
nand U27781 (N_27781,N_25753,N_25704);
nand U27782 (N_27782,N_26820,N_25970);
nor U27783 (N_27783,N_26319,N_26853);
and U27784 (N_27784,N_26896,N_25984);
xor U27785 (N_27785,N_25508,N_25721);
or U27786 (N_27786,N_26857,N_26932);
xnor U27787 (N_27787,N_26270,N_25722);
xnor U27788 (N_27788,N_26121,N_25724);
and U27789 (N_27789,N_25950,N_26795);
and U27790 (N_27790,N_26665,N_26334);
and U27791 (N_27791,N_26055,N_26806);
and U27792 (N_27792,N_26400,N_26842);
nor U27793 (N_27793,N_25728,N_26821);
xor U27794 (N_27794,N_26530,N_26677);
nand U27795 (N_27795,N_26169,N_26778);
and U27796 (N_27796,N_26400,N_25888);
or U27797 (N_27797,N_26336,N_26380);
or U27798 (N_27798,N_25667,N_25708);
xor U27799 (N_27799,N_25610,N_26459);
nor U27800 (N_27800,N_26284,N_26958);
xor U27801 (N_27801,N_26774,N_25825);
nand U27802 (N_27802,N_25921,N_25940);
and U27803 (N_27803,N_25733,N_26842);
and U27804 (N_27804,N_26922,N_26135);
xnor U27805 (N_27805,N_26907,N_26401);
and U27806 (N_27806,N_26576,N_26749);
or U27807 (N_27807,N_26853,N_26090);
xnor U27808 (N_27808,N_26670,N_25786);
nand U27809 (N_27809,N_26214,N_26870);
xnor U27810 (N_27810,N_26222,N_25822);
nand U27811 (N_27811,N_25731,N_25666);
nor U27812 (N_27812,N_25859,N_25680);
or U27813 (N_27813,N_26778,N_26258);
or U27814 (N_27814,N_25580,N_25955);
or U27815 (N_27815,N_26040,N_26340);
or U27816 (N_27816,N_26899,N_26994);
and U27817 (N_27817,N_26583,N_25799);
or U27818 (N_27818,N_26708,N_25987);
or U27819 (N_27819,N_26326,N_25951);
nand U27820 (N_27820,N_26689,N_26662);
and U27821 (N_27821,N_26796,N_26599);
nor U27822 (N_27822,N_26665,N_25570);
or U27823 (N_27823,N_26796,N_26035);
nand U27824 (N_27824,N_25772,N_26899);
nand U27825 (N_27825,N_26003,N_26773);
xor U27826 (N_27826,N_26208,N_25792);
and U27827 (N_27827,N_25762,N_26420);
xnor U27828 (N_27828,N_26404,N_26740);
or U27829 (N_27829,N_25644,N_26547);
or U27830 (N_27830,N_25514,N_26744);
nor U27831 (N_27831,N_26988,N_25953);
and U27832 (N_27832,N_26941,N_26710);
or U27833 (N_27833,N_26335,N_25944);
or U27834 (N_27834,N_26970,N_25650);
or U27835 (N_27835,N_26606,N_26586);
nand U27836 (N_27836,N_26111,N_25882);
or U27837 (N_27837,N_26987,N_25526);
xnor U27838 (N_27838,N_26056,N_26151);
and U27839 (N_27839,N_25838,N_26993);
nand U27840 (N_27840,N_26315,N_26295);
nand U27841 (N_27841,N_26326,N_26959);
xor U27842 (N_27842,N_26748,N_25522);
and U27843 (N_27843,N_26597,N_26519);
xor U27844 (N_27844,N_25697,N_26194);
or U27845 (N_27845,N_26695,N_26846);
nor U27846 (N_27846,N_26625,N_25574);
and U27847 (N_27847,N_25910,N_26593);
xor U27848 (N_27848,N_25763,N_25742);
and U27849 (N_27849,N_26755,N_25580);
and U27850 (N_27850,N_26924,N_26827);
xnor U27851 (N_27851,N_26507,N_25700);
xor U27852 (N_27852,N_26855,N_25523);
or U27853 (N_27853,N_26525,N_26146);
nand U27854 (N_27854,N_26672,N_25630);
xor U27855 (N_27855,N_26594,N_26974);
nand U27856 (N_27856,N_25522,N_25896);
or U27857 (N_27857,N_26161,N_25674);
nor U27858 (N_27858,N_25867,N_26261);
xnor U27859 (N_27859,N_25506,N_26474);
or U27860 (N_27860,N_25683,N_25840);
nand U27861 (N_27861,N_26750,N_26092);
nor U27862 (N_27862,N_25623,N_26659);
and U27863 (N_27863,N_25789,N_25512);
or U27864 (N_27864,N_26633,N_26391);
and U27865 (N_27865,N_26891,N_25733);
nand U27866 (N_27866,N_26958,N_26848);
or U27867 (N_27867,N_25715,N_26784);
nor U27868 (N_27868,N_26144,N_25641);
xor U27869 (N_27869,N_26269,N_25831);
xnor U27870 (N_27870,N_26531,N_26800);
nor U27871 (N_27871,N_25620,N_25974);
nand U27872 (N_27872,N_25736,N_25515);
and U27873 (N_27873,N_26096,N_25574);
and U27874 (N_27874,N_26144,N_26253);
and U27875 (N_27875,N_26236,N_26616);
nor U27876 (N_27876,N_26615,N_25530);
xnor U27877 (N_27877,N_25683,N_25901);
nand U27878 (N_27878,N_26999,N_26548);
or U27879 (N_27879,N_26924,N_26565);
and U27880 (N_27880,N_25595,N_26081);
xor U27881 (N_27881,N_26016,N_25576);
or U27882 (N_27882,N_26917,N_26615);
nor U27883 (N_27883,N_26240,N_25825);
nand U27884 (N_27884,N_26699,N_26338);
or U27885 (N_27885,N_26125,N_26507);
nand U27886 (N_27886,N_26451,N_26912);
nor U27887 (N_27887,N_25527,N_26700);
nor U27888 (N_27888,N_26885,N_26874);
nor U27889 (N_27889,N_25902,N_26332);
xor U27890 (N_27890,N_26358,N_26478);
xor U27891 (N_27891,N_25963,N_25695);
nor U27892 (N_27892,N_26412,N_25984);
nand U27893 (N_27893,N_26466,N_26176);
xnor U27894 (N_27894,N_25758,N_25671);
nand U27895 (N_27895,N_25829,N_25723);
nand U27896 (N_27896,N_26580,N_26997);
xnor U27897 (N_27897,N_26917,N_26049);
nand U27898 (N_27898,N_25957,N_25601);
xor U27899 (N_27899,N_25880,N_26243);
or U27900 (N_27900,N_25521,N_26816);
xor U27901 (N_27901,N_25777,N_26063);
nand U27902 (N_27902,N_25525,N_25743);
xnor U27903 (N_27903,N_26913,N_26559);
nand U27904 (N_27904,N_25914,N_25520);
nor U27905 (N_27905,N_26685,N_26775);
nor U27906 (N_27906,N_25687,N_26313);
nand U27907 (N_27907,N_26323,N_26752);
or U27908 (N_27908,N_26393,N_26216);
or U27909 (N_27909,N_25539,N_26727);
nand U27910 (N_27910,N_25541,N_26791);
nor U27911 (N_27911,N_26166,N_25590);
nand U27912 (N_27912,N_26464,N_25607);
or U27913 (N_27913,N_26143,N_26412);
nand U27914 (N_27914,N_25638,N_26209);
nor U27915 (N_27915,N_25831,N_25697);
nor U27916 (N_27916,N_26912,N_25759);
nand U27917 (N_27917,N_26990,N_25814);
and U27918 (N_27918,N_25787,N_25696);
nor U27919 (N_27919,N_26993,N_26340);
nor U27920 (N_27920,N_26369,N_25690);
nand U27921 (N_27921,N_26836,N_26251);
or U27922 (N_27922,N_26409,N_26841);
nor U27923 (N_27923,N_25713,N_25591);
and U27924 (N_27924,N_26000,N_26996);
nand U27925 (N_27925,N_26849,N_25730);
and U27926 (N_27926,N_25888,N_26130);
and U27927 (N_27927,N_26543,N_26568);
or U27928 (N_27928,N_25588,N_26584);
and U27929 (N_27929,N_26750,N_26231);
or U27930 (N_27930,N_26849,N_26097);
nand U27931 (N_27931,N_26756,N_26229);
xnor U27932 (N_27932,N_26537,N_25532);
nor U27933 (N_27933,N_26032,N_25791);
and U27934 (N_27934,N_26401,N_25679);
xor U27935 (N_27935,N_26806,N_26111);
and U27936 (N_27936,N_26896,N_26670);
nand U27937 (N_27937,N_25786,N_26847);
or U27938 (N_27938,N_25873,N_25669);
nor U27939 (N_27939,N_26759,N_26328);
and U27940 (N_27940,N_26294,N_25859);
and U27941 (N_27941,N_26957,N_26295);
xnor U27942 (N_27942,N_25693,N_26280);
xor U27943 (N_27943,N_26222,N_26227);
nand U27944 (N_27944,N_26680,N_26991);
nand U27945 (N_27945,N_26131,N_26819);
nor U27946 (N_27946,N_26368,N_25948);
and U27947 (N_27947,N_25903,N_25731);
and U27948 (N_27948,N_26335,N_25898);
or U27949 (N_27949,N_25598,N_26998);
nor U27950 (N_27950,N_26396,N_26316);
and U27951 (N_27951,N_26961,N_25754);
or U27952 (N_27952,N_26405,N_25860);
xnor U27953 (N_27953,N_25925,N_26720);
nand U27954 (N_27954,N_26655,N_26483);
nand U27955 (N_27955,N_26466,N_26639);
or U27956 (N_27956,N_26262,N_26137);
nor U27957 (N_27957,N_26337,N_26624);
and U27958 (N_27958,N_26888,N_26749);
nand U27959 (N_27959,N_26094,N_26001);
xor U27960 (N_27960,N_26501,N_25628);
nand U27961 (N_27961,N_26953,N_25671);
nor U27962 (N_27962,N_25767,N_25845);
and U27963 (N_27963,N_26933,N_26682);
or U27964 (N_27964,N_25915,N_26954);
nand U27965 (N_27965,N_26083,N_26847);
or U27966 (N_27966,N_26943,N_26966);
and U27967 (N_27967,N_25730,N_25677);
and U27968 (N_27968,N_25974,N_25866);
nand U27969 (N_27969,N_26647,N_26457);
or U27970 (N_27970,N_26249,N_25747);
nor U27971 (N_27971,N_26290,N_26531);
or U27972 (N_27972,N_26779,N_25825);
and U27973 (N_27973,N_25650,N_26583);
nor U27974 (N_27974,N_26892,N_26439);
and U27975 (N_27975,N_26364,N_25511);
nor U27976 (N_27976,N_26248,N_26977);
xor U27977 (N_27977,N_25657,N_26044);
or U27978 (N_27978,N_26449,N_26909);
and U27979 (N_27979,N_26917,N_25786);
and U27980 (N_27980,N_25940,N_26587);
or U27981 (N_27981,N_25870,N_26672);
nand U27982 (N_27982,N_25981,N_26644);
nand U27983 (N_27983,N_25888,N_25508);
nand U27984 (N_27984,N_26501,N_26144);
xnor U27985 (N_27985,N_25713,N_26178);
nand U27986 (N_27986,N_25636,N_25565);
and U27987 (N_27987,N_25747,N_26526);
nor U27988 (N_27988,N_26052,N_26835);
nand U27989 (N_27989,N_26850,N_25777);
xnor U27990 (N_27990,N_25978,N_25914);
and U27991 (N_27991,N_26743,N_26848);
nor U27992 (N_27992,N_26898,N_26799);
nor U27993 (N_27993,N_26799,N_26380);
nand U27994 (N_27994,N_26891,N_25856);
nor U27995 (N_27995,N_26385,N_25591);
nor U27996 (N_27996,N_26715,N_26349);
and U27997 (N_27997,N_26075,N_25931);
xor U27998 (N_27998,N_26080,N_26989);
nor U27999 (N_27999,N_26606,N_26783);
or U28000 (N_28000,N_26981,N_26984);
nand U28001 (N_28001,N_26428,N_26958);
and U28002 (N_28002,N_26848,N_26027);
nand U28003 (N_28003,N_25558,N_26506);
nor U28004 (N_28004,N_25708,N_25616);
or U28005 (N_28005,N_26439,N_26600);
and U28006 (N_28006,N_26806,N_25902);
nand U28007 (N_28007,N_26436,N_26195);
xnor U28008 (N_28008,N_26241,N_26640);
nand U28009 (N_28009,N_26425,N_26036);
nor U28010 (N_28010,N_26685,N_26552);
xnor U28011 (N_28011,N_25700,N_26375);
nand U28012 (N_28012,N_26174,N_25795);
and U28013 (N_28013,N_26776,N_25676);
xor U28014 (N_28014,N_26029,N_26099);
nor U28015 (N_28015,N_26093,N_26089);
and U28016 (N_28016,N_26236,N_26779);
nor U28017 (N_28017,N_25843,N_26258);
or U28018 (N_28018,N_25984,N_26250);
and U28019 (N_28019,N_25831,N_26259);
nand U28020 (N_28020,N_26331,N_26667);
xor U28021 (N_28021,N_25517,N_26194);
or U28022 (N_28022,N_25715,N_25873);
nor U28023 (N_28023,N_25793,N_26471);
nand U28024 (N_28024,N_25575,N_26826);
nor U28025 (N_28025,N_26406,N_26896);
and U28026 (N_28026,N_26325,N_26244);
and U28027 (N_28027,N_26729,N_26739);
xnor U28028 (N_28028,N_26559,N_26373);
xor U28029 (N_28029,N_25637,N_25873);
xnor U28030 (N_28030,N_26227,N_26979);
nor U28031 (N_28031,N_26771,N_25560);
or U28032 (N_28032,N_26022,N_26382);
nand U28033 (N_28033,N_25948,N_26623);
nor U28034 (N_28034,N_26654,N_26180);
xor U28035 (N_28035,N_25607,N_26245);
nor U28036 (N_28036,N_26897,N_26618);
and U28037 (N_28037,N_25647,N_26535);
or U28038 (N_28038,N_25743,N_26057);
xor U28039 (N_28039,N_25649,N_26929);
or U28040 (N_28040,N_26590,N_26899);
nand U28041 (N_28041,N_26564,N_26390);
nor U28042 (N_28042,N_26398,N_26813);
nand U28043 (N_28043,N_25753,N_26731);
nor U28044 (N_28044,N_26670,N_26191);
nand U28045 (N_28045,N_26819,N_26943);
and U28046 (N_28046,N_26194,N_25868);
nor U28047 (N_28047,N_26557,N_26098);
xor U28048 (N_28048,N_25890,N_26560);
nor U28049 (N_28049,N_26025,N_26483);
nor U28050 (N_28050,N_26515,N_25622);
or U28051 (N_28051,N_26101,N_26665);
xor U28052 (N_28052,N_26971,N_25619);
and U28053 (N_28053,N_25862,N_25791);
nor U28054 (N_28054,N_26419,N_26918);
or U28055 (N_28055,N_25764,N_26520);
nand U28056 (N_28056,N_25531,N_26298);
and U28057 (N_28057,N_26406,N_26029);
or U28058 (N_28058,N_25704,N_26281);
nor U28059 (N_28059,N_26694,N_26703);
xor U28060 (N_28060,N_26879,N_26273);
or U28061 (N_28061,N_26225,N_25733);
or U28062 (N_28062,N_26207,N_26007);
or U28063 (N_28063,N_26346,N_25962);
or U28064 (N_28064,N_25727,N_25942);
xnor U28065 (N_28065,N_25792,N_26596);
nand U28066 (N_28066,N_25583,N_26102);
nor U28067 (N_28067,N_25833,N_26251);
and U28068 (N_28068,N_26140,N_25928);
xor U28069 (N_28069,N_26957,N_26356);
and U28070 (N_28070,N_26375,N_25959);
nor U28071 (N_28071,N_26562,N_25703);
xor U28072 (N_28072,N_25652,N_25967);
or U28073 (N_28073,N_26563,N_26874);
or U28074 (N_28074,N_25669,N_25940);
and U28075 (N_28075,N_26244,N_25875);
xnor U28076 (N_28076,N_26256,N_25774);
or U28077 (N_28077,N_26263,N_26530);
nor U28078 (N_28078,N_26248,N_25600);
xor U28079 (N_28079,N_26420,N_26244);
xnor U28080 (N_28080,N_25952,N_26444);
xnor U28081 (N_28081,N_25859,N_25649);
xor U28082 (N_28082,N_26654,N_26943);
xor U28083 (N_28083,N_26355,N_25792);
and U28084 (N_28084,N_26011,N_26100);
nand U28085 (N_28085,N_25689,N_25655);
and U28086 (N_28086,N_26318,N_26313);
xnor U28087 (N_28087,N_25611,N_25631);
and U28088 (N_28088,N_26999,N_26621);
xnor U28089 (N_28089,N_25693,N_26723);
and U28090 (N_28090,N_26454,N_26734);
nand U28091 (N_28091,N_26004,N_26344);
or U28092 (N_28092,N_25968,N_26946);
and U28093 (N_28093,N_26098,N_26263);
nor U28094 (N_28094,N_26559,N_26735);
nor U28095 (N_28095,N_26442,N_26116);
or U28096 (N_28096,N_26995,N_25889);
and U28097 (N_28097,N_26764,N_25976);
or U28098 (N_28098,N_26489,N_26755);
or U28099 (N_28099,N_26941,N_26184);
or U28100 (N_28100,N_26363,N_26980);
or U28101 (N_28101,N_26448,N_26340);
and U28102 (N_28102,N_26705,N_26454);
and U28103 (N_28103,N_26848,N_26275);
or U28104 (N_28104,N_26294,N_26297);
or U28105 (N_28105,N_25807,N_26837);
and U28106 (N_28106,N_26969,N_25834);
nand U28107 (N_28107,N_26041,N_26313);
and U28108 (N_28108,N_25733,N_26668);
or U28109 (N_28109,N_26274,N_26518);
nor U28110 (N_28110,N_26090,N_26920);
and U28111 (N_28111,N_26284,N_26213);
or U28112 (N_28112,N_26493,N_26053);
nand U28113 (N_28113,N_25955,N_26282);
nand U28114 (N_28114,N_25511,N_26532);
or U28115 (N_28115,N_25964,N_26160);
nand U28116 (N_28116,N_26471,N_26531);
or U28117 (N_28117,N_26601,N_26360);
or U28118 (N_28118,N_26275,N_26508);
nand U28119 (N_28119,N_26922,N_25576);
nor U28120 (N_28120,N_26640,N_26631);
xnor U28121 (N_28121,N_26061,N_25954);
or U28122 (N_28122,N_26434,N_26503);
xor U28123 (N_28123,N_26201,N_26299);
xnor U28124 (N_28124,N_25857,N_26180);
xnor U28125 (N_28125,N_26812,N_26301);
and U28126 (N_28126,N_26956,N_26161);
nor U28127 (N_28127,N_26153,N_26373);
and U28128 (N_28128,N_25665,N_25601);
or U28129 (N_28129,N_25662,N_25613);
and U28130 (N_28130,N_26572,N_26617);
nor U28131 (N_28131,N_26471,N_25936);
nand U28132 (N_28132,N_25893,N_26925);
or U28133 (N_28133,N_26219,N_26538);
and U28134 (N_28134,N_25862,N_26384);
and U28135 (N_28135,N_25611,N_26886);
nand U28136 (N_28136,N_26777,N_26812);
nor U28137 (N_28137,N_26288,N_26965);
nand U28138 (N_28138,N_25517,N_25673);
xnor U28139 (N_28139,N_26121,N_26316);
or U28140 (N_28140,N_25935,N_26809);
xnor U28141 (N_28141,N_26575,N_25703);
and U28142 (N_28142,N_25972,N_26854);
or U28143 (N_28143,N_25717,N_25589);
xor U28144 (N_28144,N_26359,N_25592);
xnor U28145 (N_28145,N_26962,N_26295);
and U28146 (N_28146,N_26504,N_25944);
nand U28147 (N_28147,N_25993,N_26116);
or U28148 (N_28148,N_25625,N_25942);
or U28149 (N_28149,N_26047,N_25792);
nand U28150 (N_28150,N_25543,N_26679);
xor U28151 (N_28151,N_25684,N_25858);
nor U28152 (N_28152,N_26263,N_25639);
xor U28153 (N_28153,N_26387,N_26294);
or U28154 (N_28154,N_26900,N_25634);
nand U28155 (N_28155,N_25828,N_26907);
nor U28156 (N_28156,N_25502,N_26350);
nor U28157 (N_28157,N_26465,N_26568);
and U28158 (N_28158,N_26083,N_26885);
or U28159 (N_28159,N_26734,N_26002);
xnor U28160 (N_28160,N_25976,N_26690);
xor U28161 (N_28161,N_26799,N_25680);
xor U28162 (N_28162,N_25528,N_26992);
and U28163 (N_28163,N_26501,N_26072);
nor U28164 (N_28164,N_25780,N_26178);
nand U28165 (N_28165,N_26887,N_26683);
nor U28166 (N_28166,N_26404,N_26331);
xor U28167 (N_28167,N_25824,N_26340);
and U28168 (N_28168,N_26598,N_26188);
nand U28169 (N_28169,N_26022,N_26886);
nor U28170 (N_28170,N_26529,N_25617);
or U28171 (N_28171,N_26812,N_25971);
xor U28172 (N_28172,N_26462,N_25606);
nand U28173 (N_28173,N_26254,N_26765);
and U28174 (N_28174,N_26804,N_26129);
or U28175 (N_28175,N_25785,N_26661);
and U28176 (N_28176,N_26906,N_25650);
or U28177 (N_28177,N_25726,N_26806);
or U28178 (N_28178,N_26935,N_26134);
or U28179 (N_28179,N_25927,N_26384);
xor U28180 (N_28180,N_26049,N_26597);
xnor U28181 (N_28181,N_26445,N_26849);
nand U28182 (N_28182,N_26101,N_26650);
or U28183 (N_28183,N_26109,N_25757);
and U28184 (N_28184,N_25937,N_26721);
xor U28185 (N_28185,N_26892,N_26410);
and U28186 (N_28186,N_26617,N_26291);
xnor U28187 (N_28187,N_26171,N_25911);
or U28188 (N_28188,N_25847,N_25640);
nand U28189 (N_28189,N_26438,N_25750);
xor U28190 (N_28190,N_25709,N_26717);
nand U28191 (N_28191,N_26140,N_26334);
xnor U28192 (N_28192,N_26129,N_25574);
xnor U28193 (N_28193,N_26332,N_25512);
nand U28194 (N_28194,N_26170,N_26629);
and U28195 (N_28195,N_25788,N_25522);
xnor U28196 (N_28196,N_25538,N_26647);
or U28197 (N_28197,N_26443,N_26366);
and U28198 (N_28198,N_26263,N_26923);
or U28199 (N_28199,N_26926,N_25909);
and U28200 (N_28200,N_25963,N_26825);
or U28201 (N_28201,N_26970,N_26862);
nor U28202 (N_28202,N_26345,N_25617);
nor U28203 (N_28203,N_25662,N_26518);
nand U28204 (N_28204,N_25772,N_26359);
nor U28205 (N_28205,N_25871,N_26773);
nor U28206 (N_28206,N_26134,N_25724);
or U28207 (N_28207,N_25594,N_26540);
nand U28208 (N_28208,N_26196,N_26811);
nor U28209 (N_28209,N_26734,N_26554);
xnor U28210 (N_28210,N_26574,N_26971);
or U28211 (N_28211,N_25713,N_26472);
and U28212 (N_28212,N_26709,N_26774);
nand U28213 (N_28213,N_26615,N_26852);
xnor U28214 (N_28214,N_26223,N_26765);
nor U28215 (N_28215,N_26574,N_26569);
and U28216 (N_28216,N_26095,N_26764);
nand U28217 (N_28217,N_25756,N_26345);
nand U28218 (N_28218,N_26964,N_25561);
and U28219 (N_28219,N_26259,N_26640);
nand U28220 (N_28220,N_26909,N_26181);
xnor U28221 (N_28221,N_25816,N_26777);
or U28222 (N_28222,N_25790,N_25948);
nor U28223 (N_28223,N_26747,N_25622);
xnor U28224 (N_28224,N_26642,N_26659);
and U28225 (N_28225,N_26387,N_25823);
xor U28226 (N_28226,N_26286,N_26794);
nand U28227 (N_28227,N_25750,N_26748);
and U28228 (N_28228,N_26445,N_26833);
nand U28229 (N_28229,N_25672,N_26250);
nand U28230 (N_28230,N_25575,N_26115);
or U28231 (N_28231,N_26936,N_26605);
nand U28232 (N_28232,N_26376,N_26084);
xor U28233 (N_28233,N_26810,N_26873);
nand U28234 (N_28234,N_26380,N_25668);
nand U28235 (N_28235,N_26189,N_26592);
nor U28236 (N_28236,N_26751,N_25938);
xnor U28237 (N_28237,N_26470,N_26744);
xor U28238 (N_28238,N_26800,N_26956);
xnor U28239 (N_28239,N_26737,N_25885);
and U28240 (N_28240,N_26314,N_26718);
nand U28241 (N_28241,N_25794,N_26798);
nor U28242 (N_28242,N_26797,N_26482);
nand U28243 (N_28243,N_25994,N_25646);
nor U28244 (N_28244,N_26798,N_26666);
nand U28245 (N_28245,N_26650,N_25791);
xor U28246 (N_28246,N_26575,N_25573);
nand U28247 (N_28247,N_26338,N_25746);
and U28248 (N_28248,N_25528,N_25939);
xnor U28249 (N_28249,N_25713,N_26118);
nor U28250 (N_28250,N_25828,N_25942);
and U28251 (N_28251,N_25597,N_26303);
xor U28252 (N_28252,N_26737,N_26256);
or U28253 (N_28253,N_25762,N_26838);
nor U28254 (N_28254,N_25501,N_26296);
and U28255 (N_28255,N_25992,N_26640);
and U28256 (N_28256,N_25757,N_25527);
nor U28257 (N_28257,N_25739,N_26497);
or U28258 (N_28258,N_26594,N_25827);
nand U28259 (N_28259,N_26368,N_26185);
nor U28260 (N_28260,N_26178,N_26424);
or U28261 (N_28261,N_25829,N_25941);
xnor U28262 (N_28262,N_25946,N_25572);
nor U28263 (N_28263,N_26493,N_26176);
xor U28264 (N_28264,N_26831,N_26655);
xor U28265 (N_28265,N_25656,N_26340);
xnor U28266 (N_28266,N_25540,N_25802);
and U28267 (N_28267,N_25887,N_25980);
and U28268 (N_28268,N_26042,N_25838);
xnor U28269 (N_28269,N_26631,N_26655);
xnor U28270 (N_28270,N_26392,N_26163);
or U28271 (N_28271,N_25916,N_26862);
or U28272 (N_28272,N_26159,N_26680);
and U28273 (N_28273,N_26915,N_25717);
and U28274 (N_28274,N_25600,N_26437);
xor U28275 (N_28275,N_26141,N_26053);
xnor U28276 (N_28276,N_26271,N_26804);
and U28277 (N_28277,N_26370,N_26072);
xor U28278 (N_28278,N_26613,N_26993);
xor U28279 (N_28279,N_26260,N_26706);
xnor U28280 (N_28280,N_25924,N_25787);
and U28281 (N_28281,N_26754,N_26442);
or U28282 (N_28282,N_25815,N_25840);
and U28283 (N_28283,N_25869,N_26134);
and U28284 (N_28284,N_26885,N_26139);
or U28285 (N_28285,N_25959,N_26451);
nor U28286 (N_28286,N_26941,N_26970);
nor U28287 (N_28287,N_25649,N_25754);
xor U28288 (N_28288,N_25800,N_26719);
xnor U28289 (N_28289,N_25513,N_26508);
nor U28290 (N_28290,N_26512,N_26141);
and U28291 (N_28291,N_26095,N_26849);
and U28292 (N_28292,N_25717,N_26281);
xnor U28293 (N_28293,N_26824,N_25953);
or U28294 (N_28294,N_26800,N_25998);
nor U28295 (N_28295,N_26581,N_26014);
nand U28296 (N_28296,N_25705,N_25500);
xor U28297 (N_28297,N_26050,N_25549);
nand U28298 (N_28298,N_25916,N_25789);
or U28299 (N_28299,N_26270,N_25629);
and U28300 (N_28300,N_25819,N_26771);
or U28301 (N_28301,N_26253,N_26540);
nand U28302 (N_28302,N_26934,N_26502);
nand U28303 (N_28303,N_25892,N_25744);
and U28304 (N_28304,N_25787,N_26996);
and U28305 (N_28305,N_26353,N_26620);
and U28306 (N_28306,N_25505,N_26729);
xnor U28307 (N_28307,N_26839,N_26040);
nand U28308 (N_28308,N_26192,N_26950);
nor U28309 (N_28309,N_26940,N_26161);
and U28310 (N_28310,N_25985,N_26508);
nor U28311 (N_28311,N_25516,N_25636);
or U28312 (N_28312,N_26511,N_26008);
or U28313 (N_28313,N_26547,N_26074);
nor U28314 (N_28314,N_26475,N_25551);
nor U28315 (N_28315,N_26089,N_26815);
nor U28316 (N_28316,N_26127,N_26490);
xor U28317 (N_28317,N_25618,N_26353);
xor U28318 (N_28318,N_26673,N_26427);
xor U28319 (N_28319,N_25948,N_25530);
or U28320 (N_28320,N_26723,N_26917);
xnor U28321 (N_28321,N_26977,N_26098);
nand U28322 (N_28322,N_26665,N_25642);
nor U28323 (N_28323,N_25649,N_26495);
and U28324 (N_28324,N_26467,N_26632);
or U28325 (N_28325,N_26869,N_26347);
nor U28326 (N_28326,N_26282,N_26988);
nand U28327 (N_28327,N_25956,N_25643);
nand U28328 (N_28328,N_26093,N_26378);
xnor U28329 (N_28329,N_26962,N_25550);
or U28330 (N_28330,N_26554,N_26023);
or U28331 (N_28331,N_26917,N_25688);
xnor U28332 (N_28332,N_26024,N_25867);
xor U28333 (N_28333,N_26473,N_26416);
xnor U28334 (N_28334,N_25846,N_26760);
nand U28335 (N_28335,N_26786,N_26612);
nor U28336 (N_28336,N_25549,N_26420);
nor U28337 (N_28337,N_25766,N_25655);
nand U28338 (N_28338,N_26465,N_26244);
xor U28339 (N_28339,N_26904,N_26766);
nor U28340 (N_28340,N_25610,N_26737);
nand U28341 (N_28341,N_25855,N_26707);
nor U28342 (N_28342,N_25781,N_25919);
or U28343 (N_28343,N_26136,N_26842);
or U28344 (N_28344,N_26867,N_26471);
nor U28345 (N_28345,N_25872,N_25709);
or U28346 (N_28346,N_26217,N_26719);
and U28347 (N_28347,N_26023,N_25714);
xor U28348 (N_28348,N_26578,N_26594);
or U28349 (N_28349,N_25927,N_25715);
nor U28350 (N_28350,N_26459,N_25668);
xor U28351 (N_28351,N_25837,N_26766);
xor U28352 (N_28352,N_26722,N_25594);
xnor U28353 (N_28353,N_25910,N_25623);
or U28354 (N_28354,N_26421,N_26405);
nor U28355 (N_28355,N_25565,N_26314);
and U28356 (N_28356,N_25793,N_25718);
or U28357 (N_28357,N_25914,N_25629);
or U28358 (N_28358,N_26750,N_25665);
xnor U28359 (N_28359,N_26484,N_26967);
nand U28360 (N_28360,N_25574,N_26140);
and U28361 (N_28361,N_26270,N_25688);
nand U28362 (N_28362,N_25912,N_25781);
xnor U28363 (N_28363,N_26563,N_26986);
xnor U28364 (N_28364,N_26729,N_26721);
and U28365 (N_28365,N_25929,N_25655);
or U28366 (N_28366,N_26792,N_26608);
nor U28367 (N_28367,N_26554,N_26246);
nand U28368 (N_28368,N_26913,N_25847);
nand U28369 (N_28369,N_26618,N_26446);
xnor U28370 (N_28370,N_26151,N_25785);
nor U28371 (N_28371,N_25855,N_26845);
and U28372 (N_28372,N_26831,N_25939);
nand U28373 (N_28373,N_25609,N_26573);
nand U28374 (N_28374,N_26363,N_26452);
xnor U28375 (N_28375,N_25614,N_26017);
nor U28376 (N_28376,N_26651,N_26833);
or U28377 (N_28377,N_25890,N_26612);
xor U28378 (N_28378,N_26129,N_25529);
nand U28379 (N_28379,N_26371,N_26568);
xnor U28380 (N_28380,N_25756,N_25624);
and U28381 (N_28381,N_25622,N_26301);
or U28382 (N_28382,N_26437,N_26378);
nand U28383 (N_28383,N_26394,N_26274);
or U28384 (N_28384,N_25863,N_26127);
nor U28385 (N_28385,N_26719,N_26618);
nand U28386 (N_28386,N_26763,N_26918);
or U28387 (N_28387,N_26562,N_26003);
nand U28388 (N_28388,N_26442,N_26912);
or U28389 (N_28389,N_25949,N_26437);
xor U28390 (N_28390,N_26001,N_25886);
or U28391 (N_28391,N_26793,N_26186);
nand U28392 (N_28392,N_26993,N_26321);
and U28393 (N_28393,N_26437,N_26977);
nand U28394 (N_28394,N_26225,N_25801);
or U28395 (N_28395,N_25753,N_26431);
nand U28396 (N_28396,N_26490,N_26030);
nand U28397 (N_28397,N_25896,N_26583);
nor U28398 (N_28398,N_26383,N_26024);
xor U28399 (N_28399,N_26721,N_26561);
and U28400 (N_28400,N_25666,N_26151);
or U28401 (N_28401,N_26204,N_25684);
xnor U28402 (N_28402,N_26315,N_26028);
or U28403 (N_28403,N_26652,N_25780);
nor U28404 (N_28404,N_25583,N_26983);
or U28405 (N_28405,N_26034,N_25706);
nand U28406 (N_28406,N_25862,N_26465);
and U28407 (N_28407,N_26022,N_26424);
nor U28408 (N_28408,N_26106,N_26081);
nor U28409 (N_28409,N_26334,N_26824);
nand U28410 (N_28410,N_26709,N_26960);
nor U28411 (N_28411,N_25548,N_26041);
xnor U28412 (N_28412,N_26367,N_26864);
nand U28413 (N_28413,N_26456,N_26914);
nor U28414 (N_28414,N_26835,N_26471);
nand U28415 (N_28415,N_26976,N_25596);
or U28416 (N_28416,N_25936,N_26769);
and U28417 (N_28417,N_26210,N_26039);
or U28418 (N_28418,N_26178,N_26072);
and U28419 (N_28419,N_26126,N_26180);
nand U28420 (N_28420,N_25541,N_25821);
nand U28421 (N_28421,N_26746,N_26544);
xor U28422 (N_28422,N_26796,N_26981);
nand U28423 (N_28423,N_25556,N_26224);
xor U28424 (N_28424,N_26942,N_26716);
and U28425 (N_28425,N_25907,N_25777);
or U28426 (N_28426,N_25723,N_25922);
nand U28427 (N_28427,N_26631,N_26784);
nor U28428 (N_28428,N_26806,N_26968);
nand U28429 (N_28429,N_26410,N_26068);
nor U28430 (N_28430,N_26277,N_26260);
xor U28431 (N_28431,N_25992,N_26885);
nor U28432 (N_28432,N_26885,N_26030);
nand U28433 (N_28433,N_26598,N_25853);
xor U28434 (N_28434,N_26244,N_25842);
nand U28435 (N_28435,N_26310,N_25520);
and U28436 (N_28436,N_26847,N_25555);
and U28437 (N_28437,N_26540,N_25618);
or U28438 (N_28438,N_26231,N_26898);
nand U28439 (N_28439,N_26081,N_26102);
nor U28440 (N_28440,N_26701,N_25914);
nor U28441 (N_28441,N_25756,N_25595);
xnor U28442 (N_28442,N_26225,N_25697);
nor U28443 (N_28443,N_25523,N_26614);
and U28444 (N_28444,N_26465,N_26859);
xor U28445 (N_28445,N_26347,N_25757);
nand U28446 (N_28446,N_26203,N_26855);
nor U28447 (N_28447,N_26604,N_25529);
or U28448 (N_28448,N_26052,N_25740);
or U28449 (N_28449,N_25661,N_26178);
or U28450 (N_28450,N_26423,N_26112);
nor U28451 (N_28451,N_26252,N_26277);
nor U28452 (N_28452,N_26674,N_26917);
or U28453 (N_28453,N_26095,N_25692);
nand U28454 (N_28454,N_26172,N_26465);
nand U28455 (N_28455,N_25786,N_26468);
nand U28456 (N_28456,N_26843,N_26295);
nor U28457 (N_28457,N_26715,N_26194);
or U28458 (N_28458,N_25828,N_26230);
nor U28459 (N_28459,N_26415,N_26918);
and U28460 (N_28460,N_26034,N_26948);
nand U28461 (N_28461,N_25722,N_26021);
or U28462 (N_28462,N_26688,N_26930);
nand U28463 (N_28463,N_26941,N_26478);
and U28464 (N_28464,N_26307,N_26825);
and U28465 (N_28465,N_26071,N_26861);
nor U28466 (N_28466,N_26960,N_25916);
or U28467 (N_28467,N_26749,N_25972);
xor U28468 (N_28468,N_26962,N_26063);
xor U28469 (N_28469,N_26077,N_26155);
xnor U28470 (N_28470,N_26627,N_25649);
xnor U28471 (N_28471,N_26798,N_25633);
nand U28472 (N_28472,N_26589,N_25931);
and U28473 (N_28473,N_26720,N_26739);
nand U28474 (N_28474,N_25712,N_26149);
and U28475 (N_28475,N_26026,N_26795);
or U28476 (N_28476,N_25762,N_25938);
and U28477 (N_28477,N_25646,N_26077);
xor U28478 (N_28478,N_25850,N_25651);
nor U28479 (N_28479,N_25667,N_25969);
or U28480 (N_28480,N_26082,N_26522);
and U28481 (N_28481,N_26614,N_25732);
or U28482 (N_28482,N_26519,N_25834);
or U28483 (N_28483,N_25790,N_25602);
nor U28484 (N_28484,N_25549,N_25855);
or U28485 (N_28485,N_25688,N_26482);
nor U28486 (N_28486,N_26808,N_25958);
nand U28487 (N_28487,N_26978,N_26381);
or U28488 (N_28488,N_26749,N_26287);
nand U28489 (N_28489,N_26941,N_26578);
nand U28490 (N_28490,N_26905,N_25813);
or U28491 (N_28491,N_26567,N_26459);
xor U28492 (N_28492,N_25915,N_25955);
nand U28493 (N_28493,N_25924,N_25744);
or U28494 (N_28494,N_26839,N_26476);
xor U28495 (N_28495,N_26708,N_25599);
and U28496 (N_28496,N_25876,N_26276);
nand U28497 (N_28497,N_25835,N_26265);
xor U28498 (N_28498,N_26307,N_26975);
xnor U28499 (N_28499,N_26311,N_26962);
xnor U28500 (N_28500,N_27310,N_28412);
or U28501 (N_28501,N_27990,N_27216);
nand U28502 (N_28502,N_27363,N_27813);
and U28503 (N_28503,N_27064,N_28466);
and U28504 (N_28504,N_28112,N_28456);
and U28505 (N_28505,N_27308,N_28404);
nor U28506 (N_28506,N_27080,N_27034);
and U28507 (N_28507,N_28407,N_27247);
and U28508 (N_28508,N_28223,N_27858);
or U28509 (N_28509,N_27533,N_28207);
xor U28510 (N_28510,N_27014,N_27855);
and U28511 (N_28511,N_27907,N_27219);
or U28512 (N_28512,N_28353,N_27786);
xor U28513 (N_28513,N_27718,N_27576);
and U28514 (N_28514,N_27775,N_28081);
and U28515 (N_28515,N_27372,N_28137);
nor U28516 (N_28516,N_28188,N_27058);
nor U28517 (N_28517,N_27179,N_27100);
xor U28518 (N_28518,N_27838,N_27544);
nand U28519 (N_28519,N_27743,N_28428);
xor U28520 (N_28520,N_28355,N_27096);
nor U28521 (N_28521,N_28396,N_27102);
nand U28522 (N_28522,N_27202,N_28199);
nor U28523 (N_28523,N_28332,N_28113);
and U28524 (N_28524,N_27593,N_27424);
or U28525 (N_28525,N_27091,N_28493);
nand U28526 (N_28526,N_27360,N_27190);
xor U28527 (N_28527,N_28348,N_27253);
xor U28528 (N_28528,N_28044,N_28415);
xnor U28529 (N_28529,N_28279,N_27804);
nor U28530 (N_28530,N_28416,N_28383);
nor U28531 (N_28531,N_27473,N_27112);
and U28532 (N_28532,N_27975,N_27325);
nor U28533 (N_28533,N_27879,N_28234);
and U28534 (N_28534,N_28413,N_27513);
nand U28535 (N_28535,N_27146,N_27018);
and U28536 (N_28536,N_28129,N_27236);
and U28537 (N_28537,N_27688,N_27700);
and U28538 (N_28538,N_27790,N_28290);
and U28539 (N_28539,N_27303,N_27040);
and U28540 (N_28540,N_27256,N_28075);
xor U28541 (N_28541,N_28459,N_27306);
nor U28542 (N_28542,N_28489,N_27494);
or U28543 (N_28543,N_27655,N_27948);
or U28544 (N_28544,N_28121,N_27807);
xor U28545 (N_28545,N_27636,N_27368);
xnor U28546 (N_28546,N_27666,N_27892);
nand U28547 (N_28547,N_28276,N_27139);
xnor U28548 (N_28548,N_27993,N_28155);
nor U28549 (N_28549,N_28002,N_28462);
nand U28550 (N_28550,N_27489,N_27821);
nand U28551 (N_28551,N_27897,N_27152);
nand U28552 (N_28552,N_27419,N_27230);
nor U28553 (N_28553,N_27311,N_27508);
xnor U28554 (N_28554,N_27465,N_27832);
or U28555 (N_28555,N_27836,N_27931);
nor U28556 (N_28556,N_27628,N_28083);
or U28557 (N_28557,N_27232,N_27214);
and U28558 (N_28558,N_27789,N_28022);
nor U28559 (N_28559,N_27422,N_27884);
nor U28560 (N_28560,N_28449,N_28176);
nor U28561 (N_28561,N_27410,N_28340);
nor U28562 (N_28562,N_27840,N_27921);
xnor U28563 (N_28563,N_27568,N_27623);
xor U28564 (N_28564,N_27580,N_27677);
nand U28565 (N_28565,N_27449,N_27977);
nand U28566 (N_28566,N_28196,N_27564);
nand U28567 (N_28567,N_27717,N_27249);
nand U28568 (N_28568,N_27328,N_28344);
nor U28569 (N_28569,N_27397,N_27844);
nand U28570 (N_28570,N_27347,N_28209);
xor U28571 (N_28571,N_28399,N_27296);
xnor U28572 (N_28572,N_27611,N_28178);
xnor U28573 (N_28573,N_28149,N_27981);
or U28574 (N_28574,N_27209,N_27885);
and U28575 (N_28575,N_27073,N_28054);
xor U28576 (N_28576,N_28009,N_28213);
nor U28577 (N_28577,N_28485,N_27258);
nor U28578 (N_28578,N_27114,N_27367);
or U28579 (N_28579,N_27634,N_27266);
nand U28580 (N_28580,N_27778,N_27485);
or U28581 (N_28581,N_28227,N_27950);
xor U28582 (N_28582,N_27643,N_27217);
nor U28583 (N_28583,N_28319,N_27971);
xor U28584 (N_28584,N_27187,N_28088);
and U28585 (N_28585,N_28482,N_28218);
nor U28586 (N_28586,N_28401,N_28423);
and U28587 (N_28587,N_28092,N_27590);
and U28588 (N_28588,N_27183,N_27589);
nor U28589 (N_28589,N_28388,N_27346);
nand U28590 (N_28590,N_27010,N_27751);
nand U28591 (N_28591,N_27278,N_28389);
and U28592 (N_28592,N_27663,N_27859);
nor U28593 (N_28593,N_28246,N_27226);
and U28594 (N_28594,N_27326,N_27873);
and U28595 (N_28595,N_28291,N_27221);
nand U28596 (N_28596,N_27413,N_28425);
nor U28597 (N_28597,N_27733,N_28360);
nor U28598 (N_28598,N_28183,N_27127);
or U28599 (N_28599,N_27572,N_28420);
or U28600 (N_28600,N_27167,N_27758);
nand U28601 (N_28601,N_27341,N_27918);
xnor U28602 (N_28602,N_27805,N_27350);
nor U28603 (N_28603,N_27652,N_27756);
nand U28604 (N_28604,N_27160,N_27822);
and U28605 (N_28605,N_27767,N_27177);
or U28606 (N_28606,N_28241,N_27668);
nor U28607 (N_28607,N_28278,N_27357);
or U28608 (N_28608,N_27138,N_27824);
nor U28609 (N_28609,N_28451,N_27204);
xnor U28610 (N_28610,N_28032,N_28061);
nand U28611 (N_28611,N_27615,N_27358);
nor U28612 (N_28612,N_28141,N_28123);
or U28613 (N_28613,N_27366,N_27342);
and U28614 (N_28614,N_27870,N_28381);
nor U28615 (N_28615,N_27617,N_28043);
nand U28616 (N_28616,N_28023,N_27072);
and U28617 (N_28617,N_28268,N_28430);
and U28618 (N_28618,N_27452,N_27488);
nor U28619 (N_28619,N_27997,N_28496);
nand U28620 (N_28620,N_27773,N_27373);
and U28621 (N_28621,N_28358,N_27288);
and U28622 (N_28622,N_28216,N_27106);
and U28623 (N_28623,N_27588,N_28331);
or U28624 (N_28624,N_28219,N_27240);
or U28625 (N_28625,N_27047,N_27039);
or U28626 (N_28626,N_27706,N_27754);
nor U28627 (N_28627,N_27637,N_27481);
nor U28628 (N_28628,N_28439,N_27770);
or U28629 (N_28629,N_27947,N_28147);
or U28630 (N_28630,N_27168,N_27330);
or U28631 (N_28631,N_27052,N_28245);
or U28632 (N_28632,N_28136,N_28084);
xnor U28633 (N_28633,N_27888,N_28168);
nand U28634 (N_28634,N_27799,N_27672);
and U28635 (N_28635,N_27188,N_28078);
nand U28636 (N_28636,N_28217,N_27523);
nand U28637 (N_28637,N_27491,N_27430);
nor U28638 (N_28638,N_28326,N_28110);
and U28639 (N_28639,N_27548,N_28177);
xnor U28640 (N_28640,N_27131,N_27156);
or U28641 (N_28641,N_27432,N_27173);
nand U28642 (N_28642,N_28492,N_27268);
xnor U28643 (N_28643,N_28013,N_27653);
xnor U28644 (N_28644,N_27697,N_27881);
nor U28645 (N_28645,N_28247,N_27493);
nand U28646 (N_28646,N_27792,N_28214);
nand U28647 (N_28647,N_27536,N_27684);
nor U28648 (N_28648,N_27246,N_27462);
and U28649 (N_28649,N_27895,N_27283);
nand U28650 (N_28650,N_27354,N_27763);
and U28651 (N_28651,N_27999,N_27779);
xnor U28652 (N_28652,N_27293,N_27675);
nor U28653 (N_28653,N_28455,N_27798);
xor U28654 (N_28654,N_27498,N_27499);
nand U28655 (N_28655,N_27055,N_27995);
xor U28656 (N_28656,N_28488,N_27414);
nor U28657 (N_28657,N_27746,N_27864);
xnor U28658 (N_28658,N_27029,N_27049);
and U28659 (N_28659,N_27336,N_27017);
and U28660 (N_28660,N_28049,N_28060);
xor U28661 (N_28661,N_28487,N_28150);
nand U28662 (N_28662,N_27186,N_27448);
or U28663 (N_28663,N_28313,N_28342);
or U28664 (N_28664,N_27930,N_27134);
or U28665 (N_28665,N_27954,N_27126);
and U28666 (N_28666,N_27104,N_27483);
xnor U28667 (N_28667,N_27027,N_27932);
and U28668 (N_28668,N_27674,N_27043);
nand U28669 (N_28669,N_28408,N_28352);
or U28670 (N_28670,N_27551,N_27955);
nand U28671 (N_28671,N_27327,N_27915);
nor U28672 (N_28672,N_27708,N_28122);
nand U28673 (N_28673,N_28292,N_28314);
or U28674 (N_28674,N_28051,N_27871);
and U28675 (N_28675,N_27914,N_28156);
nor U28676 (N_28676,N_28167,N_28202);
or U28677 (N_28677,N_27255,N_27009);
xnor U28678 (N_28678,N_27478,N_27317);
or U28679 (N_28679,N_28484,N_27264);
or U28680 (N_28680,N_27391,N_27348);
xnor U28681 (N_28681,N_28153,N_28042);
and U28682 (N_28682,N_28180,N_27322);
xnor U28683 (N_28683,N_27776,N_27290);
nor U28684 (N_28684,N_28463,N_28095);
and U28685 (N_28685,N_27045,N_28094);
nand U28686 (N_28686,N_27678,N_27899);
or U28687 (N_28687,N_27861,N_28190);
nand U28688 (N_28688,N_27012,N_27853);
xnor U28689 (N_28689,N_28139,N_27974);
or U28690 (N_28690,N_27889,N_27111);
xor U28691 (N_28691,N_27528,N_28166);
nand U28692 (N_28692,N_27624,N_27123);
nor U28693 (N_28693,N_27951,N_27594);
xor U28694 (N_28694,N_28001,N_28034);
xor U28695 (N_28695,N_27297,N_28300);
nand U28696 (N_28696,N_28473,N_27782);
nor U28697 (N_28697,N_27978,N_27679);
or U28698 (N_28698,N_27562,N_27644);
nor U28699 (N_28699,N_27713,N_27143);
or U28700 (N_28700,N_28323,N_27845);
nand U28701 (N_28701,N_27911,N_28030);
nor U28702 (N_28702,N_28028,N_28098);
and U28703 (N_28703,N_27002,N_27965);
and U28704 (N_28704,N_28371,N_27431);
xor U28705 (N_28705,N_27570,N_27760);
and U28706 (N_28706,N_28351,N_27878);
nand U28707 (N_28707,N_27319,N_27060);
nand U28708 (N_28708,N_28441,N_27711);
nand U28709 (N_28709,N_27436,N_27400);
or U28710 (N_28710,N_27086,N_28405);
xor U28711 (N_28711,N_28363,N_28115);
nand U28712 (N_28712,N_28090,N_27969);
xnor U28713 (N_28713,N_27492,N_28382);
nand U28714 (N_28714,N_27857,N_27459);
and U28715 (N_28715,N_27231,N_28373);
and U28716 (N_28716,N_28429,N_28135);
and U28717 (N_28717,N_27817,N_27957);
nand U28718 (N_28718,N_27208,N_28179);
xor U28719 (N_28719,N_27835,N_28158);
or U28720 (N_28720,N_27116,N_27630);
or U28721 (N_28721,N_27683,N_28200);
nand U28722 (N_28722,N_27441,N_28230);
or U28723 (N_28723,N_27245,N_27834);
nor U28724 (N_28724,N_28045,N_28447);
and U28725 (N_28725,N_28187,N_27720);
and U28726 (N_28726,N_27987,N_27164);
nor U28727 (N_28727,N_27170,N_27937);
and U28728 (N_28728,N_28171,N_27385);
nand U28729 (N_28729,N_28232,N_27059);
nor U28730 (N_28730,N_28134,N_27279);
xnor U28731 (N_28731,N_27768,N_27189);
or U28732 (N_28732,N_27598,N_28008);
and U28733 (N_28733,N_27867,N_27517);
and U28734 (N_28734,N_28309,N_27178);
or U28735 (N_28735,N_28359,N_27933);
or U28736 (N_28736,N_27893,N_28233);
nor U28737 (N_28737,N_27235,N_27740);
nand U28738 (N_28738,N_28310,N_27891);
or U28739 (N_28739,N_28470,N_27090);
or U28740 (N_28740,N_27998,N_28418);
nand U28741 (N_28741,N_28080,N_27890);
and U28742 (N_28742,N_28341,N_28460);
and U28743 (N_28743,N_28469,N_28427);
or U28744 (N_28744,N_27466,N_28333);
xor U28745 (N_28745,N_28303,N_27103);
xnor U28746 (N_28746,N_28370,N_28288);
nor U28747 (N_28747,N_27607,N_28266);
xor U28748 (N_28748,N_27257,N_27613);
nand U28749 (N_28749,N_27901,N_28262);
or U28750 (N_28750,N_27145,N_28375);
and U28751 (N_28751,N_27051,N_27560);
nand U28752 (N_28752,N_27375,N_27195);
nor U28753 (N_28753,N_27712,N_27359);
and U28754 (N_28754,N_28099,N_27755);
and U28755 (N_28755,N_28283,N_27401);
and U28756 (N_28756,N_28221,N_28033);
nor U28757 (N_28757,N_27956,N_27180);
nor U28758 (N_28758,N_27693,N_28374);
nor U28759 (N_28759,N_27352,N_27622);
nand U28760 (N_28760,N_27934,N_27333);
nor U28761 (N_28761,N_27282,N_28263);
and U28762 (N_28762,N_27913,N_27816);
nand U28763 (N_28763,N_28071,N_27691);
nor U28764 (N_28764,N_27982,N_27285);
or U28765 (N_28765,N_28362,N_27984);
xor U28766 (N_28766,N_27582,N_27894);
nor U28767 (N_28767,N_28464,N_27093);
or U28768 (N_28768,N_27966,N_27004);
nand U28769 (N_28769,N_27196,N_28029);
nand U28770 (N_28770,N_27631,N_27592);
nor U28771 (N_28771,N_27815,N_28164);
nor U28772 (N_28772,N_27726,N_27062);
nand U28773 (N_28773,N_28119,N_27550);
xnor U28774 (N_28774,N_27411,N_28142);
nor U28775 (N_28775,N_27689,N_27107);
xor U28776 (N_28776,N_27554,N_27651);
xor U28777 (N_28777,N_28306,N_28105);
nor U28778 (N_28778,N_28194,N_28437);
xor U28779 (N_28779,N_28387,N_27757);
nand U28780 (N_28780,N_27722,N_27021);
or U28781 (N_28781,N_27117,N_27752);
and U28782 (N_28782,N_27862,N_27406);
and U28783 (N_28783,N_27929,N_27682);
xnor U28784 (N_28784,N_27985,N_28184);
nand U28785 (N_28785,N_28361,N_27159);
or U28786 (N_28786,N_27201,N_27670);
and U28787 (N_28787,N_27001,N_28481);
nand U28788 (N_28788,N_27353,N_27656);
xor U28789 (N_28789,N_27113,N_27181);
or U28790 (N_28790,N_27182,N_28175);
xnor U28791 (N_28791,N_28025,N_28499);
nor U28792 (N_28792,N_27587,N_27584);
nand U28793 (N_28793,N_28014,N_27785);
xor U28794 (N_28794,N_27161,N_27676);
nand U28795 (N_28795,N_27783,N_28055);
nand U28796 (N_28796,N_28458,N_28284);
nor U28797 (N_28797,N_27084,N_27166);
nor U28798 (N_28798,N_28379,N_28308);
xnor U28799 (N_28799,N_27962,N_27635);
or U28800 (N_28800,N_28229,N_27239);
and U28801 (N_28801,N_28478,N_27140);
or U28802 (N_28802,N_28311,N_28254);
nor U28803 (N_28803,N_27866,N_28243);
nor U28804 (N_28804,N_27337,N_27942);
nand U28805 (N_28805,N_28157,N_28320);
and U28806 (N_28806,N_27447,N_28063);
and U28807 (N_28807,N_27780,N_28345);
nor U28808 (N_28808,N_27271,N_27471);
and U28809 (N_28809,N_28210,N_27772);
xnor U28810 (N_28810,N_27263,N_28046);
xnor U28811 (N_28811,N_28445,N_27645);
nor U28812 (N_28812,N_27714,N_27595);
or U28813 (N_28813,N_28208,N_28047);
or U28814 (N_28814,N_27339,N_27983);
nand U28815 (N_28815,N_27837,N_27629);
xor U28816 (N_28816,N_27795,N_27527);
and U28817 (N_28817,N_27638,N_28434);
nand U28818 (N_28818,N_28402,N_27903);
xor U28819 (N_28819,N_27924,N_27900);
nor U28820 (N_28820,N_27673,N_27741);
nand U28821 (N_28821,N_27793,N_27101);
xnor U28822 (N_28822,N_27814,N_28026);
nor U28823 (N_28823,N_27203,N_28019);
or U28824 (N_28824,N_27865,N_27393);
nor U28825 (N_28825,N_27735,N_27371);
xor U28826 (N_28826,N_28397,N_27329);
and U28827 (N_28827,N_27280,N_27192);
xnor U28828 (N_28828,N_27525,N_27601);
and U28829 (N_28829,N_27136,N_28133);
nand U28830 (N_28830,N_27692,N_28440);
nor U28831 (N_28831,N_27374,N_27387);
nand U28832 (N_28832,N_27737,N_28056);
nor U28833 (N_28833,N_27273,N_27602);
nand U28834 (N_28834,N_28366,N_27380);
xnor U28835 (N_28835,N_28058,N_27571);
or U28836 (N_28836,N_27979,N_27728);
nor U28837 (N_28837,N_28421,N_28079);
xnor U28838 (N_28838,N_27575,N_28302);
xor U28839 (N_28839,N_28448,N_27088);
nand U28840 (N_28840,N_27243,N_28204);
nand U28841 (N_28841,N_27596,N_27162);
and U28842 (N_28842,N_27500,N_27515);
nand U28843 (N_28843,N_28108,N_27627);
xor U28844 (N_28844,N_28274,N_27928);
xor U28845 (N_28845,N_27825,N_27470);
xnor U28846 (N_28846,N_28050,N_27142);
xnor U28847 (N_28847,N_27830,N_27917);
xor U28848 (N_28848,N_27734,N_28074);
nor U28849 (N_28849,N_27361,N_27024);
or U28850 (N_28850,N_28003,N_27557);
or U28851 (N_28851,N_28422,N_28307);
nor U28852 (N_28852,N_28335,N_28037);
nor U28853 (N_28853,N_28189,N_27042);
xor U28854 (N_28854,N_28384,N_27313);
nor U28855 (N_28855,N_27415,N_27067);
and U28856 (N_28856,N_27632,N_27753);
nand U28857 (N_28857,N_27218,N_27662);
or U28858 (N_28858,N_28438,N_28406);
or U28859 (N_28859,N_28201,N_28472);
or U28860 (N_28860,N_27223,N_28446);
nand U28861 (N_28861,N_28226,N_27272);
and U28862 (N_28862,N_28419,N_27340);
nor U28863 (N_28863,N_28109,N_27553);
nor U28864 (N_28864,N_27125,N_28224);
or U28865 (N_28865,N_27109,N_28337);
and U28866 (N_28866,N_28474,N_27276);
nor U28867 (N_28867,N_28398,N_28298);
and U28868 (N_28868,N_27461,N_28236);
nand U28869 (N_28869,N_27210,N_27300);
nand U28870 (N_28870,N_27621,N_27658);
nand U28871 (N_28871,N_27044,N_27149);
nand U28872 (N_28872,N_28483,N_28285);
and U28873 (N_28873,N_27484,N_27988);
nand U28874 (N_28874,N_28161,N_27671);
and U28875 (N_28875,N_27241,N_28145);
or U28876 (N_28876,N_28424,N_27875);
nand U28877 (N_28877,N_27509,N_28193);
and U28878 (N_28878,N_27972,N_27665);
nand U28879 (N_28879,N_28124,N_28261);
or U28880 (N_28880,N_28457,N_27124);
and U28881 (N_28881,N_27738,N_28443);
nor U28882 (N_28882,N_27082,N_27787);
or U28883 (N_28883,N_27019,N_27633);
or U28884 (N_28884,N_27454,N_27151);
nand U28885 (N_28885,N_27370,N_27490);
and U28886 (N_28886,N_27169,N_28403);
or U28887 (N_28887,N_28380,N_28035);
and U28888 (N_28888,N_28205,N_28409);
xor U28889 (N_28889,N_27747,N_27229);
and U28890 (N_28890,N_27524,N_27991);
and U28891 (N_28891,N_28390,N_27133);
or U28892 (N_28892,N_27577,N_27952);
nand U28893 (N_28893,N_28118,N_27549);
nor U28894 (N_28894,N_28006,N_27699);
or U28895 (N_28895,N_27495,N_27334);
xor U28896 (N_28896,N_27794,N_27510);
xnor U28897 (N_28897,N_27906,N_27439);
nand U28898 (N_28898,N_27823,N_28372);
nand U28899 (N_28899,N_27421,N_27497);
xnor U28900 (N_28900,N_27573,N_27882);
or U28901 (N_28901,N_27250,N_27616);
xnor U28902 (N_28902,N_27382,N_27295);
and U28903 (N_28903,N_27725,N_27289);
xor U28904 (N_28904,N_27841,N_27154);
or U28905 (N_28905,N_28354,N_28117);
xor U28906 (N_28906,N_27158,N_27739);
and U28907 (N_28907,N_27800,N_27031);
xnor U28908 (N_28908,N_27220,N_27332);
xnor U28909 (N_28909,N_27521,N_27961);
and U28910 (N_28910,N_27868,N_27287);
nor U28911 (N_28911,N_27343,N_27355);
xor U28912 (N_28912,N_28282,N_27318);
xnor U28913 (N_28913,N_27829,N_27801);
nand U28914 (N_28914,N_27669,N_27076);
and U28915 (N_28915,N_27843,N_27398);
xnor U28916 (N_28916,N_28468,N_27854);
and U28917 (N_28917,N_27315,N_27464);
and U28918 (N_28918,N_27939,N_28338);
and U28919 (N_28919,N_28152,N_27150);
nor U28920 (N_28920,N_28299,N_28169);
or U28921 (N_28921,N_27863,N_28281);
xor U28922 (N_28922,N_27705,N_28289);
and U28923 (N_28923,N_27599,N_27277);
xnor U28924 (N_28924,N_28170,N_28138);
nand U28925 (N_28925,N_28346,N_27153);
or U28926 (N_28926,N_28085,N_28410);
and U28927 (N_28927,N_28100,N_27531);
or U28928 (N_28928,N_27135,N_28357);
or U28929 (N_28929,N_27949,N_27262);
or U28930 (N_28930,N_28329,N_28065);
xnor U28931 (N_28931,N_28400,N_27083);
and U28932 (N_28932,N_27395,N_27909);
and U28933 (N_28933,N_27877,N_28004);
xor U28934 (N_28934,N_27546,N_27946);
nor U28935 (N_28935,N_27144,N_27680);
and U28936 (N_28936,N_27392,N_27608);
nand U28937 (N_28937,N_27530,N_27455);
xnor U28938 (N_28938,N_28270,N_27943);
or U28939 (N_28939,N_28369,N_28111);
or U28940 (N_28940,N_27860,N_28296);
nor U28941 (N_28941,N_27619,N_27565);
xor U28942 (N_28942,N_28336,N_27038);
nor U28943 (N_28943,N_27284,N_27479);
xnor U28944 (N_28944,N_28154,N_27438);
nand U28945 (N_28945,N_27727,N_27070);
nor U28946 (N_28946,N_28265,N_27605);
nor U28947 (N_28947,N_27299,N_28120);
or U28948 (N_28948,N_27056,N_27960);
or U28949 (N_28949,N_27050,N_27654);
nand U28950 (N_28950,N_27482,N_27069);
xor U28951 (N_28951,N_28436,N_27033);
nor U28952 (N_28952,N_27369,N_28317);
nor U28953 (N_28953,N_27450,N_27543);
or U28954 (N_28954,N_27476,N_28432);
xor U28955 (N_28955,N_28148,N_28116);
and U28956 (N_28956,N_28259,N_27199);
xor U28957 (N_28957,N_27526,N_27444);
nand U28958 (N_28958,N_27819,N_28417);
and U28959 (N_28959,N_27407,N_27225);
or U28960 (N_28960,N_27003,N_27077);
nand U28961 (N_28961,N_28062,N_27259);
and U28962 (N_28962,N_27994,N_27556);
or U28963 (N_28963,N_28173,N_28435);
and U28964 (N_28964,N_27468,N_27791);
or U28965 (N_28965,N_28240,N_28212);
and U28966 (N_28966,N_27486,N_28377);
or U28967 (N_28967,N_28041,N_27567);
nor U28968 (N_28968,N_27206,N_27298);
xnor U28969 (N_28969,N_27079,N_28318);
xor U28970 (N_28970,N_27715,N_27496);
nand U28971 (N_28971,N_27540,N_27908);
nand U28972 (N_28972,N_28327,N_27007);
nor U28973 (N_28973,N_27011,N_27880);
or U28974 (N_28974,N_27238,N_28077);
or U28975 (N_28975,N_27944,N_27316);
xor U28976 (N_28976,N_27389,N_27659);
nand U28977 (N_28977,N_27110,N_27445);
nor U28978 (N_28978,N_27175,N_27561);
and U28979 (N_28979,N_27660,N_27518);
nor U28980 (N_28980,N_28242,N_28144);
or U28981 (N_28981,N_27852,N_27443);
xnor U28982 (N_28982,N_28159,N_27234);
and U28983 (N_28983,N_27539,N_27275);
or U28984 (N_28984,N_28163,N_27769);
xor U28985 (N_28985,N_27585,N_27320);
nor U28986 (N_28986,N_27749,N_27442);
and U28987 (N_28987,N_27227,N_28349);
xnor U28988 (N_28988,N_27477,N_27826);
or U28989 (N_28989,N_28275,N_27417);
xor U28990 (N_28990,N_27940,N_27338);
nand U28991 (N_28991,N_28101,N_27690);
nor U28992 (N_28992,N_27095,N_27061);
nand U28993 (N_28993,N_27505,N_27809);
and U28994 (N_28994,N_28271,N_27171);
and U28995 (N_28995,N_27198,N_27820);
and U28996 (N_28996,N_27764,N_27745);
nand U28997 (N_28997,N_27848,N_27475);
nor U28998 (N_28998,N_28325,N_27200);
nand U28999 (N_28999,N_27547,N_28067);
nor U29000 (N_29000,N_27312,N_28024);
nand U29001 (N_29001,N_28251,N_27771);
xor U29002 (N_29002,N_27402,N_28107);
and U29003 (N_29003,N_27657,N_27847);
nand U29004 (N_29004,N_27335,N_27097);
and U29005 (N_29005,N_27831,N_27085);
nand U29006 (N_29006,N_28491,N_27618);
and U29007 (N_29007,N_27925,N_27810);
or U29008 (N_29008,N_28350,N_27129);
nor U29009 (N_29009,N_28260,N_28235);
and U29010 (N_29010,N_27973,N_28102);
nor U29011 (N_29011,N_27394,N_27032);
or U29012 (N_29012,N_28253,N_27105);
nand U29013 (N_29013,N_27851,N_28376);
nand U29014 (N_29014,N_28494,N_27016);
nand U29015 (N_29015,N_27344,N_28316);
nor U29016 (N_29016,N_27304,N_28293);
and U29017 (N_29017,N_28272,N_27980);
nor U29018 (N_29018,N_28264,N_28495);
and U29019 (N_29019,N_27035,N_27457);
nand U29020 (N_29020,N_27435,N_27252);
nand U29021 (N_29021,N_27364,N_27945);
and U29022 (N_29022,N_27818,N_28256);
nand U29023 (N_29023,N_27716,N_28185);
and U29024 (N_29024,N_27487,N_27827);
nor U29025 (N_29025,N_27681,N_27803);
xor U29026 (N_29026,N_28066,N_27812);
nand U29027 (N_29027,N_28411,N_28461);
nand U29028 (N_29028,N_27194,N_28206);
or U29029 (N_29029,N_27744,N_27703);
nand U29030 (N_29030,N_27197,N_27132);
or U29031 (N_29031,N_27456,N_28069);
nand U29032 (N_29032,N_27883,N_27233);
nand U29033 (N_29033,N_27797,N_27451);
nor U29034 (N_29034,N_27321,N_27390);
or U29035 (N_29035,N_27609,N_27068);
or U29036 (N_29036,N_28228,N_28126);
or U29037 (N_29037,N_27405,N_28477);
and U29038 (N_29038,N_27503,N_28450);
and U29039 (N_29039,N_27641,N_27919);
or U29040 (N_29040,N_27155,N_27552);
nand U29041 (N_29041,N_27774,N_27887);
nor U29042 (N_29042,N_27428,N_27365);
or U29043 (N_29043,N_28239,N_27936);
or U29044 (N_29044,N_28497,N_27709);
nor U29045 (N_29045,N_27081,N_27356);
nor U29046 (N_29046,N_28480,N_28433);
nand U29047 (N_29047,N_28315,N_28356);
xnor U29048 (N_29048,N_27719,N_27396);
and U29049 (N_29049,N_27251,N_28073);
or U29050 (N_29050,N_28106,N_27006);
and U29051 (N_29051,N_27193,N_27078);
xor U29052 (N_29052,N_28490,N_27351);
or U29053 (N_29053,N_28057,N_27157);
and U29054 (N_29054,N_27606,N_27041);
or U29055 (N_29055,N_27028,N_28431);
or U29056 (N_29056,N_28426,N_28089);
and U29057 (N_29057,N_27964,N_27185);
or U29058 (N_29058,N_28211,N_27642);
nor U29059 (N_29059,N_28385,N_28114);
nor U29060 (N_29060,N_27579,N_28465);
xor U29061 (N_29061,N_27224,N_27507);
or U29062 (N_29062,N_27383,N_27066);
and U29063 (N_29063,N_27989,N_28127);
nand U29064 (N_29064,N_27916,N_28198);
or U29065 (N_29065,N_27412,N_28364);
nor U29066 (N_29066,N_27704,N_27664);
or U29067 (N_29067,N_27399,N_28321);
nand U29068 (N_29068,N_28244,N_27118);
nand U29069 (N_29069,N_28203,N_27846);
nor U29070 (N_29070,N_28231,N_28182);
nand U29071 (N_29071,N_27941,N_27896);
nand U29072 (N_29072,N_27759,N_27625);
nor U29073 (N_29073,N_27968,N_27089);
and U29074 (N_29074,N_28267,N_28052);
and U29075 (N_29075,N_27053,N_27030);
nor U29076 (N_29076,N_27647,N_28103);
and U29077 (N_29077,N_27661,N_27938);
nand U29078 (N_29078,N_28322,N_28082);
nand U29079 (N_29079,N_28286,N_27502);
xnor U29080 (N_29080,N_28064,N_28096);
and U29081 (N_29081,N_27723,N_27535);
xnor U29082 (N_29082,N_28442,N_28011);
and U29083 (N_29083,N_27098,N_27766);
nand U29084 (N_29084,N_27384,N_27710);
xnor U29085 (N_29085,N_27141,N_27650);
xor U29086 (N_29086,N_27781,N_28220);
nand U29087 (N_29087,N_27874,N_27425);
and U29088 (N_29088,N_28015,N_27872);
and U29089 (N_29089,N_27418,N_27057);
nor U29090 (N_29090,N_28444,N_28453);
nor U29091 (N_29091,N_27532,N_28252);
or U29092 (N_29092,N_27121,N_28343);
nor U29093 (N_29093,N_27721,N_27922);
nor U29094 (N_29094,N_27015,N_27511);
xor U29095 (N_29095,N_28174,N_28132);
nor U29096 (N_29096,N_28330,N_28130);
nand U29097 (N_29097,N_28091,N_27828);
and U29098 (N_29098,N_27434,N_27054);
nand U29099 (N_29099,N_27426,N_28165);
and U29100 (N_29100,N_27514,N_27345);
nor U29101 (N_29101,N_28020,N_27291);
xor U29102 (N_29102,N_27172,N_27472);
nor U29103 (N_29103,N_27261,N_27174);
or U29104 (N_29104,N_27099,N_27569);
nor U29105 (N_29105,N_27269,N_28076);
xor U29106 (N_29106,N_27063,N_27046);
or U29107 (N_29107,N_28191,N_27122);
nand U29108 (N_29108,N_27286,N_27750);
xor U29109 (N_29109,N_27839,N_28328);
and U29110 (N_29110,N_27378,N_28498);
nor U29111 (N_29111,N_28186,N_27501);
and U29112 (N_29112,N_27094,N_27429);
nand U29113 (N_29113,N_27211,N_28215);
nand U29114 (N_29114,N_27075,N_28471);
nand U29115 (N_29115,N_27578,N_27686);
nand U29116 (N_29116,N_27538,N_27222);
nand U29117 (N_29117,N_27205,N_27013);
or U29118 (N_29118,N_27784,N_28280);
xor U29119 (N_29119,N_27008,N_27506);
or U29120 (N_29120,N_28143,N_28027);
and U29121 (N_29121,N_27516,N_27967);
nor U29122 (N_29122,N_27504,N_27761);
and U29123 (N_29123,N_27742,N_27963);
or U29124 (N_29124,N_27996,N_27802);
and U29125 (N_29125,N_27469,N_27023);
xnor U29126 (N_29126,N_27920,N_27886);
xor U29127 (N_29127,N_28146,N_27000);
xor U29128 (N_29128,N_27260,N_28250);
nand U29129 (N_29129,N_27869,N_27408);
and U29130 (N_29130,N_27986,N_27542);
or U29131 (N_29131,N_27555,N_27905);
or U29132 (N_29132,N_28391,N_27026);
and U29133 (N_29133,N_28339,N_27036);
nor U29134 (N_29134,N_27976,N_28304);
and U29135 (N_29135,N_28452,N_27833);
nand U29136 (N_29136,N_28334,N_28048);
and U29137 (N_29137,N_27520,N_27702);
xnor U29138 (N_29138,N_28195,N_27274);
nor U29139 (N_29139,N_27381,N_27724);
and U29140 (N_29140,N_27228,N_27701);
and U29141 (N_29141,N_27696,N_27534);
and U29142 (N_29142,N_28386,N_27581);
nor U29143 (N_29143,N_27215,N_27695);
nor U29144 (N_29144,N_27856,N_28053);
or U29145 (N_29145,N_27237,N_27649);
xnor U29146 (N_29146,N_27519,N_27349);
nand U29147 (N_29147,N_27309,N_27646);
xnor U29148 (N_29148,N_28000,N_27614);
or U29149 (N_29149,N_28181,N_27281);
nand U29150 (N_29150,N_27307,N_27087);
nand U29151 (N_29151,N_27324,N_27176);
nand U29152 (N_29152,N_28070,N_28225);
xnor U29153 (N_29153,N_27458,N_27639);
and U29154 (N_29154,N_27207,N_28010);
nand U29155 (N_29155,N_27270,N_28086);
nand U29156 (N_29156,N_27294,N_27463);
or U29157 (N_29157,N_27005,N_27022);
nor U29158 (N_29158,N_27409,N_27603);
and U29159 (N_29159,N_27729,N_27137);
nor U29160 (N_29160,N_28347,N_28172);
or U29161 (N_29161,N_27648,N_27788);
nand U29162 (N_29162,N_27244,N_27707);
nand U29163 (N_29163,N_28128,N_27796);
and U29164 (N_29164,N_28222,N_27586);
nor U29165 (N_29165,N_27404,N_27147);
nand U29166 (N_29166,N_28012,N_28238);
nand U29167 (N_29167,N_28031,N_27301);
nor U29168 (N_29168,N_28248,N_27731);
nor U29169 (N_29169,N_27522,N_28068);
or U29170 (N_29170,N_27923,N_27574);
and U29171 (N_29171,N_27912,N_27927);
nand U29172 (N_29172,N_28312,N_27213);
and U29173 (N_29173,N_27037,N_27694);
and U29174 (N_29174,N_27437,N_27876);
or U29175 (N_29175,N_27610,N_27850);
xor U29176 (N_29176,N_27420,N_27842);
xnor U29177 (N_29177,N_27898,N_28038);
nand U29178 (N_29178,N_28392,N_27970);
nor U29179 (N_29179,N_28393,N_27904);
or U29180 (N_29180,N_27254,N_27376);
xor U29181 (N_29181,N_28192,N_28016);
xnor U29182 (N_29182,N_28476,N_28297);
or U29183 (N_29183,N_28160,N_27386);
xor U29184 (N_29184,N_28007,N_27808);
nor U29185 (N_29185,N_27685,N_28378);
and U29186 (N_29186,N_28414,N_28454);
and U29187 (N_29187,N_27242,N_28269);
nor U29188 (N_29188,N_27474,N_27732);
nand U29189 (N_29189,N_27377,N_27148);
or U29190 (N_29190,N_28072,N_28273);
nand U29191 (N_29191,N_28324,N_27314);
and U29192 (N_29192,N_27403,N_28097);
nor U29193 (N_29193,N_28018,N_27806);
nor U29194 (N_29194,N_27558,N_27600);
or U29195 (N_29195,N_27559,N_28394);
nor U29196 (N_29196,N_28140,N_27323);
nand U29197 (N_29197,N_27191,N_27926);
nor U29198 (N_29198,N_27302,N_27765);
or U29199 (N_29199,N_28093,N_27566);
nor U29200 (N_29200,N_28305,N_27423);
xnor U29201 (N_29201,N_27212,N_28368);
and U29202 (N_29202,N_27379,N_27331);
xor U29203 (N_29203,N_28475,N_27292);
or U29204 (N_29204,N_27115,N_27433);
or U29205 (N_29205,N_27748,N_27480);
and U29206 (N_29206,N_27762,N_27163);
xor U29207 (N_29207,N_27071,N_27467);
xor U29208 (N_29208,N_27074,N_27048);
or U29209 (N_29209,N_28125,N_28301);
or U29210 (N_29210,N_27267,N_27620);
and U29211 (N_29211,N_28036,N_27687);
xor U29212 (N_29212,N_28005,N_28162);
or U29213 (N_29213,N_28295,N_28294);
xor U29214 (N_29214,N_27184,N_27935);
or U29215 (N_29215,N_28021,N_28258);
xor U29216 (N_29216,N_27453,N_27537);
nand U29217 (N_29217,N_27902,N_27529);
and U29218 (N_29218,N_27305,N_28255);
nand U29219 (N_29219,N_28277,N_27736);
or U29220 (N_29220,N_27545,N_27612);
and U29221 (N_29221,N_28059,N_28131);
xor U29222 (N_29222,N_28237,N_27130);
nor U29223 (N_29223,N_27165,N_27604);
or U29224 (N_29224,N_28039,N_27388);
nand U29225 (N_29225,N_28479,N_27777);
nor U29226 (N_29226,N_27362,N_27626);
nand U29227 (N_29227,N_27108,N_28467);
and U29228 (N_29228,N_27446,N_27910);
and U29229 (N_29229,N_27541,N_28367);
or U29230 (N_29230,N_28197,N_27440);
nor U29231 (N_29231,N_27427,N_28257);
or U29232 (N_29232,N_27119,N_28104);
nand U29233 (N_29233,N_27120,N_28087);
and U29234 (N_29234,N_27416,N_28287);
and U29235 (N_29235,N_27591,N_27020);
nand U29236 (N_29236,N_27092,N_27248);
and U29237 (N_29237,N_27953,N_27065);
xor U29238 (N_29238,N_27958,N_28040);
xor U29239 (N_29239,N_27959,N_27460);
nor U29240 (N_29240,N_28486,N_27667);
nand U29241 (N_29241,N_27265,N_28365);
nor U29242 (N_29242,N_28249,N_27849);
or U29243 (N_29243,N_27025,N_28017);
nand U29244 (N_29244,N_27128,N_27597);
xnor U29245 (N_29245,N_28395,N_27583);
xnor U29246 (N_29246,N_27563,N_27512);
nand U29247 (N_29247,N_27730,N_27640);
and U29248 (N_29248,N_27811,N_27698);
nor U29249 (N_29249,N_28151,N_27992);
nand U29250 (N_29250,N_27937,N_27045);
nand U29251 (N_29251,N_27556,N_27895);
and U29252 (N_29252,N_28489,N_27960);
and U29253 (N_29253,N_27604,N_28269);
or U29254 (N_29254,N_28121,N_28255);
nand U29255 (N_29255,N_28128,N_28054);
nor U29256 (N_29256,N_28408,N_28033);
nor U29257 (N_29257,N_27549,N_27336);
and U29258 (N_29258,N_28086,N_27882);
or U29259 (N_29259,N_28455,N_28233);
nor U29260 (N_29260,N_28222,N_28469);
and U29261 (N_29261,N_27243,N_27188);
and U29262 (N_29262,N_27551,N_27258);
xor U29263 (N_29263,N_27738,N_28411);
xnor U29264 (N_29264,N_27500,N_27602);
and U29265 (N_29265,N_27787,N_27835);
nor U29266 (N_29266,N_27213,N_27580);
or U29267 (N_29267,N_27793,N_27461);
nand U29268 (N_29268,N_27487,N_27261);
and U29269 (N_29269,N_28025,N_28173);
nor U29270 (N_29270,N_27074,N_28424);
nor U29271 (N_29271,N_27725,N_27240);
xor U29272 (N_29272,N_27249,N_27718);
or U29273 (N_29273,N_27181,N_27757);
or U29274 (N_29274,N_28321,N_28410);
xor U29275 (N_29275,N_28085,N_28263);
nor U29276 (N_29276,N_27073,N_28499);
nor U29277 (N_29277,N_27071,N_27644);
nor U29278 (N_29278,N_27640,N_27596);
or U29279 (N_29279,N_27968,N_27803);
and U29280 (N_29280,N_28161,N_28091);
or U29281 (N_29281,N_28198,N_27881);
xnor U29282 (N_29282,N_27565,N_28268);
or U29283 (N_29283,N_27481,N_28098);
and U29284 (N_29284,N_27799,N_27552);
nand U29285 (N_29285,N_27844,N_27203);
nand U29286 (N_29286,N_27904,N_27154);
or U29287 (N_29287,N_27044,N_28284);
nand U29288 (N_29288,N_28338,N_28064);
nand U29289 (N_29289,N_28006,N_28287);
or U29290 (N_29290,N_27929,N_28405);
nor U29291 (N_29291,N_27319,N_27276);
nor U29292 (N_29292,N_27027,N_28025);
xor U29293 (N_29293,N_28368,N_27963);
or U29294 (N_29294,N_27925,N_28459);
or U29295 (N_29295,N_27645,N_27512);
and U29296 (N_29296,N_28483,N_27106);
or U29297 (N_29297,N_28194,N_28188);
and U29298 (N_29298,N_28234,N_28085);
and U29299 (N_29299,N_28318,N_28203);
nand U29300 (N_29300,N_28097,N_27678);
xor U29301 (N_29301,N_27636,N_28235);
nor U29302 (N_29302,N_27900,N_27095);
nor U29303 (N_29303,N_28469,N_28340);
nand U29304 (N_29304,N_27551,N_27461);
nand U29305 (N_29305,N_27301,N_27733);
and U29306 (N_29306,N_27826,N_27358);
xnor U29307 (N_29307,N_27990,N_27162);
xor U29308 (N_29308,N_27390,N_27597);
nand U29309 (N_29309,N_27491,N_27095);
nand U29310 (N_29310,N_27521,N_27018);
xor U29311 (N_29311,N_28087,N_28049);
or U29312 (N_29312,N_27945,N_27095);
xnor U29313 (N_29313,N_27370,N_28291);
nand U29314 (N_29314,N_27298,N_27519);
nor U29315 (N_29315,N_28136,N_28230);
nand U29316 (N_29316,N_27070,N_28229);
nor U29317 (N_29317,N_28099,N_27877);
xnor U29318 (N_29318,N_27507,N_27059);
or U29319 (N_29319,N_27509,N_27529);
xnor U29320 (N_29320,N_27670,N_27654);
or U29321 (N_29321,N_27248,N_27379);
or U29322 (N_29322,N_27802,N_28074);
and U29323 (N_29323,N_27940,N_27907);
xor U29324 (N_29324,N_27059,N_28468);
nand U29325 (N_29325,N_28441,N_28110);
nand U29326 (N_29326,N_27211,N_27624);
nand U29327 (N_29327,N_27140,N_27303);
or U29328 (N_29328,N_27277,N_27486);
or U29329 (N_29329,N_27628,N_27747);
nor U29330 (N_29330,N_27542,N_28105);
and U29331 (N_29331,N_27985,N_27099);
and U29332 (N_29332,N_28001,N_27034);
nand U29333 (N_29333,N_28020,N_27334);
and U29334 (N_29334,N_27981,N_27173);
and U29335 (N_29335,N_27737,N_28103);
nand U29336 (N_29336,N_27567,N_28334);
xor U29337 (N_29337,N_28097,N_28383);
xnor U29338 (N_29338,N_28482,N_28316);
and U29339 (N_29339,N_27996,N_28451);
nand U29340 (N_29340,N_27899,N_28183);
xnor U29341 (N_29341,N_27941,N_27834);
or U29342 (N_29342,N_27541,N_27952);
nand U29343 (N_29343,N_27957,N_28438);
nand U29344 (N_29344,N_28038,N_27045);
xnor U29345 (N_29345,N_27199,N_27066);
nor U29346 (N_29346,N_28204,N_27115);
nand U29347 (N_29347,N_27059,N_27030);
or U29348 (N_29348,N_27649,N_27501);
nor U29349 (N_29349,N_27834,N_28145);
or U29350 (N_29350,N_28017,N_27680);
xnor U29351 (N_29351,N_27906,N_27256);
xor U29352 (N_29352,N_27850,N_27426);
nor U29353 (N_29353,N_27164,N_27944);
xnor U29354 (N_29354,N_28367,N_28481);
xor U29355 (N_29355,N_27962,N_27451);
nand U29356 (N_29356,N_27640,N_27019);
nand U29357 (N_29357,N_28190,N_27306);
xor U29358 (N_29358,N_27655,N_27660);
nor U29359 (N_29359,N_27659,N_28080);
or U29360 (N_29360,N_27968,N_28168);
xor U29361 (N_29361,N_27513,N_27290);
xnor U29362 (N_29362,N_27819,N_28238);
xor U29363 (N_29363,N_27544,N_28305);
or U29364 (N_29364,N_27046,N_27425);
or U29365 (N_29365,N_28365,N_27727);
nor U29366 (N_29366,N_27370,N_28167);
or U29367 (N_29367,N_28069,N_27448);
and U29368 (N_29368,N_27107,N_27048);
nor U29369 (N_29369,N_27758,N_28318);
and U29370 (N_29370,N_27733,N_28469);
nand U29371 (N_29371,N_27312,N_27863);
and U29372 (N_29372,N_27880,N_28098);
xor U29373 (N_29373,N_27545,N_28492);
xnor U29374 (N_29374,N_27307,N_28492);
nor U29375 (N_29375,N_27957,N_27229);
or U29376 (N_29376,N_28254,N_27695);
xor U29377 (N_29377,N_28377,N_27772);
or U29378 (N_29378,N_27022,N_27858);
nand U29379 (N_29379,N_28294,N_27521);
or U29380 (N_29380,N_27760,N_27147);
or U29381 (N_29381,N_27487,N_27375);
xor U29382 (N_29382,N_28014,N_27416);
and U29383 (N_29383,N_27191,N_27104);
nand U29384 (N_29384,N_28422,N_27564);
nand U29385 (N_29385,N_28163,N_27410);
nor U29386 (N_29386,N_28206,N_27704);
nor U29387 (N_29387,N_28240,N_27094);
nor U29388 (N_29388,N_27355,N_27198);
or U29389 (N_29389,N_27787,N_28492);
nand U29390 (N_29390,N_27622,N_27204);
xor U29391 (N_29391,N_27922,N_27388);
xor U29392 (N_29392,N_27093,N_27653);
and U29393 (N_29393,N_28419,N_27714);
nand U29394 (N_29394,N_27718,N_28153);
and U29395 (N_29395,N_27886,N_27685);
and U29396 (N_29396,N_27265,N_27506);
and U29397 (N_29397,N_27249,N_27242);
nand U29398 (N_29398,N_28180,N_27246);
and U29399 (N_29399,N_27490,N_27735);
and U29400 (N_29400,N_27693,N_27213);
nor U29401 (N_29401,N_27037,N_27902);
nand U29402 (N_29402,N_28467,N_27760);
or U29403 (N_29403,N_27201,N_27512);
and U29404 (N_29404,N_27054,N_27887);
or U29405 (N_29405,N_27304,N_28285);
xor U29406 (N_29406,N_27016,N_28460);
nand U29407 (N_29407,N_27501,N_27887);
nand U29408 (N_29408,N_27081,N_28262);
and U29409 (N_29409,N_27073,N_28151);
or U29410 (N_29410,N_28476,N_27514);
xor U29411 (N_29411,N_28152,N_27111);
nand U29412 (N_29412,N_28096,N_27555);
nand U29413 (N_29413,N_27805,N_27549);
and U29414 (N_29414,N_28396,N_28259);
or U29415 (N_29415,N_28058,N_28293);
and U29416 (N_29416,N_27617,N_27227);
or U29417 (N_29417,N_27360,N_27236);
or U29418 (N_29418,N_27075,N_27877);
and U29419 (N_29419,N_27911,N_27616);
xor U29420 (N_29420,N_28127,N_27546);
or U29421 (N_29421,N_28224,N_27285);
and U29422 (N_29422,N_28343,N_27947);
xnor U29423 (N_29423,N_27249,N_27575);
nor U29424 (N_29424,N_28064,N_27575);
or U29425 (N_29425,N_28158,N_28098);
or U29426 (N_29426,N_28379,N_27282);
nand U29427 (N_29427,N_28499,N_28478);
nor U29428 (N_29428,N_27496,N_27459);
nand U29429 (N_29429,N_27019,N_28369);
nor U29430 (N_29430,N_27420,N_27312);
and U29431 (N_29431,N_28404,N_28391);
nand U29432 (N_29432,N_28148,N_28486);
nand U29433 (N_29433,N_27312,N_27076);
or U29434 (N_29434,N_27363,N_28147);
and U29435 (N_29435,N_27484,N_28433);
nor U29436 (N_29436,N_28485,N_27053);
and U29437 (N_29437,N_27024,N_27544);
nor U29438 (N_29438,N_27186,N_27019);
xor U29439 (N_29439,N_28375,N_27200);
and U29440 (N_29440,N_28284,N_27128);
and U29441 (N_29441,N_27569,N_27948);
or U29442 (N_29442,N_28464,N_27431);
xnor U29443 (N_29443,N_27694,N_27724);
nor U29444 (N_29444,N_28294,N_28079);
xor U29445 (N_29445,N_27292,N_27642);
and U29446 (N_29446,N_28471,N_28284);
and U29447 (N_29447,N_28359,N_27257);
xnor U29448 (N_29448,N_27830,N_27473);
nand U29449 (N_29449,N_27282,N_27337);
and U29450 (N_29450,N_28055,N_27892);
or U29451 (N_29451,N_27442,N_27620);
or U29452 (N_29452,N_27019,N_27566);
or U29453 (N_29453,N_27902,N_28490);
nor U29454 (N_29454,N_27778,N_28471);
nor U29455 (N_29455,N_27482,N_28211);
and U29456 (N_29456,N_27726,N_28011);
or U29457 (N_29457,N_28226,N_28405);
xnor U29458 (N_29458,N_28325,N_27756);
and U29459 (N_29459,N_27389,N_27053);
and U29460 (N_29460,N_27384,N_27150);
nor U29461 (N_29461,N_27825,N_28036);
nor U29462 (N_29462,N_28096,N_27150);
nor U29463 (N_29463,N_27387,N_27155);
and U29464 (N_29464,N_28184,N_27199);
or U29465 (N_29465,N_27256,N_27246);
xor U29466 (N_29466,N_27253,N_28240);
and U29467 (N_29467,N_27215,N_27378);
nand U29468 (N_29468,N_27161,N_27452);
nand U29469 (N_29469,N_28273,N_28439);
xnor U29470 (N_29470,N_27400,N_27179);
nand U29471 (N_29471,N_28290,N_28031);
nor U29472 (N_29472,N_27711,N_27734);
or U29473 (N_29473,N_28345,N_27000);
nor U29474 (N_29474,N_28491,N_28121);
nand U29475 (N_29475,N_27615,N_28340);
or U29476 (N_29476,N_27086,N_27990);
or U29477 (N_29477,N_27365,N_27383);
xnor U29478 (N_29478,N_28320,N_28430);
and U29479 (N_29479,N_27822,N_27872);
or U29480 (N_29480,N_27502,N_28255);
and U29481 (N_29481,N_27113,N_27994);
xor U29482 (N_29482,N_27756,N_27065);
nor U29483 (N_29483,N_27851,N_27487);
and U29484 (N_29484,N_28445,N_27291);
nor U29485 (N_29485,N_28497,N_27083);
xnor U29486 (N_29486,N_27871,N_27326);
or U29487 (N_29487,N_28482,N_27212);
and U29488 (N_29488,N_28482,N_28013);
xnor U29489 (N_29489,N_28167,N_28233);
nor U29490 (N_29490,N_27932,N_27170);
nor U29491 (N_29491,N_27111,N_27635);
xnor U29492 (N_29492,N_27600,N_27753);
nor U29493 (N_29493,N_28147,N_27810);
nor U29494 (N_29494,N_28042,N_28260);
nor U29495 (N_29495,N_27137,N_27132);
or U29496 (N_29496,N_27868,N_27394);
or U29497 (N_29497,N_27245,N_28292);
nand U29498 (N_29498,N_28034,N_27806);
nor U29499 (N_29499,N_27913,N_27708);
and U29500 (N_29500,N_27476,N_27436);
xor U29501 (N_29501,N_27111,N_27271);
xnor U29502 (N_29502,N_27307,N_28222);
or U29503 (N_29503,N_27774,N_27643);
xnor U29504 (N_29504,N_27108,N_27456);
or U29505 (N_29505,N_27807,N_27912);
or U29506 (N_29506,N_28195,N_27863);
xor U29507 (N_29507,N_27013,N_27829);
nand U29508 (N_29508,N_27276,N_28258);
xor U29509 (N_29509,N_27687,N_27707);
nor U29510 (N_29510,N_27691,N_28438);
nand U29511 (N_29511,N_27953,N_27053);
nor U29512 (N_29512,N_27691,N_28375);
and U29513 (N_29513,N_27115,N_27231);
nand U29514 (N_29514,N_27695,N_28322);
or U29515 (N_29515,N_27179,N_28169);
and U29516 (N_29516,N_28153,N_28075);
nand U29517 (N_29517,N_27257,N_28360);
xnor U29518 (N_29518,N_27254,N_27910);
nand U29519 (N_29519,N_28014,N_27958);
nand U29520 (N_29520,N_28152,N_28366);
or U29521 (N_29521,N_27502,N_28303);
or U29522 (N_29522,N_27801,N_27509);
nor U29523 (N_29523,N_28480,N_27902);
nor U29524 (N_29524,N_27255,N_27488);
or U29525 (N_29525,N_27015,N_27673);
nand U29526 (N_29526,N_27711,N_27911);
or U29527 (N_29527,N_27011,N_27095);
nand U29528 (N_29528,N_27401,N_27572);
xor U29529 (N_29529,N_27491,N_27031);
and U29530 (N_29530,N_27661,N_27698);
xnor U29531 (N_29531,N_27782,N_28228);
nor U29532 (N_29532,N_27169,N_27271);
xor U29533 (N_29533,N_28324,N_27025);
xnor U29534 (N_29534,N_28398,N_28244);
nor U29535 (N_29535,N_27297,N_27708);
nor U29536 (N_29536,N_27073,N_27242);
or U29537 (N_29537,N_28268,N_27626);
nor U29538 (N_29538,N_28197,N_27643);
nand U29539 (N_29539,N_27369,N_27322);
nor U29540 (N_29540,N_27627,N_27054);
nor U29541 (N_29541,N_28298,N_28097);
nor U29542 (N_29542,N_27374,N_27654);
nand U29543 (N_29543,N_27481,N_28208);
nand U29544 (N_29544,N_28318,N_27083);
or U29545 (N_29545,N_27429,N_28347);
nand U29546 (N_29546,N_28171,N_28300);
or U29547 (N_29547,N_27712,N_28034);
xnor U29548 (N_29548,N_28245,N_27658);
and U29549 (N_29549,N_28273,N_28124);
or U29550 (N_29550,N_28179,N_27514);
or U29551 (N_29551,N_27177,N_27926);
nor U29552 (N_29552,N_27952,N_27830);
and U29553 (N_29553,N_28476,N_27959);
or U29554 (N_29554,N_28085,N_28384);
nand U29555 (N_29555,N_27455,N_27404);
nor U29556 (N_29556,N_27223,N_27500);
xor U29557 (N_29557,N_27327,N_27883);
nand U29558 (N_29558,N_27684,N_27260);
and U29559 (N_29559,N_27212,N_28457);
or U29560 (N_29560,N_27866,N_28175);
xor U29561 (N_29561,N_28280,N_27907);
nor U29562 (N_29562,N_27726,N_28361);
or U29563 (N_29563,N_27307,N_27187);
nand U29564 (N_29564,N_28185,N_27746);
nand U29565 (N_29565,N_28208,N_28310);
and U29566 (N_29566,N_27079,N_28477);
nor U29567 (N_29567,N_28150,N_27268);
and U29568 (N_29568,N_28268,N_28192);
and U29569 (N_29569,N_27541,N_27020);
and U29570 (N_29570,N_28282,N_27619);
nor U29571 (N_29571,N_28239,N_27569);
or U29572 (N_29572,N_28490,N_27907);
or U29573 (N_29573,N_27091,N_27696);
nand U29574 (N_29574,N_27830,N_27692);
and U29575 (N_29575,N_27827,N_27355);
nand U29576 (N_29576,N_27574,N_27874);
nand U29577 (N_29577,N_27484,N_27329);
or U29578 (N_29578,N_28022,N_27661);
xnor U29579 (N_29579,N_27671,N_27004);
xnor U29580 (N_29580,N_27511,N_27988);
nand U29581 (N_29581,N_27950,N_27835);
nor U29582 (N_29582,N_27043,N_28345);
xnor U29583 (N_29583,N_27608,N_28228);
xnor U29584 (N_29584,N_28378,N_27686);
nor U29585 (N_29585,N_27971,N_28439);
nor U29586 (N_29586,N_27365,N_27691);
nand U29587 (N_29587,N_28351,N_27702);
nand U29588 (N_29588,N_27333,N_28199);
nor U29589 (N_29589,N_28396,N_27869);
or U29590 (N_29590,N_27547,N_28263);
xnor U29591 (N_29591,N_27183,N_27557);
xor U29592 (N_29592,N_28287,N_28381);
xnor U29593 (N_29593,N_27168,N_27410);
xor U29594 (N_29594,N_27629,N_28366);
xor U29595 (N_29595,N_27619,N_28072);
or U29596 (N_29596,N_28394,N_27912);
nor U29597 (N_29597,N_27417,N_27800);
or U29598 (N_29598,N_27027,N_28161);
nand U29599 (N_29599,N_28165,N_28246);
and U29600 (N_29600,N_27296,N_28155);
or U29601 (N_29601,N_27541,N_27821);
or U29602 (N_29602,N_27951,N_27849);
nand U29603 (N_29603,N_27986,N_27888);
and U29604 (N_29604,N_27885,N_27598);
nand U29605 (N_29605,N_27178,N_27624);
xnor U29606 (N_29606,N_27390,N_28119);
or U29607 (N_29607,N_28238,N_28076);
and U29608 (N_29608,N_27220,N_27557);
nand U29609 (N_29609,N_27965,N_28480);
and U29610 (N_29610,N_28258,N_27693);
and U29611 (N_29611,N_27805,N_27651);
xor U29612 (N_29612,N_27761,N_28452);
nor U29613 (N_29613,N_27844,N_27419);
nand U29614 (N_29614,N_27290,N_28148);
and U29615 (N_29615,N_27732,N_28053);
xor U29616 (N_29616,N_28093,N_28091);
and U29617 (N_29617,N_27673,N_27648);
and U29618 (N_29618,N_28295,N_28293);
and U29619 (N_29619,N_28169,N_27355);
nand U29620 (N_29620,N_27352,N_27599);
nor U29621 (N_29621,N_28465,N_27639);
and U29622 (N_29622,N_27038,N_28089);
and U29623 (N_29623,N_27096,N_28383);
nand U29624 (N_29624,N_28293,N_27872);
or U29625 (N_29625,N_27096,N_28079);
or U29626 (N_29626,N_27896,N_27863);
nor U29627 (N_29627,N_27435,N_28270);
and U29628 (N_29628,N_27263,N_28209);
nor U29629 (N_29629,N_27846,N_28248);
and U29630 (N_29630,N_27657,N_27520);
xnor U29631 (N_29631,N_27105,N_27205);
nand U29632 (N_29632,N_28168,N_28124);
nor U29633 (N_29633,N_27995,N_28317);
xor U29634 (N_29634,N_28334,N_27548);
nor U29635 (N_29635,N_28265,N_27201);
and U29636 (N_29636,N_27645,N_27592);
and U29637 (N_29637,N_28029,N_27942);
and U29638 (N_29638,N_27274,N_27595);
and U29639 (N_29639,N_28333,N_28123);
xor U29640 (N_29640,N_27275,N_28400);
nor U29641 (N_29641,N_27503,N_27786);
and U29642 (N_29642,N_28232,N_27242);
and U29643 (N_29643,N_27999,N_27861);
and U29644 (N_29644,N_27570,N_28135);
nand U29645 (N_29645,N_28428,N_27354);
and U29646 (N_29646,N_27750,N_27684);
xor U29647 (N_29647,N_28265,N_28130);
nor U29648 (N_29648,N_27741,N_27066);
nand U29649 (N_29649,N_28371,N_28378);
xor U29650 (N_29650,N_27634,N_27710);
xnor U29651 (N_29651,N_27364,N_27172);
nand U29652 (N_29652,N_27292,N_28461);
and U29653 (N_29653,N_27585,N_27538);
or U29654 (N_29654,N_27133,N_27362);
xor U29655 (N_29655,N_28016,N_28103);
nand U29656 (N_29656,N_27980,N_27355);
xor U29657 (N_29657,N_27749,N_27380);
and U29658 (N_29658,N_27951,N_28238);
nor U29659 (N_29659,N_27235,N_27199);
or U29660 (N_29660,N_28433,N_27505);
or U29661 (N_29661,N_28056,N_28448);
xnor U29662 (N_29662,N_28224,N_28408);
nor U29663 (N_29663,N_27273,N_28478);
and U29664 (N_29664,N_28341,N_28111);
nor U29665 (N_29665,N_27089,N_27558);
xor U29666 (N_29666,N_27635,N_27468);
and U29667 (N_29667,N_27278,N_27616);
and U29668 (N_29668,N_28131,N_28082);
nand U29669 (N_29669,N_27282,N_28333);
or U29670 (N_29670,N_28136,N_28296);
and U29671 (N_29671,N_27384,N_28130);
nand U29672 (N_29672,N_27067,N_27823);
xnor U29673 (N_29673,N_28164,N_27912);
nor U29674 (N_29674,N_27589,N_27080);
nand U29675 (N_29675,N_27556,N_27420);
nand U29676 (N_29676,N_27097,N_27475);
nand U29677 (N_29677,N_27831,N_27042);
and U29678 (N_29678,N_27331,N_27857);
and U29679 (N_29679,N_27456,N_28141);
nand U29680 (N_29680,N_27058,N_28491);
xnor U29681 (N_29681,N_28457,N_27134);
xnor U29682 (N_29682,N_28385,N_27796);
and U29683 (N_29683,N_27756,N_28444);
xnor U29684 (N_29684,N_28116,N_27144);
or U29685 (N_29685,N_27220,N_28163);
xnor U29686 (N_29686,N_27426,N_27776);
and U29687 (N_29687,N_28107,N_27586);
nand U29688 (N_29688,N_28013,N_27819);
and U29689 (N_29689,N_28434,N_27902);
nor U29690 (N_29690,N_27506,N_27597);
or U29691 (N_29691,N_27327,N_27064);
nor U29692 (N_29692,N_27759,N_27839);
or U29693 (N_29693,N_27038,N_27445);
xor U29694 (N_29694,N_27649,N_27048);
xnor U29695 (N_29695,N_28473,N_27190);
nand U29696 (N_29696,N_28271,N_28376);
xnor U29697 (N_29697,N_28060,N_28355);
xor U29698 (N_29698,N_27691,N_27500);
nand U29699 (N_29699,N_27277,N_27171);
or U29700 (N_29700,N_28170,N_27283);
or U29701 (N_29701,N_27724,N_27312);
xor U29702 (N_29702,N_27563,N_27183);
or U29703 (N_29703,N_27145,N_28309);
xor U29704 (N_29704,N_27003,N_27415);
or U29705 (N_29705,N_27427,N_28365);
nor U29706 (N_29706,N_28055,N_27943);
nand U29707 (N_29707,N_28165,N_27674);
and U29708 (N_29708,N_28236,N_27850);
nor U29709 (N_29709,N_27528,N_28107);
nand U29710 (N_29710,N_27137,N_28153);
and U29711 (N_29711,N_27011,N_27182);
nand U29712 (N_29712,N_27807,N_28155);
nand U29713 (N_29713,N_27237,N_28136);
or U29714 (N_29714,N_27572,N_28238);
nor U29715 (N_29715,N_28422,N_28131);
xor U29716 (N_29716,N_27559,N_27773);
nand U29717 (N_29717,N_27436,N_27503);
nand U29718 (N_29718,N_27701,N_27574);
nand U29719 (N_29719,N_27281,N_27819);
nand U29720 (N_29720,N_27850,N_27714);
and U29721 (N_29721,N_27677,N_27050);
nor U29722 (N_29722,N_28073,N_27944);
nor U29723 (N_29723,N_28067,N_27760);
and U29724 (N_29724,N_28401,N_27670);
xnor U29725 (N_29725,N_27830,N_27390);
or U29726 (N_29726,N_27360,N_27280);
nor U29727 (N_29727,N_27092,N_28069);
xor U29728 (N_29728,N_27479,N_27368);
and U29729 (N_29729,N_27418,N_28144);
nor U29730 (N_29730,N_28082,N_27938);
or U29731 (N_29731,N_27230,N_27023);
or U29732 (N_29732,N_27276,N_27342);
and U29733 (N_29733,N_27884,N_27477);
nor U29734 (N_29734,N_28417,N_28259);
or U29735 (N_29735,N_27935,N_28134);
nand U29736 (N_29736,N_27645,N_28008);
or U29737 (N_29737,N_27948,N_28175);
xor U29738 (N_29738,N_27815,N_27056);
xor U29739 (N_29739,N_28396,N_27460);
and U29740 (N_29740,N_27201,N_28297);
nor U29741 (N_29741,N_28286,N_27776);
nor U29742 (N_29742,N_28199,N_28143);
nand U29743 (N_29743,N_27474,N_27536);
and U29744 (N_29744,N_27347,N_27277);
nand U29745 (N_29745,N_28288,N_27769);
xnor U29746 (N_29746,N_27415,N_27058);
nand U29747 (N_29747,N_28330,N_28388);
or U29748 (N_29748,N_27208,N_27900);
nor U29749 (N_29749,N_28481,N_27566);
nor U29750 (N_29750,N_27017,N_28288);
xor U29751 (N_29751,N_28133,N_27648);
nor U29752 (N_29752,N_27020,N_28340);
nand U29753 (N_29753,N_28087,N_28263);
nor U29754 (N_29754,N_27942,N_27236);
and U29755 (N_29755,N_28256,N_28129);
xor U29756 (N_29756,N_27256,N_27559);
or U29757 (N_29757,N_27544,N_27770);
nand U29758 (N_29758,N_27362,N_27861);
or U29759 (N_29759,N_27041,N_27314);
xor U29760 (N_29760,N_27288,N_27679);
xor U29761 (N_29761,N_28342,N_27575);
nand U29762 (N_29762,N_28432,N_28375);
and U29763 (N_29763,N_28431,N_28217);
and U29764 (N_29764,N_27576,N_27419);
nor U29765 (N_29765,N_27267,N_28049);
or U29766 (N_29766,N_27917,N_27743);
nand U29767 (N_29767,N_27991,N_27111);
xnor U29768 (N_29768,N_27847,N_28232);
nand U29769 (N_29769,N_27918,N_27358);
or U29770 (N_29770,N_27112,N_27830);
nand U29771 (N_29771,N_28423,N_27127);
nor U29772 (N_29772,N_28188,N_28495);
nor U29773 (N_29773,N_28310,N_27000);
and U29774 (N_29774,N_27978,N_28025);
or U29775 (N_29775,N_27092,N_28311);
and U29776 (N_29776,N_27263,N_28435);
xnor U29777 (N_29777,N_28450,N_27862);
and U29778 (N_29778,N_28219,N_28406);
and U29779 (N_29779,N_27938,N_27675);
nand U29780 (N_29780,N_28466,N_27808);
nor U29781 (N_29781,N_27315,N_27211);
xnor U29782 (N_29782,N_27044,N_27438);
nor U29783 (N_29783,N_27937,N_27766);
and U29784 (N_29784,N_27920,N_27677);
or U29785 (N_29785,N_27282,N_28429);
nor U29786 (N_29786,N_28074,N_27230);
nand U29787 (N_29787,N_28013,N_28228);
or U29788 (N_29788,N_28347,N_27277);
or U29789 (N_29789,N_28056,N_27825);
and U29790 (N_29790,N_27508,N_28368);
and U29791 (N_29791,N_27324,N_27635);
xnor U29792 (N_29792,N_28380,N_28447);
nor U29793 (N_29793,N_27165,N_27260);
and U29794 (N_29794,N_28407,N_27427);
or U29795 (N_29795,N_27449,N_28440);
nor U29796 (N_29796,N_27428,N_28330);
nand U29797 (N_29797,N_28060,N_28026);
nand U29798 (N_29798,N_28120,N_27216);
xor U29799 (N_29799,N_28335,N_27596);
nand U29800 (N_29800,N_27764,N_27829);
nor U29801 (N_29801,N_27126,N_28414);
nor U29802 (N_29802,N_27275,N_27822);
and U29803 (N_29803,N_27590,N_27346);
or U29804 (N_29804,N_28297,N_27324);
nor U29805 (N_29805,N_27318,N_28469);
nor U29806 (N_29806,N_28428,N_28349);
nor U29807 (N_29807,N_28185,N_27433);
and U29808 (N_29808,N_28052,N_27904);
nor U29809 (N_29809,N_28230,N_27052);
or U29810 (N_29810,N_27506,N_28205);
or U29811 (N_29811,N_27798,N_27574);
nor U29812 (N_29812,N_27630,N_28086);
nor U29813 (N_29813,N_27179,N_27046);
nand U29814 (N_29814,N_28354,N_28375);
nor U29815 (N_29815,N_27459,N_27258);
xnor U29816 (N_29816,N_27084,N_27611);
nand U29817 (N_29817,N_27954,N_27614);
nand U29818 (N_29818,N_28169,N_27954);
xnor U29819 (N_29819,N_27950,N_27579);
xor U29820 (N_29820,N_28489,N_28243);
and U29821 (N_29821,N_28367,N_27017);
and U29822 (N_29822,N_27243,N_27720);
and U29823 (N_29823,N_28146,N_28314);
xnor U29824 (N_29824,N_28289,N_28209);
and U29825 (N_29825,N_28159,N_28372);
and U29826 (N_29826,N_28020,N_27618);
or U29827 (N_29827,N_27210,N_27920);
xor U29828 (N_29828,N_27746,N_27686);
or U29829 (N_29829,N_27608,N_27374);
xnor U29830 (N_29830,N_27376,N_27908);
nand U29831 (N_29831,N_28127,N_28455);
xnor U29832 (N_29832,N_27330,N_28016);
or U29833 (N_29833,N_27510,N_28003);
or U29834 (N_29834,N_28053,N_27057);
nor U29835 (N_29835,N_27095,N_28474);
nand U29836 (N_29836,N_27216,N_27838);
or U29837 (N_29837,N_28145,N_28025);
and U29838 (N_29838,N_27872,N_28021);
or U29839 (N_29839,N_27142,N_27683);
nand U29840 (N_29840,N_28004,N_28428);
nor U29841 (N_29841,N_27594,N_27112);
or U29842 (N_29842,N_27946,N_28048);
xnor U29843 (N_29843,N_27501,N_28027);
nand U29844 (N_29844,N_27883,N_27661);
xnor U29845 (N_29845,N_28112,N_27220);
xor U29846 (N_29846,N_27867,N_28054);
xor U29847 (N_29847,N_27426,N_27230);
or U29848 (N_29848,N_28252,N_27800);
xnor U29849 (N_29849,N_27296,N_27396);
or U29850 (N_29850,N_27227,N_27534);
and U29851 (N_29851,N_28079,N_28182);
nor U29852 (N_29852,N_27203,N_28039);
or U29853 (N_29853,N_28251,N_28370);
nor U29854 (N_29854,N_27616,N_27826);
xor U29855 (N_29855,N_27913,N_27780);
xor U29856 (N_29856,N_28254,N_27070);
and U29857 (N_29857,N_28096,N_27844);
nor U29858 (N_29858,N_28366,N_27460);
or U29859 (N_29859,N_27518,N_27595);
or U29860 (N_29860,N_28104,N_28193);
or U29861 (N_29861,N_28211,N_27271);
nand U29862 (N_29862,N_28020,N_27686);
or U29863 (N_29863,N_27089,N_27900);
nand U29864 (N_29864,N_27737,N_27189);
and U29865 (N_29865,N_28416,N_27234);
xor U29866 (N_29866,N_27457,N_28250);
xor U29867 (N_29867,N_28275,N_27848);
nor U29868 (N_29868,N_27710,N_27418);
and U29869 (N_29869,N_27163,N_27893);
nand U29870 (N_29870,N_28002,N_28049);
or U29871 (N_29871,N_27315,N_27949);
xor U29872 (N_29872,N_28375,N_28002);
and U29873 (N_29873,N_27914,N_28307);
or U29874 (N_29874,N_27848,N_27833);
or U29875 (N_29875,N_27786,N_27017);
xor U29876 (N_29876,N_27264,N_27758);
or U29877 (N_29877,N_27337,N_28216);
and U29878 (N_29878,N_27610,N_28009);
nor U29879 (N_29879,N_27108,N_28499);
and U29880 (N_29880,N_28153,N_27169);
xor U29881 (N_29881,N_27585,N_27095);
nand U29882 (N_29882,N_27719,N_28272);
and U29883 (N_29883,N_27566,N_27599);
xor U29884 (N_29884,N_27910,N_27982);
nand U29885 (N_29885,N_27960,N_27052);
xor U29886 (N_29886,N_27510,N_28493);
and U29887 (N_29887,N_27453,N_27633);
xor U29888 (N_29888,N_27033,N_28013);
nor U29889 (N_29889,N_27449,N_27446);
and U29890 (N_29890,N_28360,N_28349);
xor U29891 (N_29891,N_27806,N_28216);
and U29892 (N_29892,N_27760,N_27864);
and U29893 (N_29893,N_27844,N_27459);
nor U29894 (N_29894,N_27459,N_28160);
and U29895 (N_29895,N_27723,N_27969);
or U29896 (N_29896,N_27929,N_28268);
nor U29897 (N_29897,N_27150,N_27225);
or U29898 (N_29898,N_27031,N_28140);
xnor U29899 (N_29899,N_27219,N_27433);
and U29900 (N_29900,N_27926,N_27755);
nor U29901 (N_29901,N_27983,N_27905);
nand U29902 (N_29902,N_28235,N_27168);
xnor U29903 (N_29903,N_27272,N_27380);
and U29904 (N_29904,N_27989,N_27218);
xor U29905 (N_29905,N_27195,N_28439);
and U29906 (N_29906,N_27956,N_28247);
or U29907 (N_29907,N_28293,N_27115);
nor U29908 (N_29908,N_27047,N_28348);
or U29909 (N_29909,N_28195,N_28078);
and U29910 (N_29910,N_28164,N_27911);
nor U29911 (N_29911,N_28224,N_28406);
nor U29912 (N_29912,N_28474,N_27913);
nor U29913 (N_29913,N_27488,N_27408);
nor U29914 (N_29914,N_27053,N_28331);
or U29915 (N_29915,N_27312,N_28335);
and U29916 (N_29916,N_27440,N_28175);
xor U29917 (N_29917,N_27823,N_27808);
or U29918 (N_29918,N_28460,N_27087);
and U29919 (N_29919,N_28374,N_27782);
nand U29920 (N_29920,N_27248,N_28497);
nand U29921 (N_29921,N_28410,N_27071);
nor U29922 (N_29922,N_27647,N_27121);
nor U29923 (N_29923,N_27310,N_28261);
and U29924 (N_29924,N_28224,N_27740);
nor U29925 (N_29925,N_27564,N_28044);
xor U29926 (N_29926,N_28174,N_27995);
or U29927 (N_29927,N_28386,N_27599);
nor U29928 (N_29928,N_27008,N_28491);
nand U29929 (N_29929,N_27757,N_27855);
nand U29930 (N_29930,N_27607,N_27832);
nor U29931 (N_29931,N_28037,N_28023);
nand U29932 (N_29932,N_27477,N_28117);
xor U29933 (N_29933,N_28346,N_27160);
xnor U29934 (N_29934,N_27863,N_27071);
nand U29935 (N_29935,N_27050,N_27437);
nand U29936 (N_29936,N_27904,N_28389);
and U29937 (N_29937,N_27302,N_27784);
and U29938 (N_29938,N_27491,N_28096);
nand U29939 (N_29939,N_27510,N_27620);
nor U29940 (N_29940,N_28386,N_28272);
and U29941 (N_29941,N_27396,N_28347);
nor U29942 (N_29942,N_28025,N_27299);
nor U29943 (N_29943,N_27096,N_27065);
xor U29944 (N_29944,N_27046,N_28406);
xnor U29945 (N_29945,N_28316,N_28274);
nor U29946 (N_29946,N_27848,N_27503);
nor U29947 (N_29947,N_28297,N_27018);
or U29948 (N_29948,N_27931,N_27671);
or U29949 (N_29949,N_27060,N_28357);
nand U29950 (N_29950,N_28213,N_27047);
xor U29951 (N_29951,N_27771,N_27742);
and U29952 (N_29952,N_27713,N_27372);
or U29953 (N_29953,N_27897,N_27501);
nor U29954 (N_29954,N_27579,N_27635);
or U29955 (N_29955,N_28059,N_27795);
nor U29956 (N_29956,N_27793,N_27248);
or U29957 (N_29957,N_28210,N_27889);
nor U29958 (N_29958,N_27956,N_27077);
nor U29959 (N_29959,N_28268,N_27883);
nand U29960 (N_29960,N_28271,N_27702);
xnor U29961 (N_29961,N_27502,N_27350);
nor U29962 (N_29962,N_27604,N_28097);
nor U29963 (N_29963,N_27395,N_27544);
and U29964 (N_29964,N_27685,N_28418);
nand U29965 (N_29965,N_27069,N_27392);
xor U29966 (N_29966,N_27229,N_28273);
xor U29967 (N_29967,N_27998,N_27935);
and U29968 (N_29968,N_28245,N_27969);
or U29969 (N_29969,N_27057,N_27616);
or U29970 (N_29970,N_27436,N_27132);
nand U29971 (N_29971,N_28348,N_27081);
nor U29972 (N_29972,N_28462,N_27897);
nor U29973 (N_29973,N_27290,N_27915);
xor U29974 (N_29974,N_27063,N_27981);
xnor U29975 (N_29975,N_27109,N_27317);
xor U29976 (N_29976,N_27146,N_27260);
nor U29977 (N_29977,N_27269,N_27403);
xor U29978 (N_29978,N_27396,N_28243);
or U29979 (N_29979,N_28338,N_28366);
and U29980 (N_29980,N_27515,N_27796);
xnor U29981 (N_29981,N_27719,N_27181);
nand U29982 (N_29982,N_27128,N_27736);
nand U29983 (N_29983,N_28301,N_28412);
nand U29984 (N_29984,N_28072,N_28020);
or U29985 (N_29985,N_28057,N_27513);
nor U29986 (N_29986,N_27101,N_27285);
or U29987 (N_29987,N_27265,N_27713);
nor U29988 (N_29988,N_27536,N_27387);
or U29989 (N_29989,N_27604,N_27361);
nand U29990 (N_29990,N_27035,N_27972);
nor U29991 (N_29991,N_27570,N_28387);
xnor U29992 (N_29992,N_27771,N_27828);
nor U29993 (N_29993,N_28284,N_27802);
and U29994 (N_29994,N_27433,N_28145);
or U29995 (N_29995,N_27791,N_27572);
nand U29996 (N_29996,N_28170,N_27455);
xnor U29997 (N_29997,N_27750,N_27265);
or U29998 (N_29998,N_27186,N_28131);
or U29999 (N_29999,N_27748,N_28369);
or UO_0 (O_0,N_29359,N_28669);
xnor UO_1 (O_1,N_28765,N_29906);
and UO_2 (O_2,N_29731,N_29618);
or UO_3 (O_3,N_28720,N_29717);
nand UO_4 (O_4,N_29071,N_28627);
xnor UO_5 (O_5,N_29568,N_29084);
and UO_6 (O_6,N_29609,N_29134);
nand UO_7 (O_7,N_29829,N_29849);
and UO_8 (O_8,N_28610,N_29825);
xnor UO_9 (O_9,N_29098,N_29170);
and UO_10 (O_10,N_28626,N_29328);
or UO_11 (O_11,N_28939,N_28793);
and UO_12 (O_12,N_29574,N_29467);
nand UO_13 (O_13,N_29081,N_28919);
nand UO_14 (O_14,N_28881,N_29539);
nand UO_15 (O_15,N_29299,N_28579);
nand UO_16 (O_16,N_29482,N_29128);
and UO_17 (O_17,N_29981,N_29211);
nand UO_18 (O_18,N_29343,N_29483);
and UO_19 (O_19,N_29641,N_29632);
xor UO_20 (O_20,N_28813,N_28513);
or UO_21 (O_21,N_28582,N_29325);
and UO_22 (O_22,N_28668,N_29649);
xor UO_23 (O_23,N_29136,N_28657);
nor UO_24 (O_24,N_28860,N_28866);
and UO_25 (O_25,N_28841,N_29000);
xor UO_26 (O_26,N_28565,N_29326);
and UO_27 (O_27,N_28664,N_28570);
nand UO_28 (O_28,N_29377,N_29747);
and UO_29 (O_29,N_29012,N_28755);
nor UO_30 (O_30,N_28876,N_29104);
nand UO_31 (O_31,N_29986,N_29209);
nor UO_32 (O_32,N_29276,N_28854);
or UO_33 (O_33,N_29407,N_28549);
nand UO_34 (O_34,N_29840,N_29861);
and UO_35 (O_35,N_28955,N_29666);
nand UO_36 (O_36,N_29603,N_29199);
xor UO_37 (O_37,N_29390,N_29912);
nor UO_38 (O_38,N_28891,N_28636);
and UO_39 (O_39,N_29621,N_28943);
nor UO_40 (O_40,N_28823,N_28604);
nand UO_41 (O_41,N_29578,N_29540);
xnor UO_42 (O_42,N_28547,N_29463);
nor UO_43 (O_43,N_29980,N_28617);
xnor UO_44 (O_44,N_29113,N_29311);
or UO_45 (O_45,N_29371,N_29651);
xor UO_46 (O_46,N_29910,N_28992);
xnor UO_47 (O_47,N_28723,N_29238);
nand UO_48 (O_48,N_29530,N_29320);
nor UO_49 (O_49,N_29809,N_29634);
nand UO_50 (O_50,N_29744,N_29970);
or UO_51 (O_51,N_29039,N_29347);
and UO_52 (O_52,N_28978,N_28808);
or UO_53 (O_53,N_28994,N_28873);
xor UO_54 (O_54,N_29440,N_29333);
nor UO_55 (O_55,N_29399,N_28735);
xor UO_56 (O_56,N_29414,N_29885);
nand UO_57 (O_57,N_28971,N_28804);
and UO_58 (O_58,N_29230,N_29415);
xnor UO_59 (O_59,N_29548,N_29888);
nand UO_60 (O_60,N_28621,N_29152);
nand UO_61 (O_61,N_29727,N_29705);
nand UO_62 (O_62,N_29119,N_29898);
and UO_63 (O_63,N_29792,N_29724);
xor UO_64 (O_64,N_29524,N_28874);
nand UO_65 (O_65,N_29750,N_29254);
nand UO_66 (O_66,N_29669,N_29363);
xor UO_67 (O_67,N_29880,N_28659);
nor UO_68 (O_68,N_28806,N_28965);
nor UO_69 (O_69,N_28786,N_29674);
and UO_70 (O_70,N_28768,N_29205);
and UO_71 (O_71,N_29497,N_28908);
and UO_72 (O_72,N_28524,N_29505);
nor UO_73 (O_73,N_29197,N_29477);
xnor UO_74 (O_74,N_28799,N_29506);
or UO_75 (O_75,N_29028,N_29346);
and UO_76 (O_76,N_29257,N_28890);
nand UO_77 (O_77,N_28719,N_29266);
xor UO_78 (O_78,N_29799,N_29614);
or UO_79 (O_79,N_28661,N_28567);
and UO_80 (O_80,N_28984,N_28538);
xor UO_81 (O_81,N_28801,N_29436);
nand UO_82 (O_82,N_29408,N_28756);
nor UO_83 (O_83,N_29633,N_28686);
nor UO_84 (O_84,N_29516,N_28504);
or UO_85 (O_85,N_28949,N_29661);
nand UO_86 (O_86,N_28798,N_29720);
nand UO_87 (O_87,N_29135,N_29663);
or UO_88 (O_88,N_29817,N_29203);
xnor UO_89 (O_89,N_29573,N_28677);
nand UO_90 (O_90,N_29766,N_28746);
xor UO_91 (O_91,N_29904,N_28647);
or UO_92 (O_92,N_28597,N_29221);
or UO_93 (O_93,N_29665,N_29718);
xor UO_94 (O_94,N_28802,N_28863);
and UO_95 (O_95,N_29358,N_29962);
nand UO_96 (O_96,N_29657,N_28910);
nand UO_97 (O_97,N_29531,N_29887);
xnor UO_98 (O_98,N_28809,N_29367);
xor UO_99 (O_99,N_29590,N_28564);
nor UO_100 (O_100,N_29522,N_29575);
nor UO_101 (O_101,N_28927,N_29564);
and UO_102 (O_102,N_28999,N_28578);
or UO_103 (O_103,N_28731,N_29942);
or UO_104 (O_104,N_28847,N_29867);
xnor UO_105 (O_105,N_29046,N_29008);
xnor UO_106 (O_106,N_28775,N_28505);
or UO_107 (O_107,N_28827,N_29298);
and UO_108 (O_108,N_29340,N_29490);
nand UO_109 (O_109,N_29916,N_29097);
or UO_110 (O_110,N_28958,N_29245);
nand UO_111 (O_111,N_29033,N_28913);
nand UO_112 (O_112,N_29406,N_29389);
xor UO_113 (O_113,N_28737,N_28898);
or UO_114 (O_114,N_29294,N_29638);
or UO_115 (O_115,N_29940,N_28869);
xor UO_116 (O_116,N_29272,N_28838);
nand UO_117 (O_117,N_29421,N_29869);
and UO_118 (O_118,N_28857,N_28633);
and UO_119 (O_119,N_29220,N_29026);
or UO_120 (O_120,N_28993,N_29001);
or UO_121 (O_121,N_29581,N_29789);
or UO_122 (O_122,N_29950,N_29527);
or UO_123 (O_123,N_29570,N_28771);
and UO_124 (O_124,N_29120,N_29056);
and UO_125 (O_125,N_29379,N_28722);
nand UO_126 (O_126,N_28935,N_28629);
xor UO_127 (O_127,N_29741,N_29159);
nor UO_128 (O_128,N_29156,N_29608);
xnor UO_129 (O_129,N_28725,N_28918);
and UO_130 (O_130,N_28708,N_29819);
or UO_131 (O_131,N_29279,N_28527);
xor UO_132 (O_132,N_29895,N_28744);
nand UO_133 (O_133,N_28609,N_29019);
xnor UO_134 (O_134,N_29446,N_29429);
and UO_135 (O_135,N_29434,N_29612);
xor UO_136 (O_136,N_29443,N_28718);
or UO_137 (O_137,N_29274,N_29251);
nand UO_138 (O_138,N_28563,N_29991);
and UO_139 (O_139,N_29932,N_29773);
and UO_140 (O_140,N_29141,N_28986);
and UO_141 (O_141,N_29123,N_29957);
nand UO_142 (O_142,N_29722,N_28620);
and UO_143 (O_143,N_29528,N_29210);
nand UO_144 (O_144,N_28783,N_28551);
or UO_145 (O_145,N_28501,N_29258);
xnor UO_146 (O_146,N_28666,N_28608);
nand UO_147 (O_147,N_29402,N_29133);
xnor UO_148 (O_148,N_29743,N_29450);
nand UO_149 (O_149,N_28745,N_29316);
nor UO_150 (O_150,N_29512,N_29647);
nand UO_151 (O_151,N_29262,N_28596);
nand UO_152 (O_152,N_29395,N_29973);
or UO_153 (O_153,N_29937,N_29250);
nand UO_154 (O_154,N_29827,N_29821);
nor UO_155 (O_155,N_29546,N_28644);
nor UO_156 (O_156,N_28968,N_29112);
xnor UO_157 (O_157,N_29074,N_28820);
nor UO_158 (O_158,N_28576,N_29925);
and UO_159 (O_159,N_28946,N_28662);
and UO_160 (O_160,N_29312,N_28982);
nand UO_161 (O_161,N_28688,N_28577);
and UO_162 (O_162,N_29302,N_29783);
nand UO_163 (O_163,N_29457,N_29162);
or UO_164 (O_164,N_29810,N_28909);
nor UO_165 (O_165,N_29969,N_29561);
nor UO_166 (O_166,N_29751,N_29862);
and UO_167 (O_167,N_29968,N_29529);
and UO_168 (O_168,N_29896,N_28778);
or UO_169 (O_169,N_28936,N_29460);
and UO_170 (O_170,N_29818,N_29486);
nor UO_171 (O_171,N_29972,N_28835);
and UO_172 (O_172,N_28566,N_29853);
xnor UO_173 (O_173,N_29627,N_29671);
nor UO_174 (O_174,N_29286,N_28784);
nor UO_175 (O_175,N_29479,N_28534);
and UO_176 (O_176,N_29598,N_29858);
nor UO_177 (O_177,N_29356,N_28648);
and UO_178 (O_178,N_29719,N_28973);
and UO_179 (O_179,N_29079,N_28619);
nor UO_180 (O_180,N_29737,N_28836);
nor UO_181 (O_181,N_29922,N_28815);
and UO_182 (O_182,N_29150,N_29556);
nor UO_183 (O_183,N_28681,N_29726);
or UO_184 (O_184,N_29617,N_28700);
xor UO_185 (O_185,N_29297,N_28580);
xor UO_186 (O_186,N_28655,N_29329);
and UO_187 (O_187,N_29198,N_28638);
nand UO_188 (O_188,N_29144,N_29894);
or UO_189 (O_189,N_28675,N_29049);
nor UO_190 (O_190,N_29958,N_29161);
and UO_191 (O_191,N_28751,N_28717);
and UO_192 (O_192,N_29374,N_29448);
nand UO_193 (O_193,N_29301,N_29044);
nand UO_194 (O_194,N_29337,N_28901);
nor UO_195 (O_195,N_29029,N_28931);
and UO_196 (O_196,N_28732,N_29680);
nand UO_197 (O_197,N_29303,N_28606);
nand UO_198 (O_198,N_28998,N_28739);
xnor UO_199 (O_199,N_29283,N_29190);
nor UO_200 (O_200,N_29845,N_29721);
or UO_201 (O_201,N_28598,N_28684);
or UO_202 (O_202,N_28667,N_29015);
nor UO_203 (O_203,N_29260,N_29129);
nor UO_204 (O_204,N_29660,N_29189);
and UO_205 (O_205,N_29938,N_29105);
and UO_206 (O_206,N_29289,N_28753);
nand UO_207 (O_207,N_29403,N_29848);
nor UO_208 (O_208,N_29416,N_29735);
nor UO_209 (O_209,N_28500,N_29879);
or UO_210 (O_210,N_28941,N_28789);
xor UO_211 (O_211,N_29716,N_28800);
nand UO_212 (O_212,N_29860,N_29109);
and UO_213 (O_213,N_28589,N_29749);
nor UO_214 (O_214,N_29708,N_29077);
xor UO_215 (O_215,N_29915,N_28894);
or UO_216 (O_216,N_29936,N_29419);
xnor UO_217 (O_217,N_29075,N_28516);
xnor UO_218 (O_218,N_28856,N_29801);
and UO_219 (O_219,N_28981,N_28861);
nand UO_220 (O_220,N_28837,N_29424);
nor UO_221 (O_221,N_29375,N_28569);
or UO_222 (O_222,N_29692,N_29380);
nand UO_223 (O_223,N_28792,N_29763);
or UO_224 (O_224,N_29194,N_28780);
or UO_225 (O_225,N_29174,N_29820);
and UO_226 (O_226,N_29239,N_28523);
or UO_227 (O_227,N_29410,N_29089);
nor UO_228 (O_228,N_28715,N_28671);
nand UO_229 (O_229,N_29465,N_29370);
nand UO_230 (O_230,N_29688,N_29110);
xnor UO_231 (O_231,N_28646,N_28554);
nor UO_232 (O_232,N_29067,N_29070);
and UO_233 (O_233,N_29130,N_28911);
nor UO_234 (O_234,N_28899,N_28591);
nor UO_235 (O_235,N_29057,N_28896);
or UO_236 (O_236,N_29143,N_29300);
or UO_237 (O_237,N_28709,N_29499);
nor UO_238 (O_238,N_29226,N_29035);
and UO_239 (O_239,N_29715,N_28740);
xor UO_240 (O_240,N_29249,N_29353);
and UO_241 (O_241,N_29831,N_29814);
nor UO_242 (O_242,N_29532,N_29670);
nand UO_243 (O_243,N_29805,N_29664);
and UO_244 (O_244,N_29405,N_28512);
xor UO_245 (O_245,N_29160,N_29668);
or UO_246 (O_246,N_29914,N_29934);
nand UO_247 (O_247,N_28691,N_28782);
or UO_248 (O_248,N_29317,N_28650);
or UO_249 (O_249,N_29689,N_29882);
or UO_250 (O_250,N_28697,N_28510);
or UO_251 (O_251,N_28825,N_28665);
and UO_252 (O_252,N_29591,N_29271);
nor UO_253 (O_253,N_28588,N_28829);
xor UO_254 (O_254,N_29281,N_29489);
nor UO_255 (O_255,N_29865,N_28502);
nor UO_256 (O_256,N_29510,N_29228);
and UO_257 (O_257,N_29780,N_29439);
xnor UO_258 (O_258,N_28987,N_29182);
nand UO_259 (O_259,N_29031,N_29427);
nor UO_260 (O_260,N_29016,N_28848);
xor UO_261 (O_261,N_28678,N_29212);
nor UO_262 (O_262,N_29107,N_29856);
nand UO_263 (O_263,N_29710,N_28773);
and UO_264 (O_264,N_29058,N_28980);
nor UO_265 (O_265,N_29901,N_28517);
nor UO_266 (O_266,N_29485,N_29494);
nor UO_267 (O_267,N_29462,N_29273);
or UO_268 (O_268,N_29622,N_28628);
nand UO_269 (O_269,N_29456,N_28616);
or UO_270 (O_270,N_29218,N_28702);
xnor UO_271 (O_271,N_28673,N_28832);
xnor UO_272 (O_272,N_29559,N_28821);
and UO_273 (O_273,N_29188,N_29127);
and UO_274 (O_274,N_29225,N_29224);
or UO_275 (O_275,N_29268,N_29905);
and UO_276 (O_276,N_28590,N_29565);
nand UO_277 (O_277,N_29960,N_29315);
nand UO_278 (O_278,N_28506,N_29919);
nand UO_279 (O_279,N_29233,N_29157);
nand UO_280 (O_280,N_29392,N_29884);
xnor UO_281 (O_281,N_29642,N_29501);
xnor UO_282 (O_282,N_29760,N_28865);
nor UO_283 (O_283,N_28546,N_29562);
xnor UO_284 (O_284,N_28924,N_29053);
and UO_285 (O_285,N_29695,N_29148);
nor UO_286 (O_286,N_28733,N_29847);
and UO_287 (O_287,N_29623,N_28858);
xnor UO_288 (O_288,N_29171,N_28575);
nand UO_289 (O_289,N_28870,N_29536);
or UO_290 (O_290,N_29579,N_29338);
nor UO_291 (O_291,N_29180,N_28743);
nand UO_292 (O_292,N_29544,N_29703);
xnor UO_293 (O_293,N_29362,N_28728);
nor UO_294 (O_294,N_29437,N_29396);
xnor UO_295 (O_295,N_29132,N_28679);
nand UO_296 (O_296,N_28875,N_29247);
nor UO_297 (O_297,N_29111,N_29842);
nand UO_298 (O_298,N_28571,N_29740);
nand UO_299 (O_299,N_29386,N_29961);
or UO_300 (O_300,N_29354,N_29625);
xor UO_301 (O_301,N_29954,N_29577);
and UO_302 (O_302,N_28851,N_28692);
and UO_303 (O_303,N_28831,N_29471);
xnor UO_304 (O_304,N_29106,N_29543);
nand UO_305 (O_305,N_28964,N_29580);
or UO_306 (O_306,N_29701,N_29235);
nor UO_307 (O_307,N_29126,N_29640);
nor UO_308 (O_308,N_29401,N_29813);
xor UO_309 (O_309,N_29227,N_28921);
nand UO_310 (O_310,N_28929,N_29757);
xor UO_311 (O_311,N_28830,N_28796);
and UO_312 (O_312,N_29065,N_29868);
or UO_313 (O_313,N_29746,N_29907);
nor UO_314 (O_314,N_29576,N_29352);
or UO_315 (O_315,N_29487,N_29630);
or UO_316 (O_316,N_28788,N_28845);
xor UO_317 (O_317,N_29229,N_28952);
or UO_318 (O_318,N_28907,N_28607);
xor UO_319 (O_319,N_29890,N_28862);
nand UO_320 (O_320,N_29285,N_28940);
nand UO_321 (O_321,N_29005,N_29723);
nand UO_322 (O_322,N_28849,N_29534);
nand UO_323 (O_323,N_29096,N_29851);
nor UO_324 (O_324,N_29480,N_29038);
nor UO_325 (O_325,N_29515,N_29116);
xnor UO_326 (O_326,N_29990,N_29381);
nor UO_327 (O_327,N_29798,N_29673);
xor UO_328 (O_328,N_29214,N_28561);
or UO_329 (O_329,N_29237,N_29178);
or UO_330 (O_330,N_29877,N_28568);
nor UO_331 (O_331,N_28752,N_29378);
xor UO_332 (O_332,N_29176,N_28531);
and UO_333 (O_333,N_29142,N_28762);
nor UO_334 (O_334,N_29784,N_29411);
nor UO_335 (O_335,N_28543,N_29087);
nor UO_336 (O_336,N_28853,N_29054);
nand UO_337 (O_337,N_29796,N_28613);
or UO_338 (O_338,N_29108,N_28942);
and UO_339 (O_339,N_28558,N_29394);
nor UO_340 (O_340,N_28904,N_29832);
nor UO_341 (O_341,N_29607,N_28642);
and UO_342 (O_342,N_29491,N_28879);
and UO_343 (O_343,N_29124,N_29458);
and UO_344 (O_344,N_29500,N_29167);
or UO_345 (O_345,N_28658,N_29728);
xor UO_346 (O_346,N_28764,N_29172);
or UO_347 (O_347,N_29383,N_29777);
nand UO_348 (O_348,N_29153,N_29704);
nor UO_349 (O_349,N_29020,N_29449);
xnor UO_350 (O_350,N_29086,N_29850);
nor UO_351 (O_351,N_29733,N_28585);
nor UO_352 (O_352,N_28791,N_29983);
and UO_353 (O_353,N_29444,N_28970);
xnor UO_354 (O_354,N_28539,N_29658);
and UO_355 (O_355,N_29521,N_29770);
nor UO_356 (O_356,N_29422,N_28519);
xnor UO_357 (O_357,N_29305,N_29854);
or UO_358 (O_358,N_28701,N_29027);
and UO_359 (O_359,N_28794,N_29620);
and UO_360 (O_360,N_29208,N_28748);
nor UO_361 (O_361,N_28727,N_29324);
or UO_362 (O_362,N_29795,N_29100);
nor UO_363 (O_363,N_29547,N_29985);
or UO_364 (O_364,N_29903,N_28948);
or UO_365 (O_365,N_29287,N_28533);
nand UO_366 (O_366,N_29277,N_29837);
nor UO_367 (O_367,N_28574,N_29335);
nand UO_368 (O_368,N_29738,N_29369);
nand UO_369 (O_369,N_29115,N_28738);
nand UO_370 (O_370,N_28514,N_28541);
nor UO_371 (O_371,N_29552,N_29288);
nor UO_372 (O_372,N_29184,N_29892);
or UO_373 (O_373,N_28749,N_28611);
nand UO_374 (O_374,N_28839,N_29259);
or UO_375 (O_375,N_29899,N_28974);
or UO_376 (O_376,N_29014,N_28916);
xor UO_377 (O_377,N_29871,N_28938);
and UO_378 (O_378,N_29255,N_29822);
nor UO_379 (O_379,N_29902,N_29606);
nor UO_380 (O_380,N_29857,N_28880);
xnor UO_381 (O_381,N_29496,N_29765);
xor UO_382 (O_382,N_29654,N_29526);
or UO_383 (O_383,N_29931,N_28886);
nor UO_384 (O_384,N_29024,N_29706);
and UO_385 (O_385,N_28842,N_28819);
or UO_386 (O_386,N_29451,N_29140);
nand UO_387 (O_387,N_29196,N_28960);
and UO_388 (O_388,N_29537,N_28776);
or UO_389 (O_389,N_29385,N_29252);
nand UO_390 (O_390,N_28844,N_28925);
nand UO_391 (O_391,N_29611,N_29060);
nor UO_392 (O_392,N_29202,N_28895);
nor UO_393 (O_393,N_29586,N_29927);
nand UO_394 (O_394,N_29200,N_29447);
nand UO_395 (O_395,N_29791,N_29361);
xnor UO_396 (O_396,N_29461,N_29769);
nand UO_397 (O_397,N_29217,N_28711);
nor UO_398 (O_398,N_29920,N_29545);
nand UO_399 (O_399,N_29676,N_29322);
and UO_400 (O_400,N_28529,N_29063);
and UO_401 (O_401,N_28817,N_29730);
nor UO_402 (O_402,N_29433,N_29158);
or UO_403 (O_403,N_29987,N_29939);
nor UO_404 (O_404,N_28962,N_29846);
xnor UO_405 (O_405,N_29023,N_29691);
nand UO_406 (O_406,N_29484,N_28713);
and UO_407 (O_407,N_29678,N_28742);
xor UO_408 (O_408,N_28972,N_29165);
nand UO_409 (O_409,N_29073,N_28966);
xnor UO_410 (O_410,N_28649,N_29473);
or UO_411 (O_411,N_29808,N_29652);
and UO_412 (O_412,N_29953,N_29732);
nand UO_413 (O_413,N_29166,N_29613);
and UO_414 (O_414,N_28689,N_28548);
and UO_415 (O_415,N_29518,N_29948);
nand UO_416 (O_416,N_29707,N_28660);
nor UO_417 (O_417,N_28696,N_29048);
nor UO_418 (O_418,N_29043,N_28712);
or UO_419 (O_419,N_28805,N_28833);
nand UO_420 (O_420,N_28900,N_29185);
and UO_421 (O_421,N_28757,N_29772);
xnor UO_422 (O_422,N_28584,N_29563);
nor UO_423 (O_423,N_28915,N_29571);
nor UO_424 (O_424,N_29240,N_29125);
xnor UO_425 (O_425,N_29307,N_29149);
and UO_426 (O_426,N_29794,N_29525);
nand UO_427 (O_427,N_28790,N_29050);
or UO_428 (O_428,N_29318,N_28963);
nor UO_429 (O_429,N_28877,N_29839);
and UO_430 (O_430,N_29807,N_29684);
and UO_431 (O_431,N_29169,N_29420);
nand UO_432 (O_432,N_28716,N_29917);
nand UO_433 (O_433,N_29913,N_29041);
nand UO_434 (O_434,N_29551,N_29533);
and UO_435 (O_435,N_29030,N_28605);
or UO_436 (O_436,N_29503,N_29816);
and UO_437 (O_437,N_29959,N_29206);
or UO_438 (O_438,N_28781,N_29398);
or UO_439 (O_439,N_28828,N_29145);
nand UO_440 (O_440,N_28643,N_29683);
and UO_441 (O_441,N_28640,N_29121);
nor UO_442 (O_442,N_29011,N_29232);
nand UO_443 (O_443,N_29042,N_29223);
or UO_444 (O_444,N_29835,N_29520);
and UO_445 (O_445,N_28507,N_29267);
nand UO_446 (O_446,N_29535,N_29009);
or UO_447 (O_447,N_29872,N_28864);
nand UO_448 (O_448,N_29364,N_28540);
and UO_449 (O_449,N_29013,N_28797);
and UO_450 (O_450,N_29191,N_29253);
nor UO_451 (O_451,N_29413,N_29099);
and UO_452 (O_452,N_29874,N_29393);
nor UO_453 (O_453,N_29826,N_28846);
nand UO_454 (O_454,N_29756,N_29788);
xnor UO_455 (O_455,N_29748,N_29659);
xor UO_456 (O_456,N_29933,N_28885);
or UO_457 (O_457,N_28695,N_28511);
and UO_458 (O_458,N_28525,N_29762);
nand UO_459 (O_459,N_29092,N_29786);
or UO_460 (O_460,N_28586,N_29928);
nor UO_461 (O_461,N_28897,N_29323);
xnor UO_462 (O_462,N_29594,N_28750);
nand UO_463 (O_463,N_28622,N_29992);
and UO_464 (O_464,N_29605,N_29365);
xor UO_465 (O_465,N_29055,N_29697);
nand UO_466 (O_466,N_29975,N_29412);
nor UO_467 (O_467,N_29560,N_29059);
nor UO_468 (O_468,N_28997,N_29930);
nor UO_469 (O_469,N_29061,N_28816);
nor UO_470 (O_470,N_29442,N_29094);
and UO_471 (O_471,N_29306,N_29971);
and UO_472 (O_472,N_29682,N_28889);
xor UO_473 (O_473,N_29095,N_29790);
nor UO_474 (O_474,N_29812,N_29082);
and UO_475 (O_475,N_29690,N_29131);
nor UO_476 (O_476,N_29597,N_29332);
nand UO_477 (O_477,N_29508,N_29918);
and UO_478 (O_478,N_29834,N_29921);
nand UO_479 (O_479,N_29264,N_28683);
or UO_480 (O_480,N_28508,N_28934);
and UO_481 (O_481,N_29998,N_28956);
nor UO_482 (O_482,N_29088,N_29844);
or UO_483 (O_483,N_29215,N_28654);
and UO_484 (O_484,N_28557,N_28726);
and UO_485 (O_485,N_28693,N_29181);
and UO_486 (O_486,N_28906,N_28902);
xnor UO_487 (O_487,N_29929,N_29873);
xnor UO_488 (O_488,N_29947,N_29811);
nand UO_489 (O_489,N_29681,N_29550);
nand UO_490 (O_490,N_28653,N_29453);
nor UO_491 (O_491,N_29445,N_29068);
nand UO_492 (O_492,N_28522,N_29891);
nand UO_493 (O_493,N_29963,N_29761);
nor UO_494 (O_494,N_29327,N_28961);
and UO_495 (O_495,N_28581,N_28957);
xor UO_496 (O_496,N_29863,N_29417);
and UO_497 (O_497,N_29204,N_29781);
xor UO_498 (O_498,N_28763,N_29804);
nand UO_499 (O_499,N_28639,N_29610);
and UO_500 (O_500,N_29686,N_29295);
nor UO_501 (O_501,N_29213,N_28623);
and UO_502 (O_502,N_29889,N_28656);
and UO_503 (O_503,N_29069,N_29852);
xor UO_504 (O_504,N_29549,N_28930);
nor UO_505 (O_505,N_28587,N_28884);
or UO_506 (O_506,N_29334,N_29626);
and UO_507 (O_507,N_29256,N_29739);
nand UO_508 (O_508,N_29587,N_29179);
nor UO_509 (O_509,N_28509,N_29977);
and UO_510 (O_510,N_28953,N_28989);
nor UO_511 (O_511,N_28637,N_28600);
nand UO_512 (O_512,N_28562,N_29093);
or UO_513 (O_513,N_28706,N_29064);
nor UO_514 (O_514,N_29557,N_29999);
and UO_515 (O_515,N_29103,N_29387);
nand UO_516 (O_516,N_29976,N_28903);
xor UO_517 (O_517,N_28625,N_29996);
and UO_518 (O_518,N_29567,N_28988);
nor UO_519 (O_519,N_28944,N_28795);
nor UO_520 (O_520,N_29935,N_29045);
and UO_521 (O_521,N_29881,N_29509);
xnor UO_522 (O_522,N_28859,N_29441);
xnor UO_523 (O_523,N_29644,N_28729);
and UO_524 (O_524,N_29685,N_28612);
xor UO_525 (O_525,N_28652,N_29313);
and UO_526 (O_526,N_29513,N_28710);
and UO_527 (O_527,N_29350,N_28528);
nand UO_528 (O_528,N_29517,N_29321);
nor UO_529 (O_529,N_29409,N_29672);
nor UO_530 (O_530,N_29003,N_29219);
or UO_531 (O_531,N_28933,N_29310);
xnor UO_532 (O_532,N_28670,N_29117);
xnor UO_533 (O_533,N_29569,N_29893);
xnor UO_534 (O_534,N_28503,N_29592);
nand UO_535 (O_535,N_29875,N_28772);
and UO_536 (O_536,N_28630,N_28887);
and UO_537 (O_537,N_29924,N_29498);
nor UO_538 (O_538,N_29636,N_29582);
and UO_539 (O_539,N_29698,N_29357);
or UO_540 (O_540,N_29454,N_28811);
nand UO_541 (O_541,N_29388,N_28676);
nor UO_542 (O_542,N_29168,N_29648);
or UO_543 (O_543,N_29051,N_29366);
nor UO_544 (O_544,N_28698,N_29758);
or UO_545 (O_545,N_29432,N_29965);
nor UO_546 (O_546,N_29231,N_29308);
nor UO_547 (O_547,N_29599,N_28730);
nand UO_548 (O_548,N_29502,N_29102);
nand UO_549 (O_549,N_29776,N_29759);
or UO_550 (O_550,N_29693,N_28779);
nand UO_551 (O_551,N_29554,N_29742);
xnor UO_552 (O_552,N_29909,N_29767);
nor UO_553 (O_553,N_29886,N_29883);
xor UO_554 (O_554,N_29583,N_29650);
xnor UO_555 (O_555,N_29542,N_29687);
xor UO_556 (O_556,N_29004,N_28685);
nand UO_557 (O_557,N_28594,N_29309);
nor UO_558 (O_558,N_29787,N_28834);
nor UO_559 (O_559,N_29455,N_28893);
nand UO_560 (O_560,N_28741,N_29908);
or UO_561 (O_561,N_29662,N_28544);
nand UO_562 (O_562,N_29806,N_29425);
and UO_563 (O_563,N_29269,N_29349);
nor UO_564 (O_564,N_28945,N_28593);
nor UO_565 (O_565,N_29372,N_29507);
or UO_566 (O_566,N_29368,N_28985);
nand UO_567 (O_567,N_29519,N_29949);
nor UO_568 (O_568,N_28818,N_29943);
xor UO_569 (O_569,N_28892,N_28615);
or UO_570 (O_570,N_29714,N_29192);
nand UO_571 (O_571,N_29459,N_29146);
nand UO_572 (O_572,N_29995,N_28682);
or UO_573 (O_573,N_29155,N_29474);
nand UO_574 (O_574,N_29978,N_29034);
xor UO_575 (O_575,N_28599,N_28777);
nor UO_576 (O_576,N_29589,N_28785);
xnor UO_577 (O_577,N_29523,N_29466);
and UO_578 (O_578,N_29859,N_29709);
and UO_579 (O_579,N_29175,N_29823);
or UO_580 (O_580,N_29736,N_29566);
and UO_581 (O_581,N_28905,N_29291);
nor UO_582 (O_582,N_29122,N_28996);
or UO_583 (O_583,N_28951,N_29768);
nand UO_584 (O_584,N_28991,N_29052);
xnor UO_585 (O_585,N_29154,N_29514);
or UO_586 (O_586,N_29838,N_29675);
or UO_587 (O_587,N_29645,N_29982);
xor UO_588 (O_588,N_28822,N_28552);
nand UO_589 (O_589,N_28559,N_29800);
nand UO_590 (O_590,N_29797,N_29355);
and UO_591 (O_591,N_29677,N_28976);
nor UO_592 (O_592,N_29833,N_29336);
nor UO_593 (O_593,N_29470,N_29018);
or UO_594 (O_594,N_29195,N_28787);
or UO_595 (O_595,N_29007,N_29945);
and UO_596 (O_596,N_28672,N_29083);
and UO_597 (O_597,N_29604,N_29236);
and UO_598 (O_598,N_28983,N_29911);
nor UO_599 (O_599,N_28645,N_28618);
or UO_600 (O_600,N_28774,N_29080);
and UO_601 (O_601,N_28555,N_28758);
xnor UO_602 (O_602,N_29078,N_29022);
xor UO_603 (O_603,N_28824,N_29643);
nand UO_604 (O_604,N_29729,N_28734);
or UO_605 (O_605,N_28550,N_28922);
nand UO_606 (O_606,N_29755,N_28535);
nand UO_607 (O_607,N_28767,N_29348);
nand UO_608 (O_608,N_29006,N_29653);
and UO_609 (O_609,N_28923,N_28631);
and UO_610 (O_610,N_28807,N_28680);
nor UO_611 (O_611,N_29010,N_28967);
or UO_612 (O_612,N_28553,N_29319);
nand UO_613 (O_613,N_29595,N_28812);
nor UO_614 (O_614,N_28635,N_29187);
xnor UO_615 (O_615,N_29216,N_29468);
xor UO_616 (O_616,N_29553,N_29090);
or UO_617 (O_617,N_29384,N_29753);
nand UO_618 (O_618,N_29700,N_29679);
or UO_619 (O_619,N_29984,N_29541);
nor UO_620 (O_620,N_29032,N_28920);
nand UO_621 (O_621,N_29628,N_28624);
xnor UO_622 (O_622,N_29488,N_29778);
or UO_623 (O_623,N_29619,N_28560);
and UO_624 (O_624,N_28754,N_29376);
and UO_625 (O_625,N_28878,N_29139);
xor UO_626 (O_626,N_29431,N_29118);
and UO_627 (O_627,N_29941,N_29878);
and UO_628 (O_628,N_29397,N_28975);
nand UO_629 (O_629,N_29855,N_29278);
nand UO_630 (O_630,N_29341,N_28724);
xor UO_631 (O_631,N_28850,N_29655);
nor UO_632 (O_632,N_29234,N_29275);
or UO_633 (O_633,N_28532,N_29478);
xnor UO_634 (O_634,N_29114,N_28603);
xnor UO_635 (O_635,N_29248,N_28690);
nor UO_636 (O_636,N_28721,N_29946);
or UO_637 (O_637,N_29988,N_28888);
and UO_638 (O_638,N_28614,N_28803);
and UO_639 (O_639,N_29373,N_29472);
and UO_640 (O_640,N_29147,N_29629);
xor UO_641 (O_641,N_29764,N_28556);
or UO_642 (O_642,N_28518,N_29966);
and UO_643 (O_643,N_29774,N_28760);
nand UO_644 (O_644,N_28969,N_28699);
xor UO_645 (O_645,N_29469,N_29331);
xor UO_646 (O_646,N_29712,N_29339);
xor UO_647 (O_647,N_29292,N_29047);
nand UO_648 (O_648,N_28766,N_29639);
nor UO_649 (O_649,N_29656,N_28573);
or UO_650 (O_650,N_29994,N_28840);
xnor UO_651 (O_651,N_29423,N_29585);
nor UO_652 (O_652,N_28515,N_28704);
xor UO_653 (O_653,N_28632,N_29828);
nand UO_654 (O_654,N_29711,N_29964);
nand UO_655 (O_655,N_29284,N_29270);
nor UO_656 (O_656,N_29085,N_28979);
and UO_657 (O_657,N_29694,N_28814);
or UO_658 (O_658,N_29280,N_28770);
xnor UO_659 (O_659,N_29967,N_28914);
nor UO_660 (O_660,N_28572,N_29944);
xnor UO_661 (O_661,N_29616,N_28736);
nand UO_662 (O_662,N_29430,N_29637);
and UO_663 (O_663,N_29997,N_29435);
xnor UO_664 (O_664,N_29492,N_29584);
or UO_665 (O_665,N_29602,N_29091);
and UO_666 (O_666,N_29824,N_29438);
xor UO_667 (O_667,N_29101,N_28694);
or UO_668 (O_668,N_28521,N_28959);
nor UO_669 (O_669,N_29186,N_28545);
or UO_670 (O_670,N_29601,N_29351);
or UO_671 (O_671,N_29037,N_29866);
or UO_672 (O_672,N_29785,N_29222);
and UO_673 (O_673,N_29344,N_29667);
xnor UO_674 (O_674,N_28536,N_29775);
and UO_675 (O_675,N_29734,N_29193);
xor UO_676 (O_676,N_28526,N_28595);
nor UO_677 (O_677,N_28674,N_28826);
nor UO_678 (O_678,N_29955,N_29538);
nor UO_679 (O_679,N_28928,N_29137);
xnor UO_680 (O_680,N_29382,N_29754);
nor UO_681 (O_681,N_28990,N_29293);
nor UO_682 (O_682,N_29870,N_29713);
or UO_683 (O_683,N_29802,N_29900);
nand UO_684 (O_684,N_29615,N_29815);
and UO_685 (O_685,N_29391,N_28882);
or UO_686 (O_686,N_29261,N_29864);
nor UO_687 (O_687,N_29504,N_29696);
or UO_688 (O_688,N_29330,N_29779);
xnor UO_689 (O_689,N_29495,N_29979);
nand UO_690 (O_690,N_28592,N_29725);
and UO_691 (O_691,N_29752,N_29241);
xnor UO_692 (O_692,N_29993,N_28602);
nand UO_693 (O_693,N_28759,N_29002);
xor UO_694 (O_694,N_29452,N_28601);
xor UO_695 (O_695,N_29314,N_29076);
nand UO_696 (O_696,N_28883,N_29989);
and UO_697 (O_697,N_28937,N_29631);
or UO_698 (O_698,N_29243,N_29244);
xor UO_699 (O_699,N_29040,N_28520);
and UO_700 (O_700,N_28634,N_29476);
nor UO_701 (O_701,N_29803,N_28769);
nand UO_702 (O_702,N_28542,N_28761);
or UO_703 (O_703,N_28852,N_29173);
xor UO_704 (O_704,N_29163,N_29265);
nor UO_705 (O_705,N_28932,N_29426);
or UO_706 (O_706,N_29242,N_28912);
and UO_707 (O_707,N_28530,N_29600);
and UO_708 (O_708,N_29342,N_29177);
nand UO_709 (O_709,N_28871,N_29588);
or UO_710 (O_710,N_28947,N_29956);
xor UO_711 (O_711,N_29183,N_29974);
xor UO_712 (O_712,N_28977,N_29036);
nand UO_713 (O_713,N_29841,N_29782);
nand UO_714 (O_714,N_28843,N_28714);
xnor UO_715 (O_715,N_29793,N_28855);
xnor UO_716 (O_716,N_29464,N_28705);
nor UO_717 (O_717,N_29635,N_29296);
nor UO_718 (O_718,N_29830,N_28872);
or UO_719 (O_719,N_29593,N_28867);
nor UO_720 (O_720,N_28950,N_29290);
and UO_721 (O_721,N_29481,N_29624);
or UO_722 (O_722,N_29360,N_29771);
nand UO_723 (O_723,N_29572,N_28707);
nand UO_724 (O_724,N_29201,N_28537);
or UO_725 (O_725,N_29066,N_29151);
xor UO_726 (O_726,N_28917,N_29428);
xor UO_727 (O_727,N_29951,N_29646);
nand UO_728 (O_728,N_28687,N_28810);
xnor UO_729 (O_729,N_29304,N_28954);
nor UO_730 (O_730,N_29699,N_29345);
nor UO_731 (O_731,N_29404,N_29164);
and UO_732 (O_732,N_29418,N_29400);
and UO_733 (O_733,N_29745,N_29555);
xor UO_734 (O_734,N_29836,N_29511);
nand UO_735 (O_735,N_29558,N_29021);
nand UO_736 (O_736,N_28641,N_29207);
or UO_737 (O_737,N_29025,N_28703);
and UO_738 (O_738,N_29138,N_29475);
nor UO_739 (O_739,N_29926,N_29493);
nand UO_740 (O_740,N_29263,N_28583);
nor UO_741 (O_741,N_29897,N_28747);
nor UO_742 (O_742,N_29876,N_29923);
nor UO_743 (O_743,N_28926,N_28995);
xnor UO_744 (O_744,N_28868,N_29282);
and UO_745 (O_745,N_29952,N_29017);
and UO_746 (O_746,N_28651,N_28663);
xnor UO_747 (O_747,N_29702,N_29072);
and UO_748 (O_748,N_29246,N_29062);
nand UO_749 (O_749,N_29843,N_29596);
xnor UO_750 (O_750,N_29447,N_29331);
nand UO_751 (O_751,N_29035,N_29222);
nor UO_752 (O_752,N_29480,N_28550);
nor UO_753 (O_753,N_28835,N_28959);
xnor UO_754 (O_754,N_28587,N_29980);
or UO_755 (O_755,N_28914,N_29727);
nor UO_756 (O_756,N_29748,N_29740);
nor UO_757 (O_757,N_28599,N_29700);
xnor UO_758 (O_758,N_29938,N_28733);
nand UO_759 (O_759,N_29165,N_29392);
xnor UO_760 (O_760,N_29009,N_28599);
nor UO_761 (O_761,N_29099,N_28747);
nor UO_762 (O_762,N_29322,N_28601);
and UO_763 (O_763,N_29488,N_29893);
and UO_764 (O_764,N_28837,N_28755);
nand UO_765 (O_765,N_29119,N_29105);
nor UO_766 (O_766,N_28726,N_29848);
or UO_767 (O_767,N_29169,N_29113);
and UO_768 (O_768,N_28771,N_29354);
nand UO_769 (O_769,N_29499,N_29778);
nand UO_770 (O_770,N_29614,N_29752);
and UO_771 (O_771,N_28902,N_29831);
or UO_772 (O_772,N_28981,N_29747);
xnor UO_773 (O_773,N_29538,N_29937);
nand UO_774 (O_774,N_28699,N_29774);
xor UO_775 (O_775,N_29717,N_29895);
and UO_776 (O_776,N_28815,N_28750);
xor UO_777 (O_777,N_29273,N_28678);
xnor UO_778 (O_778,N_29567,N_29726);
nand UO_779 (O_779,N_29312,N_29113);
or UO_780 (O_780,N_29531,N_29513);
and UO_781 (O_781,N_28910,N_28710);
and UO_782 (O_782,N_29634,N_28870);
nand UO_783 (O_783,N_28761,N_28780);
nand UO_784 (O_784,N_29243,N_29863);
and UO_785 (O_785,N_28510,N_29767);
nor UO_786 (O_786,N_29794,N_28754);
nand UO_787 (O_787,N_28747,N_28931);
nor UO_788 (O_788,N_29198,N_28721);
or UO_789 (O_789,N_28592,N_28932);
or UO_790 (O_790,N_29465,N_28964);
or UO_791 (O_791,N_29869,N_28576);
and UO_792 (O_792,N_29393,N_29067);
nor UO_793 (O_793,N_29129,N_28562);
or UO_794 (O_794,N_29154,N_28685);
nor UO_795 (O_795,N_28848,N_28859);
nor UO_796 (O_796,N_29033,N_28752);
nand UO_797 (O_797,N_28657,N_29697);
xnor UO_798 (O_798,N_28919,N_29115);
nor UO_799 (O_799,N_29585,N_29567);
and UO_800 (O_800,N_29623,N_29867);
xor UO_801 (O_801,N_29063,N_29541);
and UO_802 (O_802,N_28922,N_29939);
and UO_803 (O_803,N_29209,N_28946);
and UO_804 (O_804,N_28797,N_29076);
xor UO_805 (O_805,N_29577,N_29212);
xor UO_806 (O_806,N_29883,N_28925);
nand UO_807 (O_807,N_29500,N_28587);
or UO_808 (O_808,N_29987,N_29179);
and UO_809 (O_809,N_29397,N_28619);
nor UO_810 (O_810,N_29367,N_29948);
nor UO_811 (O_811,N_28737,N_29189);
xnor UO_812 (O_812,N_28672,N_28791);
xor UO_813 (O_813,N_28583,N_29116);
nand UO_814 (O_814,N_28665,N_28544);
and UO_815 (O_815,N_29101,N_29947);
nand UO_816 (O_816,N_28859,N_28928);
nand UO_817 (O_817,N_28979,N_29882);
nand UO_818 (O_818,N_29052,N_29995);
or UO_819 (O_819,N_29583,N_29289);
and UO_820 (O_820,N_29619,N_29004);
nor UO_821 (O_821,N_29183,N_29574);
or UO_822 (O_822,N_29328,N_28934);
nor UO_823 (O_823,N_29032,N_28924);
or UO_824 (O_824,N_28935,N_28597);
and UO_825 (O_825,N_29437,N_29581);
nor UO_826 (O_826,N_29636,N_28678);
nor UO_827 (O_827,N_29633,N_29952);
nand UO_828 (O_828,N_28760,N_29534);
nand UO_829 (O_829,N_29559,N_29198);
or UO_830 (O_830,N_28923,N_29243);
nor UO_831 (O_831,N_28537,N_28518);
and UO_832 (O_832,N_29407,N_29754);
and UO_833 (O_833,N_28858,N_28773);
nand UO_834 (O_834,N_29634,N_29260);
and UO_835 (O_835,N_29327,N_29764);
and UO_836 (O_836,N_28857,N_28635);
nor UO_837 (O_837,N_29440,N_28527);
xor UO_838 (O_838,N_29089,N_29803);
nor UO_839 (O_839,N_29581,N_29965);
xor UO_840 (O_840,N_29804,N_29470);
nor UO_841 (O_841,N_29390,N_28819);
or UO_842 (O_842,N_29830,N_29820);
or UO_843 (O_843,N_29459,N_29608);
or UO_844 (O_844,N_29175,N_29573);
nand UO_845 (O_845,N_29670,N_29860);
nand UO_846 (O_846,N_29983,N_29102);
and UO_847 (O_847,N_28633,N_28928);
and UO_848 (O_848,N_29246,N_28626);
and UO_849 (O_849,N_29444,N_28974);
nand UO_850 (O_850,N_28731,N_29732);
and UO_851 (O_851,N_29592,N_29635);
nand UO_852 (O_852,N_29277,N_29015);
or UO_853 (O_853,N_29950,N_29164);
nor UO_854 (O_854,N_28884,N_29436);
nand UO_855 (O_855,N_29078,N_29164);
and UO_856 (O_856,N_28863,N_29129);
or UO_857 (O_857,N_29021,N_28640);
nand UO_858 (O_858,N_29539,N_29268);
nand UO_859 (O_859,N_29708,N_29896);
xnor UO_860 (O_860,N_29596,N_29722);
nor UO_861 (O_861,N_29353,N_29577);
xnor UO_862 (O_862,N_29159,N_28523);
nor UO_863 (O_863,N_29211,N_28688);
nor UO_864 (O_864,N_29642,N_28777);
nor UO_865 (O_865,N_29773,N_28629);
xor UO_866 (O_866,N_28818,N_28829);
nand UO_867 (O_867,N_29819,N_28905);
xnor UO_868 (O_868,N_29624,N_29039);
nor UO_869 (O_869,N_29309,N_29762);
nor UO_870 (O_870,N_28650,N_29261);
or UO_871 (O_871,N_29347,N_29636);
xnor UO_872 (O_872,N_28839,N_29048);
nand UO_873 (O_873,N_29953,N_28977);
or UO_874 (O_874,N_29189,N_28555);
nand UO_875 (O_875,N_29873,N_28933);
and UO_876 (O_876,N_29196,N_28775);
nor UO_877 (O_877,N_29267,N_29757);
or UO_878 (O_878,N_29295,N_29864);
nor UO_879 (O_879,N_29614,N_29154);
or UO_880 (O_880,N_29469,N_28904);
xor UO_881 (O_881,N_29637,N_29612);
or UO_882 (O_882,N_28506,N_29839);
nand UO_883 (O_883,N_29603,N_29282);
xnor UO_884 (O_884,N_29678,N_29150);
and UO_885 (O_885,N_29955,N_29659);
and UO_886 (O_886,N_28708,N_29612);
nand UO_887 (O_887,N_29588,N_29319);
nor UO_888 (O_888,N_29361,N_29511);
nor UO_889 (O_889,N_29531,N_28541);
or UO_890 (O_890,N_29723,N_29893);
nand UO_891 (O_891,N_28902,N_29259);
and UO_892 (O_892,N_29925,N_29001);
and UO_893 (O_893,N_28732,N_29469);
and UO_894 (O_894,N_29859,N_28710);
and UO_895 (O_895,N_29786,N_29970);
nor UO_896 (O_896,N_29348,N_28904);
and UO_897 (O_897,N_29305,N_29059);
and UO_898 (O_898,N_29329,N_28819);
or UO_899 (O_899,N_29476,N_29614);
nor UO_900 (O_900,N_28617,N_29992);
or UO_901 (O_901,N_28827,N_29149);
nor UO_902 (O_902,N_29187,N_29938);
or UO_903 (O_903,N_28759,N_29320);
xnor UO_904 (O_904,N_29845,N_29702);
nor UO_905 (O_905,N_29868,N_29626);
nor UO_906 (O_906,N_28640,N_29150);
nor UO_907 (O_907,N_29384,N_29213);
xnor UO_908 (O_908,N_29905,N_29871);
and UO_909 (O_909,N_28658,N_29197);
or UO_910 (O_910,N_29933,N_28800);
nand UO_911 (O_911,N_29357,N_29330);
xnor UO_912 (O_912,N_29800,N_29107);
nand UO_913 (O_913,N_28508,N_29448);
and UO_914 (O_914,N_29997,N_29540);
and UO_915 (O_915,N_29366,N_29462);
nand UO_916 (O_916,N_29046,N_28970);
nor UO_917 (O_917,N_28922,N_29381);
nor UO_918 (O_918,N_28507,N_29206);
nand UO_919 (O_919,N_29909,N_29750);
nor UO_920 (O_920,N_29123,N_28520);
nand UO_921 (O_921,N_29037,N_29732);
and UO_922 (O_922,N_28877,N_29577);
nand UO_923 (O_923,N_29016,N_29798);
nand UO_924 (O_924,N_29210,N_28607);
xor UO_925 (O_925,N_29580,N_28579);
nand UO_926 (O_926,N_29290,N_29589);
nor UO_927 (O_927,N_29865,N_29745);
nand UO_928 (O_928,N_29171,N_29117);
xnor UO_929 (O_929,N_29438,N_29300);
nand UO_930 (O_930,N_29859,N_29256);
or UO_931 (O_931,N_29377,N_29084);
nor UO_932 (O_932,N_29146,N_29498);
nor UO_933 (O_933,N_29648,N_29218);
nor UO_934 (O_934,N_28538,N_29827);
or UO_935 (O_935,N_29169,N_29933);
xor UO_936 (O_936,N_28591,N_29545);
and UO_937 (O_937,N_28715,N_29575);
and UO_938 (O_938,N_29265,N_29957);
and UO_939 (O_939,N_28969,N_29909);
or UO_940 (O_940,N_28718,N_29861);
or UO_941 (O_941,N_29276,N_29067);
nor UO_942 (O_942,N_29961,N_29418);
nor UO_943 (O_943,N_28897,N_28637);
xor UO_944 (O_944,N_29435,N_28965);
and UO_945 (O_945,N_28796,N_29860);
nand UO_946 (O_946,N_29245,N_29673);
or UO_947 (O_947,N_29791,N_28817);
nand UO_948 (O_948,N_28749,N_28755);
and UO_949 (O_949,N_29434,N_29075);
nor UO_950 (O_950,N_29822,N_29668);
and UO_951 (O_951,N_29963,N_28874);
nor UO_952 (O_952,N_29229,N_29612);
and UO_953 (O_953,N_29415,N_28915);
nand UO_954 (O_954,N_29020,N_29205);
or UO_955 (O_955,N_29479,N_29610);
xor UO_956 (O_956,N_29765,N_29135);
and UO_957 (O_957,N_28769,N_29452);
nor UO_958 (O_958,N_28597,N_29357);
nor UO_959 (O_959,N_29128,N_29805);
xor UO_960 (O_960,N_29153,N_28715);
nand UO_961 (O_961,N_28981,N_29112);
nand UO_962 (O_962,N_29518,N_29131);
or UO_963 (O_963,N_28608,N_28585);
or UO_964 (O_964,N_29404,N_29320);
nand UO_965 (O_965,N_28724,N_28902);
nand UO_966 (O_966,N_29185,N_28526);
or UO_967 (O_967,N_29585,N_29059);
nand UO_968 (O_968,N_29978,N_29425);
nor UO_969 (O_969,N_29926,N_29817);
nor UO_970 (O_970,N_28608,N_28562);
nand UO_971 (O_971,N_29518,N_29683);
xor UO_972 (O_972,N_28650,N_29556);
nor UO_973 (O_973,N_29280,N_28932);
xor UO_974 (O_974,N_29442,N_28809);
xor UO_975 (O_975,N_29373,N_28536);
nor UO_976 (O_976,N_29094,N_29043);
and UO_977 (O_977,N_28622,N_29184);
and UO_978 (O_978,N_29021,N_28536);
nor UO_979 (O_979,N_28705,N_29599);
and UO_980 (O_980,N_29170,N_29537);
nand UO_981 (O_981,N_29688,N_28533);
xor UO_982 (O_982,N_28519,N_28748);
nand UO_983 (O_983,N_29387,N_29579);
xor UO_984 (O_984,N_28683,N_29636);
and UO_985 (O_985,N_28614,N_28974);
nand UO_986 (O_986,N_29243,N_29130);
xnor UO_987 (O_987,N_29327,N_29486);
or UO_988 (O_988,N_29781,N_29566);
and UO_989 (O_989,N_29612,N_28559);
xor UO_990 (O_990,N_29208,N_29719);
or UO_991 (O_991,N_29904,N_29310);
or UO_992 (O_992,N_29420,N_29406);
xor UO_993 (O_993,N_29801,N_28502);
and UO_994 (O_994,N_29502,N_29007);
nor UO_995 (O_995,N_28822,N_28951);
or UO_996 (O_996,N_29134,N_28826);
xnor UO_997 (O_997,N_28787,N_29305);
nor UO_998 (O_998,N_29246,N_29636);
xnor UO_999 (O_999,N_29609,N_28620);
or UO_1000 (O_1000,N_29647,N_28943);
or UO_1001 (O_1001,N_29575,N_29659);
and UO_1002 (O_1002,N_28878,N_29037);
and UO_1003 (O_1003,N_28975,N_28641);
xor UO_1004 (O_1004,N_29516,N_29434);
nor UO_1005 (O_1005,N_29261,N_29173);
and UO_1006 (O_1006,N_29091,N_29590);
and UO_1007 (O_1007,N_28617,N_28776);
nand UO_1008 (O_1008,N_28710,N_29540);
or UO_1009 (O_1009,N_28743,N_29475);
or UO_1010 (O_1010,N_29418,N_28578);
and UO_1011 (O_1011,N_28651,N_28697);
or UO_1012 (O_1012,N_29803,N_29433);
and UO_1013 (O_1013,N_29265,N_29174);
xnor UO_1014 (O_1014,N_29483,N_29893);
xor UO_1015 (O_1015,N_29580,N_29288);
or UO_1016 (O_1016,N_28829,N_28845);
nand UO_1017 (O_1017,N_29310,N_28754);
and UO_1018 (O_1018,N_29531,N_28848);
nand UO_1019 (O_1019,N_29792,N_29485);
nor UO_1020 (O_1020,N_28921,N_29933);
or UO_1021 (O_1021,N_29723,N_29628);
nand UO_1022 (O_1022,N_29378,N_28762);
or UO_1023 (O_1023,N_29853,N_29687);
nand UO_1024 (O_1024,N_29786,N_29865);
nor UO_1025 (O_1025,N_29912,N_29746);
nand UO_1026 (O_1026,N_29258,N_29331);
and UO_1027 (O_1027,N_28691,N_29244);
nor UO_1028 (O_1028,N_29982,N_29085);
and UO_1029 (O_1029,N_29770,N_29507);
or UO_1030 (O_1030,N_29685,N_29214);
nor UO_1031 (O_1031,N_28749,N_29102);
or UO_1032 (O_1032,N_29553,N_28858);
or UO_1033 (O_1033,N_29490,N_28937);
nor UO_1034 (O_1034,N_29764,N_29803);
nand UO_1035 (O_1035,N_29459,N_29974);
and UO_1036 (O_1036,N_29710,N_28733);
nor UO_1037 (O_1037,N_29257,N_29359);
and UO_1038 (O_1038,N_29698,N_29853);
nand UO_1039 (O_1039,N_29315,N_28689);
nor UO_1040 (O_1040,N_28726,N_29743);
nand UO_1041 (O_1041,N_29548,N_29889);
nor UO_1042 (O_1042,N_29806,N_29423);
nor UO_1043 (O_1043,N_29666,N_29008);
xor UO_1044 (O_1044,N_29699,N_28816);
nor UO_1045 (O_1045,N_29001,N_28982);
nor UO_1046 (O_1046,N_29359,N_28562);
nor UO_1047 (O_1047,N_29307,N_28650);
nor UO_1048 (O_1048,N_29042,N_29999);
nand UO_1049 (O_1049,N_29079,N_28854);
nor UO_1050 (O_1050,N_29942,N_28696);
nor UO_1051 (O_1051,N_29915,N_29037);
or UO_1052 (O_1052,N_28764,N_28710);
nor UO_1053 (O_1053,N_29483,N_29756);
or UO_1054 (O_1054,N_28542,N_29859);
xor UO_1055 (O_1055,N_28941,N_28716);
xor UO_1056 (O_1056,N_29128,N_29801);
nand UO_1057 (O_1057,N_28927,N_28562);
nor UO_1058 (O_1058,N_29339,N_29472);
or UO_1059 (O_1059,N_28887,N_29718);
or UO_1060 (O_1060,N_29431,N_28794);
nor UO_1061 (O_1061,N_29462,N_29641);
nor UO_1062 (O_1062,N_29050,N_29027);
or UO_1063 (O_1063,N_29197,N_29740);
nand UO_1064 (O_1064,N_29327,N_28899);
nand UO_1065 (O_1065,N_28615,N_29333);
or UO_1066 (O_1066,N_29324,N_29060);
nor UO_1067 (O_1067,N_28975,N_29945);
xor UO_1068 (O_1068,N_29552,N_29339);
or UO_1069 (O_1069,N_28750,N_29562);
or UO_1070 (O_1070,N_28883,N_29934);
or UO_1071 (O_1071,N_28770,N_29991);
nor UO_1072 (O_1072,N_29403,N_29645);
xnor UO_1073 (O_1073,N_29105,N_29028);
nor UO_1074 (O_1074,N_29834,N_29271);
nor UO_1075 (O_1075,N_29101,N_29761);
or UO_1076 (O_1076,N_28684,N_28512);
nand UO_1077 (O_1077,N_29147,N_29019);
xnor UO_1078 (O_1078,N_28617,N_29349);
xnor UO_1079 (O_1079,N_29427,N_29585);
xor UO_1080 (O_1080,N_29104,N_29393);
xor UO_1081 (O_1081,N_28683,N_28590);
xnor UO_1082 (O_1082,N_28537,N_28649);
or UO_1083 (O_1083,N_29256,N_29148);
or UO_1084 (O_1084,N_28582,N_28911);
and UO_1085 (O_1085,N_29347,N_29527);
and UO_1086 (O_1086,N_29537,N_29514);
nor UO_1087 (O_1087,N_29024,N_29217);
or UO_1088 (O_1088,N_28687,N_28593);
and UO_1089 (O_1089,N_28528,N_29996);
and UO_1090 (O_1090,N_28788,N_29383);
nor UO_1091 (O_1091,N_28929,N_29484);
nand UO_1092 (O_1092,N_29586,N_29906);
and UO_1093 (O_1093,N_28525,N_29302);
or UO_1094 (O_1094,N_29295,N_29911);
nor UO_1095 (O_1095,N_29194,N_28552);
nand UO_1096 (O_1096,N_28609,N_29921);
nor UO_1097 (O_1097,N_29783,N_28824);
nor UO_1098 (O_1098,N_29543,N_28786);
xnor UO_1099 (O_1099,N_29203,N_29441);
nor UO_1100 (O_1100,N_29764,N_29432);
xnor UO_1101 (O_1101,N_28567,N_29933);
or UO_1102 (O_1102,N_28907,N_29241);
or UO_1103 (O_1103,N_28654,N_29217);
nand UO_1104 (O_1104,N_28728,N_28710);
nor UO_1105 (O_1105,N_29300,N_28700);
and UO_1106 (O_1106,N_29350,N_29811);
nor UO_1107 (O_1107,N_29112,N_29448);
and UO_1108 (O_1108,N_28595,N_28834);
and UO_1109 (O_1109,N_28555,N_29436);
and UO_1110 (O_1110,N_28727,N_29859);
nor UO_1111 (O_1111,N_29466,N_29560);
or UO_1112 (O_1112,N_29773,N_29739);
nor UO_1113 (O_1113,N_28981,N_28728);
or UO_1114 (O_1114,N_28839,N_29289);
nor UO_1115 (O_1115,N_29376,N_29614);
or UO_1116 (O_1116,N_28972,N_29049);
nand UO_1117 (O_1117,N_28896,N_29454);
nand UO_1118 (O_1118,N_29127,N_29624);
or UO_1119 (O_1119,N_29676,N_29677);
xor UO_1120 (O_1120,N_28793,N_29286);
xor UO_1121 (O_1121,N_28777,N_28774);
xor UO_1122 (O_1122,N_28589,N_29349);
nor UO_1123 (O_1123,N_29615,N_28618);
nand UO_1124 (O_1124,N_29681,N_29189);
or UO_1125 (O_1125,N_29024,N_29206);
xnor UO_1126 (O_1126,N_28636,N_28565);
or UO_1127 (O_1127,N_29303,N_28850);
or UO_1128 (O_1128,N_29660,N_28770);
nor UO_1129 (O_1129,N_29822,N_29760);
and UO_1130 (O_1130,N_29473,N_28702);
and UO_1131 (O_1131,N_29872,N_29489);
or UO_1132 (O_1132,N_29888,N_29687);
nand UO_1133 (O_1133,N_29793,N_29712);
nand UO_1134 (O_1134,N_29230,N_29116);
nor UO_1135 (O_1135,N_28731,N_29803);
nand UO_1136 (O_1136,N_29135,N_29035);
nand UO_1137 (O_1137,N_29316,N_29613);
nor UO_1138 (O_1138,N_29398,N_29013);
xor UO_1139 (O_1139,N_28854,N_29783);
xor UO_1140 (O_1140,N_29291,N_29868);
and UO_1141 (O_1141,N_28923,N_28621);
and UO_1142 (O_1142,N_29532,N_29221);
and UO_1143 (O_1143,N_28945,N_28732);
xnor UO_1144 (O_1144,N_28980,N_29604);
and UO_1145 (O_1145,N_28900,N_28765);
or UO_1146 (O_1146,N_29408,N_28897);
nor UO_1147 (O_1147,N_28583,N_28921);
or UO_1148 (O_1148,N_28826,N_29174);
and UO_1149 (O_1149,N_28992,N_29549);
nand UO_1150 (O_1150,N_29374,N_29971);
and UO_1151 (O_1151,N_29481,N_28545);
nand UO_1152 (O_1152,N_28561,N_29522);
and UO_1153 (O_1153,N_29336,N_28917);
nand UO_1154 (O_1154,N_28694,N_29961);
and UO_1155 (O_1155,N_29851,N_29935);
nand UO_1156 (O_1156,N_29970,N_29981);
and UO_1157 (O_1157,N_29907,N_29089);
nand UO_1158 (O_1158,N_29839,N_28655);
and UO_1159 (O_1159,N_28753,N_28519);
nor UO_1160 (O_1160,N_28823,N_29758);
or UO_1161 (O_1161,N_29567,N_28998);
nand UO_1162 (O_1162,N_29793,N_29183);
xor UO_1163 (O_1163,N_29980,N_29827);
or UO_1164 (O_1164,N_29464,N_29648);
or UO_1165 (O_1165,N_29163,N_29340);
nor UO_1166 (O_1166,N_29722,N_29941);
nand UO_1167 (O_1167,N_28847,N_29094);
nand UO_1168 (O_1168,N_29884,N_29040);
nor UO_1169 (O_1169,N_28897,N_29152);
and UO_1170 (O_1170,N_29995,N_29414);
or UO_1171 (O_1171,N_29935,N_29107);
xor UO_1172 (O_1172,N_28586,N_29585);
xnor UO_1173 (O_1173,N_28681,N_29234);
nand UO_1174 (O_1174,N_28736,N_28510);
or UO_1175 (O_1175,N_28923,N_29624);
or UO_1176 (O_1176,N_28999,N_29750);
nand UO_1177 (O_1177,N_29694,N_28579);
and UO_1178 (O_1178,N_29934,N_29472);
xor UO_1179 (O_1179,N_28766,N_28651);
or UO_1180 (O_1180,N_28774,N_29850);
nand UO_1181 (O_1181,N_29301,N_29185);
xnor UO_1182 (O_1182,N_29984,N_29136);
and UO_1183 (O_1183,N_28681,N_28753);
nor UO_1184 (O_1184,N_28688,N_28642);
and UO_1185 (O_1185,N_29246,N_28533);
or UO_1186 (O_1186,N_29141,N_29543);
nor UO_1187 (O_1187,N_29538,N_28709);
nor UO_1188 (O_1188,N_29466,N_28504);
nand UO_1189 (O_1189,N_28601,N_29430);
nand UO_1190 (O_1190,N_29386,N_28969);
and UO_1191 (O_1191,N_28584,N_29187);
nor UO_1192 (O_1192,N_29507,N_29429);
or UO_1193 (O_1193,N_28509,N_28754);
xor UO_1194 (O_1194,N_29635,N_29995);
or UO_1195 (O_1195,N_29318,N_29721);
nand UO_1196 (O_1196,N_28558,N_29121);
or UO_1197 (O_1197,N_28800,N_29106);
nor UO_1198 (O_1198,N_29896,N_28798);
xor UO_1199 (O_1199,N_28916,N_29821);
nand UO_1200 (O_1200,N_28519,N_28906);
nand UO_1201 (O_1201,N_28793,N_28886);
nand UO_1202 (O_1202,N_29749,N_28568);
nor UO_1203 (O_1203,N_29417,N_29318);
nand UO_1204 (O_1204,N_28554,N_29565);
and UO_1205 (O_1205,N_29857,N_29798);
xnor UO_1206 (O_1206,N_28852,N_29209);
or UO_1207 (O_1207,N_29213,N_29930);
or UO_1208 (O_1208,N_28921,N_29931);
nand UO_1209 (O_1209,N_29739,N_29005);
and UO_1210 (O_1210,N_28757,N_28844);
nand UO_1211 (O_1211,N_29485,N_29609);
and UO_1212 (O_1212,N_29749,N_29924);
xnor UO_1213 (O_1213,N_28774,N_29515);
and UO_1214 (O_1214,N_28538,N_28536);
xor UO_1215 (O_1215,N_29224,N_28597);
and UO_1216 (O_1216,N_29518,N_29087);
xnor UO_1217 (O_1217,N_28505,N_28587);
nor UO_1218 (O_1218,N_29527,N_29682);
nand UO_1219 (O_1219,N_29507,N_29027);
xnor UO_1220 (O_1220,N_29172,N_29745);
and UO_1221 (O_1221,N_29822,N_29770);
and UO_1222 (O_1222,N_29681,N_29297);
nand UO_1223 (O_1223,N_29407,N_29036);
nand UO_1224 (O_1224,N_29301,N_28600);
or UO_1225 (O_1225,N_29051,N_29665);
xnor UO_1226 (O_1226,N_29339,N_29213);
xor UO_1227 (O_1227,N_28661,N_29149);
and UO_1228 (O_1228,N_29265,N_29583);
and UO_1229 (O_1229,N_29241,N_29233);
and UO_1230 (O_1230,N_29488,N_29798);
nor UO_1231 (O_1231,N_29133,N_29701);
xor UO_1232 (O_1232,N_29862,N_28600);
and UO_1233 (O_1233,N_29117,N_29443);
or UO_1234 (O_1234,N_28906,N_29817);
or UO_1235 (O_1235,N_29297,N_29508);
xor UO_1236 (O_1236,N_28528,N_29371);
xnor UO_1237 (O_1237,N_28952,N_29280);
nand UO_1238 (O_1238,N_29343,N_28918);
nand UO_1239 (O_1239,N_28634,N_29134);
or UO_1240 (O_1240,N_29186,N_29750);
and UO_1241 (O_1241,N_29190,N_29748);
nand UO_1242 (O_1242,N_29624,N_28836);
nand UO_1243 (O_1243,N_28912,N_29712);
or UO_1244 (O_1244,N_29991,N_29421);
and UO_1245 (O_1245,N_29242,N_29738);
nand UO_1246 (O_1246,N_28960,N_28888);
xor UO_1247 (O_1247,N_29393,N_28751);
or UO_1248 (O_1248,N_29120,N_29426);
nor UO_1249 (O_1249,N_29889,N_28675);
xor UO_1250 (O_1250,N_29804,N_28778);
or UO_1251 (O_1251,N_29478,N_28554);
xor UO_1252 (O_1252,N_28653,N_29881);
and UO_1253 (O_1253,N_29796,N_29762);
and UO_1254 (O_1254,N_28528,N_28832);
or UO_1255 (O_1255,N_29143,N_29699);
and UO_1256 (O_1256,N_29059,N_29537);
nor UO_1257 (O_1257,N_28912,N_29193);
and UO_1258 (O_1258,N_28584,N_29489);
or UO_1259 (O_1259,N_28636,N_29832);
nand UO_1260 (O_1260,N_28644,N_28928);
and UO_1261 (O_1261,N_28650,N_29623);
nand UO_1262 (O_1262,N_29915,N_29275);
nand UO_1263 (O_1263,N_28939,N_29013);
nand UO_1264 (O_1264,N_29366,N_29021);
nand UO_1265 (O_1265,N_29905,N_29776);
xor UO_1266 (O_1266,N_29917,N_29177);
nand UO_1267 (O_1267,N_29432,N_29327);
and UO_1268 (O_1268,N_29725,N_28547);
or UO_1269 (O_1269,N_28616,N_29545);
nand UO_1270 (O_1270,N_29882,N_29903);
and UO_1271 (O_1271,N_29516,N_29888);
xnor UO_1272 (O_1272,N_28679,N_29719);
and UO_1273 (O_1273,N_29518,N_29001);
nand UO_1274 (O_1274,N_29173,N_28937);
nand UO_1275 (O_1275,N_29044,N_28899);
xnor UO_1276 (O_1276,N_28920,N_29925);
nor UO_1277 (O_1277,N_29690,N_29691);
nor UO_1278 (O_1278,N_29629,N_29212);
or UO_1279 (O_1279,N_29845,N_29523);
nand UO_1280 (O_1280,N_29964,N_28914);
and UO_1281 (O_1281,N_29536,N_28863);
or UO_1282 (O_1282,N_29627,N_29674);
or UO_1283 (O_1283,N_28676,N_29606);
xor UO_1284 (O_1284,N_29303,N_28547);
and UO_1285 (O_1285,N_29179,N_28699);
nor UO_1286 (O_1286,N_28875,N_29035);
nand UO_1287 (O_1287,N_29917,N_29503);
xnor UO_1288 (O_1288,N_29722,N_29735);
nand UO_1289 (O_1289,N_29812,N_28728);
xor UO_1290 (O_1290,N_29812,N_29957);
nor UO_1291 (O_1291,N_29827,N_28805);
nand UO_1292 (O_1292,N_29392,N_28537);
and UO_1293 (O_1293,N_28773,N_29554);
nor UO_1294 (O_1294,N_29249,N_28961);
xnor UO_1295 (O_1295,N_28958,N_29485);
xor UO_1296 (O_1296,N_29437,N_28514);
or UO_1297 (O_1297,N_29354,N_28990);
nor UO_1298 (O_1298,N_28505,N_28709);
nand UO_1299 (O_1299,N_28908,N_29171);
xnor UO_1300 (O_1300,N_29874,N_29017);
xor UO_1301 (O_1301,N_28872,N_29798);
and UO_1302 (O_1302,N_29440,N_29165);
and UO_1303 (O_1303,N_29726,N_29705);
nor UO_1304 (O_1304,N_28858,N_29364);
or UO_1305 (O_1305,N_29641,N_28780);
nand UO_1306 (O_1306,N_28501,N_29993);
xnor UO_1307 (O_1307,N_29619,N_29330);
nand UO_1308 (O_1308,N_29487,N_28613);
nand UO_1309 (O_1309,N_29771,N_28902);
and UO_1310 (O_1310,N_29338,N_28680);
or UO_1311 (O_1311,N_29423,N_28660);
nand UO_1312 (O_1312,N_29531,N_29108);
and UO_1313 (O_1313,N_29903,N_29129);
nor UO_1314 (O_1314,N_29039,N_28514);
xnor UO_1315 (O_1315,N_29701,N_28723);
nand UO_1316 (O_1316,N_28948,N_28924);
nand UO_1317 (O_1317,N_28587,N_28750);
nor UO_1318 (O_1318,N_29864,N_28533);
nor UO_1319 (O_1319,N_29450,N_29183);
or UO_1320 (O_1320,N_28525,N_29218);
xnor UO_1321 (O_1321,N_28718,N_29587);
nor UO_1322 (O_1322,N_29665,N_28644);
nor UO_1323 (O_1323,N_29918,N_29657);
and UO_1324 (O_1324,N_29436,N_28904);
nor UO_1325 (O_1325,N_29053,N_29362);
nand UO_1326 (O_1326,N_29175,N_28787);
nand UO_1327 (O_1327,N_29787,N_29223);
nand UO_1328 (O_1328,N_29690,N_28675);
nor UO_1329 (O_1329,N_28846,N_29935);
or UO_1330 (O_1330,N_29478,N_29636);
and UO_1331 (O_1331,N_29905,N_28752);
xor UO_1332 (O_1332,N_29152,N_29468);
xnor UO_1333 (O_1333,N_28759,N_28559);
nand UO_1334 (O_1334,N_29352,N_29024);
nor UO_1335 (O_1335,N_29445,N_29401);
or UO_1336 (O_1336,N_29132,N_29082);
or UO_1337 (O_1337,N_29567,N_29879);
xor UO_1338 (O_1338,N_29713,N_29749);
xnor UO_1339 (O_1339,N_28703,N_29282);
or UO_1340 (O_1340,N_28886,N_29614);
nand UO_1341 (O_1341,N_28720,N_28766);
and UO_1342 (O_1342,N_29990,N_29657);
and UO_1343 (O_1343,N_29882,N_29601);
or UO_1344 (O_1344,N_28793,N_29666);
xor UO_1345 (O_1345,N_29572,N_29347);
nor UO_1346 (O_1346,N_29272,N_29182);
xor UO_1347 (O_1347,N_29168,N_29761);
and UO_1348 (O_1348,N_29779,N_29588);
or UO_1349 (O_1349,N_29092,N_28749);
nor UO_1350 (O_1350,N_29330,N_29280);
nand UO_1351 (O_1351,N_29348,N_28627);
or UO_1352 (O_1352,N_28771,N_28881);
nand UO_1353 (O_1353,N_29422,N_29031);
or UO_1354 (O_1354,N_29199,N_29041);
or UO_1355 (O_1355,N_29605,N_29478);
or UO_1356 (O_1356,N_29627,N_28725);
or UO_1357 (O_1357,N_28511,N_28876);
or UO_1358 (O_1358,N_29595,N_29168);
and UO_1359 (O_1359,N_29385,N_29947);
xor UO_1360 (O_1360,N_29974,N_29451);
nand UO_1361 (O_1361,N_28934,N_29702);
or UO_1362 (O_1362,N_29343,N_29164);
nor UO_1363 (O_1363,N_29158,N_29873);
or UO_1364 (O_1364,N_29966,N_29567);
nor UO_1365 (O_1365,N_29826,N_29252);
nand UO_1366 (O_1366,N_29175,N_29504);
and UO_1367 (O_1367,N_29117,N_28551);
nor UO_1368 (O_1368,N_29693,N_28657);
nand UO_1369 (O_1369,N_28985,N_28872);
and UO_1370 (O_1370,N_28565,N_29340);
and UO_1371 (O_1371,N_29413,N_29227);
and UO_1372 (O_1372,N_29897,N_28875);
xnor UO_1373 (O_1373,N_28666,N_29180);
xor UO_1374 (O_1374,N_29497,N_29977);
xnor UO_1375 (O_1375,N_28714,N_29258);
nor UO_1376 (O_1376,N_29714,N_28880);
nand UO_1377 (O_1377,N_28779,N_29198);
xor UO_1378 (O_1378,N_28525,N_29624);
nor UO_1379 (O_1379,N_28935,N_29494);
and UO_1380 (O_1380,N_29921,N_29309);
xnor UO_1381 (O_1381,N_29880,N_29914);
nand UO_1382 (O_1382,N_28981,N_28757);
and UO_1383 (O_1383,N_29556,N_29912);
and UO_1384 (O_1384,N_28776,N_29678);
nor UO_1385 (O_1385,N_29156,N_29579);
xor UO_1386 (O_1386,N_28811,N_29599);
or UO_1387 (O_1387,N_29091,N_28830);
xor UO_1388 (O_1388,N_28511,N_29565);
nand UO_1389 (O_1389,N_28968,N_29908);
or UO_1390 (O_1390,N_29327,N_28882);
nor UO_1391 (O_1391,N_28833,N_29136);
and UO_1392 (O_1392,N_29255,N_28769);
nor UO_1393 (O_1393,N_29623,N_29015);
and UO_1394 (O_1394,N_28938,N_28751);
and UO_1395 (O_1395,N_28620,N_29490);
or UO_1396 (O_1396,N_29967,N_29278);
nand UO_1397 (O_1397,N_28776,N_29335);
nand UO_1398 (O_1398,N_29414,N_29627);
xor UO_1399 (O_1399,N_29305,N_29747);
or UO_1400 (O_1400,N_29856,N_28805);
and UO_1401 (O_1401,N_28667,N_28799);
nand UO_1402 (O_1402,N_29771,N_29459);
xor UO_1403 (O_1403,N_29286,N_28909);
nor UO_1404 (O_1404,N_29154,N_28820);
or UO_1405 (O_1405,N_29354,N_29852);
nor UO_1406 (O_1406,N_28802,N_29751);
nor UO_1407 (O_1407,N_28754,N_28666);
and UO_1408 (O_1408,N_29590,N_29066);
or UO_1409 (O_1409,N_29310,N_29386);
and UO_1410 (O_1410,N_28677,N_28644);
xor UO_1411 (O_1411,N_29956,N_28652);
xor UO_1412 (O_1412,N_29270,N_28935);
and UO_1413 (O_1413,N_29766,N_29081);
nor UO_1414 (O_1414,N_29037,N_29560);
xnor UO_1415 (O_1415,N_29427,N_29382);
nand UO_1416 (O_1416,N_29947,N_29150);
xnor UO_1417 (O_1417,N_28855,N_29639);
xnor UO_1418 (O_1418,N_29955,N_29562);
and UO_1419 (O_1419,N_28944,N_29331);
and UO_1420 (O_1420,N_29802,N_28512);
and UO_1421 (O_1421,N_28720,N_29527);
or UO_1422 (O_1422,N_29779,N_29450);
xor UO_1423 (O_1423,N_28879,N_29435);
or UO_1424 (O_1424,N_29013,N_28796);
and UO_1425 (O_1425,N_29960,N_29720);
nand UO_1426 (O_1426,N_29797,N_28649);
nand UO_1427 (O_1427,N_28823,N_28899);
xnor UO_1428 (O_1428,N_29266,N_29634);
nand UO_1429 (O_1429,N_29220,N_28506);
xor UO_1430 (O_1430,N_29153,N_29255);
and UO_1431 (O_1431,N_28807,N_29539);
nand UO_1432 (O_1432,N_28961,N_29124);
and UO_1433 (O_1433,N_29703,N_29199);
or UO_1434 (O_1434,N_29618,N_29728);
nor UO_1435 (O_1435,N_28664,N_28964);
nand UO_1436 (O_1436,N_29731,N_28660);
nand UO_1437 (O_1437,N_28877,N_29807);
nand UO_1438 (O_1438,N_28851,N_28884);
nor UO_1439 (O_1439,N_29698,N_29861);
and UO_1440 (O_1440,N_29103,N_29447);
nand UO_1441 (O_1441,N_28616,N_29930);
and UO_1442 (O_1442,N_29520,N_29889);
nor UO_1443 (O_1443,N_29892,N_29639);
and UO_1444 (O_1444,N_28550,N_29378);
xnor UO_1445 (O_1445,N_28519,N_28667);
nand UO_1446 (O_1446,N_29396,N_29474);
nand UO_1447 (O_1447,N_29606,N_29616);
nand UO_1448 (O_1448,N_29106,N_29311);
or UO_1449 (O_1449,N_29923,N_28813);
nand UO_1450 (O_1450,N_29568,N_29707);
nor UO_1451 (O_1451,N_29450,N_28784);
or UO_1452 (O_1452,N_28553,N_29487);
nand UO_1453 (O_1453,N_28721,N_28635);
nand UO_1454 (O_1454,N_29158,N_29117);
or UO_1455 (O_1455,N_28716,N_29710);
or UO_1456 (O_1456,N_28701,N_29670);
and UO_1457 (O_1457,N_29407,N_28565);
and UO_1458 (O_1458,N_29866,N_29296);
or UO_1459 (O_1459,N_29884,N_29449);
and UO_1460 (O_1460,N_29719,N_29665);
or UO_1461 (O_1461,N_29063,N_28820);
xor UO_1462 (O_1462,N_28997,N_29205);
nand UO_1463 (O_1463,N_29903,N_28871);
nand UO_1464 (O_1464,N_29869,N_29641);
xnor UO_1465 (O_1465,N_28845,N_29660);
xor UO_1466 (O_1466,N_28534,N_29584);
or UO_1467 (O_1467,N_29347,N_28990);
nand UO_1468 (O_1468,N_29006,N_29518);
nor UO_1469 (O_1469,N_29593,N_29524);
xor UO_1470 (O_1470,N_29275,N_28551);
or UO_1471 (O_1471,N_29058,N_28595);
xnor UO_1472 (O_1472,N_29561,N_29837);
or UO_1473 (O_1473,N_29124,N_29767);
or UO_1474 (O_1474,N_29886,N_29739);
xnor UO_1475 (O_1475,N_29299,N_29581);
nor UO_1476 (O_1476,N_29949,N_28638);
xor UO_1477 (O_1477,N_29839,N_28640);
xor UO_1478 (O_1478,N_29520,N_29010);
and UO_1479 (O_1479,N_29265,N_29420);
nor UO_1480 (O_1480,N_28922,N_29114);
nand UO_1481 (O_1481,N_29487,N_29858);
and UO_1482 (O_1482,N_29202,N_29321);
nor UO_1483 (O_1483,N_29591,N_29493);
xor UO_1484 (O_1484,N_29608,N_29823);
xor UO_1485 (O_1485,N_29294,N_29063);
or UO_1486 (O_1486,N_28829,N_29094);
or UO_1487 (O_1487,N_29436,N_29953);
nor UO_1488 (O_1488,N_29495,N_28551);
nand UO_1489 (O_1489,N_29902,N_28551);
or UO_1490 (O_1490,N_28823,N_29488);
nand UO_1491 (O_1491,N_29016,N_28698);
nand UO_1492 (O_1492,N_29361,N_28893);
xor UO_1493 (O_1493,N_29598,N_29646);
nor UO_1494 (O_1494,N_29844,N_29332);
or UO_1495 (O_1495,N_28852,N_29285);
and UO_1496 (O_1496,N_28566,N_29210);
and UO_1497 (O_1497,N_28889,N_29278);
nor UO_1498 (O_1498,N_29455,N_29174);
nor UO_1499 (O_1499,N_29533,N_28731);
nor UO_1500 (O_1500,N_28952,N_29450);
nor UO_1501 (O_1501,N_29947,N_29027);
nor UO_1502 (O_1502,N_28927,N_29688);
nand UO_1503 (O_1503,N_29792,N_29521);
or UO_1504 (O_1504,N_28883,N_28553);
and UO_1505 (O_1505,N_28843,N_29071);
or UO_1506 (O_1506,N_28501,N_29480);
nand UO_1507 (O_1507,N_29985,N_29732);
and UO_1508 (O_1508,N_28674,N_29470);
nor UO_1509 (O_1509,N_28746,N_29817);
and UO_1510 (O_1510,N_29386,N_29607);
or UO_1511 (O_1511,N_29251,N_29770);
xnor UO_1512 (O_1512,N_29032,N_29825);
nand UO_1513 (O_1513,N_29806,N_28673);
xnor UO_1514 (O_1514,N_28768,N_29654);
nand UO_1515 (O_1515,N_29985,N_28832);
and UO_1516 (O_1516,N_29395,N_29765);
nor UO_1517 (O_1517,N_29467,N_29555);
xor UO_1518 (O_1518,N_29403,N_28907);
xor UO_1519 (O_1519,N_29330,N_28867);
nand UO_1520 (O_1520,N_29562,N_28791);
nor UO_1521 (O_1521,N_29136,N_28853);
nand UO_1522 (O_1522,N_29026,N_28918);
xor UO_1523 (O_1523,N_28795,N_28727);
and UO_1524 (O_1524,N_28536,N_28682);
nand UO_1525 (O_1525,N_29585,N_28733);
or UO_1526 (O_1526,N_28718,N_29038);
nor UO_1527 (O_1527,N_29969,N_28880);
or UO_1528 (O_1528,N_29557,N_28505);
nor UO_1529 (O_1529,N_29911,N_29330);
xor UO_1530 (O_1530,N_29370,N_29585);
nand UO_1531 (O_1531,N_28880,N_29037);
nor UO_1532 (O_1532,N_29983,N_29547);
or UO_1533 (O_1533,N_28819,N_28748);
nor UO_1534 (O_1534,N_29511,N_28840);
xor UO_1535 (O_1535,N_29779,N_29488);
or UO_1536 (O_1536,N_29400,N_29641);
or UO_1537 (O_1537,N_28794,N_29907);
xor UO_1538 (O_1538,N_28821,N_29705);
or UO_1539 (O_1539,N_29326,N_29791);
xnor UO_1540 (O_1540,N_29428,N_29129);
or UO_1541 (O_1541,N_28799,N_29259);
nand UO_1542 (O_1542,N_29512,N_29810);
nand UO_1543 (O_1543,N_29767,N_29913);
and UO_1544 (O_1544,N_29158,N_29060);
or UO_1545 (O_1545,N_29978,N_29414);
or UO_1546 (O_1546,N_29840,N_29033);
xor UO_1547 (O_1547,N_28786,N_29181);
xnor UO_1548 (O_1548,N_29340,N_29472);
or UO_1549 (O_1549,N_29052,N_29181);
or UO_1550 (O_1550,N_28647,N_29630);
nor UO_1551 (O_1551,N_28764,N_29520);
or UO_1552 (O_1552,N_29911,N_29962);
xor UO_1553 (O_1553,N_28908,N_29352);
nand UO_1554 (O_1554,N_29586,N_29462);
xnor UO_1555 (O_1555,N_29257,N_29009);
xor UO_1556 (O_1556,N_29692,N_29006);
nand UO_1557 (O_1557,N_28550,N_29857);
and UO_1558 (O_1558,N_29833,N_29406);
or UO_1559 (O_1559,N_28866,N_29439);
nand UO_1560 (O_1560,N_28526,N_29657);
nor UO_1561 (O_1561,N_29281,N_28920);
xnor UO_1562 (O_1562,N_29406,N_29220);
and UO_1563 (O_1563,N_28682,N_29344);
nor UO_1564 (O_1564,N_29486,N_29986);
or UO_1565 (O_1565,N_29019,N_29673);
and UO_1566 (O_1566,N_28733,N_28866);
or UO_1567 (O_1567,N_29680,N_29093);
nand UO_1568 (O_1568,N_29425,N_28670);
or UO_1569 (O_1569,N_29936,N_28628);
or UO_1570 (O_1570,N_28976,N_29871);
nor UO_1571 (O_1571,N_29910,N_28928);
xor UO_1572 (O_1572,N_29547,N_29283);
and UO_1573 (O_1573,N_29573,N_29960);
or UO_1574 (O_1574,N_28742,N_28902);
xnor UO_1575 (O_1575,N_28690,N_29137);
nor UO_1576 (O_1576,N_28993,N_28865);
or UO_1577 (O_1577,N_29516,N_29451);
nor UO_1578 (O_1578,N_29341,N_29398);
nand UO_1579 (O_1579,N_29310,N_29981);
nand UO_1580 (O_1580,N_29638,N_28789);
xnor UO_1581 (O_1581,N_29485,N_29303);
and UO_1582 (O_1582,N_29089,N_29829);
and UO_1583 (O_1583,N_29153,N_29458);
nor UO_1584 (O_1584,N_29181,N_29658);
or UO_1585 (O_1585,N_29870,N_29705);
and UO_1586 (O_1586,N_29652,N_28505);
and UO_1587 (O_1587,N_29982,N_29119);
nor UO_1588 (O_1588,N_29535,N_29842);
nand UO_1589 (O_1589,N_29556,N_29835);
nand UO_1590 (O_1590,N_29986,N_29033);
and UO_1591 (O_1591,N_28518,N_28608);
nand UO_1592 (O_1592,N_29627,N_29690);
nand UO_1593 (O_1593,N_29110,N_28536);
and UO_1594 (O_1594,N_28528,N_29092);
xor UO_1595 (O_1595,N_29444,N_29574);
or UO_1596 (O_1596,N_28704,N_28834);
nor UO_1597 (O_1597,N_29185,N_29660);
and UO_1598 (O_1598,N_28603,N_28508);
xnor UO_1599 (O_1599,N_29137,N_29894);
and UO_1600 (O_1600,N_29637,N_29799);
xor UO_1601 (O_1601,N_29462,N_28966);
xor UO_1602 (O_1602,N_29251,N_29629);
and UO_1603 (O_1603,N_29605,N_28710);
or UO_1604 (O_1604,N_29260,N_28709);
nor UO_1605 (O_1605,N_29179,N_28789);
or UO_1606 (O_1606,N_29461,N_29861);
and UO_1607 (O_1607,N_29389,N_29315);
nand UO_1608 (O_1608,N_28704,N_29286);
and UO_1609 (O_1609,N_28954,N_29918);
or UO_1610 (O_1610,N_29460,N_29624);
nor UO_1611 (O_1611,N_29881,N_28785);
or UO_1612 (O_1612,N_28603,N_29937);
nor UO_1613 (O_1613,N_28609,N_28542);
and UO_1614 (O_1614,N_29373,N_29326);
nor UO_1615 (O_1615,N_29893,N_29506);
xor UO_1616 (O_1616,N_29797,N_29558);
and UO_1617 (O_1617,N_28542,N_28633);
nand UO_1618 (O_1618,N_29297,N_29025);
xor UO_1619 (O_1619,N_28937,N_29081);
nor UO_1620 (O_1620,N_28711,N_29043);
nor UO_1621 (O_1621,N_29566,N_28897);
nor UO_1622 (O_1622,N_29705,N_28542);
nand UO_1623 (O_1623,N_28570,N_28868);
or UO_1624 (O_1624,N_29955,N_29319);
nand UO_1625 (O_1625,N_28630,N_29628);
nand UO_1626 (O_1626,N_29846,N_29820);
nand UO_1627 (O_1627,N_29577,N_28520);
or UO_1628 (O_1628,N_29510,N_28630);
nor UO_1629 (O_1629,N_29555,N_29700);
nand UO_1630 (O_1630,N_29386,N_28923);
or UO_1631 (O_1631,N_28983,N_29004);
or UO_1632 (O_1632,N_29359,N_28919);
xor UO_1633 (O_1633,N_28622,N_29712);
and UO_1634 (O_1634,N_28865,N_29376);
xnor UO_1635 (O_1635,N_28509,N_28948);
nand UO_1636 (O_1636,N_29711,N_28635);
xor UO_1637 (O_1637,N_28966,N_29580);
nand UO_1638 (O_1638,N_29971,N_28774);
nand UO_1639 (O_1639,N_29552,N_28819);
xor UO_1640 (O_1640,N_28602,N_29545);
xor UO_1641 (O_1641,N_28785,N_29917);
nor UO_1642 (O_1642,N_29310,N_29836);
xor UO_1643 (O_1643,N_29002,N_29741);
nor UO_1644 (O_1644,N_28885,N_29627);
or UO_1645 (O_1645,N_28695,N_28946);
xor UO_1646 (O_1646,N_28804,N_28754);
xor UO_1647 (O_1647,N_29705,N_29193);
nand UO_1648 (O_1648,N_28709,N_28632);
xor UO_1649 (O_1649,N_29464,N_29248);
nand UO_1650 (O_1650,N_28671,N_29342);
xnor UO_1651 (O_1651,N_29350,N_28629);
and UO_1652 (O_1652,N_29248,N_28845);
nand UO_1653 (O_1653,N_29466,N_28964);
and UO_1654 (O_1654,N_29373,N_29250);
or UO_1655 (O_1655,N_28871,N_29535);
nand UO_1656 (O_1656,N_29192,N_29149);
xor UO_1657 (O_1657,N_28820,N_28832);
nor UO_1658 (O_1658,N_29391,N_29463);
nand UO_1659 (O_1659,N_29453,N_29451);
xor UO_1660 (O_1660,N_28592,N_28906);
nor UO_1661 (O_1661,N_29622,N_28834);
nor UO_1662 (O_1662,N_28977,N_29757);
xor UO_1663 (O_1663,N_29784,N_29030);
nand UO_1664 (O_1664,N_29407,N_28695);
nor UO_1665 (O_1665,N_29424,N_29641);
or UO_1666 (O_1666,N_29524,N_28523);
xnor UO_1667 (O_1667,N_29374,N_29432);
xor UO_1668 (O_1668,N_29470,N_28686);
or UO_1669 (O_1669,N_29429,N_29662);
xnor UO_1670 (O_1670,N_28922,N_29279);
and UO_1671 (O_1671,N_28546,N_29968);
or UO_1672 (O_1672,N_29334,N_29776);
nand UO_1673 (O_1673,N_29907,N_29687);
nor UO_1674 (O_1674,N_29694,N_28865);
nor UO_1675 (O_1675,N_28533,N_29076);
nor UO_1676 (O_1676,N_29236,N_29201);
nor UO_1677 (O_1677,N_28917,N_29402);
and UO_1678 (O_1678,N_28897,N_29754);
nor UO_1679 (O_1679,N_28932,N_29509);
nand UO_1680 (O_1680,N_29467,N_29713);
and UO_1681 (O_1681,N_28870,N_28895);
nor UO_1682 (O_1682,N_28822,N_28604);
or UO_1683 (O_1683,N_29237,N_29795);
xnor UO_1684 (O_1684,N_29250,N_29440);
nor UO_1685 (O_1685,N_29512,N_28945);
nand UO_1686 (O_1686,N_29589,N_29440);
and UO_1687 (O_1687,N_29866,N_29049);
or UO_1688 (O_1688,N_29900,N_29548);
nor UO_1689 (O_1689,N_29805,N_28689);
nand UO_1690 (O_1690,N_29275,N_29179);
nor UO_1691 (O_1691,N_28648,N_28596);
nor UO_1692 (O_1692,N_29514,N_29653);
nand UO_1693 (O_1693,N_29482,N_29466);
nor UO_1694 (O_1694,N_29982,N_28529);
or UO_1695 (O_1695,N_29378,N_29241);
nand UO_1696 (O_1696,N_29237,N_28780);
nand UO_1697 (O_1697,N_29154,N_29576);
and UO_1698 (O_1698,N_29926,N_28826);
or UO_1699 (O_1699,N_29679,N_29478);
xor UO_1700 (O_1700,N_29173,N_29406);
nor UO_1701 (O_1701,N_29075,N_29164);
and UO_1702 (O_1702,N_29052,N_29085);
or UO_1703 (O_1703,N_28989,N_29769);
nand UO_1704 (O_1704,N_28585,N_29545);
nand UO_1705 (O_1705,N_29203,N_29045);
xor UO_1706 (O_1706,N_29367,N_28866);
and UO_1707 (O_1707,N_29932,N_29238);
and UO_1708 (O_1708,N_29588,N_28718);
or UO_1709 (O_1709,N_28516,N_29089);
and UO_1710 (O_1710,N_29670,N_29271);
or UO_1711 (O_1711,N_29031,N_28682);
xor UO_1712 (O_1712,N_29183,N_29705);
nor UO_1713 (O_1713,N_29114,N_29292);
or UO_1714 (O_1714,N_29586,N_29954);
or UO_1715 (O_1715,N_29985,N_28964);
nor UO_1716 (O_1716,N_29710,N_29973);
and UO_1717 (O_1717,N_29707,N_29094);
xor UO_1718 (O_1718,N_28801,N_28765);
nand UO_1719 (O_1719,N_29711,N_29339);
or UO_1720 (O_1720,N_29302,N_28527);
and UO_1721 (O_1721,N_29887,N_28696);
and UO_1722 (O_1722,N_29941,N_29621);
and UO_1723 (O_1723,N_28942,N_29289);
nor UO_1724 (O_1724,N_29521,N_28822);
xnor UO_1725 (O_1725,N_29313,N_28826);
xnor UO_1726 (O_1726,N_28570,N_29060);
nor UO_1727 (O_1727,N_29623,N_28562);
xnor UO_1728 (O_1728,N_29592,N_28906);
and UO_1729 (O_1729,N_29449,N_29015);
or UO_1730 (O_1730,N_29371,N_28827);
xnor UO_1731 (O_1731,N_29429,N_29437);
or UO_1732 (O_1732,N_29142,N_29045);
xnor UO_1733 (O_1733,N_28552,N_29704);
nand UO_1734 (O_1734,N_29862,N_29005);
or UO_1735 (O_1735,N_28782,N_29476);
nor UO_1736 (O_1736,N_29018,N_29146);
and UO_1737 (O_1737,N_28821,N_29386);
nand UO_1738 (O_1738,N_28870,N_29837);
xnor UO_1739 (O_1739,N_28946,N_29369);
nor UO_1740 (O_1740,N_29637,N_29034);
nand UO_1741 (O_1741,N_29570,N_29064);
and UO_1742 (O_1742,N_29300,N_28558);
nor UO_1743 (O_1743,N_28570,N_28907);
or UO_1744 (O_1744,N_29776,N_29647);
or UO_1745 (O_1745,N_29694,N_29212);
nor UO_1746 (O_1746,N_29338,N_29066);
nand UO_1747 (O_1747,N_28834,N_28674);
xor UO_1748 (O_1748,N_28556,N_29039);
and UO_1749 (O_1749,N_29053,N_28995);
nor UO_1750 (O_1750,N_29631,N_28581);
and UO_1751 (O_1751,N_29507,N_28693);
xor UO_1752 (O_1752,N_29820,N_29187);
xor UO_1753 (O_1753,N_29562,N_29846);
xor UO_1754 (O_1754,N_28877,N_29067);
nand UO_1755 (O_1755,N_29412,N_29100);
and UO_1756 (O_1756,N_29988,N_29657);
nor UO_1757 (O_1757,N_29436,N_28811);
nand UO_1758 (O_1758,N_29359,N_28848);
and UO_1759 (O_1759,N_28950,N_29591);
nor UO_1760 (O_1760,N_28995,N_29729);
xor UO_1761 (O_1761,N_29431,N_28940);
or UO_1762 (O_1762,N_29534,N_28887);
or UO_1763 (O_1763,N_29104,N_29596);
nor UO_1764 (O_1764,N_28653,N_29741);
xnor UO_1765 (O_1765,N_28636,N_28651);
nand UO_1766 (O_1766,N_29359,N_29007);
and UO_1767 (O_1767,N_29479,N_29995);
nor UO_1768 (O_1768,N_29557,N_28672);
and UO_1769 (O_1769,N_29582,N_28957);
nand UO_1770 (O_1770,N_29991,N_28923);
and UO_1771 (O_1771,N_29088,N_29404);
nand UO_1772 (O_1772,N_29862,N_29971);
nand UO_1773 (O_1773,N_29356,N_28629);
or UO_1774 (O_1774,N_28826,N_29178);
and UO_1775 (O_1775,N_29166,N_29822);
nand UO_1776 (O_1776,N_28633,N_29183);
nand UO_1777 (O_1777,N_29046,N_29322);
xor UO_1778 (O_1778,N_29863,N_29859);
and UO_1779 (O_1779,N_29897,N_28569);
or UO_1780 (O_1780,N_29404,N_28897);
and UO_1781 (O_1781,N_29810,N_29395);
xnor UO_1782 (O_1782,N_29054,N_29985);
or UO_1783 (O_1783,N_29348,N_29922);
xor UO_1784 (O_1784,N_28605,N_29202);
nor UO_1785 (O_1785,N_29029,N_29527);
or UO_1786 (O_1786,N_29231,N_29027);
xnor UO_1787 (O_1787,N_29311,N_29548);
and UO_1788 (O_1788,N_29820,N_28803);
nand UO_1789 (O_1789,N_28886,N_29013);
and UO_1790 (O_1790,N_29308,N_28954);
xnor UO_1791 (O_1791,N_28924,N_29615);
xor UO_1792 (O_1792,N_28781,N_29320);
or UO_1793 (O_1793,N_29106,N_29627);
and UO_1794 (O_1794,N_29260,N_28982);
and UO_1795 (O_1795,N_29867,N_29225);
and UO_1796 (O_1796,N_29316,N_29495);
xnor UO_1797 (O_1797,N_28848,N_29548);
nand UO_1798 (O_1798,N_29247,N_28632);
and UO_1799 (O_1799,N_28524,N_29216);
or UO_1800 (O_1800,N_29408,N_28547);
xnor UO_1801 (O_1801,N_28735,N_28894);
xor UO_1802 (O_1802,N_29255,N_28720);
nor UO_1803 (O_1803,N_29852,N_29768);
and UO_1804 (O_1804,N_28567,N_28568);
nor UO_1805 (O_1805,N_29878,N_29925);
nor UO_1806 (O_1806,N_28930,N_29456);
nand UO_1807 (O_1807,N_28968,N_29541);
nand UO_1808 (O_1808,N_29783,N_29696);
xnor UO_1809 (O_1809,N_28723,N_28907);
and UO_1810 (O_1810,N_29881,N_29566);
and UO_1811 (O_1811,N_29577,N_29069);
xnor UO_1812 (O_1812,N_29978,N_29747);
nand UO_1813 (O_1813,N_28566,N_29973);
xor UO_1814 (O_1814,N_29886,N_28579);
nand UO_1815 (O_1815,N_29426,N_28523);
and UO_1816 (O_1816,N_29179,N_29292);
nor UO_1817 (O_1817,N_28590,N_28508);
nand UO_1818 (O_1818,N_29372,N_29877);
or UO_1819 (O_1819,N_28755,N_28688);
or UO_1820 (O_1820,N_29188,N_29930);
or UO_1821 (O_1821,N_29413,N_29133);
or UO_1822 (O_1822,N_29824,N_29439);
nand UO_1823 (O_1823,N_28606,N_29128);
xnor UO_1824 (O_1824,N_28628,N_28844);
xor UO_1825 (O_1825,N_29830,N_28661);
xnor UO_1826 (O_1826,N_29810,N_29411);
and UO_1827 (O_1827,N_29551,N_28796);
nand UO_1828 (O_1828,N_28945,N_29573);
nand UO_1829 (O_1829,N_28815,N_29764);
nand UO_1830 (O_1830,N_28649,N_28843);
nor UO_1831 (O_1831,N_28645,N_29828);
or UO_1832 (O_1832,N_29307,N_29099);
or UO_1833 (O_1833,N_29800,N_28578);
xor UO_1834 (O_1834,N_29381,N_28812);
and UO_1835 (O_1835,N_29301,N_28924);
and UO_1836 (O_1836,N_29615,N_28776);
nor UO_1837 (O_1837,N_29901,N_29028);
nand UO_1838 (O_1838,N_28951,N_29777);
or UO_1839 (O_1839,N_29601,N_28661);
nor UO_1840 (O_1840,N_29290,N_29205);
nand UO_1841 (O_1841,N_29064,N_29769);
and UO_1842 (O_1842,N_29132,N_28846);
and UO_1843 (O_1843,N_29824,N_28970);
and UO_1844 (O_1844,N_28681,N_29127);
nor UO_1845 (O_1845,N_29142,N_29930);
nand UO_1846 (O_1846,N_28672,N_29848);
nand UO_1847 (O_1847,N_29740,N_29154);
nor UO_1848 (O_1848,N_29540,N_29817);
nor UO_1849 (O_1849,N_29437,N_29038);
xor UO_1850 (O_1850,N_29648,N_29008);
xor UO_1851 (O_1851,N_29709,N_29459);
nand UO_1852 (O_1852,N_29983,N_29399);
or UO_1853 (O_1853,N_29864,N_29376);
nor UO_1854 (O_1854,N_28626,N_29488);
and UO_1855 (O_1855,N_28703,N_29295);
or UO_1856 (O_1856,N_28858,N_28845);
or UO_1857 (O_1857,N_28707,N_29067);
xor UO_1858 (O_1858,N_28957,N_29133);
nand UO_1859 (O_1859,N_29213,N_29180);
nand UO_1860 (O_1860,N_28969,N_29005);
or UO_1861 (O_1861,N_29107,N_29370);
nor UO_1862 (O_1862,N_29420,N_29019);
nor UO_1863 (O_1863,N_29686,N_28622);
nand UO_1864 (O_1864,N_29932,N_28729);
and UO_1865 (O_1865,N_29160,N_29346);
nand UO_1866 (O_1866,N_29156,N_29600);
or UO_1867 (O_1867,N_28691,N_29925);
nor UO_1868 (O_1868,N_29610,N_29717);
and UO_1869 (O_1869,N_28813,N_29593);
or UO_1870 (O_1870,N_29940,N_28751);
or UO_1871 (O_1871,N_28627,N_29587);
xnor UO_1872 (O_1872,N_29154,N_29803);
nand UO_1873 (O_1873,N_29512,N_29442);
xnor UO_1874 (O_1874,N_28644,N_29811);
nand UO_1875 (O_1875,N_29645,N_29963);
nand UO_1876 (O_1876,N_28542,N_29819);
or UO_1877 (O_1877,N_29542,N_28816);
nand UO_1878 (O_1878,N_29392,N_29876);
nor UO_1879 (O_1879,N_28618,N_29909);
and UO_1880 (O_1880,N_28836,N_29895);
xnor UO_1881 (O_1881,N_29327,N_29194);
nand UO_1882 (O_1882,N_28853,N_28740);
nand UO_1883 (O_1883,N_29025,N_29222);
xor UO_1884 (O_1884,N_29337,N_28917);
nor UO_1885 (O_1885,N_29499,N_29573);
and UO_1886 (O_1886,N_29015,N_29827);
and UO_1887 (O_1887,N_29461,N_29271);
xnor UO_1888 (O_1888,N_29245,N_28974);
nor UO_1889 (O_1889,N_29869,N_29698);
or UO_1890 (O_1890,N_29163,N_29927);
or UO_1891 (O_1891,N_28914,N_29764);
nand UO_1892 (O_1892,N_28899,N_29790);
or UO_1893 (O_1893,N_29778,N_29655);
xor UO_1894 (O_1894,N_29214,N_29708);
or UO_1895 (O_1895,N_28589,N_28587);
nor UO_1896 (O_1896,N_29044,N_29198);
xor UO_1897 (O_1897,N_29465,N_29802);
xor UO_1898 (O_1898,N_29503,N_28781);
nand UO_1899 (O_1899,N_29496,N_29630);
or UO_1900 (O_1900,N_29866,N_28699);
and UO_1901 (O_1901,N_29435,N_29483);
xor UO_1902 (O_1902,N_28541,N_28754);
nor UO_1903 (O_1903,N_29500,N_29039);
nor UO_1904 (O_1904,N_28743,N_29648);
or UO_1905 (O_1905,N_28847,N_29898);
nor UO_1906 (O_1906,N_28637,N_29399);
or UO_1907 (O_1907,N_28504,N_28759);
or UO_1908 (O_1908,N_29761,N_29780);
and UO_1909 (O_1909,N_29177,N_29333);
xor UO_1910 (O_1910,N_28909,N_29372);
nor UO_1911 (O_1911,N_28612,N_29371);
and UO_1912 (O_1912,N_29689,N_28650);
and UO_1913 (O_1913,N_29409,N_29173);
or UO_1914 (O_1914,N_29492,N_28534);
or UO_1915 (O_1915,N_29426,N_28689);
or UO_1916 (O_1916,N_28634,N_29948);
nor UO_1917 (O_1917,N_28874,N_29189);
xnor UO_1918 (O_1918,N_29487,N_29446);
nand UO_1919 (O_1919,N_28643,N_29497);
nor UO_1920 (O_1920,N_29256,N_29622);
nor UO_1921 (O_1921,N_29040,N_29568);
nand UO_1922 (O_1922,N_29918,N_29235);
or UO_1923 (O_1923,N_29802,N_29463);
or UO_1924 (O_1924,N_28628,N_28874);
nand UO_1925 (O_1925,N_29263,N_28727);
nor UO_1926 (O_1926,N_29792,N_29597);
and UO_1927 (O_1927,N_29799,N_29554);
xnor UO_1928 (O_1928,N_29441,N_29152);
nor UO_1929 (O_1929,N_29178,N_29335);
nand UO_1930 (O_1930,N_29712,N_29858);
nand UO_1931 (O_1931,N_28617,N_29214);
xnor UO_1932 (O_1932,N_29874,N_29551);
nand UO_1933 (O_1933,N_29066,N_29362);
nor UO_1934 (O_1934,N_29664,N_29243);
and UO_1935 (O_1935,N_28572,N_29068);
xor UO_1936 (O_1936,N_29570,N_29458);
xor UO_1937 (O_1937,N_29571,N_29272);
nor UO_1938 (O_1938,N_29671,N_28656);
and UO_1939 (O_1939,N_28902,N_28711);
or UO_1940 (O_1940,N_29578,N_28955);
or UO_1941 (O_1941,N_29957,N_29331);
and UO_1942 (O_1942,N_28547,N_28667);
xor UO_1943 (O_1943,N_29465,N_28993);
nand UO_1944 (O_1944,N_29273,N_29345);
nand UO_1945 (O_1945,N_29166,N_29057);
and UO_1946 (O_1946,N_29205,N_29055);
xor UO_1947 (O_1947,N_28664,N_29962);
nand UO_1948 (O_1948,N_29147,N_28967);
nand UO_1949 (O_1949,N_28787,N_29307);
nand UO_1950 (O_1950,N_29635,N_29868);
nand UO_1951 (O_1951,N_29715,N_29684);
nor UO_1952 (O_1952,N_29055,N_29211);
xnor UO_1953 (O_1953,N_29068,N_28837);
and UO_1954 (O_1954,N_29856,N_28851);
nor UO_1955 (O_1955,N_29800,N_29658);
and UO_1956 (O_1956,N_29459,N_29525);
xnor UO_1957 (O_1957,N_29659,N_28741);
or UO_1958 (O_1958,N_29903,N_29595);
or UO_1959 (O_1959,N_29112,N_29561);
nand UO_1960 (O_1960,N_29116,N_29676);
nand UO_1961 (O_1961,N_28801,N_28548);
and UO_1962 (O_1962,N_28944,N_28954);
nor UO_1963 (O_1963,N_28583,N_28859);
xnor UO_1964 (O_1964,N_28826,N_28887);
nor UO_1965 (O_1965,N_28501,N_28740);
and UO_1966 (O_1966,N_28826,N_29577);
and UO_1967 (O_1967,N_28526,N_29061);
xnor UO_1968 (O_1968,N_29478,N_29917);
and UO_1969 (O_1969,N_29180,N_29116);
nor UO_1970 (O_1970,N_29770,N_28844);
xor UO_1971 (O_1971,N_29525,N_29219);
nand UO_1972 (O_1972,N_28932,N_28755);
nor UO_1973 (O_1973,N_28708,N_29257);
xnor UO_1974 (O_1974,N_29615,N_29166);
and UO_1975 (O_1975,N_29462,N_29179);
or UO_1976 (O_1976,N_29015,N_29555);
nor UO_1977 (O_1977,N_29722,N_29285);
xnor UO_1978 (O_1978,N_28951,N_29977);
nand UO_1979 (O_1979,N_28625,N_28784);
and UO_1980 (O_1980,N_29636,N_29403);
or UO_1981 (O_1981,N_29493,N_28655);
or UO_1982 (O_1982,N_28828,N_29171);
nor UO_1983 (O_1983,N_28544,N_28953);
nand UO_1984 (O_1984,N_29091,N_29426);
nor UO_1985 (O_1985,N_29478,N_29687);
nand UO_1986 (O_1986,N_29611,N_29208);
or UO_1987 (O_1987,N_29125,N_29814);
and UO_1988 (O_1988,N_29403,N_29418);
nand UO_1989 (O_1989,N_29587,N_28897);
nor UO_1990 (O_1990,N_29786,N_28645);
nor UO_1991 (O_1991,N_28943,N_29145);
and UO_1992 (O_1992,N_29712,N_29232);
or UO_1993 (O_1993,N_28576,N_29403);
nor UO_1994 (O_1994,N_29400,N_29550);
nor UO_1995 (O_1995,N_29005,N_29577);
nor UO_1996 (O_1996,N_29843,N_29459);
xnor UO_1997 (O_1997,N_28610,N_29886);
nor UO_1998 (O_1998,N_29836,N_28852);
xnor UO_1999 (O_1999,N_29379,N_28728);
nor UO_2000 (O_2000,N_29425,N_28845);
nor UO_2001 (O_2001,N_29922,N_28545);
or UO_2002 (O_2002,N_29123,N_29775);
nor UO_2003 (O_2003,N_29158,N_29112);
nor UO_2004 (O_2004,N_28744,N_29621);
and UO_2005 (O_2005,N_28936,N_29404);
and UO_2006 (O_2006,N_28744,N_29704);
and UO_2007 (O_2007,N_29577,N_28848);
nor UO_2008 (O_2008,N_29701,N_29828);
and UO_2009 (O_2009,N_28861,N_29977);
xnor UO_2010 (O_2010,N_28873,N_29080);
nor UO_2011 (O_2011,N_29743,N_29031);
nand UO_2012 (O_2012,N_29037,N_29877);
nor UO_2013 (O_2013,N_29953,N_29628);
or UO_2014 (O_2014,N_29653,N_29447);
nor UO_2015 (O_2015,N_29138,N_29816);
nand UO_2016 (O_2016,N_29740,N_28860);
and UO_2017 (O_2017,N_29554,N_29671);
nand UO_2018 (O_2018,N_28500,N_28703);
xnor UO_2019 (O_2019,N_29023,N_28674);
xor UO_2020 (O_2020,N_28530,N_29227);
or UO_2021 (O_2021,N_29921,N_28773);
nand UO_2022 (O_2022,N_29527,N_28516);
and UO_2023 (O_2023,N_29665,N_29742);
or UO_2024 (O_2024,N_29572,N_29779);
and UO_2025 (O_2025,N_29644,N_29838);
nor UO_2026 (O_2026,N_28974,N_29173);
xor UO_2027 (O_2027,N_28887,N_29849);
or UO_2028 (O_2028,N_28751,N_28671);
or UO_2029 (O_2029,N_29130,N_28633);
nor UO_2030 (O_2030,N_29645,N_28609);
and UO_2031 (O_2031,N_28922,N_28831);
and UO_2032 (O_2032,N_29620,N_29188);
and UO_2033 (O_2033,N_29450,N_28642);
and UO_2034 (O_2034,N_29745,N_28734);
xnor UO_2035 (O_2035,N_29107,N_28600);
or UO_2036 (O_2036,N_28757,N_29647);
xor UO_2037 (O_2037,N_28996,N_29720);
xnor UO_2038 (O_2038,N_28989,N_28560);
xor UO_2039 (O_2039,N_29634,N_28616);
xor UO_2040 (O_2040,N_29433,N_29976);
or UO_2041 (O_2041,N_29411,N_28617);
or UO_2042 (O_2042,N_29150,N_28982);
xnor UO_2043 (O_2043,N_28561,N_29197);
nor UO_2044 (O_2044,N_28629,N_28582);
nor UO_2045 (O_2045,N_29637,N_28596);
xor UO_2046 (O_2046,N_29468,N_28723);
nand UO_2047 (O_2047,N_28855,N_29189);
xnor UO_2048 (O_2048,N_28824,N_29596);
and UO_2049 (O_2049,N_28913,N_29283);
xnor UO_2050 (O_2050,N_29273,N_28528);
or UO_2051 (O_2051,N_29250,N_29986);
and UO_2052 (O_2052,N_29393,N_28959);
or UO_2053 (O_2053,N_28628,N_28655);
nor UO_2054 (O_2054,N_29336,N_29230);
or UO_2055 (O_2055,N_29034,N_29642);
nor UO_2056 (O_2056,N_29793,N_28641);
nand UO_2057 (O_2057,N_28614,N_29392);
xnor UO_2058 (O_2058,N_28714,N_29161);
nand UO_2059 (O_2059,N_29534,N_29831);
xnor UO_2060 (O_2060,N_29743,N_29253);
xnor UO_2061 (O_2061,N_28591,N_29284);
or UO_2062 (O_2062,N_28587,N_29545);
or UO_2063 (O_2063,N_28554,N_28583);
nand UO_2064 (O_2064,N_28898,N_29147);
xnor UO_2065 (O_2065,N_29415,N_29297);
nand UO_2066 (O_2066,N_28788,N_29993);
nand UO_2067 (O_2067,N_29650,N_28503);
or UO_2068 (O_2068,N_29341,N_29215);
or UO_2069 (O_2069,N_29259,N_29069);
nor UO_2070 (O_2070,N_29703,N_28625);
nor UO_2071 (O_2071,N_28540,N_29659);
nand UO_2072 (O_2072,N_29933,N_29342);
nor UO_2073 (O_2073,N_29582,N_29337);
or UO_2074 (O_2074,N_29930,N_28858);
nor UO_2075 (O_2075,N_29673,N_29094);
nand UO_2076 (O_2076,N_29351,N_28571);
nand UO_2077 (O_2077,N_28764,N_28736);
or UO_2078 (O_2078,N_29072,N_29682);
or UO_2079 (O_2079,N_29641,N_28633);
and UO_2080 (O_2080,N_29287,N_29895);
xor UO_2081 (O_2081,N_29739,N_29781);
xnor UO_2082 (O_2082,N_28850,N_28949);
and UO_2083 (O_2083,N_29334,N_28524);
and UO_2084 (O_2084,N_28834,N_28600);
nand UO_2085 (O_2085,N_29322,N_29794);
xnor UO_2086 (O_2086,N_29380,N_28967);
nand UO_2087 (O_2087,N_28851,N_29710);
and UO_2088 (O_2088,N_29550,N_28539);
and UO_2089 (O_2089,N_29376,N_29385);
xnor UO_2090 (O_2090,N_29860,N_28671);
nor UO_2091 (O_2091,N_28826,N_29000);
xor UO_2092 (O_2092,N_29682,N_29988);
xor UO_2093 (O_2093,N_29042,N_28906);
or UO_2094 (O_2094,N_28706,N_28612);
nand UO_2095 (O_2095,N_28981,N_29763);
nand UO_2096 (O_2096,N_29890,N_29213);
xnor UO_2097 (O_2097,N_28637,N_29574);
nand UO_2098 (O_2098,N_29795,N_28556);
xnor UO_2099 (O_2099,N_28901,N_28586);
xor UO_2100 (O_2100,N_29964,N_29312);
and UO_2101 (O_2101,N_29673,N_29529);
nor UO_2102 (O_2102,N_29096,N_28594);
and UO_2103 (O_2103,N_28678,N_29079);
or UO_2104 (O_2104,N_29128,N_29717);
nand UO_2105 (O_2105,N_29649,N_29976);
xor UO_2106 (O_2106,N_28763,N_28680);
nand UO_2107 (O_2107,N_28671,N_29185);
and UO_2108 (O_2108,N_29669,N_29377);
nor UO_2109 (O_2109,N_29951,N_29027);
nand UO_2110 (O_2110,N_28596,N_29353);
or UO_2111 (O_2111,N_29064,N_29001);
or UO_2112 (O_2112,N_28799,N_29006);
nand UO_2113 (O_2113,N_29980,N_29807);
or UO_2114 (O_2114,N_29406,N_28597);
nand UO_2115 (O_2115,N_28636,N_29965);
or UO_2116 (O_2116,N_29471,N_28954);
nor UO_2117 (O_2117,N_29415,N_28611);
xnor UO_2118 (O_2118,N_29854,N_29814);
or UO_2119 (O_2119,N_29073,N_29266);
or UO_2120 (O_2120,N_28602,N_29030);
nor UO_2121 (O_2121,N_28745,N_29206);
nand UO_2122 (O_2122,N_28918,N_29014);
and UO_2123 (O_2123,N_28587,N_28763);
or UO_2124 (O_2124,N_29914,N_28503);
nand UO_2125 (O_2125,N_29837,N_28699);
xnor UO_2126 (O_2126,N_28956,N_29797);
xnor UO_2127 (O_2127,N_28752,N_28603);
and UO_2128 (O_2128,N_28597,N_28770);
xor UO_2129 (O_2129,N_29196,N_29556);
and UO_2130 (O_2130,N_28812,N_28556);
and UO_2131 (O_2131,N_28809,N_29882);
and UO_2132 (O_2132,N_29070,N_29925);
or UO_2133 (O_2133,N_28785,N_29507);
and UO_2134 (O_2134,N_29423,N_29801);
xor UO_2135 (O_2135,N_28603,N_28601);
nor UO_2136 (O_2136,N_29064,N_28840);
nand UO_2137 (O_2137,N_29435,N_29604);
and UO_2138 (O_2138,N_28974,N_29504);
xor UO_2139 (O_2139,N_28634,N_29771);
nand UO_2140 (O_2140,N_29083,N_29200);
nor UO_2141 (O_2141,N_28788,N_29870);
xor UO_2142 (O_2142,N_29836,N_29933);
or UO_2143 (O_2143,N_29839,N_28813);
and UO_2144 (O_2144,N_29598,N_29146);
and UO_2145 (O_2145,N_29561,N_28707);
or UO_2146 (O_2146,N_29962,N_29767);
xor UO_2147 (O_2147,N_28873,N_28755);
xnor UO_2148 (O_2148,N_28584,N_29000);
or UO_2149 (O_2149,N_29283,N_29017);
nor UO_2150 (O_2150,N_29803,N_29719);
and UO_2151 (O_2151,N_29565,N_28720);
and UO_2152 (O_2152,N_28676,N_29529);
nand UO_2153 (O_2153,N_28975,N_29236);
nand UO_2154 (O_2154,N_29399,N_28955);
nand UO_2155 (O_2155,N_29728,N_29482);
nand UO_2156 (O_2156,N_28891,N_29480);
nor UO_2157 (O_2157,N_28899,N_29104);
and UO_2158 (O_2158,N_29194,N_29838);
nand UO_2159 (O_2159,N_29619,N_28723);
xor UO_2160 (O_2160,N_29180,N_29795);
and UO_2161 (O_2161,N_28965,N_29052);
nor UO_2162 (O_2162,N_28863,N_29786);
or UO_2163 (O_2163,N_28615,N_29390);
or UO_2164 (O_2164,N_29612,N_29894);
or UO_2165 (O_2165,N_29813,N_29165);
and UO_2166 (O_2166,N_29538,N_29220);
xnor UO_2167 (O_2167,N_29773,N_29378);
nand UO_2168 (O_2168,N_29663,N_29112);
or UO_2169 (O_2169,N_29655,N_29509);
nand UO_2170 (O_2170,N_28736,N_29640);
or UO_2171 (O_2171,N_28665,N_28727);
or UO_2172 (O_2172,N_28920,N_28929);
or UO_2173 (O_2173,N_29972,N_28551);
nand UO_2174 (O_2174,N_29551,N_29222);
or UO_2175 (O_2175,N_28829,N_29134);
and UO_2176 (O_2176,N_29231,N_29220);
or UO_2177 (O_2177,N_29413,N_28734);
and UO_2178 (O_2178,N_29585,N_29535);
nand UO_2179 (O_2179,N_29898,N_29262);
nand UO_2180 (O_2180,N_29067,N_28746);
and UO_2181 (O_2181,N_29122,N_29697);
nor UO_2182 (O_2182,N_29525,N_29535);
nand UO_2183 (O_2183,N_29041,N_28975);
xnor UO_2184 (O_2184,N_29375,N_28775);
or UO_2185 (O_2185,N_29553,N_29969);
xnor UO_2186 (O_2186,N_29970,N_28572);
or UO_2187 (O_2187,N_29116,N_28923);
xnor UO_2188 (O_2188,N_29014,N_28746);
xor UO_2189 (O_2189,N_28867,N_28691);
nor UO_2190 (O_2190,N_29518,N_29413);
nand UO_2191 (O_2191,N_29145,N_29795);
nor UO_2192 (O_2192,N_29679,N_28761);
and UO_2193 (O_2193,N_29522,N_29264);
nand UO_2194 (O_2194,N_29932,N_29839);
and UO_2195 (O_2195,N_29124,N_28781);
xnor UO_2196 (O_2196,N_28771,N_29096);
and UO_2197 (O_2197,N_29080,N_28692);
and UO_2198 (O_2198,N_28902,N_29655);
or UO_2199 (O_2199,N_28739,N_29901);
or UO_2200 (O_2200,N_29869,N_29907);
and UO_2201 (O_2201,N_29491,N_29474);
nor UO_2202 (O_2202,N_29199,N_29692);
nand UO_2203 (O_2203,N_28908,N_29256);
and UO_2204 (O_2204,N_29547,N_29318);
and UO_2205 (O_2205,N_29880,N_29186);
or UO_2206 (O_2206,N_29795,N_29061);
or UO_2207 (O_2207,N_29084,N_29515);
or UO_2208 (O_2208,N_29938,N_29341);
and UO_2209 (O_2209,N_29290,N_29675);
nand UO_2210 (O_2210,N_29324,N_29039);
or UO_2211 (O_2211,N_29064,N_28622);
and UO_2212 (O_2212,N_29913,N_29358);
or UO_2213 (O_2213,N_28784,N_28551);
and UO_2214 (O_2214,N_28911,N_29622);
or UO_2215 (O_2215,N_29844,N_28827);
or UO_2216 (O_2216,N_28994,N_29898);
xnor UO_2217 (O_2217,N_28961,N_29426);
xor UO_2218 (O_2218,N_29621,N_29377);
and UO_2219 (O_2219,N_28914,N_28975);
nand UO_2220 (O_2220,N_29100,N_29617);
nand UO_2221 (O_2221,N_29721,N_29252);
or UO_2222 (O_2222,N_29622,N_28866);
nor UO_2223 (O_2223,N_28966,N_29825);
xnor UO_2224 (O_2224,N_29357,N_28999);
nand UO_2225 (O_2225,N_28930,N_28518);
or UO_2226 (O_2226,N_28554,N_29426);
nand UO_2227 (O_2227,N_28535,N_28657);
nand UO_2228 (O_2228,N_28659,N_29286);
or UO_2229 (O_2229,N_28732,N_28730);
nand UO_2230 (O_2230,N_28843,N_29493);
nor UO_2231 (O_2231,N_29608,N_29037);
xnor UO_2232 (O_2232,N_29395,N_29341);
nand UO_2233 (O_2233,N_29681,N_29844);
or UO_2234 (O_2234,N_28584,N_28981);
xnor UO_2235 (O_2235,N_28676,N_29659);
xor UO_2236 (O_2236,N_29329,N_29030);
or UO_2237 (O_2237,N_29126,N_29206);
and UO_2238 (O_2238,N_28999,N_29321);
xnor UO_2239 (O_2239,N_29869,N_29050);
xnor UO_2240 (O_2240,N_29119,N_29654);
nand UO_2241 (O_2241,N_28500,N_29790);
nor UO_2242 (O_2242,N_29123,N_29797);
nand UO_2243 (O_2243,N_29788,N_28663);
nand UO_2244 (O_2244,N_28690,N_29891);
or UO_2245 (O_2245,N_28788,N_28701);
xnor UO_2246 (O_2246,N_28881,N_29451);
xor UO_2247 (O_2247,N_28752,N_29262);
or UO_2248 (O_2248,N_29937,N_29493);
or UO_2249 (O_2249,N_29664,N_28540);
nor UO_2250 (O_2250,N_29497,N_28929);
nand UO_2251 (O_2251,N_29548,N_29061);
nor UO_2252 (O_2252,N_28755,N_29772);
xor UO_2253 (O_2253,N_29240,N_29889);
nand UO_2254 (O_2254,N_29999,N_28568);
nor UO_2255 (O_2255,N_29072,N_28846);
xnor UO_2256 (O_2256,N_29824,N_29683);
nand UO_2257 (O_2257,N_28549,N_29602);
nand UO_2258 (O_2258,N_29753,N_29130);
nand UO_2259 (O_2259,N_29198,N_28761);
or UO_2260 (O_2260,N_29395,N_29452);
or UO_2261 (O_2261,N_29873,N_29173);
and UO_2262 (O_2262,N_29013,N_29919);
or UO_2263 (O_2263,N_28851,N_29564);
nand UO_2264 (O_2264,N_29219,N_29289);
xnor UO_2265 (O_2265,N_28778,N_29285);
or UO_2266 (O_2266,N_28850,N_29799);
or UO_2267 (O_2267,N_28736,N_29842);
or UO_2268 (O_2268,N_29155,N_28902);
nand UO_2269 (O_2269,N_28738,N_29705);
nor UO_2270 (O_2270,N_29277,N_28986);
or UO_2271 (O_2271,N_29156,N_29097);
xor UO_2272 (O_2272,N_29157,N_28875);
or UO_2273 (O_2273,N_29011,N_28574);
xnor UO_2274 (O_2274,N_29460,N_29362);
and UO_2275 (O_2275,N_29506,N_29866);
and UO_2276 (O_2276,N_29618,N_29262);
nand UO_2277 (O_2277,N_29005,N_29526);
nand UO_2278 (O_2278,N_28532,N_29596);
and UO_2279 (O_2279,N_29840,N_29649);
xor UO_2280 (O_2280,N_29745,N_29723);
nand UO_2281 (O_2281,N_28862,N_29535);
and UO_2282 (O_2282,N_28808,N_29867);
nand UO_2283 (O_2283,N_29074,N_29101);
and UO_2284 (O_2284,N_29632,N_29040);
nand UO_2285 (O_2285,N_28725,N_29998);
nand UO_2286 (O_2286,N_28757,N_29825);
or UO_2287 (O_2287,N_29065,N_29721);
nand UO_2288 (O_2288,N_29260,N_29557);
nor UO_2289 (O_2289,N_28784,N_29348);
and UO_2290 (O_2290,N_29907,N_29473);
nor UO_2291 (O_2291,N_29771,N_28818);
and UO_2292 (O_2292,N_28619,N_29032);
xnor UO_2293 (O_2293,N_28778,N_28893);
nand UO_2294 (O_2294,N_28553,N_28591);
or UO_2295 (O_2295,N_28787,N_28635);
nand UO_2296 (O_2296,N_29187,N_29890);
xnor UO_2297 (O_2297,N_29049,N_29686);
nor UO_2298 (O_2298,N_29315,N_28974);
nand UO_2299 (O_2299,N_28634,N_29979);
xnor UO_2300 (O_2300,N_28603,N_29892);
and UO_2301 (O_2301,N_28733,N_29053);
xnor UO_2302 (O_2302,N_28539,N_29668);
or UO_2303 (O_2303,N_28952,N_29152);
nor UO_2304 (O_2304,N_29778,N_29405);
nand UO_2305 (O_2305,N_29140,N_29283);
nand UO_2306 (O_2306,N_29841,N_29381);
or UO_2307 (O_2307,N_28799,N_29488);
and UO_2308 (O_2308,N_29879,N_28636);
nand UO_2309 (O_2309,N_28658,N_29293);
nand UO_2310 (O_2310,N_29113,N_28984);
and UO_2311 (O_2311,N_29717,N_29017);
or UO_2312 (O_2312,N_29063,N_29641);
or UO_2313 (O_2313,N_29747,N_28665);
or UO_2314 (O_2314,N_29621,N_29630);
nand UO_2315 (O_2315,N_28529,N_29559);
nand UO_2316 (O_2316,N_28531,N_29106);
and UO_2317 (O_2317,N_28964,N_29153);
xnor UO_2318 (O_2318,N_28579,N_28633);
nand UO_2319 (O_2319,N_28525,N_29150);
nor UO_2320 (O_2320,N_29159,N_29999);
nand UO_2321 (O_2321,N_29689,N_28693);
or UO_2322 (O_2322,N_29049,N_28899);
nor UO_2323 (O_2323,N_29127,N_29755);
nand UO_2324 (O_2324,N_29769,N_29170);
nor UO_2325 (O_2325,N_28891,N_28673);
and UO_2326 (O_2326,N_29405,N_29458);
nand UO_2327 (O_2327,N_28507,N_28661);
xnor UO_2328 (O_2328,N_29962,N_29186);
and UO_2329 (O_2329,N_29613,N_29052);
nor UO_2330 (O_2330,N_29180,N_28888);
and UO_2331 (O_2331,N_29199,N_29095);
nand UO_2332 (O_2332,N_29408,N_29761);
or UO_2333 (O_2333,N_28575,N_29495);
nand UO_2334 (O_2334,N_29087,N_28807);
or UO_2335 (O_2335,N_29737,N_29282);
or UO_2336 (O_2336,N_29969,N_28943);
or UO_2337 (O_2337,N_29358,N_28777);
nand UO_2338 (O_2338,N_29537,N_28891);
nand UO_2339 (O_2339,N_29857,N_28752);
nand UO_2340 (O_2340,N_29683,N_28607);
xor UO_2341 (O_2341,N_29090,N_29066);
nor UO_2342 (O_2342,N_29990,N_29276);
and UO_2343 (O_2343,N_29397,N_29426);
nor UO_2344 (O_2344,N_29890,N_29957);
xor UO_2345 (O_2345,N_28737,N_28674);
and UO_2346 (O_2346,N_28628,N_29187);
and UO_2347 (O_2347,N_29065,N_29368);
xnor UO_2348 (O_2348,N_29615,N_28919);
and UO_2349 (O_2349,N_29303,N_29635);
or UO_2350 (O_2350,N_29732,N_29130);
xnor UO_2351 (O_2351,N_29883,N_29820);
nor UO_2352 (O_2352,N_28987,N_29094);
or UO_2353 (O_2353,N_29939,N_29535);
nand UO_2354 (O_2354,N_29607,N_29448);
nand UO_2355 (O_2355,N_29577,N_29839);
xnor UO_2356 (O_2356,N_28968,N_29939);
xnor UO_2357 (O_2357,N_28725,N_28840);
nand UO_2358 (O_2358,N_29313,N_29566);
nor UO_2359 (O_2359,N_29035,N_29693);
nor UO_2360 (O_2360,N_29027,N_29065);
or UO_2361 (O_2361,N_29469,N_28601);
nor UO_2362 (O_2362,N_28903,N_29908);
nand UO_2363 (O_2363,N_29491,N_28989);
xnor UO_2364 (O_2364,N_29504,N_28963);
or UO_2365 (O_2365,N_28618,N_29138);
xor UO_2366 (O_2366,N_28537,N_29409);
and UO_2367 (O_2367,N_29218,N_28677);
nor UO_2368 (O_2368,N_29555,N_28622);
nand UO_2369 (O_2369,N_29988,N_29149);
nor UO_2370 (O_2370,N_29620,N_28524);
xor UO_2371 (O_2371,N_29516,N_29078);
and UO_2372 (O_2372,N_29249,N_29701);
nor UO_2373 (O_2373,N_29003,N_28502);
xnor UO_2374 (O_2374,N_29207,N_28886);
xor UO_2375 (O_2375,N_28521,N_29605);
nand UO_2376 (O_2376,N_29131,N_29495);
nand UO_2377 (O_2377,N_29152,N_29093);
xnor UO_2378 (O_2378,N_29561,N_29525);
xnor UO_2379 (O_2379,N_29816,N_28519);
xnor UO_2380 (O_2380,N_28870,N_29580);
and UO_2381 (O_2381,N_29586,N_29094);
and UO_2382 (O_2382,N_28509,N_29965);
nor UO_2383 (O_2383,N_29617,N_29809);
or UO_2384 (O_2384,N_28913,N_29311);
nor UO_2385 (O_2385,N_28991,N_28786);
nand UO_2386 (O_2386,N_29892,N_28962);
nor UO_2387 (O_2387,N_29834,N_29761);
xor UO_2388 (O_2388,N_29698,N_29379);
or UO_2389 (O_2389,N_29865,N_29175);
nand UO_2390 (O_2390,N_28507,N_28660);
nor UO_2391 (O_2391,N_29913,N_29125);
and UO_2392 (O_2392,N_29630,N_29137);
and UO_2393 (O_2393,N_28793,N_28541);
nand UO_2394 (O_2394,N_28568,N_29531);
xor UO_2395 (O_2395,N_28540,N_28800);
nor UO_2396 (O_2396,N_29194,N_28655);
or UO_2397 (O_2397,N_29321,N_29568);
xnor UO_2398 (O_2398,N_28673,N_28974);
xnor UO_2399 (O_2399,N_28550,N_28757);
or UO_2400 (O_2400,N_28689,N_29586);
and UO_2401 (O_2401,N_29891,N_28511);
nand UO_2402 (O_2402,N_28950,N_29790);
nor UO_2403 (O_2403,N_28702,N_28731);
and UO_2404 (O_2404,N_29848,N_28702);
nor UO_2405 (O_2405,N_28659,N_29751);
or UO_2406 (O_2406,N_29758,N_28995);
or UO_2407 (O_2407,N_29960,N_28926);
xnor UO_2408 (O_2408,N_29520,N_29859);
nor UO_2409 (O_2409,N_29663,N_28959);
nand UO_2410 (O_2410,N_29050,N_28597);
or UO_2411 (O_2411,N_29538,N_29997);
xor UO_2412 (O_2412,N_29693,N_29320);
nand UO_2413 (O_2413,N_28820,N_29300);
xnor UO_2414 (O_2414,N_28830,N_29120);
nor UO_2415 (O_2415,N_29809,N_29563);
or UO_2416 (O_2416,N_29671,N_29040);
xor UO_2417 (O_2417,N_29753,N_28528);
xnor UO_2418 (O_2418,N_29246,N_29665);
and UO_2419 (O_2419,N_28756,N_29605);
nor UO_2420 (O_2420,N_29964,N_29162);
nor UO_2421 (O_2421,N_29347,N_29765);
or UO_2422 (O_2422,N_29459,N_29944);
nor UO_2423 (O_2423,N_29737,N_28830);
nor UO_2424 (O_2424,N_29565,N_29641);
nand UO_2425 (O_2425,N_28673,N_29319);
nor UO_2426 (O_2426,N_29261,N_28808);
or UO_2427 (O_2427,N_28863,N_28615);
nor UO_2428 (O_2428,N_29483,N_29847);
and UO_2429 (O_2429,N_29611,N_29067);
nor UO_2430 (O_2430,N_29136,N_29080);
or UO_2431 (O_2431,N_28668,N_29164);
nand UO_2432 (O_2432,N_29450,N_29749);
nor UO_2433 (O_2433,N_29521,N_28597);
and UO_2434 (O_2434,N_29188,N_29995);
xnor UO_2435 (O_2435,N_29059,N_29923);
nor UO_2436 (O_2436,N_29647,N_28741);
xnor UO_2437 (O_2437,N_29901,N_29689);
nor UO_2438 (O_2438,N_29156,N_29420);
and UO_2439 (O_2439,N_29610,N_29497);
nand UO_2440 (O_2440,N_29372,N_29768);
nand UO_2441 (O_2441,N_28656,N_29709);
or UO_2442 (O_2442,N_29359,N_29337);
nor UO_2443 (O_2443,N_29339,N_28540);
xor UO_2444 (O_2444,N_29105,N_28603);
nand UO_2445 (O_2445,N_29876,N_28728);
xor UO_2446 (O_2446,N_29872,N_28578);
nand UO_2447 (O_2447,N_28521,N_29345);
and UO_2448 (O_2448,N_29668,N_29940);
or UO_2449 (O_2449,N_29112,N_29191);
or UO_2450 (O_2450,N_28513,N_28930);
nor UO_2451 (O_2451,N_28966,N_29243);
xor UO_2452 (O_2452,N_29263,N_29441);
nor UO_2453 (O_2453,N_29387,N_29614);
and UO_2454 (O_2454,N_29573,N_28876);
xnor UO_2455 (O_2455,N_29159,N_28751);
nor UO_2456 (O_2456,N_29559,N_28732);
and UO_2457 (O_2457,N_29554,N_29520);
nor UO_2458 (O_2458,N_29684,N_29360);
or UO_2459 (O_2459,N_29747,N_29157);
or UO_2460 (O_2460,N_29011,N_29616);
or UO_2461 (O_2461,N_28667,N_29442);
nor UO_2462 (O_2462,N_29725,N_29492);
nand UO_2463 (O_2463,N_28758,N_29971);
nor UO_2464 (O_2464,N_28556,N_28946);
or UO_2465 (O_2465,N_29443,N_28601);
and UO_2466 (O_2466,N_29172,N_29645);
nand UO_2467 (O_2467,N_28531,N_29455);
nand UO_2468 (O_2468,N_28808,N_29404);
nor UO_2469 (O_2469,N_29193,N_28888);
nor UO_2470 (O_2470,N_28720,N_29505);
and UO_2471 (O_2471,N_28647,N_29211);
xnor UO_2472 (O_2472,N_29701,N_29825);
xnor UO_2473 (O_2473,N_28865,N_29494);
nor UO_2474 (O_2474,N_29242,N_28775);
nor UO_2475 (O_2475,N_29066,N_28550);
and UO_2476 (O_2476,N_29341,N_29781);
nor UO_2477 (O_2477,N_28612,N_29101);
and UO_2478 (O_2478,N_28824,N_28652);
or UO_2479 (O_2479,N_28778,N_28612);
xor UO_2480 (O_2480,N_29498,N_29716);
or UO_2481 (O_2481,N_29913,N_29385);
nand UO_2482 (O_2482,N_29388,N_29520);
or UO_2483 (O_2483,N_29297,N_29776);
nor UO_2484 (O_2484,N_29166,N_28559);
or UO_2485 (O_2485,N_28601,N_28728);
nand UO_2486 (O_2486,N_29395,N_28643);
xor UO_2487 (O_2487,N_28647,N_29543);
nand UO_2488 (O_2488,N_29199,N_29129);
nand UO_2489 (O_2489,N_28632,N_28653);
nor UO_2490 (O_2490,N_29224,N_29307);
and UO_2491 (O_2491,N_28515,N_28679);
and UO_2492 (O_2492,N_29638,N_28729);
xor UO_2493 (O_2493,N_29084,N_29821);
nor UO_2494 (O_2494,N_29253,N_29776);
nor UO_2495 (O_2495,N_29071,N_28740);
or UO_2496 (O_2496,N_29854,N_28593);
and UO_2497 (O_2497,N_29742,N_28864);
nand UO_2498 (O_2498,N_28600,N_29691);
or UO_2499 (O_2499,N_29731,N_28525);
xor UO_2500 (O_2500,N_29915,N_29690);
xor UO_2501 (O_2501,N_29952,N_29937);
nor UO_2502 (O_2502,N_29334,N_28926);
and UO_2503 (O_2503,N_29820,N_29900);
or UO_2504 (O_2504,N_29632,N_29877);
and UO_2505 (O_2505,N_29129,N_28799);
nand UO_2506 (O_2506,N_28787,N_29771);
nor UO_2507 (O_2507,N_29500,N_29919);
nor UO_2508 (O_2508,N_29299,N_28966);
or UO_2509 (O_2509,N_29102,N_29366);
xnor UO_2510 (O_2510,N_28981,N_28973);
or UO_2511 (O_2511,N_29472,N_29712);
and UO_2512 (O_2512,N_29630,N_29610);
nor UO_2513 (O_2513,N_29158,N_28794);
and UO_2514 (O_2514,N_29868,N_29660);
xnor UO_2515 (O_2515,N_29315,N_29987);
and UO_2516 (O_2516,N_29661,N_29570);
nor UO_2517 (O_2517,N_28874,N_28771);
nand UO_2518 (O_2518,N_29085,N_28954);
and UO_2519 (O_2519,N_29189,N_29284);
nand UO_2520 (O_2520,N_29073,N_28692);
xnor UO_2521 (O_2521,N_29602,N_29278);
and UO_2522 (O_2522,N_28593,N_28929);
and UO_2523 (O_2523,N_29529,N_28892);
nand UO_2524 (O_2524,N_29028,N_29205);
or UO_2525 (O_2525,N_28574,N_29255);
nand UO_2526 (O_2526,N_29286,N_28957);
nand UO_2527 (O_2527,N_28682,N_28920);
nor UO_2528 (O_2528,N_28530,N_28522);
or UO_2529 (O_2529,N_28797,N_29403);
or UO_2530 (O_2530,N_29077,N_29984);
xor UO_2531 (O_2531,N_29300,N_29607);
and UO_2532 (O_2532,N_28961,N_29098);
nand UO_2533 (O_2533,N_29808,N_29374);
and UO_2534 (O_2534,N_28546,N_28671);
and UO_2535 (O_2535,N_28771,N_28879);
xor UO_2536 (O_2536,N_29295,N_29269);
nor UO_2537 (O_2537,N_29935,N_28902);
nand UO_2538 (O_2538,N_28774,N_29685);
nor UO_2539 (O_2539,N_29420,N_29205);
nor UO_2540 (O_2540,N_29701,N_28787);
nor UO_2541 (O_2541,N_28814,N_29951);
and UO_2542 (O_2542,N_29166,N_29146);
xnor UO_2543 (O_2543,N_29745,N_29645);
xnor UO_2544 (O_2544,N_28537,N_29444);
and UO_2545 (O_2545,N_29491,N_29384);
nand UO_2546 (O_2546,N_28746,N_28642);
xor UO_2547 (O_2547,N_29561,N_29587);
and UO_2548 (O_2548,N_28635,N_28954);
or UO_2549 (O_2549,N_28667,N_29869);
xor UO_2550 (O_2550,N_29419,N_29450);
nand UO_2551 (O_2551,N_29509,N_28842);
nand UO_2552 (O_2552,N_29294,N_28872);
xor UO_2553 (O_2553,N_29878,N_29899);
and UO_2554 (O_2554,N_28942,N_29752);
xor UO_2555 (O_2555,N_28570,N_29454);
and UO_2556 (O_2556,N_28891,N_28555);
and UO_2557 (O_2557,N_28714,N_29076);
nor UO_2558 (O_2558,N_29991,N_28580);
xor UO_2559 (O_2559,N_29172,N_29307);
xor UO_2560 (O_2560,N_29149,N_28872);
nor UO_2561 (O_2561,N_29948,N_29738);
xor UO_2562 (O_2562,N_28849,N_28993);
xnor UO_2563 (O_2563,N_28586,N_28636);
xor UO_2564 (O_2564,N_29629,N_29036);
nor UO_2565 (O_2565,N_29062,N_28774);
nor UO_2566 (O_2566,N_29113,N_29598);
nor UO_2567 (O_2567,N_29291,N_29105);
xnor UO_2568 (O_2568,N_29385,N_28508);
nand UO_2569 (O_2569,N_29350,N_29545);
and UO_2570 (O_2570,N_29580,N_29808);
nand UO_2571 (O_2571,N_28694,N_28524);
nand UO_2572 (O_2572,N_28994,N_28691);
nor UO_2573 (O_2573,N_29999,N_29931);
nand UO_2574 (O_2574,N_28654,N_29765);
nand UO_2575 (O_2575,N_29192,N_29540);
or UO_2576 (O_2576,N_29283,N_29568);
nand UO_2577 (O_2577,N_29608,N_29634);
or UO_2578 (O_2578,N_29604,N_29291);
nor UO_2579 (O_2579,N_29894,N_29550);
xor UO_2580 (O_2580,N_29886,N_28542);
and UO_2581 (O_2581,N_29806,N_29873);
nand UO_2582 (O_2582,N_29618,N_29628);
and UO_2583 (O_2583,N_29593,N_29602);
and UO_2584 (O_2584,N_28922,N_29072);
xor UO_2585 (O_2585,N_28838,N_29191);
nor UO_2586 (O_2586,N_29318,N_29692);
and UO_2587 (O_2587,N_29328,N_28771);
xnor UO_2588 (O_2588,N_29123,N_28754);
nand UO_2589 (O_2589,N_29937,N_28862);
nor UO_2590 (O_2590,N_29587,N_29114);
nand UO_2591 (O_2591,N_29908,N_29718);
xnor UO_2592 (O_2592,N_29798,N_28580);
nand UO_2593 (O_2593,N_29097,N_29365);
nand UO_2594 (O_2594,N_28820,N_28669);
nand UO_2595 (O_2595,N_29686,N_28760);
or UO_2596 (O_2596,N_29673,N_28883);
nor UO_2597 (O_2597,N_29987,N_28792);
or UO_2598 (O_2598,N_29171,N_29120);
nand UO_2599 (O_2599,N_29203,N_29958);
and UO_2600 (O_2600,N_28822,N_29155);
xor UO_2601 (O_2601,N_29258,N_29264);
or UO_2602 (O_2602,N_28506,N_28700);
nor UO_2603 (O_2603,N_29508,N_29433);
or UO_2604 (O_2604,N_29419,N_28786);
or UO_2605 (O_2605,N_28593,N_28577);
xnor UO_2606 (O_2606,N_28923,N_29101);
nand UO_2607 (O_2607,N_29474,N_29542);
or UO_2608 (O_2608,N_28880,N_29200);
xnor UO_2609 (O_2609,N_29285,N_28567);
nand UO_2610 (O_2610,N_29565,N_29245);
or UO_2611 (O_2611,N_28755,N_29705);
nand UO_2612 (O_2612,N_29132,N_29919);
xnor UO_2613 (O_2613,N_28751,N_28863);
xnor UO_2614 (O_2614,N_29849,N_29039);
or UO_2615 (O_2615,N_28731,N_29973);
nor UO_2616 (O_2616,N_28538,N_29048);
or UO_2617 (O_2617,N_29424,N_29232);
nor UO_2618 (O_2618,N_29468,N_28617);
xor UO_2619 (O_2619,N_29811,N_29401);
or UO_2620 (O_2620,N_28516,N_29970);
nor UO_2621 (O_2621,N_29602,N_29025);
nand UO_2622 (O_2622,N_28944,N_29322);
nor UO_2623 (O_2623,N_29505,N_28535);
nand UO_2624 (O_2624,N_29354,N_28515);
nor UO_2625 (O_2625,N_29462,N_29313);
and UO_2626 (O_2626,N_29344,N_29318);
nand UO_2627 (O_2627,N_29350,N_29459);
or UO_2628 (O_2628,N_29355,N_29329);
xor UO_2629 (O_2629,N_29786,N_28906);
nand UO_2630 (O_2630,N_29042,N_28651);
and UO_2631 (O_2631,N_29522,N_28922);
nor UO_2632 (O_2632,N_29202,N_29302);
or UO_2633 (O_2633,N_28890,N_29671);
nor UO_2634 (O_2634,N_28735,N_29612);
xnor UO_2635 (O_2635,N_28761,N_29859);
nor UO_2636 (O_2636,N_28916,N_29500);
nor UO_2637 (O_2637,N_29793,N_29409);
nor UO_2638 (O_2638,N_29949,N_28755);
and UO_2639 (O_2639,N_29209,N_29911);
nor UO_2640 (O_2640,N_28974,N_28968);
nor UO_2641 (O_2641,N_28940,N_29841);
and UO_2642 (O_2642,N_28786,N_29249);
nand UO_2643 (O_2643,N_29157,N_29143);
and UO_2644 (O_2644,N_29228,N_29301);
and UO_2645 (O_2645,N_28871,N_29561);
nand UO_2646 (O_2646,N_29502,N_29482);
nand UO_2647 (O_2647,N_28746,N_28553);
or UO_2648 (O_2648,N_29443,N_29812);
xor UO_2649 (O_2649,N_29796,N_28663);
nor UO_2650 (O_2650,N_28840,N_29276);
nand UO_2651 (O_2651,N_29036,N_28582);
or UO_2652 (O_2652,N_29874,N_28866);
and UO_2653 (O_2653,N_29347,N_28886);
nor UO_2654 (O_2654,N_29478,N_29409);
or UO_2655 (O_2655,N_29882,N_29460);
nor UO_2656 (O_2656,N_28883,N_28512);
or UO_2657 (O_2657,N_28691,N_29588);
xor UO_2658 (O_2658,N_29005,N_29647);
or UO_2659 (O_2659,N_28986,N_29281);
or UO_2660 (O_2660,N_29559,N_29282);
xnor UO_2661 (O_2661,N_29097,N_28709);
xnor UO_2662 (O_2662,N_29406,N_28970);
or UO_2663 (O_2663,N_28576,N_28594);
nor UO_2664 (O_2664,N_29448,N_29491);
xor UO_2665 (O_2665,N_28949,N_29823);
nand UO_2666 (O_2666,N_29554,N_29954);
xnor UO_2667 (O_2667,N_29336,N_29839);
nand UO_2668 (O_2668,N_29142,N_29664);
nor UO_2669 (O_2669,N_29256,N_29269);
nand UO_2670 (O_2670,N_29270,N_28616);
xor UO_2671 (O_2671,N_29517,N_28980);
or UO_2672 (O_2672,N_29168,N_29364);
or UO_2673 (O_2673,N_29803,N_29097);
or UO_2674 (O_2674,N_28994,N_29869);
nand UO_2675 (O_2675,N_29935,N_29927);
or UO_2676 (O_2676,N_29350,N_29214);
xor UO_2677 (O_2677,N_28524,N_29897);
nand UO_2678 (O_2678,N_29989,N_29513);
nor UO_2679 (O_2679,N_29842,N_29173);
nor UO_2680 (O_2680,N_29847,N_29077);
xor UO_2681 (O_2681,N_29572,N_28633);
nand UO_2682 (O_2682,N_28646,N_29134);
nor UO_2683 (O_2683,N_29494,N_29454);
nor UO_2684 (O_2684,N_29559,N_28557);
nand UO_2685 (O_2685,N_29222,N_28544);
or UO_2686 (O_2686,N_29747,N_29033);
and UO_2687 (O_2687,N_28645,N_28666);
and UO_2688 (O_2688,N_28717,N_28653);
nand UO_2689 (O_2689,N_29465,N_28663);
nand UO_2690 (O_2690,N_29994,N_29796);
nor UO_2691 (O_2691,N_28549,N_28895);
nand UO_2692 (O_2692,N_29271,N_29304);
nor UO_2693 (O_2693,N_29330,N_29441);
or UO_2694 (O_2694,N_28882,N_28533);
or UO_2695 (O_2695,N_29977,N_29615);
nand UO_2696 (O_2696,N_29844,N_29083);
and UO_2697 (O_2697,N_28982,N_29109);
or UO_2698 (O_2698,N_29857,N_28898);
or UO_2699 (O_2699,N_29871,N_29042);
nor UO_2700 (O_2700,N_29921,N_29286);
and UO_2701 (O_2701,N_29363,N_29368);
or UO_2702 (O_2702,N_29022,N_28995);
or UO_2703 (O_2703,N_29876,N_28773);
nand UO_2704 (O_2704,N_29100,N_29399);
xor UO_2705 (O_2705,N_28693,N_29440);
nor UO_2706 (O_2706,N_29031,N_28593);
or UO_2707 (O_2707,N_28660,N_29496);
nand UO_2708 (O_2708,N_29707,N_29660);
and UO_2709 (O_2709,N_28553,N_29939);
xor UO_2710 (O_2710,N_29193,N_29727);
nand UO_2711 (O_2711,N_28765,N_28907);
or UO_2712 (O_2712,N_29311,N_28592);
nor UO_2713 (O_2713,N_29367,N_29501);
and UO_2714 (O_2714,N_29002,N_29767);
nor UO_2715 (O_2715,N_28899,N_28704);
nand UO_2716 (O_2716,N_29644,N_28720);
and UO_2717 (O_2717,N_29822,N_29023);
nor UO_2718 (O_2718,N_28736,N_29535);
nand UO_2719 (O_2719,N_29112,N_29052);
or UO_2720 (O_2720,N_29732,N_29951);
nor UO_2721 (O_2721,N_28518,N_29174);
or UO_2722 (O_2722,N_28913,N_29870);
nand UO_2723 (O_2723,N_29657,N_29615);
nand UO_2724 (O_2724,N_29643,N_28645);
xor UO_2725 (O_2725,N_29885,N_29770);
or UO_2726 (O_2726,N_28949,N_29321);
and UO_2727 (O_2727,N_29414,N_29881);
xor UO_2728 (O_2728,N_28601,N_28694);
nand UO_2729 (O_2729,N_29919,N_29579);
nor UO_2730 (O_2730,N_29876,N_29920);
xor UO_2731 (O_2731,N_29611,N_28948);
xor UO_2732 (O_2732,N_28758,N_29948);
and UO_2733 (O_2733,N_29988,N_29873);
xor UO_2734 (O_2734,N_28725,N_29609);
xor UO_2735 (O_2735,N_28625,N_29195);
nor UO_2736 (O_2736,N_29595,N_28666);
xor UO_2737 (O_2737,N_29561,N_29270);
nor UO_2738 (O_2738,N_28527,N_29792);
nand UO_2739 (O_2739,N_29402,N_29181);
xnor UO_2740 (O_2740,N_29617,N_29099);
nand UO_2741 (O_2741,N_28692,N_29402);
xnor UO_2742 (O_2742,N_29049,N_28528);
xnor UO_2743 (O_2743,N_29822,N_28763);
nand UO_2744 (O_2744,N_29879,N_29214);
or UO_2745 (O_2745,N_28756,N_29857);
xor UO_2746 (O_2746,N_28804,N_29958);
nand UO_2747 (O_2747,N_28565,N_29854);
nor UO_2748 (O_2748,N_28826,N_29012);
nor UO_2749 (O_2749,N_29089,N_29761);
xor UO_2750 (O_2750,N_29989,N_29516);
or UO_2751 (O_2751,N_28636,N_29917);
nand UO_2752 (O_2752,N_29167,N_29355);
nand UO_2753 (O_2753,N_29329,N_28944);
nand UO_2754 (O_2754,N_29807,N_29185);
xor UO_2755 (O_2755,N_29531,N_28544);
nor UO_2756 (O_2756,N_29299,N_29942);
xor UO_2757 (O_2757,N_29992,N_28758);
or UO_2758 (O_2758,N_28906,N_28584);
or UO_2759 (O_2759,N_29994,N_29239);
and UO_2760 (O_2760,N_29691,N_29383);
nand UO_2761 (O_2761,N_29602,N_28656);
nor UO_2762 (O_2762,N_29710,N_29351);
nor UO_2763 (O_2763,N_29577,N_29579);
nor UO_2764 (O_2764,N_28916,N_28639);
nand UO_2765 (O_2765,N_29990,N_28663);
and UO_2766 (O_2766,N_29734,N_29454);
nor UO_2767 (O_2767,N_29357,N_29300);
and UO_2768 (O_2768,N_29932,N_29717);
nor UO_2769 (O_2769,N_29557,N_29262);
nor UO_2770 (O_2770,N_28528,N_29556);
or UO_2771 (O_2771,N_29490,N_29445);
nor UO_2772 (O_2772,N_28823,N_28551);
nand UO_2773 (O_2773,N_28762,N_29855);
and UO_2774 (O_2774,N_29778,N_29482);
and UO_2775 (O_2775,N_29935,N_29487);
and UO_2776 (O_2776,N_29545,N_29373);
nand UO_2777 (O_2777,N_28731,N_29141);
or UO_2778 (O_2778,N_29546,N_29959);
nand UO_2779 (O_2779,N_29927,N_28907);
and UO_2780 (O_2780,N_29530,N_29324);
and UO_2781 (O_2781,N_29775,N_29044);
xor UO_2782 (O_2782,N_29470,N_29220);
nor UO_2783 (O_2783,N_29893,N_29646);
and UO_2784 (O_2784,N_29800,N_29092);
xnor UO_2785 (O_2785,N_28788,N_29876);
nor UO_2786 (O_2786,N_28843,N_29738);
or UO_2787 (O_2787,N_29661,N_28597);
nor UO_2788 (O_2788,N_29413,N_28973);
nor UO_2789 (O_2789,N_28595,N_29119);
or UO_2790 (O_2790,N_29066,N_29543);
nor UO_2791 (O_2791,N_29137,N_29620);
or UO_2792 (O_2792,N_29884,N_29253);
or UO_2793 (O_2793,N_28506,N_28782);
xnor UO_2794 (O_2794,N_29208,N_28754);
or UO_2795 (O_2795,N_28625,N_29972);
nand UO_2796 (O_2796,N_29752,N_29726);
or UO_2797 (O_2797,N_29350,N_29660);
nand UO_2798 (O_2798,N_29941,N_29208);
or UO_2799 (O_2799,N_28980,N_29321);
or UO_2800 (O_2800,N_29431,N_28699);
nand UO_2801 (O_2801,N_29780,N_29192);
xor UO_2802 (O_2802,N_29583,N_29661);
xnor UO_2803 (O_2803,N_29279,N_29269);
nor UO_2804 (O_2804,N_28545,N_28788);
or UO_2805 (O_2805,N_28609,N_29822);
nand UO_2806 (O_2806,N_28528,N_29125);
or UO_2807 (O_2807,N_28999,N_28911);
nor UO_2808 (O_2808,N_28644,N_28841);
or UO_2809 (O_2809,N_29825,N_29147);
xor UO_2810 (O_2810,N_29009,N_29013);
and UO_2811 (O_2811,N_29203,N_28916);
or UO_2812 (O_2812,N_29023,N_29747);
and UO_2813 (O_2813,N_28802,N_28939);
and UO_2814 (O_2814,N_28939,N_29267);
nand UO_2815 (O_2815,N_29122,N_29271);
or UO_2816 (O_2816,N_29757,N_29273);
and UO_2817 (O_2817,N_28900,N_29029);
and UO_2818 (O_2818,N_29351,N_29254);
nand UO_2819 (O_2819,N_28972,N_29322);
nand UO_2820 (O_2820,N_28777,N_28644);
and UO_2821 (O_2821,N_28787,N_28761);
or UO_2822 (O_2822,N_29999,N_29408);
and UO_2823 (O_2823,N_29255,N_29593);
nor UO_2824 (O_2824,N_29763,N_29876);
nand UO_2825 (O_2825,N_29164,N_28867);
nand UO_2826 (O_2826,N_28970,N_29728);
nand UO_2827 (O_2827,N_29640,N_29743);
xor UO_2828 (O_2828,N_29215,N_29768);
and UO_2829 (O_2829,N_29876,N_29554);
or UO_2830 (O_2830,N_28741,N_28838);
nand UO_2831 (O_2831,N_28770,N_28610);
nand UO_2832 (O_2832,N_28859,N_28624);
nand UO_2833 (O_2833,N_29747,N_29095);
nor UO_2834 (O_2834,N_29552,N_28897);
or UO_2835 (O_2835,N_29766,N_29381);
nand UO_2836 (O_2836,N_29035,N_29770);
xor UO_2837 (O_2837,N_29426,N_28738);
xnor UO_2838 (O_2838,N_29096,N_28550);
nor UO_2839 (O_2839,N_28941,N_29747);
nand UO_2840 (O_2840,N_28803,N_29658);
xor UO_2841 (O_2841,N_29638,N_29876);
nor UO_2842 (O_2842,N_29903,N_29239);
nor UO_2843 (O_2843,N_29822,N_28662);
and UO_2844 (O_2844,N_29168,N_28847);
nand UO_2845 (O_2845,N_28891,N_28996);
nor UO_2846 (O_2846,N_29526,N_29869);
xnor UO_2847 (O_2847,N_28803,N_28790);
or UO_2848 (O_2848,N_29401,N_28545);
nand UO_2849 (O_2849,N_28805,N_28605);
nand UO_2850 (O_2850,N_29043,N_28564);
xnor UO_2851 (O_2851,N_29886,N_28926);
nand UO_2852 (O_2852,N_29596,N_29769);
or UO_2853 (O_2853,N_29066,N_29415);
nor UO_2854 (O_2854,N_28802,N_29766);
nand UO_2855 (O_2855,N_29385,N_28745);
or UO_2856 (O_2856,N_28663,N_28605);
xor UO_2857 (O_2857,N_29838,N_29542);
or UO_2858 (O_2858,N_28665,N_29536);
nand UO_2859 (O_2859,N_28779,N_29805);
or UO_2860 (O_2860,N_28755,N_28867);
xor UO_2861 (O_2861,N_29453,N_28953);
xor UO_2862 (O_2862,N_29895,N_29226);
and UO_2863 (O_2863,N_29195,N_29662);
or UO_2864 (O_2864,N_29982,N_29874);
nor UO_2865 (O_2865,N_29596,N_29053);
nor UO_2866 (O_2866,N_28802,N_29151);
or UO_2867 (O_2867,N_29638,N_29969);
nor UO_2868 (O_2868,N_28835,N_28988);
and UO_2869 (O_2869,N_28650,N_28992);
nor UO_2870 (O_2870,N_29863,N_28883);
and UO_2871 (O_2871,N_28502,N_29152);
and UO_2872 (O_2872,N_29196,N_28931);
nand UO_2873 (O_2873,N_28792,N_29420);
nand UO_2874 (O_2874,N_29381,N_29166);
nand UO_2875 (O_2875,N_29537,N_29906);
or UO_2876 (O_2876,N_29037,N_29100);
nor UO_2877 (O_2877,N_29979,N_29027);
or UO_2878 (O_2878,N_29164,N_29490);
nor UO_2879 (O_2879,N_29823,N_29786);
nand UO_2880 (O_2880,N_28749,N_29058);
and UO_2881 (O_2881,N_29425,N_28924);
nor UO_2882 (O_2882,N_28909,N_29778);
nand UO_2883 (O_2883,N_29291,N_28715);
nand UO_2884 (O_2884,N_29710,N_29458);
and UO_2885 (O_2885,N_28644,N_29718);
and UO_2886 (O_2886,N_28701,N_29558);
xnor UO_2887 (O_2887,N_29568,N_28827);
nand UO_2888 (O_2888,N_28823,N_29451);
or UO_2889 (O_2889,N_29297,N_28985);
nor UO_2890 (O_2890,N_29627,N_29374);
xor UO_2891 (O_2891,N_29065,N_28604);
or UO_2892 (O_2892,N_28892,N_29334);
and UO_2893 (O_2893,N_29328,N_28530);
nand UO_2894 (O_2894,N_29284,N_29861);
nand UO_2895 (O_2895,N_28978,N_29005);
or UO_2896 (O_2896,N_29592,N_29107);
xnor UO_2897 (O_2897,N_29597,N_29357);
xnor UO_2898 (O_2898,N_29583,N_28556);
or UO_2899 (O_2899,N_29072,N_28994);
nor UO_2900 (O_2900,N_29149,N_29053);
and UO_2901 (O_2901,N_29782,N_28915);
xnor UO_2902 (O_2902,N_28715,N_29626);
nand UO_2903 (O_2903,N_29347,N_28648);
nand UO_2904 (O_2904,N_29279,N_28621);
xor UO_2905 (O_2905,N_29711,N_29888);
nor UO_2906 (O_2906,N_29622,N_29385);
or UO_2907 (O_2907,N_28755,N_29994);
xor UO_2908 (O_2908,N_28819,N_29324);
xnor UO_2909 (O_2909,N_28513,N_29285);
or UO_2910 (O_2910,N_29951,N_28770);
or UO_2911 (O_2911,N_28667,N_29793);
nor UO_2912 (O_2912,N_29798,N_28989);
nand UO_2913 (O_2913,N_29501,N_29518);
or UO_2914 (O_2914,N_29170,N_29362);
nand UO_2915 (O_2915,N_28506,N_29820);
xor UO_2916 (O_2916,N_29891,N_29666);
and UO_2917 (O_2917,N_28717,N_29164);
or UO_2918 (O_2918,N_29078,N_29428);
or UO_2919 (O_2919,N_28835,N_29411);
and UO_2920 (O_2920,N_28510,N_28792);
or UO_2921 (O_2921,N_29706,N_29578);
nand UO_2922 (O_2922,N_29229,N_29249);
nor UO_2923 (O_2923,N_29459,N_28637);
and UO_2924 (O_2924,N_28762,N_29181);
and UO_2925 (O_2925,N_29313,N_28604);
and UO_2926 (O_2926,N_29752,N_28507);
nor UO_2927 (O_2927,N_29275,N_29266);
nor UO_2928 (O_2928,N_28503,N_29301);
nand UO_2929 (O_2929,N_28734,N_29442);
or UO_2930 (O_2930,N_28637,N_29311);
xor UO_2931 (O_2931,N_29048,N_28636);
and UO_2932 (O_2932,N_29519,N_28926);
and UO_2933 (O_2933,N_29559,N_28728);
xor UO_2934 (O_2934,N_29645,N_29877);
nor UO_2935 (O_2935,N_29655,N_28612);
xor UO_2936 (O_2936,N_29016,N_29315);
and UO_2937 (O_2937,N_29573,N_29636);
nor UO_2938 (O_2938,N_29714,N_29866);
nor UO_2939 (O_2939,N_29139,N_28735);
xnor UO_2940 (O_2940,N_29047,N_29513);
nor UO_2941 (O_2941,N_29750,N_29712);
nor UO_2942 (O_2942,N_29740,N_28759);
and UO_2943 (O_2943,N_28529,N_29406);
or UO_2944 (O_2944,N_28598,N_29057);
nand UO_2945 (O_2945,N_28558,N_29361);
nand UO_2946 (O_2946,N_29125,N_29168);
or UO_2947 (O_2947,N_29858,N_28816);
nor UO_2948 (O_2948,N_29677,N_28624);
nand UO_2949 (O_2949,N_29413,N_29058);
nand UO_2950 (O_2950,N_28647,N_29800);
nand UO_2951 (O_2951,N_28650,N_29441);
or UO_2952 (O_2952,N_28946,N_29885);
or UO_2953 (O_2953,N_29003,N_28892);
xor UO_2954 (O_2954,N_29750,N_29359);
xor UO_2955 (O_2955,N_29188,N_28763);
nand UO_2956 (O_2956,N_29044,N_28613);
nand UO_2957 (O_2957,N_28653,N_28960);
nand UO_2958 (O_2958,N_29732,N_29419);
xor UO_2959 (O_2959,N_29503,N_29110);
nor UO_2960 (O_2960,N_28934,N_29910);
and UO_2961 (O_2961,N_29476,N_28700);
or UO_2962 (O_2962,N_28606,N_28990);
nor UO_2963 (O_2963,N_28873,N_29216);
nor UO_2964 (O_2964,N_29804,N_29205);
and UO_2965 (O_2965,N_29089,N_29069);
xnor UO_2966 (O_2966,N_28520,N_29541);
and UO_2967 (O_2967,N_29655,N_29251);
xor UO_2968 (O_2968,N_29096,N_29494);
nor UO_2969 (O_2969,N_28733,N_28700);
nand UO_2970 (O_2970,N_29825,N_28928);
nand UO_2971 (O_2971,N_29961,N_29689);
nor UO_2972 (O_2972,N_29967,N_29842);
or UO_2973 (O_2973,N_29950,N_28520);
or UO_2974 (O_2974,N_29160,N_29665);
or UO_2975 (O_2975,N_29120,N_29886);
or UO_2976 (O_2976,N_29220,N_28685);
nor UO_2977 (O_2977,N_29355,N_29890);
or UO_2978 (O_2978,N_29661,N_29565);
nor UO_2979 (O_2979,N_29745,N_29643);
xor UO_2980 (O_2980,N_29230,N_28947);
xor UO_2981 (O_2981,N_29494,N_28505);
xor UO_2982 (O_2982,N_29315,N_29245);
nor UO_2983 (O_2983,N_29979,N_28718);
nor UO_2984 (O_2984,N_29778,N_28637);
xnor UO_2985 (O_2985,N_29816,N_29093);
or UO_2986 (O_2986,N_28542,N_29150);
nand UO_2987 (O_2987,N_29968,N_29019);
xor UO_2988 (O_2988,N_29414,N_29768);
xnor UO_2989 (O_2989,N_28855,N_29206);
or UO_2990 (O_2990,N_29635,N_28663);
xor UO_2991 (O_2991,N_29049,N_29639);
xnor UO_2992 (O_2992,N_29970,N_29255);
or UO_2993 (O_2993,N_29527,N_28811);
nor UO_2994 (O_2994,N_28515,N_29623);
nor UO_2995 (O_2995,N_28928,N_28787);
nor UO_2996 (O_2996,N_29018,N_29418);
or UO_2997 (O_2997,N_28726,N_28797);
nor UO_2998 (O_2998,N_29927,N_29143);
or UO_2999 (O_2999,N_29536,N_28796);
nor UO_3000 (O_3000,N_29556,N_28973);
and UO_3001 (O_3001,N_29675,N_29841);
nor UO_3002 (O_3002,N_29008,N_28751);
nand UO_3003 (O_3003,N_28653,N_28737);
nor UO_3004 (O_3004,N_29890,N_29087);
or UO_3005 (O_3005,N_28684,N_29422);
xor UO_3006 (O_3006,N_29316,N_29326);
nor UO_3007 (O_3007,N_28695,N_29906);
nor UO_3008 (O_3008,N_29402,N_29928);
nor UO_3009 (O_3009,N_28545,N_28813);
nor UO_3010 (O_3010,N_28598,N_29819);
or UO_3011 (O_3011,N_29800,N_28765);
or UO_3012 (O_3012,N_29956,N_28688);
xor UO_3013 (O_3013,N_28982,N_29140);
xor UO_3014 (O_3014,N_28538,N_29026);
nand UO_3015 (O_3015,N_29953,N_28699);
xor UO_3016 (O_3016,N_29919,N_29889);
and UO_3017 (O_3017,N_29091,N_28599);
or UO_3018 (O_3018,N_29225,N_29724);
nand UO_3019 (O_3019,N_29624,N_29213);
nand UO_3020 (O_3020,N_29371,N_28664);
nand UO_3021 (O_3021,N_28582,N_28905);
nand UO_3022 (O_3022,N_29352,N_29877);
nand UO_3023 (O_3023,N_29730,N_28662);
or UO_3024 (O_3024,N_29801,N_28758);
and UO_3025 (O_3025,N_29340,N_29977);
nand UO_3026 (O_3026,N_28637,N_28854);
xor UO_3027 (O_3027,N_29617,N_28587);
nor UO_3028 (O_3028,N_29821,N_29108);
xnor UO_3029 (O_3029,N_28634,N_29965);
or UO_3030 (O_3030,N_28704,N_29399);
nand UO_3031 (O_3031,N_29256,N_29546);
or UO_3032 (O_3032,N_29016,N_29385);
or UO_3033 (O_3033,N_29307,N_29150);
nor UO_3034 (O_3034,N_29483,N_29289);
and UO_3035 (O_3035,N_29183,N_28767);
or UO_3036 (O_3036,N_29674,N_29194);
nor UO_3037 (O_3037,N_29406,N_29690);
or UO_3038 (O_3038,N_28546,N_28524);
nand UO_3039 (O_3039,N_28649,N_29266);
nor UO_3040 (O_3040,N_29659,N_28622);
and UO_3041 (O_3041,N_29673,N_29887);
nor UO_3042 (O_3042,N_29658,N_29511);
and UO_3043 (O_3043,N_29644,N_28732);
or UO_3044 (O_3044,N_28990,N_29193);
and UO_3045 (O_3045,N_28584,N_29063);
nand UO_3046 (O_3046,N_29856,N_29499);
nand UO_3047 (O_3047,N_28790,N_29119);
and UO_3048 (O_3048,N_29572,N_29867);
nor UO_3049 (O_3049,N_29181,N_29439);
and UO_3050 (O_3050,N_29000,N_28534);
nand UO_3051 (O_3051,N_29866,N_29788);
xnor UO_3052 (O_3052,N_29933,N_28543);
or UO_3053 (O_3053,N_29162,N_29244);
and UO_3054 (O_3054,N_29501,N_29551);
and UO_3055 (O_3055,N_28520,N_28794);
or UO_3056 (O_3056,N_29737,N_29228);
xor UO_3057 (O_3057,N_29624,N_29367);
nand UO_3058 (O_3058,N_29679,N_28793);
xor UO_3059 (O_3059,N_28606,N_29272);
nand UO_3060 (O_3060,N_29893,N_29663);
nand UO_3061 (O_3061,N_28841,N_29987);
nor UO_3062 (O_3062,N_29517,N_29129);
xor UO_3063 (O_3063,N_29996,N_29120);
or UO_3064 (O_3064,N_28786,N_29752);
or UO_3065 (O_3065,N_29951,N_28699);
nor UO_3066 (O_3066,N_29416,N_29004);
xnor UO_3067 (O_3067,N_28920,N_28928);
nand UO_3068 (O_3068,N_28522,N_29462);
xor UO_3069 (O_3069,N_28608,N_29033);
or UO_3070 (O_3070,N_29275,N_29368);
xor UO_3071 (O_3071,N_28931,N_29707);
nor UO_3072 (O_3072,N_28871,N_29800);
and UO_3073 (O_3073,N_28717,N_29785);
nor UO_3074 (O_3074,N_29739,N_28884);
xor UO_3075 (O_3075,N_29961,N_29409);
or UO_3076 (O_3076,N_29703,N_29811);
and UO_3077 (O_3077,N_29357,N_29423);
or UO_3078 (O_3078,N_28836,N_29404);
and UO_3079 (O_3079,N_29741,N_29440);
or UO_3080 (O_3080,N_28733,N_28651);
or UO_3081 (O_3081,N_29796,N_29297);
nor UO_3082 (O_3082,N_29280,N_29602);
nand UO_3083 (O_3083,N_28875,N_29433);
nor UO_3084 (O_3084,N_28547,N_28535);
xor UO_3085 (O_3085,N_29639,N_29185);
nand UO_3086 (O_3086,N_29036,N_28616);
nand UO_3087 (O_3087,N_28603,N_28650);
or UO_3088 (O_3088,N_29983,N_29052);
nand UO_3089 (O_3089,N_29594,N_29246);
and UO_3090 (O_3090,N_28856,N_29091);
xor UO_3091 (O_3091,N_29329,N_28775);
or UO_3092 (O_3092,N_28668,N_29523);
nand UO_3093 (O_3093,N_29628,N_29082);
nand UO_3094 (O_3094,N_29848,N_28906);
or UO_3095 (O_3095,N_29015,N_29991);
nor UO_3096 (O_3096,N_28828,N_28865);
xor UO_3097 (O_3097,N_28908,N_29844);
nand UO_3098 (O_3098,N_28776,N_29160);
nor UO_3099 (O_3099,N_29587,N_28780);
nor UO_3100 (O_3100,N_29408,N_29340);
xnor UO_3101 (O_3101,N_29127,N_29382);
xnor UO_3102 (O_3102,N_29534,N_29180);
nor UO_3103 (O_3103,N_29423,N_29626);
nand UO_3104 (O_3104,N_29031,N_29124);
and UO_3105 (O_3105,N_29033,N_28842);
and UO_3106 (O_3106,N_29557,N_28610);
nand UO_3107 (O_3107,N_29761,N_29875);
nand UO_3108 (O_3108,N_28856,N_29092);
or UO_3109 (O_3109,N_29850,N_28575);
or UO_3110 (O_3110,N_28647,N_29187);
nor UO_3111 (O_3111,N_29873,N_28869);
nor UO_3112 (O_3112,N_29596,N_29266);
and UO_3113 (O_3113,N_29369,N_29672);
nand UO_3114 (O_3114,N_29303,N_29556);
or UO_3115 (O_3115,N_29099,N_29326);
nor UO_3116 (O_3116,N_29957,N_29669);
nand UO_3117 (O_3117,N_28587,N_29497);
or UO_3118 (O_3118,N_28524,N_28891);
xor UO_3119 (O_3119,N_29969,N_28763);
or UO_3120 (O_3120,N_29479,N_28851);
and UO_3121 (O_3121,N_28912,N_29629);
nand UO_3122 (O_3122,N_28520,N_28838);
and UO_3123 (O_3123,N_28835,N_29258);
or UO_3124 (O_3124,N_29228,N_29781);
xor UO_3125 (O_3125,N_28944,N_28771);
xor UO_3126 (O_3126,N_29936,N_29075);
and UO_3127 (O_3127,N_28952,N_28951);
or UO_3128 (O_3128,N_28938,N_29720);
xor UO_3129 (O_3129,N_28750,N_28904);
nand UO_3130 (O_3130,N_28869,N_29823);
nand UO_3131 (O_3131,N_28893,N_29952);
nor UO_3132 (O_3132,N_29753,N_29334);
nor UO_3133 (O_3133,N_29479,N_28694);
nor UO_3134 (O_3134,N_29636,N_28890);
and UO_3135 (O_3135,N_28513,N_29329);
xor UO_3136 (O_3136,N_29236,N_29416);
xor UO_3137 (O_3137,N_29267,N_28530);
xnor UO_3138 (O_3138,N_29615,N_29880);
nand UO_3139 (O_3139,N_29257,N_29048);
and UO_3140 (O_3140,N_28895,N_29692);
xnor UO_3141 (O_3141,N_28781,N_28615);
or UO_3142 (O_3142,N_28746,N_29842);
nor UO_3143 (O_3143,N_29355,N_29819);
nand UO_3144 (O_3144,N_29867,N_29334);
or UO_3145 (O_3145,N_29357,N_28500);
or UO_3146 (O_3146,N_28881,N_29082);
xor UO_3147 (O_3147,N_29138,N_29252);
and UO_3148 (O_3148,N_28907,N_28954);
nor UO_3149 (O_3149,N_29648,N_29039);
nor UO_3150 (O_3150,N_28567,N_29687);
nor UO_3151 (O_3151,N_29435,N_28605);
nor UO_3152 (O_3152,N_29247,N_29911);
and UO_3153 (O_3153,N_29432,N_29619);
and UO_3154 (O_3154,N_29466,N_28670);
nor UO_3155 (O_3155,N_29406,N_29497);
xor UO_3156 (O_3156,N_28669,N_29893);
nand UO_3157 (O_3157,N_29032,N_28959);
nand UO_3158 (O_3158,N_28962,N_29857);
nor UO_3159 (O_3159,N_29764,N_29932);
nor UO_3160 (O_3160,N_29341,N_28844);
nor UO_3161 (O_3161,N_29959,N_29673);
and UO_3162 (O_3162,N_28691,N_29790);
xor UO_3163 (O_3163,N_28905,N_29660);
nor UO_3164 (O_3164,N_29970,N_29439);
and UO_3165 (O_3165,N_28865,N_29293);
xor UO_3166 (O_3166,N_29095,N_28608);
xor UO_3167 (O_3167,N_29812,N_28675);
and UO_3168 (O_3168,N_29020,N_29719);
nand UO_3169 (O_3169,N_28632,N_28672);
xor UO_3170 (O_3170,N_29657,N_29472);
or UO_3171 (O_3171,N_28685,N_28799);
nand UO_3172 (O_3172,N_28822,N_28918);
nand UO_3173 (O_3173,N_28737,N_28977);
or UO_3174 (O_3174,N_28575,N_28563);
or UO_3175 (O_3175,N_29054,N_28697);
nand UO_3176 (O_3176,N_29378,N_29010);
and UO_3177 (O_3177,N_29031,N_29936);
or UO_3178 (O_3178,N_29076,N_28960);
or UO_3179 (O_3179,N_29465,N_29708);
nor UO_3180 (O_3180,N_28986,N_29843);
nor UO_3181 (O_3181,N_29840,N_29919);
and UO_3182 (O_3182,N_28682,N_28804);
and UO_3183 (O_3183,N_29488,N_29499);
and UO_3184 (O_3184,N_29532,N_29157);
xor UO_3185 (O_3185,N_28705,N_28546);
and UO_3186 (O_3186,N_28505,N_29116);
nor UO_3187 (O_3187,N_29851,N_29691);
and UO_3188 (O_3188,N_29553,N_29432);
or UO_3189 (O_3189,N_29772,N_28949);
or UO_3190 (O_3190,N_29562,N_29348);
xnor UO_3191 (O_3191,N_29285,N_29218);
or UO_3192 (O_3192,N_29185,N_29427);
nor UO_3193 (O_3193,N_28574,N_29097);
nand UO_3194 (O_3194,N_28792,N_29472);
or UO_3195 (O_3195,N_29086,N_29568);
xor UO_3196 (O_3196,N_29882,N_29569);
or UO_3197 (O_3197,N_29198,N_28999);
nor UO_3198 (O_3198,N_28648,N_29278);
nor UO_3199 (O_3199,N_29805,N_29444);
or UO_3200 (O_3200,N_29151,N_29604);
nand UO_3201 (O_3201,N_29134,N_29383);
and UO_3202 (O_3202,N_29844,N_29493);
xnor UO_3203 (O_3203,N_29563,N_28608);
xor UO_3204 (O_3204,N_29015,N_29436);
nor UO_3205 (O_3205,N_29366,N_29648);
nor UO_3206 (O_3206,N_28942,N_29801);
and UO_3207 (O_3207,N_29016,N_29416);
and UO_3208 (O_3208,N_29877,N_29395);
xnor UO_3209 (O_3209,N_29973,N_29849);
nand UO_3210 (O_3210,N_28717,N_29040);
nand UO_3211 (O_3211,N_29804,N_29319);
nor UO_3212 (O_3212,N_29176,N_28776);
or UO_3213 (O_3213,N_29217,N_29950);
or UO_3214 (O_3214,N_29672,N_29904);
nor UO_3215 (O_3215,N_28773,N_28695);
xnor UO_3216 (O_3216,N_29073,N_29748);
nor UO_3217 (O_3217,N_29540,N_28946);
or UO_3218 (O_3218,N_28837,N_29218);
and UO_3219 (O_3219,N_28504,N_29266);
nor UO_3220 (O_3220,N_29463,N_28843);
or UO_3221 (O_3221,N_29281,N_29906);
or UO_3222 (O_3222,N_29522,N_28985);
and UO_3223 (O_3223,N_29866,N_29810);
nand UO_3224 (O_3224,N_28544,N_29003);
and UO_3225 (O_3225,N_29489,N_29848);
or UO_3226 (O_3226,N_29137,N_29959);
or UO_3227 (O_3227,N_29963,N_29828);
xnor UO_3228 (O_3228,N_29272,N_28951);
nand UO_3229 (O_3229,N_28782,N_29666);
nand UO_3230 (O_3230,N_29745,N_29304);
and UO_3231 (O_3231,N_29106,N_28853);
and UO_3232 (O_3232,N_29897,N_28722);
nand UO_3233 (O_3233,N_28730,N_29033);
nand UO_3234 (O_3234,N_28896,N_28981);
or UO_3235 (O_3235,N_29646,N_29405);
xnor UO_3236 (O_3236,N_28764,N_29993);
nor UO_3237 (O_3237,N_29459,N_28509);
and UO_3238 (O_3238,N_29762,N_28586);
xor UO_3239 (O_3239,N_29188,N_29595);
nor UO_3240 (O_3240,N_29757,N_29089);
nand UO_3241 (O_3241,N_29272,N_29296);
xnor UO_3242 (O_3242,N_28634,N_29883);
and UO_3243 (O_3243,N_29533,N_29214);
and UO_3244 (O_3244,N_28941,N_28945);
nand UO_3245 (O_3245,N_28612,N_28677);
or UO_3246 (O_3246,N_29661,N_29090);
nor UO_3247 (O_3247,N_29924,N_29410);
and UO_3248 (O_3248,N_29122,N_29368);
xor UO_3249 (O_3249,N_29342,N_29230);
nand UO_3250 (O_3250,N_29564,N_28825);
xnor UO_3251 (O_3251,N_29224,N_29696);
and UO_3252 (O_3252,N_29889,N_29992);
or UO_3253 (O_3253,N_28866,N_29103);
xnor UO_3254 (O_3254,N_29277,N_29658);
nand UO_3255 (O_3255,N_29106,N_28521);
nand UO_3256 (O_3256,N_29984,N_29965);
nor UO_3257 (O_3257,N_28890,N_28881);
nand UO_3258 (O_3258,N_29634,N_29920);
or UO_3259 (O_3259,N_29762,N_28831);
xnor UO_3260 (O_3260,N_28882,N_29350);
nand UO_3261 (O_3261,N_29186,N_28863);
and UO_3262 (O_3262,N_29386,N_29939);
nand UO_3263 (O_3263,N_28769,N_28969);
nand UO_3264 (O_3264,N_28781,N_29961);
or UO_3265 (O_3265,N_29377,N_29786);
nand UO_3266 (O_3266,N_28623,N_29812);
or UO_3267 (O_3267,N_29953,N_29871);
xor UO_3268 (O_3268,N_28799,N_29220);
and UO_3269 (O_3269,N_28931,N_29528);
or UO_3270 (O_3270,N_29498,N_29798);
nand UO_3271 (O_3271,N_29223,N_28954);
nor UO_3272 (O_3272,N_28807,N_28933);
xnor UO_3273 (O_3273,N_29681,N_29836);
nand UO_3274 (O_3274,N_29443,N_28677);
or UO_3275 (O_3275,N_29687,N_29842);
nor UO_3276 (O_3276,N_28756,N_29821);
and UO_3277 (O_3277,N_29787,N_29341);
xor UO_3278 (O_3278,N_29313,N_29321);
and UO_3279 (O_3279,N_29165,N_29208);
or UO_3280 (O_3280,N_29200,N_29189);
and UO_3281 (O_3281,N_28967,N_29347);
or UO_3282 (O_3282,N_28532,N_28735);
nand UO_3283 (O_3283,N_28677,N_29700);
xor UO_3284 (O_3284,N_29999,N_28592);
nor UO_3285 (O_3285,N_29369,N_29981);
or UO_3286 (O_3286,N_29164,N_29733);
or UO_3287 (O_3287,N_28596,N_29896);
xnor UO_3288 (O_3288,N_28910,N_29704);
and UO_3289 (O_3289,N_28848,N_29828);
nor UO_3290 (O_3290,N_29765,N_29757);
nor UO_3291 (O_3291,N_29555,N_29407);
or UO_3292 (O_3292,N_28712,N_29788);
xnor UO_3293 (O_3293,N_29532,N_28832);
or UO_3294 (O_3294,N_28976,N_28561);
nor UO_3295 (O_3295,N_29123,N_29713);
or UO_3296 (O_3296,N_28932,N_29626);
nor UO_3297 (O_3297,N_29489,N_29980);
nand UO_3298 (O_3298,N_28897,N_29261);
nor UO_3299 (O_3299,N_28733,N_28718);
nor UO_3300 (O_3300,N_29967,N_29819);
or UO_3301 (O_3301,N_28557,N_28933);
nor UO_3302 (O_3302,N_28593,N_29186);
nand UO_3303 (O_3303,N_29853,N_28651);
and UO_3304 (O_3304,N_29725,N_29653);
nor UO_3305 (O_3305,N_29622,N_29346);
and UO_3306 (O_3306,N_29516,N_29481);
nor UO_3307 (O_3307,N_29473,N_29084);
xor UO_3308 (O_3308,N_28559,N_29868);
xnor UO_3309 (O_3309,N_28681,N_29143);
nor UO_3310 (O_3310,N_29378,N_29149);
or UO_3311 (O_3311,N_29537,N_29801);
nand UO_3312 (O_3312,N_28642,N_29470);
nor UO_3313 (O_3313,N_29477,N_29028);
nor UO_3314 (O_3314,N_28501,N_28811);
and UO_3315 (O_3315,N_29839,N_29183);
and UO_3316 (O_3316,N_28679,N_28899);
nor UO_3317 (O_3317,N_28560,N_29919);
xnor UO_3318 (O_3318,N_29612,N_29704);
xnor UO_3319 (O_3319,N_29014,N_29765);
and UO_3320 (O_3320,N_29030,N_28921);
or UO_3321 (O_3321,N_29168,N_29936);
nand UO_3322 (O_3322,N_29681,N_29241);
nand UO_3323 (O_3323,N_29953,N_28540);
and UO_3324 (O_3324,N_29823,N_29752);
and UO_3325 (O_3325,N_29142,N_29459);
nor UO_3326 (O_3326,N_28850,N_28667);
xnor UO_3327 (O_3327,N_29288,N_29247);
xnor UO_3328 (O_3328,N_28855,N_28579);
and UO_3329 (O_3329,N_29859,N_29483);
or UO_3330 (O_3330,N_29580,N_28581);
nand UO_3331 (O_3331,N_29203,N_29787);
nor UO_3332 (O_3332,N_29521,N_29836);
nand UO_3333 (O_3333,N_29650,N_29929);
or UO_3334 (O_3334,N_29875,N_28757);
and UO_3335 (O_3335,N_28556,N_29223);
and UO_3336 (O_3336,N_29896,N_28949);
and UO_3337 (O_3337,N_28572,N_29475);
nand UO_3338 (O_3338,N_29033,N_29541);
xor UO_3339 (O_3339,N_29540,N_29901);
and UO_3340 (O_3340,N_28927,N_28659);
xnor UO_3341 (O_3341,N_28962,N_29830);
xnor UO_3342 (O_3342,N_29020,N_28860);
nor UO_3343 (O_3343,N_29222,N_28763);
and UO_3344 (O_3344,N_29176,N_28657);
and UO_3345 (O_3345,N_29976,N_29845);
or UO_3346 (O_3346,N_29907,N_29317);
nor UO_3347 (O_3347,N_28892,N_29658);
xor UO_3348 (O_3348,N_29632,N_29708);
nor UO_3349 (O_3349,N_29335,N_29063);
xor UO_3350 (O_3350,N_29193,N_29569);
and UO_3351 (O_3351,N_28518,N_28951);
or UO_3352 (O_3352,N_29930,N_28738);
nor UO_3353 (O_3353,N_28855,N_29551);
and UO_3354 (O_3354,N_29554,N_29327);
nor UO_3355 (O_3355,N_29181,N_28690);
xor UO_3356 (O_3356,N_29590,N_29824);
or UO_3357 (O_3357,N_29681,N_29440);
nand UO_3358 (O_3358,N_29818,N_29582);
nand UO_3359 (O_3359,N_29036,N_29018);
xnor UO_3360 (O_3360,N_29141,N_28817);
nor UO_3361 (O_3361,N_29868,N_28847);
xnor UO_3362 (O_3362,N_28867,N_28608);
and UO_3363 (O_3363,N_29535,N_29918);
and UO_3364 (O_3364,N_28923,N_29197);
nand UO_3365 (O_3365,N_29798,N_29764);
nand UO_3366 (O_3366,N_29195,N_28851);
nor UO_3367 (O_3367,N_29347,N_29266);
or UO_3368 (O_3368,N_28892,N_28625);
nor UO_3369 (O_3369,N_28828,N_29725);
nand UO_3370 (O_3370,N_29998,N_29581);
nand UO_3371 (O_3371,N_29946,N_29234);
or UO_3372 (O_3372,N_29900,N_29670);
nand UO_3373 (O_3373,N_28658,N_29908);
xnor UO_3374 (O_3374,N_28802,N_29752);
nor UO_3375 (O_3375,N_28791,N_29361);
and UO_3376 (O_3376,N_29930,N_29273);
or UO_3377 (O_3377,N_29751,N_28867);
nor UO_3378 (O_3378,N_29214,N_28884);
xnor UO_3379 (O_3379,N_29460,N_29751);
nand UO_3380 (O_3380,N_29286,N_28683);
nor UO_3381 (O_3381,N_29307,N_29462);
xnor UO_3382 (O_3382,N_28720,N_28722);
or UO_3383 (O_3383,N_29574,N_29394);
or UO_3384 (O_3384,N_29243,N_29247);
nand UO_3385 (O_3385,N_29152,N_29213);
nand UO_3386 (O_3386,N_29471,N_29032);
or UO_3387 (O_3387,N_28682,N_29786);
xnor UO_3388 (O_3388,N_29070,N_29432);
and UO_3389 (O_3389,N_29077,N_28815);
and UO_3390 (O_3390,N_29315,N_29349);
or UO_3391 (O_3391,N_28888,N_29629);
and UO_3392 (O_3392,N_29969,N_29384);
nor UO_3393 (O_3393,N_29102,N_28556);
nor UO_3394 (O_3394,N_29973,N_29046);
or UO_3395 (O_3395,N_28904,N_28922);
or UO_3396 (O_3396,N_29795,N_28679);
nor UO_3397 (O_3397,N_28873,N_29501);
and UO_3398 (O_3398,N_28541,N_29580);
nand UO_3399 (O_3399,N_29559,N_29865);
nor UO_3400 (O_3400,N_29110,N_29150);
or UO_3401 (O_3401,N_28857,N_29737);
and UO_3402 (O_3402,N_29355,N_28612);
or UO_3403 (O_3403,N_28544,N_29589);
and UO_3404 (O_3404,N_29945,N_29924);
xor UO_3405 (O_3405,N_29779,N_29944);
nand UO_3406 (O_3406,N_29367,N_28765);
nor UO_3407 (O_3407,N_29070,N_29716);
xnor UO_3408 (O_3408,N_28509,N_29849);
nor UO_3409 (O_3409,N_28851,N_28959);
nor UO_3410 (O_3410,N_29553,N_29050);
nor UO_3411 (O_3411,N_29019,N_29997);
or UO_3412 (O_3412,N_29538,N_28905);
or UO_3413 (O_3413,N_29957,N_29437);
or UO_3414 (O_3414,N_29968,N_29987);
and UO_3415 (O_3415,N_28642,N_28899);
or UO_3416 (O_3416,N_28643,N_29684);
and UO_3417 (O_3417,N_29076,N_29461);
or UO_3418 (O_3418,N_28582,N_28761);
nand UO_3419 (O_3419,N_29150,N_28705);
xnor UO_3420 (O_3420,N_28809,N_29140);
nor UO_3421 (O_3421,N_29029,N_29848);
or UO_3422 (O_3422,N_29841,N_29996);
or UO_3423 (O_3423,N_29306,N_28808);
and UO_3424 (O_3424,N_28700,N_28858);
nor UO_3425 (O_3425,N_29608,N_29741);
xnor UO_3426 (O_3426,N_29013,N_29774);
and UO_3427 (O_3427,N_29383,N_29506);
nor UO_3428 (O_3428,N_29997,N_29572);
xnor UO_3429 (O_3429,N_29064,N_28944);
nand UO_3430 (O_3430,N_29928,N_29373);
nand UO_3431 (O_3431,N_28562,N_28857);
nor UO_3432 (O_3432,N_29392,N_28913);
and UO_3433 (O_3433,N_29776,N_28990);
and UO_3434 (O_3434,N_29869,N_29555);
nand UO_3435 (O_3435,N_28641,N_29074);
or UO_3436 (O_3436,N_29442,N_28948);
nor UO_3437 (O_3437,N_28663,N_29769);
nand UO_3438 (O_3438,N_29789,N_29889);
xor UO_3439 (O_3439,N_28616,N_28797);
xor UO_3440 (O_3440,N_29737,N_29630);
xnor UO_3441 (O_3441,N_29596,N_29307);
nand UO_3442 (O_3442,N_28529,N_28772);
xor UO_3443 (O_3443,N_29226,N_29242);
nor UO_3444 (O_3444,N_28651,N_29997);
and UO_3445 (O_3445,N_29774,N_28517);
nor UO_3446 (O_3446,N_29102,N_29458);
xnor UO_3447 (O_3447,N_28526,N_29456);
nor UO_3448 (O_3448,N_29749,N_29017);
xnor UO_3449 (O_3449,N_29485,N_29597);
nor UO_3450 (O_3450,N_28630,N_28661);
nand UO_3451 (O_3451,N_28508,N_29035);
or UO_3452 (O_3452,N_29907,N_28819);
or UO_3453 (O_3453,N_29409,N_28874);
or UO_3454 (O_3454,N_28735,N_28715);
and UO_3455 (O_3455,N_29017,N_29711);
xor UO_3456 (O_3456,N_28984,N_29690);
and UO_3457 (O_3457,N_29015,N_28555);
nand UO_3458 (O_3458,N_29502,N_29628);
nor UO_3459 (O_3459,N_29952,N_28506);
and UO_3460 (O_3460,N_29557,N_28972);
and UO_3461 (O_3461,N_29188,N_29003);
xor UO_3462 (O_3462,N_29265,N_29985);
nand UO_3463 (O_3463,N_29310,N_29590);
xor UO_3464 (O_3464,N_29394,N_29469);
nor UO_3465 (O_3465,N_29195,N_29136);
and UO_3466 (O_3466,N_28842,N_29472);
nor UO_3467 (O_3467,N_28579,N_28593);
xor UO_3468 (O_3468,N_29484,N_29669);
nand UO_3469 (O_3469,N_28722,N_28728);
nand UO_3470 (O_3470,N_29813,N_29708);
or UO_3471 (O_3471,N_28787,N_29311);
and UO_3472 (O_3472,N_29000,N_29402);
nor UO_3473 (O_3473,N_28537,N_29934);
or UO_3474 (O_3474,N_28705,N_28820);
xnor UO_3475 (O_3475,N_28770,N_29132);
or UO_3476 (O_3476,N_29688,N_28862);
nand UO_3477 (O_3477,N_29204,N_28829);
xnor UO_3478 (O_3478,N_29458,N_29680);
nor UO_3479 (O_3479,N_29254,N_29242);
xor UO_3480 (O_3480,N_29032,N_29488);
nand UO_3481 (O_3481,N_29014,N_29067);
nor UO_3482 (O_3482,N_28587,N_29517);
xor UO_3483 (O_3483,N_29243,N_29133);
xor UO_3484 (O_3484,N_29263,N_29530);
nor UO_3485 (O_3485,N_29064,N_28600);
xnor UO_3486 (O_3486,N_29474,N_29809);
or UO_3487 (O_3487,N_29572,N_29903);
and UO_3488 (O_3488,N_29600,N_29973);
nand UO_3489 (O_3489,N_28749,N_29210);
nor UO_3490 (O_3490,N_29619,N_29022);
and UO_3491 (O_3491,N_29899,N_28922);
xnor UO_3492 (O_3492,N_29373,N_29122);
nand UO_3493 (O_3493,N_29606,N_29135);
or UO_3494 (O_3494,N_28897,N_29879);
or UO_3495 (O_3495,N_29344,N_29819);
nand UO_3496 (O_3496,N_29609,N_29133);
and UO_3497 (O_3497,N_29849,N_29160);
and UO_3498 (O_3498,N_29133,N_28984);
nand UO_3499 (O_3499,N_28764,N_29692);
endmodule