module basic_500_3000_500_30_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_436,In_468);
nor U1 (N_1,In_236,In_452);
or U2 (N_2,In_247,In_217);
or U3 (N_3,In_259,In_199);
and U4 (N_4,In_284,In_22);
or U5 (N_5,In_435,In_234);
nand U6 (N_6,In_201,In_464);
nor U7 (N_7,In_7,In_386);
nor U8 (N_8,In_81,In_161);
or U9 (N_9,In_180,In_278);
nand U10 (N_10,In_208,In_343);
nor U11 (N_11,In_494,In_32);
nor U12 (N_12,In_258,In_159);
nand U13 (N_13,In_203,In_366);
and U14 (N_14,In_354,In_313);
nor U15 (N_15,In_391,In_415);
nor U16 (N_16,In_91,In_426);
and U17 (N_17,In_268,In_407);
and U18 (N_18,In_277,In_175);
and U19 (N_19,In_498,In_205);
nand U20 (N_20,In_177,In_427);
nand U21 (N_21,In_384,In_163);
nor U22 (N_22,In_10,In_342);
nand U23 (N_23,In_275,In_198);
and U24 (N_24,In_228,In_256);
and U25 (N_25,In_491,In_309);
and U26 (N_26,In_145,In_230);
and U27 (N_27,In_191,In_476);
or U28 (N_28,In_458,In_314);
or U29 (N_29,In_467,In_190);
and U30 (N_30,In_434,In_227);
nand U31 (N_31,In_385,In_167);
and U32 (N_32,In_403,In_94);
nand U33 (N_33,In_148,In_80);
nand U34 (N_34,In_388,In_14);
nand U35 (N_35,In_95,In_404);
nand U36 (N_36,In_33,In_419);
nand U37 (N_37,In_484,In_340);
nand U38 (N_38,In_413,In_67);
nor U39 (N_39,In_15,In_399);
and U40 (N_40,In_302,In_474);
xnor U41 (N_41,In_363,In_308);
and U42 (N_42,In_371,In_237);
and U43 (N_43,In_471,In_74);
nand U44 (N_44,In_357,In_6);
nand U45 (N_45,In_4,In_374);
or U46 (N_46,In_345,In_2);
nor U47 (N_47,In_486,In_96);
nor U48 (N_48,In_333,In_144);
nand U49 (N_49,In_331,In_249);
nand U50 (N_50,In_183,In_323);
or U51 (N_51,In_478,In_348);
and U52 (N_52,In_493,In_253);
nor U53 (N_53,In_410,In_315);
nand U54 (N_54,In_186,In_267);
nand U55 (N_55,In_117,In_54);
or U56 (N_56,In_383,In_179);
and U57 (N_57,In_396,In_143);
nand U58 (N_58,In_127,In_152);
nor U59 (N_59,In_335,In_424);
and U60 (N_60,In_176,In_84);
and U61 (N_61,In_245,In_35);
and U62 (N_62,In_114,In_64);
and U63 (N_63,In_111,In_166);
nor U64 (N_64,In_328,In_5);
or U65 (N_65,In_189,In_178);
nor U66 (N_66,In_206,In_330);
or U67 (N_67,In_241,In_25);
or U68 (N_68,In_125,In_266);
xnor U69 (N_69,In_27,In_450);
or U70 (N_70,In_104,In_57);
nor U71 (N_71,In_394,In_157);
nor U72 (N_72,In_16,In_400);
nor U73 (N_73,In_250,In_350);
and U74 (N_74,In_212,In_8);
or U75 (N_75,In_360,In_90);
nand U76 (N_76,In_246,In_115);
nand U77 (N_77,In_257,In_12);
nand U78 (N_78,In_233,In_221);
nand U79 (N_79,In_306,In_214);
xor U80 (N_80,In_172,In_365);
or U81 (N_81,In_232,In_136);
nor U82 (N_82,In_325,In_20);
and U83 (N_83,In_356,In_359);
nand U84 (N_84,In_171,In_310);
nor U85 (N_85,In_77,In_283);
and U86 (N_86,In_287,In_106);
or U87 (N_87,In_155,In_377);
or U88 (N_88,In_102,In_489);
nand U89 (N_89,In_76,In_289);
or U90 (N_90,In_272,In_222);
nor U91 (N_91,In_300,In_69);
and U92 (N_92,In_83,In_320);
and U93 (N_93,In_238,In_137);
and U94 (N_94,In_122,In_472);
nand U95 (N_95,In_274,In_279);
nor U96 (N_96,In_30,In_497);
or U97 (N_97,In_226,In_88);
or U98 (N_98,In_321,In_251);
and U99 (N_99,In_239,In_496);
nor U100 (N_100,In_454,N_59);
nor U101 (N_101,In_409,In_193);
nand U102 (N_102,N_34,In_26);
and U103 (N_103,N_2,In_92);
and U104 (N_104,N_19,In_291);
nor U105 (N_105,In_52,In_215);
or U106 (N_106,In_202,N_25);
or U107 (N_107,N_31,N_15);
nand U108 (N_108,In_499,In_75);
and U109 (N_109,In_466,In_139);
and U110 (N_110,In_301,In_105);
xor U111 (N_111,N_12,N_93);
nand U112 (N_112,In_142,In_68);
nor U113 (N_113,In_270,In_432);
or U114 (N_114,In_197,N_88);
or U115 (N_115,N_51,In_381);
and U116 (N_116,In_112,N_50);
and U117 (N_117,In_229,N_63);
or U118 (N_118,N_35,In_393);
and U119 (N_119,In_60,In_444);
or U120 (N_120,In_368,In_174);
or U121 (N_121,N_47,In_460);
or U122 (N_122,In_82,N_38);
nor U123 (N_123,In_101,In_446);
or U124 (N_124,N_89,N_57);
or U125 (N_125,In_73,In_131);
and U126 (N_126,In_319,N_28);
and U127 (N_127,In_107,N_74);
xor U128 (N_128,In_322,In_36);
nor U129 (N_129,In_378,In_477);
and U130 (N_130,In_406,In_329);
nor U131 (N_131,In_207,In_294);
or U132 (N_132,In_318,N_20);
nor U133 (N_133,In_341,N_42);
nor U134 (N_134,In_408,In_185);
or U135 (N_135,N_13,In_367);
xnor U136 (N_136,In_305,In_169);
or U137 (N_137,In_445,In_462);
nand U138 (N_138,N_79,In_37);
or U139 (N_139,N_77,N_48);
nand U140 (N_140,In_13,In_182);
nand U141 (N_141,In_431,N_94);
or U142 (N_142,In_344,In_100);
nor U143 (N_143,In_412,In_273);
xnor U144 (N_144,In_451,In_485);
and U145 (N_145,In_269,N_24);
nand U146 (N_146,In_120,In_240);
and U147 (N_147,In_418,In_128);
or U148 (N_148,N_65,In_126);
or U149 (N_149,In_17,N_16);
nand U150 (N_150,In_252,In_422);
and U151 (N_151,In_298,In_53);
and U152 (N_152,In_420,In_213);
or U153 (N_153,N_68,In_286);
xor U154 (N_154,In_153,N_80);
and U155 (N_155,N_83,In_150);
xor U156 (N_156,N_37,In_282);
nand U157 (N_157,In_395,In_181);
and U158 (N_158,N_92,In_254);
nand U159 (N_159,In_487,In_162);
nand U160 (N_160,N_23,In_71);
nor U161 (N_161,N_41,In_87);
and U162 (N_162,N_98,In_392);
nor U163 (N_163,N_61,In_43);
and U164 (N_164,In_483,In_447);
and U165 (N_165,In_479,In_370);
nand U166 (N_166,N_32,In_264);
xnor U167 (N_167,N_73,In_39);
nand U168 (N_168,In_297,N_11);
nand U169 (N_169,N_62,N_8);
or U170 (N_170,In_376,In_244);
nand U171 (N_171,N_95,N_97);
nand U172 (N_172,In_265,In_78);
xnor U173 (N_173,In_347,N_99);
or U174 (N_174,In_327,In_86);
xnor U175 (N_175,In_248,In_352);
nor U176 (N_176,In_132,In_98);
or U177 (N_177,In_387,In_380);
or U178 (N_178,In_56,N_96);
nor U179 (N_179,In_124,In_361);
nor U180 (N_180,In_324,In_443);
nor U181 (N_181,In_164,In_255);
and U182 (N_182,N_21,N_71);
nor U183 (N_183,In_147,In_192);
nand U184 (N_184,In_261,In_149);
nor U185 (N_185,In_337,In_24);
xor U186 (N_186,In_364,In_417);
nand U187 (N_187,In_349,In_303);
nand U188 (N_188,N_33,In_113);
xor U189 (N_189,N_66,In_47);
nor U190 (N_190,In_441,In_219);
nor U191 (N_191,N_75,N_0);
and U192 (N_192,N_56,N_49);
xnor U193 (N_193,In_482,In_61);
nor U194 (N_194,In_156,N_46);
or U195 (N_195,In_168,In_38);
or U196 (N_196,In_118,N_3);
xnor U197 (N_197,In_1,In_50);
or U198 (N_198,In_316,In_196);
and U199 (N_199,In_332,In_480);
and U200 (N_200,In_260,In_79);
nand U201 (N_201,N_170,In_45);
or U202 (N_202,In_421,N_101);
xnor U203 (N_203,N_6,In_293);
xnor U204 (N_204,In_495,In_51);
nand U205 (N_205,In_3,N_67);
and U206 (N_206,N_102,In_389);
or U207 (N_207,In_194,N_4);
nor U208 (N_208,N_54,N_147);
and U209 (N_209,N_185,In_373);
xnor U210 (N_210,N_193,N_164);
and U211 (N_211,In_416,In_290);
nor U212 (N_212,In_46,N_130);
nand U213 (N_213,N_159,N_69);
and U214 (N_214,N_137,N_168);
and U215 (N_215,N_58,N_161);
xnor U216 (N_216,N_121,In_351);
nor U217 (N_217,N_53,N_176);
or U218 (N_218,N_138,In_437);
nor U219 (N_219,In_41,In_429);
nor U220 (N_220,In_49,In_85);
nand U221 (N_221,N_14,N_105);
or U222 (N_222,N_103,N_17);
and U223 (N_223,In_141,In_281);
nor U224 (N_224,N_86,In_209);
or U225 (N_225,N_10,In_346);
nand U226 (N_226,In_242,N_119);
nand U227 (N_227,N_191,N_39);
nand U228 (N_228,In_42,In_138);
nor U229 (N_229,In_225,In_492);
or U230 (N_230,In_271,N_182);
nand U231 (N_231,N_160,N_120);
or U232 (N_232,In_72,N_29);
nor U233 (N_233,In_184,N_189);
nand U234 (N_234,N_135,N_196);
nand U235 (N_235,In_146,In_288);
nand U236 (N_236,N_115,N_108);
xnor U237 (N_237,N_43,In_438);
or U238 (N_238,In_430,N_36);
nor U239 (N_239,N_7,In_397);
nand U240 (N_240,N_30,In_488);
xnor U241 (N_241,N_167,In_449);
or U242 (N_242,N_124,N_148);
or U243 (N_243,In_173,In_481);
and U244 (N_244,In_470,N_144);
nand U245 (N_245,In_220,In_130);
nor U246 (N_246,In_243,In_490);
and U247 (N_247,In_299,In_204);
nor U248 (N_248,In_411,In_40);
nand U249 (N_249,In_58,In_292);
and U250 (N_250,In_218,N_186);
and U251 (N_251,In_440,N_169);
nor U252 (N_252,In_295,N_163);
or U253 (N_253,In_336,N_27);
and U254 (N_254,In_31,N_198);
nor U255 (N_255,In_338,In_457);
nor U256 (N_256,N_26,N_117);
nand U257 (N_257,In_461,In_103);
or U258 (N_258,N_143,In_475);
nor U259 (N_259,In_134,N_118);
and U260 (N_260,In_34,N_145);
nand U261 (N_261,In_160,In_119);
or U262 (N_262,N_190,N_178);
nor U263 (N_263,In_235,N_171);
nor U264 (N_264,N_188,In_262);
nor U265 (N_265,In_280,N_109);
and U266 (N_266,In_97,In_433);
xnor U267 (N_267,N_146,N_136);
xor U268 (N_268,N_1,N_76);
nand U269 (N_269,In_398,In_99);
xnor U270 (N_270,In_401,N_100);
and U271 (N_271,In_390,N_60);
or U272 (N_272,N_110,N_162);
and U273 (N_273,In_334,In_358);
nor U274 (N_274,In_44,N_140);
nor U275 (N_275,N_139,In_263);
nor U276 (N_276,N_9,In_109);
and U277 (N_277,In_369,N_111);
nor U278 (N_278,N_113,In_48);
and U279 (N_279,N_129,In_121);
nand U280 (N_280,N_165,In_425);
nand U281 (N_281,N_183,In_405);
and U282 (N_282,N_104,In_11);
and U283 (N_283,In_151,In_140);
or U284 (N_284,N_154,In_307);
xor U285 (N_285,N_40,In_339);
nand U286 (N_286,N_114,In_18);
and U287 (N_287,In_442,In_70);
nor U288 (N_288,In_428,In_414);
nor U289 (N_289,In_129,N_153);
nand U290 (N_290,N_116,In_224);
nand U291 (N_291,N_133,In_158);
or U292 (N_292,In_55,N_84);
or U293 (N_293,N_131,In_195);
nand U294 (N_294,In_62,N_184);
nand U295 (N_295,In_89,In_108);
nand U296 (N_296,In_93,In_187);
nand U297 (N_297,N_150,In_9);
nor U298 (N_298,In_448,In_135);
nand U299 (N_299,N_45,In_465);
nand U300 (N_300,N_90,N_226);
nor U301 (N_301,N_149,N_126);
nand U302 (N_302,N_158,In_123);
and U303 (N_303,N_174,N_205);
and U304 (N_304,N_268,N_112);
nor U305 (N_305,N_287,N_220);
xor U306 (N_306,N_230,N_81);
nor U307 (N_307,N_225,In_439);
and U308 (N_308,N_290,N_229);
and U309 (N_309,In_326,In_312);
or U310 (N_310,In_456,In_473);
nand U311 (N_311,N_213,In_116);
and U312 (N_312,N_85,N_125);
xor U313 (N_313,In_402,N_271);
or U314 (N_314,N_264,N_249);
nor U315 (N_315,N_283,N_238);
nor U316 (N_316,N_204,N_234);
and U317 (N_317,N_245,N_247);
or U318 (N_318,In_382,N_151);
nor U319 (N_319,N_18,N_277);
or U320 (N_320,N_228,In_28);
nor U321 (N_321,In_133,In_463);
nand U322 (N_322,N_207,N_199);
xnor U323 (N_323,N_107,N_127);
and U324 (N_324,N_261,N_260);
nor U325 (N_325,N_221,N_248);
or U326 (N_326,N_250,In_317);
xnor U327 (N_327,N_254,In_29);
or U328 (N_328,N_194,N_142);
nand U329 (N_329,In_423,N_232);
nand U330 (N_330,In_21,N_233);
nor U331 (N_331,N_217,N_273);
xnor U332 (N_332,In_379,In_65);
and U333 (N_333,N_202,N_258);
or U334 (N_334,N_180,N_224);
or U335 (N_335,N_289,N_253);
nor U336 (N_336,N_239,N_5);
and U337 (N_337,N_251,In_23);
nor U338 (N_338,N_270,N_235);
nor U339 (N_339,N_91,In_223);
nand U340 (N_340,N_192,N_288);
nand U341 (N_341,N_44,N_210);
and U342 (N_342,N_280,N_285);
nor U343 (N_343,N_297,N_215);
and U344 (N_344,N_175,N_22);
and U345 (N_345,N_179,In_355);
and U346 (N_346,N_243,In_165);
nand U347 (N_347,In_375,N_197);
nor U348 (N_348,In_66,N_298);
or U349 (N_349,N_240,In_296);
nand U350 (N_350,N_203,N_292);
xor U351 (N_351,N_172,N_155);
nand U352 (N_352,N_281,N_208);
or U353 (N_353,N_286,N_294);
or U354 (N_354,In_285,N_227);
or U355 (N_355,N_279,N_187);
nand U356 (N_356,N_284,N_252);
and U357 (N_357,N_269,N_70);
xnor U358 (N_358,N_128,N_141);
or U359 (N_359,In_231,N_293);
nand U360 (N_360,N_299,In_453);
nand U361 (N_361,In_276,N_55);
nor U362 (N_362,N_222,In_188);
nand U363 (N_363,N_218,In_362);
and U364 (N_364,In_210,N_266);
xor U365 (N_365,N_157,N_156);
nand U366 (N_366,N_209,N_259);
xor U367 (N_367,N_231,N_64);
nor U368 (N_368,In_455,N_274);
or U369 (N_369,In_372,In_63);
and U370 (N_370,N_152,N_257);
nor U371 (N_371,N_132,N_106);
nand U372 (N_372,N_122,In_459);
or U373 (N_373,In_170,N_216);
nand U374 (N_374,N_82,N_166);
nor U375 (N_375,In_19,N_177);
nor U376 (N_376,N_267,N_255);
nand U377 (N_377,In_0,N_282);
nor U378 (N_378,N_223,In_304);
or U379 (N_379,N_123,N_296);
and U380 (N_380,N_173,In_353);
xnor U381 (N_381,N_211,N_195);
nand U382 (N_382,N_242,N_52);
or U383 (N_383,In_469,N_244);
nor U384 (N_384,N_212,In_154);
nor U385 (N_385,N_200,N_256);
and U386 (N_386,N_295,N_246);
nor U387 (N_387,N_275,N_241);
or U388 (N_388,N_134,N_78);
nor U389 (N_389,N_262,N_206);
nor U390 (N_390,N_236,N_265);
or U391 (N_391,In_110,In_211);
or U392 (N_392,In_59,N_219);
xor U393 (N_393,N_291,N_181);
nor U394 (N_394,N_87,N_201);
or U395 (N_395,N_72,N_276);
nor U396 (N_396,N_214,In_200);
and U397 (N_397,N_263,N_272);
and U398 (N_398,In_216,In_311);
nor U399 (N_399,N_278,N_237);
nand U400 (N_400,N_380,N_335);
nand U401 (N_401,N_348,N_310);
nand U402 (N_402,N_399,N_395);
nand U403 (N_403,N_305,N_398);
nand U404 (N_404,N_315,N_336);
or U405 (N_405,N_381,N_387);
and U406 (N_406,N_379,N_321);
and U407 (N_407,N_372,N_303);
or U408 (N_408,N_370,N_312);
or U409 (N_409,N_374,N_316);
or U410 (N_410,N_361,N_328);
or U411 (N_411,N_389,N_349);
or U412 (N_412,N_377,N_344);
or U413 (N_413,N_388,N_325);
nor U414 (N_414,N_383,N_307);
and U415 (N_415,N_364,N_371);
nor U416 (N_416,N_326,N_347);
and U417 (N_417,N_350,N_331);
and U418 (N_418,N_324,N_369);
or U419 (N_419,N_355,N_309);
and U420 (N_420,N_365,N_356);
and U421 (N_421,N_373,N_366);
nand U422 (N_422,N_341,N_352);
or U423 (N_423,N_334,N_354);
and U424 (N_424,N_306,N_311);
or U425 (N_425,N_332,N_360);
or U426 (N_426,N_337,N_330);
nand U427 (N_427,N_319,N_339);
or U428 (N_428,N_357,N_394);
xnor U429 (N_429,N_368,N_327);
and U430 (N_430,N_391,N_323);
nand U431 (N_431,N_363,N_346);
and U432 (N_432,N_386,N_351);
nor U433 (N_433,N_313,N_362);
and U434 (N_434,N_358,N_397);
and U435 (N_435,N_340,N_320);
or U436 (N_436,N_375,N_382);
xor U437 (N_437,N_385,N_302);
or U438 (N_438,N_353,N_392);
and U439 (N_439,N_390,N_345);
xnor U440 (N_440,N_393,N_329);
nand U441 (N_441,N_338,N_378);
nand U442 (N_442,N_314,N_376);
and U443 (N_443,N_300,N_367);
nand U444 (N_444,N_359,N_396);
and U445 (N_445,N_342,N_308);
nor U446 (N_446,N_384,N_333);
and U447 (N_447,N_304,N_343);
or U448 (N_448,N_317,N_318);
or U449 (N_449,N_322,N_301);
nor U450 (N_450,N_398,N_326);
nor U451 (N_451,N_372,N_391);
nor U452 (N_452,N_379,N_328);
nor U453 (N_453,N_300,N_311);
or U454 (N_454,N_301,N_349);
or U455 (N_455,N_352,N_389);
or U456 (N_456,N_385,N_308);
or U457 (N_457,N_361,N_340);
nand U458 (N_458,N_350,N_393);
nand U459 (N_459,N_301,N_345);
xor U460 (N_460,N_393,N_330);
nor U461 (N_461,N_356,N_315);
xor U462 (N_462,N_339,N_309);
nand U463 (N_463,N_371,N_329);
nand U464 (N_464,N_372,N_304);
and U465 (N_465,N_397,N_307);
nor U466 (N_466,N_377,N_376);
or U467 (N_467,N_321,N_363);
and U468 (N_468,N_335,N_327);
or U469 (N_469,N_387,N_312);
nor U470 (N_470,N_377,N_354);
or U471 (N_471,N_317,N_323);
xor U472 (N_472,N_391,N_353);
nor U473 (N_473,N_353,N_345);
nor U474 (N_474,N_310,N_326);
nand U475 (N_475,N_323,N_367);
nor U476 (N_476,N_334,N_386);
xnor U477 (N_477,N_324,N_336);
nor U478 (N_478,N_328,N_302);
and U479 (N_479,N_311,N_368);
and U480 (N_480,N_390,N_398);
nor U481 (N_481,N_344,N_384);
or U482 (N_482,N_359,N_311);
and U483 (N_483,N_348,N_334);
nor U484 (N_484,N_385,N_311);
and U485 (N_485,N_363,N_311);
nor U486 (N_486,N_326,N_329);
nand U487 (N_487,N_323,N_346);
nor U488 (N_488,N_343,N_331);
and U489 (N_489,N_395,N_368);
nor U490 (N_490,N_309,N_352);
nand U491 (N_491,N_340,N_332);
nand U492 (N_492,N_328,N_381);
and U493 (N_493,N_381,N_317);
or U494 (N_494,N_365,N_351);
nor U495 (N_495,N_335,N_346);
and U496 (N_496,N_361,N_356);
nor U497 (N_497,N_310,N_328);
nand U498 (N_498,N_383,N_335);
xor U499 (N_499,N_348,N_309);
nand U500 (N_500,N_455,N_479);
or U501 (N_501,N_423,N_445);
nor U502 (N_502,N_452,N_412);
nand U503 (N_503,N_417,N_461);
and U504 (N_504,N_480,N_401);
nor U505 (N_505,N_442,N_408);
and U506 (N_506,N_487,N_473);
or U507 (N_507,N_447,N_419);
or U508 (N_508,N_486,N_464);
xnor U509 (N_509,N_409,N_482);
or U510 (N_510,N_474,N_407);
xnor U511 (N_511,N_457,N_415);
or U512 (N_512,N_427,N_490);
nor U513 (N_513,N_481,N_463);
and U514 (N_514,N_430,N_488);
nand U515 (N_515,N_448,N_456);
or U516 (N_516,N_436,N_429);
and U517 (N_517,N_469,N_485);
or U518 (N_518,N_446,N_439);
nor U519 (N_519,N_449,N_476);
nand U520 (N_520,N_450,N_424);
nor U521 (N_521,N_451,N_497);
and U522 (N_522,N_493,N_428);
or U523 (N_523,N_435,N_475);
or U524 (N_524,N_410,N_431);
nand U525 (N_525,N_468,N_472);
or U526 (N_526,N_416,N_413);
or U527 (N_527,N_492,N_420);
and U528 (N_528,N_499,N_438);
or U529 (N_529,N_494,N_400);
nor U530 (N_530,N_496,N_498);
or U531 (N_531,N_437,N_470);
nor U532 (N_532,N_460,N_402);
nand U533 (N_533,N_467,N_459);
nand U534 (N_534,N_421,N_477);
xnor U535 (N_535,N_454,N_483);
and U536 (N_536,N_462,N_406);
or U537 (N_537,N_489,N_440);
xnor U538 (N_538,N_495,N_418);
nand U539 (N_539,N_403,N_478);
and U540 (N_540,N_433,N_425);
or U541 (N_541,N_422,N_465);
or U542 (N_542,N_458,N_444);
or U543 (N_543,N_411,N_405);
nor U544 (N_544,N_484,N_471);
nand U545 (N_545,N_414,N_466);
xnor U546 (N_546,N_434,N_432);
and U547 (N_547,N_443,N_441);
or U548 (N_548,N_453,N_491);
nand U549 (N_549,N_426,N_404);
or U550 (N_550,N_479,N_476);
or U551 (N_551,N_465,N_402);
nor U552 (N_552,N_461,N_471);
and U553 (N_553,N_462,N_479);
or U554 (N_554,N_496,N_410);
or U555 (N_555,N_409,N_401);
nand U556 (N_556,N_490,N_444);
xor U557 (N_557,N_434,N_479);
or U558 (N_558,N_439,N_496);
and U559 (N_559,N_498,N_465);
nor U560 (N_560,N_479,N_486);
nor U561 (N_561,N_434,N_483);
xnor U562 (N_562,N_478,N_456);
or U563 (N_563,N_487,N_417);
and U564 (N_564,N_408,N_485);
or U565 (N_565,N_423,N_455);
nor U566 (N_566,N_466,N_483);
nand U567 (N_567,N_417,N_430);
xor U568 (N_568,N_455,N_482);
or U569 (N_569,N_446,N_485);
nand U570 (N_570,N_413,N_417);
xor U571 (N_571,N_474,N_406);
or U572 (N_572,N_433,N_438);
nor U573 (N_573,N_462,N_417);
nand U574 (N_574,N_413,N_469);
or U575 (N_575,N_429,N_451);
or U576 (N_576,N_419,N_492);
or U577 (N_577,N_480,N_421);
and U578 (N_578,N_423,N_474);
nor U579 (N_579,N_482,N_436);
nand U580 (N_580,N_406,N_439);
or U581 (N_581,N_436,N_464);
nor U582 (N_582,N_449,N_428);
nor U583 (N_583,N_483,N_479);
and U584 (N_584,N_466,N_456);
and U585 (N_585,N_462,N_495);
and U586 (N_586,N_439,N_490);
or U587 (N_587,N_499,N_432);
and U588 (N_588,N_498,N_403);
nand U589 (N_589,N_464,N_444);
xnor U590 (N_590,N_458,N_482);
nand U591 (N_591,N_441,N_428);
xor U592 (N_592,N_441,N_415);
or U593 (N_593,N_402,N_400);
nand U594 (N_594,N_446,N_450);
and U595 (N_595,N_459,N_432);
or U596 (N_596,N_482,N_424);
and U597 (N_597,N_462,N_473);
and U598 (N_598,N_480,N_469);
or U599 (N_599,N_490,N_475);
nand U600 (N_600,N_533,N_504);
or U601 (N_601,N_547,N_510);
nand U602 (N_602,N_546,N_560);
nor U603 (N_603,N_542,N_562);
or U604 (N_604,N_500,N_570);
nor U605 (N_605,N_543,N_555);
xnor U606 (N_606,N_569,N_590);
or U607 (N_607,N_535,N_579);
xnor U608 (N_608,N_518,N_589);
xor U609 (N_609,N_506,N_526);
or U610 (N_610,N_573,N_537);
nor U611 (N_611,N_519,N_580);
and U612 (N_612,N_557,N_565);
nor U613 (N_613,N_551,N_503);
xnor U614 (N_614,N_571,N_507);
and U615 (N_615,N_585,N_534);
and U616 (N_616,N_539,N_567);
and U617 (N_617,N_577,N_595);
or U618 (N_618,N_572,N_536);
or U619 (N_619,N_576,N_575);
nand U620 (N_620,N_561,N_550);
nand U621 (N_621,N_514,N_538);
and U622 (N_622,N_554,N_599);
and U623 (N_623,N_516,N_544);
nor U624 (N_624,N_588,N_568);
or U625 (N_625,N_566,N_552);
nand U626 (N_626,N_531,N_521);
nor U627 (N_627,N_517,N_564);
and U628 (N_628,N_593,N_524);
and U629 (N_629,N_591,N_505);
and U630 (N_630,N_582,N_556);
xor U631 (N_631,N_596,N_511);
nand U632 (N_632,N_549,N_501);
nor U633 (N_633,N_559,N_584);
or U634 (N_634,N_522,N_527);
nor U635 (N_635,N_586,N_515);
nor U636 (N_636,N_540,N_530);
and U637 (N_637,N_520,N_563);
nand U638 (N_638,N_558,N_594);
and U639 (N_639,N_523,N_574);
nand U640 (N_640,N_545,N_532);
nand U641 (N_641,N_597,N_528);
and U642 (N_642,N_541,N_509);
or U643 (N_643,N_502,N_583);
and U644 (N_644,N_512,N_513);
and U645 (N_645,N_578,N_581);
or U646 (N_646,N_508,N_592);
nor U647 (N_647,N_587,N_598);
or U648 (N_648,N_553,N_548);
nor U649 (N_649,N_525,N_529);
nand U650 (N_650,N_563,N_518);
nor U651 (N_651,N_591,N_598);
and U652 (N_652,N_530,N_599);
or U653 (N_653,N_533,N_517);
and U654 (N_654,N_513,N_561);
nor U655 (N_655,N_581,N_562);
nand U656 (N_656,N_579,N_531);
nand U657 (N_657,N_512,N_593);
or U658 (N_658,N_539,N_594);
xnor U659 (N_659,N_550,N_599);
or U660 (N_660,N_514,N_599);
nand U661 (N_661,N_559,N_503);
or U662 (N_662,N_502,N_576);
nor U663 (N_663,N_538,N_598);
or U664 (N_664,N_509,N_526);
or U665 (N_665,N_570,N_529);
nand U666 (N_666,N_524,N_522);
or U667 (N_667,N_585,N_569);
nor U668 (N_668,N_525,N_591);
and U669 (N_669,N_542,N_537);
xnor U670 (N_670,N_546,N_504);
or U671 (N_671,N_582,N_549);
and U672 (N_672,N_597,N_535);
nor U673 (N_673,N_523,N_581);
or U674 (N_674,N_590,N_534);
and U675 (N_675,N_591,N_515);
xnor U676 (N_676,N_543,N_509);
xor U677 (N_677,N_594,N_543);
xnor U678 (N_678,N_571,N_595);
nor U679 (N_679,N_537,N_511);
or U680 (N_680,N_515,N_574);
and U681 (N_681,N_551,N_528);
nand U682 (N_682,N_579,N_540);
nand U683 (N_683,N_577,N_563);
nor U684 (N_684,N_519,N_564);
nand U685 (N_685,N_577,N_565);
and U686 (N_686,N_570,N_503);
nor U687 (N_687,N_582,N_553);
nor U688 (N_688,N_542,N_561);
and U689 (N_689,N_503,N_592);
or U690 (N_690,N_515,N_521);
or U691 (N_691,N_516,N_578);
xor U692 (N_692,N_539,N_599);
or U693 (N_693,N_554,N_524);
or U694 (N_694,N_502,N_573);
and U695 (N_695,N_517,N_594);
xnor U696 (N_696,N_533,N_576);
xnor U697 (N_697,N_529,N_532);
nand U698 (N_698,N_569,N_586);
nand U699 (N_699,N_595,N_529);
or U700 (N_700,N_667,N_664);
or U701 (N_701,N_653,N_678);
xor U702 (N_702,N_616,N_636);
and U703 (N_703,N_668,N_686);
nand U704 (N_704,N_601,N_619);
nand U705 (N_705,N_639,N_621);
nor U706 (N_706,N_698,N_606);
and U707 (N_707,N_675,N_681);
or U708 (N_708,N_645,N_697);
and U709 (N_709,N_660,N_610);
or U710 (N_710,N_600,N_674);
nand U711 (N_711,N_632,N_617);
nand U712 (N_712,N_669,N_622);
or U713 (N_713,N_685,N_696);
nor U714 (N_714,N_623,N_680);
nand U715 (N_715,N_671,N_654);
xnor U716 (N_716,N_670,N_604);
or U717 (N_717,N_633,N_687);
nand U718 (N_718,N_673,N_620);
and U719 (N_719,N_627,N_672);
and U720 (N_720,N_689,N_666);
nand U721 (N_721,N_649,N_658);
nand U722 (N_722,N_650,N_661);
and U723 (N_723,N_634,N_613);
and U724 (N_724,N_607,N_642);
and U725 (N_725,N_676,N_637);
nand U726 (N_726,N_628,N_631);
nand U727 (N_727,N_605,N_682);
nor U728 (N_728,N_677,N_618);
nor U729 (N_729,N_693,N_630);
and U730 (N_730,N_626,N_603);
or U731 (N_731,N_657,N_641);
and U732 (N_732,N_611,N_694);
nand U733 (N_733,N_683,N_640);
and U734 (N_734,N_608,N_699);
nor U735 (N_735,N_692,N_656);
nor U736 (N_736,N_638,N_691);
or U737 (N_737,N_651,N_602);
or U738 (N_738,N_646,N_644);
xnor U739 (N_739,N_612,N_688);
or U740 (N_740,N_648,N_690);
or U741 (N_741,N_662,N_643);
and U742 (N_742,N_665,N_684);
nand U743 (N_743,N_624,N_659);
and U744 (N_744,N_655,N_625);
nor U745 (N_745,N_663,N_635);
or U746 (N_746,N_695,N_647);
and U747 (N_747,N_629,N_614);
xor U748 (N_748,N_609,N_615);
and U749 (N_749,N_652,N_679);
and U750 (N_750,N_638,N_631);
or U751 (N_751,N_688,N_651);
and U752 (N_752,N_640,N_690);
nor U753 (N_753,N_634,N_617);
and U754 (N_754,N_624,N_677);
xnor U755 (N_755,N_688,N_669);
xnor U756 (N_756,N_601,N_632);
or U757 (N_757,N_679,N_658);
or U758 (N_758,N_601,N_655);
xnor U759 (N_759,N_674,N_678);
or U760 (N_760,N_641,N_664);
nand U761 (N_761,N_603,N_637);
or U762 (N_762,N_602,N_605);
nand U763 (N_763,N_639,N_623);
nor U764 (N_764,N_683,N_633);
xnor U765 (N_765,N_603,N_688);
nand U766 (N_766,N_674,N_625);
or U767 (N_767,N_686,N_672);
or U768 (N_768,N_657,N_606);
xor U769 (N_769,N_638,N_667);
nor U770 (N_770,N_657,N_663);
nor U771 (N_771,N_652,N_615);
nand U772 (N_772,N_608,N_690);
nor U773 (N_773,N_629,N_697);
xnor U774 (N_774,N_689,N_691);
or U775 (N_775,N_662,N_692);
nor U776 (N_776,N_635,N_692);
nand U777 (N_777,N_633,N_648);
or U778 (N_778,N_639,N_641);
xnor U779 (N_779,N_626,N_617);
xnor U780 (N_780,N_673,N_629);
xor U781 (N_781,N_646,N_698);
nand U782 (N_782,N_678,N_692);
or U783 (N_783,N_627,N_649);
and U784 (N_784,N_697,N_670);
and U785 (N_785,N_681,N_649);
nor U786 (N_786,N_620,N_619);
nor U787 (N_787,N_631,N_660);
nor U788 (N_788,N_623,N_650);
and U789 (N_789,N_699,N_686);
or U790 (N_790,N_687,N_640);
nor U791 (N_791,N_611,N_658);
and U792 (N_792,N_650,N_636);
xor U793 (N_793,N_656,N_603);
or U794 (N_794,N_613,N_682);
xnor U795 (N_795,N_643,N_632);
nor U796 (N_796,N_647,N_606);
nand U797 (N_797,N_650,N_642);
nand U798 (N_798,N_610,N_602);
nand U799 (N_799,N_693,N_682);
nor U800 (N_800,N_775,N_766);
and U801 (N_801,N_794,N_721);
xor U802 (N_802,N_768,N_785);
and U803 (N_803,N_744,N_786);
nand U804 (N_804,N_787,N_734);
nor U805 (N_805,N_751,N_770);
and U806 (N_806,N_749,N_717);
nand U807 (N_807,N_756,N_716);
or U808 (N_808,N_752,N_740);
nor U809 (N_809,N_723,N_729);
nor U810 (N_810,N_760,N_780);
nand U811 (N_811,N_736,N_792);
or U812 (N_812,N_735,N_769);
nor U813 (N_813,N_789,N_754);
nand U814 (N_814,N_777,N_706);
nand U815 (N_815,N_759,N_725);
nand U816 (N_816,N_713,N_793);
or U817 (N_817,N_762,N_722);
nand U818 (N_818,N_747,N_748);
nand U819 (N_819,N_743,N_788);
or U820 (N_820,N_778,N_755);
nand U821 (N_821,N_764,N_703);
or U822 (N_822,N_799,N_745);
nor U823 (N_823,N_738,N_783);
nand U824 (N_824,N_776,N_705);
or U825 (N_825,N_746,N_704);
nor U826 (N_826,N_771,N_720);
or U827 (N_827,N_797,N_790);
or U828 (N_828,N_730,N_714);
nand U829 (N_829,N_750,N_758);
or U830 (N_830,N_795,N_781);
xor U831 (N_831,N_765,N_733);
nor U832 (N_832,N_737,N_772);
or U833 (N_833,N_767,N_761);
nor U834 (N_834,N_774,N_728);
nor U835 (N_835,N_798,N_702);
and U836 (N_836,N_726,N_791);
nand U837 (N_837,N_739,N_757);
nor U838 (N_838,N_712,N_701);
nor U839 (N_839,N_708,N_724);
or U840 (N_840,N_731,N_741);
nor U841 (N_841,N_784,N_782);
nand U842 (N_842,N_732,N_763);
and U843 (N_843,N_707,N_710);
xnor U844 (N_844,N_796,N_709);
nor U845 (N_845,N_715,N_773);
nor U846 (N_846,N_742,N_700);
nor U847 (N_847,N_719,N_753);
or U848 (N_848,N_779,N_711);
or U849 (N_849,N_718,N_727);
nand U850 (N_850,N_748,N_759);
or U851 (N_851,N_711,N_796);
or U852 (N_852,N_753,N_765);
nor U853 (N_853,N_700,N_768);
nor U854 (N_854,N_792,N_777);
or U855 (N_855,N_711,N_725);
or U856 (N_856,N_715,N_781);
or U857 (N_857,N_795,N_738);
nor U858 (N_858,N_793,N_717);
nand U859 (N_859,N_752,N_756);
or U860 (N_860,N_791,N_709);
nor U861 (N_861,N_731,N_716);
or U862 (N_862,N_799,N_758);
and U863 (N_863,N_788,N_725);
and U864 (N_864,N_732,N_762);
nor U865 (N_865,N_720,N_768);
nor U866 (N_866,N_705,N_760);
nor U867 (N_867,N_757,N_761);
and U868 (N_868,N_724,N_712);
nor U869 (N_869,N_711,N_733);
xnor U870 (N_870,N_762,N_789);
nor U871 (N_871,N_710,N_729);
xnor U872 (N_872,N_792,N_735);
and U873 (N_873,N_728,N_711);
nand U874 (N_874,N_782,N_748);
nand U875 (N_875,N_722,N_734);
nor U876 (N_876,N_708,N_768);
nor U877 (N_877,N_775,N_723);
xnor U878 (N_878,N_741,N_772);
nand U879 (N_879,N_748,N_725);
nand U880 (N_880,N_760,N_759);
nand U881 (N_881,N_714,N_704);
xnor U882 (N_882,N_779,N_770);
nand U883 (N_883,N_775,N_798);
nor U884 (N_884,N_778,N_751);
and U885 (N_885,N_769,N_774);
nand U886 (N_886,N_720,N_779);
nand U887 (N_887,N_737,N_712);
and U888 (N_888,N_755,N_737);
nand U889 (N_889,N_798,N_706);
nor U890 (N_890,N_709,N_736);
nand U891 (N_891,N_752,N_742);
and U892 (N_892,N_709,N_761);
nor U893 (N_893,N_722,N_761);
and U894 (N_894,N_705,N_726);
and U895 (N_895,N_723,N_735);
or U896 (N_896,N_788,N_763);
nor U897 (N_897,N_700,N_712);
or U898 (N_898,N_743,N_754);
nand U899 (N_899,N_739,N_730);
and U900 (N_900,N_874,N_807);
nor U901 (N_901,N_829,N_803);
nand U902 (N_902,N_815,N_865);
and U903 (N_903,N_859,N_891);
or U904 (N_904,N_858,N_845);
and U905 (N_905,N_894,N_863);
nand U906 (N_906,N_840,N_866);
and U907 (N_907,N_820,N_827);
or U908 (N_908,N_818,N_879);
and U909 (N_909,N_875,N_881);
and U910 (N_910,N_855,N_837);
nand U911 (N_911,N_842,N_887);
and U912 (N_912,N_850,N_852);
nor U913 (N_913,N_817,N_832);
or U914 (N_914,N_888,N_847);
and U915 (N_915,N_825,N_839);
xor U916 (N_916,N_857,N_802);
nand U917 (N_917,N_836,N_890);
nor U918 (N_918,N_819,N_862);
and U919 (N_919,N_899,N_892);
nand U920 (N_920,N_877,N_868);
nand U921 (N_921,N_872,N_876);
and U922 (N_922,N_816,N_864);
and U923 (N_923,N_885,N_860);
nand U924 (N_924,N_886,N_898);
nand U925 (N_925,N_800,N_856);
xnor U926 (N_926,N_804,N_897);
or U927 (N_927,N_844,N_853);
nand U928 (N_928,N_851,N_896);
nor U929 (N_929,N_846,N_806);
nor U930 (N_930,N_895,N_828);
and U931 (N_931,N_811,N_883);
nand U932 (N_932,N_809,N_884);
nand U933 (N_933,N_830,N_805);
nor U934 (N_934,N_821,N_882);
nand U935 (N_935,N_824,N_843);
nor U936 (N_936,N_810,N_869);
nand U937 (N_937,N_831,N_834);
nand U938 (N_938,N_848,N_822);
nand U939 (N_939,N_814,N_871);
xnor U940 (N_940,N_812,N_854);
and U941 (N_941,N_823,N_889);
nor U942 (N_942,N_813,N_841);
nand U943 (N_943,N_870,N_833);
nand U944 (N_944,N_808,N_849);
nand U945 (N_945,N_893,N_873);
or U946 (N_946,N_838,N_801);
and U947 (N_947,N_880,N_835);
nor U948 (N_948,N_826,N_861);
or U949 (N_949,N_867,N_878);
nor U950 (N_950,N_873,N_802);
nand U951 (N_951,N_855,N_830);
or U952 (N_952,N_864,N_815);
nand U953 (N_953,N_880,N_884);
or U954 (N_954,N_855,N_899);
nand U955 (N_955,N_861,N_801);
and U956 (N_956,N_878,N_819);
or U957 (N_957,N_838,N_844);
and U958 (N_958,N_886,N_843);
or U959 (N_959,N_838,N_825);
or U960 (N_960,N_864,N_896);
and U961 (N_961,N_851,N_813);
nor U962 (N_962,N_883,N_881);
xor U963 (N_963,N_887,N_891);
nor U964 (N_964,N_806,N_813);
nand U965 (N_965,N_852,N_897);
xnor U966 (N_966,N_891,N_850);
nand U967 (N_967,N_857,N_895);
xor U968 (N_968,N_890,N_852);
and U969 (N_969,N_814,N_837);
nand U970 (N_970,N_813,N_848);
nand U971 (N_971,N_829,N_840);
nand U972 (N_972,N_811,N_861);
nor U973 (N_973,N_866,N_883);
nand U974 (N_974,N_866,N_881);
and U975 (N_975,N_876,N_854);
and U976 (N_976,N_898,N_862);
nand U977 (N_977,N_862,N_899);
and U978 (N_978,N_833,N_869);
xor U979 (N_979,N_843,N_894);
and U980 (N_980,N_895,N_813);
nand U981 (N_981,N_883,N_887);
and U982 (N_982,N_874,N_858);
or U983 (N_983,N_849,N_800);
and U984 (N_984,N_867,N_879);
and U985 (N_985,N_847,N_880);
nor U986 (N_986,N_889,N_840);
nand U987 (N_987,N_806,N_811);
or U988 (N_988,N_864,N_823);
nand U989 (N_989,N_869,N_853);
and U990 (N_990,N_885,N_804);
or U991 (N_991,N_869,N_819);
and U992 (N_992,N_858,N_866);
nand U993 (N_993,N_865,N_825);
or U994 (N_994,N_864,N_801);
and U995 (N_995,N_806,N_879);
nand U996 (N_996,N_821,N_829);
or U997 (N_997,N_805,N_836);
or U998 (N_998,N_870,N_827);
nand U999 (N_999,N_828,N_809);
nand U1000 (N_1000,N_970,N_995);
or U1001 (N_1001,N_997,N_920);
nor U1002 (N_1002,N_934,N_912);
or U1003 (N_1003,N_992,N_948);
nand U1004 (N_1004,N_956,N_936);
nor U1005 (N_1005,N_908,N_923);
xor U1006 (N_1006,N_949,N_961);
or U1007 (N_1007,N_944,N_921);
nor U1008 (N_1008,N_933,N_993);
or U1009 (N_1009,N_957,N_979);
nand U1010 (N_1010,N_951,N_931);
and U1011 (N_1011,N_969,N_975);
and U1012 (N_1012,N_950,N_930);
xnor U1013 (N_1013,N_935,N_916);
and U1014 (N_1014,N_966,N_945);
and U1015 (N_1015,N_953,N_985);
nand U1016 (N_1016,N_977,N_980);
nor U1017 (N_1017,N_976,N_938);
and U1018 (N_1018,N_971,N_947);
nor U1019 (N_1019,N_918,N_915);
or U1020 (N_1020,N_974,N_932);
nor U1021 (N_1021,N_942,N_958);
nand U1022 (N_1022,N_954,N_994);
or U1023 (N_1023,N_987,N_968);
nand U1024 (N_1024,N_909,N_982);
and U1025 (N_1025,N_991,N_913);
xnor U1026 (N_1026,N_999,N_941);
and U1027 (N_1027,N_911,N_960);
and U1028 (N_1028,N_907,N_972);
nand U1029 (N_1029,N_925,N_996);
or U1030 (N_1030,N_955,N_900);
or U1031 (N_1031,N_910,N_940);
xnor U1032 (N_1032,N_978,N_919);
nand U1033 (N_1033,N_990,N_981);
and U1034 (N_1034,N_904,N_924);
or U1035 (N_1035,N_901,N_903);
xnor U1036 (N_1036,N_905,N_998);
xnor U1037 (N_1037,N_952,N_917);
xnor U1038 (N_1038,N_986,N_927);
xor U1039 (N_1039,N_964,N_963);
nor U1040 (N_1040,N_962,N_939);
or U1041 (N_1041,N_914,N_973);
xnor U1042 (N_1042,N_965,N_906);
nor U1043 (N_1043,N_926,N_922);
or U1044 (N_1044,N_988,N_984);
nor U1045 (N_1045,N_937,N_967);
xor U1046 (N_1046,N_928,N_902);
xnor U1047 (N_1047,N_983,N_946);
nor U1048 (N_1048,N_929,N_989);
nand U1049 (N_1049,N_959,N_943);
and U1050 (N_1050,N_937,N_935);
and U1051 (N_1051,N_917,N_909);
and U1052 (N_1052,N_950,N_989);
nand U1053 (N_1053,N_996,N_979);
or U1054 (N_1054,N_971,N_978);
xnor U1055 (N_1055,N_942,N_906);
or U1056 (N_1056,N_998,N_910);
nand U1057 (N_1057,N_938,N_923);
nor U1058 (N_1058,N_933,N_999);
or U1059 (N_1059,N_919,N_942);
nand U1060 (N_1060,N_939,N_966);
nor U1061 (N_1061,N_993,N_947);
or U1062 (N_1062,N_925,N_902);
nor U1063 (N_1063,N_918,N_910);
or U1064 (N_1064,N_975,N_945);
or U1065 (N_1065,N_987,N_940);
or U1066 (N_1066,N_977,N_949);
and U1067 (N_1067,N_940,N_950);
nor U1068 (N_1068,N_994,N_988);
or U1069 (N_1069,N_919,N_953);
and U1070 (N_1070,N_926,N_943);
xnor U1071 (N_1071,N_956,N_941);
nand U1072 (N_1072,N_913,N_932);
or U1073 (N_1073,N_956,N_915);
nor U1074 (N_1074,N_963,N_999);
or U1075 (N_1075,N_901,N_960);
xnor U1076 (N_1076,N_952,N_971);
nor U1077 (N_1077,N_996,N_931);
and U1078 (N_1078,N_914,N_987);
and U1079 (N_1079,N_904,N_986);
nand U1080 (N_1080,N_919,N_971);
nand U1081 (N_1081,N_965,N_998);
and U1082 (N_1082,N_985,N_989);
and U1083 (N_1083,N_950,N_984);
nor U1084 (N_1084,N_995,N_938);
nand U1085 (N_1085,N_970,N_987);
or U1086 (N_1086,N_906,N_979);
nand U1087 (N_1087,N_932,N_920);
xnor U1088 (N_1088,N_960,N_923);
or U1089 (N_1089,N_948,N_911);
and U1090 (N_1090,N_980,N_962);
or U1091 (N_1091,N_927,N_980);
or U1092 (N_1092,N_994,N_993);
nand U1093 (N_1093,N_923,N_917);
xnor U1094 (N_1094,N_960,N_952);
and U1095 (N_1095,N_947,N_939);
xnor U1096 (N_1096,N_909,N_986);
nor U1097 (N_1097,N_913,N_965);
xor U1098 (N_1098,N_992,N_958);
nor U1099 (N_1099,N_967,N_932);
nor U1100 (N_1100,N_1020,N_1049);
and U1101 (N_1101,N_1096,N_1073);
and U1102 (N_1102,N_1068,N_1043);
nor U1103 (N_1103,N_1084,N_1009);
nand U1104 (N_1104,N_1010,N_1003);
or U1105 (N_1105,N_1026,N_1023);
nand U1106 (N_1106,N_1051,N_1055);
nand U1107 (N_1107,N_1045,N_1041);
xor U1108 (N_1108,N_1065,N_1044);
nand U1109 (N_1109,N_1088,N_1025);
nor U1110 (N_1110,N_1001,N_1091);
nor U1111 (N_1111,N_1040,N_1004);
nor U1112 (N_1112,N_1069,N_1059);
nand U1113 (N_1113,N_1075,N_1000);
xor U1114 (N_1114,N_1082,N_1080);
nand U1115 (N_1115,N_1032,N_1047);
and U1116 (N_1116,N_1095,N_1076);
nand U1117 (N_1117,N_1031,N_1024);
nor U1118 (N_1118,N_1067,N_1021);
and U1119 (N_1119,N_1036,N_1070);
or U1120 (N_1120,N_1083,N_1050);
xnor U1121 (N_1121,N_1077,N_1099);
nor U1122 (N_1122,N_1092,N_1046);
nand U1123 (N_1123,N_1060,N_1028);
and U1124 (N_1124,N_1094,N_1017);
and U1125 (N_1125,N_1062,N_1042);
xnor U1126 (N_1126,N_1011,N_1007);
nor U1127 (N_1127,N_1034,N_1014);
nor U1128 (N_1128,N_1012,N_1029);
nor U1129 (N_1129,N_1058,N_1086);
nor U1130 (N_1130,N_1027,N_1035);
nand U1131 (N_1131,N_1089,N_1087);
and U1132 (N_1132,N_1006,N_1090);
or U1133 (N_1133,N_1078,N_1097);
xnor U1134 (N_1134,N_1085,N_1033);
and U1135 (N_1135,N_1074,N_1019);
nor U1136 (N_1136,N_1022,N_1053);
xnor U1137 (N_1137,N_1054,N_1016);
nor U1138 (N_1138,N_1037,N_1063);
and U1139 (N_1139,N_1008,N_1005);
or U1140 (N_1140,N_1038,N_1052);
nand U1141 (N_1141,N_1002,N_1048);
or U1142 (N_1142,N_1061,N_1015);
and U1143 (N_1143,N_1081,N_1056);
xor U1144 (N_1144,N_1030,N_1072);
and U1145 (N_1145,N_1098,N_1039);
nor U1146 (N_1146,N_1093,N_1079);
nor U1147 (N_1147,N_1071,N_1018);
nand U1148 (N_1148,N_1013,N_1066);
or U1149 (N_1149,N_1064,N_1057);
and U1150 (N_1150,N_1003,N_1094);
and U1151 (N_1151,N_1052,N_1029);
nand U1152 (N_1152,N_1065,N_1057);
or U1153 (N_1153,N_1015,N_1044);
or U1154 (N_1154,N_1073,N_1055);
nand U1155 (N_1155,N_1019,N_1021);
and U1156 (N_1156,N_1076,N_1018);
xor U1157 (N_1157,N_1097,N_1017);
nor U1158 (N_1158,N_1086,N_1081);
nor U1159 (N_1159,N_1090,N_1012);
nand U1160 (N_1160,N_1083,N_1026);
xnor U1161 (N_1161,N_1029,N_1077);
nor U1162 (N_1162,N_1024,N_1038);
nand U1163 (N_1163,N_1026,N_1093);
or U1164 (N_1164,N_1048,N_1037);
nor U1165 (N_1165,N_1011,N_1047);
and U1166 (N_1166,N_1045,N_1046);
and U1167 (N_1167,N_1011,N_1071);
nand U1168 (N_1168,N_1041,N_1051);
and U1169 (N_1169,N_1013,N_1024);
xnor U1170 (N_1170,N_1049,N_1015);
nor U1171 (N_1171,N_1046,N_1051);
nor U1172 (N_1172,N_1040,N_1045);
and U1173 (N_1173,N_1022,N_1043);
nand U1174 (N_1174,N_1063,N_1075);
nand U1175 (N_1175,N_1040,N_1094);
and U1176 (N_1176,N_1003,N_1005);
nand U1177 (N_1177,N_1043,N_1024);
nand U1178 (N_1178,N_1059,N_1018);
and U1179 (N_1179,N_1000,N_1010);
nand U1180 (N_1180,N_1014,N_1023);
or U1181 (N_1181,N_1042,N_1074);
nand U1182 (N_1182,N_1019,N_1098);
nand U1183 (N_1183,N_1085,N_1086);
or U1184 (N_1184,N_1098,N_1067);
nor U1185 (N_1185,N_1081,N_1039);
or U1186 (N_1186,N_1006,N_1075);
and U1187 (N_1187,N_1068,N_1094);
or U1188 (N_1188,N_1089,N_1009);
or U1189 (N_1189,N_1025,N_1089);
nor U1190 (N_1190,N_1017,N_1002);
nand U1191 (N_1191,N_1026,N_1046);
nand U1192 (N_1192,N_1098,N_1027);
nand U1193 (N_1193,N_1067,N_1053);
nor U1194 (N_1194,N_1001,N_1088);
xnor U1195 (N_1195,N_1051,N_1010);
nand U1196 (N_1196,N_1089,N_1070);
nand U1197 (N_1197,N_1068,N_1071);
or U1198 (N_1198,N_1003,N_1096);
or U1199 (N_1199,N_1039,N_1067);
nand U1200 (N_1200,N_1142,N_1137);
or U1201 (N_1201,N_1154,N_1130);
nand U1202 (N_1202,N_1149,N_1136);
nand U1203 (N_1203,N_1148,N_1197);
nand U1204 (N_1204,N_1157,N_1170);
xor U1205 (N_1205,N_1163,N_1172);
nand U1206 (N_1206,N_1160,N_1164);
and U1207 (N_1207,N_1169,N_1111);
nand U1208 (N_1208,N_1113,N_1127);
nor U1209 (N_1209,N_1139,N_1117);
nor U1210 (N_1210,N_1159,N_1176);
nand U1211 (N_1211,N_1181,N_1193);
and U1212 (N_1212,N_1116,N_1146);
and U1213 (N_1213,N_1175,N_1186);
and U1214 (N_1214,N_1112,N_1135);
nand U1215 (N_1215,N_1198,N_1119);
or U1216 (N_1216,N_1162,N_1124);
nor U1217 (N_1217,N_1104,N_1153);
or U1218 (N_1218,N_1188,N_1141);
nor U1219 (N_1219,N_1121,N_1144);
and U1220 (N_1220,N_1174,N_1182);
nor U1221 (N_1221,N_1147,N_1133);
nand U1222 (N_1222,N_1109,N_1118);
and U1223 (N_1223,N_1134,N_1190);
nand U1224 (N_1224,N_1199,N_1131);
nor U1225 (N_1225,N_1122,N_1140);
nor U1226 (N_1226,N_1179,N_1177);
nor U1227 (N_1227,N_1107,N_1115);
and U1228 (N_1228,N_1105,N_1100);
or U1229 (N_1229,N_1156,N_1103);
or U1230 (N_1230,N_1167,N_1123);
nor U1231 (N_1231,N_1168,N_1180);
nor U1232 (N_1232,N_1155,N_1158);
nand U1233 (N_1233,N_1194,N_1138);
and U1234 (N_1234,N_1128,N_1145);
or U1235 (N_1235,N_1192,N_1152);
or U1236 (N_1236,N_1184,N_1178);
or U1237 (N_1237,N_1102,N_1129);
or U1238 (N_1238,N_1165,N_1196);
nand U1239 (N_1239,N_1183,N_1166);
or U1240 (N_1240,N_1161,N_1173);
nor U1241 (N_1241,N_1126,N_1108);
nand U1242 (N_1242,N_1120,N_1191);
nand U1243 (N_1243,N_1125,N_1151);
and U1244 (N_1244,N_1150,N_1106);
xnor U1245 (N_1245,N_1185,N_1114);
or U1246 (N_1246,N_1187,N_1101);
and U1247 (N_1247,N_1195,N_1171);
and U1248 (N_1248,N_1189,N_1143);
nor U1249 (N_1249,N_1110,N_1132);
nand U1250 (N_1250,N_1196,N_1189);
or U1251 (N_1251,N_1177,N_1109);
xor U1252 (N_1252,N_1101,N_1141);
or U1253 (N_1253,N_1122,N_1172);
nor U1254 (N_1254,N_1191,N_1155);
nand U1255 (N_1255,N_1186,N_1106);
nand U1256 (N_1256,N_1130,N_1121);
and U1257 (N_1257,N_1171,N_1149);
and U1258 (N_1258,N_1123,N_1161);
and U1259 (N_1259,N_1140,N_1181);
and U1260 (N_1260,N_1160,N_1171);
or U1261 (N_1261,N_1151,N_1123);
and U1262 (N_1262,N_1177,N_1187);
and U1263 (N_1263,N_1109,N_1124);
nor U1264 (N_1264,N_1118,N_1149);
xnor U1265 (N_1265,N_1194,N_1191);
or U1266 (N_1266,N_1112,N_1127);
and U1267 (N_1267,N_1100,N_1113);
xnor U1268 (N_1268,N_1129,N_1136);
or U1269 (N_1269,N_1102,N_1190);
nand U1270 (N_1270,N_1168,N_1157);
nor U1271 (N_1271,N_1171,N_1111);
and U1272 (N_1272,N_1113,N_1199);
and U1273 (N_1273,N_1191,N_1160);
and U1274 (N_1274,N_1190,N_1165);
nor U1275 (N_1275,N_1146,N_1175);
or U1276 (N_1276,N_1113,N_1138);
nor U1277 (N_1277,N_1116,N_1101);
nand U1278 (N_1278,N_1155,N_1104);
or U1279 (N_1279,N_1101,N_1107);
or U1280 (N_1280,N_1174,N_1118);
or U1281 (N_1281,N_1175,N_1185);
and U1282 (N_1282,N_1156,N_1171);
nand U1283 (N_1283,N_1196,N_1172);
nand U1284 (N_1284,N_1154,N_1165);
or U1285 (N_1285,N_1111,N_1186);
or U1286 (N_1286,N_1174,N_1172);
nand U1287 (N_1287,N_1119,N_1177);
xnor U1288 (N_1288,N_1104,N_1177);
xnor U1289 (N_1289,N_1133,N_1143);
nor U1290 (N_1290,N_1110,N_1179);
nor U1291 (N_1291,N_1162,N_1160);
nand U1292 (N_1292,N_1105,N_1139);
nand U1293 (N_1293,N_1112,N_1167);
nor U1294 (N_1294,N_1174,N_1163);
or U1295 (N_1295,N_1199,N_1177);
or U1296 (N_1296,N_1160,N_1194);
xnor U1297 (N_1297,N_1157,N_1151);
and U1298 (N_1298,N_1173,N_1142);
nand U1299 (N_1299,N_1178,N_1103);
or U1300 (N_1300,N_1242,N_1235);
nand U1301 (N_1301,N_1246,N_1263);
nand U1302 (N_1302,N_1277,N_1247);
or U1303 (N_1303,N_1221,N_1282);
or U1304 (N_1304,N_1290,N_1202);
nand U1305 (N_1305,N_1206,N_1233);
nand U1306 (N_1306,N_1201,N_1257);
xor U1307 (N_1307,N_1266,N_1225);
nand U1308 (N_1308,N_1248,N_1244);
nor U1309 (N_1309,N_1265,N_1214);
nand U1310 (N_1310,N_1258,N_1203);
nor U1311 (N_1311,N_1292,N_1228);
and U1312 (N_1312,N_1216,N_1276);
and U1313 (N_1313,N_1283,N_1281);
nor U1314 (N_1314,N_1284,N_1234);
and U1315 (N_1315,N_1294,N_1252);
or U1316 (N_1316,N_1270,N_1241);
and U1317 (N_1317,N_1256,N_1259);
or U1318 (N_1318,N_1213,N_1279);
and U1319 (N_1319,N_1223,N_1238);
and U1320 (N_1320,N_1211,N_1229);
and U1321 (N_1321,N_1271,N_1226);
xor U1322 (N_1322,N_1296,N_1204);
xor U1323 (N_1323,N_1245,N_1222);
xnor U1324 (N_1324,N_1289,N_1207);
and U1325 (N_1325,N_1208,N_1236);
and U1326 (N_1326,N_1269,N_1274);
and U1327 (N_1327,N_1215,N_1219);
nand U1328 (N_1328,N_1237,N_1231);
nand U1329 (N_1329,N_1285,N_1268);
xor U1330 (N_1330,N_1261,N_1288);
and U1331 (N_1331,N_1278,N_1249);
nor U1332 (N_1332,N_1232,N_1267);
nand U1333 (N_1333,N_1286,N_1220);
nor U1334 (N_1334,N_1240,N_1293);
nand U1335 (N_1335,N_1200,N_1253);
xor U1336 (N_1336,N_1239,N_1297);
and U1337 (N_1337,N_1218,N_1260);
nand U1338 (N_1338,N_1262,N_1250);
nand U1339 (N_1339,N_1217,N_1212);
nor U1340 (N_1340,N_1272,N_1243);
nor U1341 (N_1341,N_1230,N_1287);
nand U1342 (N_1342,N_1227,N_1280);
nor U1343 (N_1343,N_1275,N_1255);
or U1344 (N_1344,N_1299,N_1264);
and U1345 (N_1345,N_1224,N_1273);
and U1346 (N_1346,N_1210,N_1251);
nor U1347 (N_1347,N_1205,N_1209);
or U1348 (N_1348,N_1291,N_1295);
nand U1349 (N_1349,N_1298,N_1254);
and U1350 (N_1350,N_1262,N_1265);
nor U1351 (N_1351,N_1233,N_1240);
and U1352 (N_1352,N_1244,N_1243);
or U1353 (N_1353,N_1249,N_1281);
nand U1354 (N_1354,N_1205,N_1262);
and U1355 (N_1355,N_1254,N_1282);
and U1356 (N_1356,N_1238,N_1208);
or U1357 (N_1357,N_1277,N_1222);
or U1358 (N_1358,N_1276,N_1262);
nor U1359 (N_1359,N_1272,N_1202);
and U1360 (N_1360,N_1295,N_1294);
nor U1361 (N_1361,N_1201,N_1241);
or U1362 (N_1362,N_1292,N_1266);
or U1363 (N_1363,N_1210,N_1295);
nand U1364 (N_1364,N_1291,N_1212);
and U1365 (N_1365,N_1208,N_1283);
nor U1366 (N_1366,N_1290,N_1226);
and U1367 (N_1367,N_1233,N_1215);
nor U1368 (N_1368,N_1251,N_1258);
xnor U1369 (N_1369,N_1240,N_1210);
or U1370 (N_1370,N_1246,N_1289);
and U1371 (N_1371,N_1200,N_1246);
or U1372 (N_1372,N_1234,N_1244);
nand U1373 (N_1373,N_1274,N_1201);
or U1374 (N_1374,N_1205,N_1258);
or U1375 (N_1375,N_1294,N_1285);
and U1376 (N_1376,N_1224,N_1237);
nand U1377 (N_1377,N_1288,N_1255);
and U1378 (N_1378,N_1262,N_1267);
nand U1379 (N_1379,N_1256,N_1297);
and U1380 (N_1380,N_1241,N_1242);
xnor U1381 (N_1381,N_1259,N_1243);
nor U1382 (N_1382,N_1221,N_1238);
nor U1383 (N_1383,N_1255,N_1287);
and U1384 (N_1384,N_1234,N_1263);
nand U1385 (N_1385,N_1267,N_1268);
and U1386 (N_1386,N_1215,N_1251);
or U1387 (N_1387,N_1268,N_1205);
and U1388 (N_1388,N_1220,N_1273);
or U1389 (N_1389,N_1292,N_1250);
nor U1390 (N_1390,N_1280,N_1251);
nor U1391 (N_1391,N_1270,N_1208);
and U1392 (N_1392,N_1255,N_1254);
nand U1393 (N_1393,N_1289,N_1229);
nand U1394 (N_1394,N_1299,N_1213);
nand U1395 (N_1395,N_1294,N_1205);
and U1396 (N_1396,N_1230,N_1233);
or U1397 (N_1397,N_1255,N_1240);
nor U1398 (N_1398,N_1233,N_1232);
nor U1399 (N_1399,N_1225,N_1203);
and U1400 (N_1400,N_1398,N_1364);
nor U1401 (N_1401,N_1304,N_1320);
nor U1402 (N_1402,N_1325,N_1397);
nand U1403 (N_1403,N_1376,N_1302);
nand U1404 (N_1404,N_1350,N_1394);
and U1405 (N_1405,N_1363,N_1386);
or U1406 (N_1406,N_1372,N_1389);
and U1407 (N_1407,N_1382,N_1315);
and U1408 (N_1408,N_1318,N_1338);
nor U1409 (N_1409,N_1303,N_1335);
or U1410 (N_1410,N_1307,N_1322);
nor U1411 (N_1411,N_1396,N_1301);
and U1412 (N_1412,N_1388,N_1378);
or U1413 (N_1413,N_1373,N_1371);
nand U1414 (N_1414,N_1392,N_1351);
and U1415 (N_1415,N_1365,N_1317);
nand U1416 (N_1416,N_1349,N_1336);
nand U1417 (N_1417,N_1334,N_1379);
nand U1418 (N_1418,N_1359,N_1331);
nand U1419 (N_1419,N_1311,N_1374);
nand U1420 (N_1420,N_1310,N_1381);
nor U1421 (N_1421,N_1362,N_1300);
nand U1422 (N_1422,N_1324,N_1370);
nor U1423 (N_1423,N_1312,N_1393);
xnor U1424 (N_1424,N_1354,N_1326);
nand U1425 (N_1425,N_1314,N_1390);
nor U1426 (N_1426,N_1348,N_1305);
xnor U1427 (N_1427,N_1369,N_1368);
nor U1428 (N_1428,N_1306,N_1356);
and U1429 (N_1429,N_1341,N_1319);
nor U1430 (N_1430,N_1377,N_1399);
and U1431 (N_1431,N_1357,N_1367);
nand U1432 (N_1432,N_1327,N_1340);
and U1433 (N_1433,N_1391,N_1353);
nor U1434 (N_1434,N_1316,N_1352);
nor U1435 (N_1435,N_1358,N_1395);
nand U1436 (N_1436,N_1330,N_1347);
xor U1437 (N_1437,N_1355,N_1313);
and U1438 (N_1438,N_1384,N_1345);
and U1439 (N_1439,N_1329,N_1360);
xnor U1440 (N_1440,N_1383,N_1366);
nand U1441 (N_1441,N_1337,N_1361);
nor U1442 (N_1442,N_1323,N_1380);
nand U1443 (N_1443,N_1343,N_1344);
nand U1444 (N_1444,N_1346,N_1339);
or U1445 (N_1445,N_1308,N_1342);
or U1446 (N_1446,N_1387,N_1333);
nand U1447 (N_1447,N_1309,N_1328);
and U1448 (N_1448,N_1321,N_1375);
nand U1449 (N_1449,N_1385,N_1332);
and U1450 (N_1450,N_1389,N_1377);
or U1451 (N_1451,N_1355,N_1362);
nor U1452 (N_1452,N_1387,N_1356);
nand U1453 (N_1453,N_1331,N_1308);
nor U1454 (N_1454,N_1345,N_1343);
and U1455 (N_1455,N_1353,N_1376);
nor U1456 (N_1456,N_1324,N_1372);
and U1457 (N_1457,N_1333,N_1355);
nand U1458 (N_1458,N_1312,N_1307);
and U1459 (N_1459,N_1305,N_1350);
nand U1460 (N_1460,N_1319,N_1361);
nor U1461 (N_1461,N_1305,N_1336);
nor U1462 (N_1462,N_1363,N_1376);
nand U1463 (N_1463,N_1369,N_1332);
nor U1464 (N_1464,N_1389,N_1344);
xor U1465 (N_1465,N_1399,N_1373);
and U1466 (N_1466,N_1397,N_1308);
or U1467 (N_1467,N_1385,N_1326);
nor U1468 (N_1468,N_1362,N_1341);
nor U1469 (N_1469,N_1305,N_1349);
and U1470 (N_1470,N_1344,N_1302);
or U1471 (N_1471,N_1370,N_1361);
or U1472 (N_1472,N_1368,N_1320);
and U1473 (N_1473,N_1396,N_1387);
nand U1474 (N_1474,N_1304,N_1337);
and U1475 (N_1475,N_1309,N_1374);
or U1476 (N_1476,N_1385,N_1383);
nor U1477 (N_1477,N_1389,N_1347);
xnor U1478 (N_1478,N_1331,N_1347);
or U1479 (N_1479,N_1356,N_1386);
xor U1480 (N_1480,N_1399,N_1306);
nor U1481 (N_1481,N_1353,N_1364);
or U1482 (N_1482,N_1314,N_1327);
and U1483 (N_1483,N_1350,N_1386);
and U1484 (N_1484,N_1387,N_1307);
nor U1485 (N_1485,N_1310,N_1330);
or U1486 (N_1486,N_1379,N_1349);
xnor U1487 (N_1487,N_1346,N_1375);
nor U1488 (N_1488,N_1311,N_1383);
nand U1489 (N_1489,N_1382,N_1321);
nor U1490 (N_1490,N_1323,N_1353);
or U1491 (N_1491,N_1330,N_1341);
or U1492 (N_1492,N_1311,N_1317);
nand U1493 (N_1493,N_1332,N_1351);
and U1494 (N_1494,N_1357,N_1384);
and U1495 (N_1495,N_1365,N_1368);
nand U1496 (N_1496,N_1300,N_1355);
nor U1497 (N_1497,N_1316,N_1399);
or U1498 (N_1498,N_1383,N_1352);
or U1499 (N_1499,N_1339,N_1373);
nor U1500 (N_1500,N_1405,N_1446);
xor U1501 (N_1501,N_1491,N_1479);
and U1502 (N_1502,N_1439,N_1425);
and U1503 (N_1503,N_1492,N_1459);
xnor U1504 (N_1504,N_1403,N_1462);
nand U1505 (N_1505,N_1493,N_1400);
nor U1506 (N_1506,N_1488,N_1418);
nor U1507 (N_1507,N_1453,N_1447);
or U1508 (N_1508,N_1430,N_1489);
nor U1509 (N_1509,N_1428,N_1407);
and U1510 (N_1510,N_1474,N_1431);
nand U1511 (N_1511,N_1499,N_1477);
or U1512 (N_1512,N_1461,N_1454);
or U1513 (N_1513,N_1448,N_1427);
and U1514 (N_1514,N_1498,N_1436);
nor U1515 (N_1515,N_1424,N_1438);
and U1516 (N_1516,N_1402,N_1412);
and U1517 (N_1517,N_1470,N_1467);
nor U1518 (N_1518,N_1455,N_1443);
nand U1519 (N_1519,N_1476,N_1457);
xnor U1520 (N_1520,N_1435,N_1450);
nand U1521 (N_1521,N_1495,N_1415);
nor U1522 (N_1522,N_1475,N_1440);
and U1523 (N_1523,N_1401,N_1496);
nor U1524 (N_1524,N_1497,N_1458);
nor U1525 (N_1525,N_1421,N_1411);
xor U1526 (N_1526,N_1445,N_1406);
or U1527 (N_1527,N_1444,N_1449);
nor U1528 (N_1528,N_1451,N_1464);
and U1529 (N_1529,N_1441,N_1490);
nand U1530 (N_1530,N_1478,N_1442);
nand U1531 (N_1531,N_1466,N_1423);
nor U1532 (N_1532,N_1416,N_1486);
nor U1533 (N_1533,N_1433,N_1460);
nand U1534 (N_1534,N_1463,N_1484);
xnor U1535 (N_1535,N_1409,N_1465);
or U1536 (N_1536,N_1422,N_1429);
xnor U1537 (N_1537,N_1452,N_1414);
nor U1538 (N_1538,N_1408,N_1437);
nor U1539 (N_1539,N_1413,N_1404);
nor U1540 (N_1540,N_1471,N_1483);
nand U1541 (N_1541,N_1410,N_1469);
nor U1542 (N_1542,N_1419,N_1432);
nand U1543 (N_1543,N_1434,N_1485);
and U1544 (N_1544,N_1487,N_1481);
or U1545 (N_1545,N_1482,N_1417);
and U1546 (N_1546,N_1473,N_1472);
nand U1547 (N_1547,N_1426,N_1468);
nor U1548 (N_1548,N_1420,N_1456);
nand U1549 (N_1549,N_1480,N_1494);
nor U1550 (N_1550,N_1473,N_1402);
or U1551 (N_1551,N_1448,N_1472);
nand U1552 (N_1552,N_1441,N_1405);
and U1553 (N_1553,N_1463,N_1406);
nor U1554 (N_1554,N_1463,N_1421);
nand U1555 (N_1555,N_1446,N_1401);
nand U1556 (N_1556,N_1425,N_1459);
xnor U1557 (N_1557,N_1454,N_1456);
nand U1558 (N_1558,N_1442,N_1424);
and U1559 (N_1559,N_1461,N_1492);
or U1560 (N_1560,N_1472,N_1483);
nand U1561 (N_1561,N_1400,N_1421);
nor U1562 (N_1562,N_1455,N_1414);
nand U1563 (N_1563,N_1434,N_1419);
xor U1564 (N_1564,N_1420,N_1458);
nor U1565 (N_1565,N_1476,N_1444);
or U1566 (N_1566,N_1426,N_1460);
xor U1567 (N_1567,N_1423,N_1412);
or U1568 (N_1568,N_1473,N_1457);
and U1569 (N_1569,N_1432,N_1465);
or U1570 (N_1570,N_1480,N_1478);
xor U1571 (N_1571,N_1433,N_1484);
nand U1572 (N_1572,N_1483,N_1412);
or U1573 (N_1573,N_1412,N_1455);
or U1574 (N_1574,N_1465,N_1496);
or U1575 (N_1575,N_1464,N_1453);
xor U1576 (N_1576,N_1432,N_1453);
nand U1577 (N_1577,N_1415,N_1494);
nand U1578 (N_1578,N_1476,N_1478);
nor U1579 (N_1579,N_1434,N_1448);
or U1580 (N_1580,N_1469,N_1494);
nand U1581 (N_1581,N_1413,N_1416);
nor U1582 (N_1582,N_1457,N_1472);
nor U1583 (N_1583,N_1458,N_1445);
and U1584 (N_1584,N_1477,N_1439);
xnor U1585 (N_1585,N_1433,N_1409);
nor U1586 (N_1586,N_1477,N_1474);
or U1587 (N_1587,N_1431,N_1470);
or U1588 (N_1588,N_1452,N_1427);
or U1589 (N_1589,N_1484,N_1408);
xnor U1590 (N_1590,N_1492,N_1423);
nor U1591 (N_1591,N_1466,N_1464);
and U1592 (N_1592,N_1420,N_1453);
nand U1593 (N_1593,N_1483,N_1414);
nor U1594 (N_1594,N_1483,N_1463);
xor U1595 (N_1595,N_1413,N_1467);
and U1596 (N_1596,N_1428,N_1489);
nor U1597 (N_1597,N_1406,N_1456);
nand U1598 (N_1598,N_1438,N_1456);
or U1599 (N_1599,N_1445,N_1430);
or U1600 (N_1600,N_1552,N_1544);
nor U1601 (N_1601,N_1515,N_1537);
nor U1602 (N_1602,N_1581,N_1592);
nand U1603 (N_1603,N_1571,N_1531);
nand U1604 (N_1604,N_1587,N_1597);
and U1605 (N_1605,N_1559,N_1555);
nor U1606 (N_1606,N_1577,N_1586);
nor U1607 (N_1607,N_1504,N_1560);
xor U1608 (N_1608,N_1599,N_1510);
nand U1609 (N_1609,N_1520,N_1532);
xnor U1610 (N_1610,N_1543,N_1512);
nor U1611 (N_1611,N_1536,N_1516);
or U1612 (N_1612,N_1524,N_1598);
or U1613 (N_1613,N_1527,N_1562);
nor U1614 (N_1614,N_1549,N_1538);
nor U1615 (N_1615,N_1548,N_1566);
or U1616 (N_1616,N_1564,N_1593);
or U1617 (N_1617,N_1541,N_1584);
or U1618 (N_1618,N_1530,N_1525);
and U1619 (N_1619,N_1579,N_1568);
nand U1620 (N_1620,N_1570,N_1569);
nor U1621 (N_1621,N_1540,N_1589);
and U1622 (N_1622,N_1526,N_1563);
or U1623 (N_1623,N_1500,N_1539);
nor U1624 (N_1624,N_1523,N_1521);
or U1625 (N_1625,N_1561,N_1573);
and U1626 (N_1626,N_1575,N_1533);
and U1627 (N_1627,N_1535,N_1580);
and U1628 (N_1628,N_1576,N_1553);
nor U1629 (N_1629,N_1517,N_1519);
or U1630 (N_1630,N_1550,N_1578);
nand U1631 (N_1631,N_1583,N_1596);
and U1632 (N_1632,N_1514,N_1547);
nand U1633 (N_1633,N_1502,N_1545);
or U1634 (N_1634,N_1501,N_1585);
or U1635 (N_1635,N_1529,N_1542);
nand U1636 (N_1636,N_1591,N_1518);
nand U1637 (N_1637,N_1594,N_1511);
nor U1638 (N_1638,N_1590,N_1513);
xnor U1639 (N_1639,N_1509,N_1522);
or U1640 (N_1640,N_1506,N_1558);
or U1641 (N_1641,N_1505,N_1588);
or U1642 (N_1642,N_1546,N_1565);
and U1643 (N_1643,N_1534,N_1528);
and U1644 (N_1644,N_1557,N_1595);
and U1645 (N_1645,N_1554,N_1556);
nor U1646 (N_1646,N_1503,N_1582);
nor U1647 (N_1647,N_1572,N_1551);
nor U1648 (N_1648,N_1508,N_1567);
nand U1649 (N_1649,N_1574,N_1507);
and U1650 (N_1650,N_1527,N_1572);
nand U1651 (N_1651,N_1506,N_1593);
and U1652 (N_1652,N_1577,N_1516);
nand U1653 (N_1653,N_1503,N_1505);
nor U1654 (N_1654,N_1575,N_1523);
or U1655 (N_1655,N_1577,N_1539);
and U1656 (N_1656,N_1512,N_1535);
nand U1657 (N_1657,N_1579,N_1502);
and U1658 (N_1658,N_1584,N_1521);
or U1659 (N_1659,N_1532,N_1501);
nor U1660 (N_1660,N_1583,N_1540);
and U1661 (N_1661,N_1523,N_1551);
nor U1662 (N_1662,N_1527,N_1595);
and U1663 (N_1663,N_1504,N_1519);
and U1664 (N_1664,N_1516,N_1568);
xnor U1665 (N_1665,N_1508,N_1557);
or U1666 (N_1666,N_1599,N_1595);
and U1667 (N_1667,N_1553,N_1557);
nor U1668 (N_1668,N_1562,N_1569);
and U1669 (N_1669,N_1582,N_1535);
and U1670 (N_1670,N_1528,N_1552);
nor U1671 (N_1671,N_1514,N_1517);
nand U1672 (N_1672,N_1597,N_1512);
nand U1673 (N_1673,N_1566,N_1504);
or U1674 (N_1674,N_1548,N_1509);
or U1675 (N_1675,N_1536,N_1507);
xor U1676 (N_1676,N_1513,N_1524);
nand U1677 (N_1677,N_1557,N_1554);
nand U1678 (N_1678,N_1539,N_1511);
xnor U1679 (N_1679,N_1598,N_1517);
xnor U1680 (N_1680,N_1573,N_1553);
nand U1681 (N_1681,N_1519,N_1558);
nor U1682 (N_1682,N_1518,N_1550);
nor U1683 (N_1683,N_1512,N_1518);
nand U1684 (N_1684,N_1567,N_1594);
and U1685 (N_1685,N_1506,N_1553);
and U1686 (N_1686,N_1510,N_1568);
nand U1687 (N_1687,N_1590,N_1548);
or U1688 (N_1688,N_1589,N_1556);
nor U1689 (N_1689,N_1512,N_1510);
xnor U1690 (N_1690,N_1501,N_1503);
or U1691 (N_1691,N_1564,N_1540);
nand U1692 (N_1692,N_1553,N_1523);
and U1693 (N_1693,N_1596,N_1589);
and U1694 (N_1694,N_1555,N_1591);
or U1695 (N_1695,N_1557,N_1591);
xor U1696 (N_1696,N_1532,N_1552);
or U1697 (N_1697,N_1597,N_1582);
and U1698 (N_1698,N_1547,N_1597);
nor U1699 (N_1699,N_1568,N_1547);
or U1700 (N_1700,N_1682,N_1608);
nor U1701 (N_1701,N_1640,N_1670);
nand U1702 (N_1702,N_1607,N_1642);
nor U1703 (N_1703,N_1666,N_1684);
or U1704 (N_1704,N_1664,N_1652);
and U1705 (N_1705,N_1659,N_1648);
and U1706 (N_1706,N_1650,N_1634);
or U1707 (N_1707,N_1625,N_1658);
nor U1708 (N_1708,N_1679,N_1602);
and U1709 (N_1709,N_1606,N_1690);
or U1710 (N_1710,N_1691,N_1605);
xnor U1711 (N_1711,N_1636,N_1647);
or U1712 (N_1712,N_1678,N_1693);
or U1713 (N_1713,N_1614,N_1622);
or U1714 (N_1714,N_1694,N_1609);
nand U1715 (N_1715,N_1676,N_1600);
or U1716 (N_1716,N_1681,N_1621);
xor U1717 (N_1717,N_1677,N_1698);
or U1718 (N_1718,N_1637,N_1649);
nor U1719 (N_1719,N_1657,N_1692);
and U1720 (N_1720,N_1631,N_1624);
or U1721 (N_1721,N_1669,N_1687);
or U1722 (N_1722,N_1653,N_1633);
nand U1723 (N_1723,N_1645,N_1685);
nand U1724 (N_1724,N_1689,N_1641);
nor U1725 (N_1725,N_1663,N_1601);
or U1726 (N_1726,N_1646,N_1654);
or U1727 (N_1727,N_1617,N_1628);
and U1728 (N_1728,N_1632,N_1688);
or U1729 (N_1729,N_1630,N_1629);
nor U1730 (N_1730,N_1662,N_1644);
xor U1731 (N_1731,N_1620,N_1613);
nand U1732 (N_1732,N_1635,N_1603);
or U1733 (N_1733,N_1626,N_1699);
nor U1734 (N_1734,N_1667,N_1643);
nand U1735 (N_1735,N_1623,N_1673);
and U1736 (N_1736,N_1638,N_1672);
nand U1737 (N_1737,N_1619,N_1615);
nor U1738 (N_1738,N_1661,N_1627);
nor U1739 (N_1739,N_1695,N_1651);
nand U1740 (N_1740,N_1668,N_1610);
nand U1741 (N_1741,N_1686,N_1618);
or U1742 (N_1742,N_1655,N_1604);
and U1743 (N_1743,N_1697,N_1683);
nor U1744 (N_1744,N_1639,N_1674);
nor U1745 (N_1745,N_1696,N_1665);
or U1746 (N_1746,N_1660,N_1675);
nor U1747 (N_1747,N_1616,N_1671);
and U1748 (N_1748,N_1656,N_1611);
nor U1749 (N_1749,N_1612,N_1680);
or U1750 (N_1750,N_1619,N_1648);
and U1751 (N_1751,N_1656,N_1627);
nand U1752 (N_1752,N_1658,N_1663);
nand U1753 (N_1753,N_1660,N_1656);
or U1754 (N_1754,N_1640,N_1666);
or U1755 (N_1755,N_1676,N_1601);
and U1756 (N_1756,N_1676,N_1686);
and U1757 (N_1757,N_1618,N_1651);
and U1758 (N_1758,N_1658,N_1661);
or U1759 (N_1759,N_1650,N_1601);
and U1760 (N_1760,N_1681,N_1612);
xnor U1761 (N_1761,N_1677,N_1651);
and U1762 (N_1762,N_1687,N_1666);
nand U1763 (N_1763,N_1687,N_1683);
nand U1764 (N_1764,N_1630,N_1656);
and U1765 (N_1765,N_1638,N_1631);
nor U1766 (N_1766,N_1673,N_1664);
nor U1767 (N_1767,N_1618,N_1605);
and U1768 (N_1768,N_1668,N_1633);
nand U1769 (N_1769,N_1637,N_1611);
nand U1770 (N_1770,N_1624,N_1622);
and U1771 (N_1771,N_1671,N_1600);
and U1772 (N_1772,N_1657,N_1624);
nor U1773 (N_1773,N_1687,N_1697);
or U1774 (N_1774,N_1676,N_1652);
or U1775 (N_1775,N_1639,N_1679);
xnor U1776 (N_1776,N_1664,N_1626);
nor U1777 (N_1777,N_1616,N_1668);
nor U1778 (N_1778,N_1637,N_1679);
nand U1779 (N_1779,N_1641,N_1620);
nand U1780 (N_1780,N_1672,N_1668);
and U1781 (N_1781,N_1610,N_1632);
and U1782 (N_1782,N_1609,N_1633);
nor U1783 (N_1783,N_1659,N_1699);
or U1784 (N_1784,N_1676,N_1655);
nor U1785 (N_1785,N_1699,N_1619);
or U1786 (N_1786,N_1622,N_1665);
nand U1787 (N_1787,N_1669,N_1686);
nand U1788 (N_1788,N_1697,N_1615);
and U1789 (N_1789,N_1677,N_1609);
nor U1790 (N_1790,N_1623,N_1685);
or U1791 (N_1791,N_1601,N_1677);
nor U1792 (N_1792,N_1627,N_1684);
or U1793 (N_1793,N_1670,N_1644);
and U1794 (N_1794,N_1691,N_1684);
or U1795 (N_1795,N_1623,N_1644);
and U1796 (N_1796,N_1606,N_1669);
nand U1797 (N_1797,N_1697,N_1668);
nor U1798 (N_1798,N_1610,N_1641);
nor U1799 (N_1799,N_1647,N_1677);
nand U1800 (N_1800,N_1710,N_1723);
or U1801 (N_1801,N_1798,N_1712);
nor U1802 (N_1802,N_1794,N_1775);
xor U1803 (N_1803,N_1792,N_1726);
nor U1804 (N_1804,N_1790,N_1753);
nor U1805 (N_1805,N_1749,N_1709);
nand U1806 (N_1806,N_1740,N_1788);
nor U1807 (N_1807,N_1799,N_1724);
nand U1808 (N_1808,N_1744,N_1786);
xor U1809 (N_1809,N_1774,N_1751);
nand U1810 (N_1810,N_1702,N_1785);
or U1811 (N_1811,N_1787,N_1730);
and U1812 (N_1812,N_1720,N_1756);
or U1813 (N_1813,N_1797,N_1791);
nor U1814 (N_1814,N_1779,N_1731);
and U1815 (N_1815,N_1728,N_1732);
or U1816 (N_1816,N_1765,N_1700);
or U1817 (N_1817,N_1754,N_1736);
nand U1818 (N_1818,N_1750,N_1703);
nand U1819 (N_1819,N_1705,N_1752);
nand U1820 (N_1820,N_1721,N_1704);
and U1821 (N_1821,N_1738,N_1739);
xor U1822 (N_1822,N_1711,N_1745);
nor U1823 (N_1823,N_1769,N_1729);
or U1824 (N_1824,N_1773,N_1784);
nand U1825 (N_1825,N_1735,N_1718);
xor U1826 (N_1826,N_1757,N_1776);
or U1827 (N_1827,N_1717,N_1782);
nand U1828 (N_1828,N_1768,N_1734);
or U1829 (N_1829,N_1772,N_1715);
or U1830 (N_1830,N_1741,N_1793);
and U1831 (N_1831,N_1755,N_1746);
nor U1832 (N_1832,N_1771,N_1796);
or U1833 (N_1833,N_1789,N_1701);
or U1834 (N_1834,N_1707,N_1742);
nand U1835 (N_1835,N_1777,N_1708);
nor U1836 (N_1836,N_1780,N_1747);
xor U1837 (N_1837,N_1781,N_1763);
nand U1838 (N_1838,N_1758,N_1748);
xnor U1839 (N_1839,N_1743,N_1795);
nor U1840 (N_1840,N_1767,N_1783);
nand U1841 (N_1841,N_1766,N_1716);
nor U1842 (N_1842,N_1759,N_1727);
or U1843 (N_1843,N_1761,N_1762);
xnor U1844 (N_1844,N_1764,N_1733);
or U1845 (N_1845,N_1719,N_1760);
and U1846 (N_1846,N_1706,N_1714);
and U1847 (N_1847,N_1722,N_1725);
nand U1848 (N_1848,N_1778,N_1713);
nor U1849 (N_1849,N_1737,N_1770);
or U1850 (N_1850,N_1725,N_1775);
nor U1851 (N_1851,N_1790,N_1740);
or U1852 (N_1852,N_1787,N_1794);
and U1853 (N_1853,N_1789,N_1730);
and U1854 (N_1854,N_1756,N_1715);
or U1855 (N_1855,N_1739,N_1761);
xnor U1856 (N_1856,N_1799,N_1717);
and U1857 (N_1857,N_1760,N_1733);
and U1858 (N_1858,N_1764,N_1719);
nand U1859 (N_1859,N_1719,N_1780);
or U1860 (N_1860,N_1727,N_1799);
nor U1861 (N_1861,N_1738,N_1796);
and U1862 (N_1862,N_1763,N_1704);
nand U1863 (N_1863,N_1715,N_1781);
nor U1864 (N_1864,N_1739,N_1716);
or U1865 (N_1865,N_1766,N_1712);
nand U1866 (N_1866,N_1700,N_1781);
nor U1867 (N_1867,N_1757,N_1752);
nand U1868 (N_1868,N_1759,N_1765);
nand U1869 (N_1869,N_1770,N_1740);
or U1870 (N_1870,N_1743,N_1717);
nand U1871 (N_1871,N_1740,N_1774);
nand U1872 (N_1872,N_1764,N_1798);
nand U1873 (N_1873,N_1726,N_1771);
nand U1874 (N_1874,N_1758,N_1730);
and U1875 (N_1875,N_1703,N_1772);
nand U1876 (N_1876,N_1738,N_1708);
or U1877 (N_1877,N_1757,N_1726);
or U1878 (N_1878,N_1703,N_1738);
nor U1879 (N_1879,N_1720,N_1749);
or U1880 (N_1880,N_1710,N_1737);
and U1881 (N_1881,N_1734,N_1784);
or U1882 (N_1882,N_1718,N_1720);
or U1883 (N_1883,N_1775,N_1735);
and U1884 (N_1884,N_1760,N_1711);
nand U1885 (N_1885,N_1760,N_1752);
nand U1886 (N_1886,N_1794,N_1706);
or U1887 (N_1887,N_1798,N_1739);
xor U1888 (N_1888,N_1754,N_1739);
nor U1889 (N_1889,N_1766,N_1742);
nand U1890 (N_1890,N_1790,N_1774);
nand U1891 (N_1891,N_1789,N_1756);
xnor U1892 (N_1892,N_1786,N_1797);
nor U1893 (N_1893,N_1781,N_1745);
and U1894 (N_1894,N_1729,N_1773);
nand U1895 (N_1895,N_1755,N_1783);
nor U1896 (N_1896,N_1729,N_1757);
xor U1897 (N_1897,N_1789,N_1712);
nor U1898 (N_1898,N_1717,N_1735);
or U1899 (N_1899,N_1740,N_1748);
and U1900 (N_1900,N_1805,N_1865);
xor U1901 (N_1901,N_1836,N_1881);
and U1902 (N_1902,N_1835,N_1840);
and U1903 (N_1903,N_1863,N_1882);
and U1904 (N_1904,N_1801,N_1866);
or U1905 (N_1905,N_1878,N_1856);
xnor U1906 (N_1906,N_1834,N_1850);
or U1907 (N_1907,N_1817,N_1853);
and U1908 (N_1908,N_1864,N_1831);
nor U1909 (N_1909,N_1854,N_1852);
nand U1910 (N_1910,N_1898,N_1824);
or U1911 (N_1911,N_1875,N_1803);
or U1912 (N_1912,N_1812,N_1883);
nor U1913 (N_1913,N_1804,N_1847);
xor U1914 (N_1914,N_1820,N_1855);
nand U1915 (N_1915,N_1838,N_1891);
or U1916 (N_1916,N_1877,N_1825);
nor U1917 (N_1917,N_1844,N_1816);
xnor U1918 (N_1918,N_1833,N_1897);
nand U1919 (N_1919,N_1813,N_1887);
and U1920 (N_1920,N_1886,N_1841);
xor U1921 (N_1921,N_1879,N_1807);
or U1922 (N_1922,N_1873,N_1839);
xnor U1923 (N_1923,N_1815,N_1861);
or U1924 (N_1924,N_1823,N_1806);
and U1925 (N_1925,N_1858,N_1848);
or U1926 (N_1926,N_1888,N_1880);
nor U1927 (N_1927,N_1829,N_1872);
or U1928 (N_1928,N_1862,N_1890);
xor U1929 (N_1929,N_1859,N_1899);
nand U1930 (N_1930,N_1828,N_1892);
xnor U1931 (N_1931,N_1822,N_1893);
or U1932 (N_1932,N_1811,N_1837);
xnor U1933 (N_1933,N_1800,N_1867);
nor U1934 (N_1934,N_1849,N_1819);
xnor U1935 (N_1935,N_1871,N_1896);
or U1936 (N_1936,N_1832,N_1826);
nand U1937 (N_1937,N_1814,N_1851);
nand U1938 (N_1938,N_1860,N_1885);
or U1939 (N_1939,N_1857,N_1870);
nor U1940 (N_1940,N_1808,N_1869);
or U1941 (N_1941,N_1846,N_1845);
nand U1942 (N_1942,N_1868,N_1810);
and U1943 (N_1943,N_1884,N_1874);
nor U1944 (N_1944,N_1818,N_1802);
nand U1945 (N_1945,N_1895,N_1876);
or U1946 (N_1946,N_1889,N_1843);
nor U1947 (N_1947,N_1827,N_1842);
nand U1948 (N_1948,N_1894,N_1821);
and U1949 (N_1949,N_1809,N_1830);
nor U1950 (N_1950,N_1867,N_1812);
or U1951 (N_1951,N_1852,N_1882);
nor U1952 (N_1952,N_1809,N_1831);
and U1953 (N_1953,N_1895,N_1817);
nor U1954 (N_1954,N_1823,N_1852);
or U1955 (N_1955,N_1824,N_1833);
or U1956 (N_1956,N_1897,N_1818);
nand U1957 (N_1957,N_1808,N_1867);
nand U1958 (N_1958,N_1844,N_1804);
nand U1959 (N_1959,N_1885,N_1846);
xnor U1960 (N_1960,N_1899,N_1890);
nor U1961 (N_1961,N_1856,N_1821);
or U1962 (N_1962,N_1806,N_1836);
and U1963 (N_1963,N_1828,N_1885);
nor U1964 (N_1964,N_1868,N_1833);
or U1965 (N_1965,N_1827,N_1882);
nand U1966 (N_1966,N_1807,N_1816);
nor U1967 (N_1967,N_1897,N_1877);
nor U1968 (N_1968,N_1807,N_1868);
and U1969 (N_1969,N_1837,N_1801);
or U1970 (N_1970,N_1821,N_1846);
nand U1971 (N_1971,N_1848,N_1838);
xnor U1972 (N_1972,N_1813,N_1817);
nand U1973 (N_1973,N_1884,N_1821);
or U1974 (N_1974,N_1874,N_1853);
and U1975 (N_1975,N_1823,N_1870);
nand U1976 (N_1976,N_1863,N_1883);
and U1977 (N_1977,N_1825,N_1835);
or U1978 (N_1978,N_1808,N_1874);
nand U1979 (N_1979,N_1845,N_1824);
and U1980 (N_1980,N_1808,N_1895);
and U1981 (N_1981,N_1814,N_1865);
and U1982 (N_1982,N_1892,N_1800);
xnor U1983 (N_1983,N_1896,N_1848);
and U1984 (N_1984,N_1813,N_1819);
or U1985 (N_1985,N_1873,N_1895);
nor U1986 (N_1986,N_1876,N_1801);
or U1987 (N_1987,N_1877,N_1813);
or U1988 (N_1988,N_1821,N_1886);
nor U1989 (N_1989,N_1871,N_1856);
nand U1990 (N_1990,N_1833,N_1886);
nand U1991 (N_1991,N_1845,N_1893);
and U1992 (N_1992,N_1803,N_1834);
and U1993 (N_1993,N_1843,N_1849);
nor U1994 (N_1994,N_1829,N_1843);
nor U1995 (N_1995,N_1831,N_1827);
nand U1996 (N_1996,N_1816,N_1899);
nand U1997 (N_1997,N_1813,N_1897);
nand U1998 (N_1998,N_1876,N_1846);
and U1999 (N_1999,N_1898,N_1813);
nor U2000 (N_2000,N_1971,N_1920);
or U2001 (N_2001,N_1927,N_1906);
and U2002 (N_2002,N_1910,N_1938);
nor U2003 (N_2003,N_1999,N_1909);
nand U2004 (N_2004,N_1961,N_1980);
nor U2005 (N_2005,N_1977,N_1953);
or U2006 (N_2006,N_1929,N_1955);
or U2007 (N_2007,N_1922,N_1900);
or U2008 (N_2008,N_1939,N_1950);
or U2009 (N_2009,N_1990,N_1930);
and U2010 (N_2010,N_1926,N_1985);
or U2011 (N_2011,N_1937,N_1905);
nand U2012 (N_2012,N_1951,N_1936);
or U2013 (N_2013,N_1989,N_1991);
and U2014 (N_2014,N_1981,N_1923);
nand U2015 (N_2015,N_1996,N_1988);
nor U2016 (N_2016,N_1946,N_1995);
or U2017 (N_2017,N_1944,N_1931);
nor U2018 (N_2018,N_1948,N_1998);
or U2019 (N_2019,N_1960,N_1984);
nor U2020 (N_2020,N_1940,N_1997);
or U2021 (N_2021,N_1916,N_1902);
nor U2022 (N_2022,N_1943,N_1915);
nand U2023 (N_2023,N_1970,N_1954);
nor U2024 (N_2024,N_1913,N_1963);
xor U2025 (N_2025,N_1982,N_1908);
nand U2026 (N_2026,N_1921,N_1952);
nand U2027 (N_2027,N_1945,N_1935);
and U2028 (N_2028,N_1966,N_1976);
nor U2029 (N_2029,N_1983,N_1975);
and U2030 (N_2030,N_1974,N_1912);
nor U2031 (N_2031,N_1919,N_1973);
and U2032 (N_2032,N_1965,N_1949);
and U2033 (N_2033,N_1993,N_1911);
nor U2034 (N_2034,N_1986,N_1928);
and U2035 (N_2035,N_1959,N_1957);
nand U2036 (N_2036,N_1958,N_1903);
or U2037 (N_2037,N_1901,N_1967);
xnor U2038 (N_2038,N_1994,N_1917);
and U2039 (N_2039,N_1969,N_1914);
nor U2040 (N_2040,N_1968,N_1956);
xnor U2041 (N_2041,N_1992,N_1932);
or U2042 (N_2042,N_1918,N_1962);
or U2043 (N_2043,N_1979,N_1987);
nand U2044 (N_2044,N_1934,N_1904);
and U2045 (N_2045,N_1907,N_1947);
nand U2046 (N_2046,N_1942,N_1925);
or U2047 (N_2047,N_1972,N_1924);
nand U2048 (N_2048,N_1964,N_1941);
or U2049 (N_2049,N_1978,N_1933);
nor U2050 (N_2050,N_1924,N_1908);
and U2051 (N_2051,N_1979,N_1968);
and U2052 (N_2052,N_1921,N_1965);
nor U2053 (N_2053,N_1977,N_1964);
nand U2054 (N_2054,N_1905,N_1966);
and U2055 (N_2055,N_1929,N_1950);
nor U2056 (N_2056,N_1978,N_1913);
and U2057 (N_2057,N_1990,N_1905);
xor U2058 (N_2058,N_1970,N_1956);
and U2059 (N_2059,N_1941,N_1952);
or U2060 (N_2060,N_1998,N_1987);
and U2061 (N_2061,N_1956,N_1997);
nand U2062 (N_2062,N_1924,N_1991);
nand U2063 (N_2063,N_1922,N_1955);
and U2064 (N_2064,N_1977,N_1900);
nor U2065 (N_2065,N_1936,N_1919);
nand U2066 (N_2066,N_1900,N_1956);
nand U2067 (N_2067,N_1999,N_1940);
xor U2068 (N_2068,N_1935,N_1926);
or U2069 (N_2069,N_1957,N_1932);
or U2070 (N_2070,N_1936,N_1913);
and U2071 (N_2071,N_1960,N_1969);
nor U2072 (N_2072,N_1980,N_1981);
nand U2073 (N_2073,N_1937,N_1900);
xor U2074 (N_2074,N_1909,N_1974);
nand U2075 (N_2075,N_1994,N_1982);
or U2076 (N_2076,N_1981,N_1933);
nand U2077 (N_2077,N_1986,N_1946);
nor U2078 (N_2078,N_1952,N_1949);
or U2079 (N_2079,N_1935,N_1938);
nand U2080 (N_2080,N_1989,N_1964);
or U2081 (N_2081,N_1927,N_1948);
nor U2082 (N_2082,N_1915,N_1917);
xnor U2083 (N_2083,N_1991,N_1944);
or U2084 (N_2084,N_1926,N_1964);
or U2085 (N_2085,N_1937,N_1918);
nand U2086 (N_2086,N_1960,N_1959);
nand U2087 (N_2087,N_1928,N_1930);
and U2088 (N_2088,N_1938,N_1968);
nor U2089 (N_2089,N_1951,N_1948);
or U2090 (N_2090,N_1917,N_1925);
or U2091 (N_2091,N_1991,N_1971);
nand U2092 (N_2092,N_1907,N_1954);
nor U2093 (N_2093,N_1911,N_1968);
xnor U2094 (N_2094,N_1925,N_1997);
or U2095 (N_2095,N_1974,N_1941);
xnor U2096 (N_2096,N_1950,N_1953);
and U2097 (N_2097,N_1908,N_1938);
and U2098 (N_2098,N_1912,N_1952);
nand U2099 (N_2099,N_1946,N_1971);
nand U2100 (N_2100,N_2053,N_2071);
xnor U2101 (N_2101,N_2091,N_2058);
or U2102 (N_2102,N_2040,N_2046);
nand U2103 (N_2103,N_2056,N_2067);
or U2104 (N_2104,N_2032,N_2083);
nand U2105 (N_2105,N_2015,N_2059);
nor U2106 (N_2106,N_2068,N_2024);
and U2107 (N_2107,N_2051,N_2026);
or U2108 (N_2108,N_2061,N_2044);
and U2109 (N_2109,N_2092,N_2094);
nor U2110 (N_2110,N_2084,N_2076);
nand U2111 (N_2111,N_2002,N_2037);
nand U2112 (N_2112,N_2004,N_2035);
nor U2113 (N_2113,N_2078,N_2020);
nor U2114 (N_2114,N_2033,N_2003);
xnor U2115 (N_2115,N_2077,N_2013);
nor U2116 (N_2116,N_2036,N_2034);
or U2117 (N_2117,N_2066,N_2018);
and U2118 (N_2118,N_2014,N_2050);
nand U2119 (N_2119,N_2049,N_2043);
nor U2120 (N_2120,N_2028,N_2087);
or U2121 (N_2121,N_2021,N_2027);
nor U2122 (N_2122,N_2069,N_2093);
or U2123 (N_2123,N_2081,N_2030);
nand U2124 (N_2124,N_2029,N_2011);
nor U2125 (N_2125,N_2047,N_2060);
nand U2126 (N_2126,N_2096,N_2086);
or U2127 (N_2127,N_2023,N_2007);
or U2128 (N_2128,N_2006,N_2089);
or U2129 (N_2129,N_2064,N_2097);
nand U2130 (N_2130,N_2005,N_2070);
nor U2131 (N_2131,N_2012,N_2016);
nor U2132 (N_2132,N_2079,N_2042);
and U2133 (N_2133,N_2055,N_2080);
and U2134 (N_2134,N_2065,N_2031);
and U2135 (N_2135,N_2038,N_2045);
and U2136 (N_2136,N_2075,N_2095);
nor U2137 (N_2137,N_2009,N_2039);
and U2138 (N_2138,N_2054,N_2022);
nand U2139 (N_2139,N_2017,N_2085);
and U2140 (N_2140,N_2073,N_2010);
nand U2141 (N_2141,N_2000,N_2041);
nor U2142 (N_2142,N_2062,N_2074);
nor U2143 (N_2143,N_2082,N_2099);
nor U2144 (N_2144,N_2008,N_2057);
nor U2145 (N_2145,N_2063,N_2072);
nor U2146 (N_2146,N_2052,N_2019);
or U2147 (N_2147,N_2001,N_2098);
nor U2148 (N_2148,N_2090,N_2025);
or U2149 (N_2149,N_2088,N_2048);
or U2150 (N_2150,N_2011,N_2071);
nand U2151 (N_2151,N_2027,N_2069);
xnor U2152 (N_2152,N_2015,N_2054);
nand U2153 (N_2153,N_2077,N_2042);
xnor U2154 (N_2154,N_2019,N_2099);
or U2155 (N_2155,N_2079,N_2064);
nand U2156 (N_2156,N_2015,N_2009);
nor U2157 (N_2157,N_2034,N_2061);
and U2158 (N_2158,N_2074,N_2040);
and U2159 (N_2159,N_2095,N_2090);
xnor U2160 (N_2160,N_2011,N_2056);
nor U2161 (N_2161,N_2018,N_2080);
nor U2162 (N_2162,N_2089,N_2031);
xor U2163 (N_2163,N_2096,N_2022);
nor U2164 (N_2164,N_2006,N_2090);
nor U2165 (N_2165,N_2031,N_2028);
and U2166 (N_2166,N_2061,N_2089);
nor U2167 (N_2167,N_2071,N_2062);
or U2168 (N_2168,N_2048,N_2085);
nor U2169 (N_2169,N_2008,N_2034);
or U2170 (N_2170,N_2011,N_2092);
and U2171 (N_2171,N_2007,N_2075);
or U2172 (N_2172,N_2090,N_2084);
xnor U2173 (N_2173,N_2024,N_2057);
or U2174 (N_2174,N_2088,N_2021);
nand U2175 (N_2175,N_2093,N_2083);
and U2176 (N_2176,N_2002,N_2044);
nor U2177 (N_2177,N_2005,N_2050);
or U2178 (N_2178,N_2050,N_2029);
nor U2179 (N_2179,N_2064,N_2004);
and U2180 (N_2180,N_2071,N_2084);
nor U2181 (N_2181,N_2034,N_2027);
and U2182 (N_2182,N_2044,N_2028);
nor U2183 (N_2183,N_2016,N_2067);
nand U2184 (N_2184,N_2043,N_2034);
nor U2185 (N_2185,N_2077,N_2016);
and U2186 (N_2186,N_2090,N_2052);
xnor U2187 (N_2187,N_2014,N_2064);
nand U2188 (N_2188,N_2096,N_2026);
or U2189 (N_2189,N_2066,N_2084);
nor U2190 (N_2190,N_2089,N_2062);
or U2191 (N_2191,N_2098,N_2050);
or U2192 (N_2192,N_2006,N_2030);
and U2193 (N_2193,N_2021,N_2024);
and U2194 (N_2194,N_2093,N_2007);
and U2195 (N_2195,N_2049,N_2073);
xor U2196 (N_2196,N_2095,N_2008);
nand U2197 (N_2197,N_2004,N_2087);
and U2198 (N_2198,N_2009,N_2002);
nor U2199 (N_2199,N_2023,N_2032);
nor U2200 (N_2200,N_2132,N_2165);
or U2201 (N_2201,N_2163,N_2109);
or U2202 (N_2202,N_2199,N_2171);
and U2203 (N_2203,N_2145,N_2197);
or U2204 (N_2204,N_2164,N_2184);
nand U2205 (N_2205,N_2162,N_2127);
nor U2206 (N_2206,N_2156,N_2123);
xor U2207 (N_2207,N_2181,N_2129);
or U2208 (N_2208,N_2153,N_2144);
or U2209 (N_2209,N_2125,N_2108);
and U2210 (N_2210,N_2169,N_2140);
nor U2211 (N_2211,N_2102,N_2170);
and U2212 (N_2212,N_2186,N_2150);
nand U2213 (N_2213,N_2159,N_2126);
nor U2214 (N_2214,N_2101,N_2158);
xor U2215 (N_2215,N_2106,N_2152);
and U2216 (N_2216,N_2183,N_2138);
nor U2217 (N_2217,N_2139,N_2118);
or U2218 (N_2218,N_2133,N_2180);
xor U2219 (N_2219,N_2122,N_2105);
or U2220 (N_2220,N_2148,N_2188);
or U2221 (N_2221,N_2185,N_2187);
or U2222 (N_2222,N_2117,N_2111);
or U2223 (N_2223,N_2104,N_2137);
nand U2224 (N_2224,N_2174,N_2113);
nor U2225 (N_2225,N_2179,N_2114);
or U2226 (N_2226,N_2120,N_2190);
nand U2227 (N_2227,N_2124,N_2131);
nor U2228 (N_2228,N_2154,N_2119);
and U2229 (N_2229,N_2167,N_2130);
and U2230 (N_2230,N_2166,N_2110);
xor U2231 (N_2231,N_2193,N_2178);
or U2232 (N_2232,N_2182,N_2142);
nand U2233 (N_2233,N_2146,N_2191);
nand U2234 (N_2234,N_2161,N_2189);
or U2235 (N_2235,N_2115,N_2112);
or U2236 (N_2236,N_2177,N_2151);
xor U2237 (N_2237,N_2135,N_2196);
and U2238 (N_2238,N_2195,N_2116);
and U2239 (N_2239,N_2141,N_2149);
and U2240 (N_2240,N_2128,N_2168);
or U2241 (N_2241,N_2107,N_2198);
nand U2242 (N_2242,N_2194,N_2172);
xor U2243 (N_2243,N_2121,N_2175);
nand U2244 (N_2244,N_2103,N_2160);
nor U2245 (N_2245,N_2143,N_2176);
nor U2246 (N_2246,N_2136,N_2173);
or U2247 (N_2247,N_2155,N_2147);
and U2248 (N_2248,N_2100,N_2192);
nor U2249 (N_2249,N_2134,N_2157);
or U2250 (N_2250,N_2199,N_2110);
xor U2251 (N_2251,N_2131,N_2110);
and U2252 (N_2252,N_2189,N_2101);
or U2253 (N_2253,N_2183,N_2123);
and U2254 (N_2254,N_2161,N_2156);
nor U2255 (N_2255,N_2191,N_2108);
or U2256 (N_2256,N_2171,N_2151);
nor U2257 (N_2257,N_2164,N_2144);
and U2258 (N_2258,N_2164,N_2151);
and U2259 (N_2259,N_2173,N_2119);
or U2260 (N_2260,N_2151,N_2168);
and U2261 (N_2261,N_2162,N_2172);
nor U2262 (N_2262,N_2186,N_2163);
nand U2263 (N_2263,N_2146,N_2120);
and U2264 (N_2264,N_2110,N_2156);
nand U2265 (N_2265,N_2173,N_2157);
or U2266 (N_2266,N_2114,N_2123);
nand U2267 (N_2267,N_2169,N_2124);
nand U2268 (N_2268,N_2157,N_2183);
nand U2269 (N_2269,N_2107,N_2160);
nand U2270 (N_2270,N_2138,N_2120);
xor U2271 (N_2271,N_2131,N_2121);
nor U2272 (N_2272,N_2145,N_2134);
nand U2273 (N_2273,N_2117,N_2184);
and U2274 (N_2274,N_2111,N_2155);
or U2275 (N_2275,N_2132,N_2136);
nand U2276 (N_2276,N_2119,N_2179);
and U2277 (N_2277,N_2191,N_2110);
or U2278 (N_2278,N_2103,N_2182);
or U2279 (N_2279,N_2159,N_2138);
or U2280 (N_2280,N_2177,N_2198);
and U2281 (N_2281,N_2175,N_2176);
nand U2282 (N_2282,N_2133,N_2184);
or U2283 (N_2283,N_2155,N_2149);
or U2284 (N_2284,N_2151,N_2154);
xor U2285 (N_2285,N_2145,N_2180);
or U2286 (N_2286,N_2180,N_2164);
and U2287 (N_2287,N_2141,N_2116);
or U2288 (N_2288,N_2105,N_2155);
xor U2289 (N_2289,N_2164,N_2115);
nor U2290 (N_2290,N_2159,N_2134);
and U2291 (N_2291,N_2184,N_2120);
or U2292 (N_2292,N_2122,N_2120);
or U2293 (N_2293,N_2180,N_2161);
or U2294 (N_2294,N_2158,N_2128);
and U2295 (N_2295,N_2159,N_2164);
nand U2296 (N_2296,N_2197,N_2120);
nand U2297 (N_2297,N_2138,N_2179);
xnor U2298 (N_2298,N_2174,N_2118);
and U2299 (N_2299,N_2144,N_2148);
xor U2300 (N_2300,N_2217,N_2203);
nor U2301 (N_2301,N_2278,N_2293);
nand U2302 (N_2302,N_2290,N_2231);
nand U2303 (N_2303,N_2291,N_2210);
and U2304 (N_2304,N_2219,N_2224);
and U2305 (N_2305,N_2202,N_2258);
and U2306 (N_2306,N_2286,N_2280);
xor U2307 (N_2307,N_2226,N_2213);
nand U2308 (N_2308,N_2241,N_2297);
nand U2309 (N_2309,N_2264,N_2296);
nand U2310 (N_2310,N_2265,N_2223);
or U2311 (N_2311,N_2272,N_2228);
nand U2312 (N_2312,N_2220,N_2222);
or U2313 (N_2313,N_2232,N_2242);
and U2314 (N_2314,N_2263,N_2214);
or U2315 (N_2315,N_2225,N_2256);
and U2316 (N_2316,N_2234,N_2235);
nand U2317 (N_2317,N_2243,N_2211);
nand U2318 (N_2318,N_2245,N_2298);
xor U2319 (N_2319,N_2246,N_2215);
or U2320 (N_2320,N_2287,N_2244);
nor U2321 (N_2321,N_2257,N_2294);
xnor U2322 (N_2322,N_2201,N_2284);
xor U2323 (N_2323,N_2255,N_2292);
and U2324 (N_2324,N_2285,N_2208);
nand U2325 (N_2325,N_2206,N_2249);
nand U2326 (N_2326,N_2299,N_2267);
and U2327 (N_2327,N_2227,N_2262);
or U2328 (N_2328,N_2248,N_2200);
nor U2329 (N_2329,N_2282,N_2266);
and U2330 (N_2330,N_2271,N_2261);
or U2331 (N_2331,N_2279,N_2295);
xor U2332 (N_2332,N_2221,N_2288);
nor U2333 (N_2333,N_2273,N_2270);
nand U2334 (N_2334,N_2269,N_2230);
and U2335 (N_2335,N_2229,N_2268);
and U2336 (N_2336,N_2274,N_2216);
nand U2337 (N_2337,N_2233,N_2239);
or U2338 (N_2338,N_2250,N_2275);
and U2339 (N_2339,N_2283,N_2251);
nor U2340 (N_2340,N_2207,N_2212);
nand U2341 (N_2341,N_2277,N_2238);
nand U2342 (N_2342,N_2253,N_2205);
nor U2343 (N_2343,N_2276,N_2240);
nor U2344 (N_2344,N_2218,N_2254);
nor U2345 (N_2345,N_2252,N_2237);
nand U2346 (N_2346,N_2236,N_2247);
nand U2347 (N_2347,N_2289,N_2259);
or U2348 (N_2348,N_2204,N_2260);
or U2349 (N_2349,N_2281,N_2209);
nor U2350 (N_2350,N_2274,N_2276);
nand U2351 (N_2351,N_2271,N_2206);
or U2352 (N_2352,N_2234,N_2201);
nand U2353 (N_2353,N_2244,N_2216);
and U2354 (N_2354,N_2278,N_2205);
or U2355 (N_2355,N_2267,N_2283);
and U2356 (N_2356,N_2274,N_2272);
nand U2357 (N_2357,N_2254,N_2223);
nor U2358 (N_2358,N_2275,N_2235);
nor U2359 (N_2359,N_2284,N_2217);
and U2360 (N_2360,N_2210,N_2248);
and U2361 (N_2361,N_2234,N_2262);
and U2362 (N_2362,N_2293,N_2273);
nor U2363 (N_2363,N_2283,N_2213);
and U2364 (N_2364,N_2258,N_2288);
nor U2365 (N_2365,N_2246,N_2248);
nor U2366 (N_2366,N_2216,N_2269);
nand U2367 (N_2367,N_2228,N_2243);
nand U2368 (N_2368,N_2220,N_2294);
or U2369 (N_2369,N_2225,N_2269);
or U2370 (N_2370,N_2201,N_2264);
nor U2371 (N_2371,N_2286,N_2299);
nand U2372 (N_2372,N_2224,N_2211);
or U2373 (N_2373,N_2259,N_2234);
nor U2374 (N_2374,N_2287,N_2261);
nor U2375 (N_2375,N_2265,N_2296);
nand U2376 (N_2376,N_2276,N_2217);
or U2377 (N_2377,N_2206,N_2229);
and U2378 (N_2378,N_2293,N_2248);
nand U2379 (N_2379,N_2254,N_2243);
nand U2380 (N_2380,N_2214,N_2269);
nor U2381 (N_2381,N_2269,N_2209);
nand U2382 (N_2382,N_2208,N_2232);
or U2383 (N_2383,N_2223,N_2252);
and U2384 (N_2384,N_2211,N_2244);
nand U2385 (N_2385,N_2278,N_2274);
or U2386 (N_2386,N_2220,N_2261);
and U2387 (N_2387,N_2284,N_2224);
xnor U2388 (N_2388,N_2271,N_2258);
nand U2389 (N_2389,N_2254,N_2238);
and U2390 (N_2390,N_2257,N_2255);
and U2391 (N_2391,N_2245,N_2201);
or U2392 (N_2392,N_2234,N_2243);
nor U2393 (N_2393,N_2288,N_2263);
nor U2394 (N_2394,N_2223,N_2245);
nand U2395 (N_2395,N_2214,N_2295);
nor U2396 (N_2396,N_2207,N_2233);
and U2397 (N_2397,N_2250,N_2247);
nor U2398 (N_2398,N_2291,N_2267);
nor U2399 (N_2399,N_2222,N_2265);
or U2400 (N_2400,N_2343,N_2383);
xnor U2401 (N_2401,N_2360,N_2374);
or U2402 (N_2402,N_2317,N_2396);
nand U2403 (N_2403,N_2369,N_2395);
and U2404 (N_2404,N_2361,N_2332);
nor U2405 (N_2405,N_2398,N_2375);
nand U2406 (N_2406,N_2384,N_2393);
and U2407 (N_2407,N_2337,N_2351);
and U2408 (N_2408,N_2391,N_2344);
and U2409 (N_2409,N_2304,N_2379);
and U2410 (N_2410,N_2311,N_2368);
and U2411 (N_2411,N_2365,N_2328);
nand U2412 (N_2412,N_2370,N_2386);
and U2413 (N_2413,N_2373,N_2363);
and U2414 (N_2414,N_2346,N_2308);
or U2415 (N_2415,N_2339,N_2342);
nand U2416 (N_2416,N_2358,N_2348);
xor U2417 (N_2417,N_2335,N_2338);
xnor U2418 (N_2418,N_2330,N_2366);
nor U2419 (N_2419,N_2359,N_2319);
and U2420 (N_2420,N_2322,N_2385);
or U2421 (N_2421,N_2301,N_2313);
nor U2422 (N_2422,N_2323,N_2307);
or U2423 (N_2423,N_2310,N_2325);
or U2424 (N_2424,N_2312,N_2371);
or U2425 (N_2425,N_2390,N_2336);
and U2426 (N_2426,N_2340,N_2354);
and U2427 (N_2427,N_2389,N_2353);
and U2428 (N_2428,N_2372,N_2394);
nor U2429 (N_2429,N_2352,N_2388);
and U2430 (N_2430,N_2318,N_2300);
or U2431 (N_2431,N_2324,N_2347);
or U2432 (N_2432,N_2349,N_2397);
nand U2433 (N_2433,N_2376,N_2320);
nand U2434 (N_2434,N_2355,N_2305);
and U2435 (N_2435,N_2333,N_2327);
or U2436 (N_2436,N_2326,N_2381);
nand U2437 (N_2437,N_2399,N_2331);
or U2438 (N_2438,N_2367,N_2314);
nor U2439 (N_2439,N_2334,N_2306);
nor U2440 (N_2440,N_2303,N_2380);
and U2441 (N_2441,N_2321,N_2382);
nor U2442 (N_2442,N_2302,N_2357);
and U2443 (N_2443,N_2341,N_2364);
or U2444 (N_2444,N_2378,N_2315);
nand U2445 (N_2445,N_2387,N_2345);
nand U2446 (N_2446,N_2316,N_2350);
nand U2447 (N_2447,N_2362,N_2329);
nand U2448 (N_2448,N_2392,N_2377);
nand U2449 (N_2449,N_2356,N_2309);
nor U2450 (N_2450,N_2349,N_2395);
and U2451 (N_2451,N_2323,N_2321);
or U2452 (N_2452,N_2340,N_2362);
nand U2453 (N_2453,N_2315,N_2342);
nand U2454 (N_2454,N_2331,N_2342);
or U2455 (N_2455,N_2371,N_2311);
or U2456 (N_2456,N_2309,N_2322);
or U2457 (N_2457,N_2306,N_2302);
or U2458 (N_2458,N_2368,N_2354);
nor U2459 (N_2459,N_2398,N_2368);
and U2460 (N_2460,N_2307,N_2368);
and U2461 (N_2461,N_2346,N_2377);
nor U2462 (N_2462,N_2391,N_2341);
nor U2463 (N_2463,N_2378,N_2325);
nor U2464 (N_2464,N_2312,N_2311);
nand U2465 (N_2465,N_2385,N_2390);
or U2466 (N_2466,N_2373,N_2379);
or U2467 (N_2467,N_2351,N_2310);
xnor U2468 (N_2468,N_2337,N_2370);
nor U2469 (N_2469,N_2338,N_2385);
or U2470 (N_2470,N_2388,N_2379);
or U2471 (N_2471,N_2320,N_2347);
nand U2472 (N_2472,N_2377,N_2313);
xnor U2473 (N_2473,N_2372,N_2351);
and U2474 (N_2474,N_2324,N_2367);
or U2475 (N_2475,N_2314,N_2362);
nor U2476 (N_2476,N_2379,N_2369);
or U2477 (N_2477,N_2365,N_2300);
xor U2478 (N_2478,N_2325,N_2353);
nor U2479 (N_2479,N_2355,N_2327);
nor U2480 (N_2480,N_2373,N_2388);
or U2481 (N_2481,N_2375,N_2347);
and U2482 (N_2482,N_2380,N_2365);
and U2483 (N_2483,N_2316,N_2343);
nand U2484 (N_2484,N_2321,N_2362);
and U2485 (N_2485,N_2371,N_2321);
nor U2486 (N_2486,N_2375,N_2323);
nor U2487 (N_2487,N_2343,N_2368);
nor U2488 (N_2488,N_2351,N_2369);
nand U2489 (N_2489,N_2328,N_2321);
nor U2490 (N_2490,N_2343,N_2397);
or U2491 (N_2491,N_2380,N_2399);
or U2492 (N_2492,N_2322,N_2362);
nor U2493 (N_2493,N_2374,N_2358);
nand U2494 (N_2494,N_2348,N_2321);
or U2495 (N_2495,N_2387,N_2300);
and U2496 (N_2496,N_2364,N_2388);
nand U2497 (N_2497,N_2340,N_2320);
and U2498 (N_2498,N_2311,N_2367);
or U2499 (N_2499,N_2387,N_2303);
or U2500 (N_2500,N_2463,N_2489);
or U2501 (N_2501,N_2421,N_2494);
nor U2502 (N_2502,N_2444,N_2441);
xor U2503 (N_2503,N_2453,N_2423);
and U2504 (N_2504,N_2499,N_2473);
xnor U2505 (N_2505,N_2480,N_2497);
nand U2506 (N_2506,N_2433,N_2440);
nand U2507 (N_2507,N_2483,N_2430);
nand U2508 (N_2508,N_2488,N_2446);
and U2509 (N_2509,N_2474,N_2486);
nor U2510 (N_2510,N_2451,N_2434);
nand U2511 (N_2511,N_2449,N_2475);
or U2512 (N_2512,N_2470,N_2407);
xnor U2513 (N_2513,N_2478,N_2448);
and U2514 (N_2514,N_2476,N_2471);
xor U2515 (N_2515,N_2435,N_2443);
or U2516 (N_2516,N_2415,N_2469);
nor U2517 (N_2517,N_2456,N_2481);
nand U2518 (N_2518,N_2418,N_2411);
nor U2519 (N_2519,N_2465,N_2436);
nor U2520 (N_2520,N_2439,N_2485);
or U2521 (N_2521,N_2419,N_2438);
nor U2522 (N_2522,N_2400,N_2424);
xnor U2523 (N_2523,N_2472,N_2468);
and U2524 (N_2524,N_2402,N_2461);
nand U2525 (N_2525,N_2409,N_2417);
xor U2526 (N_2526,N_2408,N_2445);
and U2527 (N_2527,N_2427,N_2492);
or U2528 (N_2528,N_2447,N_2425);
nor U2529 (N_2529,N_2413,N_2498);
nand U2530 (N_2530,N_2404,N_2490);
nor U2531 (N_2531,N_2477,N_2432);
and U2532 (N_2532,N_2403,N_2414);
nor U2533 (N_2533,N_2479,N_2457);
or U2534 (N_2534,N_2493,N_2455);
or U2535 (N_2535,N_2467,N_2452);
and U2536 (N_2536,N_2437,N_2462);
or U2537 (N_2537,N_2410,N_2450);
or U2538 (N_2538,N_2431,N_2406);
or U2539 (N_2539,N_2458,N_2495);
nor U2540 (N_2540,N_2428,N_2487);
nor U2541 (N_2541,N_2459,N_2416);
nand U2542 (N_2542,N_2496,N_2401);
xnor U2543 (N_2543,N_2429,N_2464);
nand U2544 (N_2544,N_2460,N_2426);
nor U2545 (N_2545,N_2412,N_2466);
nand U2546 (N_2546,N_2422,N_2442);
or U2547 (N_2547,N_2482,N_2484);
nand U2548 (N_2548,N_2405,N_2420);
and U2549 (N_2549,N_2454,N_2491);
nor U2550 (N_2550,N_2423,N_2408);
and U2551 (N_2551,N_2489,N_2473);
nand U2552 (N_2552,N_2442,N_2408);
nor U2553 (N_2553,N_2480,N_2430);
nor U2554 (N_2554,N_2459,N_2437);
and U2555 (N_2555,N_2445,N_2422);
nand U2556 (N_2556,N_2404,N_2425);
or U2557 (N_2557,N_2420,N_2409);
xnor U2558 (N_2558,N_2475,N_2422);
or U2559 (N_2559,N_2477,N_2461);
and U2560 (N_2560,N_2441,N_2488);
nand U2561 (N_2561,N_2498,N_2466);
and U2562 (N_2562,N_2414,N_2452);
xnor U2563 (N_2563,N_2435,N_2461);
and U2564 (N_2564,N_2415,N_2487);
nand U2565 (N_2565,N_2461,N_2407);
xnor U2566 (N_2566,N_2453,N_2426);
nor U2567 (N_2567,N_2416,N_2432);
and U2568 (N_2568,N_2403,N_2415);
nor U2569 (N_2569,N_2423,N_2431);
or U2570 (N_2570,N_2418,N_2402);
or U2571 (N_2571,N_2496,N_2473);
nor U2572 (N_2572,N_2482,N_2466);
nor U2573 (N_2573,N_2416,N_2465);
and U2574 (N_2574,N_2403,N_2496);
or U2575 (N_2575,N_2416,N_2435);
nand U2576 (N_2576,N_2462,N_2419);
and U2577 (N_2577,N_2476,N_2462);
and U2578 (N_2578,N_2460,N_2439);
xnor U2579 (N_2579,N_2458,N_2494);
and U2580 (N_2580,N_2429,N_2400);
and U2581 (N_2581,N_2481,N_2413);
and U2582 (N_2582,N_2450,N_2453);
nor U2583 (N_2583,N_2449,N_2429);
nand U2584 (N_2584,N_2406,N_2470);
or U2585 (N_2585,N_2437,N_2400);
nand U2586 (N_2586,N_2495,N_2451);
and U2587 (N_2587,N_2434,N_2405);
nand U2588 (N_2588,N_2445,N_2480);
nand U2589 (N_2589,N_2411,N_2404);
nand U2590 (N_2590,N_2426,N_2428);
nor U2591 (N_2591,N_2437,N_2451);
and U2592 (N_2592,N_2450,N_2422);
and U2593 (N_2593,N_2452,N_2426);
or U2594 (N_2594,N_2458,N_2497);
and U2595 (N_2595,N_2449,N_2430);
and U2596 (N_2596,N_2497,N_2447);
and U2597 (N_2597,N_2448,N_2486);
or U2598 (N_2598,N_2438,N_2463);
or U2599 (N_2599,N_2468,N_2417);
nand U2600 (N_2600,N_2591,N_2539);
or U2601 (N_2601,N_2523,N_2573);
and U2602 (N_2602,N_2555,N_2524);
or U2603 (N_2603,N_2547,N_2537);
and U2604 (N_2604,N_2504,N_2503);
nor U2605 (N_2605,N_2592,N_2567);
nor U2606 (N_2606,N_2559,N_2540);
nor U2607 (N_2607,N_2560,N_2581);
nand U2608 (N_2608,N_2585,N_2561);
nand U2609 (N_2609,N_2557,N_2522);
or U2610 (N_2610,N_2502,N_2514);
and U2611 (N_2611,N_2530,N_2551);
or U2612 (N_2612,N_2593,N_2521);
xor U2613 (N_2613,N_2541,N_2511);
or U2614 (N_2614,N_2507,N_2509);
or U2615 (N_2615,N_2594,N_2572);
and U2616 (N_2616,N_2558,N_2534);
and U2617 (N_2617,N_2549,N_2583);
nor U2618 (N_2618,N_2579,N_2597);
nor U2619 (N_2619,N_2556,N_2535);
xnor U2620 (N_2620,N_2562,N_2518);
nand U2621 (N_2621,N_2505,N_2577);
or U2622 (N_2622,N_2515,N_2517);
or U2623 (N_2623,N_2506,N_2529);
nand U2624 (N_2624,N_2590,N_2595);
and U2625 (N_2625,N_2589,N_2516);
or U2626 (N_2626,N_2553,N_2565);
or U2627 (N_2627,N_2548,N_2576);
nand U2628 (N_2628,N_2520,N_2570);
and U2629 (N_2629,N_2546,N_2510);
or U2630 (N_2630,N_2525,N_2574);
or U2631 (N_2631,N_2588,N_2580);
xnor U2632 (N_2632,N_2545,N_2519);
nor U2633 (N_2633,N_2513,N_2533);
and U2634 (N_2634,N_2550,N_2532);
or U2635 (N_2635,N_2531,N_2586);
nor U2636 (N_2636,N_2575,N_2571);
and U2637 (N_2637,N_2528,N_2526);
and U2638 (N_2638,N_2500,N_2566);
xnor U2639 (N_2639,N_2598,N_2599);
xor U2640 (N_2640,N_2543,N_2564);
nor U2641 (N_2641,N_2501,N_2554);
and U2642 (N_2642,N_2578,N_2527);
nor U2643 (N_2643,N_2563,N_2552);
and U2644 (N_2644,N_2584,N_2508);
nor U2645 (N_2645,N_2544,N_2582);
and U2646 (N_2646,N_2587,N_2536);
or U2647 (N_2647,N_2568,N_2542);
nand U2648 (N_2648,N_2596,N_2538);
nand U2649 (N_2649,N_2512,N_2569);
and U2650 (N_2650,N_2583,N_2572);
nor U2651 (N_2651,N_2524,N_2503);
nor U2652 (N_2652,N_2568,N_2528);
xor U2653 (N_2653,N_2578,N_2563);
and U2654 (N_2654,N_2528,N_2548);
and U2655 (N_2655,N_2598,N_2533);
nand U2656 (N_2656,N_2507,N_2566);
or U2657 (N_2657,N_2599,N_2554);
and U2658 (N_2658,N_2564,N_2501);
xnor U2659 (N_2659,N_2547,N_2540);
and U2660 (N_2660,N_2555,N_2580);
nor U2661 (N_2661,N_2516,N_2500);
or U2662 (N_2662,N_2590,N_2530);
nand U2663 (N_2663,N_2518,N_2514);
or U2664 (N_2664,N_2570,N_2588);
nor U2665 (N_2665,N_2568,N_2565);
or U2666 (N_2666,N_2577,N_2565);
nand U2667 (N_2667,N_2538,N_2526);
or U2668 (N_2668,N_2599,N_2540);
nor U2669 (N_2669,N_2530,N_2525);
nand U2670 (N_2670,N_2565,N_2548);
or U2671 (N_2671,N_2511,N_2507);
or U2672 (N_2672,N_2501,N_2557);
or U2673 (N_2673,N_2567,N_2545);
and U2674 (N_2674,N_2518,N_2521);
and U2675 (N_2675,N_2520,N_2531);
or U2676 (N_2676,N_2506,N_2547);
nand U2677 (N_2677,N_2548,N_2593);
or U2678 (N_2678,N_2542,N_2545);
and U2679 (N_2679,N_2567,N_2500);
or U2680 (N_2680,N_2544,N_2534);
nor U2681 (N_2681,N_2588,N_2512);
and U2682 (N_2682,N_2579,N_2561);
nand U2683 (N_2683,N_2554,N_2538);
nand U2684 (N_2684,N_2597,N_2563);
xor U2685 (N_2685,N_2548,N_2573);
or U2686 (N_2686,N_2562,N_2551);
nand U2687 (N_2687,N_2512,N_2547);
xor U2688 (N_2688,N_2590,N_2532);
nand U2689 (N_2689,N_2565,N_2575);
or U2690 (N_2690,N_2523,N_2506);
and U2691 (N_2691,N_2541,N_2571);
nand U2692 (N_2692,N_2522,N_2524);
or U2693 (N_2693,N_2560,N_2533);
nand U2694 (N_2694,N_2577,N_2541);
xnor U2695 (N_2695,N_2537,N_2589);
or U2696 (N_2696,N_2586,N_2500);
or U2697 (N_2697,N_2589,N_2535);
nand U2698 (N_2698,N_2540,N_2581);
or U2699 (N_2699,N_2539,N_2534);
and U2700 (N_2700,N_2694,N_2675);
nor U2701 (N_2701,N_2668,N_2631);
or U2702 (N_2702,N_2652,N_2655);
or U2703 (N_2703,N_2663,N_2618);
nor U2704 (N_2704,N_2621,N_2606);
and U2705 (N_2705,N_2678,N_2667);
nor U2706 (N_2706,N_2600,N_2684);
or U2707 (N_2707,N_2628,N_2697);
xnor U2708 (N_2708,N_2601,N_2645);
nand U2709 (N_2709,N_2613,N_2644);
or U2710 (N_2710,N_2633,N_2636);
nor U2711 (N_2711,N_2676,N_2669);
nand U2712 (N_2712,N_2620,N_2605);
xor U2713 (N_2713,N_2693,N_2680);
nand U2714 (N_2714,N_2674,N_2685);
xor U2715 (N_2715,N_2608,N_2673);
or U2716 (N_2716,N_2639,N_2687);
nand U2717 (N_2717,N_2607,N_2660);
and U2718 (N_2718,N_2683,N_2614);
or U2719 (N_2719,N_2696,N_2690);
and U2720 (N_2720,N_2666,N_2698);
or U2721 (N_2721,N_2659,N_2686);
nand U2722 (N_2722,N_2647,N_2637);
and U2723 (N_2723,N_2646,N_2612);
nor U2724 (N_2724,N_2615,N_2671);
or U2725 (N_2725,N_2692,N_2625);
or U2726 (N_2726,N_2661,N_2695);
nor U2727 (N_2727,N_2632,N_2677);
and U2728 (N_2728,N_2689,N_2616);
or U2729 (N_2729,N_2650,N_2624);
xor U2730 (N_2730,N_2649,N_2609);
nor U2731 (N_2731,N_2688,N_2623);
nand U2732 (N_2732,N_2657,N_2626);
nor U2733 (N_2733,N_2619,N_2662);
nor U2734 (N_2734,N_2658,N_2653);
xnor U2735 (N_2735,N_2638,N_2665);
nor U2736 (N_2736,N_2682,N_2611);
xor U2737 (N_2737,N_2656,N_2640);
nor U2738 (N_2738,N_2699,N_2681);
nor U2739 (N_2739,N_2654,N_2691);
and U2740 (N_2740,N_2602,N_2627);
or U2741 (N_2741,N_2648,N_2622);
xnor U2742 (N_2742,N_2617,N_2634);
xnor U2743 (N_2743,N_2672,N_2641);
nor U2744 (N_2744,N_2642,N_2651);
or U2745 (N_2745,N_2643,N_2629);
or U2746 (N_2746,N_2664,N_2679);
nand U2747 (N_2747,N_2604,N_2630);
nand U2748 (N_2748,N_2670,N_2610);
nor U2749 (N_2749,N_2635,N_2603);
xor U2750 (N_2750,N_2637,N_2692);
nand U2751 (N_2751,N_2667,N_2657);
or U2752 (N_2752,N_2601,N_2620);
nor U2753 (N_2753,N_2617,N_2627);
and U2754 (N_2754,N_2630,N_2655);
nor U2755 (N_2755,N_2694,N_2614);
nand U2756 (N_2756,N_2688,N_2600);
and U2757 (N_2757,N_2644,N_2678);
or U2758 (N_2758,N_2623,N_2603);
nor U2759 (N_2759,N_2636,N_2666);
and U2760 (N_2760,N_2620,N_2655);
xnor U2761 (N_2761,N_2678,N_2638);
and U2762 (N_2762,N_2621,N_2636);
and U2763 (N_2763,N_2659,N_2661);
nand U2764 (N_2764,N_2684,N_2612);
or U2765 (N_2765,N_2661,N_2656);
nor U2766 (N_2766,N_2600,N_2665);
nor U2767 (N_2767,N_2689,N_2629);
and U2768 (N_2768,N_2602,N_2657);
nand U2769 (N_2769,N_2637,N_2620);
nor U2770 (N_2770,N_2685,N_2681);
nand U2771 (N_2771,N_2650,N_2644);
xnor U2772 (N_2772,N_2650,N_2684);
nor U2773 (N_2773,N_2625,N_2697);
nor U2774 (N_2774,N_2600,N_2663);
or U2775 (N_2775,N_2631,N_2603);
nor U2776 (N_2776,N_2612,N_2629);
and U2777 (N_2777,N_2683,N_2633);
nand U2778 (N_2778,N_2680,N_2661);
nand U2779 (N_2779,N_2612,N_2623);
or U2780 (N_2780,N_2609,N_2627);
or U2781 (N_2781,N_2673,N_2604);
or U2782 (N_2782,N_2673,N_2695);
nand U2783 (N_2783,N_2601,N_2608);
nand U2784 (N_2784,N_2630,N_2676);
nor U2785 (N_2785,N_2660,N_2667);
xnor U2786 (N_2786,N_2652,N_2673);
nand U2787 (N_2787,N_2694,N_2648);
nor U2788 (N_2788,N_2658,N_2659);
nand U2789 (N_2789,N_2690,N_2666);
nor U2790 (N_2790,N_2619,N_2614);
xor U2791 (N_2791,N_2661,N_2626);
or U2792 (N_2792,N_2643,N_2630);
nand U2793 (N_2793,N_2668,N_2678);
nand U2794 (N_2794,N_2654,N_2612);
or U2795 (N_2795,N_2648,N_2640);
and U2796 (N_2796,N_2689,N_2603);
nor U2797 (N_2797,N_2650,N_2699);
nand U2798 (N_2798,N_2670,N_2628);
nor U2799 (N_2799,N_2622,N_2669);
nor U2800 (N_2800,N_2781,N_2744);
nand U2801 (N_2801,N_2796,N_2749);
and U2802 (N_2802,N_2748,N_2773);
and U2803 (N_2803,N_2731,N_2784);
and U2804 (N_2804,N_2750,N_2793);
nor U2805 (N_2805,N_2715,N_2762);
and U2806 (N_2806,N_2797,N_2764);
xor U2807 (N_2807,N_2724,N_2725);
or U2808 (N_2808,N_2766,N_2734);
and U2809 (N_2809,N_2794,N_2702);
and U2810 (N_2810,N_2712,N_2701);
nor U2811 (N_2811,N_2765,N_2758);
or U2812 (N_2812,N_2798,N_2710);
or U2813 (N_2813,N_2775,N_2787);
nor U2814 (N_2814,N_2771,N_2769);
and U2815 (N_2815,N_2738,N_2780);
and U2816 (N_2816,N_2791,N_2768);
and U2817 (N_2817,N_2760,N_2792);
or U2818 (N_2818,N_2753,N_2782);
and U2819 (N_2819,N_2703,N_2717);
or U2820 (N_2820,N_2726,N_2776);
xor U2821 (N_2821,N_2763,N_2785);
and U2822 (N_2822,N_2790,N_2718);
or U2823 (N_2823,N_2745,N_2779);
or U2824 (N_2824,N_2737,N_2729);
nor U2825 (N_2825,N_2789,N_2786);
nor U2826 (N_2826,N_2774,N_2728);
and U2827 (N_2827,N_2740,N_2727);
xor U2828 (N_2828,N_2709,N_2742);
nor U2829 (N_2829,N_2770,N_2711);
nor U2830 (N_2830,N_2708,N_2759);
xnor U2831 (N_2831,N_2700,N_2714);
nor U2832 (N_2832,N_2722,N_2747);
or U2833 (N_2833,N_2739,N_2755);
nor U2834 (N_2834,N_2772,N_2777);
nand U2835 (N_2835,N_2733,N_2795);
xnor U2836 (N_2836,N_2713,N_2721);
xor U2837 (N_2837,N_2732,N_2723);
nand U2838 (N_2838,N_2743,N_2783);
and U2839 (N_2839,N_2757,N_2741);
nand U2840 (N_2840,N_2767,N_2799);
or U2841 (N_2841,N_2730,N_2707);
or U2842 (N_2842,N_2788,N_2752);
or U2843 (N_2843,N_2761,N_2756);
nor U2844 (N_2844,N_2704,N_2736);
or U2845 (N_2845,N_2735,N_2706);
nor U2846 (N_2846,N_2716,N_2705);
xor U2847 (N_2847,N_2751,N_2754);
or U2848 (N_2848,N_2719,N_2778);
xor U2849 (N_2849,N_2746,N_2720);
nor U2850 (N_2850,N_2764,N_2794);
nor U2851 (N_2851,N_2703,N_2791);
nand U2852 (N_2852,N_2713,N_2788);
or U2853 (N_2853,N_2789,N_2702);
nand U2854 (N_2854,N_2776,N_2789);
nor U2855 (N_2855,N_2718,N_2716);
nor U2856 (N_2856,N_2771,N_2779);
nor U2857 (N_2857,N_2728,N_2705);
nor U2858 (N_2858,N_2728,N_2722);
or U2859 (N_2859,N_2706,N_2702);
nor U2860 (N_2860,N_2756,N_2734);
xnor U2861 (N_2861,N_2730,N_2797);
or U2862 (N_2862,N_2772,N_2779);
and U2863 (N_2863,N_2780,N_2712);
or U2864 (N_2864,N_2766,N_2747);
nand U2865 (N_2865,N_2741,N_2709);
nor U2866 (N_2866,N_2761,N_2703);
and U2867 (N_2867,N_2726,N_2779);
nor U2868 (N_2868,N_2772,N_2762);
and U2869 (N_2869,N_2714,N_2772);
nor U2870 (N_2870,N_2752,N_2726);
xor U2871 (N_2871,N_2793,N_2714);
nand U2872 (N_2872,N_2747,N_2742);
nor U2873 (N_2873,N_2755,N_2783);
nor U2874 (N_2874,N_2731,N_2799);
nor U2875 (N_2875,N_2773,N_2707);
and U2876 (N_2876,N_2757,N_2795);
or U2877 (N_2877,N_2784,N_2768);
nand U2878 (N_2878,N_2727,N_2719);
or U2879 (N_2879,N_2777,N_2783);
nand U2880 (N_2880,N_2730,N_2712);
xor U2881 (N_2881,N_2723,N_2730);
xnor U2882 (N_2882,N_2721,N_2756);
and U2883 (N_2883,N_2718,N_2759);
xnor U2884 (N_2884,N_2798,N_2722);
and U2885 (N_2885,N_2754,N_2762);
or U2886 (N_2886,N_2700,N_2750);
nor U2887 (N_2887,N_2773,N_2737);
nand U2888 (N_2888,N_2795,N_2779);
nand U2889 (N_2889,N_2764,N_2708);
nor U2890 (N_2890,N_2744,N_2768);
and U2891 (N_2891,N_2743,N_2764);
or U2892 (N_2892,N_2737,N_2772);
nor U2893 (N_2893,N_2767,N_2778);
or U2894 (N_2894,N_2717,N_2720);
nor U2895 (N_2895,N_2786,N_2709);
nand U2896 (N_2896,N_2796,N_2773);
xnor U2897 (N_2897,N_2780,N_2719);
or U2898 (N_2898,N_2751,N_2776);
nand U2899 (N_2899,N_2781,N_2751);
and U2900 (N_2900,N_2816,N_2893);
or U2901 (N_2901,N_2886,N_2847);
xor U2902 (N_2902,N_2889,N_2875);
and U2903 (N_2903,N_2824,N_2872);
or U2904 (N_2904,N_2856,N_2869);
or U2905 (N_2905,N_2863,N_2867);
or U2906 (N_2906,N_2838,N_2835);
and U2907 (N_2907,N_2873,N_2853);
nor U2908 (N_2908,N_2864,N_2888);
xor U2909 (N_2909,N_2859,N_2841);
nand U2910 (N_2910,N_2866,N_2832);
or U2911 (N_2911,N_2865,N_2807);
nand U2912 (N_2912,N_2879,N_2897);
nor U2913 (N_2913,N_2833,N_2858);
xnor U2914 (N_2914,N_2837,N_2850);
nor U2915 (N_2915,N_2899,N_2870);
nor U2916 (N_2916,N_2822,N_2878);
nand U2917 (N_2917,N_2840,N_2823);
nand U2918 (N_2918,N_2874,N_2855);
nand U2919 (N_2919,N_2880,N_2882);
and U2920 (N_2920,N_2806,N_2877);
nand U2921 (N_2921,N_2817,N_2808);
nand U2922 (N_2922,N_2842,N_2839);
nor U2923 (N_2923,N_2827,N_2881);
or U2924 (N_2924,N_2814,N_2868);
or U2925 (N_2925,N_2885,N_2845);
and U2926 (N_2926,N_2819,N_2815);
nand U2927 (N_2927,N_2896,N_2854);
xnor U2928 (N_2928,N_2829,N_2860);
nor U2929 (N_2929,N_2834,N_2801);
nand U2930 (N_2930,N_2828,N_2821);
or U2931 (N_2931,N_2862,N_2800);
xor U2932 (N_2932,N_2805,N_2846);
nand U2933 (N_2933,N_2887,N_2843);
and U2934 (N_2934,N_2809,N_2810);
nand U2935 (N_2935,N_2803,N_2883);
nand U2936 (N_2936,N_2890,N_2830);
nand U2937 (N_2937,N_2825,N_2876);
nor U2938 (N_2938,N_2894,N_2861);
nand U2939 (N_2939,N_2826,N_2871);
and U2940 (N_2940,N_2802,N_2820);
xor U2941 (N_2941,N_2848,N_2812);
or U2942 (N_2942,N_2844,N_2811);
nand U2943 (N_2943,N_2857,N_2895);
nor U2944 (N_2944,N_2892,N_2836);
and U2945 (N_2945,N_2813,N_2804);
and U2946 (N_2946,N_2852,N_2831);
nor U2947 (N_2947,N_2898,N_2851);
nor U2948 (N_2948,N_2891,N_2884);
nor U2949 (N_2949,N_2818,N_2849);
or U2950 (N_2950,N_2878,N_2823);
and U2951 (N_2951,N_2815,N_2848);
or U2952 (N_2952,N_2856,N_2895);
nand U2953 (N_2953,N_2811,N_2865);
and U2954 (N_2954,N_2879,N_2865);
and U2955 (N_2955,N_2839,N_2848);
nor U2956 (N_2956,N_2805,N_2882);
or U2957 (N_2957,N_2804,N_2817);
nor U2958 (N_2958,N_2879,N_2857);
nor U2959 (N_2959,N_2892,N_2852);
nor U2960 (N_2960,N_2840,N_2865);
nor U2961 (N_2961,N_2821,N_2806);
nor U2962 (N_2962,N_2862,N_2804);
nor U2963 (N_2963,N_2845,N_2877);
or U2964 (N_2964,N_2853,N_2875);
xnor U2965 (N_2965,N_2868,N_2888);
nor U2966 (N_2966,N_2835,N_2819);
or U2967 (N_2967,N_2874,N_2804);
and U2968 (N_2968,N_2879,N_2803);
nor U2969 (N_2969,N_2826,N_2844);
xor U2970 (N_2970,N_2846,N_2876);
or U2971 (N_2971,N_2898,N_2860);
nand U2972 (N_2972,N_2819,N_2870);
and U2973 (N_2973,N_2847,N_2863);
and U2974 (N_2974,N_2855,N_2890);
nand U2975 (N_2975,N_2861,N_2868);
and U2976 (N_2976,N_2820,N_2807);
or U2977 (N_2977,N_2878,N_2866);
or U2978 (N_2978,N_2896,N_2897);
and U2979 (N_2979,N_2805,N_2872);
or U2980 (N_2980,N_2835,N_2878);
or U2981 (N_2981,N_2819,N_2881);
nand U2982 (N_2982,N_2880,N_2806);
nand U2983 (N_2983,N_2826,N_2831);
and U2984 (N_2984,N_2851,N_2840);
nor U2985 (N_2985,N_2806,N_2828);
nand U2986 (N_2986,N_2884,N_2811);
nor U2987 (N_2987,N_2803,N_2898);
nand U2988 (N_2988,N_2862,N_2838);
nand U2989 (N_2989,N_2845,N_2881);
nor U2990 (N_2990,N_2876,N_2809);
nand U2991 (N_2991,N_2879,N_2848);
or U2992 (N_2992,N_2859,N_2865);
and U2993 (N_2993,N_2875,N_2818);
or U2994 (N_2994,N_2857,N_2843);
and U2995 (N_2995,N_2815,N_2856);
xnor U2996 (N_2996,N_2891,N_2871);
nor U2997 (N_2997,N_2843,N_2813);
nand U2998 (N_2998,N_2812,N_2819);
xnor U2999 (N_2999,N_2864,N_2831);
nand UO_0 (O_0,N_2970,N_2902);
and UO_1 (O_1,N_2954,N_2939);
nand UO_2 (O_2,N_2967,N_2955);
and UO_3 (O_3,N_2977,N_2992);
and UO_4 (O_4,N_2986,N_2972);
nor UO_5 (O_5,N_2926,N_2982);
and UO_6 (O_6,N_2931,N_2969);
nand UO_7 (O_7,N_2958,N_2973);
or UO_8 (O_8,N_2976,N_2963);
nand UO_9 (O_9,N_2984,N_2929);
nor UO_10 (O_10,N_2971,N_2925);
nand UO_11 (O_11,N_2993,N_2946);
nor UO_12 (O_12,N_2900,N_2983);
nor UO_13 (O_13,N_2951,N_2980);
nor UO_14 (O_14,N_2942,N_2943);
and UO_15 (O_15,N_2957,N_2913);
nand UO_16 (O_16,N_2948,N_2910);
nor UO_17 (O_17,N_2906,N_2932);
nor UO_18 (O_18,N_2994,N_2999);
or UO_19 (O_19,N_2914,N_2949);
and UO_20 (O_20,N_2921,N_2919);
nand UO_21 (O_21,N_2978,N_2947);
or UO_22 (O_22,N_2997,N_2924);
nor UO_23 (O_23,N_2933,N_2920);
nor UO_24 (O_24,N_2908,N_2915);
nand UO_25 (O_25,N_2998,N_2991);
and UO_26 (O_26,N_2944,N_2912);
nand UO_27 (O_27,N_2918,N_2968);
nand UO_28 (O_28,N_2981,N_2960);
or UO_29 (O_29,N_2974,N_2916);
or UO_30 (O_30,N_2996,N_2904);
and UO_31 (O_31,N_2909,N_2953);
nor UO_32 (O_32,N_2917,N_2907);
nand UO_33 (O_33,N_2911,N_2935);
xnor UO_34 (O_34,N_2934,N_2961);
nor UO_35 (O_35,N_2985,N_2941);
and UO_36 (O_36,N_2930,N_2922);
or UO_37 (O_37,N_2956,N_2950);
and UO_38 (O_38,N_2965,N_2995);
nand UO_39 (O_39,N_2989,N_2927);
nand UO_40 (O_40,N_2964,N_2987);
nor UO_41 (O_41,N_2959,N_2979);
nor UO_42 (O_42,N_2962,N_2945);
and UO_43 (O_43,N_2966,N_2988);
and UO_44 (O_44,N_2937,N_2990);
nor UO_45 (O_45,N_2936,N_2938);
and UO_46 (O_46,N_2901,N_2940);
nor UO_47 (O_47,N_2975,N_2952);
xor UO_48 (O_48,N_2928,N_2923);
or UO_49 (O_49,N_2905,N_2903);
and UO_50 (O_50,N_2907,N_2969);
nor UO_51 (O_51,N_2904,N_2927);
nand UO_52 (O_52,N_2917,N_2987);
nand UO_53 (O_53,N_2968,N_2948);
nand UO_54 (O_54,N_2985,N_2971);
or UO_55 (O_55,N_2953,N_2960);
or UO_56 (O_56,N_2917,N_2989);
nor UO_57 (O_57,N_2966,N_2935);
nand UO_58 (O_58,N_2950,N_2973);
or UO_59 (O_59,N_2912,N_2942);
nor UO_60 (O_60,N_2999,N_2955);
nor UO_61 (O_61,N_2961,N_2958);
or UO_62 (O_62,N_2984,N_2925);
nor UO_63 (O_63,N_2945,N_2902);
xor UO_64 (O_64,N_2957,N_2998);
nor UO_65 (O_65,N_2916,N_2917);
nand UO_66 (O_66,N_2921,N_2938);
nand UO_67 (O_67,N_2957,N_2964);
nor UO_68 (O_68,N_2966,N_2932);
xnor UO_69 (O_69,N_2958,N_2978);
and UO_70 (O_70,N_2918,N_2987);
and UO_71 (O_71,N_2948,N_2916);
nor UO_72 (O_72,N_2900,N_2984);
and UO_73 (O_73,N_2965,N_2979);
nand UO_74 (O_74,N_2920,N_2949);
nand UO_75 (O_75,N_2910,N_2913);
and UO_76 (O_76,N_2921,N_2900);
nand UO_77 (O_77,N_2942,N_2926);
and UO_78 (O_78,N_2929,N_2926);
nor UO_79 (O_79,N_2998,N_2917);
nor UO_80 (O_80,N_2992,N_2947);
or UO_81 (O_81,N_2973,N_2913);
xor UO_82 (O_82,N_2936,N_2978);
nand UO_83 (O_83,N_2923,N_2918);
and UO_84 (O_84,N_2962,N_2984);
or UO_85 (O_85,N_2924,N_2982);
xor UO_86 (O_86,N_2956,N_2932);
and UO_87 (O_87,N_2949,N_2958);
or UO_88 (O_88,N_2942,N_2976);
or UO_89 (O_89,N_2930,N_2967);
and UO_90 (O_90,N_2935,N_2942);
nand UO_91 (O_91,N_2917,N_2976);
or UO_92 (O_92,N_2923,N_2903);
nand UO_93 (O_93,N_2975,N_2969);
xor UO_94 (O_94,N_2931,N_2974);
or UO_95 (O_95,N_2900,N_2978);
or UO_96 (O_96,N_2973,N_2949);
nor UO_97 (O_97,N_2983,N_2960);
and UO_98 (O_98,N_2960,N_2906);
and UO_99 (O_99,N_2906,N_2946);
or UO_100 (O_100,N_2940,N_2914);
or UO_101 (O_101,N_2933,N_2967);
and UO_102 (O_102,N_2941,N_2965);
nand UO_103 (O_103,N_2911,N_2943);
nand UO_104 (O_104,N_2972,N_2923);
nor UO_105 (O_105,N_2946,N_2977);
nor UO_106 (O_106,N_2950,N_2909);
nor UO_107 (O_107,N_2972,N_2921);
xor UO_108 (O_108,N_2923,N_2956);
nor UO_109 (O_109,N_2949,N_2976);
nand UO_110 (O_110,N_2914,N_2969);
nand UO_111 (O_111,N_2992,N_2955);
nand UO_112 (O_112,N_2990,N_2942);
and UO_113 (O_113,N_2971,N_2909);
and UO_114 (O_114,N_2932,N_2980);
or UO_115 (O_115,N_2997,N_2983);
or UO_116 (O_116,N_2960,N_2924);
nor UO_117 (O_117,N_2995,N_2907);
or UO_118 (O_118,N_2932,N_2936);
or UO_119 (O_119,N_2933,N_2984);
nor UO_120 (O_120,N_2992,N_2971);
or UO_121 (O_121,N_2945,N_2984);
nor UO_122 (O_122,N_2901,N_2982);
or UO_123 (O_123,N_2968,N_2915);
nand UO_124 (O_124,N_2918,N_2912);
or UO_125 (O_125,N_2990,N_2970);
or UO_126 (O_126,N_2991,N_2914);
or UO_127 (O_127,N_2961,N_2935);
or UO_128 (O_128,N_2978,N_2992);
xnor UO_129 (O_129,N_2995,N_2968);
nor UO_130 (O_130,N_2928,N_2991);
or UO_131 (O_131,N_2921,N_2946);
nand UO_132 (O_132,N_2968,N_2965);
nor UO_133 (O_133,N_2910,N_2901);
nor UO_134 (O_134,N_2920,N_2936);
and UO_135 (O_135,N_2993,N_2919);
and UO_136 (O_136,N_2930,N_2993);
and UO_137 (O_137,N_2980,N_2931);
and UO_138 (O_138,N_2916,N_2956);
and UO_139 (O_139,N_2966,N_2954);
nand UO_140 (O_140,N_2992,N_2943);
nor UO_141 (O_141,N_2957,N_2926);
or UO_142 (O_142,N_2964,N_2991);
and UO_143 (O_143,N_2960,N_2980);
nand UO_144 (O_144,N_2900,N_2908);
nor UO_145 (O_145,N_2973,N_2934);
and UO_146 (O_146,N_2913,N_2962);
and UO_147 (O_147,N_2955,N_2909);
and UO_148 (O_148,N_2983,N_2905);
nor UO_149 (O_149,N_2917,N_2959);
and UO_150 (O_150,N_2916,N_2965);
nor UO_151 (O_151,N_2924,N_2974);
nand UO_152 (O_152,N_2931,N_2973);
or UO_153 (O_153,N_2975,N_2970);
nor UO_154 (O_154,N_2958,N_2924);
or UO_155 (O_155,N_2954,N_2920);
nor UO_156 (O_156,N_2928,N_2907);
or UO_157 (O_157,N_2918,N_2917);
or UO_158 (O_158,N_2991,N_2924);
nand UO_159 (O_159,N_2991,N_2980);
nor UO_160 (O_160,N_2928,N_2946);
or UO_161 (O_161,N_2924,N_2948);
or UO_162 (O_162,N_2970,N_2979);
xnor UO_163 (O_163,N_2904,N_2969);
nor UO_164 (O_164,N_2928,N_2902);
nand UO_165 (O_165,N_2909,N_2923);
and UO_166 (O_166,N_2905,N_2924);
nor UO_167 (O_167,N_2943,N_2931);
and UO_168 (O_168,N_2959,N_2934);
and UO_169 (O_169,N_2927,N_2916);
nand UO_170 (O_170,N_2913,N_2982);
or UO_171 (O_171,N_2943,N_2988);
nand UO_172 (O_172,N_2935,N_2946);
nor UO_173 (O_173,N_2992,N_2942);
and UO_174 (O_174,N_2946,N_2974);
nand UO_175 (O_175,N_2961,N_2988);
and UO_176 (O_176,N_2968,N_2914);
nor UO_177 (O_177,N_2986,N_2916);
nor UO_178 (O_178,N_2967,N_2983);
nor UO_179 (O_179,N_2977,N_2924);
and UO_180 (O_180,N_2947,N_2998);
nand UO_181 (O_181,N_2978,N_2956);
or UO_182 (O_182,N_2989,N_2949);
or UO_183 (O_183,N_2963,N_2936);
nor UO_184 (O_184,N_2983,N_2974);
or UO_185 (O_185,N_2940,N_2906);
and UO_186 (O_186,N_2900,N_2925);
nand UO_187 (O_187,N_2967,N_2974);
nor UO_188 (O_188,N_2939,N_2950);
nor UO_189 (O_189,N_2961,N_2950);
nand UO_190 (O_190,N_2970,N_2988);
nand UO_191 (O_191,N_2972,N_2968);
nand UO_192 (O_192,N_2907,N_2956);
nand UO_193 (O_193,N_2975,N_2964);
and UO_194 (O_194,N_2910,N_2926);
nor UO_195 (O_195,N_2904,N_2966);
and UO_196 (O_196,N_2917,N_2932);
and UO_197 (O_197,N_2999,N_2907);
and UO_198 (O_198,N_2972,N_2904);
or UO_199 (O_199,N_2996,N_2987);
or UO_200 (O_200,N_2939,N_2942);
and UO_201 (O_201,N_2927,N_2939);
or UO_202 (O_202,N_2911,N_2903);
nor UO_203 (O_203,N_2941,N_2994);
or UO_204 (O_204,N_2948,N_2953);
xor UO_205 (O_205,N_2971,N_2977);
nand UO_206 (O_206,N_2924,N_2919);
nor UO_207 (O_207,N_2975,N_2974);
nor UO_208 (O_208,N_2912,N_2923);
or UO_209 (O_209,N_2950,N_2945);
nand UO_210 (O_210,N_2925,N_2933);
xor UO_211 (O_211,N_2924,N_2901);
or UO_212 (O_212,N_2972,N_2943);
nor UO_213 (O_213,N_2958,N_2930);
and UO_214 (O_214,N_2912,N_2965);
nand UO_215 (O_215,N_2938,N_2946);
or UO_216 (O_216,N_2938,N_2952);
and UO_217 (O_217,N_2963,N_2926);
nand UO_218 (O_218,N_2931,N_2952);
nand UO_219 (O_219,N_2944,N_2968);
nand UO_220 (O_220,N_2905,N_2950);
and UO_221 (O_221,N_2918,N_2949);
and UO_222 (O_222,N_2907,N_2980);
nand UO_223 (O_223,N_2958,N_2922);
nand UO_224 (O_224,N_2902,N_2967);
or UO_225 (O_225,N_2987,N_2961);
and UO_226 (O_226,N_2954,N_2913);
nor UO_227 (O_227,N_2908,N_2936);
nor UO_228 (O_228,N_2970,N_2994);
or UO_229 (O_229,N_2955,N_2964);
nor UO_230 (O_230,N_2974,N_2962);
and UO_231 (O_231,N_2938,N_2904);
nor UO_232 (O_232,N_2900,N_2957);
or UO_233 (O_233,N_2977,N_2901);
or UO_234 (O_234,N_2982,N_2909);
nor UO_235 (O_235,N_2995,N_2940);
and UO_236 (O_236,N_2968,N_2947);
and UO_237 (O_237,N_2992,N_2975);
nor UO_238 (O_238,N_2901,N_2980);
nand UO_239 (O_239,N_2960,N_2951);
or UO_240 (O_240,N_2914,N_2925);
xnor UO_241 (O_241,N_2962,N_2977);
nand UO_242 (O_242,N_2990,N_2980);
or UO_243 (O_243,N_2916,N_2926);
nor UO_244 (O_244,N_2994,N_2945);
and UO_245 (O_245,N_2900,N_2901);
xnor UO_246 (O_246,N_2933,N_2945);
nor UO_247 (O_247,N_2970,N_2993);
and UO_248 (O_248,N_2955,N_2927);
or UO_249 (O_249,N_2927,N_2962);
and UO_250 (O_250,N_2904,N_2915);
and UO_251 (O_251,N_2983,N_2912);
nand UO_252 (O_252,N_2966,N_2959);
or UO_253 (O_253,N_2942,N_2916);
nor UO_254 (O_254,N_2979,N_2958);
and UO_255 (O_255,N_2929,N_2914);
and UO_256 (O_256,N_2985,N_2950);
and UO_257 (O_257,N_2919,N_2971);
and UO_258 (O_258,N_2963,N_2978);
nand UO_259 (O_259,N_2993,N_2999);
xnor UO_260 (O_260,N_2981,N_2924);
nor UO_261 (O_261,N_2905,N_2960);
nand UO_262 (O_262,N_2952,N_2922);
nand UO_263 (O_263,N_2920,N_2951);
nand UO_264 (O_264,N_2982,N_2984);
or UO_265 (O_265,N_2941,N_2968);
or UO_266 (O_266,N_2907,N_2950);
nand UO_267 (O_267,N_2926,N_2993);
or UO_268 (O_268,N_2992,N_2929);
xnor UO_269 (O_269,N_2986,N_2968);
nand UO_270 (O_270,N_2915,N_2943);
nand UO_271 (O_271,N_2958,N_2908);
nor UO_272 (O_272,N_2950,N_2974);
or UO_273 (O_273,N_2917,N_2968);
nor UO_274 (O_274,N_2911,N_2957);
and UO_275 (O_275,N_2964,N_2951);
and UO_276 (O_276,N_2901,N_2932);
and UO_277 (O_277,N_2966,N_2908);
and UO_278 (O_278,N_2933,N_2990);
nand UO_279 (O_279,N_2945,N_2959);
or UO_280 (O_280,N_2966,N_2980);
nor UO_281 (O_281,N_2909,N_2906);
nor UO_282 (O_282,N_2913,N_2914);
or UO_283 (O_283,N_2967,N_2912);
nand UO_284 (O_284,N_2997,N_2984);
nor UO_285 (O_285,N_2958,N_2959);
and UO_286 (O_286,N_2946,N_2954);
nand UO_287 (O_287,N_2904,N_2901);
nor UO_288 (O_288,N_2933,N_2946);
and UO_289 (O_289,N_2987,N_2903);
or UO_290 (O_290,N_2932,N_2907);
and UO_291 (O_291,N_2929,N_2941);
xnor UO_292 (O_292,N_2909,N_2916);
xnor UO_293 (O_293,N_2968,N_2950);
nand UO_294 (O_294,N_2925,N_2946);
and UO_295 (O_295,N_2918,N_2921);
or UO_296 (O_296,N_2959,N_2949);
nor UO_297 (O_297,N_2919,N_2966);
nor UO_298 (O_298,N_2952,N_2978);
xnor UO_299 (O_299,N_2913,N_2947);
nor UO_300 (O_300,N_2903,N_2927);
nand UO_301 (O_301,N_2957,N_2929);
nand UO_302 (O_302,N_2935,N_2996);
and UO_303 (O_303,N_2991,N_2919);
nor UO_304 (O_304,N_2981,N_2979);
nor UO_305 (O_305,N_2972,N_2909);
nand UO_306 (O_306,N_2976,N_2940);
nand UO_307 (O_307,N_2921,N_2937);
nor UO_308 (O_308,N_2938,N_2903);
nor UO_309 (O_309,N_2968,N_2997);
nand UO_310 (O_310,N_2982,N_2956);
nand UO_311 (O_311,N_2910,N_2969);
and UO_312 (O_312,N_2965,N_2958);
or UO_313 (O_313,N_2987,N_2963);
or UO_314 (O_314,N_2943,N_2965);
or UO_315 (O_315,N_2976,N_2945);
and UO_316 (O_316,N_2969,N_2979);
or UO_317 (O_317,N_2900,N_2916);
and UO_318 (O_318,N_2946,N_2947);
nor UO_319 (O_319,N_2959,N_2969);
or UO_320 (O_320,N_2949,N_2900);
nand UO_321 (O_321,N_2977,N_2916);
or UO_322 (O_322,N_2922,N_2957);
nor UO_323 (O_323,N_2970,N_2928);
xor UO_324 (O_324,N_2973,N_2924);
xor UO_325 (O_325,N_2937,N_2914);
nor UO_326 (O_326,N_2917,N_2996);
and UO_327 (O_327,N_2982,N_2949);
and UO_328 (O_328,N_2977,N_2989);
nand UO_329 (O_329,N_2932,N_2919);
nor UO_330 (O_330,N_2951,N_2962);
and UO_331 (O_331,N_2970,N_2918);
and UO_332 (O_332,N_2981,N_2938);
or UO_333 (O_333,N_2939,N_2956);
nor UO_334 (O_334,N_2985,N_2945);
nand UO_335 (O_335,N_2961,N_2984);
nand UO_336 (O_336,N_2960,N_2907);
xor UO_337 (O_337,N_2915,N_2998);
nor UO_338 (O_338,N_2914,N_2911);
or UO_339 (O_339,N_2914,N_2997);
nor UO_340 (O_340,N_2935,N_2988);
xnor UO_341 (O_341,N_2991,N_2911);
xor UO_342 (O_342,N_2931,N_2965);
nand UO_343 (O_343,N_2933,N_2951);
or UO_344 (O_344,N_2931,N_2977);
or UO_345 (O_345,N_2904,N_2958);
or UO_346 (O_346,N_2960,N_2989);
or UO_347 (O_347,N_2925,N_2905);
or UO_348 (O_348,N_2932,N_2991);
xnor UO_349 (O_349,N_2902,N_2976);
nor UO_350 (O_350,N_2930,N_2994);
or UO_351 (O_351,N_2995,N_2980);
xor UO_352 (O_352,N_2937,N_2952);
and UO_353 (O_353,N_2938,N_2996);
and UO_354 (O_354,N_2986,N_2998);
or UO_355 (O_355,N_2928,N_2978);
or UO_356 (O_356,N_2915,N_2900);
or UO_357 (O_357,N_2916,N_2907);
and UO_358 (O_358,N_2926,N_2906);
nand UO_359 (O_359,N_2936,N_2986);
or UO_360 (O_360,N_2965,N_2974);
nor UO_361 (O_361,N_2954,N_2911);
and UO_362 (O_362,N_2908,N_2918);
nand UO_363 (O_363,N_2956,N_2983);
xnor UO_364 (O_364,N_2970,N_2983);
nand UO_365 (O_365,N_2934,N_2944);
and UO_366 (O_366,N_2952,N_2924);
xnor UO_367 (O_367,N_2977,N_2943);
xnor UO_368 (O_368,N_2978,N_2999);
xnor UO_369 (O_369,N_2905,N_2972);
nand UO_370 (O_370,N_2936,N_2970);
xor UO_371 (O_371,N_2900,N_2967);
and UO_372 (O_372,N_2970,N_2933);
or UO_373 (O_373,N_2965,N_2956);
nand UO_374 (O_374,N_2952,N_2963);
and UO_375 (O_375,N_2920,N_2907);
nor UO_376 (O_376,N_2979,N_2921);
nand UO_377 (O_377,N_2939,N_2941);
nor UO_378 (O_378,N_2900,N_2905);
or UO_379 (O_379,N_2933,N_2987);
xnor UO_380 (O_380,N_2932,N_2986);
and UO_381 (O_381,N_2940,N_2939);
or UO_382 (O_382,N_2918,N_2910);
or UO_383 (O_383,N_2900,N_2911);
or UO_384 (O_384,N_2961,N_2974);
and UO_385 (O_385,N_2995,N_2993);
and UO_386 (O_386,N_2964,N_2925);
or UO_387 (O_387,N_2917,N_2978);
nand UO_388 (O_388,N_2905,N_2931);
xor UO_389 (O_389,N_2956,N_2970);
nor UO_390 (O_390,N_2956,N_2951);
nand UO_391 (O_391,N_2945,N_2907);
nand UO_392 (O_392,N_2907,N_2934);
nor UO_393 (O_393,N_2966,N_2939);
or UO_394 (O_394,N_2967,N_2938);
or UO_395 (O_395,N_2931,N_2910);
or UO_396 (O_396,N_2994,N_2981);
nor UO_397 (O_397,N_2971,N_2902);
or UO_398 (O_398,N_2967,N_2945);
or UO_399 (O_399,N_2960,N_2991);
nand UO_400 (O_400,N_2985,N_2948);
xnor UO_401 (O_401,N_2952,N_2989);
nand UO_402 (O_402,N_2929,N_2938);
or UO_403 (O_403,N_2950,N_2901);
nand UO_404 (O_404,N_2918,N_2939);
and UO_405 (O_405,N_2934,N_2949);
and UO_406 (O_406,N_2980,N_2944);
nor UO_407 (O_407,N_2964,N_2928);
or UO_408 (O_408,N_2998,N_2945);
and UO_409 (O_409,N_2968,N_2996);
or UO_410 (O_410,N_2944,N_2982);
or UO_411 (O_411,N_2968,N_2946);
or UO_412 (O_412,N_2923,N_2950);
nor UO_413 (O_413,N_2910,N_2934);
nand UO_414 (O_414,N_2920,N_2986);
or UO_415 (O_415,N_2939,N_2975);
and UO_416 (O_416,N_2976,N_2929);
or UO_417 (O_417,N_2914,N_2943);
or UO_418 (O_418,N_2925,N_2994);
nor UO_419 (O_419,N_2959,N_2923);
and UO_420 (O_420,N_2926,N_2966);
and UO_421 (O_421,N_2913,N_2920);
nand UO_422 (O_422,N_2946,N_2913);
and UO_423 (O_423,N_2964,N_2976);
and UO_424 (O_424,N_2930,N_2928);
nor UO_425 (O_425,N_2909,N_2949);
or UO_426 (O_426,N_2993,N_2940);
and UO_427 (O_427,N_2936,N_2979);
and UO_428 (O_428,N_2973,N_2962);
and UO_429 (O_429,N_2979,N_2984);
nor UO_430 (O_430,N_2960,N_2992);
or UO_431 (O_431,N_2985,N_2923);
xnor UO_432 (O_432,N_2940,N_2903);
nor UO_433 (O_433,N_2922,N_2920);
nor UO_434 (O_434,N_2928,N_2908);
or UO_435 (O_435,N_2971,N_2944);
or UO_436 (O_436,N_2929,N_2989);
xnor UO_437 (O_437,N_2903,N_2949);
or UO_438 (O_438,N_2980,N_2918);
nand UO_439 (O_439,N_2980,N_2976);
nand UO_440 (O_440,N_2987,N_2959);
or UO_441 (O_441,N_2946,N_2944);
and UO_442 (O_442,N_2931,N_2957);
nand UO_443 (O_443,N_2961,N_2928);
or UO_444 (O_444,N_2942,N_2940);
nand UO_445 (O_445,N_2912,N_2924);
or UO_446 (O_446,N_2928,N_2926);
nor UO_447 (O_447,N_2950,N_2967);
nor UO_448 (O_448,N_2925,N_2966);
and UO_449 (O_449,N_2933,N_2922);
and UO_450 (O_450,N_2905,N_2939);
or UO_451 (O_451,N_2943,N_2921);
nor UO_452 (O_452,N_2962,N_2948);
or UO_453 (O_453,N_2986,N_2988);
and UO_454 (O_454,N_2932,N_2971);
nand UO_455 (O_455,N_2916,N_2995);
nand UO_456 (O_456,N_2990,N_2947);
xor UO_457 (O_457,N_2995,N_2961);
nor UO_458 (O_458,N_2991,N_2921);
nand UO_459 (O_459,N_2940,N_2999);
nand UO_460 (O_460,N_2900,N_2910);
and UO_461 (O_461,N_2909,N_2933);
nand UO_462 (O_462,N_2929,N_2927);
nor UO_463 (O_463,N_2962,N_2905);
nand UO_464 (O_464,N_2902,N_2919);
and UO_465 (O_465,N_2972,N_2956);
nor UO_466 (O_466,N_2906,N_2983);
nand UO_467 (O_467,N_2945,N_2941);
nor UO_468 (O_468,N_2977,N_2900);
nand UO_469 (O_469,N_2987,N_2986);
or UO_470 (O_470,N_2908,N_2955);
xor UO_471 (O_471,N_2992,N_2963);
xnor UO_472 (O_472,N_2938,N_2998);
or UO_473 (O_473,N_2998,N_2977);
nand UO_474 (O_474,N_2939,N_2919);
or UO_475 (O_475,N_2944,N_2958);
and UO_476 (O_476,N_2916,N_2921);
nand UO_477 (O_477,N_2960,N_2927);
nor UO_478 (O_478,N_2990,N_2908);
and UO_479 (O_479,N_2943,N_2999);
or UO_480 (O_480,N_2983,N_2952);
nand UO_481 (O_481,N_2990,N_2977);
nand UO_482 (O_482,N_2995,N_2905);
nor UO_483 (O_483,N_2928,N_2916);
and UO_484 (O_484,N_2958,N_2974);
nor UO_485 (O_485,N_2934,N_2939);
xnor UO_486 (O_486,N_2953,N_2989);
or UO_487 (O_487,N_2903,N_2919);
nor UO_488 (O_488,N_2957,N_2944);
or UO_489 (O_489,N_2998,N_2987);
nor UO_490 (O_490,N_2922,N_2941);
nand UO_491 (O_491,N_2903,N_2910);
nor UO_492 (O_492,N_2914,N_2988);
or UO_493 (O_493,N_2926,N_2977);
or UO_494 (O_494,N_2983,N_2922);
nor UO_495 (O_495,N_2991,N_2982);
and UO_496 (O_496,N_2912,N_2976);
nand UO_497 (O_497,N_2955,N_2985);
nand UO_498 (O_498,N_2935,N_2948);
nand UO_499 (O_499,N_2968,N_2911);
endmodule