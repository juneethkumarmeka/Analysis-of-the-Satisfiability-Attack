module basic_2000_20000_2500_125_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_1124,In_88);
nand U1 (N_1,In_107,In_1199);
nor U2 (N_2,In_457,In_1262);
xor U3 (N_3,In_1518,In_335);
xor U4 (N_4,In_917,In_329);
nor U5 (N_5,In_161,In_634);
nand U6 (N_6,In_1,In_754);
and U7 (N_7,In_652,In_228);
nand U8 (N_8,In_1464,In_940);
or U9 (N_9,In_1070,In_56);
nor U10 (N_10,In_1308,In_1782);
or U11 (N_11,In_1783,In_784);
or U12 (N_12,In_1526,In_1077);
xnor U13 (N_13,In_23,In_909);
nor U14 (N_14,In_958,In_1395);
nand U15 (N_15,In_355,In_1964);
xor U16 (N_16,In_362,In_226);
and U17 (N_17,In_1313,In_404);
nand U18 (N_18,In_912,In_1867);
or U19 (N_19,In_1791,In_1509);
nand U20 (N_20,In_64,In_955);
nor U21 (N_21,In_207,In_1855);
nor U22 (N_22,In_734,In_1127);
and U23 (N_23,In_1414,In_1546);
or U24 (N_24,In_910,In_1117);
xnor U25 (N_25,In_735,In_243);
and U26 (N_26,In_129,In_898);
nand U27 (N_27,In_126,In_1829);
or U28 (N_28,In_1762,In_792);
and U29 (N_29,In_371,In_302);
or U30 (N_30,In_1008,In_1873);
and U31 (N_31,In_514,In_655);
nor U32 (N_32,In_264,In_1358);
xnor U33 (N_33,In_1031,In_320);
nand U34 (N_34,In_163,In_1667);
nand U35 (N_35,In_221,In_767);
and U36 (N_36,In_643,In_1610);
xor U37 (N_37,In_1534,In_1214);
xnor U38 (N_38,In_1076,In_1251);
nand U39 (N_39,In_990,In_595);
or U40 (N_40,In_262,In_706);
xnor U41 (N_41,In_540,In_1084);
or U42 (N_42,In_1805,In_1780);
nand U43 (N_43,In_446,In_1836);
or U44 (N_44,In_560,In_114);
nor U45 (N_45,In_1774,In_988);
or U46 (N_46,In_775,In_1926);
xor U47 (N_47,In_1682,In_1496);
and U48 (N_48,In_469,In_1644);
and U49 (N_49,In_1955,In_997);
nand U50 (N_50,In_290,In_1068);
nor U51 (N_51,In_1156,In_1179);
and U52 (N_52,In_1723,In_1589);
nand U53 (N_53,In_478,In_1275);
and U54 (N_54,In_47,In_1286);
nor U55 (N_55,In_144,In_1093);
nor U56 (N_56,In_1029,In_1011);
and U57 (N_57,In_570,In_1971);
and U58 (N_58,In_1298,In_1902);
and U59 (N_59,In_1520,In_434);
or U60 (N_60,In_1134,In_51);
nand U61 (N_61,In_1843,In_1990);
nor U62 (N_62,In_99,In_522);
and U63 (N_63,In_877,In_919);
nand U64 (N_64,In_1916,In_659);
or U65 (N_65,In_504,In_1104);
and U66 (N_66,In_1492,In_170);
or U67 (N_67,In_1892,In_394);
nand U68 (N_68,In_1003,In_893);
xnor U69 (N_69,In_710,In_785);
or U70 (N_70,In_384,In_1842);
or U71 (N_71,In_856,In_285);
nand U72 (N_72,In_196,In_1352);
or U73 (N_73,In_1261,In_1638);
and U74 (N_74,In_970,In_93);
and U75 (N_75,In_1121,In_1670);
or U76 (N_76,In_800,In_1229);
xnor U77 (N_77,In_690,In_12);
and U78 (N_78,In_980,In_1972);
xnor U79 (N_79,In_24,In_1514);
and U80 (N_80,In_1795,In_389);
xnor U81 (N_81,In_1116,In_1436);
or U82 (N_82,In_1254,In_700);
nand U83 (N_83,In_1437,In_7);
nand U84 (N_84,In_120,In_626);
xor U85 (N_85,In_1541,In_1797);
xnor U86 (N_86,In_598,In_1624);
xor U87 (N_87,In_744,In_564);
nor U88 (N_88,In_1089,In_1167);
or U89 (N_89,In_766,In_798);
or U90 (N_90,In_294,In_1497);
nor U91 (N_91,In_1367,In_77);
nor U92 (N_92,In_675,In_1649);
and U93 (N_93,In_1694,In_410);
nand U94 (N_94,In_353,In_820);
nand U95 (N_95,In_533,In_968);
nor U96 (N_96,In_1151,In_923);
and U97 (N_97,In_1960,In_1345);
xor U98 (N_98,In_455,In_198);
and U99 (N_99,In_1391,In_1653);
and U100 (N_100,In_1082,In_489);
nand U101 (N_101,In_109,In_1641);
xnor U102 (N_102,In_1221,In_319);
or U103 (N_103,In_1635,In_730);
xnor U104 (N_104,In_1302,In_166);
and U105 (N_105,In_1161,In_366);
nor U106 (N_106,In_1525,In_1264);
nor U107 (N_107,In_1023,In_1461);
and U108 (N_108,In_1877,In_202);
xor U109 (N_109,In_1574,In_1714);
nor U110 (N_110,In_527,In_270);
or U111 (N_111,In_433,In_1890);
and U112 (N_112,In_1809,In_908);
nand U113 (N_113,In_1051,In_795);
or U114 (N_114,In_1681,In_760);
and U115 (N_115,In_1028,In_1561);
or U116 (N_116,In_1899,In_176);
and U117 (N_117,In_855,In_1773);
xor U118 (N_118,In_1096,In_9);
nor U119 (N_119,In_1118,In_344);
nor U120 (N_120,In_367,In_1612);
and U121 (N_121,In_1450,In_1249);
or U122 (N_122,In_804,In_45);
nand U123 (N_123,In_1476,In_1383);
nor U124 (N_124,In_1999,In_1713);
and U125 (N_125,In_1552,In_580);
and U126 (N_126,In_1283,In_991);
nor U127 (N_127,In_1236,In_1136);
xor U128 (N_128,In_1152,In_397);
or U129 (N_129,In_903,In_1691);
or U130 (N_130,In_587,In_697);
and U131 (N_131,In_551,In_76);
nor U132 (N_132,In_1884,In_897);
nand U133 (N_133,In_405,In_1591);
nor U134 (N_134,In_379,In_1353);
nor U135 (N_135,In_1812,In_509);
nor U136 (N_136,In_423,In_180);
xnor U137 (N_137,In_776,In_1252);
and U138 (N_138,In_1471,In_1961);
nor U139 (N_139,In_783,In_1906);
nand U140 (N_140,In_1386,In_722);
or U141 (N_141,In_484,In_1223);
xor U142 (N_142,In_496,In_918);
and U143 (N_143,In_688,In_439);
nand U144 (N_144,In_1431,In_289);
nor U145 (N_145,In_920,In_122);
or U146 (N_146,In_1138,In_1172);
and U147 (N_147,In_78,In_1241);
and U148 (N_148,In_1322,In_1778);
and U149 (N_149,In_57,In_470);
nand U150 (N_150,In_1922,In_1398);
xor U151 (N_151,In_138,In_542);
or U152 (N_152,In_1666,In_924);
nor U153 (N_153,In_696,In_1763);
or U154 (N_154,In_1711,In_1754);
nand U155 (N_155,In_1382,In_1366);
nand U156 (N_156,In_1558,In_773);
nand U157 (N_157,In_1122,In_1689);
and U158 (N_158,In_1072,In_812);
xnor U159 (N_159,In_1942,In_86);
nand U160 (N_160,In_83,In_177);
nand U161 (N_161,In_284,In_195);
and U162 (N_162,In_1732,In_1976);
and U163 (N_163,In_1129,In_1542);
or U164 (N_164,In_1365,In_664);
and U165 (N_165,In_333,In_1311);
and U166 (N_166,In_507,In_1397);
and U167 (N_167,In_913,In_1602);
and U168 (N_168,In_565,In_1086);
or U169 (N_169,In_233,In_1177);
nor U170 (N_170,In_1060,In_975);
and U171 (N_171,In_590,N_158);
nand U172 (N_172,In_318,In_1193);
xor U173 (N_173,In_1941,In_1688);
xor U174 (N_174,In_463,N_127);
nand U175 (N_175,In_1348,In_653);
and U176 (N_176,In_838,In_2);
nor U177 (N_177,In_1384,In_407);
nor U178 (N_178,In_21,In_1339);
or U179 (N_179,In_1936,In_577);
nor U180 (N_180,In_181,In_673);
nor U181 (N_181,In_1055,In_963);
xnor U182 (N_182,In_1253,N_61);
nand U183 (N_183,In_1769,In_998);
xnor U184 (N_184,In_375,In_1473);
xnor U185 (N_185,In_1278,In_1297);
or U186 (N_186,In_1043,In_497);
nand U187 (N_187,In_826,In_513);
xnor U188 (N_188,In_191,In_1149);
and U189 (N_189,N_96,In_135);
or U190 (N_190,In_1547,N_12);
nor U191 (N_191,In_1631,In_1826);
xnor U192 (N_192,In_1914,In_1176);
xor U193 (N_193,In_203,In_1881);
or U194 (N_194,In_52,In_1393);
nand U195 (N_195,In_1065,In_1833);
nand U196 (N_196,In_1701,In_452);
and U197 (N_197,In_1355,In_837);
or U198 (N_198,N_84,In_1731);
xor U199 (N_199,In_1108,In_1946);
xnor U200 (N_200,In_746,In_1952);
nand U201 (N_201,In_505,In_483);
or U202 (N_202,In_677,In_1284);
and U203 (N_203,In_737,In_831);
xor U204 (N_204,In_1604,In_1417);
xor U205 (N_205,In_1370,In_1927);
or U206 (N_206,In_1343,In_1664);
nand U207 (N_207,In_945,In_1672);
xnor U208 (N_208,In_1832,N_33);
and U209 (N_209,In_969,In_1066);
xor U210 (N_210,In_1968,In_235);
xor U211 (N_211,In_1636,In_1412);
nand U212 (N_212,In_1059,In_747);
nor U213 (N_213,In_1037,In_836);
nor U214 (N_214,In_1354,In_1537);
nor U215 (N_215,In_865,In_658);
nand U216 (N_216,In_1027,In_1105);
nor U217 (N_217,In_292,In_703);
nand U218 (N_218,In_538,In_806);
xnor U219 (N_219,In_633,In_1803);
nand U220 (N_220,N_23,In_1741);
nand U221 (N_221,In_101,N_11);
xnor U222 (N_222,N_95,In_486);
nor U223 (N_223,In_571,In_383);
or U224 (N_224,In_588,In_946);
nor U225 (N_225,In_1577,In_89);
nor U226 (N_226,In_479,In_840);
nand U227 (N_227,In_451,In_871);
and U228 (N_228,In_1539,In_751);
nand U229 (N_229,In_1827,In_1523);
nor U230 (N_230,In_857,In_667);
or U231 (N_231,N_76,In_1771);
nor U232 (N_232,In_293,In_1777);
xor U233 (N_233,In_589,In_761);
and U234 (N_234,In_1446,In_1310);
and U235 (N_235,N_141,In_686);
or U236 (N_236,In_448,In_1690);
xor U237 (N_237,In_584,N_4);
nand U238 (N_238,In_1620,In_715);
xor U239 (N_239,In_949,In_1106);
and U240 (N_240,In_1119,In_549);
nor U241 (N_241,In_1265,In_327);
nor U242 (N_242,In_989,In_905);
and U243 (N_243,In_1957,In_454);
nor U244 (N_244,N_135,In_1841);
nor U245 (N_245,In_38,In_115);
nand U246 (N_246,In_844,In_234);
nor U247 (N_247,In_1991,In_600);
nor U248 (N_248,In_627,In_17);
and U249 (N_249,In_1553,In_1719);
xor U250 (N_250,In_880,In_1042);
nor U251 (N_251,N_32,In_890);
xor U252 (N_252,In_1875,N_36);
nand U253 (N_253,N_13,In_1882);
nor U254 (N_254,In_1204,In_1988);
nor U255 (N_255,In_1317,In_1013);
nand U256 (N_256,In_1718,In_1704);
or U257 (N_257,N_137,In_834);
nor U258 (N_258,N_107,In_1901);
or U259 (N_259,N_153,In_1513);
or U260 (N_260,In_331,In_1734);
nand U261 (N_261,In_1462,In_1341);
nand U262 (N_262,In_16,In_681);
nand U263 (N_263,In_1715,In_94);
nand U264 (N_264,In_1818,In_780);
and U265 (N_265,In_79,In_252);
nand U266 (N_266,In_885,In_105);
and U267 (N_267,In_1846,In_1220);
and U268 (N_268,In_435,In_1894);
and U269 (N_269,In_324,In_541);
and U270 (N_270,In_1793,In_561);
nand U271 (N_271,In_92,In_743);
or U272 (N_272,In_466,N_34);
or U273 (N_273,In_1493,In_543);
xor U274 (N_274,In_733,In_1056);
xnor U275 (N_275,In_1000,In_1075);
and U276 (N_276,In_1614,In_15);
and U277 (N_277,In_552,In_1592);
or U278 (N_278,In_1259,In_498);
or U279 (N_279,In_1987,In_1433);
xnor U280 (N_280,In_1344,In_683);
nor U281 (N_281,In_1565,In_1325);
or U282 (N_282,N_25,In_340);
or U283 (N_283,In_53,In_412);
nand U284 (N_284,In_1909,In_174);
or U285 (N_285,In_1814,In_310);
nor U286 (N_286,In_637,N_131);
nor U287 (N_287,In_1137,In_22);
xnor U288 (N_288,In_240,In_1652);
and U289 (N_289,In_473,In_1184);
xor U290 (N_290,In_139,In_1218);
and U291 (N_291,In_1730,In_485);
nand U292 (N_292,In_583,In_1182);
and U293 (N_293,In_654,In_833);
xnor U294 (N_294,In_1373,In_558);
nand U295 (N_295,In_406,In_611);
xor U296 (N_296,In_1584,In_1187);
xor U297 (N_297,In_1939,In_1896);
xor U298 (N_298,In_227,In_1870);
xnor U299 (N_299,In_1237,In_1212);
nor U300 (N_300,In_1616,In_568);
xor U301 (N_301,N_48,In_644);
xor U302 (N_302,In_35,In_612);
or U303 (N_303,In_160,In_511);
and U304 (N_304,In_1443,In_1851);
and U305 (N_305,In_1989,In_71);
and U306 (N_306,In_212,In_1510);
xor U307 (N_307,In_54,In_1956);
and U308 (N_308,In_420,In_1717);
xor U309 (N_309,In_1621,In_432);
nor U310 (N_310,In_1396,In_41);
or U311 (N_311,In_188,In_1063);
nor U312 (N_312,In_326,In_1048);
nor U313 (N_313,In_1394,In_1665);
nor U314 (N_314,In_698,In_927);
xnor U315 (N_315,In_1727,In_272);
xnor U316 (N_316,N_105,In_1796);
and U317 (N_317,In_569,In_875);
or U318 (N_318,In_1675,In_1128);
or U319 (N_319,In_847,In_253);
nor U320 (N_320,In_1292,N_251);
nand U321 (N_321,N_0,In_1656);
nor U322 (N_322,In_621,N_63);
or U323 (N_323,In_1570,N_225);
or U324 (N_324,In_199,In_167);
and U325 (N_325,In_1905,In_217);
nor U326 (N_326,In_291,In_1811);
and U327 (N_327,In_154,In_849);
or U328 (N_328,In_721,In_332);
xor U329 (N_329,In_745,N_267);
and U330 (N_330,In_1248,N_192);
and U331 (N_331,In_186,In_870);
and U332 (N_332,In_887,In_1329);
xor U333 (N_333,N_151,In_308);
or U334 (N_334,In_1052,In_815);
nor U335 (N_335,In_720,N_204);
nand U336 (N_336,In_1937,In_1921);
xnor U337 (N_337,In_1678,In_1757);
or U338 (N_338,N_118,In_449);
or U339 (N_339,In_1180,In_1560);
xor U340 (N_340,N_145,In_829);
and U341 (N_341,In_1502,In_192);
or U342 (N_342,In_1556,In_299);
nand U343 (N_343,In_1073,In_793);
nor U344 (N_344,In_1406,N_38);
or U345 (N_345,N_53,In_594);
and U346 (N_346,N_302,In_1965);
and U347 (N_347,In_1005,N_314);
xnor U348 (N_348,In_1387,N_57);
nor U349 (N_349,In_471,In_628);
xor U350 (N_350,In_1423,In_649);
or U351 (N_351,In_1157,In_1874);
xnor U352 (N_352,In_387,In_750);
and U353 (N_353,In_100,N_17);
nor U354 (N_354,In_1611,In_1369);
nand U355 (N_355,In_953,In_1181);
xnor U356 (N_356,N_232,N_266);
or U357 (N_357,In_1444,In_430);
and U358 (N_358,In_368,In_1661);
and U359 (N_359,In_593,N_171);
or U360 (N_360,In_1974,N_257);
or U361 (N_361,In_245,In_1654);
nand U362 (N_362,In_1239,In_1872);
or U363 (N_363,In_605,In_1679);
or U364 (N_364,In_1538,In_1529);
nor U365 (N_365,In_977,In_1798);
nor U366 (N_366,In_1573,In_1848);
or U367 (N_367,In_1947,In_1500);
nand U368 (N_368,In_528,In_1575);
and U369 (N_369,In_307,In_1153);
and U370 (N_370,In_55,N_189);
xor U371 (N_371,In_1954,In_1183);
xor U372 (N_372,In_1943,In_853);
and U373 (N_373,In_98,In_1865);
or U374 (N_374,In_1629,In_1676);
nor U375 (N_375,In_1256,In_692);
nand U376 (N_376,In_492,In_1021);
xnor U377 (N_377,In_1687,In_821);
nand U378 (N_378,N_161,In_599);
nor U379 (N_379,In_1897,N_75);
nor U380 (N_380,In_1390,In_396);
nor U381 (N_381,In_614,In_1931);
and U382 (N_382,In_390,In_685);
nor U383 (N_383,In_91,In_1505);
or U384 (N_384,In_823,In_1985);
and U385 (N_385,In_481,In_846);
nand U386 (N_386,N_262,In_493);
nor U387 (N_387,N_176,In_345);
nand U388 (N_388,In_889,In_805);
and U389 (N_389,In_157,N_9);
nor U390 (N_390,In_1871,N_183);
xor U391 (N_391,In_1162,In_250);
nand U392 (N_392,In_881,In_1996);
or U393 (N_393,N_27,In_1634);
or U394 (N_394,In_445,In_322);
nand U395 (N_395,In_786,In_380);
nand U396 (N_396,In_1306,In_125);
nand U397 (N_397,In_851,N_213);
and U398 (N_398,In_1904,In_1448);
xnor U399 (N_399,N_264,N_284);
xnor U400 (N_400,In_1247,In_1113);
nand U401 (N_401,In_297,In_629);
or U402 (N_402,In_1053,In_211);
xnor U403 (N_403,In_475,N_205);
and U404 (N_404,N_224,In_1145);
nor U405 (N_405,In_687,In_1545);
or U406 (N_406,In_1001,In_638);
or U407 (N_407,In_777,In_0);
or U408 (N_408,In_1411,In_1222);
and U409 (N_409,N_50,N_293);
nor U410 (N_410,In_1766,In_1095);
nor U411 (N_411,In_1720,N_256);
nand U412 (N_412,In_431,In_1879);
xor U413 (N_413,In_461,N_211);
and U414 (N_414,In_1615,In_650);
xnor U415 (N_415,In_1950,N_190);
xor U416 (N_416,In_1637,In_1737);
nand U417 (N_417,N_258,In_361);
xnor U418 (N_418,In_518,In_69);
or U419 (N_419,N_274,In_1663);
and U420 (N_420,In_480,In_632);
or U421 (N_421,In_925,In_1456);
xor U422 (N_422,In_693,In_1765);
nand U423 (N_423,In_935,In_392);
nor U424 (N_424,In_864,N_111);
and U425 (N_425,In_1126,In_1405);
xnor U426 (N_426,In_1932,In_194);
xor U427 (N_427,In_708,In_1824);
or U428 (N_428,N_203,In_1728);
or U429 (N_429,In_1958,In_618);
or U430 (N_430,N_228,In_520);
and U431 (N_431,In_1421,In_794);
nand U432 (N_432,In_811,N_282);
and U433 (N_433,In_269,In_136);
or U434 (N_434,In_950,In_1282);
and U435 (N_435,N_310,In_1244);
or U436 (N_436,In_258,In_75);
or U437 (N_437,N_248,In_1756);
xor U438 (N_438,In_1170,In_539);
xor U439 (N_439,In_1944,In_1736);
and U440 (N_440,In_352,In_1069);
nor U441 (N_441,In_399,In_1300);
and U442 (N_442,In_364,In_1019);
nand U443 (N_443,In_1609,In_1058);
nor U444 (N_444,N_167,N_212);
and U445 (N_445,In_182,In_1619);
xor U446 (N_446,In_1074,In_1362);
xor U447 (N_447,In_348,In_1740);
xor U448 (N_448,In_641,N_92);
xnor U449 (N_449,In_516,In_1594);
or U450 (N_450,In_1238,N_303);
and U451 (N_451,In_848,In_1357);
xor U452 (N_452,In_1430,In_763);
or U453 (N_453,In_462,In_278);
or U454 (N_454,In_1071,In_774);
and U455 (N_455,In_358,In_1685);
and U456 (N_456,In_1830,In_1330);
or U457 (N_457,In_133,In_1198);
or U458 (N_458,In_961,In_158);
nor U459 (N_459,In_97,In_1439);
nor U460 (N_460,In_309,In_678);
nor U461 (N_461,N_116,In_70);
nand U462 (N_462,In_1760,In_1503);
or U463 (N_463,In_296,In_427);
or U464 (N_464,In_315,In_741);
nand U465 (N_465,In_952,In_13);
nor U466 (N_466,In_1288,In_1318);
nor U467 (N_467,In_1210,N_41);
xnor U468 (N_468,In_1478,In_1512);
nor U469 (N_469,In_797,In_1572);
and U470 (N_470,In_1536,In_323);
and U471 (N_471,In_689,In_1643);
or U472 (N_472,In_828,In_738);
xnor U473 (N_473,N_271,In_1992);
nand U474 (N_474,In_1331,In_1016);
xnor U475 (N_475,In_305,N_234);
xnor U476 (N_476,In_1840,In_1915);
nor U477 (N_477,In_172,N_163);
nand U478 (N_478,In_824,In_1605);
nand U479 (N_479,In_537,N_114);
xor U480 (N_480,In_261,In_1401);
and U481 (N_481,In_117,In_1191);
nor U482 (N_482,N_320,In_534);
and U483 (N_483,N_368,In_388);
nand U484 (N_484,In_408,N_438);
or U485 (N_485,In_1091,In_317);
or U486 (N_486,In_657,In_209);
xnor U487 (N_487,In_1721,N_97);
xor U488 (N_488,N_410,In_957);
xor U489 (N_489,In_242,In_251);
xnor U490 (N_490,In_1981,N_24);
nand U491 (N_491,In_58,N_462);
nand U492 (N_492,N_359,In_546);
nand U493 (N_493,In_557,N_477);
nand U494 (N_494,In_1133,In_1208);
or U495 (N_495,N_338,N_62);
nand U496 (N_496,In_1750,In_506);
nand U497 (N_497,In_1789,In_1213);
nor U498 (N_498,In_339,In_1227);
xor U499 (N_499,In_349,In_842);
xor U500 (N_500,In_525,N_450);
or U501 (N_501,N_235,N_309);
nand U502 (N_502,In_576,N_129);
and U503 (N_503,In_1869,In_1039);
nor U504 (N_504,In_1289,In_694);
xnor U505 (N_505,In_1579,In_1655);
nand U506 (N_506,In_1438,In_1868);
and U507 (N_507,In_1806,N_2);
xnor U508 (N_508,In_378,In_1938);
xor U509 (N_509,In_146,In_1810);
nor U510 (N_510,In_799,N_89);
nand U511 (N_511,In_30,In_1372);
and U512 (N_512,In_403,In_521);
nor U513 (N_513,N_83,In_1844);
or U514 (N_514,In_1408,In_1078);
xor U515 (N_515,In_559,In_1114);
or U516 (N_516,N_290,In_1695);
nor U517 (N_517,In_1995,N_125);
and U518 (N_518,In_1242,In_642);
nor U519 (N_519,N_369,In_802);
xnor U520 (N_520,In_10,In_458);
and U521 (N_521,In_303,N_191);
and U522 (N_522,In_27,In_1034);
nor U523 (N_523,In_1794,N_130);
or U524 (N_524,In_1379,In_1268);
nand U525 (N_525,In_1522,In_1361);
and U526 (N_526,In_1432,In_1628);
nand U527 (N_527,In_33,In_947);
nor U528 (N_528,In_1142,In_1115);
xor U529 (N_529,In_347,In_1823);
or U530 (N_530,In_996,In_1920);
nor U531 (N_531,N_221,In_183);
xnor U532 (N_532,In_586,In_1969);
and U533 (N_533,In_1451,In_956);
and U534 (N_534,In_112,In_59);
nor U535 (N_535,In_544,In_869);
nor U536 (N_536,In_1800,In_1693);
and U537 (N_537,In_610,N_383);
xor U538 (N_538,In_1758,In_922);
nand U539 (N_539,In_1385,In_1626);
nand U540 (N_540,In_271,In_1404);
or U541 (N_541,In_1983,In_732);
or U542 (N_542,In_550,In_554);
or U543 (N_543,In_416,N_401);
and U544 (N_544,In_1279,N_345);
or U545 (N_545,In_453,In_902);
or U546 (N_546,N_449,N_119);
and U547 (N_547,In_400,In_789);
or U548 (N_548,N_73,In_960);
or U549 (N_549,N_458,In_357);
nor U550 (N_550,In_1186,In_300);
nand U551 (N_551,In_1440,N_260);
or U552 (N_552,In_1257,N_79);
nand U553 (N_553,In_959,In_862);
and U554 (N_554,In_1535,In_1099);
and U555 (N_555,In_1784,N_21);
and U556 (N_556,In_85,In_441);
nand U557 (N_557,In_225,In_450);
or U558 (N_558,N_297,In_356);
xor U559 (N_559,In_1967,In_531);
and U560 (N_560,N_467,In_563);
nand U561 (N_561,In_1164,In_1792);
and U562 (N_562,In_1776,In_1650);
nor U563 (N_563,N_132,In_801);
xor U564 (N_564,N_279,In_1903);
xnor U565 (N_565,In_1017,In_343);
or U566 (N_566,N_328,In_1441);
and U567 (N_567,In_1576,In_939);
and U568 (N_568,In_273,N_268);
and U569 (N_569,N_373,In_1601);
or U570 (N_570,In_636,In_1524);
xor U571 (N_571,In_899,In_1231);
or U572 (N_572,In_338,In_1603);
and U573 (N_573,In_1360,In_1966);
xor U574 (N_574,In_861,In_175);
nor U575 (N_575,In_34,N_98);
nor U576 (N_576,In_742,N_378);
nand U577 (N_577,In_20,In_1010);
nor U578 (N_578,N_300,In_915);
or U579 (N_579,In_1569,In_287);
xor U580 (N_580,In_860,N_87);
nor U581 (N_581,In_1554,In_1209);
or U582 (N_582,In_169,In_656);
and U583 (N_583,N_22,In_1340);
xor U584 (N_584,In_503,In_911);
and U585 (N_585,In_1640,N_387);
or U586 (N_586,N_15,In_1080);
or U587 (N_587,In_1266,In_1024);
nor U588 (N_588,In_1913,N_296);
and U589 (N_589,In_415,N_331);
and U590 (N_590,In_137,N_403);
and U591 (N_591,In_1599,In_8);
or U592 (N_592,In_1808,In_867);
nand U593 (N_593,N_289,In_1817);
nor U594 (N_594,N_216,In_419);
nand U595 (N_595,In_1980,In_1738);
or U596 (N_596,N_377,In_369);
nor U597 (N_597,N_7,N_18);
and U598 (N_598,In_1551,N_444);
nor U599 (N_599,In_1004,N_6);
nor U600 (N_600,In_1315,In_1998);
xnor U601 (N_601,In_943,In_37);
nand U602 (N_602,In_200,In_36);
or U603 (N_603,In_547,In_1562);
nand U604 (N_604,In_46,In_131);
nand U605 (N_605,N_391,In_1898);
xnor U606 (N_606,In_1356,N_287);
and U607 (N_607,In_671,In_421);
nor U608 (N_608,In_938,In_825);
or U609 (N_609,In_1363,N_194);
or U610 (N_610,In_1725,In_1131);
nor U611 (N_611,N_374,N_174);
nand U612 (N_612,In_515,In_1853);
or U613 (N_613,In_365,In_204);
and U614 (N_614,In_280,N_121);
nor U615 (N_615,In_1467,In_1907);
nor U616 (N_616,In_1984,In_680);
nand U617 (N_617,In_640,In_311);
or U618 (N_618,N_440,In_1657);
nor U619 (N_619,In_26,In_124);
and U620 (N_620,In_1767,In_153);
nand U621 (N_621,In_1332,In_414);
xnor U622 (N_622,In_426,In_972);
nand U623 (N_623,In_1413,In_354);
or U624 (N_624,N_336,N_366);
or U625 (N_625,N_101,In_467);
nand U626 (N_626,In_246,N_360);
or U627 (N_627,N_350,In_1735);
nor U628 (N_628,In_1169,In_948);
or U629 (N_629,N_406,In_602);
or U630 (N_630,In_1759,N_179);
nand U631 (N_631,In_1324,In_1158);
or U632 (N_632,In_106,N_173);
nor U633 (N_633,In_84,In_1595);
xnor U634 (N_634,In_1895,In_476);
nor U635 (N_635,In_1276,In_1111);
nand U636 (N_636,In_1951,In_438);
and U637 (N_637,In_1683,In_429);
nand U638 (N_638,N_445,In_306);
nor U639 (N_639,In_762,In_1886);
and U640 (N_640,In_1081,In_113);
or U641 (N_641,In_1726,In_1224);
nor U642 (N_642,In_1930,N_496);
nand U643 (N_643,N_56,In_208);
xnor U644 (N_644,In_1140,N_522);
xnor U645 (N_645,In_376,In_87);
nor U646 (N_646,N_10,In_1240);
or U647 (N_647,In_68,N_115);
xnor U648 (N_648,N_292,N_277);
or U649 (N_649,N_143,In_1540);
and U650 (N_650,N_609,In_128);
nor U651 (N_651,In_1703,In_1761);
nor U652 (N_652,N_611,N_100);
nor U653 (N_653,In_896,In_401);
or U654 (N_654,In_1531,In_1087);
xnor U655 (N_655,N_589,N_498);
and U656 (N_656,N_459,In_907);
nand U657 (N_657,In_647,In_1346);
xnor U658 (N_658,In_1854,In_814);
or U659 (N_659,In_1802,In_1488);
nand U660 (N_660,In_1770,In_1350);
or U661 (N_661,In_1608,In_74);
and U662 (N_662,In_1790,In_1532);
nor U663 (N_663,In_1219,In_1516);
or U664 (N_664,N_424,N_329);
xor U665 (N_665,In_1094,In_80);
xnor U666 (N_666,N_446,In_1216);
and U667 (N_667,In_474,N_586);
nor U668 (N_668,N_353,In_1729);
or U669 (N_669,In_65,In_1303);
nand U670 (N_670,N_480,N_570);
or U671 (N_671,N_283,In_32);
or U672 (N_672,In_1020,In_346);
or U673 (N_673,N_263,In_1660);
nand U674 (N_674,In_645,In_1747);
nand U675 (N_675,In_1739,N_604);
or U676 (N_676,N_217,N_616);
and U677 (N_677,In_148,N_415);
or U678 (N_678,N_605,N_428);
nor U679 (N_679,In_1470,In_661);
nor U680 (N_680,In_1155,In_108);
nor U681 (N_681,N_506,In_104);
xnor U682 (N_682,In_809,In_1975);
and U683 (N_683,In_1215,N_321);
xor U684 (N_684,N_51,In_145);
nor U685 (N_685,N_470,N_516);
nand U686 (N_686,N_270,In_1389);
xor U687 (N_687,In_622,In_724);
xnor U688 (N_688,In_1494,In_42);
nor U689 (N_689,In_1856,N_394);
and U690 (N_690,In_428,In_1112);
or U691 (N_691,In_440,In_937);
and U692 (N_692,In_1045,In_676);
xnor U693 (N_693,N_479,N_575);
nand U694 (N_694,N_304,N_307);
nor U695 (N_695,In_1548,N_491);
and U696 (N_696,In_819,In_134);
nand U697 (N_697,In_249,In_548);
or U698 (N_698,In_402,N_222);
nand U699 (N_699,N_511,In_223);
and U700 (N_700,N_247,In_1933);
xnor U701 (N_701,N_156,N_399);
nand U702 (N_702,N_45,In_702);
or U703 (N_703,In_1376,In_491);
and U704 (N_704,N_39,In_152);
nor U705 (N_705,In_994,N_411);
and U706 (N_706,In_1293,In_1934);
xnor U707 (N_707,N_324,N_568);
xnor U708 (N_708,In_1359,In_276);
or U709 (N_709,In_1410,N_578);
xnor U710 (N_710,N_31,In_731);
xnor U711 (N_711,N_405,In_1527);
nor U712 (N_712,N_562,In_845);
nor U713 (N_713,In_572,In_1477);
nand U714 (N_714,In_1092,In_1375);
xor U715 (N_715,In_718,N_313);
or U716 (N_716,In_609,N_237);
or U717 (N_717,In_895,In_1409);
nor U718 (N_718,In_1722,N_486);
or U719 (N_719,N_457,In_350);
xor U720 (N_720,In_1630,N_124);
and U721 (N_721,In_1588,In_1335);
nor U722 (N_722,N_574,In_1173);
or U723 (N_723,N_177,N_613);
xnor U724 (N_724,In_1692,In_1197);
xnor U725 (N_725,In_684,In_312);
nor U726 (N_726,In_524,In_238);
xnor U727 (N_727,In_132,In_764);
xnor U728 (N_728,In_1466,N_133);
nor U729 (N_729,N_59,N_291);
xnor U730 (N_730,N_612,N_197);
xnor U731 (N_731,In_987,In_360);
nand U732 (N_732,In_1007,In_95);
or U733 (N_733,In_1334,N_342);
nor U734 (N_734,In_1490,N_514);
nor U735 (N_735,In_695,In_29);
and U736 (N_736,In_1495,In_1600);
xnor U737 (N_737,N_358,N_219);
nand U738 (N_738,In_1949,In_1098);
xor U739 (N_739,N_255,N_599);
or U740 (N_740,In_502,N_372);
xnor U741 (N_741,N_561,In_1491);
nor U742 (N_742,In_635,In_1751);
or U743 (N_743,In_48,In_1319);
nor U744 (N_744,N_242,In_1243);
and U745 (N_745,In_1154,N_594);
and U746 (N_746,In_1696,In_140);
nand U747 (N_747,In_281,In_1233);
or U748 (N_748,In_1280,In_232);
nor U749 (N_749,In_1813,N_233);
nand U750 (N_750,N_241,In_879);
nand U751 (N_751,In_1633,In_1508);
xnor U752 (N_752,In_1018,In_1659);
and U753 (N_753,In_1123,In_1507);
nand U754 (N_754,In_90,N_476);
nor U755 (N_755,N_117,N_37);
or U756 (N_756,In_382,In_321);
nor U757 (N_757,N_103,In_61);
and U758 (N_758,N_597,In_983);
and U759 (N_759,N_364,N_223);
xor U760 (N_760,In_316,In_119);
nor U761 (N_761,In_1911,In_1642);
or U762 (N_762,In_941,In_719);
nand U763 (N_763,N_558,N_272);
or U764 (N_764,N_207,In_67);
nor U765 (N_765,In_1891,In_1141);
nand U766 (N_766,In_1710,In_526);
or U767 (N_767,In_73,In_1578);
or U768 (N_768,In_1860,In_1501);
or U769 (N_769,In_218,N_351);
nor U770 (N_770,In_759,N_499);
xor U771 (N_771,In_974,N_346);
and U772 (N_772,N_508,N_261);
nor U773 (N_773,N_226,In_359);
nor U774 (N_774,In_1465,In_1787);
or U775 (N_775,N_639,In_951);
xnor U776 (N_776,In_1838,In_1305);
nand U777 (N_777,In_1863,In_606);
xor U778 (N_778,In_1320,In_1563);
nand U779 (N_779,In_1684,N_567);
xnor U780 (N_780,N_531,In_1295);
or U781 (N_781,N_465,N_231);
nand U782 (N_782,In_778,In_1880);
and U783 (N_783,N_482,In_1940);
xor U784 (N_784,N_99,In_472);
nand U785 (N_785,In_1165,In_337);
nand U786 (N_786,In_1607,In_237);
and U787 (N_787,In_43,In_1864);
and U788 (N_788,In_1668,In_872);
xnor U789 (N_789,In_31,In_1698);
nand U790 (N_790,In_1900,N_572);
and U791 (N_791,In_1712,In_1674);
and U792 (N_792,In_1371,In_40);
or U793 (N_793,N_635,N_240);
or U794 (N_794,In_442,N_162);
or U795 (N_795,N_543,In_1646);
nand U796 (N_796,In_82,In_224);
nor U797 (N_797,In_341,N_182);
nor U798 (N_798,N_454,N_427);
xor U799 (N_799,N_434,N_281);
or U800 (N_800,N_52,In_1449);
or U801 (N_801,In_418,In_1296);
xor U802 (N_802,N_566,In_1566);
and U803 (N_803,N_761,In_765);
xnor U804 (N_804,In_1716,In_1742);
or U805 (N_805,In_1147,N_8);
or U806 (N_806,In_1474,In_810);
nand U807 (N_807,N_538,N_325);
nor U808 (N_808,In_1203,In_1807);
xor U809 (N_809,N_710,In_863);
and U810 (N_810,In_1030,In_1006);
or U811 (N_811,N_333,In_1801);
or U812 (N_812,In_1707,In_682);
and U813 (N_813,N_745,In_523);
nor U814 (N_814,In_156,In_1733);
xnor U815 (N_815,N_593,N_706);
or U816 (N_816,In_1945,N_573);
nand U817 (N_817,In_1143,N_585);
and U818 (N_818,In_729,In_1057);
xnor U819 (N_819,In_336,N_308);
nand U820 (N_820,In_1651,In_1230);
or U821 (N_821,In_1400,In_1709);
and U822 (N_822,N_20,N_627);
and U823 (N_823,N_759,In_892);
nand U824 (N_824,In_1953,N_793);
and U825 (N_825,In_1580,N_670);
nor U826 (N_826,In_1973,In_63);
xor U827 (N_827,In_1418,In_1487);
nand U828 (N_828,N_713,In_1658);
nor U829 (N_829,In_1861,In_298);
and U830 (N_830,In_130,In_884);
or U831 (N_831,N_532,In_772);
xnor U832 (N_832,In_1174,In_1135);
nand U833 (N_833,In_1032,N_72);
xnor U834 (N_834,N_708,N_741);
nor U835 (N_835,N_199,N_348);
nand U836 (N_836,N_412,N_697);
xor U837 (N_837,N_792,In_28);
nor U838 (N_838,In_965,N_649);
or U839 (N_839,N_400,In_758);
or U840 (N_840,N_452,N_344);
nor U841 (N_841,N_484,In_1571);
nor U842 (N_842,N_28,N_764);
nand U843 (N_843,In_179,N_341);
nor U844 (N_844,In_1272,N_494);
xnor U845 (N_845,N_109,In_1847);
nor U846 (N_846,In_459,In_822);
or U847 (N_847,In_1468,In_111);
nand U848 (N_848,In_1482,N_664);
and U849 (N_849,In_1917,In_1918);
xnor U850 (N_850,N_563,N_738);
nand U851 (N_851,N_230,In_1309);
nor U852 (N_852,In_263,In_1831);
or U853 (N_853,In_1815,N_487);
and U854 (N_854,N_58,In_984);
or U855 (N_855,In_736,In_816);
nand U856 (N_856,N_789,In_1912);
nor U857 (N_857,In_1351,In_1764);
nor U858 (N_858,In_256,N_610);
xnor U859 (N_859,N_390,N_652);
nor U860 (N_860,In_582,In_162);
xor U861 (N_861,N_417,N_744);
xor U862 (N_862,In_646,N_726);
xnor U863 (N_863,In_372,In_1997);
nor U864 (N_864,N_743,N_544);
xnor U865 (N_865,In_4,In_934);
nor U866 (N_866,In_1434,In_1403);
and U867 (N_867,In_1110,N_278);
nand U868 (N_868,In_999,N_413);
xnor U869 (N_869,N_16,N_674);
nor U870 (N_870,In_1299,In_1277);
nor U871 (N_871,In_254,N_535);
nor U872 (N_872,N_724,N_259);
xor U873 (N_873,N_667,In_782);
xnor U874 (N_874,In_510,N_769);
nor U875 (N_875,In_769,In_1050);
and U876 (N_876,In_1928,In_1910);
and U877 (N_877,N_335,In_717);
nand U878 (N_878,In_1550,In_81);
or U879 (N_879,In_1582,In_283);
nor U880 (N_880,In_1677,In_1959);
nand U881 (N_881,In_1090,N_196);
nor U882 (N_882,N_437,In_1100);
or U883 (N_883,N_632,N_316);
xor U884 (N_884,In_1312,In_1217);
nor U885 (N_885,N_776,In_1103);
or U886 (N_886,N_763,N_500);
nand U887 (N_887,N_633,In_295);
nor U888 (N_888,In_1316,N_766);
and U889 (N_889,N_598,In_159);
or U890 (N_890,N_206,In_932);
or U891 (N_891,N_799,In_1067);
xnor U892 (N_892,N_775,In_1786);
xor U893 (N_893,In_1205,N_638);
nand U894 (N_894,N_729,In_330);
nor U895 (N_895,In_916,N_541);
xor U896 (N_896,N_788,In_1194);
nor U897 (N_897,N_576,In_1779);
xnor U898 (N_898,N_489,In_1304);
nor U899 (N_899,N_402,In_1225);
nand U900 (N_900,In_60,In_660);
and U901 (N_901,N_779,N_557);
and U902 (N_902,In_1260,In_617);
xnor U903 (N_903,N_363,In_1862);
xor U904 (N_904,N_507,In_370);
nand U905 (N_905,In_1012,In_1889);
nand U906 (N_906,In_1392,In_1544);
and U907 (N_907,N_634,N_306);
nor U908 (N_908,N_407,N_110);
and U909 (N_909,In_944,In_488);
nand U910 (N_910,N_154,N_43);
and U911 (N_911,N_108,N_551);
or U912 (N_912,N_679,N_720);
nor U913 (N_913,In_1517,In_1185);
and U914 (N_914,In_279,N_601);
xor U915 (N_915,N_185,N_317);
or U916 (N_916,In_1327,In_495);
nor U917 (N_917,In_1825,In_147);
xor U918 (N_918,N_501,In_669);
nand U919 (N_919,N_187,N_517);
or U920 (N_920,In_536,N_644);
xnor U921 (N_921,In_1235,In_1189);
and U922 (N_922,In_149,N_448);
nor U923 (N_923,In_592,N_134);
xnor U924 (N_924,In_978,In_1107);
and U925 (N_925,In_118,N_425);
xnor U926 (N_926,In_301,N_787);
nand U927 (N_927,In_1533,N_748);
and U928 (N_928,N_85,In_791);
nand U929 (N_929,In_1125,N_523);
and U930 (N_930,N_188,In_121);
xnor U931 (N_931,In_906,In_142);
xor U932 (N_932,In_444,N_530);
nand U933 (N_933,In_501,N_343);
nor U934 (N_934,N_687,In_672);
nor U935 (N_935,N_695,In_854);
and U936 (N_936,In_1994,In_1294);
and U937 (N_937,In_44,In_265);
and U938 (N_938,In_1908,N_160);
nor U939 (N_939,N_128,N_614);
and U940 (N_940,N_379,In_241);
and U941 (N_941,N_54,In_215);
nand U942 (N_942,N_752,N_701);
or U943 (N_943,In_1835,In_630);
or U944 (N_944,N_723,In_1378);
nor U945 (N_945,In_193,N_643);
and U946 (N_946,N_136,N_104);
and U947 (N_947,N_640,N_629);
nand U948 (N_948,N_165,In_674);
nand U949 (N_949,In_986,N_3);
and U950 (N_950,N_209,In_286);
nand U951 (N_951,N_149,N_584);
xnor U952 (N_952,N_354,In_190);
nand U953 (N_953,N_636,In_1374);
and U954 (N_954,In_1852,N_1);
and U955 (N_955,In_1593,In_62);
nand U956 (N_956,N_388,N_138);
or U957 (N_957,In_1705,N_442);
xor U958 (N_958,N_698,N_739);
xnor U959 (N_959,N_751,In_1772);
nand U960 (N_960,In_1314,N_675);
xor U961 (N_961,N_275,N_529);
nand U962 (N_962,N_880,In_1047);
or U963 (N_963,N_848,In_1267);
xor U964 (N_964,In_992,N_460);
and U965 (N_965,N_483,In_841);
nor U966 (N_966,In_229,N_772);
nand U967 (N_967,In_1680,N_229);
xor U968 (N_968,N_478,N_386);
xnor U969 (N_969,In_878,N_542);
xor U970 (N_970,In_116,N_921);
xnor U971 (N_971,In_573,In_748);
xor U972 (N_972,In_665,N_862);
nand U973 (N_973,In_711,N_932);
nand U974 (N_974,N_942,N_653);
nand U975 (N_975,N_365,In_11);
nor U976 (N_976,In_1130,N_953);
nand U977 (N_977,In_1479,In_1402);
nor U978 (N_978,In_756,N_665);
xor U979 (N_979,In_1061,N_829);
or U980 (N_980,N_615,In_257);
nand U981 (N_981,In_1481,In_771);
and U982 (N_982,In_740,N_835);
xnor U983 (N_983,In_1040,In_1083);
nor U984 (N_984,N_80,In_770);
or U985 (N_985,In_275,In_436);
or U986 (N_986,In_1752,In_1424);
nor U987 (N_987,In_1469,N_721);
xor U988 (N_988,In_411,In_1755);
nor U989 (N_989,N_463,N_590);
and U990 (N_990,In_6,In_494);
nor U991 (N_991,N_493,N_944);
or U992 (N_992,In_601,N_822);
or U993 (N_993,In_1515,N_931);
and U994 (N_994,N_436,In_259);
xnor U995 (N_995,In_1543,N_423);
xnor U996 (N_996,In_859,N_870);
nand U997 (N_997,N_801,N_503);
and U998 (N_998,N_936,N_901);
or U999 (N_999,In_1459,In_216);
and U1000 (N_1000,N_14,In_1035);
xor U1001 (N_1001,N_181,N_803);
nand U1002 (N_1002,N_794,In_1887);
and U1003 (N_1003,N_361,N_510);
xnor U1004 (N_1004,In_1036,N_347);
and U1005 (N_1005,N_550,N_672);
nand U1006 (N_1006,In_817,N_250);
and U1007 (N_1007,In_1109,N_805);
and U1008 (N_1008,N_758,N_774);
xor U1009 (N_1009,N_844,In_1673);
nand U1010 (N_1010,N_628,N_252);
and U1011 (N_1011,N_81,In_490);
xor U1012 (N_1012,N_461,In_830);
and U1013 (N_1013,In_1380,N_797);
nor U1014 (N_1014,In_712,N_655);
or U1015 (N_1015,In_704,N_126);
xnor U1016 (N_1016,N_265,N_700);
nand U1017 (N_1017,N_750,In_72);
nand U1018 (N_1018,In_425,N_330);
xnor U1019 (N_1019,N_814,N_874);
and U1020 (N_1020,In_1555,In_818);
nor U1021 (N_1021,N_184,In_1749);
nor U1022 (N_1022,N_868,In_50);
xor U1023 (N_1023,In_173,N_474);
nor U1024 (N_1024,In_578,In_535);
or U1025 (N_1025,N_294,In_447);
nand U1026 (N_1026,N_624,N_148);
xor U1027 (N_1027,N_236,In_381);
or U1028 (N_1028,In_1804,In_662);
nor U1029 (N_1029,N_783,In_1743);
and U1030 (N_1030,In_942,N_846);
and U1031 (N_1031,In_1377,N_946);
xnor U1032 (N_1032,In_1883,N_908);
nand U1033 (N_1033,In_1463,In_1708);
or U1034 (N_1034,N_273,N_332);
xor U1035 (N_1035,N_569,In_1336);
or U1036 (N_1036,N_899,N_747);
xor U1037 (N_1037,N_714,In_1144);
xnor U1038 (N_1038,In_1195,In_832);
nor U1039 (N_1039,In_96,In_1407);
or U1040 (N_1040,N_582,In_1178);
and U1041 (N_1041,In_1026,In_1590);
and U1042 (N_1042,N_898,N_902);
or U1043 (N_1043,N_220,N_276);
nand U1044 (N_1044,In_189,N_548);
nand U1045 (N_1045,In_624,N_785);
xnor U1046 (N_1046,In_468,N_488);
nor U1047 (N_1047,N_676,N_917);
nand U1048 (N_1048,N_715,In_512);
nand U1049 (N_1049,In_808,N_923);
or U1050 (N_1050,In_220,In_604);
nor U1051 (N_1051,N_429,In_1484);
xnor U1052 (N_1052,N_102,N_186);
nor U1053 (N_1053,N_784,In_409);
xor U1054 (N_1054,N_883,N_736);
nor U1055 (N_1055,In_1291,In_1671);
nand U1056 (N_1056,In_1273,In_1475);
and U1057 (N_1057,N_879,N_866);
nand U1058 (N_1058,In_603,In_1748);
xor U1059 (N_1059,In_277,N_208);
nor U1060 (N_1060,In_313,N_957);
nor U1061 (N_1061,N_680,In_651);
and U1062 (N_1062,In_66,N_757);
nor U1063 (N_1063,In_1419,N_646);
nand U1064 (N_1064,In_187,N_847);
nor U1065 (N_1065,In_579,In_1489);
nand U1066 (N_1066,In_1885,N_897);
nand U1067 (N_1067,N_941,N_88);
and U1068 (N_1068,N_737,N_725);
nand U1069 (N_1069,In_1062,N_245);
xnor U1070 (N_1070,N_370,N_389);
or U1071 (N_1071,N_888,N_854);
xor U1072 (N_1072,In_596,In_500);
xnor U1073 (N_1073,N_311,In_981);
nand U1074 (N_1074,In_1850,N_727);
nor U1075 (N_1075,N_711,In_1226);
or U1076 (N_1076,In_723,N_735);
nor U1077 (N_1077,N_765,In_709);
nor U1078 (N_1078,In_668,In_1639);
nor U1079 (N_1079,N_684,In_236);
xnor U1080 (N_1080,N_238,N_855);
nand U1081 (N_1081,In_1648,N_592);
nand U1082 (N_1082,N_831,In_530);
or U1083 (N_1083,N_853,N_762);
nand U1084 (N_1084,In_1427,N_950);
nor U1085 (N_1085,N_707,N_352);
nor U1086 (N_1086,N_907,N_69);
nand U1087 (N_1087,N_334,In_567);
nor U1088 (N_1088,In_1559,N_754);
nand U1089 (N_1089,N_397,N_820);
and U1090 (N_1090,N_671,In_1557);
and U1091 (N_1091,N_617,N_945);
or U1092 (N_1092,In_555,N_159);
or U1093 (N_1093,In_873,N_367);
xor U1094 (N_1094,In_1702,N_786);
and U1095 (N_1095,N_398,N_288);
and U1096 (N_1096,In_1858,In_701);
xor U1097 (N_1097,N_914,N_693);
or U1098 (N_1098,N_804,In_843);
and U1099 (N_1099,N_851,N_660);
and U1100 (N_1100,In_954,N_692);
xnor U1101 (N_1101,N_852,N_580);
or U1102 (N_1102,N_419,In_1416);
or U1103 (N_1103,N_889,In_1049);
and U1104 (N_1104,In_691,In_1700);
nand U1105 (N_1105,In_1923,In_1828);
and U1106 (N_1106,In_1285,N_928);
and U1107 (N_1107,In_178,In_936);
nor U1108 (N_1108,N_473,In_752);
nand U1109 (N_1109,N_553,N_526);
nor U1110 (N_1110,N_677,N_893);
and U1111 (N_1111,In_566,N_689);
xnor U1112 (N_1112,In_1697,N_170);
or U1113 (N_1113,In_835,In_1935);
nand U1114 (N_1114,In_1422,N_832);
and U1115 (N_1115,N_305,N_869);
nand U1116 (N_1116,N_834,N_524);
xnor U1117 (N_1117,In_574,In_900);
and U1118 (N_1118,In_639,N_951);
and U1119 (N_1119,N_139,In_931);
nor U1120 (N_1120,N_685,N_495);
xnor U1121 (N_1121,N_155,N_591);
nand U1122 (N_1122,N_481,N_767);
and U1123 (N_1123,N_625,N_356);
xnor U1124 (N_1124,N_896,N_285);
and U1125 (N_1125,N_362,N_968);
xor U1126 (N_1126,N_65,In_982);
nand U1127 (N_1127,N_1114,N_1060);
or U1128 (N_1128,N_74,N_1037);
xor U1129 (N_1129,In_852,N_1040);
xor U1130 (N_1130,In_532,N_475);
and U1131 (N_1131,N_618,N_843);
xor U1132 (N_1132,N_1119,In_979);
nand U1133 (N_1133,N_647,In_282);
nand U1134 (N_1134,N_837,N_817);
nor U1135 (N_1135,N_702,In_230);
or U1136 (N_1136,In_508,N_863);
nand U1137 (N_1137,N_120,In_1521);
nand U1138 (N_1138,In_1201,In_1472);
and U1139 (N_1139,In_1506,N_818);
and U1140 (N_1140,N_299,N_825);
xnor U1141 (N_1141,N_443,N_215);
or U1142 (N_1142,In_1775,N_1085);
nand U1143 (N_1143,N_552,N_520);
nand U1144 (N_1144,N_960,N_1102);
nor U1145 (N_1145,In_1033,N_392);
or U1146 (N_1146,N_905,In_705);
and U1147 (N_1147,In_1202,In_1586);
xor U1148 (N_1148,N_430,N_768);
or U1149 (N_1149,In_102,In_1839);
and U1150 (N_1150,In_904,N_169);
nor U1151 (N_1151,In_1452,In_395);
nor U1152 (N_1152,N_433,In_1645);
or U1153 (N_1153,In_1627,N_1029);
nor U1154 (N_1154,In_1420,In_1102);
and U1155 (N_1155,N_934,N_546);
and U1156 (N_1156,N_886,N_900);
nor U1157 (N_1157,N_980,In_1623);
and U1158 (N_1158,In_1866,N_795);
xor U1159 (N_1159,In_1568,N_534);
nand U1160 (N_1160,In_213,In_739);
xnor U1161 (N_1161,In_562,N_521);
nor U1162 (N_1162,In_1948,N_645);
or U1163 (N_1163,N_431,N_409);
nor U1164 (N_1164,N_731,In_1290);
or U1165 (N_1165,In_868,In_1498);
nand U1166 (N_1166,N_1076,N_547);
nor U1167 (N_1167,In_385,N_987);
xor U1168 (N_1168,N_180,N_1090);
xnor U1169 (N_1169,N_630,N_77);
or U1170 (N_1170,In_1009,N_404);
nand U1171 (N_1171,In_1120,N_1093);
nor U1172 (N_1172,N_540,N_1100);
nor U1173 (N_1173,N_286,N_1003);
and U1174 (N_1174,In_625,In_787);
nand U1175 (N_1175,In_1647,N_940);
or U1176 (N_1176,N_1010,In_894);
nor U1177 (N_1177,N_327,N_64);
nor U1178 (N_1178,N_1075,N_875);
and U1179 (N_1179,N_812,N_1030);
xor U1180 (N_1180,In_247,N_631);
nand U1181 (N_1181,N_536,N_1098);
nand U1182 (N_1182,N_1041,In_914);
xnor U1183 (N_1183,N_1116,In_1982);
nor U1184 (N_1184,N_1069,N_808);
nor U1185 (N_1185,N_864,In_623);
or U1186 (N_1186,N_796,In_631);
or U1187 (N_1187,N_823,N_1015);
xnor U1188 (N_1188,N_600,In_888);
nor U1189 (N_1189,N_1109,N_778);
xnor U1190 (N_1190,N_68,N_682);
nor U1191 (N_1191,N_1059,N_906);
or U1192 (N_1192,In_1200,N_933);
xnor U1193 (N_1193,N_918,In_1428);
and U1194 (N_1194,N_696,In_155);
and U1195 (N_1195,In_398,In_49);
xnor U1196 (N_1196,In_608,N_654);
xor U1197 (N_1197,N_746,N_962);
and U1198 (N_1198,N_919,N_44);
nor U1199 (N_1199,In_1617,In_1876);
nand U1200 (N_1200,In_1258,In_973);
and U1201 (N_1201,N_935,N_668);
nor U1202 (N_1202,N_298,N_1081);
or U1203 (N_1203,N_1017,N_318);
or U1204 (N_1204,N_1101,In_556);
nor U1205 (N_1205,N_661,In_1271);
xnor U1206 (N_1206,N_504,In_477);
and U1207 (N_1207,N_858,N_1047);
and U1208 (N_1208,N_381,N_86);
nand U1209 (N_1209,N_142,In_1924);
or U1210 (N_1210,In_966,In_391);
and U1211 (N_1211,In_1925,N_349);
nand U1212 (N_1212,In_1250,In_268);
nand U1213 (N_1213,In_813,N_730);
nand U1214 (N_1214,N_254,N_1024);
nor U1215 (N_1215,N_505,N_1012);
and U1216 (N_1216,N_833,N_1048);
nand U1217 (N_1217,N_1057,N_26);
nand U1218 (N_1218,N_152,In_239);
nor U1219 (N_1219,N_910,N_810);
xor U1220 (N_1220,N_773,In_1785);
nand U1221 (N_1221,N_865,In_1768);
or U1222 (N_1222,N_967,In_1425);
nor U1223 (N_1223,In_779,N_1027);
nor U1224 (N_1224,In_1132,In_244);
nor U1225 (N_1225,In_1849,N_619);
or U1226 (N_1226,N_924,In_1962);
and U1227 (N_1227,N_421,N_1110);
nor U1228 (N_1228,N_94,In_288);
or U1229 (N_1229,In_995,In_1234);
xnor U1230 (N_1230,N_1080,N_1088);
nor U1231 (N_1231,N_842,In_437);
or U1232 (N_1232,In_1046,In_1447);
and U1233 (N_1233,N_588,N_1050);
nand U1234 (N_1234,N_798,In_1044);
or U1235 (N_1235,In_1038,N_1072);
xnor U1236 (N_1236,In_933,In_231);
and U1237 (N_1237,In_1528,N_91);
and U1238 (N_1238,N_1062,In_1442);
nand U1239 (N_1239,N_1105,In_1263);
xnor U1240 (N_1240,In_1686,N_1094);
or U1241 (N_1241,N_712,In_1821);
or U1242 (N_1242,N_49,N_1099);
nand U1243 (N_1243,N_301,In_127);
nor U1244 (N_1244,In_807,N_657);
and U1245 (N_1245,In_1753,In_314);
and U1246 (N_1246,In_1364,In_197);
nand U1247 (N_1247,N_420,In_928);
nor U1248 (N_1248,N_466,N_382);
xnor U1249 (N_1249,In_1857,N_66);
nor U1250 (N_1250,In_1978,N_82);
or U1251 (N_1251,N_157,N_1018);
nor U1252 (N_1252,N_1011,N_581);
nand U1253 (N_1253,N_948,In_1415);
nand U1254 (N_1254,In_1970,N_29);
or U1255 (N_1255,N_371,In_1368);
xnor U1256 (N_1256,N_911,N_678);
and U1257 (N_1257,N_1035,In_1166);
or U1258 (N_1258,N_512,In_1613);
and U1259 (N_1259,N_35,N_533);
xnor U1260 (N_1260,In_1326,N_472);
nor U1261 (N_1261,N_1028,N_1083);
or U1262 (N_1262,N_1031,In_1159);
xor U1263 (N_1263,N_995,N_755);
nand U1264 (N_1264,In_1993,N_656);
nor U1265 (N_1265,N_651,N_1049);
or U1266 (N_1266,N_122,In_1381);
and U1267 (N_1267,N_857,In_607);
nor U1268 (N_1268,N_824,N_525);
nand U1269 (N_1269,In_648,N_269);
nand U1270 (N_1270,N_1104,In_164);
or U1271 (N_1271,In_886,In_206);
and U1272 (N_1272,In_205,In_1598);
nor U1273 (N_1273,N_67,In_757);
xnor U1274 (N_1274,In_1929,In_519);
nand U1275 (N_1275,N_202,In_930);
and U1276 (N_1276,N_867,In_1188);
or U1277 (N_1277,N_861,In_1175);
nor U1278 (N_1278,In_487,N_717);
xor U1279 (N_1279,N_841,N_1008);
nor U1280 (N_1280,N_1111,In_210);
and U1281 (N_1281,N_315,N_1178);
xnor U1282 (N_1282,N_719,In_1977);
xnor U1283 (N_1283,N_1218,N_1126);
or U1284 (N_1284,N_1179,In_248);
xnor U1285 (N_1285,N_1086,N_1089);
nor U1286 (N_1286,N_559,N_435);
nand U1287 (N_1287,In_1834,N_451);
nor U1288 (N_1288,In_1002,N_1279);
nor U1289 (N_1289,N_537,In_1101);
and U1290 (N_1290,N_5,N_147);
xor U1291 (N_1291,N_1264,N_1107);
nor U1292 (N_1292,N_683,In_1746);
nor U1293 (N_1293,In_1025,In_1816);
nor U1294 (N_1294,In_123,N_1092);
nand U1295 (N_1295,In_499,N_753);
nand U1296 (N_1296,N_528,In_255);
nand U1297 (N_1297,N_1124,In_1255);
xnor U1298 (N_1298,N_123,N_519);
xnor U1299 (N_1299,In_1618,In_363);
nand U1300 (N_1300,N_1265,N_19);
xnor U1301 (N_1301,In_1347,In_796);
nand U1302 (N_1302,N_966,In_1564);
nor U1303 (N_1303,N_648,In_168);
or U1304 (N_1304,N_175,N_728);
and U1305 (N_1305,N_422,N_704);
or U1306 (N_1306,In_1190,N_882);
or U1307 (N_1307,In_1146,N_227);
and U1308 (N_1308,N_1065,N_596);
nor U1309 (N_1309,N_1153,In_1455);
nor U1310 (N_1310,N_891,N_485);
and U1311 (N_1311,N_856,In_443);
nand U1312 (N_1312,In_1625,N_1212);
and U1313 (N_1313,N_828,N_821);
xnor U1314 (N_1314,N_515,In_5);
xnor U1315 (N_1315,N_603,N_239);
or U1316 (N_1316,In_1820,N_916);
or U1317 (N_1317,In_1504,N_691);
or U1318 (N_1318,In_377,N_1246);
and U1319 (N_1319,N_60,N_560);
xnor U1320 (N_1320,N_892,In_699);
and U1321 (N_1321,N_1054,N_969);
or U1322 (N_1322,N_790,N_927);
or U1323 (N_1323,In_304,N_539);
and U1324 (N_1324,In_591,N_164);
or U1325 (N_1325,In_184,N_1096);
nor U1326 (N_1326,N_1134,N_992);
or U1327 (N_1327,N_718,N_1034);
xnor U1328 (N_1328,In_373,N_1000);
xnor U1329 (N_1329,N_1164,N_244);
and U1330 (N_1330,N_1020,N_694);
nor U1331 (N_1331,N_146,N_1147);
nor U1332 (N_1332,N_1066,N_1159);
nor U1333 (N_1333,N_414,N_1023);
and U1334 (N_1334,N_1187,N_172);
xnor U1335 (N_1335,N_1239,N_178);
nor U1336 (N_1336,In_1349,N_920);
or U1337 (N_1337,N_979,N_1176);
nor U1338 (N_1338,N_985,N_666);
or U1339 (N_1339,N_497,N_637);
nand U1340 (N_1340,In_929,N_1122);
nor U1341 (N_1341,N_895,N_663);
and U1342 (N_1342,In_342,N_1204);
and U1343 (N_1343,N_1158,N_1112);
xor U1344 (N_1344,In_1519,N_970);
nor U1345 (N_1345,N_1195,N_1013);
nor U1346 (N_1346,N_990,N_1200);
nand U1347 (N_1347,N_1274,In_1622);
nor U1348 (N_1348,N_662,N_811);
nor U1349 (N_1349,N_716,N_802);
or U1350 (N_1350,N_1238,N_1262);
and U1351 (N_1351,In_716,N_1268);
nand U1352 (N_1352,N_872,N_469);
nand U1353 (N_1353,N_384,N_1273);
xor U1354 (N_1354,In_1859,N_545);
or U1355 (N_1355,N_564,In_1486);
nor U1356 (N_1356,N_1058,N_46);
xnor U1357 (N_1357,N_1056,N_1002);
xor U1358 (N_1358,In_790,N_819);
or U1359 (N_1359,In_464,N_1247);
or U1360 (N_1360,N_887,In_1567);
or U1361 (N_1361,In_201,N_1130);
nand U1362 (N_1362,N_722,N_1231);
xnor U1363 (N_1363,N_1137,N_1192);
nand U1364 (N_1364,N_490,N_1221);
or U1365 (N_1365,N_1266,N_791);
and U1366 (N_1366,In_1337,In_749);
and U1367 (N_1367,In_424,N_1148);
nand U1368 (N_1368,N_830,N_620);
or U1369 (N_1369,N_1103,N_1120);
and U1370 (N_1370,N_1194,N_492);
xor U1371 (N_1371,N_977,In_1888);
and U1372 (N_1372,N_999,N_1078);
and U1373 (N_1373,In_1274,N_1087);
nand U1374 (N_1374,In_417,N_195);
xor U1375 (N_1375,N_1210,N_1129);
nand U1376 (N_1376,N_839,In_1245);
nand U1377 (N_1377,N_1245,N_1278);
xnor U1378 (N_1378,N_1074,In_971);
nand U1379 (N_1379,N_395,N_732);
xor U1380 (N_1380,In_613,In_143);
nand U1381 (N_1381,N_1260,N_1225);
nor U1382 (N_1382,In_1301,N_1019);
xnor U1383 (N_1383,In_1781,N_904);
and U1384 (N_1384,In_529,In_882);
and U1385 (N_1385,N_1036,N_1052);
or U1386 (N_1386,N_659,In_993);
or U1387 (N_1387,In_1088,In_1015);
and U1388 (N_1388,In_1460,N_1097);
nand U1389 (N_1389,In_1585,N_1004);
or U1390 (N_1390,In_1426,N_1166);
or U1391 (N_1391,N_322,N_249);
nor U1392 (N_1392,In_985,N_860);
nor U1393 (N_1393,N_1146,N_1230);
xnor U1394 (N_1394,N_1154,N_909);
nor U1395 (N_1395,In_1338,N_1033);
nor U1396 (N_1396,N_577,N_622);
nand U1397 (N_1397,N_602,N_937);
nand U1398 (N_1398,In_171,N_1113);
or U1399 (N_1399,In_1014,N_623);
xnor U1400 (N_1400,N_1151,N_1121);
nand U1401 (N_1401,N_337,N_112);
xor U1402 (N_1402,N_871,In_1388);
nand U1403 (N_1403,N_319,In_768);
nor U1404 (N_1404,N_1079,In_1064);
and U1405 (N_1405,N_681,N_973);
xnor U1406 (N_1406,N_380,In_1399);
or U1407 (N_1407,N_1253,In_374);
and U1408 (N_1408,N_1149,N_218);
xor U1409 (N_1409,N_913,In_1328);
nand U1410 (N_1410,In_753,N_1188);
and U1411 (N_1411,N_838,N_1071);
or U1412 (N_1412,N_1001,N_709);
or U1413 (N_1413,In_620,N_780);
xnor U1414 (N_1414,N_959,N_513);
and U1415 (N_1415,N_1167,In_1160);
nor U1416 (N_1416,N_1138,N_1220);
and U1417 (N_1417,In_1148,N_996);
or U1418 (N_1418,N_1228,N_965);
or U1419 (N_1419,N_1203,N_1135);
and U1420 (N_1420,In_1457,In_1281);
or U1421 (N_1421,In_1054,N_954);
nand U1422 (N_1422,In_1669,N_579);
nor U1423 (N_1423,In_876,N_1155);
nor U1424 (N_1424,N_690,N_1132);
xnor U1425 (N_1425,N_393,In_1597);
nor U1426 (N_1426,N_986,In_1530);
nor U1427 (N_1427,In_141,N_699);
or U1428 (N_1428,N_1235,N_1162);
nor U1429 (N_1429,In_962,N_978);
nor U1430 (N_1430,In_1745,N_93);
nor U1431 (N_1431,N_982,N_1095);
nand U1432 (N_1432,N_1181,N_1250);
nor U1433 (N_1433,N_464,N_1263);
and U1434 (N_1434,In_1483,N_673);
or U1435 (N_1435,N_949,N_1209);
xor U1436 (N_1436,N_777,N_78);
xnor U1437 (N_1437,In_1435,N_807);
nand U1438 (N_1438,In_1837,In_103);
and U1439 (N_1439,In_334,In_663);
nand U1440 (N_1440,In_1196,In_1211);
nand U1441 (N_1441,In_456,N_1258);
or U1442 (N_1442,N_1142,N_1325);
nand U1443 (N_1443,N_1302,N_214);
nor U1444 (N_1444,N_1319,N_1419);
nand U1445 (N_1445,N_1172,N_1217);
nand U1446 (N_1446,N_1044,N_42);
xnor U1447 (N_1447,N_1276,In_1596);
nand U1448 (N_1448,N_1417,N_441);
nor U1449 (N_1449,N_1042,N_1385);
or U1450 (N_1450,N_168,In_266);
nand U1451 (N_1451,In_788,N_742);
and U1452 (N_1452,In_1287,N_502);
xor U1453 (N_1453,N_658,N_1389);
xor U1454 (N_1454,N_1367,N_193);
or U1455 (N_1455,N_1039,N_1401);
nor U1456 (N_1456,N_1261,In_1583);
or U1457 (N_1457,N_1369,N_878);
nand U1458 (N_1458,N_915,N_565);
nand U1459 (N_1459,N_607,In_803);
nor U1460 (N_1460,In_1963,N_688);
and U1461 (N_1461,N_1371,N_1428);
and U1462 (N_1462,N_991,In_1581);
nand U1463 (N_1463,N_1377,N_1334);
nor U1464 (N_1464,In_39,In_413);
nor U1465 (N_1465,N_922,N_1084);
nor U1466 (N_1466,N_1287,N_1414);
and U1467 (N_1467,N_1277,N_894);
xnor U1468 (N_1468,In_351,N_1421);
and U1469 (N_1469,N_1418,N_885);
xor U1470 (N_1470,N_1310,N_1393);
nor U1471 (N_1471,N_686,N_1182);
xnor U1472 (N_1472,N_1390,N_749);
nand U1473 (N_1473,N_1423,N_375);
nor U1474 (N_1474,N_1222,N_806);
nor U1475 (N_1475,N_1395,In_1307);
xor U1476 (N_1476,In_151,N_850);
or U1477 (N_1477,N_1205,N_1254);
nor U1478 (N_1478,N_626,In_755);
xor U1479 (N_1479,N_549,N_1244);
xor U1480 (N_1480,N_1366,N_1326);
nand U1481 (N_1481,N_357,N_1282);
and U1482 (N_1482,N_981,In_670);
and U1483 (N_1483,N_816,N_1236);
or U1484 (N_1484,N_1297,N_201);
nor U1485 (N_1485,In_482,In_581);
or U1486 (N_1486,N_1295,N_1387);
or U1487 (N_1487,In_1744,In_185);
xnor U1488 (N_1488,N_1354,N_1426);
xor U1489 (N_1489,N_1160,N_200);
or U1490 (N_1490,N_340,In_545);
xnor U1491 (N_1491,In_219,N_1343);
nor U1492 (N_1492,N_947,N_1193);
nor U1493 (N_1493,N_1317,N_210);
or U1494 (N_1494,N_1070,N_1284);
and U1495 (N_1495,N_952,N_1352);
or U1496 (N_1496,N_1180,N_1198);
nand U1497 (N_1497,N_1345,N_1252);
xor U1498 (N_1498,N_1067,N_1373);
or U1499 (N_1499,N_1073,In_839);
xor U1500 (N_1500,N_1234,N_1398);
or U1501 (N_1501,N_554,N_1270);
xnor U1502 (N_1502,N_770,N_964);
and U1503 (N_1503,In_1323,N_955);
nand U1504 (N_1504,In_1699,N_1108);
nand U1505 (N_1505,N_1427,N_1143);
nor U1506 (N_1506,N_903,In_422);
and U1507 (N_1507,N_971,N_1305);
xnor U1508 (N_1508,In_19,N_800);
or U1509 (N_1509,N_1171,N_1224);
or U1510 (N_1510,N_930,N_929);
nand U1511 (N_1511,N_418,In_1207);
or U1512 (N_1512,N_740,N_1063);
or U1513 (N_1513,N_1243,N_1051);
xnor U1514 (N_1514,N_106,N_1006);
nor U1515 (N_1515,In_713,N_555);
or U1516 (N_1516,N_243,N_1301);
nand U1517 (N_1517,N_1360,N_1077);
xor U1518 (N_1518,In_222,In_1919);
and U1519 (N_1519,N_439,N_1351);
or U1520 (N_1520,In_575,N_984);
nand U1521 (N_1521,In_781,N_1370);
nor U1522 (N_1522,In_1163,N_705);
nor U1523 (N_1523,N_1242,N_1123);
xor U1524 (N_1524,N_1091,N_669);
or U1525 (N_1525,N_939,N_1420);
and U1526 (N_1526,N_40,N_1163);
nand U1527 (N_1527,N_974,N_1437);
and U1528 (N_1528,N_1196,N_253);
or U1529 (N_1529,N_376,N_1005);
or U1530 (N_1530,N_1299,N_1298);
or U1531 (N_1531,N_1237,N_1206);
or U1532 (N_1532,N_1410,N_1207);
and U1533 (N_1533,In_1321,N_1378);
xnor U1534 (N_1534,N_1346,In_1168);
nor U1535 (N_1535,N_1199,N_1140);
nor U1536 (N_1536,N_312,N_1332);
or U1537 (N_1537,N_1355,In_25);
or U1538 (N_1538,N_993,In_1706);
or U1539 (N_1539,In_726,N_1311);
and U1540 (N_1540,N_1251,N_1328);
nor U1541 (N_1541,N_1304,In_18);
nand U1542 (N_1542,N_1053,N_1292);
xor U1543 (N_1543,N_1327,N_1359);
xor U1544 (N_1544,N_1032,N_1406);
or U1545 (N_1545,N_1394,N_1358);
and U1546 (N_1546,N_71,In_1246);
nor U1547 (N_1547,N_1318,N_1061);
and U1548 (N_1548,N_1380,In_1485);
nor U1549 (N_1549,N_1430,In_14);
nand U1550 (N_1550,N_1021,In_901);
nand U1551 (N_1551,In_1606,In_110);
nor U1552 (N_1552,N_1339,N_1342);
and U1553 (N_1553,N_1240,N_1219);
nor U1554 (N_1554,N_1141,N_1347);
or U1555 (N_1555,N_326,N_988);
nor U1556 (N_1556,In_1150,N_782);
nand U1557 (N_1557,N_1055,N_827);
or U1558 (N_1558,N_1333,N_1300);
and U1559 (N_1559,N_1381,In_3);
xnor U1560 (N_1560,N_1214,N_1232);
nor U1561 (N_1561,N_1257,N_471);
nand U1562 (N_1562,N_1431,N_1226);
nand U1563 (N_1563,In_1454,N_983);
xnor U1564 (N_1564,In_1269,N_1173);
xor U1565 (N_1565,N_760,N_1127);
and U1566 (N_1566,N_1115,In_714);
nor U1567 (N_1567,In_1085,N_1014);
xor U1568 (N_1568,N_606,N_1269);
and U1569 (N_1569,In_926,N_1405);
or U1570 (N_1570,N_1324,N_1275);
nor U1571 (N_1571,In_1139,In_1986);
nand U1572 (N_1572,In_850,N_1227);
nor U1573 (N_1573,N_144,N_1336);
xnor U1574 (N_1574,N_961,In_1097);
nor U1575 (N_1575,N_845,In_1333);
or U1576 (N_1576,In_1342,N_1280);
nor U1577 (N_1577,N_1335,N_1329);
or U1578 (N_1578,N_280,N_1384);
and U1579 (N_1579,N_1314,N_1357);
xor U1580 (N_1580,N_1285,N_1043);
nand U1581 (N_1581,N_1216,N_455);
xnor U1582 (N_1582,N_1286,N_1340);
or U1583 (N_1583,In_585,N_1185);
nand U1584 (N_1584,N_963,N_339);
xnor U1585 (N_1585,In_967,In_328);
xor U1586 (N_1586,In_883,In_517);
nor U1587 (N_1587,N_1296,N_1368);
xor U1588 (N_1588,N_1408,N_571);
nor U1589 (N_1589,N_587,In_1171);
or U1590 (N_1590,In_725,N_912);
nand U1591 (N_1591,N_456,N_1293);
and U1592 (N_1592,N_447,N_518);
nand U1593 (N_1593,In_1979,In_1724);
nor U1594 (N_1594,N_1190,N_1372);
nand U1595 (N_1595,In_165,N_1241);
xnor U1596 (N_1596,In_866,In_214);
xor U1597 (N_1597,N_881,N_1379);
nand U1598 (N_1598,N_509,N_1399);
nand U1599 (N_1599,N_1400,N_1392);
nand U1600 (N_1600,In_728,N_1169);
nand U1601 (N_1601,In_1480,N_1566);
nor U1602 (N_1602,N_1315,N_1575);
or U1603 (N_1603,N_1466,N_1559);
xnor U1604 (N_1604,N_295,N_1561);
nor U1605 (N_1605,In_1228,N_70);
or U1606 (N_1606,N_1552,N_1579);
nand U1607 (N_1607,N_1474,N_1525);
or U1608 (N_1608,N_1568,N_1223);
or U1609 (N_1609,N_432,In_1453);
or U1610 (N_1610,In_553,N_1007);
nor U1611 (N_1611,N_1567,N_1521);
and U1612 (N_1612,N_1577,N_1433);
or U1613 (N_1613,N_1551,N_621);
nand U1614 (N_1614,N_1152,N_1547);
xor U1615 (N_1615,N_1183,N_1350);
and U1616 (N_1616,N_1288,N_1593);
nor U1617 (N_1617,N_1344,N_140);
nor U1618 (N_1618,N_1524,In_150);
nand U1619 (N_1619,N_385,N_198);
nor U1620 (N_1620,N_1233,N_1449);
nand U1621 (N_1621,N_1177,N_938);
nor U1622 (N_1622,N_1541,N_1469);
nand U1623 (N_1623,N_1313,N_997);
xor U1624 (N_1624,N_30,N_1571);
xnor U1625 (N_1625,N_809,N_246);
xnor U1626 (N_1626,N_1538,N_1503);
nand U1627 (N_1627,N_1478,N_1506);
nor U1628 (N_1628,N_1184,N_1249);
nor U1629 (N_1629,N_355,N_1492);
nand U1630 (N_1630,N_1472,N_583);
or U1631 (N_1631,N_884,In_325);
and U1632 (N_1632,N_1505,N_1479);
nand U1633 (N_1633,N_1527,N_1386);
nor U1634 (N_1634,N_1026,N_1404);
xnor U1635 (N_1635,N_958,N_1485);
nor U1636 (N_1636,In_1079,N_1501);
nor U1637 (N_1637,N_1553,N_1022);
and U1638 (N_1638,N_1482,N_1533);
xnor U1639 (N_1639,In_1499,N_1499);
xnor U1640 (N_1640,N_1403,N_840);
or U1641 (N_1641,N_1460,N_1434);
and U1642 (N_1642,N_1570,In_1458);
and U1643 (N_1643,In_679,N_1082);
nor U1644 (N_1644,N_1563,N_1374);
xor U1645 (N_1645,N_1530,N_396);
nand U1646 (N_1646,N_1456,N_989);
xor U1647 (N_1647,N_1397,N_813);
or U1648 (N_1648,In_1893,N_608);
nor U1649 (N_1649,N_956,N_1496);
xor U1650 (N_1650,N_1586,N_1450);
xor U1651 (N_1651,N_1560,N_1463);
or U1652 (N_1652,N_1447,N_925);
or U1653 (N_1653,In_465,N_849);
nand U1654 (N_1654,N_1536,In_1587);
nand U1655 (N_1655,N_1520,N_1145);
nand U1656 (N_1656,N_1045,N_733);
or U1657 (N_1657,N_1307,N_1451);
nand U1658 (N_1658,N_650,N_1136);
nor U1659 (N_1659,N_1489,N_1556);
and U1660 (N_1660,In_615,N_1259);
or U1661 (N_1661,In_1822,N_1457);
and U1662 (N_1662,N_1539,N_1375);
nand U1663 (N_1663,N_90,N_1446);
xor U1664 (N_1664,N_1133,N_1312);
nor U1665 (N_1665,N_1455,In_260);
xnor U1666 (N_1666,N_1581,In_1429);
and U1667 (N_1667,N_1550,In_460);
or U1668 (N_1668,N_1522,N_1445);
and U1669 (N_1669,N_1598,N_1439);
or U1670 (N_1670,N_1046,N_1510);
nand U1671 (N_1671,N_1583,N_1519);
nor U1672 (N_1672,N_1321,N_1558);
nor U1673 (N_1673,N_1412,In_1662);
and U1674 (N_1674,N_1248,N_408);
xor U1675 (N_1675,N_1511,N_1118);
and U1676 (N_1676,N_468,N_1106);
or U1677 (N_1677,N_1376,N_972);
nand U1678 (N_1678,N_1415,N_1442);
or U1679 (N_1679,N_1125,N_1497);
nand U1680 (N_1680,N_1201,N_1425);
nor U1681 (N_1681,N_1599,N_1330);
nand U1682 (N_1682,N_1576,N_1422);
or U1683 (N_1683,N_1544,N_975);
nor U1684 (N_1684,N_556,N_1471);
and U1685 (N_1685,N_1349,In_1878);
and U1686 (N_1686,N_1453,N_1484);
or U1687 (N_1687,N_166,In_1041);
xnor U1688 (N_1688,N_1543,N_1208);
and U1689 (N_1689,N_55,N_1267);
nor U1690 (N_1690,N_1476,N_1498);
or U1691 (N_1691,N_642,N_1131);
nor U1692 (N_1692,N_1585,In_1819);
and U1693 (N_1693,N_998,N_943);
nor U1694 (N_1694,N_1435,N_1569);
and U1695 (N_1695,N_595,N_1488);
nand U1696 (N_1696,N_976,N_1564);
or U1697 (N_1697,N_1362,N_1572);
xor U1698 (N_1698,N_1391,In_1232);
nor U1699 (N_1699,N_1490,N_1416);
xor U1700 (N_1700,N_1500,N_1363);
xnor U1701 (N_1701,N_826,N_1483);
xor U1702 (N_1702,N_1429,N_1465);
and U1703 (N_1703,N_876,In_727);
nand U1704 (N_1704,N_1454,N_1139);
or U1705 (N_1705,N_1117,N_1331);
and U1706 (N_1706,N_1215,N_1441);
nor U1707 (N_1707,N_1150,N_926);
xnor U1708 (N_1708,In_393,N_1555);
and U1709 (N_1709,N_1170,N_1409);
xor U1710 (N_1710,N_1495,N_1588);
and U1711 (N_1711,N_1291,N_1283);
nand U1712 (N_1712,N_1502,N_527);
nor U1713 (N_1713,N_1303,N_1591);
or U1714 (N_1714,N_1597,N_1548);
and U1715 (N_1715,N_1316,N_1144);
nand U1716 (N_1716,N_1481,In_921);
xnor U1717 (N_1717,N_1068,N_1475);
nand U1718 (N_1718,N_1213,N_1595);
xor U1719 (N_1719,N_1573,N_1348);
or U1720 (N_1720,N_1534,N_1168);
and U1721 (N_1721,N_1590,N_1229);
nor U1722 (N_1722,N_1290,N_323);
and U1723 (N_1723,In_619,N_1289);
and U1724 (N_1724,In_1206,N_1424);
and U1725 (N_1725,N_1594,N_1523);
xor U1726 (N_1726,In_597,N_1353);
xnor U1727 (N_1727,N_1516,N_1540);
and U1728 (N_1728,N_1582,N_1584);
or U1729 (N_1729,In_858,N_1322);
nand U1730 (N_1730,N_877,N_1128);
and U1731 (N_1731,N_1197,In_274);
nor U1732 (N_1732,N_1535,N_1512);
and U1733 (N_1733,N_1477,N_1459);
nor U1734 (N_1734,N_781,N_1514);
nand U1735 (N_1735,N_1191,N_1009);
nand U1736 (N_1736,N_1596,N_1356);
nand U1737 (N_1737,N_1526,N_150);
xnor U1738 (N_1738,N_1281,In_1632);
and U1739 (N_1739,N_1562,N_1407);
or U1740 (N_1740,In_1549,N_1271);
nor U1741 (N_1741,N_1411,N_1388);
and U1742 (N_1742,N_1189,N_1532);
or U1743 (N_1743,N_836,N_1383);
nand U1744 (N_1744,N_1473,N_1175);
and U1745 (N_1745,N_1491,N_1578);
nor U1746 (N_1746,N_1587,N_1468);
xor U1747 (N_1747,N_1504,N_1323);
xor U1748 (N_1748,N_1557,N_1529);
nor U1749 (N_1749,N_771,N_1507);
nand U1750 (N_1750,In_1799,In_891);
nand U1751 (N_1751,N_1306,N_1309);
and U1752 (N_1752,N_815,N_113);
or U1753 (N_1753,N_1444,N_1546);
xnor U1754 (N_1754,N_859,In_976);
and U1755 (N_1755,N_1493,N_1574);
and U1756 (N_1756,N_1438,N_1589);
nand U1757 (N_1757,In_386,In_1511);
xnor U1758 (N_1758,N_1016,N_1025);
xnor U1759 (N_1759,N_873,N_1487);
xnor U1760 (N_1760,N_1674,N_1687);
nand U1761 (N_1761,N_1600,N_1699);
or U1762 (N_1762,N_1714,N_1645);
xor U1763 (N_1763,N_1603,In_616);
and U1764 (N_1764,N_1663,N_1727);
or U1765 (N_1765,N_1725,N_1402);
nor U1766 (N_1766,In_666,N_1542);
and U1767 (N_1767,N_1676,N_1662);
or U1768 (N_1768,N_1700,N_1728);
or U1769 (N_1769,N_1604,N_1580);
nand U1770 (N_1770,N_1341,N_1664);
and U1771 (N_1771,N_1462,N_1592);
xnor U1772 (N_1772,N_1684,N_1528);
nor U1773 (N_1773,N_1517,N_1156);
or U1774 (N_1774,N_1690,N_1165);
or U1775 (N_1775,N_1461,N_1622);
nor U1776 (N_1776,N_1448,N_1659);
xnor U1777 (N_1777,N_1643,N_1753);
and U1778 (N_1778,N_1670,N_1715);
nor U1779 (N_1779,N_1513,N_1733);
nand U1780 (N_1780,N_1653,N_1726);
nor U1781 (N_1781,N_641,N_1689);
and U1782 (N_1782,N_1480,N_1731);
or U1783 (N_1783,N_1612,N_1458);
and U1784 (N_1784,N_1703,N_1706);
nand U1785 (N_1785,N_1618,N_734);
or U1786 (N_1786,N_1470,N_1629);
nand U1787 (N_1787,N_1382,N_1364);
nor U1788 (N_1788,N_1650,N_1695);
nor U1789 (N_1789,N_1337,In_707);
xor U1790 (N_1790,N_1632,N_1320);
or U1791 (N_1791,N_1038,N_1696);
and U1792 (N_1792,N_1735,N_994);
nor U1793 (N_1793,In_964,N_1608);
or U1794 (N_1794,N_1723,N_1759);
or U1795 (N_1795,N_1744,N_1758);
nor U1796 (N_1796,N_1606,N_1702);
or U1797 (N_1797,N_1602,N_1338);
nand U1798 (N_1798,N_1736,N_1644);
xnor U1799 (N_1799,N_1657,N_1634);
nor U1800 (N_1800,N_1742,N_1646);
nand U1801 (N_1801,In_1445,N_1545);
nand U1802 (N_1802,N_1671,N_1704);
and U1803 (N_1803,N_1623,N_1620);
nand U1804 (N_1804,N_1617,N_1722);
and U1805 (N_1805,N_1494,N_1294);
nand U1806 (N_1806,N_1636,N_1633);
and U1807 (N_1807,In_827,N_1724);
and U1808 (N_1808,N_1607,N_1256);
nand U1809 (N_1809,N_1751,N_1668);
nor U1810 (N_1810,N_1440,N_1713);
xor U1811 (N_1811,N_1716,N_1443);
nand U1812 (N_1812,In_1788,N_1486);
xnor U1813 (N_1813,N_1202,N_1752);
or U1814 (N_1814,N_1757,N_1211);
nand U1815 (N_1815,N_1616,N_1665);
nand U1816 (N_1816,N_1549,N_1678);
nand U1817 (N_1817,N_1515,In_267);
or U1818 (N_1818,N_1452,N_1749);
xor U1819 (N_1819,N_1648,N_1693);
or U1820 (N_1820,N_1565,N_1747);
xnor U1821 (N_1821,N_1614,N_1732);
or U1822 (N_1822,N_1756,In_874);
or U1823 (N_1823,N_1365,N_1729);
nor U1824 (N_1824,N_1673,N_1709);
nand U1825 (N_1825,N_1361,N_1755);
and U1826 (N_1826,N_416,N_1711);
nand U1827 (N_1827,N_1682,N_1750);
nor U1828 (N_1828,N_1683,N_703);
or U1829 (N_1829,N_1675,N_1672);
xor U1830 (N_1830,N_1660,N_1619);
nand U1831 (N_1831,N_1688,N_1685);
xnor U1832 (N_1832,N_1679,N_1649);
xnor U1833 (N_1833,N_1677,N_1720);
and U1834 (N_1834,N_1705,N_1509);
nand U1835 (N_1835,N_1638,N_1694);
xnor U1836 (N_1836,N_1508,N_1743);
nand U1837 (N_1837,In_1192,N_1748);
and U1838 (N_1838,N_1698,N_1681);
xor U1839 (N_1839,N_1719,N_1745);
and U1840 (N_1840,N_1746,N_1654);
nor U1841 (N_1841,N_1413,N_1436);
or U1842 (N_1842,N_1717,N_1655);
nor U1843 (N_1843,N_1186,N_1721);
nor U1844 (N_1844,N_1624,N_1628);
xnor U1845 (N_1845,N_1064,N_1531);
xnor U1846 (N_1846,N_1272,N_1641);
or U1847 (N_1847,N_1601,N_1635);
and U1848 (N_1848,N_1626,N_1396);
nand U1849 (N_1849,N_1518,N_426);
and U1850 (N_1850,N_1710,N_1652);
nand U1851 (N_1851,N_1308,In_1022);
nand U1852 (N_1852,N_1537,N_1692);
xor U1853 (N_1853,N_1754,N_1464);
or U1854 (N_1854,N_1707,N_1730);
xor U1855 (N_1855,N_1432,N_1609);
nor U1856 (N_1856,N_1630,N_1627);
nand U1857 (N_1857,N_1467,N_1738);
xor U1858 (N_1858,N_1554,N_1691);
nand U1859 (N_1859,N_1640,N_1610);
nor U1860 (N_1860,N_1686,N_1680);
and U1861 (N_1861,N_756,N_1157);
xnor U1862 (N_1862,N_1712,N_1697);
nand U1863 (N_1863,N_1611,N_1613);
nand U1864 (N_1864,N_1666,N_1631);
and U1865 (N_1865,In_1845,N_1642);
xor U1866 (N_1866,N_1708,N_1161);
or U1867 (N_1867,N_1174,N_1647);
xnor U1868 (N_1868,N_1255,N_1637);
nor U1869 (N_1869,N_1737,N_1625);
nand U1870 (N_1870,N_1734,N_1615);
nand U1871 (N_1871,N_1669,N_1605);
nand U1872 (N_1872,N_47,N_1661);
or U1873 (N_1873,N_890,N_1621);
nand U1874 (N_1874,N_1656,N_1701);
xnor U1875 (N_1875,N_1651,N_1718);
or U1876 (N_1876,N_453,N_1658);
or U1877 (N_1877,N_1667,N_1741);
nand U1878 (N_1878,In_1270,N_1740);
nor U1879 (N_1879,N_1639,N_1739);
xor U1880 (N_1880,N_1718,N_1721);
or U1881 (N_1881,N_1625,N_1655);
nor U1882 (N_1882,N_1592,N_1744);
nor U1883 (N_1883,N_1341,N_1726);
nand U1884 (N_1884,N_1448,N_1720);
and U1885 (N_1885,N_1622,N_1757);
nor U1886 (N_1886,N_1754,N_1618);
xor U1887 (N_1887,N_1722,N_1620);
nor U1888 (N_1888,N_1537,N_1161);
or U1889 (N_1889,N_1432,N_1703);
nand U1890 (N_1890,N_1756,N_1436);
or U1891 (N_1891,N_1635,N_1670);
nor U1892 (N_1892,N_47,N_1629);
and U1893 (N_1893,N_1687,N_1692);
xnor U1894 (N_1894,N_1683,N_1165);
and U1895 (N_1895,In_827,In_707);
nor U1896 (N_1896,N_1461,N_47);
xnor U1897 (N_1897,N_1648,N_1629);
or U1898 (N_1898,N_1608,N_1565);
and U1899 (N_1899,N_1634,N_1627);
or U1900 (N_1900,N_1724,N_1611);
or U1901 (N_1901,N_1664,N_1636);
xnor U1902 (N_1902,N_1613,N_1698);
nor U1903 (N_1903,N_1681,N_1643);
xor U1904 (N_1904,N_1732,N_1753);
nand U1905 (N_1905,N_1718,N_1186);
xnor U1906 (N_1906,N_1725,N_1732);
or U1907 (N_1907,N_1338,N_1657);
nand U1908 (N_1908,N_1603,N_1174);
or U1909 (N_1909,N_1724,N_1630);
xnor U1910 (N_1910,N_1565,N_1715);
and U1911 (N_1911,N_1728,N_47);
nand U1912 (N_1912,N_1660,N_1255);
xor U1913 (N_1913,N_1679,N_1639);
xnor U1914 (N_1914,N_1679,N_1211);
nand U1915 (N_1915,N_1639,N_1742);
nand U1916 (N_1916,N_1650,N_1704);
xor U1917 (N_1917,N_1681,N_1739);
nor U1918 (N_1918,N_1666,N_1733);
nor U1919 (N_1919,N_1713,N_1755);
and U1920 (N_1920,N_1829,N_1854);
and U1921 (N_1921,N_1910,N_1819);
or U1922 (N_1922,N_1785,N_1846);
and U1923 (N_1923,N_1885,N_1868);
and U1924 (N_1924,N_1828,N_1840);
and U1925 (N_1925,N_1895,N_1864);
or U1926 (N_1926,N_1769,N_1865);
nor U1927 (N_1927,N_1914,N_1781);
or U1928 (N_1928,N_1812,N_1842);
nor U1929 (N_1929,N_1909,N_1847);
or U1930 (N_1930,N_1918,N_1782);
nand U1931 (N_1931,N_1815,N_1900);
nor U1932 (N_1932,N_1867,N_1818);
nor U1933 (N_1933,N_1904,N_1767);
xor U1934 (N_1934,N_1859,N_1771);
or U1935 (N_1935,N_1795,N_1858);
xor U1936 (N_1936,N_1913,N_1882);
nor U1937 (N_1937,N_1830,N_1856);
and U1938 (N_1938,N_1894,N_1853);
xnor U1939 (N_1939,N_1765,N_1899);
and U1940 (N_1940,N_1779,N_1902);
nor U1941 (N_1941,N_1878,N_1788);
or U1942 (N_1942,N_1875,N_1850);
nor U1943 (N_1943,N_1898,N_1763);
nand U1944 (N_1944,N_1770,N_1778);
nand U1945 (N_1945,N_1766,N_1820);
or U1946 (N_1946,N_1863,N_1896);
or U1947 (N_1947,N_1805,N_1857);
or U1948 (N_1948,N_1794,N_1919);
or U1949 (N_1949,N_1883,N_1817);
nor U1950 (N_1950,N_1762,N_1816);
or U1951 (N_1951,N_1844,N_1912);
nor U1952 (N_1952,N_1821,N_1905);
and U1953 (N_1953,N_1803,N_1790);
or U1954 (N_1954,N_1903,N_1824);
xnor U1955 (N_1955,N_1814,N_1907);
nor U1956 (N_1956,N_1887,N_1897);
and U1957 (N_1957,N_1901,N_1884);
nand U1958 (N_1958,N_1841,N_1836);
nor U1959 (N_1959,N_1825,N_1906);
and U1960 (N_1960,N_1873,N_1775);
nor U1961 (N_1961,N_1862,N_1843);
or U1962 (N_1962,N_1886,N_1776);
nor U1963 (N_1963,N_1800,N_1796);
nand U1964 (N_1964,N_1813,N_1806);
xnor U1965 (N_1965,N_1772,N_1768);
nand U1966 (N_1966,N_1877,N_1879);
nand U1967 (N_1967,N_1789,N_1801);
or U1968 (N_1968,N_1872,N_1783);
xor U1969 (N_1969,N_1845,N_1874);
or U1970 (N_1970,N_1798,N_1786);
and U1971 (N_1971,N_1797,N_1791);
or U1972 (N_1972,N_1881,N_1851);
xor U1973 (N_1973,N_1871,N_1861);
and U1974 (N_1974,N_1826,N_1852);
xor U1975 (N_1975,N_1823,N_1911);
nor U1976 (N_1976,N_1839,N_1793);
xor U1977 (N_1977,N_1833,N_1869);
or U1978 (N_1978,N_1774,N_1827);
and U1979 (N_1979,N_1888,N_1804);
or U1980 (N_1980,N_1811,N_1761);
or U1981 (N_1981,N_1870,N_1822);
and U1982 (N_1982,N_1908,N_1838);
nand U1983 (N_1983,N_1809,N_1834);
xor U1984 (N_1984,N_1917,N_1889);
nor U1985 (N_1985,N_1835,N_1777);
or U1986 (N_1986,N_1915,N_1837);
nand U1987 (N_1987,N_1876,N_1807);
or U1988 (N_1988,N_1784,N_1773);
or U1989 (N_1989,N_1848,N_1810);
nor U1990 (N_1990,N_1891,N_1832);
nor U1991 (N_1991,N_1808,N_1799);
nor U1992 (N_1992,N_1890,N_1764);
or U1993 (N_1993,N_1892,N_1831);
or U1994 (N_1994,N_1760,N_1860);
and U1995 (N_1995,N_1866,N_1792);
and U1996 (N_1996,N_1787,N_1916);
and U1997 (N_1997,N_1802,N_1880);
nand U1998 (N_1998,N_1893,N_1780);
nand U1999 (N_1999,N_1849,N_1855);
and U2000 (N_2000,N_1774,N_1877);
nand U2001 (N_2001,N_1844,N_1868);
and U2002 (N_2002,N_1878,N_1835);
and U2003 (N_2003,N_1877,N_1893);
nand U2004 (N_2004,N_1894,N_1918);
or U2005 (N_2005,N_1880,N_1799);
or U2006 (N_2006,N_1900,N_1791);
or U2007 (N_2007,N_1846,N_1889);
xor U2008 (N_2008,N_1781,N_1883);
or U2009 (N_2009,N_1881,N_1850);
and U2010 (N_2010,N_1775,N_1815);
and U2011 (N_2011,N_1893,N_1816);
nor U2012 (N_2012,N_1903,N_1891);
or U2013 (N_2013,N_1869,N_1804);
xnor U2014 (N_2014,N_1806,N_1837);
nand U2015 (N_2015,N_1892,N_1846);
nand U2016 (N_2016,N_1826,N_1772);
nor U2017 (N_2017,N_1775,N_1795);
nand U2018 (N_2018,N_1825,N_1782);
nand U2019 (N_2019,N_1803,N_1786);
xor U2020 (N_2020,N_1877,N_1790);
nand U2021 (N_2021,N_1763,N_1901);
or U2022 (N_2022,N_1798,N_1902);
nand U2023 (N_2023,N_1789,N_1848);
nor U2024 (N_2024,N_1892,N_1903);
and U2025 (N_2025,N_1872,N_1794);
and U2026 (N_2026,N_1880,N_1861);
and U2027 (N_2027,N_1867,N_1842);
nand U2028 (N_2028,N_1798,N_1763);
nor U2029 (N_2029,N_1909,N_1813);
or U2030 (N_2030,N_1844,N_1864);
xor U2031 (N_2031,N_1852,N_1818);
nor U2032 (N_2032,N_1893,N_1807);
xor U2033 (N_2033,N_1883,N_1787);
and U2034 (N_2034,N_1900,N_1777);
nand U2035 (N_2035,N_1887,N_1777);
xnor U2036 (N_2036,N_1899,N_1808);
or U2037 (N_2037,N_1805,N_1790);
nor U2038 (N_2038,N_1827,N_1895);
nand U2039 (N_2039,N_1805,N_1854);
xnor U2040 (N_2040,N_1799,N_1810);
xnor U2041 (N_2041,N_1905,N_1808);
or U2042 (N_2042,N_1827,N_1897);
xnor U2043 (N_2043,N_1892,N_1911);
or U2044 (N_2044,N_1777,N_1765);
and U2045 (N_2045,N_1824,N_1852);
and U2046 (N_2046,N_1902,N_1919);
nor U2047 (N_2047,N_1814,N_1904);
or U2048 (N_2048,N_1843,N_1795);
and U2049 (N_2049,N_1902,N_1847);
xor U2050 (N_2050,N_1883,N_1914);
and U2051 (N_2051,N_1770,N_1915);
nand U2052 (N_2052,N_1794,N_1867);
nor U2053 (N_2053,N_1871,N_1815);
nand U2054 (N_2054,N_1832,N_1833);
nand U2055 (N_2055,N_1786,N_1897);
and U2056 (N_2056,N_1889,N_1833);
or U2057 (N_2057,N_1760,N_1787);
or U2058 (N_2058,N_1772,N_1867);
xnor U2059 (N_2059,N_1861,N_1856);
xnor U2060 (N_2060,N_1842,N_1832);
xnor U2061 (N_2061,N_1814,N_1801);
or U2062 (N_2062,N_1848,N_1879);
xor U2063 (N_2063,N_1833,N_1843);
nand U2064 (N_2064,N_1828,N_1887);
xnor U2065 (N_2065,N_1789,N_1790);
xnor U2066 (N_2066,N_1878,N_1786);
nor U2067 (N_2067,N_1868,N_1850);
and U2068 (N_2068,N_1790,N_1899);
or U2069 (N_2069,N_1877,N_1917);
or U2070 (N_2070,N_1843,N_1821);
and U2071 (N_2071,N_1912,N_1807);
xnor U2072 (N_2072,N_1795,N_1875);
xor U2073 (N_2073,N_1779,N_1804);
nand U2074 (N_2074,N_1790,N_1881);
xor U2075 (N_2075,N_1830,N_1771);
and U2076 (N_2076,N_1833,N_1845);
nor U2077 (N_2077,N_1820,N_1772);
and U2078 (N_2078,N_1849,N_1782);
nor U2079 (N_2079,N_1889,N_1882);
xor U2080 (N_2080,N_1982,N_2042);
xor U2081 (N_2081,N_2051,N_2014);
and U2082 (N_2082,N_1931,N_1999);
xnor U2083 (N_2083,N_2011,N_1928);
xnor U2084 (N_2084,N_2038,N_1973);
or U2085 (N_2085,N_2069,N_2039);
nor U2086 (N_2086,N_1950,N_2046);
xor U2087 (N_2087,N_2008,N_2076);
nor U2088 (N_2088,N_1972,N_2077);
nand U2089 (N_2089,N_2033,N_1995);
nand U2090 (N_2090,N_2067,N_1951);
xor U2091 (N_2091,N_1942,N_1921);
and U2092 (N_2092,N_1996,N_1974);
or U2093 (N_2093,N_2041,N_2032);
or U2094 (N_2094,N_1939,N_1932);
xnor U2095 (N_2095,N_2023,N_1936);
nand U2096 (N_2096,N_2026,N_1965);
or U2097 (N_2097,N_1933,N_1947);
and U2098 (N_2098,N_2015,N_1971);
and U2099 (N_2099,N_1945,N_1980);
xnor U2100 (N_2100,N_1935,N_1976);
or U2101 (N_2101,N_1987,N_2055);
nand U2102 (N_2102,N_1957,N_1963);
nor U2103 (N_2103,N_2056,N_2057);
and U2104 (N_2104,N_1954,N_2017);
nand U2105 (N_2105,N_2074,N_2024);
or U2106 (N_2106,N_2013,N_2079);
xnor U2107 (N_2107,N_1920,N_1927);
or U2108 (N_2108,N_1926,N_2001);
nor U2109 (N_2109,N_2061,N_1997);
and U2110 (N_2110,N_2044,N_2070);
or U2111 (N_2111,N_1966,N_2052);
nor U2112 (N_2112,N_1993,N_2027);
xor U2113 (N_2113,N_1981,N_2066);
nor U2114 (N_2114,N_2040,N_2016);
nand U2115 (N_2115,N_2078,N_1924);
or U2116 (N_2116,N_1994,N_1961);
nand U2117 (N_2117,N_2002,N_1977);
xor U2118 (N_2118,N_2006,N_1941);
and U2119 (N_2119,N_1985,N_1934);
xor U2120 (N_2120,N_1969,N_2007);
and U2121 (N_2121,N_1938,N_1937);
nor U2122 (N_2122,N_1922,N_1949);
and U2123 (N_2123,N_1988,N_2003);
or U2124 (N_2124,N_1955,N_2031);
xor U2125 (N_2125,N_2020,N_2029);
nand U2126 (N_2126,N_2049,N_1943);
nor U2127 (N_2127,N_1948,N_1970);
or U2128 (N_2128,N_2037,N_1992);
and U2129 (N_2129,N_1962,N_2064);
and U2130 (N_2130,N_2058,N_2050);
or U2131 (N_2131,N_2054,N_1952);
nor U2132 (N_2132,N_2048,N_2025);
nand U2133 (N_2133,N_1944,N_1925);
nand U2134 (N_2134,N_1967,N_2035);
or U2135 (N_2135,N_1960,N_1953);
nand U2136 (N_2136,N_1923,N_2021);
and U2137 (N_2137,N_2068,N_2019);
xnor U2138 (N_2138,N_1940,N_1978);
nor U2139 (N_2139,N_2030,N_1983);
nor U2140 (N_2140,N_1946,N_2009);
or U2141 (N_2141,N_2022,N_2043);
nor U2142 (N_2142,N_2073,N_2028);
nand U2143 (N_2143,N_2060,N_1956);
and U2144 (N_2144,N_2036,N_2072);
xor U2145 (N_2145,N_2010,N_1989);
xnor U2146 (N_2146,N_1986,N_2059);
nand U2147 (N_2147,N_1998,N_2005);
nand U2148 (N_2148,N_1930,N_1959);
xor U2149 (N_2149,N_1968,N_2063);
or U2150 (N_2150,N_2045,N_2075);
xor U2151 (N_2151,N_1979,N_2018);
nor U2152 (N_2152,N_2047,N_2000);
or U2153 (N_2153,N_2004,N_2012);
and U2154 (N_2154,N_1964,N_1984);
and U2155 (N_2155,N_1991,N_2062);
or U2156 (N_2156,N_1990,N_2053);
and U2157 (N_2157,N_2034,N_2071);
and U2158 (N_2158,N_1975,N_1958);
and U2159 (N_2159,N_2065,N_1929);
or U2160 (N_2160,N_2070,N_2034);
nor U2161 (N_2161,N_2014,N_2008);
nand U2162 (N_2162,N_1931,N_1992);
nand U2163 (N_2163,N_1947,N_2032);
and U2164 (N_2164,N_2047,N_2050);
nand U2165 (N_2165,N_2050,N_1923);
and U2166 (N_2166,N_2003,N_1957);
and U2167 (N_2167,N_2021,N_2038);
and U2168 (N_2168,N_1984,N_2047);
or U2169 (N_2169,N_2013,N_1956);
xor U2170 (N_2170,N_2028,N_2050);
nand U2171 (N_2171,N_1947,N_1984);
nor U2172 (N_2172,N_1923,N_1956);
or U2173 (N_2173,N_2020,N_1968);
nand U2174 (N_2174,N_2022,N_1928);
nand U2175 (N_2175,N_1931,N_1962);
and U2176 (N_2176,N_1939,N_1924);
nor U2177 (N_2177,N_2045,N_2020);
and U2178 (N_2178,N_1925,N_2021);
nor U2179 (N_2179,N_1996,N_1922);
nor U2180 (N_2180,N_2008,N_2073);
and U2181 (N_2181,N_1995,N_2024);
nor U2182 (N_2182,N_1971,N_1995);
or U2183 (N_2183,N_1995,N_2045);
nor U2184 (N_2184,N_1940,N_1959);
xor U2185 (N_2185,N_1934,N_1980);
xnor U2186 (N_2186,N_1932,N_1987);
nor U2187 (N_2187,N_2079,N_2059);
and U2188 (N_2188,N_1970,N_2013);
or U2189 (N_2189,N_2060,N_1949);
and U2190 (N_2190,N_2019,N_2026);
or U2191 (N_2191,N_1980,N_2037);
xnor U2192 (N_2192,N_1947,N_1945);
nor U2193 (N_2193,N_1975,N_2028);
or U2194 (N_2194,N_2020,N_1964);
xnor U2195 (N_2195,N_2070,N_1944);
or U2196 (N_2196,N_2077,N_2011);
nor U2197 (N_2197,N_2075,N_2042);
or U2198 (N_2198,N_2074,N_2018);
or U2199 (N_2199,N_1934,N_1999);
nand U2200 (N_2200,N_1941,N_2008);
nor U2201 (N_2201,N_2074,N_1940);
xor U2202 (N_2202,N_2021,N_1988);
nand U2203 (N_2203,N_2000,N_2017);
and U2204 (N_2204,N_1974,N_1975);
xnor U2205 (N_2205,N_2015,N_1921);
nor U2206 (N_2206,N_2017,N_2020);
and U2207 (N_2207,N_1934,N_2068);
xor U2208 (N_2208,N_2076,N_2035);
nand U2209 (N_2209,N_1968,N_1934);
and U2210 (N_2210,N_1950,N_1940);
or U2211 (N_2211,N_2042,N_1971);
nand U2212 (N_2212,N_1962,N_2053);
nor U2213 (N_2213,N_2010,N_1931);
nand U2214 (N_2214,N_2026,N_2046);
and U2215 (N_2215,N_2070,N_2064);
and U2216 (N_2216,N_1977,N_1926);
xor U2217 (N_2217,N_2021,N_1929);
nand U2218 (N_2218,N_1920,N_2067);
nand U2219 (N_2219,N_1956,N_2078);
xor U2220 (N_2220,N_1940,N_1981);
nand U2221 (N_2221,N_1940,N_2079);
nand U2222 (N_2222,N_1987,N_2067);
and U2223 (N_2223,N_2029,N_1974);
xor U2224 (N_2224,N_1961,N_1939);
xnor U2225 (N_2225,N_1943,N_2058);
nor U2226 (N_2226,N_2031,N_2057);
nand U2227 (N_2227,N_1958,N_2026);
and U2228 (N_2228,N_1998,N_2068);
or U2229 (N_2229,N_2028,N_2034);
xor U2230 (N_2230,N_2048,N_1928);
or U2231 (N_2231,N_2059,N_1960);
and U2232 (N_2232,N_1921,N_1987);
xor U2233 (N_2233,N_1972,N_1960);
nand U2234 (N_2234,N_2051,N_1964);
nand U2235 (N_2235,N_1959,N_2004);
and U2236 (N_2236,N_1935,N_1997);
nand U2237 (N_2237,N_2013,N_1966);
nor U2238 (N_2238,N_1945,N_1962);
and U2239 (N_2239,N_1993,N_1935);
or U2240 (N_2240,N_2088,N_2167);
and U2241 (N_2241,N_2164,N_2124);
or U2242 (N_2242,N_2138,N_2228);
or U2243 (N_2243,N_2161,N_2203);
nand U2244 (N_2244,N_2159,N_2239);
xor U2245 (N_2245,N_2162,N_2095);
or U2246 (N_2246,N_2105,N_2112);
and U2247 (N_2247,N_2233,N_2227);
xor U2248 (N_2248,N_2219,N_2107);
and U2249 (N_2249,N_2178,N_2204);
and U2250 (N_2250,N_2185,N_2237);
nand U2251 (N_2251,N_2222,N_2142);
xnor U2252 (N_2252,N_2089,N_2118);
nand U2253 (N_2253,N_2209,N_2192);
xor U2254 (N_2254,N_2195,N_2086);
xnor U2255 (N_2255,N_2188,N_2187);
xnor U2256 (N_2256,N_2200,N_2184);
or U2257 (N_2257,N_2189,N_2135);
or U2258 (N_2258,N_2151,N_2202);
or U2259 (N_2259,N_2104,N_2176);
nand U2260 (N_2260,N_2208,N_2119);
and U2261 (N_2261,N_2157,N_2173);
xnor U2262 (N_2262,N_2220,N_2133);
nor U2263 (N_2263,N_2103,N_2090);
and U2264 (N_2264,N_2102,N_2175);
or U2265 (N_2265,N_2206,N_2120);
nor U2266 (N_2266,N_2110,N_2224);
xnor U2267 (N_2267,N_2087,N_2180);
or U2268 (N_2268,N_2137,N_2143);
xor U2269 (N_2269,N_2109,N_2210);
and U2270 (N_2270,N_2199,N_2198);
xor U2271 (N_2271,N_2217,N_2232);
and U2272 (N_2272,N_2153,N_2136);
or U2273 (N_2273,N_2235,N_2230);
nand U2274 (N_2274,N_2094,N_2111);
nand U2275 (N_2275,N_2160,N_2080);
nor U2276 (N_2276,N_2129,N_2238);
nor U2277 (N_2277,N_2196,N_2211);
and U2278 (N_2278,N_2130,N_2144);
or U2279 (N_2279,N_2158,N_2213);
xor U2280 (N_2280,N_2174,N_2098);
xor U2281 (N_2281,N_2122,N_2081);
nand U2282 (N_2282,N_2131,N_2152);
or U2283 (N_2283,N_2236,N_2155);
nand U2284 (N_2284,N_2225,N_2085);
and U2285 (N_2285,N_2108,N_2127);
xnor U2286 (N_2286,N_2092,N_2150);
xor U2287 (N_2287,N_2207,N_2170);
and U2288 (N_2288,N_2212,N_2117);
nor U2289 (N_2289,N_2234,N_2083);
or U2290 (N_2290,N_2154,N_2183);
or U2291 (N_2291,N_2191,N_2139);
nor U2292 (N_2292,N_2226,N_2190);
nor U2293 (N_2293,N_2121,N_2216);
nor U2294 (N_2294,N_2201,N_2194);
nor U2295 (N_2295,N_2214,N_2197);
nor U2296 (N_2296,N_2113,N_2128);
and U2297 (N_2297,N_2163,N_2186);
xnor U2298 (N_2298,N_2114,N_2166);
xor U2299 (N_2299,N_2101,N_2097);
or U2300 (N_2300,N_2082,N_2165);
or U2301 (N_2301,N_2169,N_2096);
nand U2302 (N_2302,N_2149,N_2100);
nand U2303 (N_2303,N_2215,N_2125);
nor U2304 (N_2304,N_2181,N_2099);
xor U2305 (N_2305,N_2116,N_2221);
nand U2306 (N_2306,N_2141,N_2193);
nand U2307 (N_2307,N_2084,N_2156);
xnor U2308 (N_2308,N_2123,N_2179);
or U2309 (N_2309,N_2177,N_2145);
xor U2310 (N_2310,N_2132,N_2126);
or U2311 (N_2311,N_2168,N_2205);
nor U2312 (N_2312,N_2140,N_2182);
nor U2313 (N_2313,N_2229,N_2106);
or U2314 (N_2314,N_2148,N_2134);
nand U2315 (N_2315,N_2218,N_2231);
nor U2316 (N_2316,N_2093,N_2147);
xnor U2317 (N_2317,N_2223,N_2115);
xnor U2318 (N_2318,N_2171,N_2146);
and U2319 (N_2319,N_2172,N_2091);
and U2320 (N_2320,N_2233,N_2152);
and U2321 (N_2321,N_2129,N_2205);
nor U2322 (N_2322,N_2151,N_2148);
nand U2323 (N_2323,N_2235,N_2238);
nand U2324 (N_2324,N_2174,N_2138);
nand U2325 (N_2325,N_2229,N_2236);
nand U2326 (N_2326,N_2201,N_2092);
nand U2327 (N_2327,N_2151,N_2234);
nand U2328 (N_2328,N_2164,N_2106);
xnor U2329 (N_2329,N_2238,N_2143);
xor U2330 (N_2330,N_2223,N_2114);
or U2331 (N_2331,N_2142,N_2161);
xnor U2332 (N_2332,N_2102,N_2088);
nor U2333 (N_2333,N_2105,N_2224);
and U2334 (N_2334,N_2090,N_2164);
xnor U2335 (N_2335,N_2081,N_2204);
and U2336 (N_2336,N_2104,N_2168);
or U2337 (N_2337,N_2227,N_2148);
nor U2338 (N_2338,N_2085,N_2095);
xnor U2339 (N_2339,N_2120,N_2212);
and U2340 (N_2340,N_2119,N_2120);
nand U2341 (N_2341,N_2163,N_2081);
nor U2342 (N_2342,N_2186,N_2100);
xnor U2343 (N_2343,N_2183,N_2086);
nor U2344 (N_2344,N_2186,N_2185);
nor U2345 (N_2345,N_2094,N_2212);
xor U2346 (N_2346,N_2082,N_2101);
nand U2347 (N_2347,N_2129,N_2200);
nand U2348 (N_2348,N_2220,N_2101);
nand U2349 (N_2349,N_2212,N_2229);
xor U2350 (N_2350,N_2090,N_2162);
nor U2351 (N_2351,N_2110,N_2118);
nand U2352 (N_2352,N_2199,N_2109);
and U2353 (N_2353,N_2095,N_2092);
and U2354 (N_2354,N_2174,N_2108);
nand U2355 (N_2355,N_2173,N_2146);
and U2356 (N_2356,N_2128,N_2136);
or U2357 (N_2357,N_2225,N_2092);
or U2358 (N_2358,N_2237,N_2232);
or U2359 (N_2359,N_2214,N_2137);
or U2360 (N_2360,N_2080,N_2192);
xor U2361 (N_2361,N_2190,N_2131);
xnor U2362 (N_2362,N_2096,N_2218);
xor U2363 (N_2363,N_2095,N_2091);
nor U2364 (N_2364,N_2129,N_2236);
and U2365 (N_2365,N_2171,N_2127);
or U2366 (N_2366,N_2135,N_2232);
or U2367 (N_2367,N_2230,N_2108);
nand U2368 (N_2368,N_2211,N_2183);
or U2369 (N_2369,N_2223,N_2119);
and U2370 (N_2370,N_2116,N_2154);
nand U2371 (N_2371,N_2183,N_2164);
xor U2372 (N_2372,N_2170,N_2126);
or U2373 (N_2373,N_2098,N_2227);
and U2374 (N_2374,N_2141,N_2126);
nand U2375 (N_2375,N_2174,N_2225);
xor U2376 (N_2376,N_2229,N_2179);
and U2377 (N_2377,N_2201,N_2184);
nor U2378 (N_2378,N_2228,N_2238);
and U2379 (N_2379,N_2172,N_2130);
nand U2380 (N_2380,N_2133,N_2199);
xnor U2381 (N_2381,N_2138,N_2126);
nor U2382 (N_2382,N_2094,N_2188);
xnor U2383 (N_2383,N_2181,N_2234);
and U2384 (N_2384,N_2221,N_2121);
nand U2385 (N_2385,N_2229,N_2125);
xor U2386 (N_2386,N_2154,N_2200);
nand U2387 (N_2387,N_2197,N_2160);
or U2388 (N_2388,N_2125,N_2082);
nor U2389 (N_2389,N_2090,N_2086);
xnor U2390 (N_2390,N_2140,N_2230);
and U2391 (N_2391,N_2133,N_2232);
nand U2392 (N_2392,N_2238,N_2209);
and U2393 (N_2393,N_2196,N_2152);
and U2394 (N_2394,N_2200,N_2163);
xor U2395 (N_2395,N_2181,N_2210);
and U2396 (N_2396,N_2192,N_2197);
and U2397 (N_2397,N_2128,N_2167);
nand U2398 (N_2398,N_2099,N_2131);
xor U2399 (N_2399,N_2186,N_2237);
and U2400 (N_2400,N_2267,N_2344);
and U2401 (N_2401,N_2367,N_2342);
xor U2402 (N_2402,N_2280,N_2394);
and U2403 (N_2403,N_2347,N_2326);
nor U2404 (N_2404,N_2360,N_2269);
xnor U2405 (N_2405,N_2318,N_2365);
xor U2406 (N_2406,N_2366,N_2249);
and U2407 (N_2407,N_2262,N_2272);
xor U2408 (N_2408,N_2327,N_2387);
xor U2409 (N_2409,N_2264,N_2321);
nor U2410 (N_2410,N_2339,N_2313);
and U2411 (N_2411,N_2240,N_2244);
or U2412 (N_2412,N_2384,N_2337);
or U2413 (N_2413,N_2277,N_2390);
nand U2414 (N_2414,N_2274,N_2292);
or U2415 (N_2415,N_2260,N_2349);
nand U2416 (N_2416,N_2383,N_2317);
nand U2417 (N_2417,N_2351,N_2301);
or U2418 (N_2418,N_2379,N_2364);
nand U2419 (N_2419,N_2346,N_2281);
and U2420 (N_2420,N_2333,N_2319);
nand U2421 (N_2421,N_2376,N_2380);
nor U2422 (N_2422,N_2282,N_2389);
or U2423 (N_2423,N_2320,N_2359);
or U2424 (N_2424,N_2293,N_2328);
xor U2425 (N_2425,N_2361,N_2378);
nor U2426 (N_2426,N_2279,N_2370);
xnor U2427 (N_2427,N_2248,N_2373);
or U2428 (N_2428,N_2371,N_2278);
and U2429 (N_2429,N_2246,N_2354);
xor U2430 (N_2430,N_2398,N_2275);
or U2431 (N_2431,N_2307,N_2309);
xnor U2432 (N_2432,N_2287,N_2306);
and U2433 (N_2433,N_2391,N_2256);
or U2434 (N_2434,N_2255,N_2352);
or U2435 (N_2435,N_2334,N_2345);
or U2436 (N_2436,N_2312,N_2304);
xor U2437 (N_2437,N_2392,N_2263);
xnor U2438 (N_2438,N_2314,N_2310);
nor U2439 (N_2439,N_2395,N_2266);
and U2440 (N_2440,N_2386,N_2315);
and U2441 (N_2441,N_2316,N_2368);
xor U2442 (N_2442,N_2363,N_2348);
nor U2443 (N_2443,N_2323,N_2338);
or U2444 (N_2444,N_2289,N_2343);
nand U2445 (N_2445,N_2276,N_2286);
nand U2446 (N_2446,N_2299,N_2329);
or U2447 (N_2447,N_2388,N_2270);
and U2448 (N_2448,N_2268,N_2285);
xnor U2449 (N_2449,N_2302,N_2295);
xor U2450 (N_2450,N_2294,N_2261);
xor U2451 (N_2451,N_2340,N_2300);
and U2452 (N_2452,N_2357,N_2247);
or U2453 (N_2453,N_2265,N_2399);
and U2454 (N_2454,N_2396,N_2397);
and U2455 (N_2455,N_2374,N_2324);
or U2456 (N_2456,N_2377,N_2335);
xnor U2457 (N_2457,N_2273,N_2336);
nor U2458 (N_2458,N_2382,N_2353);
nor U2459 (N_2459,N_2251,N_2350);
and U2460 (N_2460,N_2356,N_2369);
nor U2461 (N_2461,N_2291,N_2245);
or U2462 (N_2462,N_2259,N_2393);
nor U2463 (N_2463,N_2372,N_2322);
or U2464 (N_2464,N_2331,N_2242);
xor U2465 (N_2465,N_2290,N_2298);
or U2466 (N_2466,N_2241,N_2305);
nor U2467 (N_2467,N_2381,N_2258);
or U2468 (N_2468,N_2283,N_2254);
nor U2469 (N_2469,N_2288,N_2311);
or U2470 (N_2470,N_2308,N_2252);
nor U2471 (N_2471,N_2257,N_2362);
nor U2472 (N_2472,N_2385,N_2250);
xnor U2473 (N_2473,N_2296,N_2243);
and U2474 (N_2474,N_2325,N_2271);
nand U2475 (N_2475,N_2375,N_2303);
nand U2476 (N_2476,N_2355,N_2284);
and U2477 (N_2477,N_2341,N_2330);
nor U2478 (N_2478,N_2297,N_2253);
nand U2479 (N_2479,N_2332,N_2358);
xor U2480 (N_2480,N_2369,N_2390);
xnor U2481 (N_2481,N_2323,N_2393);
nand U2482 (N_2482,N_2359,N_2276);
and U2483 (N_2483,N_2338,N_2283);
or U2484 (N_2484,N_2362,N_2259);
nor U2485 (N_2485,N_2253,N_2274);
xor U2486 (N_2486,N_2394,N_2253);
xnor U2487 (N_2487,N_2242,N_2284);
xor U2488 (N_2488,N_2321,N_2299);
or U2489 (N_2489,N_2315,N_2355);
and U2490 (N_2490,N_2392,N_2347);
and U2491 (N_2491,N_2260,N_2398);
or U2492 (N_2492,N_2240,N_2315);
or U2493 (N_2493,N_2297,N_2331);
xor U2494 (N_2494,N_2354,N_2271);
xor U2495 (N_2495,N_2354,N_2259);
nand U2496 (N_2496,N_2345,N_2264);
xor U2497 (N_2497,N_2322,N_2305);
nor U2498 (N_2498,N_2399,N_2252);
or U2499 (N_2499,N_2347,N_2385);
xor U2500 (N_2500,N_2345,N_2262);
nand U2501 (N_2501,N_2254,N_2320);
and U2502 (N_2502,N_2296,N_2386);
xor U2503 (N_2503,N_2325,N_2353);
nor U2504 (N_2504,N_2255,N_2344);
xor U2505 (N_2505,N_2251,N_2259);
or U2506 (N_2506,N_2337,N_2314);
and U2507 (N_2507,N_2319,N_2335);
or U2508 (N_2508,N_2383,N_2396);
nor U2509 (N_2509,N_2358,N_2250);
or U2510 (N_2510,N_2256,N_2367);
nand U2511 (N_2511,N_2288,N_2360);
xor U2512 (N_2512,N_2293,N_2318);
xnor U2513 (N_2513,N_2240,N_2267);
nor U2514 (N_2514,N_2320,N_2347);
xor U2515 (N_2515,N_2314,N_2306);
nand U2516 (N_2516,N_2313,N_2256);
or U2517 (N_2517,N_2270,N_2361);
nor U2518 (N_2518,N_2332,N_2371);
nor U2519 (N_2519,N_2304,N_2342);
and U2520 (N_2520,N_2356,N_2361);
or U2521 (N_2521,N_2249,N_2311);
nand U2522 (N_2522,N_2287,N_2309);
nor U2523 (N_2523,N_2308,N_2360);
or U2524 (N_2524,N_2244,N_2386);
nand U2525 (N_2525,N_2363,N_2295);
nor U2526 (N_2526,N_2270,N_2305);
xor U2527 (N_2527,N_2269,N_2340);
and U2528 (N_2528,N_2348,N_2352);
xor U2529 (N_2529,N_2251,N_2269);
and U2530 (N_2530,N_2388,N_2277);
or U2531 (N_2531,N_2371,N_2347);
and U2532 (N_2532,N_2352,N_2369);
nor U2533 (N_2533,N_2316,N_2264);
and U2534 (N_2534,N_2261,N_2292);
xnor U2535 (N_2535,N_2342,N_2242);
nand U2536 (N_2536,N_2240,N_2270);
xor U2537 (N_2537,N_2313,N_2336);
and U2538 (N_2538,N_2375,N_2359);
or U2539 (N_2539,N_2368,N_2331);
and U2540 (N_2540,N_2328,N_2324);
and U2541 (N_2541,N_2300,N_2336);
nor U2542 (N_2542,N_2358,N_2345);
or U2543 (N_2543,N_2301,N_2324);
and U2544 (N_2544,N_2368,N_2324);
nand U2545 (N_2545,N_2358,N_2252);
nor U2546 (N_2546,N_2262,N_2322);
and U2547 (N_2547,N_2319,N_2323);
nor U2548 (N_2548,N_2311,N_2354);
and U2549 (N_2549,N_2363,N_2284);
xnor U2550 (N_2550,N_2371,N_2399);
nand U2551 (N_2551,N_2371,N_2266);
nor U2552 (N_2552,N_2248,N_2348);
nor U2553 (N_2553,N_2249,N_2391);
and U2554 (N_2554,N_2267,N_2249);
or U2555 (N_2555,N_2385,N_2321);
xnor U2556 (N_2556,N_2328,N_2268);
or U2557 (N_2557,N_2242,N_2283);
or U2558 (N_2558,N_2375,N_2282);
nor U2559 (N_2559,N_2349,N_2387);
or U2560 (N_2560,N_2403,N_2559);
nand U2561 (N_2561,N_2424,N_2474);
nand U2562 (N_2562,N_2518,N_2452);
xor U2563 (N_2563,N_2539,N_2463);
and U2564 (N_2564,N_2470,N_2489);
xnor U2565 (N_2565,N_2483,N_2555);
nor U2566 (N_2566,N_2472,N_2544);
xor U2567 (N_2567,N_2462,N_2407);
or U2568 (N_2568,N_2511,N_2520);
or U2569 (N_2569,N_2538,N_2537);
xnor U2570 (N_2570,N_2449,N_2439);
nor U2571 (N_2571,N_2540,N_2557);
or U2572 (N_2572,N_2400,N_2482);
or U2573 (N_2573,N_2554,N_2534);
nand U2574 (N_2574,N_2519,N_2517);
and U2575 (N_2575,N_2434,N_2455);
nor U2576 (N_2576,N_2451,N_2546);
nor U2577 (N_2577,N_2499,N_2543);
xnor U2578 (N_2578,N_2440,N_2551);
and U2579 (N_2579,N_2530,N_2525);
nand U2580 (N_2580,N_2526,N_2421);
nand U2581 (N_2581,N_2453,N_2497);
nor U2582 (N_2582,N_2429,N_2535);
or U2583 (N_2583,N_2406,N_2408);
nand U2584 (N_2584,N_2418,N_2524);
or U2585 (N_2585,N_2523,N_2512);
and U2586 (N_2586,N_2416,N_2420);
nor U2587 (N_2587,N_2491,N_2481);
and U2588 (N_2588,N_2466,N_2488);
or U2589 (N_2589,N_2505,N_2558);
nor U2590 (N_2590,N_2446,N_2441);
or U2591 (N_2591,N_2405,N_2553);
xor U2592 (N_2592,N_2552,N_2486);
and U2593 (N_2593,N_2431,N_2454);
xnor U2594 (N_2594,N_2461,N_2509);
nand U2595 (N_2595,N_2542,N_2442);
and U2596 (N_2596,N_2469,N_2521);
and U2597 (N_2597,N_2471,N_2450);
nor U2598 (N_2598,N_2548,N_2508);
and U2599 (N_2599,N_2513,N_2432);
nor U2600 (N_2600,N_2550,N_2506);
or U2601 (N_2601,N_2504,N_2448);
and U2602 (N_2602,N_2468,N_2467);
nor U2603 (N_2603,N_2425,N_2479);
nor U2604 (N_2604,N_2484,N_2547);
nand U2605 (N_2605,N_2444,N_2430);
xnor U2606 (N_2606,N_2414,N_2541);
nand U2607 (N_2607,N_2495,N_2502);
xor U2608 (N_2608,N_2445,N_2447);
nand U2609 (N_2609,N_2428,N_2435);
nand U2610 (N_2610,N_2480,N_2487);
xor U2611 (N_2611,N_2423,N_2527);
or U2612 (N_2612,N_2503,N_2404);
nand U2613 (N_2613,N_2417,N_2473);
and U2614 (N_2614,N_2464,N_2556);
and U2615 (N_2615,N_2443,N_2401);
and U2616 (N_2616,N_2476,N_2426);
xnor U2617 (N_2617,N_2477,N_2536);
and U2618 (N_2618,N_2409,N_2419);
xnor U2619 (N_2619,N_2410,N_2516);
and U2620 (N_2620,N_2531,N_2510);
xor U2621 (N_2621,N_2427,N_2485);
or U2622 (N_2622,N_2545,N_2413);
or U2623 (N_2623,N_2515,N_2422);
or U2624 (N_2624,N_2465,N_2475);
or U2625 (N_2625,N_2460,N_2522);
or U2626 (N_2626,N_2501,N_2498);
xnor U2627 (N_2627,N_2549,N_2433);
nor U2628 (N_2628,N_2436,N_2507);
and U2629 (N_2629,N_2514,N_2402);
and U2630 (N_2630,N_2412,N_2458);
nor U2631 (N_2631,N_2437,N_2478);
nor U2632 (N_2632,N_2490,N_2500);
and U2633 (N_2633,N_2459,N_2528);
xnor U2634 (N_2634,N_2493,N_2496);
xor U2635 (N_2635,N_2415,N_2533);
and U2636 (N_2636,N_2456,N_2411);
nor U2637 (N_2637,N_2492,N_2438);
nor U2638 (N_2638,N_2529,N_2457);
xor U2639 (N_2639,N_2494,N_2532);
and U2640 (N_2640,N_2554,N_2522);
nor U2641 (N_2641,N_2485,N_2547);
and U2642 (N_2642,N_2483,N_2460);
or U2643 (N_2643,N_2406,N_2423);
or U2644 (N_2644,N_2488,N_2483);
xor U2645 (N_2645,N_2454,N_2408);
and U2646 (N_2646,N_2498,N_2411);
nor U2647 (N_2647,N_2402,N_2521);
nand U2648 (N_2648,N_2522,N_2410);
nor U2649 (N_2649,N_2507,N_2491);
or U2650 (N_2650,N_2477,N_2411);
or U2651 (N_2651,N_2534,N_2552);
nand U2652 (N_2652,N_2493,N_2506);
nand U2653 (N_2653,N_2526,N_2522);
and U2654 (N_2654,N_2426,N_2479);
xnor U2655 (N_2655,N_2503,N_2538);
nand U2656 (N_2656,N_2441,N_2519);
and U2657 (N_2657,N_2554,N_2486);
xor U2658 (N_2658,N_2505,N_2516);
or U2659 (N_2659,N_2418,N_2413);
or U2660 (N_2660,N_2505,N_2518);
nand U2661 (N_2661,N_2457,N_2430);
nor U2662 (N_2662,N_2423,N_2542);
xor U2663 (N_2663,N_2451,N_2449);
nor U2664 (N_2664,N_2480,N_2406);
and U2665 (N_2665,N_2505,N_2423);
or U2666 (N_2666,N_2447,N_2430);
and U2667 (N_2667,N_2509,N_2475);
nand U2668 (N_2668,N_2517,N_2460);
nor U2669 (N_2669,N_2446,N_2551);
and U2670 (N_2670,N_2459,N_2411);
or U2671 (N_2671,N_2439,N_2506);
xnor U2672 (N_2672,N_2467,N_2444);
nand U2673 (N_2673,N_2439,N_2464);
nor U2674 (N_2674,N_2416,N_2451);
xnor U2675 (N_2675,N_2473,N_2490);
xnor U2676 (N_2676,N_2514,N_2404);
nor U2677 (N_2677,N_2402,N_2537);
and U2678 (N_2678,N_2436,N_2490);
and U2679 (N_2679,N_2545,N_2511);
nand U2680 (N_2680,N_2549,N_2540);
nor U2681 (N_2681,N_2551,N_2422);
xor U2682 (N_2682,N_2552,N_2450);
and U2683 (N_2683,N_2440,N_2524);
xnor U2684 (N_2684,N_2513,N_2524);
and U2685 (N_2685,N_2436,N_2527);
nand U2686 (N_2686,N_2553,N_2459);
or U2687 (N_2687,N_2514,N_2537);
nand U2688 (N_2688,N_2500,N_2486);
nand U2689 (N_2689,N_2556,N_2419);
xor U2690 (N_2690,N_2494,N_2497);
nand U2691 (N_2691,N_2513,N_2530);
xnor U2692 (N_2692,N_2410,N_2528);
and U2693 (N_2693,N_2545,N_2453);
nor U2694 (N_2694,N_2486,N_2412);
and U2695 (N_2695,N_2416,N_2542);
nor U2696 (N_2696,N_2422,N_2477);
nor U2697 (N_2697,N_2438,N_2403);
or U2698 (N_2698,N_2461,N_2540);
and U2699 (N_2699,N_2482,N_2542);
nor U2700 (N_2700,N_2523,N_2450);
nor U2701 (N_2701,N_2553,N_2449);
xnor U2702 (N_2702,N_2551,N_2511);
nor U2703 (N_2703,N_2544,N_2447);
or U2704 (N_2704,N_2529,N_2486);
nand U2705 (N_2705,N_2520,N_2504);
nor U2706 (N_2706,N_2484,N_2407);
or U2707 (N_2707,N_2493,N_2467);
nand U2708 (N_2708,N_2519,N_2503);
xnor U2709 (N_2709,N_2436,N_2419);
nor U2710 (N_2710,N_2499,N_2483);
nor U2711 (N_2711,N_2481,N_2528);
or U2712 (N_2712,N_2541,N_2510);
and U2713 (N_2713,N_2467,N_2559);
or U2714 (N_2714,N_2496,N_2414);
and U2715 (N_2715,N_2478,N_2474);
xnor U2716 (N_2716,N_2543,N_2523);
nand U2717 (N_2717,N_2499,N_2501);
or U2718 (N_2718,N_2458,N_2479);
nand U2719 (N_2719,N_2519,N_2495);
xor U2720 (N_2720,N_2602,N_2611);
xnor U2721 (N_2721,N_2673,N_2567);
nand U2722 (N_2722,N_2682,N_2649);
xor U2723 (N_2723,N_2675,N_2654);
or U2724 (N_2724,N_2686,N_2570);
or U2725 (N_2725,N_2688,N_2580);
nand U2726 (N_2726,N_2685,N_2614);
and U2727 (N_2727,N_2565,N_2592);
and U2728 (N_2728,N_2698,N_2695);
and U2729 (N_2729,N_2705,N_2662);
or U2730 (N_2730,N_2615,N_2708);
nand U2731 (N_2731,N_2588,N_2669);
and U2732 (N_2732,N_2598,N_2563);
nand U2733 (N_2733,N_2648,N_2640);
xor U2734 (N_2734,N_2576,N_2634);
xnor U2735 (N_2735,N_2719,N_2633);
or U2736 (N_2736,N_2694,N_2653);
nor U2737 (N_2737,N_2652,N_2595);
or U2738 (N_2738,N_2693,N_2582);
or U2739 (N_2739,N_2572,N_2617);
xnor U2740 (N_2740,N_2667,N_2616);
nand U2741 (N_2741,N_2701,N_2679);
nand U2742 (N_2742,N_2594,N_2586);
xor U2743 (N_2743,N_2658,N_2626);
nor U2744 (N_2744,N_2700,N_2678);
nand U2745 (N_2745,N_2560,N_2601);
and U2746 (N_2746,N_2587,N_2624);
or U2747 (N_2747,N_2618,N_2574);
nor U2748 (N_2748,N_2564,N_2645);
xor U2749 (N_2749,N_2610,N_2646);
nand U2750 (N_2750,N_2597,N_2650);
or U2751 (N_2751,N_2627,N_2643);
nor U2752 (N_2752,N_2609,N_2684);
xor U2753 (N_2753,N_2629,N_2668);
xnor U2754 (N_2754,N_2680,N_2583);
nor U2755 (N_2755,N_2561,N_2607);
xor U2756 (N_2756,N_2579,N_2704);
nand U2757 (N_2757,N_2562,N_2659);
and U2758 (N_2758,N_2655,N_2712);
and U2759 (N_2759,N_2608,N_2620);
and U2760 (N_2760,N_2656,N_2638);
nor U2761 (N_2761,N_2585,N_2622);
xor U2762 (N_2762,N_2670,N_2687);
xor U2763 (N_2763,N_2591,N_2718);
and U2764 (N_2764,N_2664,N_2642);
and U2765 (N_2765,N_2710,N_2577);
nand U2766 (N_2766,N_2674,N_2630);
and U2767 (N_2767,N_2593,N_2636);
nand U2768 (N_2768,N_2621,N_2702);
xor U2769 (N_2769,N_2663,N_2717);
xor U2770 (N_2770,N_2683,N_2677);
nor U2771 (N_2771,N_2632,N_2709);
and U2772 (N_2772,N_2714,N_2651);
nand U2773 (N_2773,N_2566,N_2691);
or U2774 (N_2774,N_2665,N_2639);
xor U2775 (N_2775,N_2690,N_2573);
nor U2776 (N_2776,N_2713,N_2599);
nand U2777 (N_2777,N_2637,N_2671);
nor U2778 (N_2778,N_2703,N_2715);
xor U2779 (N_2779,N_2666,N_2625);
nor U2780 (N_2780,N_2681,N_2706);
nor U2781 (N_2781,N_2613,N_2605);
xnor U2782 (N_2782,N_2635,N_2612);
or U2783 (N_2783,N_2568,N_2676);
and U2784 (N_2784,N_2600,N_2606);
nor U2785 (N_2785,N_2692,N_2628);
and U2786 (N_2786,N_2569,N_2603);
and U2787 (N_2787,N_2672,N_2661);
nand U2788 (N_2788,N_2699,N_2641);
nor U2789 (N_2789,N_2689,N_2578);
or U2790 (N_2790,N_2707,N_2619);
or U2791 (N_2791,N_2631,N_2647);
nor U2792 (N_2792,N_2696,N_2711);
and U2793 (N_2793,N_2644,N_2596);
nor U2794 (N_2794,N_2581,N_2604);
xnor U2795 (N_2795,N_2697,N_2657);
or U2796 (N_2796,N_2571,N_2589);
or U2797 (N_2797,N_2716,N_2575);
nor U2798 (N_2798,N_2660,N_2590);
and U2799 (N_2799,N_2584,N_2623);
xor U2800 (N_2800,N_2635,N_2701);
nor U2801 (N_2801,N_2694,N_2699);
nor U2802 (N_2802,N_2584,N_2596);
nor U2803 (N_2803,N_2688,N_2572);
xnor U2804 (N_2804,N_2608,N_2640);
or U2805 (N_2805,N_2589,N_2663);
nor U2806 (N_2806,N_2628,N_2648);
and U2807 (N_2807,N_2691,N_2649);
xnor U2808 (N_2808,N_2579,N_2633);
xnor U2809 (N_2809,N_2590,N_2717);
nand U2810 (N_2810,N_2696,N_2588);
nand U2811 (N_2811,N_2710,N_2599);
nor U2812 (N_2812,N_2632,N_2673);
nand U2813 (N_2813,N_2582,N_2664);
nor U2814 (N_2814,N_2636,N_2586);
or U2815 (N_2815,N_2647,N_2645);
nor U2816 (N_2816,N_2596,N_2605);
nor U2817 (N_2817,N_2687,N_2653);
or U2818 (N_2818,N_2617,N_2638);
nand U2819 (N_2819,N_2580,N_2633);
and U2820 (N_2820,N_2688,N_2574);
or U2821 (N_2821,N_2610,N_2579);
xnor U2822 (N_2822,N_2690,N_2696);
nand U2823 (N_2823,N_2651,N_2653);
xor U2824 (N_2824,N_2704,N_2687);
and U2825 (N_2825,N_2644,N_2698);
nand U2826 (N_2826,N_2588,N_2674);
or U2827 (N_2827,N_2576,N_2572);
nand U2828 (N_2828,N_2577,N_2606);
xor U2829 (N_2829,N_2590,N_2595);
nor U2830 (N_2830,N_2613,N_2680);
nor U2831 (N_2831,N_2675,N_2561);
nand U2832 (N_2832,N_2675,N_2586);
and U2833 (N_2833,N_2661,N_2659);
nand U2834 (N_2834,N_2657,N_2589);
xnor U2835 (N_2835,N_2609,N_2570);
xor U2836 (N_2836,N_2719,N_2652);
nor U2837 (N_2837,N_2659,N_2605);
nor U2838 (N_2838,N_2585,N_2697);
nand U2839 (N_2839,N_2710,N_2680);
or U2840 (N_2840,N_2689,N_2628);
xnor U2841 (N_2841,N_2716,N_2579);
or U2842 (N_2842,N_2572,N_2669);
and U2843 (N_2843,N_2693,N_2650);
xor U2844 (N_2844,N_2704,N_2636);
nor U2845 (N_2845,N_2652,N_2676);
xor U2846 (N_2846,N_2672,N_2575);
and U2847 (N_2847,N_2578,N_2661);
xor U2848 (N_2848,N_2576,N_2671);
nor U2849 (N_2849,N_2593,N_2675);
nand U2850 (N_2850,N_2657,N_2614);
xor U2851 (N_2851,N_2665,N_2560);
nor U2852 (N_2852,N_2566,N_2649);
nand U2853 (N_2853,N_2603,N_2718);
nand U2854 (N_2854,N_2652,N_2582);
nor U2855 (N_2855,N_2582,N_2563);
or U2856 (N_2856,N_2647,N_2695);
and U2857 (N_2857,N_2569,N_2649);
nor U2858 (N_2858,N_2682,N_2650);
and U2859 (N_2859,N_2608,N_2652);
or U2860 (N_2860,N_2585,N_2657);
nor U2861 (N_2861,N_2653,N_2631);
and U2862 (N_2862,N_2609,N_2595);
nor U2863 (N_2863,N_2590,N_2587);
nand U2864 (N_2864,N_2644,N_2585);
xnor U2865 (N_2865,N_2614,N_2712);
nor U2866 (N_2866,N_2638,N_2640);
nand U2867 (N_2867,N_2689,N_2623);
or U2868 (N_2868,N_2590,N_2711);
xor U2869 (N_2869,N_2593,N_2652);
nand U2870 (N_2870,N_2671,N_2703);
or U2871 (N_2871,N_2676,N_2614);
nor U2872 (N_2872,N_2603,N_2571);
xor U2873 (N_2873,N_2633,N_2714);
xor U2874 (N_2874,N_2599,N_2637);
or U2875 (N_2875,N_2598,N_2699);
nor U2876 (N_2876,N_2590,N_2569);
nor U2877 (N_2877,N_2688,N_2655);
and U2878 (N_2878,N_2708,N_2642);
or U2879 (N_2879,N_2667,N_2640);
xor U2880 (N_2880,N_2835,N_2858);
nand U2881 (N_2881,N_2823,N_2739);
nand U2882 (N_2882,N_2820,N_2806);
and U2883 (N_2883,N_2736,N_2748);
xnor U2884 (N_2884,N_2734,N_2731);
or U2885 (N_2885,N_2879,N_2798);
nor U2886 (N_2886,N_2814,N_2792);
and U2887 (N_2887,N_2830,N_2872);
nor U2888 (N_2888,N_2747,N_2825);
nand U2889 (N_2889,N_2828,N_2876);
and U2890 (N_2890,N_2754,N_2757);
nor U2891 (N_2891,N_2766,N_2837);
nor U2892 (N_2892,N_2818,N_2730);
nand U2893 (N_2893,N_2850,N_2860);
nand U2894 (N_2894,N_2782,N_2811);
nand U2895 (N_2895,N_2765,N_2834);
and U2896 (N_2896,N_2870,N_2821);
or U2897 (N_2897,N_2787,N_2775);
nor U2898 (N_2898,N_2854,N_2848);
xnor U2899 (N_2899,N_2836,N_2774);
or U2900 (N_2900,N_2790,N_2722);
xor U2901 (N_2901,N_2857,N_2742);
xor U2902 (N_2902,N_2874,N_2789);
and U2903 (N_2903,N_2878,N_2786);
xor U2904 (N_2904,N_2824,N_2737);
nor U2905 (N_2905,N_2738,N_2759);
or U2906 (N_2906,N_2780,N_2802);
nor U2907 (N_2907,N_2760,N_2867);
xnor U2908 (N_2908,N_2800,N_2862);
or U2909 (N_2909,N_2749,N_2843);
xnor U2910 (N_2910,N_2752,N_2859);
nor U2911 (N_2911,N_2866,N_2793);
or U2912 (N_2912,N_2829,N_2788);
xnor U2913 (N_2913,N_2846,N_2772);
or U2914 (N_2914,N_2764,N_2784);
or U2915 (N_2915,N_2761,N_2855);
xnor U2916 (N_2916,N_2763,N_2847);
and U2917 (N_2917,N_2840,N_2804);
nor U2918 (N_2918,N_2724,N_2732);
xor U2919 (N_2919,N_2868,N_2838);
xor U2920 (N_2920,N_2781,N_2726);
nand U2921 (N_2921,N_2767,N_2805);
and U2922 (N_2922,N_2809,N_2841);
nand U2923 (N_2923,N_2791,N_2826);
and U2924 (N_2924,N_2743,N_2796);
and U2925 (N_2925,N_2770,N_2729);
nor U2926 (N_2926,N_2865,N_2777);
or U2927 (N_2927,N_2799,N_2771);
nand U2928 (N_2928,N_2773,N_2839);
nand U2929 (N_2929,N_2727,N_2861);
or U2930 (N_2930,N_2776,N_2723);
nor U2931 (N_2931,N_2801,N_2842);
xor U2932 (N_2932,N_2762,N_2813);
nand U2933 (N_2933,N_2873,N_2808);
and U2934 (N_2934,N_2733,N_2783);
xor U2935 (N_2935,N_2810,N_2785);
nand U2936 (N_2936,N_2853,N_2812);
nand U2937 (N_2937,N_2864,N_2856);
nor U2938 (N_2938,N_2750,N_2725);
or U2939 (N_2939,N_2833,N_2852);
nor U2940 (N_2940,N_2720,N_2721);
nand U2941 (N_2941,N_2849,N_2807);
xnor U2942 (N_2942,N_2755,N_2741);
nor U2943 (N_2943,N_2728,N_2877);
and U2944 (N_2944,N_2769,N_2803);
and U2945 (N_2945,N_2871,N_2822);
and U2946 (N_2946,N_2779,N_2740);
and U2947 (N_2947,N_2815,N_2863);
nand U2948 (N_2948,N_2735,N_2844);
nor U2949 (N_2949,N_2758,N_2845);
nand U2950 (N_2950,N_2744,N_2797);
or U2951 (N_2951,N_2816,N_2753);
and U2952 (N_2952,N_2756,N_2778);
nand U2953 (N_2953,N_2768,N_2751);
nand U2954 (N_2954,N_2795,N_2832);
nor U2955 (N_2955,N_2875,N_2745);
or U2956 (N_2956,N_2794,N_2817);
nor U2957 (N_2957,N_2746,N_2827);
xnor U2958 (N_2958,N_2869,N_2831);
or U2959 (N_2959,N_2851,N_2819);
or U2960 (N_2960,N_2725,N_2855);
or U2961 (N_2961,N_2786,N_2726);
and U2962 (N_2962,N_2814,N_2831);
and U2963 (N_2963,N_2856,N_2720);
and U2964 (N_2964,N_2877,N_2879);
nand U2965 (N_2965,N_2865,N_2878);
xnor U2966 (N_2966,N_2730,N_2878);
or U2967 (N_2967,N_2725,N_2732);
nor U2968 (N_2968,N_2835,N_2815);
and U2969 (N_2969,N_2808,N_2736);
xor U2970 (N_2970,N_2742,N_2808);
xor U2971 (N_2971,N_2741,N_2790);
and U2972 (N_2972,N_2840,N_2783);
or U2973 (N_2973,N_2854,N_2822);
or U2974 (N_2974,N_2879,N_2730);
and U2975 (N_2975,N_2774,N_2769);
or U2976 (N_2976,N_2783,N_2828);
xor U2977 (N_2977,N_2783,N_2750);
nor U2978 (N_2978,N_2864,N_2743);
or U2979 (N_2979,N_2839,N_2764);
nand U2980 (N_2980,N_2858,N_2761);
xor U2981 (N_2981,N_2766,N_2794);
nand U2982 (N_2982,N_2748,N_2767);
nand U2983 (N_2983,N_2848,N_2780);
or U2984 (N_2984,N_2732,N_2737);
or U2985 (N_2985,N_2720,N_2830);
nor U2986 (N_2986,N_2774,N_2766);
xor U2987 (N_2987,N_2839,N_2849);
and U2988 (N_2988,N_2810,N_2761);
and U2989 (N_2989,N_2728,N_2742);
or U2990 (N_2990,N_2767,N_2870);
or U2991 (N_2991,N_2764,N_2828);
nor U2992 (N_2992,N_2858,N_2748);
nand U2993 (N_2993,N_2767,N_2877);
nand U2994 (N_2994,N_2804,N_2831);
and U2995 (N_2995,N_2814,N_2723);
or U2996 (N_2996,N_2798,N_2853);
nand U2997 (N_2997,N_2792,N_2864);
nor U2998 (N_2998,N_2827,N_2724);
and U2999 (N_2999,N_2844,N_2825);
nor U3000 (N_3000,N_2750,N_2819);
nand U3001 (N_3001,N_2836,N_2847);
nand U3002 (N_3002,N_2756,N_2843);
xnor U3003 (N_3003,N_2760,N_2853);
xnor U3004 (N_3004,N_2766,N_2809);
nand U3005 (N_3005,N_2862,N_2857);
xnor U3006 (N_3006,N_2844,N_2780);
or U3007 (N_3007,N_2824,N_2791);
nand U3008 (N_3008,N_2724,N_2759);
and U3009 (N_3009,N_2742,N_2844);
or U3010 (N_3010,N_2864,N_2780);
nand U3011 (N_3011,N_2842,N_2868);
nand U3012 (N_3012,N_2857,N_2773);
and U3013 (N_3013,N_2749,N_2741);
xor U3014 (N_3014,N_2753,N_2720);
nand U3015 (N_3015,N_2867,N_2872);
nor U3016 (N_3016,N_2723,N_2754);
nor U3017 (N_3017,N_2818,N_2756);
xor U3018 (N_3018,N_2732,N_2797);
and U3019 (N_3019,N_2873,N_2806);
xnor U3020 (N_3020,N_2769,N_2757);
xnor U3021 (N_3021,N_2723,N_2793);
nand U3022 (N_3022,N_2815,N_2775);
and U3023 (N_3023,N_2772,N_2844);
or U3024 (N_3024,N_2876,N_2867);
and U3025 (N_3025,N_2733,N_2767);
nand U3026 (N_3026,N_2720,N_2724);
xnor U3027 (N_3027,N_2809,N_2811);
nand U3028 (N_3028,N_2773,N_2871);
or U3029 (N_3029,N_2792,N_2838);
nand U3030 (N_3030,N_2751,N_2766);
xor U3031 (N_3031,N_2853,N_2773);
nor U3032 (N_3032,N_2765,N_2729);
or U3033 (N_3033,N_2774,N_2832);
and U3034 (N_3034,N_2743,N_2769);
or U3035 (N_3035,N_2821,N_2753);
nand U3036 (N_3036,N_2820,N_2730);
and U3037 (N_3037,N_2872,N_2832);
and U3038 (N_3038,N_2829,N_2839);
or U3039 (N_3039,N_2801,N_2774);
and U3040 (N_3040,N_2916,N_2898);
and U3041 (N_3041,N_2880,N_2910);
and U3042 (N_3042,N_3037,N_2964);
nand U3043 (N_3043,N_3020,N_3032);
or U3044 (N_3044,N_3005,N_2935);
nand U3045 (N_3045,N_2933,N_2989);
and U3046 (N_3046,N_2953,N_2958);
nor U3047 (N_3047,N_2905,N_2939);
or U3048 (N_3048,N_2886,N_2940);
nor U3049 (N_3049,N_2899,N_2948);
xor U3050 (N_3050,N_2982,N_2894);
and U3051 (N_3051,N_2957,N_3023);
and U3052 (N_3052,N_2895,N_2904);
xor U3053 (N_3053,N_2972,N_2896);
xnor U3054 (N_3054,N_2975,N_2963);
or U3055 (N_3055,N_2938,N_2967);
nand U3056 (N_3056,N_2888,N_2913);
nor U3057 (N_3057,N_3036,N_2900);
or U3058 (N_3058,N_2928,N_2947);
nor U3059 (N_3059,N_2934,N_3001);
and U3060 (N_3060,N_2922,N_3019);
nor U3061 (N_3061,N_2981,N_2907);
xor U3062 (N_3062,N_2974,N_3003);
nand U3063 (N_3063,N_3004,N_2927);
nand U3064 (N_3064,N_2909,N_2911);
nor U3065 (N_3065,N_2931,N_2987);
and U3066 (N_3066,N_2986,N_2978);
nand U3067 (N_3067,N_3033,N_2889);
or U3068 (N_3068,N_2932,N_2906);
xor U3069 (N_3069,N_2956,N_2892);
and U3070 (N_3070,N_3035,N_2992);
and U3071 (N_3071,N_2965,N_2969);
nand U3072 (N_3072,N_2951,N_2885);
and U3073 (N_3073,N_2977,N_3031);
and U3074 (N_3074,N_2998,N_2897);
xor U3075 (N_3075,N_2995,N_2971);
and U3076 (N_3076,N_2961,N_2944);
and U3077 (N_3077,N_2884,N_3030);
nor U3078 (N_3078,N_2976,N_3021);
or U3079 (N_3079,N_2979,N_3029);
and U3080 (N_3080,N_2887,N_3013);
nor U3081 (N_3081,N_2960,N_2925);
nor U3082 (N_3082,N_3027,N_3006);
nand U3083 (N_3083,N_2924,N_2881);
nor U3084 (N_3084,N_2980,N_2917);
nor U3085 (N_3085,N_3022,N_2983);
and U3086 (N_3086,N_3009,N_3000);
nor U3087 (N_3087,N_2999,N_2942);
nand U3088 (N_3088,N_2901,N_2936);
and U3089 (N_3089,N_2993,N_2890);
nand U3090 (N_3090,N_2954,N_3002);
nand U3091 (N_3091,N_2930,N_2882);
nand U3092 (N_3092,N_2984,N_3039);
or U3093 (N_3093,N_2985,N_2908);
and U3094 (N_3094,N_2970,N_2893);
or U3095 (N_3095,N_3038,N_2973);
xor U3096 (N_3096,N_3007,N_2996);
and U3097 (N_3097,N_2988,N_2990);
or U3098 (N_3098,N_2968,N_2891);
and U3099 (N_3099,N_2952,N_2918);
nor U3100 (N_3100,N_2941,N_3015);
xor U3101 (N_3101,N_3026,N_2949);
or U3102 (N_3102,N_3025,N_2937);
nor U3103 (N_3103,N_2955,N_2943);
nand U3104 (N_3104,N_2914,N_2920);
xnor U3105 (N_3105,N_2997,N_3008);
and U3106 (N_3106,N_2921,N_3018);
or U3107 (N_3107,N_2912,N_2946);
and U3108 (N_3108,N_2902,N_2945);
nand U3109 (N_3109,N_2959,N_3010);
nand U3110 (N_3110,N_2991,N_2919);
and U3111 (N_3111,N_2903,N_2929);
nor U3112 (N_3112,N_3011,N_3014);
nand U3113 (N_3113,N_2915,N_2950);
nand U3114 (N_3114,N_3016,N_2926);
nand U3115 (N_3115,N_3028,N_3024);
and U3116 (N_3116,N_2883,N_2966);
nand U3117 (N_3117,N_2923,N_3034);
nand U3118 (N_3118,N_3017,N_3012);
and U3119 (N_3119,N_2962,N_2994);
xor U3120 (N_3120,N_2888,N_2898);
and U3121 (N_3121,N_2932,N_2952);
or U3122 (N_3122,N_2999,N_2989);
nor U3123 (N_3123,N_2994,N_2930);
xor U3124 (N_3124,N_2887,N_2898);
nor U3125 (N_3125,N_3016,N_2968);
xnor U3126 (N_3126,N_2890,N_2999);
nand U3127 (N_3127,N_2913,N_2886);
and U3128 (N_3128,N_2932,N_2908);
xnor U3129 (N_3129,N_2910,N_2890);
or U3130 (N_3130,N_2888,N_2963);
nor U3131 (N_3131,N_2930,N_2964);
and U3132 (N_3132,N_3015,N_2912);
xor U3133 (N_3133,N_2892,N_2960);
nor U3134 (N_3134,N_2937,N_2890);
or U3135 (N_3135,N_2893,N_2906);
nand U3136 (N_3136,N_2937,N_2934);
or U3137 (N_3137,N_2954,N_2955);
and U3138 (N_3138,N_3017,N_2936);
nor U3139 (N_3139,N_2983,N_2925);
and U3140 (N_3140,N_2908,N_2938);
nand U3141 (N_3141,N_2996,N_2983);
xnor U3142 (N_3142,N_2931,N_2988);
or U3143 (N_3143,N_2931,N_2890);
or U3144 (N_3144,N_2922,N_3016);
xnor U3145 (N_3145,N_2882,N_2914);
and U3146 (N_3146,N_3037,N_2901);
or U3147 (N_3147,N_2904,N_2896);
nand U3148 (N_3148,N_3038,N_2933);
nor U3149 (N_3149,N_2895,N_3010);
or U3150 (N_3150,N_2991,N_2911);
and U3151 (N_3151,N_2944,N_2979);
or U3152 (N_3152,N_2919,N_2895);
xnor U3153 (N_3153,N_3012,N_3034);
nor U3154 (N_3154,N_2901,N_2981);
and U3155 (N_3155,N_2985,N_2942);
and U3156 (N_3156,N_2895,N_2950);
xor U3157 (N_3157,N_2904,N_2917);
and U3158 (N_3158,N_2971,N_3001);
nor U3159 (N_3159,N_3015,N_2961);
xor U3160 (N_3160,N_3037,N_2945);
nand U3161 (N_3161,N_2890,N_2897);
and U3162 (N_3162,N_2888,N_2989);
nand U3163 (N_3163,N_2881,N_2972);
nand U3164 (N_3164,N_3033,N_2992);
nand U3165 (N_3165,N_2893,N_2901);
nor U3166 (N_3166,N_2969,N_2991);
nand U3167 (N_3167,N_2888,N_2933);
and U3168 (N_3168,N_2978,N_2934);
and U3169 (N_3169,N_2940,N_2932);
nand U3170 (N_3170,N_2882,N_2894);
nand U3171 (N_3171,N_2886,N_2963);
and U3172 (N_3172,N_2946,N_2997);
nor U3173 (N_3173,N_2995,N_3011);
xor U3174 (N_3174,N_3031,N_2983);
and U3175 (N_3175,N_3039,N_2891);
or U3176 (N_3176,N_2963,N_2924);
nand U3177 (N_3177,N_3013,N_2997);
and U3178 (N_3178,N_2981,N_3036);
nor U3179 (N_3179,N_3035,N_3036);
nand U3180 (N_3180,N_2991,N_3004);
nand U3181 (N_3181,N_2962,N_2946);
nand U3182 (N_3182,N_2985,N_3014);
or U3183 (N_3183,N_3011,N_3027);
xor U3184 (N_3184,N_3005,N_2897);
nand U3185 (N_3185,N_2951,N_2983);
and U3186 (N_3186,N_2910,N_2966);
nand U3187 (N_3187,N_2954,N_2953);
and U3188 (N_3188,N_3008,N_3035);
xnor U3189 (N_3189,N_2978,N_2977);
nor U3190 (N_3190,N_2911,N_2955);
and U3191 (N_3191,N_2964,N_2956);
or U3192 (N_3192,N_2982,N_2971);
nand U3193 (N_3193,N_2922,N_2950);
xnor U3194 (N_3194,N_2953,N_2881);
or U3195 (N_3195,N_3038,N_3030);
nand U3196 (N_3196,N_2943,N_3038);
or U3197 (N_3197,N_2959,N_3022);
and U3198 (N_3198,N_2946,N_2882);
xnor U3199 (N_3199,N_2962,N_2926);
nand U3200 (N_3200,N_3193,N_3122);
xor U3201 (N_3201,N_3171,N_3121);
nand U3202 (N_3202,N_3042,N_3199);
or U3203 (N_3203,N_3164,N_3183);
or U3204 (N_3204,N_3114,N_3085);
and U3205 (N_3205,N_3111,N_3173);
nor U3206 (N_3206,N_3151,N_3092);
nand U3207 (N_3207,N_3153,N_3103);
xnor U3208 (N_3208,N_3090,N_3132);
xor U3209 (N_3209,N_3155,N_3146);
nor U3210 (N_3210,N_3108,N_3054);
or U3211 (N_3211,N_3165,N_3185);
nor U3212 (N_3212,N_3118,N_3190);
xor U3213 (N_3213,N_3158,N_3142);
xor U3214 (N_3214,N_3074,N_3091);
nor U3215 (N_3215,N_3077,N_3167);
nand U3216 (N_3216,N_3128,N_3063);
nand U3217 (N_3217,N_3044,N_3130);
xor U3218 (N_3218,N_3041,N_3160);
or U3219 (N_3219,N_3046,N_3127);
nor U3220 (N_3220,N_3186,N_3178);
or U3221 (N_3221,N_3194,N_3116);
or U3222 (N_3222,N_3048,N_3043);
xnor U3223 (N_3223,N_3064,N_3180);
and U3224 (N_3224,N_3135,N_3052);
xnor U3225 (N_3225,N_3073,N_3101);
and U3226 (N_3226,N_3159,N_3176);
nor U3227 (N_3227,N_3120,N_3079);
nor U3228 (N_3228,N_3088,N_3154);
or U3229 (N_3229,N_3124,N_3181);
or U3230 (N_3230,N_3060,N_3191);
or U3231 (N_3231,N_3126,N_3096);
and U3232 (N_3232,N_3104,N_3058);
nand U3233 (N_3233,N_3156,N_3189);
or U3234 (N_3234,N_3197,N_3087);
xor U3235 (N_3235,N_3145,N_3075);
and U3236 (N_3236,N_3070,N_3061);
nand U3237 (N_3237,N_3182,N_3047);
or U3238 (N_3238,N_3097,N_3098);
nand U3239 (N_3239,N_3134,N_3068);
nand U3240 (N_3240,N_3175,N_3066);
and U3241 (N_3241,N_3188,N_3187);
nor U3242 (N_3242,N_3112,N_3131);
nand U3243 (N_3243,N_3071,N_3081);
nor U3244 (N_3244,N_3067,N_3080);
and U3245 (N_3245,N_3051,N_3196);
or U3246 (N_3246,N_3105,N_3065);
and U3247 (N_3247,N_3109,N_3177);
xnor U3248 (N_3248,N_3136,N_3141);
and U3249 (N_3249,N_3082,N_3094);
nor U3250 (N_3250,N_3195,N_3119);
xnor U3251 (N_3251,N_3040,N_3138);
nor U3252 (N_3252,N_3139,N_3133);
nand U3253 (N_3253,N_3099,N_3117);
nor U3254 (N_3254,N_3129,N_3140);
nand U3255 (N_3255,N_3095,N_3059);
or U3256 (N_3256,N_3144,N_3053);
nor U3257 (N_3257,N_3115,N_3056);
and U3258 (N_3258,N_3161,N_3149);
and U3259 (N_3259,N_3107,N_3069);
nand U3260 (N_3260,N_3078,N_3062);
nor U3261 (N_3261,N_3152,N_3106);
nand U3262 (N_3262,N_3093,N_3162);
or U3263 (N_3263,N_3086,N_3166);
and U3264 (N_3264,N_3125,N_3147);
nor U3265 (N_3265,N_3198,N_3137);
xnor U3266 (N_3266,N_3172,N_3057);
or U3267 (N_3267,N_3163,N_3174);
or U3268 (N_3268,N_3169,N_3168);
nor U3269 (N_3269,N_3076,N_3084);
nor U3270 (N_3270,N_3102,N_3055);
xor U3271 (N_3271,N_3192,N_3049);
xnor U3272 (N_3272,N_3184,N_3050);
or U3273 (N_3273,N_3110,N_3089);
nand U3274 (N_3274,N_3143,N_3072);
xor U3275 (N_3275,N_3083,N_3148);
xor U3276 (N_3276,N_3123,N_3113);
nor U3277 (N_3277,N_3170,N_3045);
nor U3278 (N_3278,N_3100,N_3150);
and U3279 (N_3279,N_3179,N_3157);
or U3280 (N_3280,N_3131,N_3094);
nand U3281 (N_3281,N_3177,N_3142);
and U3282 (N_3282,N_3157,N_3165);
and U3283 (N_3283,N_3142,N_3049);
and U3284 (N_3284,N_3198,N_3111);
and U3285 (N_3285,N_3086,N_3199);
or U3286 (N_3286,N_3170,N_3049);
xor U3287 (N_3287,N_3077,N_3047);
or U3288 (N_3288,N_3105,N_3162);
or U3289 (N_3289,N_3166,N_3116);
nand U3290 (N_3290,N_3096,N_3114);
nor U3291 (N_3291,N_3113,N_3170);
and U3292 (N_3292,N_3050,N_3055);
and U3293 (N_3293,N_3081,N_3087);
or U3294 (N_3294,N_3134,N_3194);
nand U3295 (N_3295,N_3132,N_3040);
and U3296 (N_3296,N_3075,N_3135);
or U3297 (N_3297,N_3195,N_3124);
or U3298 (N_3298,N_3133,N_3062);
or U3299 (N_3299,N_3118,N_3076);
nand U3300 (N_3300,N_3144,N_3158);
nand U3301 (N_3301,N_3132,N_3126);
or U3302 (N_3302,N_3170,N_3150);
nand U3303 (N_3303,N_3125,N_3150);
nand U3304 (N_3304,N_3142,N_3120);
and U3305 (N_3305,N_3045,N_3118);
or U3306 (N_3306,N_3164,N_3123);
nor U3307 (N_3307,N_3069,N_3155);
and U3308 (N_3308,N_3110,N_3171);
and U3309 (N_3309,N_3115,N_3068);
nor U3310 (N_3310,N_3068,N_3091);
nand U3311 (N_3311,N_3131,N_3121);
nand U3312 (N_3312,N_3088,N_3196);
and U3313 (N_3313,N_3047,N_3106);
and U3314 (N_3314,N_3196,N_3152);
and U3315 (N_3315,N_3153,N_3113);
or U3316 (N_3316,N_3063,N_3152);
or U3317 (N_3317,N_3170,N_3138);
or U3318 (N_3318,N_3044,N_3094);
nor U3319 (N_3319,N_3136,N_3109);
xor U3320 (N_3320,N_3157,N_3113);
nand U3321 (N_3321,N_3056,N_3073);
nand U3322 (N_3322,N_3193,N_3183);
xnor U3323 (N_3323,N_3075,N_3121);
xnor U3324 (N_3324,N_3089,N_3043);
xor U3325 (N_3325,N_3167,N_3163);
and U3326 (N_3326,N_3069,N_3186);
nor U3327 (N_3327,N_3045,N_3110);
xor U3328 (N_3328,N_3134,N_3159);
and U3329 (N_3329,N_3155,N_3179);
xor U3330 (N_3330,N_3145,N_3098);
xnor U3331 (N_3331,N_3195,N_3157);
and U3332 (N_3332,N_3150,N_3081);
nor U3333 (N_3333,N_3172,N_3091);
nor U3334 (N_3334,N_3048,N_3058);
and U3335 (N_3335,N_3052,N_3143);
xor U3336 (N_3336,N_3069,N_3065);
nand U3337 (N_3337,N_3194,N_3075);
and U3338 (N_3338,N_3167,N_3192);
nand U3339 (N_3339,N_3151,N_3156);
nor U3340 (N_3340,N_3152,N_3093);
or U3341 (N_3341,N_3048,N_3067);
xor U3342 (N_3342,N_3077,N_3123);
xnor U3343 (N_3343,N_3148,N_3114);
xor U3344 (N_3344,N_3174,N_3078);
and U3345 (N_3345,N_3083,N_3117);
and U3346 (N_3346,N_3062,N_3114);
xnor U3347 (N_3347,N_3122,N_3053);
nor U3348 (N_3348,N_3087,N_3098);
nor U3349 (N_3349,N_3153,N_3076);
nor U3350 (N_3350,N_3114,N_3118);
nand U3351 (N_3351,N_3196,N_3054);
xnor U3352 (N_3352,N_3152,N_3199);
nor U3353 (N_3353,N_3121,N_3172);
nor U3354 (N_3354,N_3142,N_3066);
and U3355 (N_3355,N_3060,N_3089);
and U3356 (N_3356,N_3189,N_3082);
nand U3357 (N_3357,N_3053,N_3064);
nor U3358 (N_3358,N_3151,N_3070);
nor U3359 (N_3359,N_3107,N_3045);
nor U3360 (N_3360,N_3274,N_3218);
and U3361 (N_3361,N_3284,N_3254);
nand U3362 (N_3362,N_3246,N_3241);
xnor U3363 (N_3363,N_3237,N_3203);
nand U3364 (N_3364,N_3344,N_3224);
and U3365 (N_3365,N_3209,N_3325);
and U3366 (N_3366,N_3334,N_3291);
xor U3367 (N_3367,N_3299,N_3302);
nor U3368 (N_3368,N_3264,N_3339);
or U3369 (N_3369,N_3326,N_3307);
or U3370 (N_3370,N_3309,N_3261);
and U3371 (N_3371,N_3270,N_3243);
xor U3372 (N_3372,N_3280,N_3257);
nor U3373 (N_3373,N_3358,N_3315);
xnor U3374 (N_3374,N_3319,N_3204);
xor U3375 (N_3375,N_3245,N_3226);
xor U3376 (N_3376,N_3217,N_3355);
or U3377 (N_3377,N_3260,N_3324);
and U3378 (N_3378,N_3342,N_3286);
nor U3379 (N_3379,N_3287,N_3275);
and U3380 (N_3380,N_3357,N_3253);
or U3381 (N_3381,N_3303,N_3350);
nor U3382 (N_3382,N_3231,N_3346);
and U3383 (N_3383,N_3262,N_3304);
xnor U3384 (N_3384,N_3297,N_3250);
nor U3385 (N_3385,N_3340,N_3244);
nand U3386 (N_3386,N_3320,N_3322);
nor U3387 (N_3387,N_3249,N_3239);
or U3388 (N_3388,N_3265,N_3290);
nand U3389 (N_3389,N_3356,N_3314);
nand U3390 (N_3390,N_3220,N_3232);
xor U3391 (N_3391,N_3258,N_3269);
or U3392 (N_3392,N_3301,N_3327);
and U3393 (N_3393,N_3343,N_3277);
nand U3394 (N_3394,N_3348,N_3312);
xnor U3395 (N_3395,N_3345,N_3352);
nor U3396 (N_3396,N_3271,N_3347);
xor U3397 (N_3397,N_3201,N_3323);
or U3398 (N_3398,N_3341,N_3294);
nand U3399 (N_3399,N_3272,N_3295);
or U3400 (N_3400,N_3211,N_3238);
xnor U3401 (N_3401,N_3332,N_3227);
and U3402 (N_3402,N_3279,N_3205);
nor U3403 (N_3403,N_3316,N_3317);
nor U3404 (N_3404,N_3285,N_3236);
nor U3405 (N_3405,N_3300,N_3359);
nor U3406 (N_3406,N_3255,N_3206);
nor U3407 (N_3407,N_3251,N_3252);
xnor U3408 (N_3408,N_3235,N_3208);
xnor U3409 (N_3409,N_3336,N_3228);
and U3410 (N_3410,N_3282,N_3328);
xor U3411 (N_3411,N_3331,N_3335);
nand U3412 (N_3412,N_3221,N_3278);
nor U3413 (N_3413,N_3321,N_3276);
nand U3414 (N_3414,N_3259,N_3306);
nand U3415 (N_3415,N_3215,N_3247);
xor U3416 (N_3416,N_3330,N_3256);
and U3417 (N_3417,N_3283,N_3213);
xnor U3418 (N_3418,N_3216,N_3289);
nor U3419 (N_3419,N_3308,N_3296);
and U3420 (N_3420,N_3222,N_3333);
nor U3421 (N_3421,N_3338,N_3329);
or U3422 (N_3422,N_3349,N_3305);
xor U3423 (N_3423,N_3292,N_3293);
nand U3424 (N_3424,N_3230,N_3353);
and U3425 (N_3425,N_3225,N_3219);
xor U3426 (N_3426,N_3229,N_3240);
and U3427 (N_3427,N_3311,N_3212);
and U3428 (N_3428,N_3200,N_3268);
nand U3429 (N_3429,N_3234,N_3288);
and U3430 (N_3430,N_3210,N_3298);
nor U3431 (N_3431,N_3310,N_3273);
nor U3432 (N_3432,N_3318,N_3207);
or U3433 (N_3433,N_3281,N_3266);
xnor U3434 (N_3434,N_3233,N_3267);
nor U3435 (N_3435,N_3242,N_3202);
nor U3436 (N_3436,N_3223,N_3354);
and U3437 (N_3437,N_3214,N_3337);
xor U3438 (N_3438,N_3351,N_3248);
nor U3439 (N_3439,N_3313,N_3263);
nor U3440 (N_3440,N_3219,N_3232);
nand U3441 (N_3441,N_3351,N_3225);
nand U3442 (N_3442,N_3227,N_3349);
nand U3443 (N_3443,N_3269,N_3291);
nand U3444 (N_3444,N_3282,N_3241);
nor U3445 (N_3445,N_3278,N_3242);
and U3446 (N_3446,N_3348,N_3359);
xnor U3447 (N_3447,N_3208,N_3332);
and U3448 (N_3448,N_3341,N_3232);
xnor U3449 (N_3449,N_3204,N_3258);
nand U3450 (N_3450,N_3222,N_3206);
xor U3451 (N_3451,N_3306,N_3208);
xor U3452 (N_3452,N_3203,N_3278);
xor U3453 (N_3453,N_3219,N_3218);
and U3454 (N_3454,N_3233,N_3323);
nand U3455 (N_3455,N_3245,N_3252);
xor U3456 (N_3456,N_3337,N_3319);
nand U3457 (N_3457,N_3293,N_3242);
or U3458 (N_3458,N_3225,N_3359);
or U3459 (N_3459,N_3302,N_3278);
xor U3460 (N_3460,N_3200,N_3326);
xnor U3461 (N_3461,N_3230,N_3224);
and U3462 (N_3462,N_3241,N_3249);
nor U3463 (N_3463,N_3230,N_3333);
and U3464 (N_3464,N_3214,N_3205);
xnor U3465 (N_3465,N_3302,N_3214);
nand U3466 (N_3466,N_3331,N_3318);
or U3467 (N_3467,N_3213,N_3299);
xnor U3468 (N_3468,N_3243,N_3226);
nand U3469 (N_3469,N_3260,N_3264);
nand U3470 (N_3470,N_3317,N_3249);
nand U3471 (N_3471,N_3289,N_3259);
nand U3472 (N_3472,N_3255,N_3272);
or U3473 (N_3473,N_3294,N_3285);
nand U3474 (N_3474,N_3287,N_3210);
nor U3475 (N_3475,N_3299,N_3228);
nor U3476 (N_3476,N_3271,N_3351);
and U3477 (N_3477,N_3239,N_3326);
nor U3478 (N_3478,N_3225,N_3226);
or U3479 (N_3479,N_3356,N_3359);
nand U3480 (N_3480,N_3271,N_3276);
or U3481 (N_3481,N_3290,N_3336);
nand U3482 (N_3482,N_3301,N_3276);
nor U3483 (N_3483,N_3271,N_3309);
nand U3484 (N_3484,N_3260,N_3331);
nor U3485 (N_3485,N_3202,N_3271);
nor U3486 (N_3486,N_3304,N_3353);
and U3487 (N_3487,N_3290,N_3251);
xnor U3488 (N_3488,N_3319,N_3354);
and U3489 (N_3489,N_3309,N_3203);
or U3490 (N_3490,N_3200,N_3222);
and U3491 (N_3491,N_3278,N_3206);
xnor U3492 (N_3492,N_3234,N_3317);
nand U3493 (N_3493,N_3232,N_3228);
or U3494 (N_3494,N_3239,N_3230);
xor U3495 (N_3495,N_3240,N_3210);
nor U3496 (N_3496,N_3282,N_3318);
and U3497 (N_3497,N_3306,N_3264);
and U3498 (N_3498,N_3215,N_3349);
xor U3499 (N_3499,N_3303,N_3211);
xnor U3500 (N_3500,N_3263,N_3353);
or U3501 (N_3501,N_3255,N_3249);
or U3502 (N_3502,N_3208,N_3287);
nor U3503 (N_3503,N_3266,N_3271);
or U3504 (N_3504,N_3245,N_3243);
nand U3505 (N_3505,N_3307,N_3227);
nand U3506 (N_3506,N_3205,N_3268);
nand U3507 (N_3507,N_3255,N_3298);
xnor U3508 (N_3508,N_3353,N_3288);
and U3509 (N_3509,N_3249,N_3252);
nor U3510 (N_3510,N_3259,N_3218);
nand U3511 (N_3511,N_3348,N_3307);
nand U3512 (N_3512,N_3286,N_3312);
and U3513 (N_3513,N_3294,N_3334);
and U3514 (N_3514,N_3207,N_3323);
nor U3515 (N_3515,N_3217,N_3319);
and U3516 (N_3516,N_3235,N_3334);
nor U3517 (N_3517,N_3280,N_3287);
nor U3518 (N_3518,N_3328,N_3344);
xor U3519 (N_3519,N_3351,N_3285);
nor U3520 (N_3520,N_3505,N_3496);
and U3521 (N_3521,N_3471,N_3454);
nor U3522 (N_3522,N_3400,N_3442);
nand U3523 (N_3523,N_3374,N_3409);
nand U3524 (N_3524,N_3497,N_3446);
or U3525 (N_3525,N_3369,N_3390);
xor U3526 (N_3526,N_3510,N_3416);
nand U3527 (N_3527,N_3451,N_3418);
or U3528 (N_3528,N_3372,N_3440);
or U3529 (N_3529,N_3377,N_3476);
and U3530 (N_3530,N_3421,N_3452);
nor U3531 (N_3531,N_3439,N_3443);
nand U3532 (N_3532,N_3507,N_3455);
nand U3533 (N_3533,N_3495,N_3463);
nor U3534 (N_3534,N_3519,N_3477);
nand U3535 (N_3535,N_3387,N_3444);
xor U3536 (N_3536,N_3436,N_3386);
and U3537 (N_3537,N_3489,N_3474);
and U3538 (N_3538,N_3504,N_3405);
nand U3539 (N_3539,N_3457,N_3514);
and U3540 (N_3540,N_3399,N_3373);
or U3541 (N_3541,N_3517,N_3368);
nand U3542 (N_3542,N_3434,N_3461);
and U3543 (N_3543,N_3376,N_3473);
and U3544 (N_3544,N_3388,N_3422);
or U3545 (N_3545,N_3509,N_3435);
nand U3546 (N_3546,N_3484,N_3415);
and U3547 (N_3547,N_3396,N_3441);
xnor U3548 (N_3548,N_3429,N_3459);
and U3549 (N_3549,N_3375,N_3449);
nor U3550 (N_3550,N_3410,N_3472);
nor U3551 (N_3551,N_3382,N_3408);
or U3552 (N_3552,N_3391,N_3456);
and U3553 (N_3553,N_3469,N_3478);
xnor U3554 (N_3554,N_3402,N_3448);
xor U3555 (N_3555,N_3498,N_3501);
and U3556 (N_3556,N_3508,N_3423);
or U3557 (N_3557,N_3503,N_3512);
xor U3558 (N_3558,N_3383,N_3481);
and U3559 (N_3559,N_3379,N_3371);
xnor U3560 (N_3560,N_3483,N_3370);
xor U3561 (N_3561,N_3419,N_3381);
or U3562 (N_3562,N_3482,N_3360);
or U3563 (N_3563,N_3404,N_3426);
and U3564 (N_3564,N_3516,N_3465);
or U3565 (N_3565,N_3367,N_3427);
and U3566 (N_3566,N_3458,N_3395);
xor U3567 (N_3567,N_3398,N_3500);
xnor U3568 (N_3568,N_3362,N_3513);
nor U3569 (N_3569,N_3361,N_3453);
nand U3570 (N_3570,N_3475,N_3406);
xnor U3571 (N_3571,N_3394,N_3397);
or U3572 (N_3572,N_3417,N_3403);
xor U3573 (N_3573,N_3420,N_3413);
and U3574 (N_3574,N_3438,N_3506);
xor U3575 (N_3575,N_3502,N_3380);
and U3576 (N_3576,N_3462,N_3437);
xnor U3577 (N_3577,N_3493,N_3384);
and U3578 (N_3578,N_3490,N_3450);
or U3579 (N_3579,N_3491,N_3431);
or U3580 (N_3580,N_3494,N_3414);
xnor U3581 (N_3581,N_3385,N_3433);
and U3582 (N_3582,N_3515,N_3468);
xnor U3583 (N_3583,N_3378,N_3460);
or U3584 (N_3584,N_3487,N_3428);
nor U3585 (N_3585,N_3393,N_3485);
xor U3586 (N_3586,N_3412,N_3464);
xor U3587 (N_3587,N_3407,N_3480);
and U3588 (N_3588,N_3364,N_3389);
nor U3589 (N_3589,N_3479,N_3432);
xnor U3590 (N_3590,N_3499,N_3518);
or U3591 (N_3591,N_3401,N_3366);
xor U3592 (N_3592,N_3511,N_3392);
and U3593 (N_3593,N_3365,N_3466);
nor U3594 (N_3594,N_3486,N_3425);
xor U3595 (N_3595,N_3467,N_3470);
nor U3596 (N_3596,N_3430,N_3447);
nor U3597 (N_3597,N_3363,N_3488);
nor U3598 (N_3598,N_3424,N_3411);
nor U3599 (N_3599,N_3492,N_3445);
or U3600 (N_3600,N_3502,N_3459);
or U3601 (N_3601,N_3400,N_3384);
nand U3602 (N_3602,N_3456,N_3444);
and U3603 (N_3603,N_3389,N_3519);
and U3604 (N_3604,N_3474,N_3519);
nor U3605 (N_3605,N_3516,N_3368);
nand U3606 (N_3606,N_3425,N_3436);
and U3607 (N_3607,N_3376,N_3364);
nor U3608 (N_3608,N_3517,N_3429);
nand U3609 (N_3609,N_3419,N_3472);
nor U3610 (N_3610,N_3506,N_3374);
or U3611 (N_3611,N_3469,N_3468);
nand U3612 (N_3612,N_3386,N_3425);
or U3613 (N_3613,N_3372,N_3450);
and U3614 (N_3614,N_3453,N_3401);
nand U3615 (N_3615,N_3491,N_3420);
or U3616 (N_3616,N_3504,N_3470);
nor U3617 (N_3617,N_3511,N_3385);
xnor U3618 (N_3618,N_3448,N_3409);
or U3619 (N_3619,N_3408,N_3510);
nand U3620 (N_3620,N_3423,N_3396);
and U3621 (N_3621,N_3364,N_3386);
nor U3622 (N_3622,N_3443,N_3457);
xor U3623 (N_3623,N_3381,N_3445);
xor U3624 (N_3624,N_3411,N_3377);
xnor U3625 (N_3625,N_3518,N_3506);
and U3626 (N_3626,N_3382,N_3463);
xor U3627 (N_3627,N_3494,N_3481);
or U3628 (N_3628,N_3401,N_3515);
nor U3629 (N_3629,N_3492,N_3382);
nand U3630 (N_3630,N_3424,N_3469);
and U3631 (N_3631,N_3462,N_3407);
nand U3632 (N_3632,N_3486,N_3493);
and U3633 (N_3633,N_3503,N_3422);
or U3634 (N_3634,N_3386,N_3389);
and U3635 (N_3635,N_3443,N_3514);
and U3636 (N_3636,N_3368,N_3407);
nor U3637 (N_3637,N_3379,N_3391);
or U3638 (N_3638,N_3378,N_3436);
or U3639 (N_3639,N_3453,N_3393);
and U3640 (N_3640,N_3440,N_3389);
nor U3641 (N_3641,N_3403,N_3449);
and U3642 (N_3642,N_3476,N_3431);
xnor U3643 (N_3643,N_3483,N_3445);
xnor U3644 (N_3644,N_3382,N_3511);
xor U3645 (N_3645,N_3474,N_3386);
nor U3646 (N_3646,N_3421,N_3453);
nor U3647 (N_3647,N_3393,N_3472);
and U3648 (N_3648,N_3367,N_3511);
and U3649 (N_3649,N_3400,N_3518);
nand U3650 (N_3650,N_3494,N_3371);
nor U3651 (N_3651,N_3382,N_3409);
nor U3652 (N_3652,N_3402,N_3391);
nand U3653 (N_3653,N_3510,N_3473);
xor U3654 (N_3654,N_3392,N_3426);
nand U3655 (N_3655,N_3486,N_3481);
or U3656 (N_3656,N_3366,N_3437);
nand U3657 (N_3657,N_3439,N_3391);
xnor U3658 (N_3658,N_3456,N_3505);
xnor U3659 (N_3659,N_3399,N_3503);
nand U3660 (N_3660,N_3413,N_3487);
or U3661 (N_3661,N_3408,N_3460);
or U3662 (N_3662,N_3495,N_3485);
and U3663 (N_3663,N_3450,N_3501);
xor U3664 (N_3664,N_3423,N_3472);
or U3665 (N_3665,N_3430,N_3455);
or U3666 (N_3666,N_3460,N_3389);
nand U3667 (N_3667,N_3404,N_3387);
xor U3668 (N_3668,N_3365,N_3426);
nand U3669 (N_3669,N_3453,N_3510);
and U3670 (N_3670,N_3384,N_3465);
xor U3671 (N_3671,N_3390,N_3361);
or U3672 (N_3672,N_3471,N_3503);
xor U3673 (N_3673,N_3489,N_3387);
nand U3674 (N_3674,N_3472,N_3507);
and U3675 (N_3675,N_3473,N_3472);
and U3676 (N_3676,N_3389,N_3498);
and U3677 (N_3677,N_3519,N_3379);
nand U3678 (N_3678,N_3516,N_3472);
or U3679 (N_3679,N_3437,N_3420);
or U3680 (N_3680,N_3629,N_3626);
nor U3681 (N_3681,N_3574,N_3651);
xor U3682 (N_3682,N_3543,N_3594);
nor U3683 (N_3683,N_3585,N_3531);
nand U3684 (N_3684,N_3654,N_3567);
or U3685 (N_3685,N_3613,N_3592);
and U3686 (N_3686,N_3527,N_3614);
xnor U3687 (N_3687,N_3587,N_3663);
xnor U3688 (N_3688,N_3617,N_3646);
xor U3689 (N_3689,N_3598,N_3642);
nor U3690 (N_3690,N_3677,N_3607);
xnor U3691 (N_3691,N_3673,N_3652);
nand U3692 (N_3692,N_3618,N_3657);
nand U3693 (N_3693,N_3612,N_3643);
xnor U3694 (N_3694,N_3628,N_3552);
or U3695 (N_3695,N_3635,N_3671);
xnor U3696 (N_3696,N_3610,N_3522);
xor U3697 (N_3697,N_3524,N_3597);
nand U3698 (N_3698,N_3529,N_3633);
or U3699 (N_3699,N_3542,N_3559);
or U3700 (N_3700,N_3655,N_3631);
or U3701 (N_3701,N_3666,N_3622);
and U3702 (N_3702,N_3554,N_3530);
or U3703 (N_3703,N_3596,N_3539);
and U3704 (N_3704,N_3624,N_3611);
xor U3705 (N_3705,N_3545,N_3541);
xnor U3706 (N_3706,N_3636,N_3647);
nand U3707 (N_3707,N_3606,N_3672);
nor U3708 (N_3708,N_3679,N_3645);
or U3709 (N_3709,N_3667,N_3579);
nand U3710 (N_3710,N_3548,N_3537);
xnor U3711 (N_3711,N_3555,N_3589);
and U3712 (N_3712,N_3550,N_3544);
xnor U3713 (N_3713,N_3678,N_3656);
and U3714 (N_3714,N_3572,N_3532);
nand U3715 (N_3715,N_3573,N_3595);
nor U3716 (N_3716,N_3650,N_3604);
nand U3717 (N_3717,N_3648,N_3533);
nand U3718 (N_3718,N_3615,N_3670);
nand U3719 (N_3719,N_3602,N_3546);
and U3720 (N_3720,N_3570,N_3520);
or U3721 (N_3721,N_3560,N_3561);
xor U3722 (N_3722,N_3575,N_3526);
nand U3723 (N_3723,N_3662,N_3659);
nor U3724 (N_3724,N_3534,N_3630);
and U3725 (N_3725,N_3535,N_3660);
nor U3726 (N_3726,N_3523,N_3649);
nand U3727 (N_3727,N_3599,N_3538);
or U3728 (N_3728,N_3584,N_3571);
nor U3729 (N_3729,N_3603,N_3582);
or U3730 (N_3730,N_3558,N_3521);
nor U3731 (N_3731,N_3556,N_3676);
and U3732 (N_3732,N_3664,N_3593);
nor U3733 (N_3733,N_3581,N_3632);
nor U3734 (N_3734,N_3641,N_3564);
or U3735 (N_3735,N_3621,N_3600);
or U3736 (N_3736,N_3590,N_3661);
xor U3737 (N_3737,N_3591,N_3568);
xor U3738 (N_3738,N_3565,N_3605);
nor U3739 (N_3739,N_3563,N_3578);
nand U3740 (N_3740,N_3525,N_3644);
nor U3741 (N_3741,N_3586,N_3576);
or U3742 (N_3742,N_3577,N_3583);
and U3743 (N_3743,N_3551,N_3580);
nor U3744 (N_3744,N_3623,N_3637);
nand U3745 (N_3745,N_3609,N_3665);
or U3746 (N_3746,N_3620,N_3569);
and U3747 (N_3747,N_3625,N_3634);
and U3748 (N_3748,N_3638,N_3549);
and U3749 (N_3749,N_3640,N_3608);
xor U3750 (N_3750,N_3627,N_3653);
or U3751 (N_3751,N_3601,N_3619);
xor U3752 (N_3752,N_3616,N_3553);
nand U3753 (N_3753,N_3540,N_3566);
xor U3754 (N_3754,N_3528,N_3658);
nor U3755 (N_3755,N_3669,N_3674);
nor U3756 (N_3756,N_3536,N_3639);
and U3757 (N_3757,N_3547,N_3588);
and U3758 (N_3758,N_3668,N_3557);
xor U3759 (N_3759,N_3675,N_3562);
nor U3760 (N_3760,N_3672,N_3528);
nor U3761 (N_3761,N_3673,N_3594);
xor U3762 (N_3762,N_3624,N_3564);
or U3763 (N_3763,N_3591,N_3659);
nand U3764 (N_3764,N_3645,N_3634);
or U3765 (N_3765,N_3675,N_3661);
or U3766 (N_3766,N_3531,N_3555);
and U3767 (N_3767,N_3666,N_3558);
nand U3768 (N_3768,N_3560,N_3613);
nor U3769 (N_3769,N_3543,N_3650);
or U3770 (N_3770,N_3635,N_3561);
nand U3771 (N_3771,N_3595,N_3654);
nand U3772 (N_3772,N_3576,N_3575);
and U3773 (N_3773,N_3586,N_3614);
nor U3774 (N_3774,N_3580,N_3525);
nor U3775 (N_3775,N_3583,N_3601);
nand U3776 (N_3776,N_3584,N_3627);
xnor U3777 (N_3777,N_3542,N_3586);
or U3778 (N_3778,N_3544,N_3607);
or U3779 (N_3779,N_3539,N_3670);
nand U3780 (N_3780,N_3586,N_3532);
nand U3781 (N_3781,N_3547,N_3596);
xnor U3782 (N_3782,N_3564,N_3639);
nand U3783 (N_3783,N_3562,N_3619);
xor U3784 (N_3784,N_3649,N_3653);
and U3785 (N_3785,N_3575,N_3548);
nand U3786 (N_3786,N_3652,N_3642);
nand U3787 (N_3787,N_3584,N_3576);
and U3788 (N_3788,N_3562,N_3527);
and U3789 (N_3789,N_3584,N_3645);
and U3790 (N_3790,N_3612,N_3550);
xnor U3791 (N_3791,N_3627,N_3529);
nor U3792 (N_3792,N_3679,N_3627);
and U3793 (N_3793,N_3627,N_3525);
nand U3794 (N_3794,N_3621,N_3520);
and U3795 (N_3795,N_3564,N_3648);
or U3796 (N_3796,N_3665,N_3558);
or U3797 (N_3797,N_3574,N_3674);
or U3798 (N_3798,N_3613,N_3627);
xor U3799 (N_3799,N_3661,N_3531);
and U3800 (N_3800,N_3522,N_3577);
xnor U3801 (N_3801,N_3628,N_3569);
or U3802 (N_3802,N_3587,N_3665);
or U3803 (N_3803,N_3619,N_3644);
and U3804 (N_3804,N_3609,N_3550);
xor U3805 (N_3805,N_3544,N_3577);
or U3806 (N_3806,N_3522,N_3638);
or U3807 (N_3807,N_3596,N_3553);
nand U3808 (N_3808,N_3635,N_3611);
and U3809 (N_3809,N_3642,N_3528);
nand U3810 (N_3810,N_3594,N_3622);
nor U3811 (N_3811,N_3583,N_3568);
nand U3812 (N_3812,N_3567,N_3673);
nor U3813 (N_3813,N_3675,N_3536);
or U3814 (N_3814,N_3610,N_3635);
xor U3815 (N_3815,N_3650,N_3593);
nand U3816 (N_3816,N_3534,N_3613);
or U3817 (N_3817,N_3549,N_3540);
nand U3818 (N_3818,N_3605,N_3560);
nand U3819 (N_3819,N_3599,N_3610);
and U3820 (N_3820,N_3619,N_3599);
nand U3821 (N_3821,N_3657,N_3645);
nor U3822 (N_3822,N_3638,N_3634);
and U3823 (N_3823,N_3586,N_3574);
or U3824 (N_3824,N_3547,N_3549);
nor U3825 (N_3825,N_3670,N_3620);
nand U3826 (N_3826,N_3609,N_3658);
nand U3827 (N_3827,N_3639,N_3671);
and U3828 (N_3828,N_3633,N_3552);
xnor U3829 (N_3829,N_3535,N_3537);
nor U3830 (N_3830,N_3621,N_3559);
xor U3831 (N_3831,N_3616,N_3617);
and U3832 (N_3832,N_3624,N_3546);
or U3833 (N_3833,N_3539,N_3662);
xnor U3834 (N_3834,N_3636,N_3549);
nor U3835 (N_3835,N_3541,N_3576);
or U3836 (N_3836,N_3524,N_3532);
and U3837 (N_3837,N_3593,N_3582);
and U3838 (N_3838,N_3520,N_3551);
nand U3839 (N_3839,N_3598,N_3525);
nand U3840 (N_3840,N_3781,N_3687);
or U3841 (N_3841,N_3772,N_3692);
nand U3842 (N_3842,N_3723,N_3708);
xnor U3843 (N_3843,N_3799,N_3763);
and U3844 (N_3844,N_3804,N_3783);
xnor U3845 (N_3845,N_3739,N_3764);
nand U3846 (N_3846,N_3757,N_3812);
xnor U3847 (N_3847,N_3777,N_3750);
or U3848 (N_3848,N_3742,N_3730);
xor U3849 (N_3849,N_3823,N_3817);
nor U3850 (N_3850,N_3788,N_3731);
nor U3851 (N_3851,N_3787,N_3743);
or U3852 (N_3852,N_3814,N_3695);
or U3853 (N_3853,N_3829,N_3683);
and U3854 (N_3854,N_3694,N_3724);
nor U3855 (N_3855,N_3688,N_3700);
or U3856 (N_3856,N_3719,N_3824);
or U3857 (N_3857,N_3831,N_3782);
nand U3858 (N_3858,N_3690,N_3749);
xnor U3859 (N_3859,N_3734,N_3778);
and U3860 (N_3860,N_3769,N_3789);
xnor U3861 (N_3861,N_3786,N_3755);
nor U3862 (N_3862,N_3818,N_3811);
and U3863 (N_3863,N_3810,N_3702);
nor U3864 (N_3864,N_3830,N_3681);
nor U3865 (N_3865,N_3802,N_3745);
and U3866 (N_3866,N_3725,N_3714);
nor U3867 (N_3867,N_3837,N_3751);
nand U3868 (N_3868,N_3835,N_3758);
xnor U3869 (N_3869,N_3754,N_3806);
or U3870 (N_3870,N_3697,N_3765);
or U3871 (N_3871,N_3791,N_3716);
or U3872 (N_3872,N_3834,N_3720);
and U3873 (N_3873,N_3691,N_3826);
xor U3874 (N_3874,N_3775,N_3798);
nor U3875 (N_3875,N_3762,N_3746);
xnor U3876 (N_3876,N_3760,N_3767);
xor U3877 (N_3877,N_3686,N_3693);
nand U3878 (N_3878,N_3827,N_3759);
nand U3879 (N_3879,N_3795,N_3771);
nand U3880 (N_3880,N_3822,N_3753);
xor U3881 (N_3881,N_3785,N_3705);
nand U3882 (N_3882,N_3717,N_3684);
nand U3883 (N_3883,N_3722,N_3709);
and U3884 (N_3884,N_3809,N_3706);
nor U3885 (N_3885,N_3729,N_3680);
nor U3886 (N_3886,N_3735,N_3728);
nand U3887 (N_3887,N_3793,N_3825);
and U3888 (N_3888,N_3805,N_3710);
nand U3889 (N_3889,N_3707,N_3713);
or U3890 (N_3890,N_3770,N_3721);
xnor U3891 (N_3891,N_3696,N_3801);
or U3892 (N_3892,N_3807,N_3813);
xor U3893 (N_3893,N_3780,N_3833);
or U3894 (N_3894,N_3816,N_3790);
or U3895 (N_3895,N_3838,N_3828);
nor U3896 (N_3896,N_3752,N_3726);
or U3897 (N_3897,N_3727,N_3685);
and U3898 (N_3898,N_3732,N_3711);
or U3899 (N_3899,N_3718,N_3794);
and U3900 (N_3900,N_3699,N_3747);
nand U3901 (N_3901,N_3748,N_3701);
nand U3902 (N_3902,N_3740,N_3766);
xor U3903 (N_3903,N_3839,N_3761);
or U3904 (N_3904,N_3689,N_3797);
nand U3905 (N_3905,N_3792,N_3776);
and U3906 (N_3906,N_3736,N_3808);
nand U3907 (N_3907,N_3820,N_3796);
nor U3908 (N_3908,N_3744,N_3768);
or U3909 (N_3909,N_3698,N_3779);
nand U3910 (N_3910,N_3800,N_3784);
nor U3911 (N_3911,N_3803,N_3819);
or U3912 (N_3912,N_3756,N_3774);
nor U3913 (N_3913,N_3704,N_3821);
nor U3914 (N_3914,N_3715,N_3737);
and U3915 (N_3915,N_3682,N_3836);
nand U3916 (N_3916,N_3832,N_3703);
xor U3917 (N_3917,N_3738,N_3733);
xnor U3918 (N_3918,N_3773,N_3815);
nor U3919 (N_3919,N_3712,N_3741);
xor U3920 (N_3920,N_3726,N_3742);
or U3921 (N_3921,N_3813,N_3714);
xnor U3922 (N_3922,N_3829,N_3701);
nor U3923 (N_3923,N_3806,N_3703);
or U3924 (N_3924,N_3686,N_3807);
nor U3925 (N_3925,N_3681,N_3702);
nand U3926 (N_3926,N_3754,N_3765);
or U3927 (N_3927,N_3770,N_3759);
nor U3928 (N_3928,N_3700,N_3709);
xnor U3929 (N_3929,N_3813,N_3684);
nor U3930 (N_3930,N_3738,N_3721);
xor U3931 (N_3931,N_3814,N_3724);
and U3932 (N_3932,N_3821,N_3820);
nand U3933 (N_3933,N_3683,N_3715);
and U3934 (N_3934,N_3696,N_3681);
xnor U3935 (N_3935,N_3746,N_3823);
nand U3936 (N_3936,N_3698,N_3695);
and U3937 (N_3937,N_3817,N_3809);
and U3938 (N_3938,N_3707,N_3800);
and U3939 (N_3939,N_3815,N_3812);
and U3940 (N_3940,N_3791,N_3758);
and U3941 (N_3941,N_3835,N_3739);
or U3942 (N_3942,N_3799,N_3794);
xor U3943 (N_3943,N_3702,N_3709);
and U3944 (N_3944,N_3800,N_3683);
xnor U3945 (N_3945,N_3770,N_3680);
nand U3946 (N_3946,N_3736,N_3689);
nor U3947 (N_3947,N_3817,N_3766);
nand U3948 (N_3948,N_3733,N_3820);
or U3949 (N_3949,N_3798,N_3711);
or U3950 (N_3950,N_3696,N_3831);
and U3951 (N_3951,N_3715,N_3734);
or U3952 (N_3952,N_3781,N_3838);
and U3953 (N_3953,N_3811,N_3826);
and U3954 (N_3954,N_3792,N_3760);
nand U3955 (N_3955,N_3768,N_3739);
and U3956 (N_3956,N_3786,N_3713);
or U3957 (N_3957,N_3694,N_3761);
and U3958 (N_3958,N_3793,N_3716);
or U3959 (N_3959,N_3743,N_3720);
nor U3960 (N_3960,N_3711,N_3754);
nor U3961 (N_3961,N_3723,N_3787);
nor U3962 (N_3962,N_3727,N_3705);
nand U3963 (N_3963,N_3814,N_3699);
and U3964 (N_3964,N_3743,N_3827);
xor U3965 (N_3965,N_3689,N_3743);
and U3966 (N_3966,N_3820,N_3772);
and U3967 (N_3967,N_3800,N_3786);
xor U3968 (N_3968,N_3682,N_3717);
and U3969 (N_3969,N_3708,N_3795);
nand U3970 (N_3970,N_3743,N_3680);
nand U3971 (N_3971,N_3813,N_3819);
nand U3972 (N_3972,N_3782,N_3837);
nor U3973 (N_3973,N_3685,N_3830);
nor U3974 (N_3974,N_3799,N_3766);
or U3975 (N_3975,N_3758,N_3767);
and U3976 (N_3976,N_3781,N_3763);
or U3977 (N_3977,N_3758,N_3733);
xnor U3978 (N_3978,N_3828,N_3708);
nor U3979 (N_3979,N_3683,N_3781);
or U3980 (N_3980,N_3743,N_3835);
or U3981 (N_3981,N_3795,N_3797);
nand U3982 (N_3982,N_3806,N_3752);
and U3983 (N_3983,N_3783,N_3684);
xor U3984 (N_3984,N_3692,N_3761);
xor U3985 (N_3985,N_3807,N_3701);
nor U3986 (N_3986,N_3788,N_3837);
or U3987 (N_3987,N_3799,N_3714);
xor U3988 (N_3988,N_3816,N_3807);
nand U3989 (N_3989,N_3811,N_3761);
or U3990 (N_3990,N_3754,N_3710);
nor U3991 (N_3991,N_3744,N_3793);
and U3992 (N_3992,N_3787,N_3806);
xor U3993 (N_3993,N_3727,N_3799);
or U3994 (N_3994,N_3718,N_3764);
xnor U3995 (N_3995,N_3691,N_3789);
nand U3996 (N_3996,N_3749,N_3827);
or U3997 (N_3997,N_3702,N_3746);
or U3998 (N_3998,N_3785,N_3763);
or U3999 (N_3999,N_3690,N_3772);
and U4000 (N_4000,N_3976,N_3989);
nand U4001 (N_4001,N_3974,N_3932);
nor U4002 (N_4002,N_3852,N_3985);
nor U4003 (N_4003,N_3999,N_3895);
and U4004 (N_4004,N_3862,N_3975);
and U4005 (N_4005,N_3906,N_3868);
nor U4006 (N_4006,N_3936,N_3948);
xnor U4007 (N_4007,N_3917,N_3848);
nor U4008 (N_4008,N_3981,N_3882);
or U4009 (N_4009,N_3877,N_3865);
or U4010 (N_4010,N_3899,N_3901);
nand U4011 (N_4011,N_3893,N_3897);
nor U4012 (N_4012,N_3855,N_3902);
or U4013 (N_4013,N_3968,N_3870);
nand U4014 (N_4014,N_3886,N_3973);
or U4015 (N_4015,N_3876,N_3997);
or U4016 (N_4016,N_3841,N_3950);
nand U4017 (N_4017,N_3982,N_3941);
xnor U4018 (N_4018,N_3866,N_3990);
and U4019 (N_4019,N_3892,N_3919);
nand U4020 (N_4020,N_3861,N_3924);
or U4021 (N_4021,N_3942,N_3935);
xor U4022 (N_4022,N_3938,N_3878);
xor U4023 (N_4023,N_3977,N_3995);
nand U4024 (N_4024,N_3916,N_3884);
xnor U4025 (N_4025,N_3954,N_3983);
nand U4026 (N_4026,N_3996,N_3898);
and U4027 (N_4027,N_3856,N_3854);
xor U4028 (N_4028,N_3900,N_3987);
nand U4029 (N_4029,N_3970,N_3962);
and U4030 (N_4030,N_3993,N_3859);
and U4031 (N_4031,N_3958,N_3921);
nand U4032 (N_4032,N_3915,N_3953);
and U4033 (N_4033,N_3943,N_3903);
nand U4034 (N_4034,N_3929,N_3879);
nor U4035 (N_4035,N_3951,N_3858);
or U4036 (N_4036,N_3928,N_3869);
or U4037 (N_4037,N_3907,N_3890);
nor U4038 (N_4038,N_3918,N_3991);
and U4039 (N_4039,N_3933,N_3966);
and U4040 (N_4040,N_3863,N_3988);
nor U4041 (N_4041,N_3912,N_3969);
and U4042 (N_4042,N_3875,N_3923);
and U4043 (N_4043,N_3940,N_3872);
nand U4044 (N_4044,N_3920,N_3843);
xnor U4045 (N_4045,N_3959,N_3930);
nor U4046 (N_4046,N_3994,N_3927);
nor U4047 (N_4047,N_3847,N_3937);
or U4048 (N_4048,N_3967,N_3910);
xnor U4049 (N_4049,N_3880,N_3961);
or U4050 (N_4050,N_3911,N_3842);
xnor U4051 (N_4051,N_3957,N_3925);
and U4052 (N_4052,N_3873,N_3984);
xnor U4053 (N_4053,N_3846,N_3955);
or U4054 (N_4054,N_3871,N_3964);
and U4055 (N_4055,N_3888,N_3844);
nand U4056 (N_4056,N_3887,N_3939);
xor U4057 (N_4057,N_3909,N_3881);
nand U4058 (N_4058,N_3891,N_3860);
nand U4059 (N_4059,N_3889,N_3931);
and U4060 (N_4060,N_3905,N_3867);
nand U4061 (N_4061,N_3978,N_3914);
nand U4062 (N_4062,N_3922,N_3949);
and U4063 (N_4063,N_3864,N_3908);
xnor U4064 (N_4064,N_3904,N_3883);
nand U4065 (N_4065,N_3979,N_3986);
or U4066 (N_4066,N_3971,N_3874);
or U4067 (N_4067,N_3851,N_3857);
nor U4068 (N_4068,N_3850,N_3972);
or U4069 (N_4069,N_3963,N_3960);
and U4070 (N_4070,N_3926,N_3913);
nand U4071 (N_4071,N_3956,N_3896);
nand U4072 (N_4072,N_3845,N_3965);
and U4073 (N_4073,N_3992,N_3947);
or U4074 (N_4074,N_3944,N_3980);
nand U4075 (N_4075,N_3952,N_3840);
and U4076 (N_4076,N_3945,N_3998);
nor U4077 (N_4077,N_3853,N_3894);
nand U4078 (N_4078,N_3934,N_3885);
nand U4079 (N_4079,N_3849,N_3946);
xor U4080 (N_4080,N_3969,N_3970);
xnor U4081 (N_4081,N_3847,N_3880);
nand U4082 (N_4082,N_3856,N_3845);
and U4083 (N_4083,N_3882,N_3871);
or U4084 (N_4084,N_3899,N_3936);
nand U4085 (N_4085,N_3988,N_3905);
and U4086 (N_4086,N_3902,N_3856);
nor U4087 (N_4087,N_3939,N_3873);
or U4088 (N_4088,N_3922,N_3850);
xnor U4089 (N_4089,N_3842,N_3991);
nand U4090 (N_4090,N_3972,N_3875);
or U4091 (N_4091,N_3924,N_3872);
nor U4092 (N_4092,N_3878,N_3974);
xor U4093 (N_4093,N_3976,N_3876);
and U4094 (N_4094,N_3860,N_3896);
nor U4095 (N_4095,N_3921,N_3929);
and U4096 (N_4096,N_3988,N_3997);
nor U4097 (N_4097,N_3926,N_3868);
nand U4098 (N_4098,N_3887,N_3957);
or U4099 (N_4099,N_3971,N_3924);
and U4100 (N_4100,N_3859,N_3880);
and U4101 (N_4101,N_3999,N_3994);
xnor U4102 (N_4102,N_3991,N_3902);
nand U4103 (N_4103,N_3922,N_3858);
or U4104 (N_4104,N_3931,N_3984);
nor U4105 (N_4105,N_3973,N_3905);
nand U4106 (N_4106,N_3951,N_3886);
or U4107 (N_4107,N_3977,N_3935);
nand U4108 (N_4108,N_3888,N_3855);
and U4109 (N_4109,N_3961,N_3990);
and U4110 (N_4110,N_3938,N_3963);
xnor U4111 (N_4111,N_3913,N_3901);
or U4112 (N_4112,N_3995,N_3855);
and U4113 (N_4113,N_3902,N_3984);
nor U4114 (N_4114,N_3904,N_3866);
and U4115 (N_4115,N_3943,N_3888);
or U4116 (N_4116,N_3864,N_3846);
nor U4117 (N_4117,N_3859,N_3969);
and U4118 (N_4118,N_3886,N_3987);
xnor U4119 (N_4119,N_3968,N_3965);
nand U4120 (N_4120,N_3890,N_3904);
xnor U4121 (N_4121,N_3930,N_3936);
nor U4122 (N_4122,N_3942,N_3913);
nand U4123 (N_4123,N_3843,N_3944);
nor U4124 (N_4124,N_3917,N_3921);
nand U4125 (N_4125,N_3910,N_3948);
or U4126 (N_4126,N_3840,N_3915);
xor U4127 (N_4127,N_3985,N_3993);
or U4128 (N_4128,N_3893,N_3967);
nand U4129 (N_4129,N_3867,N_3876);
nor U4130 (N_4130,N_3848,N_3892);
xor U4131 (N_4131,N_3846,N_3853);
xnor U4132 (N_4132,N_3912,N_3935);
and U4133 (N_4133,N_3878,N_3882);
and U4134 (N_4134,N_3957,N_3911);
and U4135 (N_4135,N_3963,N_3998);
or U4136 (N_4136,N_3852,N_3984);
nand U4137 (N_4137,N_3953,N_3875);
xnor U4138 (N_4138,N_3878,N_3987);
and U4139 (N_4139,N_3892,N_3844);
or U4140 (N_4140,N_3854,N_3859);
nor U4141 (N_4141,N_3933,N_3949);
xor U4142 (N_4142,N_3969,N_3968);
and U4143 (N_4143,N_3955,N_3967);
and U4144 (N_4144,N_3924,N_3922);
nand U4145 (N_4145,N_3942,N_3891);
and U4146 (N_4146,N_3948,N_3898);
and U4147 (N_4147,N_3844,N_3980);
nor U4148 (N_4148,N_3976,N_3903);
or U4149 (N_4149,N_3925,N_3967);
and U4150 (N_4150,N_3867,N_3980);
or U4151 (N_4151,N_3971,N_3897);
nor U4152 (N_4152,N_3882,N_3962);
and U4153 (N_4153,N_3849,N_3969);
xor U4154 (N_4154,N_3877,N_3860);
or U4155 (N_4155,N_3948,N_3974);
nor U4156 (N_4156,N_3928,N_3948);
xnor U4157 (N_4157,N_3960,N_3991);
or U4158 (N_4158,N_3929,N_3906);
xor U4159 (N_4159,N_3908,N_3871);
xnor U4160 (N_4160,N_4147,N_4029);
or U4161 (N_4161,N_4129,N_4090);
xor U4162 (N_4162,N_4036,N_4049);
nor U4163 (N_4163,N_4098,N_4118);
xnor U4164 (N_4164,N_4048,N_4103);
nand U4165 (N_4165,N_4088,N_4019);
nor U4166 (N_4166,N_4153,N_4051);
nor U4167 (N_4167,N_4137,N_4035);
nand U4168 (N_4168,N_4031,N_4007);
nand U4169 (N_4169,N_4058,N_4010);
xor U4170 (N_4170,N_4092,N_4075);
nand U4171 (N_4171,N_4000,N_4022);
nand U4172 (N_4172,N_4130,N_4099);
xnor U4173 (N_4173,N_4043,N_4121);
or U4174 (N_4174,N_4131,N_4003);
or U4175 (N_4175,N_4025,N_4152);
nor U4176 (N_4176,N_4158,N_4068);
nand U4177 (N_4177,N_4042,N_4021);
xor U4178 (N_4178,N_4083,N_4159);
xor U4179 (N_4179,N_4104,N_4034);
nand U4180 (N_4180,N_4116,N_4028);
nand U4181 (N_4181,N_4038,N_4120);
and U4182 (N_4182,N_4117,N_4061);
and U4183 (N_4183,N_4111,N_4125);
and U4184 (N_4184,N_4100,N_4027);
xor U4185 (N_4185,N_4157,N_4074);
nand U4186 (N_4186,N_4062,N_4143);
and U4187 (N_4187,N_4097,N_4144);
nand U4188 (N_4188,N_4089,N_4107);
nor U4189 (N_4189,N_4145,N_4046);
and U4190 (N_4190,N_4053,N_4087);
xnor U4191 (N_4191,N_4073,N_4095);
xor U4192 (N_4192,N_4023,N_4066);
nand U4193 (N_4193,N_4070,N_4064);
nor U4194 (N_4194,N_4085,N_4102);
nor U4195 (N_4195,N_4126,N_4093);
and U4196 (N_4196,N_4026,N_4105);
nor U4197 (N_4197,N_4050,N_4094);
or U4198 (N_4198,N_4012,N_4124);
and U4199 (N_4199,N_4109,N_4149);
and U4200 (N_4200,N_4054,N_4024);
nand U4201 (N_4201,N_4065,N_4141);
xor U4202 (N_4202,N_4148,N_4030);
and U4203 (N_4203,N_4057,N_4077);
xor U4204 (N_4204,N_4004,N_4071);
nor U4205 (N_4205,N_4142,N_4009);
or U4206 (N_4206,N_4108,N_4072);
nor U4207 (N_4207,N_4013,N_4115);
nor U4208 (N_4208,N_4146,N_4091);
and U4209 (N_4209,N_4018,N_4081);
and U4210 (N_4210,N_4123,N_4084);
xor U4211 (N_4211,N_4060,N_4156);
and U4212 (N_4212,N_4006,N_4134);
nand U4213 (N_4213,N_4080,N_4106);
and U4214 (N_4214,N_4079,N_4020);
nor U4215 (N_4215,N_4014,N_4059);
xor U4216 (N_4216,N_4154,N_4037);
nor U4217 (N_4217,N_4033,N_4016);
nand U4218 (N_4218,N_4128,N_4135);
or U4219 (N_4219,N_4151,N_4101);
or U4220 (N_4220,N_4155,N_4133);
nor U4221 (N_4221,N_4017,N_4076);
xor U4222 (N_4222,N_4140,N_4132);
xor U4223 (N_4223,N_4055,N_4001);
or U4224 (N_4224,N_4032,N_4096);
xnor U4225 (N_4225,N_4127,N_4011);
or U4226 (N_4226,N_4082,N_4015);
or U4227 (N_4227,N_4041,N_4150);
and U4228 (N_4228,N_4139,N_4069);
nand U4229 (N_4229,N_4119,N_4110);
and U4230 (N_4230,N_4114,N_4056);
or U4231 (N_4231,N_4047,N_4078);
nor U4232 (N_4232,N_4040,N_4044);
xor U4233 (N_4233,N_4112,N_4045);
nor U4234 (N_4234,N_4067,N_4052);
nand U4235 (N_4235,N_4039,N_4113);
xor U4236 (N_4236,N_4086,N_4138);
nor U4237 (N_4237,N_4008,N_4005);
xnor U4238 (N_4238,N_4002,N_4122);
nor U4239 (N_4239,N_4063,N_4136);
nor U4240 (N_4240,N_4055,N_4113);
and U4241 (N_4241,N_4066,N_4006);
or U4242 (N_4242,N_4117,N_4130);
xnor U4243 (N_4243,N_4019,N_4067);
xnor U4244 (N_4244,N_4005,N_4030);
nand U4245 (N_4245,N_4043,N_4100);
nand U4246 (N_4246,N_4097,N_4159);
xor U4247 (N_4247,N_4017,N_4075);
and U4248 (N_4248,N_4097,N_4001);
or U4249 (N_4249,N_4157,N_4080);
nand U4250 (N_4250,N_4098,N_4115);
xnor U4251 (N_4251,N_4099,N_4063);
nor U4252 (N_4252,N_4119,N_4129);
nand U4253 (N_4253,N_4067,N_4062);
and U4254 (N_4254,N_4088,N_4146);
and U4255 (N_4255,N_4043,N_4144);
xnor U4256 (N_4256,N_4029,N_4057);
nor U4257 (N_4257,N_4043,N_4155);
nor U4258 (N_4258,N_4061,N_4076);
nor U4259 (N_4259,N_4086,N_4028);
or U4260 (N_4260,N_4076,N_4025);
and U4261 (N_4261,N_4101,N_4074);
nand U4262 (N_4262,N_4145,N_4018);
xnor U4263 (N_4263,N_4004,N_4009);
nor U4264 (N_4264,N_4042,N_4105);
nand U4265 (N_4265,N_4079,N_4024);
nand U4266 (N_4266,N_4069,N_4066);
nor U4267 (N_4267,N_4075,N_4006);
and U4268 (N_4268,N_4046,N_4140);
nor U4269 (N_4269,N_4139,N_4003);
xor U4270 (N_4270,N_4105,N_4074);
xnor U4271 (N_4271,N_4063,N_4055);
nor U4272 (N_4272,N_4103,N_4060);
nor U4273 (N_4273,N_4146,N_4039);
nand U4274 (N_4274,N_4089,N_4154);
nand U4275 (N_4275,N_4063,N_4139);
and U4276 (N_4276,N_4117,N_4016);
nand U4277 (N_4277,N_4048,N_4127);
nor U4278 (N_4278,N_4018,N_4074);
or U4279 (N_4279,N_4079,N_4028);
nand U4280 (N_4280,N_4031,N_4098);
or U4281 (N_4281,N_4071,N_4028);
or U4282 (N_4282,N_4148,N_4081);
and U4283 (N_4283,N_4158,N_4029);
nor U4284 (N_4284,N_4158,N_4083);
or U4285 (N_4285,N_4012,N_4083);
or U4286 (N_4286,N_4059,N_4095);
and U4287 (N_4287,N_4083,N_4119);
nor U4288 (N_4288,N_4124,N_4126);
nor U4289 (N_4289,N_4098,N_4084);
or U4290 (N_4290,N_4094,N_4039);
or U4291 (N_4291,N_4013,N_4000);
nand U4292 (N_4292,N_4043,N_4046);
and U4293 (N_4293,N_4096,N_4142);
nor U4294 (N_4294,N_4056,N_4017);
or U4295 (N_4295,N_4069,N_4146);
nand U4296 (N_4296,N_4153,N_4062);
or U4297 (N_4297,N_4123,N_4144);
nor U4298 (N_4298,N_4096,N_4120);
nor U4299 (N_4299,N_4097,N_4156);
and U4300 (N_4300,N_4146,N_4122);
nand U4301 (N_4301,N_4007,N_4071);
xnor U4302 (N_4302,N_4049,N_4014);
nand U4303 (N_4303,N_4121,N_4064);
or U4304 (N_4304,N_4013,N_4044);
nand U4305 (N_4305,N_4101,N_4031);
nand U4306 (N_4306,N_4042,N_4114);
nor U4307 (N_4307,N_4099,N_4089);
xor U4308 (N_4308,N_4083,N_4142);
or U4309 (N_4309,N_4055,N_4126);
and U4310 (N_4310,N_4132,N_4096);
nand U4311 (N_4311,N_4051,N_4063);
or U4312 (N_4312,N_4107,N_4072);
and U4313 (N_4313,N_4036,N_4029);
xor U4314 (N_4314,N_4060,N_4144);
nand U4315 (N_4315,N_4151,N_4026);
or U4316 (N_4316,N_4104,N_4149);
and U4317 (N_4317,N_4125,N_4092);
xnor U4318 (N_4318,N_4093,N_4039);
and U4319 (N_4319,N_4007,N_4063);
nand U4320 (N_4320,N_4316,N_4246);
and U4321 (N_4321,N_4280,N_4228);
nor U4322 (N_4322,N_4162,N_4262);
or U4323 (N_4323,N_4239,N_4266);
and U4324 (N_4324,N_4309,N_4179);
nand U4325 (N_4325,N_4185,N_4221);
nor U4326 (N_4326,N_4304,N_4210);
nor U4327 (N_4327,N_4283,N_4197);
or U4328 (N_4328,N_4271,N_4289);
xor U4329 (N_4329,N_4302,N_4214);
nand U4330 (N_4330,N_4178,N_4171);
xor U4331 (N_4331,N_4298,N_4256);
nor U4332 (N_4332,N_4174,N_4232);
or U4333 (N_4333,N_4223,N_4258);
nand U4334 (N_4334,N_4255,N_4269);
nor U4335 (N_4335,N_4181,N_4166);
or U4336 (N_4336,N_4234,N_4248);
or U4337 (N_4337,N_4273,N_4199);
nand U4338 (N_4338,N_4237,N_4203);
nor U4339 (N_4339,N_4188,N_4284);
nand U4340 (N_4340,N_4296,N_4169);
nand U4341 (N_4341,N_4263,N_4279);
nand U4342 (N_4342,N_4305,N_4196);
nand U4343 (N_4343,N_4227,N_4236);
xnor U4344 (N_4344,N_4164,N_4213);
nor U4345 (N_4345,N_4191,N_4173);
or U4346 (N_4346,N_4319,N_4315);
xnor U4347 (N_4347,N_4267,N_4295);
xnor U4348 (N_4348,N_4290,N_4308);
nor U4349 (N_4349,N_4209,N_4270);
nor U4350 (N_4350,N_4165,N_4310);
or U4351 (N_4351,N_4194,N_4241);
xor U4352 (N_4352,N_4230,N_4233);
or U4353 (N_4353,N_4238,N_4161);
or U4354 (N_4354,N_4176,N_4276);
nand U4355 (N_4355,N_4317,N_4243);
and U4356 (N_4356,N_4278,N_4211);
or U4357 (N_4357,N_4291,N_4307);
and U4358 (N_4358,N_4252,N_4250);
and U4359 (N_4359,N_4167,N_4160);
and U4360 (N_4360,N_4272,N_4260);
xnor U4361 (N_4361,N_4311,N_4300);
nand U4362 (N_4362,N_4299,N_4207);
nand U4363 (N_4363,N_4265,N_4189);
xnor U4364 (N_4364,N_4240,N_4288);
nor U4365 (N_4365,N_4306,N_4303);
or U4366 (N_4366,N_4215,N_4195);
nand U4367 (N_4367,N_4200,N_4225);
xnor U4368 (N_4368,N_4163,N_4259);
nand U4369 (N_4369,N_4261,N_4190);
xnor U4370 (N_4370,N_4175,N_4168);
and U4371 (N_4371,N_4205,N_4257);
nor U4372 (N_4372,N_4193,N_4187);
or U4373 (N_4373,N_4206,N_4281);
and U4374 (N_4374,N_4253,N_4219);
xnor U4375 (N_4375,N_4216,N_4314);
nand U4376 (N_4376,N_4286,N_4274);
xnor U4377 (N_4377,N_4287,N_4229);
xnor U4378 (N_4378,N_4202,N_4268);
nor U4379 (N_4379,N_4170,N_4212);
or U4380 (N_4380,N_4282,N_4297);
or U4381 (N_4381,N_4172,N_4277);
nand U4382 (N_4382,N_4245,N_4275);
xor U4383 (N_4383,N_4226,N_4285);
nor U4384 (N_4384,N_4318,N_4201);
and U4385 (N_4385,N_4312,N_4254);
or U4386 (N_4386,N_4313,N_4192);
xor U4387 (N_4387,N_4184,N_4177);
and U4388 (N_4388,N_4208,N_4231);
nor U4389 (N_4389,N_4217,N_4244);
nand U4390 (N_4390,N_4224,N_4220);
nor U4391 (N_4391,N_4294,N_4292);
nor U4392 (N_4392,N_4293,N_4249);
xnor U4393 (N_4393,N_4264,N_4235);
nand U4394 (N_4394,N_4180,N_4251);
xor U4395 (N_4395,N_4218,N_4198);
nor U4396 (N_4396,N_4247,N_4222);
or U4397 (N_4397,N_4301,N_4182);
nor U4398 (N_4398,N_4204,N_4186);
and U4399 (N_4399,N_4242,N_4183);
or U4400 (N_4400,N_4236,N_4210);
and U4401 (N_4401,N_4313,N_4220);
and U4402 (N_4402,N_4279,N_4228);
xnor U4403 (N_4403,N_4239,N_4269);
or U4404 (N_4404,N_4306,N_4171);
xor U4405 (N_4405,N_4248,N_4191);
and U4406 (N_4406,N_4185,N_4303);
and U4407 (N_4407,N_4175,N_4237);
nand U4408 (N_4408,N_4276,N_4225);
nor U4409 (N_4409,N_4173,N_4293);
nor U4410 (N_4410,N_4245,N_4291);
or U4411 (N_4411,N_4294,N_4176);
nand U4412 (N_4412,N_4226,N_4273);
nor U4413 (N_4413,N_4166,N_4255);
nor U4414 (N_4414,N_4247,N_4195);
or U4415 (N_4415,N_4315,N_4230);
xor U4416 (N_4416,N_4201,N_4235);
and U4417 (N_4417,N_4241,N_4263);
and U4418 (N_4418,N_4287,N_4195);
or U4419 (N_4419,N_4265,N_4314);
nand U4420 (N_4420,N_4232,N_4227);
xor U4421 (N_4421,N_4314,N_4207);
nand U4422 (N_4422,N_4281,N_4312);
or U4423 (N_4423,N_4276,N_4278);
nor U4424 (N_4424,N_4211,N_4217);
nor U4425 (N_4425,N_4289,N_4262);
nor U4426 (N_4426,N_4174,N_4198);
and U4427 (N_4427,N_4167,N_4291);
nor U4428 (N_4428,N_4276,N_4214);
xor U4429 (N_4429,N_4247,N_4244);
or U4430 (N_4430,N_4226,N_4262);
or U4431 (N_4431,N_4229,N_4181);
or U4432 (N_4432,N_4260,N_4253);
nor U4433 (N_4433,N_4318,N_4160);
nand U4434 (N_4434,N_4259,N_4307);
or U4435 (N_4435,N_4282,N_4178);
nand U4436 (N_4436,N_4291,N_4264);
or U4437 (N_4437,N_4268,N_4266);
xor U4438 (N_4438,N_4312,N_4292);
nor U4439 (N_4439,N_4254,N_4229);
and U4440 (N_4440,N_4284,N_4165);
and U4441 (N_4441,N_4237,N_4254);
and U4442 (N_4442,N_4206,N_4212);
nor U4443 (N_4443,N_4181,N_4259);
nor U4444 (N_4444,N_4186,N_4232);
or U4445 (N_4445,N_4237,N_4311);
and U4446 (N_4446,N_4225,N_4273);
and U4447 (N_4447,N_4230,N_4277);
nand U4448 (N_4448,N_4221,N_4269);
nor U4449 (N_4449,N_4163,N_4309);
and U4450 (N_4450,N_4273,N_4231);
xor U4451 (N_4451,N_4265,N_4245);
or U4452 (N_4452,N_4174,N_4239);
or U4453 (N_4453,N_4296,N_4243);
and U4454 (N_4454,N_4178,N_4166);
nand U4455 (N_4455,N_4285,N_4263);
or U4456 (N_4456,N_4296,N_4278);
nand U4457 (N_4457,N_4295,N_4186);
and U4458 (N_4458,N_4219,N_4301);
xnor U4459 (N_4459,N_4295,N_4247);
and U4460 (N_4460,N_4193,N_4260);
xor U4461 (N_4461,N_4247,N_4245);
nor U4462 (N_4462,N_4255,N_4282);
xor U4463 (N_4463,N_4235,N_4215);
nor U4464 (N_4464,N_4239,N_4201);
xor U4465 (N_4465,N_4200,N_4172);
and U4466 (N_4466,N_4250,N_4219);
xor U4467 (N_4467,N_4200,N_4220);
and U4468 (N_4468,N_4238,N_4226);
nand U4469 (N_4469,N_4241,N_4223);
xor U4470 (N_4470,N_4172,N_4209);
or U4471 (N_4471,N_4266,N_4290);
nand U4472 (N_4472,N_4289,N_4227);
and U4473 (N_4473,N_4220,N_4318);
nor U4474 (N_4474,N_4223,N_4212);
xor U4475 (N_4475,N_4233,N_4272);
nand U4476 (N_4476,N_4307,N_4317);
or U4477 (N_4477,N_4312,N_4214);
and U4478 (N_4478,N_4242,N_4174);
xnor U4479 (N_4479,N_4213,N_4174);
nand U4480 (N_4480,N_4376,N_4352);
xnor U4481 (N_4481,N_4477,N_4393);
nand U4482 (N_4482,N_4429,N_4459);
nand U4483 (N_4483,N_4435,N_4367);
nor U4484 (N_4484,N_4433,N_4354);
or U4485 (N_4485,N_4457,N_4344);
or U4486 (N_4486,N_4335,N_4343);
xnor U4487 (N_4487,N_4424,N_4360);
xor U4488 (N_4488,N_4448,N_4405);
nor U4489 (N_4489,N_4413,N_4466);
xor U4490 (N_4490,N_4361,N_4420);
nand U4491 (N_4491,N_4451,N_4323);
and U4492 (N_4492,N_4342,N_4359);
nand U4493 (N_4493,N_4390,N_4437);
nor U4494 (N_4494,N_4467,N_4465);
and U4495 (N_4495,N_4442,N_4398);
or U4496 (N_4496,N_4409,N_4368);
or U4497 (N_4497,N_4415,N_4410);
or U4498 (N_4498,N_4421,N_4454);
and U4499 (N_4499,N_4345,N_4356);
xnor U4500 (N_4500,N_4436,N_4463);
nor U4501 (N_4501,N_4375,N_4461);
or U4502 (N_4502,N_4419,N_4432);
xnor U4503 (N_4503,N_4453,N_4380);
xor U4504 (N_4504,N_4418,N_4423);
and U4505 (N_4505,N_4358,N_4408);
nor U4506 (N_4506,N_4383,N_4384);
xnor U4507 (N_4507,N_4329,N_4417);
and U4508 (N_4508,N_4425,N_4353);
nor U4509 (N_4509,N_4450,N_4386);
or U4510 (N_4510,N_4445,N_4388);
nand U4511 (N_4511,N_4462,N_4362);
xnor U4512 (N_4512,N_4325,N_4411);
or U4513 (N_4513,N_4395,N_4391);
and U4514 (N_4514,N_4439,N_4476);
nand U4515 (N_4515,N_4458,N_4469);
xor U4516 (N_4516,N_4399,N_4455);
and U4517 (N_4517,N_4334,N_4414);
xnor U4518 (N_4518,N_4404,N_4427);
nor U4519 (N_4519,N_4392,N_4441);
nor U4520 (N_4520,N_4444,N_4397);
nor U4521 (N_4521,N_4389,N_4479);
nand U4522 (N_4522,N_4348,N_4412);
or U4523 (N_4523,N_4456,N_4327);
nor U4524 (N_4524,N_4403,N_4370);
or U4525 (N_4525,N_4470,N_4336);
nor U4526 (N_4526,N_4449,N_4401);
and U4527 (N_4527,N_4446,N_4333);
xnor U4528 (N_4528,N_4350,N_4330);
nor U4529 (N_4529,N_4394,N_4357);
and U4530 (N_4530,N_4474,N_4349);
and U4531 (N_4531,N_4452,N_4468);
xnor U4532 (N_4532,N_4472,N_4363);
nor U4533 (N_4533,N_4346,N_4426);
xnor U4534 (N_4534,N_4416,N_4400);
and U4535 (N_4535,N_4374,N_4460);
nor U4536 (N_4536,N_4378,N_4428);
or U4537 (N_4537,N_4321,N_4369);
xnor U4538 (N_4538,N_4338,N_4475);
or U4539 (N_4539,N_4351,N_4396);
or U4540 (N_4540,N_4324,N_4443);
nor U4541 (N_4541,N_4402,N_4337);
and U4542 (N_4542,N_4366,N_4434);
or U4543 (N_4543,N_4377,N_4431);
xnor U4544 (N_4544,N_4332,N_4372);
xor U4545 (N_4545,N_4373,N_4341);
xnor U4546 (N_4546,N_4447,N_4331);
nor U4547 (N_4547,N_4322,N_4407);
xnor U4548 (N_4548,N_4365,N_4355);
nor U4549 (N_4549,N_4320,N_4381);
xnor U4550 (N_4550,N_4364,N_4430);
xor U4551 (N_4551,N_4326,N_4464);
or U4552 (N_4552,N_4385,N_4328);
or U4553 (N_4553,N_4478,N_4471);
and U4554 (N_4554,N_4340,N_4387);
xor U4555 (N_4555,N_4371,N_4339);
nor U4556 (N_4556,N_4440,N_4379);
nor U4557 (N_4557,N_4347,N_4382);
nand U4558 (N_4558,N_4473,N_4438);
and U4559 (N_4559,N_4406,N_4422);
xnor U4560 (N_4560,N_4337,N_4327);
and U4561 (N_4561,N_4435,N_4354);
nor U4562 (N_4562,N_4452,N_4456);
and U4563 (N_4563,N_4416,N_4445);
nand U4564 (N_4564,N_4369,N_4341);
and U4565 (N_4565,N_4386,N_4381);
or U4566 (N_4566,N_4403,N_4335);
or U4567 (N_4567,N_4449,N_4467);
nand U4568 (N_4568,N_4445,N_4434);
and U4569 (N_4569,N_4435,N_4454);
or U4570 (N_4570,N_4338,N_4347);
nor U4571 (N_4571,N_4352,N_4347);
nand U4572 (N_4572,N_4478,N_4404);
nor U4573 (N_4573,N_4441,N_4323);
or U4574 (N_4574,N_4413,N_4322);
nand U4575 (N_4575,N_4341,N_4447);
nand U4576 (N_4576,N_4324,N_4338);
nor U4577 (N_4577,N_4391,N_4452);
or U4578 (N_4578,N_4475,N_4413);
nand U4579 (N_4579,N_4320,N_4406);
or U4580 (N_4580,N_4360,N_4478);
or U4581 (N_4581,N_4354,N_4377);
and U4582 (N_4582,N_4327,N_4412);
nand U4583 (N_4583,N_4442,N_4344);
nand U4584 (N_4584,N_4424,N_4467);
xnor U4585 (N_4585,N_4445,N_4361);
nor U4586 (N_4586,N_4412,N_4340);
nor U4587 (N_4587,N_4407,N_4437);
nand U4588 (N_4588,N_4387,N_4346);
nand U4589 (N_4589,N_4363,N_4360);
xnor U4590 (N_4590,N_4447,N_4358);
and U4591 (N_4591,N_4415,N_4432);
or U4592 (N_4592,N_4411,N_4367);
xnor U4593 (N_4593,N_4420,N_4439);
and U4594 (N_4594,N_4390,N_4360);
nand U4595 (N_4595,N_4408,N_4472);
xor U4596 (N_4596,N_4341,N_4443);
nor U4597 (N_4597,N_4426,N_4404);
xor U4598 (N_4598,N_4394,N_4465);
or U4599 (N_4599,N_4462,N_4383);
xnor U4600 (N_4600,N_4381,N_4357);
xnor U4601 (N_4601,N_4351,N_4459);
nor U4602 (N_4602,N_4447,N_4456);
nor U4603 (N_4603,N_4322,N_4375);
xor U4604 (N_4604,N_4351,N_4328);
or U4605 (N_4605,N_4383,N_4444);
xor U4606 (N_4606,N_4461,N_4352);
xnor U4607 (N_4607,N_4375,N_4430);
nand U4608 (N_4608,N_4393,N_4352);
nor U4609 (N_4609,N_4344,N_4459);
nand U4610 (N_4610,N_4442,N_4428);
nor U4611 (N_4611,N_4470,N_4339);
nor U4612 (N_4612,N_4337,N_4434);
nor U4613 (N_4613,N_4360,N_4455);
or U4614 (N_4614,N_4354,N_4394);
xor U4615 (N_4615,N_4366,N_4335);
and U4616 (N_4616,N_4438,N_4379);
and U4617 (N_4617,N_4419,N_4473);
nor U4618 (N_4618,N_4411,N_4391);
xor U4619 (N_4619,N_4453,N_4366);
nand U4620 (N_4620,N_4468,N_4478);
nor U4621 (N_4621,N_4465,N_4320);
and U4622 (N_4622,N_4454,N_4386);
nor U4623 (N_4623,N_4380,N_4361);
nor U4624 (N_4624,N_4419,N_4336);
or U4625 (N_4625,N_4323,N_4326);
nor U4626 (N_4626,N_4466,N_4461);
xor U4627 (N_4627,N_4387,N_4337);
or U4628 (N_4628,N_4373,N_4461);
and U4629 (N_4629,N_4387,N_4361);
nand U4630 (N_4630,N_4345,N_4435);
nand U4631 (N_4631,N_4419,N_4369);
nand U4632 (N_4632,N_4460,N_4444);
and U4633 (N_4633,N_4403,N_4478);
and U4634 (N_4634,N_4435,N_4323);
or U4635 (N_4635,N_4339,N_4461);
and U4636 (N_4636,N_4471,N_4359);
nand U4637 (N_4637,N_4462,N_4393);
xor U4638 (N_4638,N_4438,N_4375);
nor U4639 (N_4639,N_4385,N_4471);
nand U4640 (N_4640,N_4497,N_4551);
or U4641 (N_4641,N_4518,N_4571);
or U4642 (N_4642,N_4535,N_4582);
or U4643 (N_4643,N_4558,N_4591);
nand U4644 (N_4644,N_4512,N_4519);
or U4645 (N_4645,N_4505,N_4619);
and U4646 (N_4646,N_4576,N_4536);
nand U4647 (N_4647,N_4483,N_4574);
or U4648 (N_4648,N_4547,N_4527);
or U4649 (N_4649,N_4623,N_4542);
nand U4650 (N_4650,N_4639,N_4584);
or U4651 (N_4651,N_4595,N_4612);
or U4652 (N_4652,N_4570,N_4564);
and U4653 (N_4653,N_4525,N_4601);
and U4654 (N_4654,N_4482,N_4572);
nor U4655 (N_4655,N_4569,N_4605);
or U4656 (N_4656,N_4524,N_4626);
xnor U4657 (N_4657,N_4538,N_4603);
xor U4658 (N_4658,N_4609,N_4622);
or U4659 (N_4659,N_4490,N_4568);
nor U4660 (N_4660,N_4631,N_4621);
or U4661 (N_4661,N_4526,N_4579);
nor U4662 (N_4662,N_4592,N_4606);
nand U4663 (N_4663,N_4607,N_4593);
xor U4664 (N_4664,N_4540,N_4509);
or U4665 (N_4665,N_4585,N_4562);
and U4666 (N_4666,N_4630,N_4628);
nand U4667 (N_4667,N_4629,N_4638);
nor U4668 (N_4668,N_4632,N_4545);
xor U4669 (N_4669,N_4517,N_4557);
nor U4670 (N_4670,N_4559,N_4531);
xnor U4671 (N_4671,N_4481,N_4523);
or U4672 (N_4672,N_4549,N_4598);
and U4673 (N_4673,N_4560,N_4521);
nand U4674 (N_4674,N_4501,N_4548);
nor U4675 (N_4675,N_4590,N_4533);
xor U4676 (N_4676,N_4508,N_4596);
nor U4677 (N_4677,N_4513,N_4600);
nor U4678 (N_4678,N_4495,N_4633);
nand U4679 (N_4679,N_4511,N_4520);
xnor U4680 (N_4680,N_4502,N_4565);
nor U4681 (N_4681,N_4615,N_4566);
nand U4682 (N_4682,N_4496,N_4494);
and U4683 (N_4683,N_4581,N_4586);
xnor U4684 (N_4684,N_4516,N_4594);
nand U4685 (N_4685,N_4627,N_4580);
nor U4686 (N_4686,N_4563,N_4550);
nand U4687 (N_4687,N_4561,N_4634);
xor U4688 (N_4688,N_4489,N_4553);
xor U4689 (N_4689,N_4539,N_4491);
nor U4690 (N_4690,N_4500,N_4487);
or U4691 (N_4691,N_4556,N_4537);
and U4692 (N_4692,N_4578,N_4493);
or U4693 (N_4693,N_4552,N_4546);
and U4694 (N_4694,N_4617,N_4602);
or U4695 (N_4695,N_4583,N_4543);
xor U4696 (N_4696,N_4503,N_4624);
nand U4697 (N_4697,N_4588,N_4530);
and U4698 (N_4698,N_4504,N_4589);
nor U4699 (N_4699,N_4604,N_4485);
nor U4700 (N_4700,N_4488,N_4573);
and U4701 (N_4701,N_4567,N_4534);
xor U4702 (N_4702,N_4610,N_4613);
and U4703 (N_4703,N_4544,N_4541);
nand U4704 (N_4704,N_4486,N_4528);
or U4705 (N_4705,N_4532,N_4611);
or U4706 (N_4706,N_4492,N_4554);
nor U4707 (N_4707,N_4635,N_4484);
and U4708 (N_4708,N_4480,N_4587);
nand U4709 (N_4709,N_4510,N_4618);
xor U4710 (N_4710,N_4636,N_4575);
and U4711 (N_4711,N_4507,N_4616);
and U4712 (N_4712,N_4515,N_4625);
and U4713 (N_4713,N_4506,N_4620);
nor U4714 (N_4714,N_4514,N_4637);
nor U4715 (N_4715,N_4577,N_4498);
nor U4716 (N_4716,N_4529,N_4555);
xnor U4717 (N_4717,N_4499,N_4597);
xor U4718 (N_4718,N_4614,N_4599);
or U4719 (N_4719,N_4522,N_4608);
xnor U4720 (N_4720,N_4607,N_4532);
nand U4721 (N_4721,N_4563,N_4534);
or U4722 (N_4722,N_4543,N_4518);
xnor U4723 (N_4723,N_4527,N_4495);
or U4724 (N_4724,N_4589,N_4522);
xor U4725 (N_4725,N_4632,N_4565);
xnor U4726 (N_4726,N_4580,N_4608);
nand U4727 (N_4727,N_4562,N_4506);
or U4728 (N_4728,N_4631,N_4517);
xor U4729 (N_4729,N_4637,N_4517);
and U4730 (N_4730,N_4610,N_4547);
xor U4731 (N_4731,N_4483,N_4502);
and U4732 (N_4732,N_4534,N_4621);
xnor U4733 (N_4733,N_4579,N_4520);
and U4734 (N_4734,N_4626,N_4501);
or U4735 (N_4735,N_4639,N_4563);
nor U4736 (N_4736,N_4639,N_4512);
nor U4737 (N_4737,N_4624,N_4637);
xor U4738 (N_4738,N_4620,N_4592);
xnor U4739 (N_4739,N_4506,N_4624);
nor U4740 (N_4740,N_4584,N_4506);
nor U4741 (N_4741,N_4638,N_4570);
nor U4742 (N_4742,N_4544,N_4558);
or U4743 (N_4743,N_4570,N_4550);
nor U4744 (N_4744,N_4523,N_4485);
xor U4745 (N_4745,N_4571,N_4558);
or U4746 (N_4746,N_4549,N_4556);
and U4747 (N_4747,N_4493,N_4615);
and U4748 (N_4748,N_4557,N_4604);
nor U4749 (N_4749,N_4554,N_4568);
xor U4750 (N_4750,N_4515,N_4495);
nand U4751 (N_4751,N_4578,N_4597);
nand U4752 (N_4752,N_4617,N_4529);
and U4753 (N_4753,N_4569,N_4483);
xnor U4754 (N_4754,N_4568,N_4630);
xor U4755 (N_4755,N_4535,N_4529);
nor U4756 (N_4756,N_4613,N_4540);
xnor U4757 (N_4757,N_4521,N_4610);
nor U4758 (N_4758,N_4559,N_4574);
xnor U4759 (N_4759,N_4553,N_4523);
or U4760 (N_4760,N_4551,N_4480);
nand U4761 (N_4761,N_4619,N_4512);
xnor U4762 (N_4762,N_4528,N_4571);
nor U4763 (N_4763,N_4485,N_4631);
xor U4764 (N_4764,N_4525,N_4570);
xor U4765 (N_4765,N_4620,N_4582);
nand U4766 (N_4766,N_4484,N_4500);
xor U4767 (N_4767,N_4543,N_4620);
and U4768 (N_4768,N_4509,N_4563);
nand U4769 (N_4769,N_4584,N_4589);
nand U4770 (N_4770,N_4569,N_4628);
nor U4771 (N_4771,N_4586,N_4538);
xor U4772 (N_4772,N_4513,N_4618);
or U4773 (N_4773,N_4634,N_4560);
xnor U4774 (N_4774,N_4561,N_4569);
and U4775 (N_4775,N_4502,N_4638);
xnor U4776 (N_4776,N_4490,N_4636);
and U4777 (N_4777,N_4620,N_4635);
or U4778 (N_4778,N_4520,N_4532);
nand U4779 (N_4779,N_4580,N_4521);
nor U4780 (N_4780,N_4550,N_4591);
or U4781 (N_4781,N_4513,N_4575);
and U4782 (N_4782,N_4625,N_4612);
nand U4783 (N_4783,N_4585,N_4615);
nor U4784 (N_4784,N_4574,N_4491);
and U4785 (N_4785,N_4491,N_4486);
or U4786 (N_4786,N_4572,N_4575);
or U4787 (N_4787,N_4595,N_4511);
nand U4788 (N_4788,N_4536,N_4583);
nor U4789 (N_4789,N_4495,N_4618);
nand U4790 (N_4790,N_4498,N_4635);
nand U4791 (N_4791,N_4611,N_4519);
xor U4792 (N_4792,N_4524,N_4570);
xnor U4793 (N_4793,N_4597,N_4608);
xnor U4794 (N_4794,N_4523,N_4623);
nor U4795 (N_4795,N_4555,N_4539);
xnor U4796 (N_4796,N_4577,N_4499);
nor U4797 (N_4797,N_4594,N_4508);
nand U4798 (N_4798,N_4590,N_4559);
or U4799 (N_4799,N_4571,N_4593);
and U4800 (N_4800,N_4668,N_4716);
or U4801 (N_4801,N_4659,N_4739);
or U4802 (N_4802,N_4752,N_4732);
nand U4803 (N_4803,N_4669,N_4718);
nand U4804 (N_4804,N_4652,N_4783);
xor U4805 (N_4805,N_4726,N_4684);
and U4806 (N_4806,N_4683,N_4706);
nand U4807 (N_4807,N_4772,N_4787);
xnor U4808 (N_4808,N_4790,N_4743);
and U4809 (N_4809,N_4670,N_4774);
nand U4810 (N_4810,N_4646,N_4736);
nand U4811 (N_4811,N_4758,N_4711);
and U4812 (N_4812,N_4773,N_4696);
and U4813 (N_4813,N_4740,N_4678);
and U4814 (N_4814,N_4697,N_4738);
xnor U4815 (N_4815,N_4653,N_4782);
nor U4816 (N_4816,N_4685,N_4650);
and U4817 (N_4817,N_4759,N_4780);
xor U4818 (N_4818,N_4657,N_4798);
and U4819 (N_4819,N_4680,N_4709);
or U4820 (N_4820,N_4717,N_4761);
xor U4821 (N_4821,N_4705,N_4742);
and U4822 (N_4822,N_4785,N_4745);
nand U4823 (N_4823,N_4640,N_4727);
nor U4824 (N_4824,N_4751,N_4797);
or U4825 (N_4825,N_4651,N_4691);
nand U4826 (N_4826,N_4700,N_4675);
nand U4827 (N_4827,N_4791,N_4744);
nand U4828 (N_4828,N_4710,N_4799);
and U4829 (N_4829,N_4788,N_4704);
xor U4830 (N_4830,N_4663,N_4687);
or U4831 (N_4831,N_4690,N_4676);
or U4832 (N_4832,N_4701,N_4654);
nor U4833 (N_4833,N_4724,N_4768);
xnor U4834 (N_4834,N_4715,N_4760);
and U4835 (N_4835,N_4674,N_4671);
xor U4836 (N_4836,N_4794,N_4689);
nor U4837 (N_4837,N_4703,N_4641);
or U4838 (N_4838,N_4649,N_4725);
nor U4839 (N_4839,N_4757,N_4770);
nand U4840 (N_4840,N_4719,N_4741);
xor U4841 (N_4841,N_4766,N_4664);
nand U4842 (N_4842,N_4686,N_4731);
and U4843 (N_4843,N_4694,N_4655);
xor U4844 (N_4844,N_4765,N_4643);
nor U4845 (N_4845,N_4688,N_4776);
or U4846 (N_4846,N_4793,N_4795);
nand U4847 (N_4847,N_4734,N_4658);
nor U4848 (N_4848,N_4777,N_4660);
xnor U4849 (N_4849,N_4729,N_4702);
xor U4850 (N_4850,N_4707,N_4667);
xor U4851 (N_4851,N_4764,N_4661);
or U4852 (N_4852,N_4728,N_4673);
xor U4853 (N_4853,N_4792,N_4784);
or U4854 (N_4854,N_4642,N_4692);
nand U4855 (N_4855,N_4748,N_4775);
or U4856 (N_4856,N_4763,N_4781);
or U4857 (N_4857,N_4755,N_4698);
and U4858 (N_4858,N_4682,N_4767);
nor U4859 (N_4859,N_4713,N_4665);
nor U4860 (N_4860,N_4722,N_4699);
nand U4861 (N_4861,N_4754,N_4779);
nand U4862 (N_4862,N_4730,N_4747);
nor U4863 (N_4863,N_4693,N_4647);
nand U4864 (N_4864,N_4708,N_4733);
nor U4865 (N_4865,N_4714,N_4662);
and U4866 (N_4866,N_4672,N_4778);
or U4867 (N_4867,N_4771,N_4721);
nor U4868 (N_4868,N_4750,N_4746);
xor U4869 (N_4869,N_4756,N_4679);
nor U4870 (N_4870,N_4645,N_4712);
or U4871 (N_4871,N_4723,N_4695);
or U4872 (N_4872,N_4749,N_4737);
nand U4873 (N_4873,N_4720,N_4644);
or U4874 (N_4874,N_4735,N_4656);
nand U4875 (N_4875,N_4769,N_4789);
nand U4876 (N_4876,N_4786,N_4648);
nor U4877 (N_4877,N_4753,N_4762);
xnor U4878 (N_4878,N_4796,N_4681);
and U4879 (N_4879,N_4677,N_4666);
and U4880 (N_4880,N_4749,N_4644);
or U4881 (N_4881,N_4674,N_4746);
xor U4882 (N_4882,N_4683,N_4653);
nand U4883 (N_4883,N_4747,N_4723);
nand U4884 (N_4884,N_4653,N_4705);
nand U4885 (N_4885,N_4737,N_4697);
xor U4886 (N_4886,N_4665,N_4750);
xnor U4887 (N_4887,N_4714,N_4641);
or U4888 (N_4888,N_4709,N_4696);
and U4889 (N_4889,N_4766,N_4693);
and U4890 (N_4890,N_4719,N_4676);
nand U4891 (N_4891,N_4746,N_4787);
nor U4892 (N_4892,N_4770,N_4666);
nor U4893 (N_4893,N_4688,N_4648);
or U4894 (N_4894,N_4728,N_4799);
xor U4895 (N_4895,N_4747,N_4774);
nor U4896 (N_4896,N_4746,N_4723);
nand U4897 (N_4897,N_4720,N_4665);
or U4898 (N_4898,N_4679,N_4746);
or U4899 (N_4899,N_4744,N_4797);
nand U4900 (N_4900,N_4734,N_4732);
and U4901 (N_4901,N_4737,N_4710);
and U4902 (N_4902,N_4659,N_4692);
or U4903 (N_4903,N_4745,N_4787);
nand U4904 (N_4904,N_4645,N_4702);
or U4905 (N_4905,N_4783,N_4657);
xnor U4906 (N_4906,N_4735,N_4765);
xnor U4907 (N_4907,N_4771,N_4786);
or U4908 (N_4908,N_4742,N_4645);
and U4909 (N_4909,N_4673,N_4698);
and U4910 (N_4910,N_4767,N_4794);
nor U4911 (N_4911,N_4790,N_4708);
nor U4912 (N_4912,N_4667,N_4660);
nand U4913 (N_4913,N_4781,N_4795);
and U4914 (N_4914,N_4710,N_4773);
xor U4915 (N_4915,N_4792,N_4650);
and U4916 (N_4916,N_4796,N_4728);
nor U4917 (N_4917,N_4790,N_4726);
or U4918 (N_4918,N_4743,N_4703);
and U4919 (N_4919,N_4667,N_4709);
or U4920 (N_4920,N_4659,N_4780);
nand U4921 (N_4921,N_4768,N_4682);
xor U4922 (N_4922,N_4658,N_4657);
or U4923 (N_4923,N_4677,N_4744);
xnor U4924 (N_4924,N_4753,N_4771);
nand U4925 (N_4925,N_4650,N_4728);
nand U4926 (N_4926,N_4664,N_4758);
and U4927 (N_4927,N_4749,N_4642);
and U4928 (N_4928,N_4731,N_4659);
nor U4929 (N_4929,N_4754,N_4721);
or U4930 (N_4930,N_4681,N_4722);
and U4931 (N_4931,N_4691,N_4790);
nor U4932 (N_4932,N_4666,N_4651);
or U4933 (N_4933,N_4781,N_4687);
nor U4934 (N_4934,N_4754,N_4648);
nor U4935 (N_4935,N_4680,N_4797);
nor U4936 (N_4936,N_4745,N_4775);
nor U4937 (N_4937,N_4726,N_4718);
nor U4938 (N_4938,N_4745,N_4740);
or U4939 (N_4939,N_4707,N_4746);
nor U4940 (N_4940,N_4770,N_4696);
and U4941 (N_4941,N_4799,N_4742);
or U4942 (N_4942,N_4798,N_4779);
or U4943 (N_4943,N_4738,N_4754);
or U4944 (N_4944,N_4766,N_4792);
and U4945 (N_4945,N_4795,N_4728);
nand U4946 (N_4946,N_4699,N_4798);
and U4947 (N_4947,N_4723,N_4754);
xor U4948 (N_4948,N_4686,N_4657);
nor U4949 (N_4949,N_4640,N_4682);
or U4950 (N_4950,N_4762,N_4679);
or U4951 (N_4951,N_4750,N_4653);
or U4952 (N_4952,N_4662,N_4690);
xnor U4953 (N_4953,N_4695,N_4657);
xor U4954 (N_4954,N_4651,N_4653);
or U4955 (N_4955,N_4785,N_4640);
nor U4956 (N_4956,N_4778,N_4640);
xor U4957 (N_4957,N_4681,N_4797);
xnor U4958 (N_4958,N_4664,N_4656);
and U4959 (N_4959,N_4714,N_4752);
nand U4960 (N_4960,N_4857,N_4820);
or U4961 (N_4961,N_4817,N_4924);
nand U4962 (N_4962,N_4930,N_4811);
and U4963 (N_4963,N_4807,N_4844);
nor U4964 (N_4964,N_4947,N_4867);
nand U4965 (N_4965,N_4821,N_4878);
nor U4966 (N_4966,N_4804,N_4923);
nor U4967 (N_4967,N_4941,N_4819);
nand U4968 (N_4968,N_4866,N_4861);
and U4969 (N_4969,N_4925,N_4939);
nor U4970 (N_4970,N_4943,N_4920);
or U4971 (N_4971,N_4829,N_4928);
nand U4972 (N_4972,N_4934,N_4802);
xnor U4973 (N_4973,N_4892,N_4904);
or U4974 (N_4974,N_4942,N_4810);
or U4975 (N_4975,N_4908,N_4872);
nor U4976 (N_4976,N_4822,N_4956);
nand U4977 (N_4977,N_4880,N_4842);
nand U4978 (N_4978,N_4865,N_4826);
xnor U4979 (N_4979,N_4903,N_4834);
xnor U4980 (N_4980,N_4839,N_4882);
or U4981 (N_4981,N_4851,N_4937);
nand U4982 (N_4982,N_4877,N_4957);
xnor U4983 (N_4983,N_4843,N_4800);
or U4984 (N_4984,N_4899,N_4913);
nor U4985 (N_4985,N_4894,N_4909);
and U4986 (N_4986,N_4838,N_4900);
nand U4987 (N_4987,N_4863,N_4806);
or U4988 (N_4988,N_4835,N_4938);
and U4989 (N_4989,N_4832,N_4946);
and U4990 (N_4990,N_4907,N_4801);
nand U4991 (N_4991,N_4836,N_4849);
xnor U4992 (N_4992,N_4953,N_4933);
nor U4993 (N_4993,N_4911,N_4895);
nand U4994 (N_4994,N_4809,N_4935);
and U4995 (N_4995,N_4927,N_4860);
and U4996 (N_4996,N_4846,N_4855);
xor U4997 (N_4997,N_4958,N_4897);
and U4998 (N_4998,N_4869,N_4827);
xor U4999 (N_4999,N_4856,N_4906);
nand U5000 (N_5000,N_4959,N_4887);
or U5001 (N_5001,N_4875,N_4944);
nand U5002 (N_5002,N_4954,N_4814);
nand U5003 (N_5003,N_4929,N_4818);
nand U5004 (N_5004,N_4837,N_4828);
or U5005 (N_5005,N_4902,N_4864);
and U5006 (N_5006,N_4841,N_4884);
nor U5007 (N_5007,N_4888,N_4830);
nor U5008 (N_5008,N_4850,N_4910);
xor U5009 (N_5009,N_4840,N_4813);
and U5010 (N_5010,N_4881,N_4912);
and U5011 (N_5011,N_4896,N_4859);
or U5012 (N_5012,N_4917,N_4803);
nand U5013 (N_5013,N_4868,N_4948);
and U5014 (N_5014,N_4916,N_4808);
or U5015 (N_5015,N_4858,N_4815);
nand U5016 (N_5016,N_4898,N_4883);
or U5017 (N_5017,N_4833,N_4873);
xor U5018 (N_5018,N_4870,N_4845);
or U5019 (N_5019,N_4812,N_4891);
nand U5020 (N_5020,N_4874,N_4950);
and U5021 (N_5021,N_4848,N_4852);
nand U5022 (N_5022,N_4952,N_4862);
or U5023 (N_5023,N_4879,N_4876);
nor U5024 (N_5024,N_4805,N_4932);
xor U5025 (N_5025,N_4914,N_4936);
nor U5026 (N_5026,N_4824,N_4940);
nand U5027 (N_5027,N_4945,N_4893);
or U5028 (N_5028,N_4816,N_4853);
and U5029 (N_5029,N_4955,N_4915);
nand U5030 (N_5030,N_4922,N_4951);
or U5031 (N_5031,N_4889,N_4918);
nand U5032 (N_5032,N_4949,N_4886);
or U5033 (N_5033,N_4854,N_4905);
nand U5034 (N_5034,N_4831,N_4871);
xor U5035 (N_5035,N_4919,N_4890);
and U5036 (N_5036,N_4823,N_4847);
nor U5037 (N_5037,N_4885,N_4931);
nor U5038 (N_5038,N_4921,N_4825);
xor U5039 (N_5039,N_4926,N_4901);
xor U5040 (N_5040,N_4813,N_4822);
nand U5041 (N_5041,N_4941,N_4812);
nand U5042 (N_5042,N_4837,N_4890);
xnor U5043 (N_5043,N_4811,N_4946);
or U5044 (N_5044,N_4809,N_4806);
nor U5045 (N_5045,N_4939,N_4841);
nor U5046 (N_5046,N_4821,N_4943);
nand U5047 (N_5047,N_4844,N_4817);
nor U5048 (N_5048,N_4927,N_4899);
and U5049 (N_5049,N_4943,N_4822);
nand U5050 (N_5050,N_4927,N_4834);
nor U5051 (N_5051,N_4926,N_4955);
nand U5052 (N_5052,N_4956,N_4904);
xnor U5053 (N_5053,N_4826,N_4831);
xor U5054 (N_5054,N_4804,N_4848);
and U5055 (N_5055,N_4880,N_4873);
nor U5056 (N_5056,N_4886,N_4921);
and U5057 (N_5057,N_4841,N_4803);
nor U5058 (N_5058,N_4930,N_4912);
nand U5059 (N_5059,N_4832,N_4918);
nand U5060 (N_5060,N_4837,N_4929);
nor U5061 (N_5061,N_4891,N_4892);
and U5062 (N_5062,N_4847,N_4886);
or U5063 (N_5063,N_4820,N_4851);
or U5064 (N_5064,N_4903,N_4803);
or U5065 (N_5065,N_4957,N_4856);
xnor U5066 (N_5066,N_4812,N_4871);
xor U5067 (N_5067,N_4856,N_4953);
or U5068 (N_5068,N_4864,N_4954);
nor U5069 (N_5069,N_4833,N_4893);
xor U5070 (N_5070,N_4906,N_4894);
xnor U5071 (N_5071,N_4875,N_4924);
xor U5072 (N_5072,N_4954,N_4877);
or U5073 (N_5073,N_4804,N_4864);
xor U5074 (N_5074,N_4801,N_4869);
nand U5075 (N_5075,N_4947,N_4912);
or U5076 (N_5076,N_4875,N_4804);
nand U5077 (N_5077,N_4893,N_4950);
or U5078 (N_5078,N_4833,N_4897);
and U5079 (N_5079,N_4853,N_4900);
nand U5080 (N_5080,N_4907,N_4822);
nor U5081 (N_5081,N_4936,N_4822);
nor U5082 (N_5082,N_4957,N_4834);
xor U5083 (N_5083,N_4805,N_4905);
or U5084 (N_5084,N_4840,N_4810);
nor U5085 (N_5085,N_4913,N_4917);
xnor U5086 (N_5086,N_4854,N_4927);
nor U5087 (N_5087,N_4915,N_4936);
xor U5088 (N_5088,N_4914,N_4938);
or U5089 (N_5089,N_4864,N_4858);
xnor U5090 (N_5090,N_4876,N_4816);
nor U5091 (N_5091,N_4944,N_4824);
xor U5092 (N_5092,N_4931,N_4865);
and U5093 (N_5093,N_4851,N_4880);
nand U5094 (N_5094,N_4946,N_4939);
nor U5095 (N_5095,N_4871,N_4803);
or U5096 (N_5096,N_4805,N_4921);
nand U5097 (N_5097,N_4950,N_4869);
or U5098 (N_5098,N_4940,N_4959);
and U5099 (N_5099,N_4921,N_4873);
or U5100 (N_5100,N_4850,N_4826);
nand U5101 (N_5101,N_4941,N_4944);
nor U5102 (N_5102,N_4878,N_4854);
xor U5103 (N_5103,N_4948,N_4917);
and U5104 (N_5104,N_4912,N_4889);
and U5105 (N_5105,N_4872,N_4876);
or U5106 (N_5106,N_4947,N_4875);
nand U5107 (N_5107,N_4897,N_4926);
xnor U5108 (N_5108,N_4926,N_4833);
and U5109 (N_5109,N_4920,N_4870);
nor U5110 (N_5110,N_4871,N_4865);
nor U5111 (N_5111,N_4906,N_4832);
and U5112 (N_5112,N_4903,N_4816);
xnor U5113 (N_5113,N_4849,N_4801);
xor U5114 (N_5114,N_4841,N_4850);
nand U5115 (N_5115,N_4856,N_4946);
xnor U5116 (N_5116,N_4896,N_4807);
nor U5117 (N_5117,N_4813,N_4958);
or U5118 (N_5118,N_4939,N_4902);
and U5119 (N_5119,N_4954,N_4842);
xor U5120 (N_5120,N_5049,N_4997);
nor U5121 (N_5121,N_5050,N_5089);
nor U5122 (N_5122,N_5001,N_5067);
nand U5123 (N_5123,N_5097,N_5042);
and U5124 (N_5124,N_5044,N_4963);
xnor U5125 (N_5125,N_5118,N_5002);
and U5126 (N_5126,N_5052,N_5039);
or U5127 (N_5127,N_5034,N_5032);
nand U5128 (N_5128,N_4965,N_5104);
or U5129 (N_5129,N_4967,N_4994);
nor U5130 (N_5130,N_5054,N_5110);
nand U5131 (N_5131,N_4983,N_4981);
and U5132 (N_5132,N_5017,N_5005);
nor U5133 (N_5133,N_5011,N_4999);
nor U5134 (N_5134,N_4996,N_4987);
nor U5135 (N_5135,N_5091,N_5012);
nor U5136 (N_5136,N_5101,N_5087);
or U5137 (N_5137,N_5098,N_5119);
and U5138 (N_5138,N_4986,N_5023);
nor U5139 (N_5139,N_5053,N_5024);
xor U5140 (N_5140,N_5021,N_5056);
xor U5141 (N_5141,N_5106,N_4998);
nand U5142 (N_5142,N_4974,N_4979);
xnor U5143 (N_5143,N_5060,N_4973);
nor U5144 (N_5144,N_4975,N_4992);
nand U5145 (N_5145,N_5033,N_5057);
xnor U5146 (N_5146,N_5006,N_5111);
nor U5147 (N_5147,N_5070,N_4988);
xnor U5148 (N_5148,N_5018,N_5061);
xnor U5149 (N_5149,N_5048,N_5062);
and U5150 (N_5150,N_5108,N_5051);
nor U5151 (N_5151,N_4978,N_5043);
nand U5152 (N_5152,N_5115,N_5113);
xor U5153 (N_5153,N_5093,N_5112);
nor U5154 (N_5154,N_5016,N_4982);
and U5155 (N_5155,N_5007,N_5027);
or U5156 (N_5156,N_5000,N_5028);
and U5157 (N_5157,N_5038,N_4966);
or U5158 (N_5158,N_4991,N_5102);
nor U5159 (N_5159,N_5019,N_5073);
nand U5160 (N_5160,N_5059,N_5014);
xor U5161 (N_5161,N_5058,N_5114);
nand U5162 (N_5162,N_4969,N_5013);
and U5163 (N_5163,N_4968,N_4984);
or U5164 (N_5164,N_5090,N_4990);
and U5165 (N_5165,N_5015,N_5008);
and U5166 (N_5166,N_5096,N_5035);
and U5167 (N_5167,N_5076,N_5109);
nor U5168 (N_5168,N_4995,N_5009);
nand U5169 (N_5169,N_4964,N_5105);
and U5170 (N_5170,N_4970,N_4977);
nor U5171 (N_5171,N_5074,N_5065);
nand U5172 (N_5172,N_5045,N_4985);
xor U5173 (N_5173,N_5010,N_5063);
nor U5174 (N_5174,N_5037,N_5020);
nand U5175 (N_5175,N_5066,N_5003);
xor U5176 (N_5176,N_4976,N_5031);
nor U5177 (N_5177,N_5069,N_5085);
nor U5178 (N_5178,N_5022,N_4962);
and U5179 (N_5179,N_4972,N_5092);
or U5180 (N_5180,N_5075,N_5036);
nand U5181 (N_5181,N_5083,N_5026);
xnor U5182 (N_5182,N_5099,N_5068);
xor U5183 (N_5183,N_5055,N_5094);
and U5184 (N_5184,N_5116,N_5072);
nand U5185 (N_5185,N_4989,N_5117);
or U5186 (N_5186,N_5046,N_4961);
xnor U5187 (N_5187,N_5004,N_4971);
or U5188 (N_5188,N_5064,N_4980);
nor U5189 (N_5189,N_5107,N_5030);
nor U5190 (N_5190,N_5071,N_5100);
nand U5191 (N_5191,N_5080,N_5029);
nand U5192 (N_5192,N_4960,N_5103);
xor U5193 (N_5193,N_4993,N_5088);
and U5194 (N_5194,N_5041,N_5095);
and U5195 (N_5195,N_5086,N_5040);
xnor U5196 (N_5196,N_5047,N_5084);
or U5197 (N_5197,N_5078,N_5082);
and U5198 (N_5198,N_5077,N_5079);
and U5199 (N_5199,N_5081,N_5025);
nor U5200 (N_5200,N_5004,N_5082);
or U5201 (N_5201,N_5057,N_5064);
nor U5202 (N_5202,N_5109,N_5088);
or U5203 (N_5203,N_5078,N_4987);
nand U5204 (N_5204,N_5097,N_5104);
xnor U5205 (N_5205,N_5007,N_5002);
nand U5206 (N_5206,N_5112,N_5069);
nor U5207 (N_5207,N_4973,N_5003);
or U5208 (N_5208,N_5086,N_5085);
and U5209 (N_5209,N_5098,N_5100);
nor U5210 (N_5210,N_5101,N_5085);
or U5211 (N_5211,N_5070,N_5096);
and U5212 (N_5212,N_5040,N_5057);
and U5213 (N_5213,N_5102,N_5071);
xnor U5214 (N_5214,N_4982,N_5081);
and U5215 (N_5215,N_4981,N_5049);
xnor U5216 (N_5216,N_4968,N_5068);
nor U5217 (N_5217,N_5088,N_5028);
nand U5218 (N_5218,N_5073,N_5059);
and U5219 (N_5219,N_5046,N_5017);
and U5220 (N_5220,N_5109,N_5040);
xnor U5221 (N_5221,N_5091,N_5045);
xnor U5222 (N_5222,N_5054,N_4977);
nor U5223 (N_5223,N_5009,N_4980);
and U5224 (N_5224,N_5098,N_5004);
nor U5225 (N_5225,N_4966,N_5105);
or U5226 (N_5226,N_5098,N_5057);
nor U5227 (N_5227,N_5052,N_5053);
or U5228 (N_5228,N_5118,N_5094);
nand U5229 (N_5229,N_5081,N_5002);
nor U5230 (N_5230,N_5014,N_5008);
and U5231 (N_5231,N_5099,N_4991);
nand U5232 (N_5232,N_5101,N_5032);
or U5233 (N_5233,N_5119,N_5036);
xnor U5234 (N_5234,N_5042,N_5053);
or U5235 (N_5235,N_5038,N_4988);
nor U5236 (N_5236,N_4997,N_5033);
nand U5237 (N_5237,N_5078,N_5095);
xor U5238 (N_5238,N_5083,N_4974);
nand U5239 (N_5239,N_5017,N_5011);
and U5240 (N_5240,N_4966,N_5113);
xor U5241 (N_5241,N_5105,N_5001);
xnor U5242 (N_5242,N_5084,N_5071);
nor U5243 (N_5243,N_4989,N_5116);
xor U5244 (N_5244,N_4999,N_4979);
xor U5245 (N_5245,N_4973,N_5086);
and U5246 (N_5246,N_5055,N_5063);
nor U5247 (N_5247,N_5017,N_4962);
xnor U5248 (N_5248,N_5041,N_5002);
nand U5249 (N_5249,N_4988,N_5101);
nand U5250 (N_5250,N_5115,N_5031);
nand U5251 (N_5251,N_5029,N_5010);
or U5252 (N_5252,N_4971,N_5007);
and U5253 (N_5253,N_5073,N_5070);
xnor U5254 (N_5254,N_4978,N_5001);
xnor U5255 (N_5255,N_5050,N_5067);
nor U5256 (N_5256,N_5104,N_5071);
or U5257 (N_5257,N_5086,N_5084);
or U5258 (N_5258,N_4967,N_5112);
nand U5259 (N_5259,N_5035,N_4983);
nand U5260 (N_5260,N_5096,N_5012);
or U5261 (N_5261,N_5002,N_5058);
nor U5262 (N_5262,N_5058,N_4961);
nand U5263 (N_5263,N_5110,N_5030);
xor U5264 (N_5264,N_5049,N_5004);
nor U5265 (N_5265,N_5023,N_4988);
nand U5266 (N_5266,N_4962,N_4971);
nor U5267 (N_5267,N_4962,N_5051);
nand U5268 (N_5268,N_5039,N_5054);
nor U5269 (N_5269,N_5075,N_5064);
and U5270 (N_5270,N_5011,N_5048);
and U5271 (N_5271,N_5097,N_5079);
or U5272 (N_5272,N_4962,N_5068);
and U5273 (N_5273,N_5091,N_5054);
nor U5274 (N_5274,N_5008,N_5021);
or U5275 (N_5275,N_4960,N_5039);
or U5276 (N_5276,N_5037,N_5041);
nor U5277 (N_5277,N_5116,N_5060);
and U5278 (N_5278,N_5025,N_5080);
nand U5279 (N_5279,N_5078,N_5092);
and U5280 (N_5280,N_5223,N_5202);
and U5281 (N_5281,N_5169,N_5271);
nor U5282 (N_5282,N_5132,N_5150);
and U5283 (N_5283,N_5253,N_5221);
or U5284 (N_5284,N_5252,N_5120);
and U5285 (N_5285,N_5213,N_5224);
nand U5286 (N_5286,N_5207,N_5197);
xor U5287 (N_5287,N_5265,N_5159);
nand U5288 (N_5288,N_5270,N_5130);
nand U5289 (N_5289,N_5277,N_5240);
and U5290 (N_5290,N_5235,N_5145);
and U5291 (N_5291,N_5186,N_5239);
nand U5292 (N_5292,N_5243,N_5218);
nor U5293 (N_5293,N_5185,N_5173);
nand U5294 (N_5294,N_5268,N_5234);
or U5295 (N_5295,N_5216,N_5155);
xor U5296 (N_5296,N_5236,N_5175);
nor U5297 (N_5297,N_5212,N_5248);
xnor U5298 (N_5298,N_5238,N_5228);
or U5299 (N_5299,N_5188,N_5262);
or U5300 (N_5300,N_5138,N_5184);
nor U5301 (N_5301,N_5269,N_5136);
and U5302 (N_5302,N_5220,N_5249);
and U5303 (N_5303,N_5140,N_5133);
and U5304 (N_5304,N_5166,N_5196);
nand U5305 (N_5305,N_5122,N_5247);
or U5306 (N_5306,N_5199,N_5137);
or U5307 (N_5307,N_5205,N_5215);
xnor U5308 (N_5308,N_5135,N_5172);
nand U5309 (N_5309,N_5255,N_5210);
nor U5310 (N_5310,N_5161,N_5157);
nor U5311 (N_5311,N_5274,N_5171);
or U5312 (N_5312,N_5192,N_5273);
or U5313 (N_5313,N_5148,N_5194);
nor U5314 (N_5314,N_5127,N_5260);
nand U5315 (N_5315,N_5214,N_5151);
and U5316 (N_5316,N_5183,N_5144);
and U5317 (N_5317,N_5208,N_5230);
or U5318 (N_5318,N_5142,N_5168);
xor U5319 (N_5319,N_5164,N_5272);
nand U5320 (N_5320,N_5242,N_5254);
and U5321 (N_5321,N_5229,N_5258);
and U5322 (N_5322,N_5162,N_5227);
or U5323 (N_5323,N_5189,N_5134);
xor U5324 (N_5324,N_5178,N_5206);
or U5325 (N_5325,N_5126,N_5129);
or U5326 (N_5326,N_5200,N_5244);
xor U5327 (N_5327,N_5225,N_5222);
and U5328 (N_5328,N_5267,N_5232);
and U5329 (N_5329,N_5190,N_5279);
and U5330 (N_5330,N_5211,N_5245);
and U5331 (N_5331,N_5198,N_5191);
and U5332 (N_5332,N_5201,N_5124);
nor U5333 (N_5333,N_5193,N_5147);
or U5334 (N_5334,N_5231,N_5219);
nor U5335 (N_5335,N_5176,N_5264);
nor U5336 (N_5336,N_5123,N_5180);
xor U5337 (N_5337,N_5275,N_5257);
and U5338 (N_5338,N_5182,N_5163);
and U5339 (N_5339,N_5156,N_5165);
nor U5340 (N_5340,N_5278,N_5246);
and U5341 (N_5341,N_5146,N_5204);
nor U5342 (N_5342,N_5167,N_5251);
nand U5343 (N_5343,N_5143,N_5263);
xor U5344 (N_5344,N_5152,N_5259);
xor U5345 (N_5345,N_5217,N_5226);
or U5346 (N_5346,N_5177,N_5153);
and U5347 (N_5347,N_5256,N_5170);
xor U5348 (N_5348,N_5128,N_5241);
nand U5349 (N_5349,N_5250,N_5174);
nand U5350 (N_5350,N_5179,N_5266);
and U5351 (N_5351,N_5209,N_5187);
nand U5352 (N_5352,N_5261,N_5237);
nand U5353 (N_5353,N_5121,N_5141);
or U5354 (N_5354,N_5203,N_5276);
and U5355 (N_5355,N_5149,N_5154);
and U5356 (N_5356,N_5181,N_5233);
xnor U5357 (N_5357,N_5139,N_5158);
nor U5358 (N_5358,N_5125,N_5131);
or U5359 (N_5359,N_5160,N_5195);
xor U5360 (N_5360,N_5151,N_5195);
and U5361 (N_5361,N_5206,N_5251);
or U5362 (N_5362,N_5251,N_5267);
or U5363 (N_5363,N_5245,N_5182);
nand U5364 (N_5364,N_5238,N_5142);
nand U5365 (N_5365,N_5176,N_5228);
or U5366 (N_5366,N_5141,N_5266);
xor U5367 (N_5367,N_5211,N_5195);
xnor U5368 (N_5368,N_5184,N_5200);
xnor U5369 (N_5369,N_5205,N_5155);
xnor U5370 (N_5370,N_5147,N_5272);
xnor U5371 (N_5371,N_5257,N_5152);
nor U5372 (N_5372,N_5236,N_5246);
xnor U5373 (N_5373,N_5239,N_5170);
xor U5374 (N_5374,N_5166,N_5126);
nor U5375 (N_5375,N_5140,N_5234);
nor U5376 (N_5376,N_5217,N_5227);
or U5377 (N_5377,N_5265,N_5151);
xnor U5378 (N_5378,N_5141,N_5175);
nand U5379 (N_5379,N_5176,N_5144);
nand U5380 (N_5380,N_5218,N_5131);
nand U5381 (N_5381,N_5251,N_5210);
nand U5382 (N_5382,N_5181,N_5212);
nand U5383 (N_5383,N_5256,N_5180);
and U5384 (N_5384,N_5134,N_5163);
and U5385 (N_5385,N_5161,N_5162);
or U5386 (N_5386,N_5208,N_5139);
nor U5387 (N_5387,N_5266,N_5202);
nand U5388 (N_5388,N_5262,N_5155);
nor U5389 (N_5389,N_5179,N_5157);
nand U5390 (N_5390,N_5150,N_5210);
nand U5391 (N_5391,N_5203,N_5262);
nand U5392 (N_5392,N_5120,N_5169);
nand U5393 (N_5393,N_5159,N_5156);
or U5394 (N_5394,N_5207,N_5138);
nor U5395 (N_5395,N_5152,N_5127);
xnor U5396 (N_5396,N_5266,N_5132);
nor U5397 (N_5397,N_5201,N_5142);
nor U5398 (N_5398,N_5126,N_5151);
and U5399 (N_5399,N_5253,N_5163);
xnor U5400 (N_5400,N_5188,N_5212);
or U5401 (N_5401,N_5271,N_5232);
xor U5402 (N_5402,N_5198,N_5174);
or U5403 (N_5403,N_5206,N_5209);
or U5404 (N_5404,N_5142,N_5191);
and U5405 (N_5405,N_5159,N_5224);
or U5406 (N_5406,N_5159,N_5212);
and U5407 (N_5407,N_5244,N_5192);
nor U5408 (N_5408,N_5208,N_5239);
nand U5409 (N_5409,N_5229,N_5223);
nand U5410 (N_5410,N_5173,N_5270);
nand U5411 (N_5411,N_5155,N_5217);
and U5412 (N_5412,N_5171,N_5149);
nor U5413 (N_5413,N_5205,N_5199);
and U5414 (N_5414,N_5246,N_5224);
and U5415 (N_5415,N_5245,N_5176);
and U5416 (N_5416,N_5248,N_5151);
or U5417 (N_5417,N_5222,N_5123);
and U5418 (N_5418,N_5161,N_5242);
and U5419 (N_5419,N_5207,N_5145);
nor U5420 (N_5420,N_5186,N_5195);
nand U5421 (N_5421,N_5175,N_5152);
xnor U5422 (N_5422,N_5161,N_5221);
and U5423 (N_5423,N_5265,N_5198);
or U5424 (N_5424,N_5224,N_5197);
xor U5425 (N_5425,N_5123,N_5251);
or U5426 (N_5426,N_5264,N_5165);
nand U5427 (N_5427,N_5263,N_5278);
nor U5428 (N_5428,N_5266,N_5215);
or U5429 (N_5429,N_5176,N_5208);
or U5430 (N_5430,N_5239,N_5176);
or U5431 (N_5431,N_5260,N_5238);
and U5432 (N_5432,N_5196,N_5182);
nand U5433 (N_5433,N_5274,N_5129);
nor U5434 (N_5434,N_5125,N_5124);
xor U5435 (N_5435,N_5154,N_5279);
xnor U5436 (N_5436,N_5184,N_5237);
nand U5437 (N_5437,N_5140,N_5225);
and U5438 (N_5438,N_5206,N_5210);
or U5439 (N_5439,N_5156,N_5188);
nand U5440 (N_5440,N_5429,N_5410);
or U5441 (N_5441,N_5414,N_5357);
nand U5442 (N_5442,N_5289,N_5363);
nand U5443 (N_5443,N_5333,N_5374);
or U5444 (N_5444,N_5425,N_5337);
xor U5445 (N_5445,N_5399,N_5283);
nor U5446 (N_5446,N_5313,N_5325);
nor U5447 (N_5447,N_5411,N_5372);
nor U5448 (N_5448,N_5323,N_5307);
nor U5449 (N_5449,N_5324,N_5382);
or U5450 (N_5450,N_5364,N_5360);
xnor U5451 (N_5451,N_5409,N_5348);
xor U5452 (N_5452,N_5412,N_5401);
and U5453 (N_5453,N_5424,N_5315);
and U5454 (N_5454,N_5303,N_5297);
xnor U5455 (N_5455,N_5370,N_5292);
xor U5456 (N_5456,N_5295,N_5285);
nor U5457 (N_5457,N_5395,N_5334);
and U5458 (N_5458,N_5280,N_5316);
xor U5459 (N_5459,N_5352,N_5415);
nand U5460 (N_5460,N_5435,N_5320);
xor U5461 (N_5461,N_5413,N_5340);
or U5462 (N_5462,N_5419,N_5317);
or U5463 (N_5463,N_5436,N_5390);
xnor U5464 (N_5464,N_5293,N_5304);
or U5465 (N_5465,N_5300,N_5281);
nor U5466 (N_5466,N_5314,N_5329);
nand U5467 (N_5467,N_5383,N_5335);
nand U5468 (N_5468,N_5355,N_5336);
xnor U5469 (N_5469,N_5373,N_5384);
or U5470 (N_5470,N_5402,N_5327);
or U5471 (N_5471,N_5392,N_5438);
xnor U5472 (N_5472,N_5319,N_5432);
xor U5473 (N_5473,N_5321,N_5385);
nand U5474 (N_5474,N_5381,N_5301);
and U5475 (N_5475,N_5408,N_5326);
nor U5476 (N_5476,N_5362,N_5397);
nand U5477 (N_5477,N_5391,N_5369);
and U5478 (N_5478,N_5306,N_5379);
nand U5479 (N_5479,N_5403,N_5430);
nand U5480 (N_5480,N_5346,N_5296);
xor U5481 (N_5481,N_5368,N_5416);
nand U5482 (N_5482,N_5354,N_5349);
nor U5483 (N_5483,N_5387,N_5312);
or U5484 (N_5484,N_5342,N_5339);
nor U5485 (N_5485,N_5291,N_5393);
or U5486 (N_5486,N_5378,N_5328);
or U5487 (N_5487,N_5361,N_5284);
nand U5488 (N_5488,N_5287,N_5431);
and U5489 (N_5489,N_5330,N_5371);
or U5490 (N_5490,N_5418,N_5420);
nand U5491 (N_5491,N_5332,N_5311);
or U5492 (N_5492,N_5400,N_5341);
or U5493 (N_5493,N_5433,N_5437);
or U5494 (N_5494,N_5298,N_5310);
or U5495 (N_5495,N_5439,N_5286);
nand U5496 (N_5496,N_5375,N_5406);
xor U5497 (N_5497,N_5365,N_5318);
nor U5498 (N_5498,N_5396,N_5282);
nor U5499 (N_5499,N_5356,N_5338);
and U5500 (N_5500,N_5343,N_5359);
nor U5501 (N_5501,N_5421,N_5305);
nor U5502 (N_5502,N_5308,N_5350);
nor U5503 (N_5503,N_5377,N_5426);
nor U5504 (N_5504,N_5398,N_5388);
nor U5505 (N_5505,N_5389,N_5331);
nor U5506 (N_5506,N_5347,N_5322);
and U5507 (N_5507,N_5434,N_5376);
nand U5508 (N_5508,N_5344,N_5423);
nand U5509 (N_5509,N_5358,N_5380);
or U5510 (N_5510,N_5394,N_5345);
nand U5511 (N_5511,N_5353,N_5427);
or U5512 (N_5512,N_5367,N_5290);
nand U5513 (N_5513,N_5294,N_5351);
nor U5514 (N_5514,N_5417,N_5309);
and U5515 (N_5515,N_5288,N_5428);
xor U5516 (N_5516,N_5422,N_5302);
and U5517 (N_5517,N_5407,N_5386);
nor U5518 (N_5518,N_5299,N_5404);
nand U5519 (N_5519,N_5405,N_5366);
or U5520 (N_5520,N_5412,N_5292);
nor U5521 (N_5521,N_5394,N_5333);
and U5522 (N_5522,N_5328,N_5399);
nor U5523 (N_5523,N_5395,N_5359);
xor U5524 (N_5524,N_5355,N_5285);
and U5525 (N_5525,N_5393,N_5346);
and U5526 (N_5526,N_5339,N_5416);
nor U5527 (N_5527,N_5302,N_5429);
nor U5528 (N_5528,N_5362,N_5352);
xnor U5529 (N_5529,N_5406,N_5307);
and U5530 (N_5530,N_5379,N_5310);
and U5531 (N_5531,N_5294,N_5281);
and U5532 (N_5532,N_5434,N_5405);
and U5533 (N_5533,N_5379,N_5383);
nor U5534 (N_5534,N_5403,N_5439);
nor U5535 (N_5535,N_5418,N_5343);
or U5536 (N_5536,N_5328,N_5368);
nand U5537 (N_5537,N_5348,N_5282);
or U5538 (N_5538,N_5344,N_5410);
xnor U5539 (N_5539,N_5394,N_5335);
nand U5540 (N_5540,N_5378,N_5301);
and U5541 (N_5541,N_5281,N_5332);
and U5542 (N_5542,N_5336,N_5365);
and U5543 (N_5543,N_5431,N_5337);
xnor U5544 (N_5544,N_5291,N_5420);
or U5545 (N_5545,N_5371,N_5397);
and U5546 (N_5546,N_5413,N_5377);
nand U5547 (N_5547,N_5364,N_5397);
nor U5548 (N_5548,N_5358,N_5367);
xor U5549 (N_5549,N_5327,N_5361);
or U5550 (N_5550,N_5375,N_5408);
or U5551 (N_5551,N_5371,N_5315);
nor U5552 (N_5552,N_5283,N_5426);
nand U5553 (N_5553,N_5428,N_5333);
nand U5554 (N_5554,N_5317,N_5356);
and U5555 (N_5555,N_5321,N_5421);
and U5556 (N_5556,N_5314,N_5323);
xor U5557 (N_5557,N_5342,N_5415);
or U5558 (N_5558,N_5416,N_5335);
or U5559 (N_5559,N_5394,N_5392);
xnor U5560 (N_5560,N_5398,N_5325);
and U5561 (N_5561,N_5321,N_5412);
and U5562 (N_5562,N_5308,N_5329);
and U5563 (N_5563,N_5365,N_5435);
nand U5564 (N_5564,N_5401,N_5303);
or U5565 (N_5565,N_5402,N_5336);
and U5566 (N_5566,N_5283,N_5367);
and U5567 (N_5567,N_5402,N_5365);
or U5568 (N_5568,N_5431,N_5383);
nor U5569 (N_5569,N_5286,N_5415);
nor U5570 (N_5570,N_5403,N_5373);
and U5571 (N_5571,N_5313,N_5332);
nand U5572 (N_5572,N_5300,N_5416);
nor U5573 (N_5573,N_5380,N_5330);
or U5574 (N_5574,N_5355,N_5288);
nand U5575 (N_5575,N_5439,N_5320);
or U5576 (N_5576,N_5370,N_5390);
nor U5577 (N_5577,N_5374,N_5305);
nor U5578 (N_5578,N_5389,N_5422);
or U5579 (N_5579,N_5409,N_5399);
xor U5580 (N_5580,N_5420,N_5417);
nor U5581 (N_5581,N_5376,N_5314);
nand U5582 (N_5582,N_5331,N_5286);
nor U5583 (N_5583,N_5302,N_5357);
or U5584 (N_5584,N_5437,N_5344);
xor U5585 (N_5585,N_5306,N_5311);
nand U5586 (N_5586,N_5281,N_5417);
or U5587 (N_5587,N_5411,N_5409);
and U5588 (N_5588,N_5433,N_5285);
or U5589 (N_5589,N_5320,N_5415);
nand U5590 (N_5590,N_5280,N_5387);
nand U5591 (N_5591,N_5358,N_5439);
and U5592 (N_5592,N_5324,N_5378);
xnor U5593 (N_5593,N_5324,N_5361);
xnor U5594 (N_5594,N_5381,N_5435);
nor U5595 (N_5595,N_5280,N_5412);
or U5596 (N_5596,N_5290,N_5318);
nor U5597 (N_5597,N_5294,N_5320);
and U5598 (N_5598,N_5400,N_5295);
and U5599 (N_5599,N_5296,N_5325);
xnor U5600 (N_5600,N_5522,N_5549);
nor U5601 (N_5601,N_5570,N_5561);
or U5602 (N_5602,N_5445,N_5457);
nor U5603 (N_5603,N_5582,N_5494);
xor U5604 (N_5604,N_5528,N_5507);
nor U5605 (N_5605,N_5444,N_5550);
or U5606 (N_5606,N_5486,N_5474);
or U5607 (N_5607,N_5586,N_5490);
nand U5608 (N_5608,N_5455,N_5594);
nand U5609 (N_5609,N_5502,N_5590);
and U5610 (N_5610,N_5596,N_5511);
nor U5611 (N_5611,N_5534,N_5532);
nand U5612 (N_5612,N_5493,N_5525);
and U5613 (N_5613,N_5524,N_5589);
or U5614 (N_5614,N_5574,N_5446);
xnor U5615 (N_5615,N_5587,N_5479);
nor U5616 (N_5616,N_5488,N_5536);
or U5617 (N_5617,N_5468,N_5461);
or U5618 (N_5618,N_5505,N_5448);
or U5619 (N_5619,N_5471,N_5571);
or U5620 (N_5620,N_5500,N_5492);
xnor U5621 (N_5621,N_5575,N_5567);
xnor U5622 (N_5622,N_5538,N_5593);
and U5623 (N_5623,N_5526,N_5579);
xnor U5624 (N_5624,N_5592,N_5501);
xor U5625 (N_5625,N_5581,N_5520);
or U5626 (N_5626,N_5459,N_5475);
or U5627 (N_5627,N_5460,N_5515);
and U5628 (N_5628,N_5476,N_5449);
or U5629 (N_5629,N_5440,N_5477);
xor U5630 (N_5630,N_5481,N_5518);
or U5631 (N_5631,N_5497,N_5458);
and U5632 (N_5632,N_5566,N_5578);
nor U5633 (N_5633,N_5463,N_5441);
nand U5634 (N_5634,N_5531,N_5560);
nand U5635 (N_5635,N_5558,N_5473);
or U5636 (N_5636,N_5495,N_5591);
xnor U5637 (N_5637,N_5484,N_5453);
and U5638 (N_5638,N_5553,N_5509);
nor U5639 (N_5639,N_5510,N_5521);
or U5640 (N_5640,N_5530,N_5583);
or U5641 (N_5641,N_5540,N_5564);
nand U5642 (N_5642,N_5454,N_5491);
nor U5643 (N_5643,N_5548,N_5537);
nand U5644 (N_5644,N_5506,N_5523);
nor U5645 (N_5645,N_5563,N_5466);
nor U5646 (N_5646,N_5576,N_5513);
and U5647 (N_5647,N_5512,N_5485);
nor U5648 (N_5648,N_5456,N_5464);
nand U5649 (N_5649,N_5562,N_5472);
or U5650 (N_5650,N_5547,N_5541);
and U5651 (N_5651,N_5483,N_5443);
nand U5652 (N_5652,N_5465,N_5551);
xor U5653 (N_5653,N_5482,N_5543);
and U5654 (N_5654,N_5470,N_5544);
or U5655 (N_5655,N_5556,N_5469);
nor U5656 (N_5656,N_5569,N_5462);
xnor U5657 (N_5657,N_5489,N_5584);
xnor U5658 (N_5658,N_5452,N_5572);
xor U5659 (N_5659,N_5504,N_5442);
xor U5660 (N_5660,N_5598,N_5498);
xnor U5661 (N_5661,N_5499,N_5546);
xnor U5662 (N_5662,N_5552,N_5542);
nor U5663 (N_5663,N_5447,N_5554);
nor U5664 (N_5664,N_5478,N_5496);
nor U5665 (N_5665,N_5565,N_5577);
or U5666 (N_5666,N_5508,N_5573);
nor U5667 (N_5667,N_5451,N_5559);
nand U5668 (N_5668,N_5533,N_5555);
and U5669 (N_5669,N_5514,N_5568);
nor U5670 (N_5670,N_5450,N_5557);
nand U5671 (N_5671,N_5503,N_5599);
nor U5672 (N_5672,N_5467,N_5487);
and U5673 (N_5673,N_5597,N_5527);
nor U5674 (N_5674,N_5580,N_5588);
xnor U5675 (N_5675,N_5585,N_5519);
nand U5676 (N_5676,N_5480,N_5595);
nor U5677 (N_5677,N_5535,N_5545);
nor U5678 (N_5678,N_5529,N_5517);
nor U5679 (N_5679,N_5539,N_5516);
nand U5680 (N_5680,N_5563,N_5573);
and U5681 (N_5681,N_5587,N_5450);
nand U5682 (N_5682,N_5535,N_5504);
or U5683 (N_5683,N_5521,N_5475);
nor U5684 (N_5684,N_5532,N_5558);
nor U5685 (N_5685,N_5502,N_5450);
or U5686 (N_5686,N_5475,N_5479);
and U5687 (N_5687,N_5549,N_5504);
nor U5688 (N_5688,N_5549,N_5516);
nor U5689 (N_5689,N_5519,N_5454);
nand U5690 (N_5690,N_5461,N_5558);
nor U5691 (N_5691,N_5586,N_5481);
and U5692 (N_5692,N_5521,N_5593);
or U5693 (N_5693,N_5492,N_5443);
nor U5694 (N_5694,N_5586,N_5477);
xor U5695 (N_5695,N_5570,N_5508);
or U5696 (N_5696,N_5586,N_5474);
and U5697 (N_5697,N_5576,N_5521);
nor U5698 (N_5698,N_5564,N_5535);
nand U5699 (N_5699,N_5468,N_5583);
nor U5700 (N_5700,N_5521,N_5496);
nor U5701 (N_5701,N_5582,N_5593);
xnor U5702 (N_5702,N_5551,N_5547);
nand U5703 (N_5703,N_5599,N_5533);
nor U5704 (N_5704,N_5558,N_5513);
nor U5705 (N_5705,N_5536,N_5463);
xor U5706 (N_5706,N_5480,N_5521);
and U5707 (N_5707,N_5593,N_5491);
nor U5708 (N_5708,N_5466,N_5498);
nand U5709 (N_5709,N_5561,N_5546);
xor U5710 (N_5710,N_5563,N_5511);
nand U5711 (N_5711,N_5498,N_5461);
nand U5712 (N_5712,N_5545,N_5550);
or U5713 (N_5713,N_5467,N_5582);
xor U5714 (N_5714,N_5515,N_5520);
and U5715 (N_5715,N_5489,N_5590);
nor U5716 (N_5716,N_5538,N_5445);
or U5717 (N_5717,N_5556,N_5444);
nor U5718 (N_5718,N_5577,N_5559);
xnor U5719 (N_5719,N_5581,N_5531);
nand U5720 (N_5720,N_5565,N_5514);
xor U5721 (N_5721,N_5576,N_5580);
nand U5722 (N_5722,N_5536,N_5518);
nor U5723 (N_5723,N_5464,N_5455);
nand U5724 (N_5724,N_5507,N_5544);
nand U5725 (N_5725,N_5567,N_5550);
and U5726 (N_5726,N_5550,N_5469);
xor U5727 (N_5727,N_5572,N_5488);
nand U5728 (N_5728,N_5577,N_5461);
nor U5729 (N_5729,N_5562,N_5530);
or U5730 (N_5730,N_5467,N_5500);
nor U5731 (N_5731,N_5510,N_5596);
or U5732 (N_5732,N_5483,N_5569);
xor U5733 (N_5733,N_5519,N_5596);
nand U5734 (N_5734,N_5442,N_5479);
or U5735 (N_5735,N_5477,N_5473);
nor U5736 (N_5736,N_5548,N_5523);
xnor U5737 (N_5737,N_5510,N_5481);
nor U5738 (N_5738,N_5580,N_5581);
nor U5739 (N_5739,N_5543,N_5469);
and U5740 (N_5740,N_5526,N_5561);
or U5741 (N_5741,N_5487,N_5477);
and U5742 (N_5742,N_5539,N_5593);
and U5743 (N_5743,N_5486,N_5529);
nand U5744 (N_5744,N_5484,N_5488);
and U5745 (N_5745,N_5449,N_5510);
nor U5746 (N_5746,N_5462,N_5499);
nand U5747 (N_5747,N_5495,N_5452);
or U5748 (N_5748,N_5575,N_5463);
nor U5749 (N_5749,N_5570,N_5539);
and U5750 (N_5750,N_5586,N_5576);
or U5751 (N_5751,N_5466,N_5458);
xor U5752 (N_5752,N_5590,N_5598);
nand U5753 (N_5753,N_5580,N_5532);
nor U5754 (N_5754,N_5475,N_5526);
and U5755 (N_5755,N_5525,N_5495);
xor U5756 (N_5756,N_5535,N_5533);
xnor U5757 (N_5757,N_5553,N_5577);
xor U5758 (N_5758,N_5440,N_5533);
nand U5759 (N_5759,N_5542,N_5570);
xnor U5760 (N_5760,N_5704,N_5727);
nor U5761 (N_5761,N_5759,N_5643);
nand U5762 (N_5762,N_5758,N_5736);
or U5763 (N_5763,N_5624,N_5601);
and U5764 (N_5764,N_5635,N_5669);
or U5765 (N_5765,N_5725,N_5737);
nand U5766 (N_5766,N_5667,N_5753);
nand U5767 (N_5767,N_5612,N_5710);
or U5768 (N_5768,N_5700,N_5637);
xor U5769 (N_5769,N_5757,N_5672);
nor U5770 (N_5770,N_5619,N_5680);
nand U5771 (N_5771,N_5653,N_5686);
and U5772 (N_5772,N_5606,N_5638);
nor U5773 (N_5773,N_5731,N_5752);
xnor U5774 (N_5774,N_5675,N_5716);
nand U5775 (N_5775,N_5665,N_5640);
or U5776 (N_5776,N_5683,N_5629);
xor U5777 (N_5777,N_5614,N_5735);
xnor U5778 (N_5778,N_5728,N_5699);
and U5779 (N_5779,N_5655,N_5718);
nor U5780 (N_5780,N_5642,N_5645);
and U5781 (N_5781,N_5673,N_5691);
xnor U5782 (N_5782,N_5600,N_5621);
and U5783 (N_5783,N_5628,N_5715);
or U5784 (N_5784,N_5662,N_5692);
nand U5785 (N_5785,N_5739,N_5751);
and U5786 (N_5786,N_5698,N_5647);
xnor U5787 (N_5787,N_5634,N_5664);
and U5788 (N_5788,N_5663,N_5609);
or U5789 (N_5789,N_5605,N_5616);
xnor U5790 (N_5790,N_5677,N_5696);
or U5791 (N_5791,N_5633,N_5630);
xnor U5792 (N_5792,N_5740,N_5732);
or U5793 (N_5793,N_5738,N_5695);
and U5794 (N_5794,N_5702,N_5742);
or U5795 (N_5795,N_5658,N_5656);
nor U5796 (N_5796,N_5744,N_5730);
xnor U5797 (N_5797,N_5701,N_5615);
and U5798 (N_5798,N_5743,N_5666);
nand U5799 (N_5799,N_5604,N_5703);
or U5800 (N_5800,N_5709,N_5613);
or U5801 (N_5801,N_5706,N_5657);
nand U5802 (N_5802,N_5639,N_5631);
nor U5803 (N_5803,N_5651,N_5741);
nor U5804 (N_5804,N_5652,N_5688);
xnor U5805 (N_5805,N_5754,N_5659);
and U5806 (N_5806,N_5636,N_5712);
and U5807 (N_5807,N_5746,N_5602);
and U5808 (N_5808,N_5722,N_5711);
xnor U5809 (N_5809,N_5755,N_5644);
xnor U5810 (N_5810,N_5697,N_5610);
nand U5811 (N_5811,N_5649,N_5734);
xor U5812 (N_5812,N_5745,N_5622);
nand U5813 (N_5813,N_5607,N_5707);
or U5814 (N_5814,N_5747,N_5717);
and U5815 (N_5815,N_5648,N_5671);
xnor U5816 (N_5816,N_5617,N_5689);
and U5817 (N_5817,N_5650,N_5708);
nand U5818 (N_5818,N_5750,N_5611);
xor U5819 (N_5819,N_5679,N_5719);
and U5820 (N_5820,N_5681,N_5661);
and U5821 (N_5821,N_5678,N_5690);
xor U5822 (N_5822,N_5632,N_5687);
nand U5823 (N_5823,N_5721,N_5684);
xnor U5824 (N_5824,N_5608,N_5660);
and U5825 (N_5825,N_5748,N_5674);
xor U5826 (N_5826,N_5729,N_5723);
nor U5827 (N_5827,N_5693,N_5618);
nand U5828 (N_5828,N_5627,N_5694);
and U5829 (N_5829,N_5749,N_5756);
xor U5830 (N_5830,N_5733,N_5676);
xnor U5831 (N_5831,N_5668,N_5714);
nand U5832 (N_5832,N_5641,N_5682);
or U5833 (N_5833,N_5654,N_5705);
and U5834 (N_5834,N_5726,N_5670);
and U5835 (N_5835,N_5724,N_5620);
or U5836 (N_5836,N_5625,N_5713);
nor U5837 (N_5837,N_5623,N_5603);
and U5838 (N_5838,N_5626,N_5720);
xor U5839 (N_5839,N_5646,N_5685);
nand U5840 (N_5840,N_5683,N_5723);
or U5841 (N_5841,N_5640,N_5726);
or U5842 (N_5842,N_5711,N_5651);
nand U5843 (N_5843,N_5623,N_5688);
or U5844 (N_5844,N_5603,N_5721);
nor U5845 (N_5845,N_5733,N_5661);
and U5846 (N_5846,N_5757,N_5654);
and U5847 (N_5847,N_5630,N_5614);
or U5848 (N_5848,N_5610,N_5718);
nand U5849 (N_5849,N_5667,N_5664);
or U5850 (N_5850,N_5690,N_5674);
nand U5851 (N_5851,N_5641,N_5613);
xor U5852 (N_5852,N_5702,N_5724);
nand U5853 (N_5853,N_5694,N_5729);
and U5854 (N_5854,N_5757,N_5733);
or U5855 (N_5855,N_5671,N_5625);
nor U5856 (N_5856,N_5659,N_5732);
nor U5857 (N_5857,N_5720,N_5695);
nor U5858 (N_5858,N_5635,N_5608);
xor U5859 (N_5859,N_5710,N_5623);
or U5860 (N_5860,N_5736,N_5737);
nor U5861 (N_5861,N_5713,N_5716);
and U5862 (N_5862,N_5604,N_5752);
xnor U5863 (N_5863,N_5732,N_5676);
nand U5864 (N_5864,N_5647,N_5639);
nand U5865 (N_5865,N_5671,N_5708);
nand U5866 (N_5866,N_5700,N_5755);
or U5867 (N_5867,N_5636,N_5688);
or U5868 (N_5868,N_5725,N_5758);
xor U5869 (N_5869,N_5669,N_5693);
or U5870 (N_5870,N_5749,N_5715);
nor U5871 (N_5871,N_5684,N_5692);
nor U5872 (N_5872,N_5691,N_5698);
nand U5873 (N_5873,N_5707,N_5619);
or U5874 (N_5874,N_5632,N_5720);
or U5875 (N_5875,N_5703,N_5733);
xnor U5876 (N_5876,N_5639,N_5638);
and U5877 (N_5877,N_5641,N_5752);
and U5878 (N_5878,N_5705,N_5723);
nor U5879 (N_5879,N_5601,N_5611);
nor U5880 (N_5880,N_5712,N_5729);
xor U5881 (N_5881,N_5731,N_5617);
nand U5882 (N_5882,N_5626,N_5692);
nor U5883 (N_5883,N_5712,N_5698);
or U5884 (N_5884,N_5699,N_5610);
xor U5885 (N_5885,N_5687,N_5721);
nor U5886 (N_5886,N_5663,N_5605);
xor U5887 (N_5887,N_5625,N_5698);
xnor U5888 (N_5888,N_5617,N_5725);
nand U5889 (N_5889,N_5692,N_5697);
nand U5890 (N_5890,N_5710,N_5602);
nor U5891 (N_5891,N_5657,N_5640);
or U5892 (N_5892,N_5629,N_5700);
and U5893 (N_5893,N_5707,N_5653);
xor U5894 (N_5894,N_5684,N_5683);
and U5895 (N_5895,N_5703,N_5748);
nor U5896 (N_5896,N_5675,N_5747);
nor U5897 (N_5897,N_5658,N_5650);
xnor U5898 (N_5898,N_5756,N_5696);
or U5899 (N_5899,N_5633,N_5743);
nand U5900 (N_5900,N_5700,N_5627);
nor U5901 (N_5901,N_5664,N_5624);
and U5902 (N_5902,N_5707,N_5665);
or U5903 (N_5903,N_5704,N_5713);
xor U5904 (N_5904,N_5651,N_5759);
nor U5905 (N_5905,N_5711,N_5756);
or U5906 (N_5906,N_5746,N_5614);
xnor U5907 (N_5907,N_5625,N_5646);
nand U5908 (N_5908,N_5644,N_5736);
xnor U5909 (N_5909,N_5686,N_5663);
nand U5910 (N_5910,N_5711,N_5623);
or U5911 (N_5911,N_5713,N_5724);
and U5912 (N_5912,N_5649,N_5684);
nor U5913 (N_5913,N_5709,N_5655);
xnor U5914 (N_5914,N_5734,N_5652);
nor U5915 (N_5915,N_5611,N_5630);
and U5916 (N_5916,N_5619,N_5611);
or U5917 (N_5917,N_5651,N_5683);
nand U5918 (N_5918,N_5638,N_5720);
xnor U5919 (N_5919,N_5621,N_5614);
nor U5920 (N_5920,N_5768,N_5802);
nand U5921 (N_5921,N_5792,N_5809);
nor U5922 (N_5922,N_5899,N_5901);
xnor U5923 (N_5923,N_5827,N_5775);
nor U5924 (N_5924,N_5785,N_5893);
nor U5925 (N_5925,N_5797,N_5877);
or U5926 (N_5926,N_5862,N_5823);
nand U5927 (N_5927,N_5790,N_5833);
nand U5928 (N_5928,N_5867,N_5885);
or U5929 (N_5929,N_5883,N_5819);
nor U5930 (N_5930,N_5892,N_5804);
nor U5931 (N_5931,N_5858,N_5842);
and U5932 (N_5932,N_5845,N_5848);
xor U5933 (N_5933,N_5846,N_5808);
xor U5934 (N_5934,N_5840,N_5830);
or U5935 (N_5935,N_5795,N_5884);
xnor U5936 (N_5936,N_5767,N_5905);
xor U5937 (N_5937,N_5794,N_5838);
nand U5938 (N_5938,N_5839,N_5769);
nor U5939 (N_5939,N_5910,N_5875);
and U5940 (N_5940,N_5816,N_5890);
xnor U5941 (N_5941,N_5817,N_5881);
xor U5942 (N_5942,N_5843,N_5876);
xor U5943 (N_5943,N_5859,N_5865);
and U5944 (N_5944,N_5909,N_5776);
and U5945 (N_5945,N_5900,N_5853);
xnor U5946 (N_5946,N_5878,N_5903);
nand U5947 (N_5947,N_5798,N_5874);
nor U5948 (N_5948,N_5837,N_5762);
nand U5949 (N_5949,N_5908,N_5844);
nand U5950 (N_5950,N_5836,N_5824);
and U5951 (N_5951,N_5780,N_5902);
nor U5952 (N_5952,N_5891,N_5784);
and U5953 (N_5953,N_5799,N_5820);
nand U5954 (N_5954,N_5773,N_5826);
nor U5955 (N_5955,N_5821,N_5871);
and U5956 (N_5956,N_5919,N_5764);
nor U5957 (N_5957,N_5894,N_5860);
xor U5958 (N_5958,N_5806,N_5818);
and U5959 (N_5959,N_5914,N_5872);
xor U5960 (N_5960,N_5814,N_5813);
nand U5961 (N_5961,N_5760,N_5832);
nand U5962 (N_5962,N_5796,N_5800);
or U5963 (N_5963,N_5898,N_5805);
or U5964 (N_5964,N_5783,N_5918);
or U5965 (N_5965,N_5788,N_5801);
and U5966 (N_5966,N_5879,N_5791);
nand U5967 (N_5967,N_5906,N_5774);
and U5968 (N_5968,N_5825,N_5828);
and U5969 (N_5969,N_5831,N_5789);
or U5970 (N_5970,N_5861,N_5811);
nor U5971 (N_5971,N_5772,N_5763);
nand U5972 (N_5972,N_5851,N_5886);
and U5973 (N_5973,N_5904,N_5835);
nand U5974 (N_5974,N_5778,N_5847);
xor U5975 (N_5975,N_5793,N_5766);
xor U5976 (N_5976,N_5761,N_5807);
xnor U5977 (N_5977,N_5770,N_5889);
nand U5978 (N_5978,N_5834,N_5822);
nor U5979 (N_5979,N_5771,N_5787);
nand U5980 (N_5980,N_5896,N_5849);
nand U5981 (N_5981,N_5863,N_5854);
xor U5982 (N_5982,N_5857,N_5781);
or U5983 (N_5983,N_5812,N_5915);
or U5984 (N_5984,N_5868,N_5850);
xor U5985 (N_5985,N_5765,N_5815);
xor U5986 (N_5986,N_5888,N_5897);
xnor U5987 (N_5987,N_5777,N_5856);
and U5988 (N_5988,N_5852,N_5855);
xnor U5989 (N_5989,N_5803,N_5887);
or U5990 (N_5990,N_5917,N_5829);
xor U5991 (N_5991,N_5895,N_5779);
or U5992 (N_5992,N_5864,N_5912);
xor U5993 (N_5993,N_5869,N_5916);
and U5994 (N_5994,N_5841,N_5810);
xnor U5995 (N_5995,N_5907,N_5782);
xnor U5996 (N_5996,N_5882,N_5911);
nand U5997 (N_5997,N_5866,N_5880);
nor U5998 (N_5998,N_5913,N_5870);
xor U5999 (N_5999,N_5786,N_5873);
nand U6000 (N_6000,N_5913,N_5873);
xor U6001 (N_6001,N_5788,N_5824);
and U6002 (N_6002,N_5773,N_5840);
nor U6003 (N_6003,N_5870,N_5773);
or U6004 (N_6004,N_5899,N_5764);
xor U6005 (N_6005,N_5830,N_5815);
and U6006 (N_6006,N_5794,N_5828);
or U6007 (N_6007,N_5846,N_5910);
xnor U6008 (N_6008,N_5908,N_5903);
and U6009 (N_6009,N_5808,N_5815);
and U6010 (N_6010,N_5829,N_5816);
nand U6011 (N_6011,N_5907,N_5814);
nand U6012 (N_6012,N_5761,N_5854);
or U6013 (N_6013,N_5843,N_5896);
nand U6014 (N_6014,N_5846,N_5889);
xnor U6015 (N_6015,N_5792,N_5905);
nand U6016 (N_6016,N_5902,N_5887);
nand U6017 (N_6017,N_5894,N_5880);
nand U6018 (N_6018,N_5823,N_5829);
nor U6019 (N_6019,N_5764,N_5858);
nor U6020 (N_6020,N_5801,N_5802);
nor U6021 (N_6021,N_5824,N_5821);
and U6022 (N_6022,N_5801,N_5765);
nor U6023 (N_6023,N_5857,N_5842);
nand U6024 (N_6024,N_5766,N_5813);
xor U6025 (N_6025,N_5860,N_5805);
nor U6026 (N_6026,N_5784,N_5760);
nor U6027 (N_6027,N_5831,N_5794);
xor U6028 (N_6028,N_5837,N_5841);
and U6029 (N_6029,N_5838,N_5914);
nor U6030 (N_6030,N_5808,N_5798);
nand U6031 (N_6031,N_5774,N_5904);
nor U6032 (N_6032,N_5836,N_5874);
nor U6033 (N_6033,N_5877,N_5871);
xor U6034 (N_6034,N_5822,N_5895);
or U6035 (N_6035,N_5799,N_5767);
and U6036 (N_6036,N_5841,N_5794);
and U6037 (N_6037,N_5812,N_5894);
nor U6038 (N_6038,N_5776,N_5918);
nor U6039 (N_6039,N_5825,N_5896);
or U6040 (N_6040,N_5801,N_5846);
xor U6041 (N_6041,N_5894,N_5817);
nand U6042 (N_6042,N_5844,N_5826);
xor U6043 (N_6043,N_5907,N_5849);
xor U6044 (N_6044,N_5814,N_5852);
nor U6045 (N_6045,N_5827,N_5832);
xnor U6046 (N_6046,N_5789,N_5845);
or U6047 (N_6047,N_5912,N_5853);
and U6048 (N_6048,N_5819,N_5767);
nor U6049 (N_6049,N_5856,N_5898);
nor U6050 (N_6050,N_5918,N_5828);
xnor U6051 (N_6051,N_5869,N_5787);
xor U6052 (N_6052,N_5852,N_5845);
nor U6053 (N_6053,N_5880,N_5911);
xnor U6054 (N_6054,N_5905,N_5907);
or U6055 (N_6055,N_5853,N_5783);
and U6056 (N_6056,N_5891,N_5918);
nor U6057 (N_6057,N_5811,N_5821);
nand U6058 (N_6058,N_5855,N_5910);
or U6059 (N_6059,N_5776,N_5847);
nor U6060 (N_6060,N_5796,N_5872);
or U6061 (N_6061,N_5911,N_5767);
xnor U6062 (N_6062,N_5883,N_5905);
and U6063 (N_6063,N_5825,N_5875);
or U6064 (N_6064,N_5862,N_5803);
xor U6065 (N_6065,N_5791,N_5901);
or U6066 (N_6066,N_5809,N_5770);
nand U6067 (N_6067,N_5883,N_5772);
or U6068 (N_6068,N_5784,N_5826);
xor U6069 (N_6069,N_5865,N_5802);
and U6070 (N_6070,N_5829,N_5801);
xor U6071 (N_6071,N_5892,N_5801);
xor U6072 (N_6072,N_5787,N_5879);
or U6073 (N_6073,N_5823,N_5901);
or U6074 (N_6074,N_5913,N_5899);
and U6075 (N_6075,N_5825,N_5813);
and U6076 (N_6076,N_5896,N_5917);
nor U6077 (N_6077,N_5777,N_5880);
nand U6078 (N_6078,N_5895,N_5894);
nand U6079 (N_6079,N_5775,N_5811);
xor U6080 (N_6080,N_5955,N_5951);
and U6081 (N_6081,N_6052,N_6058);
nor U6082 (N_6082,N_6040,N_5962);
and U6083 (N_6083,N_5943,N_6068);
nor U6084 (N_6084,N_6056,N_6010);
and U6085 (N_6085,N_6023,N_5946);
nor U6086 (N_6086,N_6050,N_6026);
and U6087 (N_6087,N_5971,N_6006);
nor U6088 (N_6088,N_6033,N_5924);
nor U6089 (N_6089,N_5928,N_6008);
and U6090 (N_6090,N_5976,N_5983);
xor U6091 (N_6091,N_5926,N_6045);
nor U6092 (N_6092,N_6012,N_6001);
nor U6093 (N_6093,N_5966,N_5941);
nand U6094 (N_6094,N_6038,N_5985);
or U6095 (N_6095,N_6076,N_5927);
xor U6096 (N_6096,N_6030,N_6054);
and U6097 (N_6097,N_6059,N_6011);
or U6098 (N_6098,N_6061,N_6049);
nor U6099 (N_6099,N_5925,N_6077);
or U6100 (N_6100,N_5932,N_6070);
or U6101 (N_6101,N_6004,N_6073);
nor U6102 (N_6102,N_6002,N_6079);
and U6103 (N_6103,N_6016,N_6018);
and U6104 (N_6104,N_6019,N_5987);
nor U6105 (N_6105,N_5965,N_6032);
or U6106 (N_6106,N_5999,N_5939);
nor U6107 (N_6107,N_6031,N_5997);
xor U6108 (N_6108,N_6041,N_6053);
nand U6109 (N_6109,N_6072,N_5988);
or U6110 (N_6110,N_5996,N_5993);
nor U6111 (N_6111,N_5989,N_6022);
or U6112 (N_6112,N_5934,N_5936);
nor U6113 (N_6113,N_5929,N_5935);
or U6114 (N_6114,N_6048,N_6025);
or U6115 (N_6115,N_5972,N_6024);
or U6116 (N_6116,N_5950,N_5949);
nor U6117 (N_6117,N_6013,N_6034);
xor U6118 (N_6118,N_6028,N_6067);
nand U6119 (N_6119,N_5952,N_6029);
xnor U6120 (N_6120,N_5979,N_5942);
or U6121 (N_6121,N_6044,N_6057);
nand U6122 (N_6122,N_5981,N_5940);
and U6123 (N_6123,N_5954,N_5973);
and U6124 (N_6124,N_5990,N_6003);
and U6125 (N_6125,N_5984,N_6020);
nor U6126 (N_6126,N_5933,N_6039);
nand U6127 (N_6127,N_5931,N_5964);
or U6128 (N_6128,N_5953,N_5995);
nor U6129 (N_6129,N_5994,N_5937);
or U6130 (N_6130,N_5963,N_6046);
nor U6131 (N_6131,N_6074,N_5930);
xor U6132 (N_6132,N_5982,N_5961);
xnor U6133 (N_6133,N_6021,N_5922);
and U6134 (N_6134,N_5977,N_6071);
and U6135 (N_6135,N_5956,N_6007);
nor U6136 (N_6136,N_5921,N_5975);
nand U6137 (N_6137,N_6027,N_6017);
nand U6138 (N_6138,N_6005,N_5970);
nand U6139 (N_6139,N_6037,N_6078);
xnor U6140 (N_6140,N_5938,N_6069);
nor U6141 (N_6141,N_5945,N_5944);
and U6142 (N_6142,N_6060,N_6065);
or U6143 (N_6143,N_5960,N_6047);
xnor U6144 (N_6144,N_6051,N_5947);
xnor U6145 (N_6145,N_6075,N_5974);
or U6146 (N_6146,N_5969,N_6066);
or U6147 (N_6147,N_5967,N_6000);
nor U6148 (N_6148,N_5998,N_6055);
nor U6149 (N_6149,N_5986,N_5957);
xnor U6150 (N_6150,N_6014,N_5980);
xor U6151 (N_6151,N_5978,N_5958);
and U6152 (N_6152,N_6042,N_6035);
xnor U6153 (N_6153,N_6043,N_6063);
or U6154 (N_6154,N_5968,N_5959);
xor U6155 (N_6155,N_5948,N_5923);
nand U6156 (N_6156,N_6015,N_5992);
nand U6157 (N_6157,N_6036,N_5991);
nand U6158 (N_6158,N_6064,N_6009);
xnor U6159 (N_6159,N_5920,N_6062);
or U6160 (N_6160,N_6066,N_5990);
and U6161 (N_6161,N_5960,N_6072);
nand U6162 (N_6162,N_5933,N_6010);
and U6163 (N_6163,N_5948,N_6017);
nand U6164 (N_6164,N_5948,N_5952);
or U6165 (N_6165,N_6046,N_6011);
or U6166 (N_6166,N_6051,N_6072);
xnor U6167 (N_6167,N_5998,N_6010);
or U6168 (N_6168,N_6020,N_5931);
nand U6169 (N_6169,N_6067,N_5937);
xor U6170 (N_6170,N_5990,N_5952);
and U6171 (N_6171,N_6058,N_5932);
xnor U6172 (N_6172,N_6037,N_6023);
or U6173 (N_6173,N_6078,N_6029);
xnor U6174 (N_6174,N_6075,N_5960);
and U6175 (N_6175,N_5974,N_6055);
nand U6176 (N_6176,N_6002,N_5931);
xnor U6177 (N_6177,N_5934,N_6063);
nand U6178 (N_6178,N_5972,N_6017);
nor U6179 (N_6179,N_6051,N_6076);
and U6180 (N_6180,N_6076,N_5978);
nand U6181 (N_6181,N_5928,N_5987);
xnor U6182 (N_6182,N_6001,N_5980);
nand U6183 (N_6183,N_6017,N_5992);
xor U6184 (N_6184,N_5941,N_6009);
xnor U6185 (N_6185,N_5929,N_6070);
xor U6186 (N_6186,N_5944,N_5931);
nor U6187 (N_6187,N_5977,N_5970);
nand U6188 (N_6188,N_5982,N_6039);
or U6189 (N_6189,N_5945,N_5936);
or U6190 (N_6190,N_5922,N_5920);
or U6191 (N_6191,N_6031,N_6066);
and U6192 (N_6192,N_5987,N_5990);
nand U6193 (N_6193,N_6012,N_6020);
xnor U6194 (N_6194,N_6024,N_6040);
xor U6195 (N_6195,N_5994,N_5976);
xnor U6196 (N_6196,N_5969,N_5981);
or U6197 (N_6197,N_6002,N_5994);
nand U6198 (N_6198,N_6001,N_6038);
nand U6199 (N_6199,N_5998,N_6069);
or U6200 (N_6200,N_5939,N_6006);
nor U6201 (N_6201,N_6077,N_5954);
or U6202 (N_6202,N_6027,N_6067);
or U6203 (N_6203,N_5981,N_6066);
and U6204 (N_6204,N_5986,N_5969);
nand U6205 (N_6205,N_6060,N_6004);
nor U6206 (N_6206,N_6038,N_6013);
xor U6207 (N_6207,N_5979,N_5921);
or U6208 (N_6208,N_6069,N_6000);
or U6209 (N_6209,N_6077,N_6079);
nand U6210 (N_6210,N_6030,N_6058);
or U6211 (N_6211,N_5994,N_6010);
nor U6212 (N_6212,N_5988,N_5975);
or U6213 (N_6213,N_5930,N_6068);
xnor U6214 (N_6214,N_5965,N_6067);
xor U6215 (N_6215,N_6019,N_5928);
xnor U6216 (N_6216,N_5959,N_5946);
or U6217 (N_6217,N_6007,N_5921);
or U6218 (N_6218,N_6001,N_5981);
or U6219 (N_6219,N_6072,N_6073);
or U6220 (N_6220,N_6008,N_6014);
nand U6221 (N_6221,N_5968,N_5946);
or U6222 (N_6222,N_6007,N_5965);
nor U6223 (N_6223,N_6037,N_6036);
or U6224 (N_6224,N_5978,N_5936);
nand U6225 (N_6225,N_6065,N_6013);
and U6226 (N_6226,N_6066,N_6034);
or U6227 (N_6227,N_6076,N_6056);
or U6228 (N_6228,N_6034,N_6071);
xor U6229 (N_6229,N_5946,N_6069);
xor U6230 (N_6230,N_5944,N_5957);
nor U6231 (N_6231,N_6067,N_6046);
or U6232 (N_6232,N_5962,N_6024);
and U6233 (N_6233,N_5925,N_5997);
or U6234 (N_6234,N_5943,N_5966);
nor U6235 (N_6235,N_5997,N_6021);
xnor U6236 (N_6236,N_6070,N_5944);
nand U6237 (N_6237,N_6043,N_5983);
xnor U6238 (N_6238,N_6003,N_5969);
nand U6239 (N_6239,N_6016,N_5985);
nor U6240 (N_6240,N_6227,N_6182);
xor U6241 (N_6241,N_6162,N_6123);
nand U6242 (N_6242,N_6088,N_6164);
or U6243 (N_6243,N_6201,N_6193);
nor U6244 (N_6244,N_6122,N_6234);
xor U6245 (N_6245,N_6178,N_6085);
xor U6246 (N_6246,N_6215,N_6149);
nand U6247 (N_6247,N_6140,N_6097);
nor U6248 (N_6248,N_6237,N_6128);
or U6249 (N_6249,N_6161,N_6184);
nor U6250 (N_6250,N_6239,N_6197);
and U6251 (N_6251,N_6146,N_6118);
xor U6252 (N_6252,N_6133,N_6102);
xnor U6253 (N_6253,N_6174,N_6169);
and U6254 (N_6254,N_6176,N_6222);
nor U6255 (N_6255,N_6080,N_6171);
nand U6256 (N_6256,N_6155,N_6132);
and U6257 (N_6257,N_6233,N_6108);
or U6258 (N_6258,N_6094,N_6236);
nor U6259 (N_6259,N_6121,N_6163);
or U6260 (N_6260,N_6101,N_6114);
xor U6261 (N_6261,N_6100,N_6156);
and U6262 (N_6262,N_6189,N_6158);
or U6263 (N_6263,N_6136,N_6130);
and U6264 (N_6264,N_6177,N_6084);
and U6265 (N_6265,N_6205,N_6220);
and U6266 (N_6266,N_6134,N_6127);
xor U6267 (N_6267,N_6148,N_6212);
xnor U6268 (N_6268,N_6141,N_6124);
nor U6269 (N_6269,N_6204,N_6190);
xnor U6270 (N_6270,N_6235,N_6112);
nand U6271 (N_6271,N_6230,N_6159);
xor U6272 (N_6272,N_6172,N_6194);
and U6273 (N_6273,N_6231,N_6086);
nand U6274 (N_6274,N_6083,N_6151);
nor U6275 (N_6275,N_6228,N_6223);
and U6276 (N_6276,N_6091,N_6082);
nand U6277 (N_6277,N_6135,N_6219);
or U6278 (N_6278,N_6131,N_6196);
xnor U6279 (N_6279,N_6166,N_6160);
nor U6280 (N_6280,N_6186,N_6216);
xor U6281 (N_6281,N_6202,N_6126);
nand U6282 (N_6282,N_6217,N_6183);
or U6283 (N_6283,N_6208,N_6081);
nor U6284 (N_6284,N_6116,N_6209);
or U6285 (N_6285,N_6117,N_6211);
nor U6286 (N_6286,N_6206,N_6125);
nor U6287 (N_6287,N_6170,N_6089);
xnor U6288 (N_6288,N_6095,N_6113);
xor U6289 (N_6289,N_6120,N_6092);
nor U6290 (N_6290,N_6185,N_6137);
or U6291 (N_6291,N_6104,N_6099);
nor U6292 (N_6292,N_6105,N_6096);
or U6293 (N_6293,N_6144,N_6213);
and U6294 (N_6294,N_6138,N_6200);
or U6295 (N_6295,N_6181,N_6167);
xnor U6296 (N_6296,N_6152,N_6110);
nor U6297 (N_6297,N_6179,N_6154);
nor U6298 (N_6298,N_6225,N_6107);
and U6299 (N_6299,N_6106,N_6218);
or U6300 (N_6300,N_6168,N_6145);
xor U6301 (N_6301,N_6157,N_6191);
or U6302 (N_6302,N_6198,N_6173);
nand U6303 (N_6303,N_6221,N_6090);
nand U6304 (N_6304,N_6224,N_6232);
xnor U6305 (N_6305,N_6188,N_6226);
nand U6306 (N_6306,N_6153,N_6093);
nor U6307 (N_6307,N_6143,N_6087);
xor U6308 (N_6308,N_6139,N_6192);
xor U6309 (N_6309,N_6129,N_6195);
nand U6310 (N_6310,N_6115,N_6109);
nand U6311 (N_6311,N_6210,N_6103);
nor U6312 (N_6312,N_6098,N_6238);
nand U6313 (N_6313,N_6187,N_6229);
or U6314 (N_6314,N_6111,N_6214);
xnor U6315 (N_6315,N_6150,N_6199);
nand U6316 (N_6316,N_6180,N_6203);
nor U6317 (N_6317,N_6147,N_6165);
xor U6318 (N_6318,N_6207,N_6175);
and U6319 (N_6319,N_6119,N_6142);
or U6320 (N_6320,N_6197,N_6096);
nor U6321 (N_6321,N_6122,N_6132);
xnor U6322 (N_6322,N_6204,N_6237);
xnor U6323 (N_6323,N_6116,N_6099);
nand U6324 (N_6324,N_6216,N_6233);
nand U6325 (N_6325,N_6089,N_6195);
xnor U6326 (N_6326,N_6233,N_6129);
xnor U6327 (N_6327,N_6081,N_6094);
nand U6328 (N_6328,N_6171,N_6115);
nand U6329 (N_6329,N_6143,N_6199);
or U6330 (N_6330,N_6189,N_6200);
nor U6331 (N_6331,N_6194,N_6211);
xor U6332 (N_6332,N_6201,N_6171);
nor U6333 (N_6333,N_6123,N_6170);
xnor U6334 (N_6334,N_6217,N_6221);
or U6335 (N_6335,N_6104,N_6146);
xor U6336 (N_6336,N_6123,N_6177);
or U6337 (N_6337,N_6172,N_6236);
or U6338 (N_6338,N_6113,N_6127);
or U6339 (N_6339,N_6091,N_6086);
nand U6340 (N_6340,N_6146,N_6209);
nor U6341 (N_6341,N_6228,N_6166);
or U6342 (N_6342,N_6147,N_6174);
xor U6343 (N_6343,N_6104,N_6232);
nor U6344 (N_6344,N_6194,N_6200);
or U6345 (N_6345,N_6210,N_6167);
nor U6346 (N_6346,N_6093,N_6167);
nor U6347 (N_6347,N_6096,N_6150);
nand U6348 (N_6348,N_6163,N_6145);
nand U6349 (N_6349,N_6193,N_6191);
nor U6350 (N_6350,N_6234,N_6103);
and U6351 (N_6351,N_6147,N_6227);
and U6352 (N_6352,N_6214,N_6150);
and U6353 (N_6353,N_6213,N_6116);
nor U6354 (N_6354,N_6164,N_6175);
xnor U6355 (N_6355,N_6115,N_6199);
nor U6356 (N_6356,N_6088,N_6178);
nand U6357 (N_6357,N_6110,N_6098);
xnor U6358 (N_6358,N_6224,N_6105);
xor U6359 (N_6359,N_6133,N_6108);
or U6360 (N_6360,N_6194,N_6113);
or U6361 (N_6361,N_6184,N_6194);
nor U6362 (N_6362,N_6237,N_6181);
nor U6363 (N_6363,N_6099,N_6207);
or U6364 (N_6364,N_6162,N_6224);
nand U6365 (N_6365,N_6096,N_6212);
nand U6366 (N_6366,N_6203,N_6122);
nand U6367 (N_6367,N_6162,N_6229);
nor U6368 (N_6368,N_6130,N_6107);
xnor U6369 (N_6369,N_6147,N_6204);
nand U6370 (N_6370,N_6110,N_6190);
or U6371 (N_6371,N_6207,N_6158);
or U6372 (N_6372,N_6225,N_6132);
xor U6373 (N_6373,N_6227,N_6238);
or U6374 (N_6374,N_6089,N_6224);
nor U6375 (N_6375,N_6157,N_6090);
nor U6376 (N_6376,N_6209,N_6151);
xnor U6377 (N_6377,N_6214,N_6229);
and U6378 (N_6378,N_6231,N_6198);
nand U6379 (N_6379,N_6205,N_6158);
nor U6380 (N_6380,N_6124,N_6112);
nor U6381 (N_6381,N_6162,N_6175);
nor U6382 (N_6382,N_6196,N_6092);
nand U6383 (N_6383,N_6192,N_6203);
nor U6384 (N_6384,N_6186,N_6151);
and U6385 (N_6385,N_6107,N_6172);
nand U6386 (N_6386,N_6151,N_6183);
xnor U6387 (N_6387,N_6111,N_6159);
nor U6388 (N_6388,N_6145,N_6157);
and U6389 (N_6389,N_6229,N_6147);
nand U6390 (N_6390,N_6141,N_6151);
xnor U6391 (N_6391,N_6233,N_6170);
or U6392 (N_6392,N_6217,N_6192);
or U6393 (N_6393,N_6164,N_6118);
or U6394 (N_6394,N_6172,N_6186);
and U6395 (N_6395,N_6201,N_6138);
and U6396 (N_6396,N_6220,N_6135);
nor U6397 (N_6397,N_6112,N_6155);
xor U6398 (N_6398,N_6225,N_6102);
nor U6399 (N_6399,N_6144,N_6122);
or U6400 (N_6400,N_6292,N_6248);
and U6401 (N_6401,N_6241,N_6349);
and U6402 (N_6402,N_6270,N_6323);
or U6403 (N_6403,N_6275,N_6330);
or U6404 (N_6404,N_6251,N_6395);
xnor U6405 (N_6405,N_6268,N_6335);
and U6406 (N_6406,N_6358,N_6301);
nand U6407 (N_6407,N_6398,N_6283);
nor U6408 (N_6408,N_6372,N_6286);
nand U6409 (N_6409,N_6346,N_6375);
nor U6410 (N_6410,N_6307,N_6256);
or U6411 (N_6411,N_6336,N_6290);
and U6412 (N_6412,N_6303,N_6363);
xnor U6413 (N_6413,N_6355,N_6388);
or U6414 (N_6414,N_6392,N_6261);
nor U6415 (N_6415,N_6273,N_6353);
or U6416 (N_6416,N_6377,N_6271);
nor U6417 (N_6417,N_6312,N_6337);
and U6418 (N_6418,N_6340,N_6313);
nand U6419 (N_6419,N_6318,N_6352);
xnor U6420 (N_6420,N_6255,N_6245);
xnor U6421 (N_6421,N_6305,N_6317);
xnor U6422 (N_6422,N_6279,N_6396);
nor U6423 (N_6423,N_6378,N_6380);
xor U6424 (N_6424,N_6263,N_6285);
nand U6425 (N_6425,N_6280,N_6276);
or U6426 (N_6426,N_6385,N_6266);
or U6427 (N_6427,N_6287,N_6295);
nor U6428 (N_6428,N_6302,N_6265);
nor U6429 (N_6429,N_6272,N_6397);
nor U6430 (N_6430,N_6343,N_6379);
nand U6431 (N_6431,N_6257,N_6326);
and U6432 (N_6432,N_6274,N_6247);
nand U6433 (N_6433,N_6310,N_6339);
nor U6434 (N_6434,N_6327,N_6364);
xnor U6435 (N_6435,N_6370,N_6382);
nand U6436 (N_6436,N_6365,N_6391);
or U6437 (N_6437,N_6338,N_6291);
or U6438 (N_6438,N_6259,N_6319);
nand U6439 (N_6439,N_6306,N_6240);
and U6440 (N_6440,N_6333,N_6350);
and U6441 (N_6441,N_6399,N_6250);
and U6442 (N_6442,N_6298,N_6309);
or U6443 (N_6443,N_6371,N_6311);
nor U6444 (N_6444,N_6367,N_6374);
and U6445 (N_6445,N_6308,N_6253);
nor U6446 (N_6446,N_6289,N_6389);
nand U6447 (N_6447,N_6341,N_6293);
and U6448 (N_6448,N_6315,N_6356);
xor U6449 (N_6449,N_6277,N_6316);
nor U6450 (N_6450,N_6260,N_6394);
xor U6451 (N_6451,N_6329,N_6386);
or U6452 (N_6452,N_6368,N_6357);
or U6453 (N_6453,N_6332,N_6258);
and U6454 (N_6454,N_6269,N_6296);
nor U6455 (N_6455,N_6383,N_6366);
and U6456 (N_6456,N_6354,N_6242);
nand U6457 (N_6457,N_6376,N_6249);
and U6458 (N_6458,N_6369,N_6267);
nand U6459 (N_6459,N_6254,N_6328);
xnor U6460 (N_6460,N_6322,N_6246);
or U6461 (N_6461,N_6387,N_6297);
xor U6462 (N_6462,N_6345,N_6300);
xnor U6463 (N_6463,N_6331,N_6373);
or U6464 (N_6464,N_6264,N_6320);
xnor U6465 (N_6465,N_6244,N_6252);
nor U6466 (N_6466,N_6284,N_6321);
nand U6467 (N_6467,N_6334,N_6262);
or U6468 (N_6468,N_6360,N_6324);
nor U6469 (N_6469,N_6359,N_6351);
nor U6470 (N_6470,N_6325,N_6384);
or U6471 (N_6471,N_6314,N_6278);
nor U6472 (N_6472,N_6361,N_6381);
nor U6473 (N_6473,N_6243,N_6342);
or U6474 (N_6474,N_6288,N_6362);
or U6475 (N_6475,N_6344,N_6299);
xnor U6476 (N_6476,N_6390,N_6348);
nand U6477 (N_6477,N_6281,N_6282);
xor U6478 (N_6478,N_6304,N_6347);
nand U6479 (N_6479,N_6294,N_6393);
nor U6480 (N_6480,N_6378,N_6360);
xnor U6481 (N_6481,N_6382,N_6257);
nand U6482 (N_6482,N_6248,N_6291);
nor U6483 (N_6483,N_6323,N_6349);
xor U6484 (N_6484,N_6252,N_6270);
nand U6485 (N_6485,N_6355,N_6376);
or U6486 (N_6486,N_6267,N_6248);
nor U6487 (N_6487,N_6279,N_6334);
and U6488 (N_6488,N_6311,N_6355);
nand U6489 (N_6489,N_6357,N_6373);
xnor U6490 (N_6490,N_6335,N_6353);
and U6491 (N_6491,N_6393,N_6285);
nor U6492 (N_6492,N_6376,N_6288);
nand U6493 (N_6493,N_6346,N_6299);
xor U6494 (N_6494,N_6347,N_6321);
xnor U6495 (N_6495,N_6325,N_6304);
xnor U6496 (N_6496,N_6291,N_6303);
and U6497 (N_6497,N_6265,N_6279);
xnor U6498 (N_6498,N_6300,N_6380);
nor U6499 (N_6499,N_6308,N_6248);
nand U6500 (N_6500,N_6253,N_6258);
nand U6501 (N_6501,N_6294,N_6251);
and U6502 (N_6502,N_6368,N_6299);
and U6503 (N_6503,N_6377,N_6287);
and U6504 (N_6504,N_6280,N_6376);
nand U6505 (N_6505,N_6347,N_6286);
nor U6506 (N_6506,N_6376,N_6384);
nand U6507 (N_6507,N_6320,N_6248);
nor U6508 (N_6508,N_6372,N_6295);
and U6509 (N_6509,N_6315,N_6254);
nand U6510 (N_6510,N_6254,N_6293);
nor U6511 (N_6511,N_6333,N_6259);
and U6512 (N_6512,N_6392,N_6292);
nor U6513 (N_6513,N_6351,N_6342);
and U6514 (N_6514,N_6240,N_6352);
and U6515 (N_6515,N_6250,N_6299);
or U6516 (N_6516,N_6302,N_6339);
or U6517 (N_6517,N_6383,N_6340);
xnor U6518 (N_6518,N_6350,N_6345);
nand U6519 (N_6519,N_6361,N_6358);
or U6520 (N_6520,N_6337,N_6340);
nand U6521 (N_6521,N_6264,N_6283);
nor U6522 (N_6522,N_6294,N_6285);
and U6523 (N_6523,N_6349,N_6356);
nand U6524 (N_6524,N_6394,N_6383);
xor U6525 (N_6525,N_6391,N_6287);
nand U6526 (N_6526,N_6371,N_6265);
or U6527 (N_6527,N_6399,N_6372);
and U6528 (N_6528,N_6339,N_6312);
xor U6529 (N_6529,N_6375,N_6366);
or U6530 (N_6530,N_6330,N_6309);
nor U6531 (N_6531,N_6331,N_6304);
or U6532 (N_6532,N_6367,N_6285);
nand U6533 (N_6533,N_6272,N_6367);
or U6534 (N_6534,N_6263,N_6392);
or U6535 (N_6535,N_6373,N_6279);
and U6536 (N_6536,N_6258,N_6263);
and U6537 (N_6537,N_6388,N_6359);
xnor U6538 (N_6538,N_6322,N_6302);
or U6539 (N_6539,N_6306,N_6242);
xnor U6540 (N_6540,N_6320,N_6289);
and U6541 (N_6541,N_6292,N_6369);
or U6542 (N_6542,N_6359,N_6387);
and U6543 (N_6543,N_6379,N_6370);
nand U6544 (N_6544,N_6317,N_6240);
or U6545 (N_6545,N_6293,N_6331);
nand U6546 (N_6546,N_6290,N_6291);
nor U6547 (N_6547,N_6298,N_6339);
nor U6548 (N_6548,N_6344,N_6322);
nor U6549 (N_6549,N_6291,N_6240);
xnor U6550 (N_6550,N_6313,N_6359);
nor U6551 (N_6551,N_6263,N_6394);
or U6552 (N_6552,N_6338,N_6389);
and U6553 (N_6553,N_6255,N_6265);
and U6554 (N_6554,N_6381,N_6244);
xnor U6555 (N_6555,N_6286,N_6345);
and U6556 (N_6556,N_6243,N_6267);
or U6557 (N_6557,N_6289,N_6378);
xor U6558 (N_6558,N_6324,N_6374);
and U6559 (N_6559,N_6242,N_6381);
nor U6560 (N_6560,N_6541,N_6477);
nor U6561 (N_6561,N_6500,N_6425);
or U6562 (N_6562,N_6455,N_6515);
and U6563 (N_6563,N_6441,N_6496);
nand U6564 (N_6564,N_6497,N_6454);
xnor U6565 (N_6565,N_6526,N_6432);
and U6566 (N_6566,N_6486,N_6531);
nor U6567 (N_6567,N_6523,N_6406);
xor U6568 (N_6568,N_6549,N_6545);
and U6569 (N_6569,N_6527,N_6536);
xor U6570 (N_6570,N_6539,N_6411);
or U6571 (N_6571,N_6471,N_6493);
nand U6572 (N_6572,N_6479,N_6473);
nand U6573 (N_6573,N_6439,N_6467);
nand U6574 (N_6574,N_6413,N_6405);
nand U6575 (N_6575,N_6516,N_6459);
xnor U6576 (N_6576,N_6416,N_6519);
or U6577 (N_6577,N_6437,N_6449);
nand U6578 (N_6578,N_6442,N_6468);
nand U6579 (N_6579,N_6457,N_6401);
nor U6580 (N_6580,N_6470,N_6535);
and U6581 (N_6581,N_6420,N_6445);
nor U6582 (N_6582,N_6422,N_6517);
nand U6583 (N_6583,N_6408,N_6458);
nand U6584 (N_6584,N_6498,N_6475);
nand U6585 (N_6585,N_6551,N_6513);
xor U6586 (N_6586,N_6537,N_6407);
xor U6587 (N_6587,N_6469,N_6488);
nand U6588 (N_6588,N_6426,N_6438);
nor U6589 (N_6589,N_6553,N_6460);
nor U6590 (N_6590,N_6522,N_6533);
nor U6591 (N_6591,N_6446,N_6546);
nor U6592 (N_6592,N_6487,N_6521);
and U6593 (N_6593,N_6483,N_6409);
nor U6594 (N_6594,N_6489,N_6421);
xnor U6595 (N_6595,N_6404,N_6538);
or U6596 (N_6596,N_6429,N_6417);
nand U6597 (N_6597,N_6492,N_6532);
or U6598 (N_6598,N_6463,N_6472);
and U6599 (N_6599,N_6554,N_6501);
or U6600 (N_6600,N_6412,N_6507);
xnor U6601 (N_6601,N_6450,N_6414);
and U6602 (N_6602,N_6529,N_6444);
xor U6603 (N_6603,N_6540,N_6547);
xnor U6604 (N_6604,N_6559,N_6552);
or U6605 (N_6605,N_6504,N_6510);
or U6606 (N_6606,N_6506,N_6435);
and U6607 (N_6607,N_6490,N_6402);
or U6608 (N_6608,N_6419,N_6434);
nand U6609 (N_6609,N_6485,N_6528);
nand U6610 (N_6610,N_6474,N_6518);
xor U6611 (N_6611,N_6481,N_6415);
xnor U6612 (N_6612,N_6502,N_6466);
and U6613 (N_6613,N_6555,N_6428);
nand U6614 (N_6614,N_6440,N_6525);
nand U6615 (N_6615,N_6410,N_6512);
nand U6616 (N_6616,N_6558,N_6430);
or U6617 (N_6617,N_6403,N_6509);
or U6618 (N_6618,N_6461,N_6448);
and U6619 (N_6619,N_6436,N_6548);
nor U6620 (N_6620,N_6443,N_6480);
xnor U6621 (N_6621,N_6514,N_6534);
or U6622 (N_6622,N_6433,N_6499);
nand U6623 (N_6623,N_6542,N_6464);
and U6624 (N_6624,N_6556,N_6465);
and U6625 (N_6625,N_6495,N_6508);
nand U6626 (N_6626,N_6462,N_6505);
nor U6627 (N_6627,N_6478,N_6503);
nor U6628 (N_6628,N_6453,N_6494);
xor U6629 (N_6629,N_6550,N_6400);
and U6630 (N_6630,N_6451,N_6530);
nand U6631 (N_6631,N_6524,N_6456);
or U6632 (N_6632,N_6557,N_6543);
xor U6633 (N_6633,N_6427,N_6476);
nand U6634 (N_6634,N_6423,N_6418);
nor U6635 (N_6635,N_6511,N_6452);
xor U6636 (N_6636,N_6424,N_6484);
or U6637 (N_6637,N_6491,N_6447);
xnor U6638 (N_6638,N_6482,N_6520);
or U6639 (N_6639,N_6431,N_6544);
nand U6640 (N_6640,N_6450,N_6514);
xor U6641 (N_6641,N_6486,N_6495);
xnor U6642 (N_6642,N_6553,N_6540);
nand U6643 (N_6643,N_6439,N_6427);
and U6644 (N_6644,N_6452,N_6516);
or U6645 (N_6645,N_6553,N_6551);
xnor U6646 (N_6646,N_6400,N_6423);
nand U6647 (N_6647,N_6557,N_6440);
or U6648 (N_6648,N_6414,N_6559);
or U6649 (N_6649,N_6434,N_6428);
nor U6650 (N_6650,N_6493,N_6552);
xnor U6651 (N_6651,N_6457,N_6484);
or U6652 (N_6652,N_6434,N_6422);
nor U6653 (N_6653,N_6479,N_6423);
and U6654 (N_6654,N_6523,N_6545);
and U6655 (N_6655,N_6539,N_6444);
or U6656 (N_6656,N_6444,N_6550);
nand U6657 (N_6657,N_6443,N_6409);
or U6658 (N_6658,N_6461,N_6557);
or U6659 (N_6659,N_6546,N_6491);
or U6660 (N_6660,N_6527,N_6421);
and U6661 (N_6661,N_6476,N_6542);
nor U6662 (N_6662,N_6413,N_6542);
xor U6663 (N_6663,N_6448,N_6539);
nand U6664 (N_6664,N_6418,N_6554);
or U6665 (N_6665,N_6515,N_6405);
nand U6666 (N_6666,N_6548,N_6541);
xnor U6667 (N_6667,N_6420,N_6535);
and U6668 (N_6668,N_6544,N_6409);
or U6669 (N_6669,N_6422,N_6477);
nand U6670 (N_6670,N_6460,N_6559);
nand U6671 (N_6671,N_6453,N_6465);
and U6672 (N_6672,N_6434,N_6467);
and U6673 (N_6673,N_6467,N_6483);
or U6674 (N_6674,N_6428,N_6499);
and U6675 (N_6675,N_6412,N_6467);
and U6676 (N_6676,N_6496,N_6521);
nor U6677 (N_6677,N_6433,N_6421);
and U6678 (N_6678,N_6409,N_6471);
nand U6679 (N_6679,N_6434,N_6470);
and U6680 (N_6680,N_6478,N_6406);
nand U6681 (N_6681,N_6445,N_6527);
and U6682 (N_6682,N_6448,N_6525);
nor U6683 (N_6683,N_6473,N_6510);
nor U6684 (N_6684,N_6437,N_6451);
and U6685 (N_6685,N_6492,N_6459);
or U6686 (N_6686,N_6463,N_6541);
or U6687 (N_6687,N_6545,N_6426);
xor U6688 (N_6688,N_6528,N_6482);
and U6689 (N_6689,N_6431,N_6401);
and U6690 (N_6690,N_6448,N_6464);
or U6691 (N_6691,N_6504,N_6421);
xnor U6692 (N_6692,N_6514,N_6473);
nand U6693 (N_6693,N_6530,N_6440);
xnor U6694 (N_6694,N_6535,N_6501);
nor U6695 (N_6695,N_6528,N_6493);
and U6696 (N_6696,N_6511,N_6520);
and U6697 (N_6697,N_6419,N_6432);
and U6698 (N_6698,N_6554,N_6512);
and U6699 (N_6699,N_6533,N_6468);
or U6700 (N_6700,N_6505,N_6415);
nor U6701 (N_6701,N_6548,N_6527);
nand U6702 (N_6702,N_6553,N_6427);
xor U6703 (N_6703,N_6423,N_6520);
xnor U6704 (N_6704,N_6558,N_6503);
xor U6705 (N_6705,N_6506,N_6551);
and U6706 (N_6706,N_6510,N_6461);
nand U6707 (N_6707,N_6413,N_6449);
nor U6708 (N_6708,N_6505,N_6453);
nor U6709 (N_6709,N_6404,N_6534);
nand U6710 (N_6710,N_6473,N_6433);
nand U6711 (N_6711,N_6467,N_6535);
xor U6712 (N_6712,N_6465,N_6489);
nor U6713 (N_6713,N_6457,N_6525);
nand U6714 (N_6714,N_6502,N_6406);
xor U6715 (N_6715,N_6430,N_6414);
or U6716 (N_6716,N_6483,N_6459);
xor U6717 (N_6717,N_6509,N_6485);
xnor U6718 (N_6718,N_6443,N_6545);
nor U6719 (N_6719,N_6448,N_6552);
nor U6720 (N_6720,N_6651,N_6610);
or U6721 (N_6721,N_6690,N_6560);
or U6722 (N_6722,N_6619,N_6598);
xor U6723 (N_6723,N_6652,N_6631);
xor U6724 (N_6724,N_6580,N_6707);
nor U6725 (N_6725,N_6679,N_6589);
nor U6726 (N_6726,N_6562,N_6620);
and U6727 (N_6727,N_6622,N_6612);
nor U6728 (N_6728,N_6643,N_6606);
xor U6729 (N_6729,N_6693,N_6570);
or U6730 (N_6730,N_6705,N_6648);
nand U6731 (N_6731,N_6680,N_6624);
nor U6732 (N_6732,N_6710,N_6711);
xnor U6733 (N_6733,N_6607,N_6682);
nor U6734 (N_6734,N_6563,N_6657);
nand U6735 (N_6735,N_6715,N_6568);
or U6736 (N_6736,N_6654,N_6684);
nand U6737 (N_6737,N_6669,N_6655);
nor U6738 (N_6738,N_6592,N_6694);
and U6739 (N_6739,N_6660,N_6681);
nor U6740 (N_6740,N_6659,N_6646);
or U6741 (N_6741,N_6676,N_6617);
nor U6742 (N_6742,N_6675,N_6637);
or U6743 (N_6743,N_6701,N_6674);
and U6744 (N_6744,N_6582,N_6639);
nand U6745 (N_6745,N_6633,N_6621);
nand U6746 (N_6746,N_6644,N_6709);
nor U6747 (N_6747,N_6689,N_6708);
nand U6748 (N_6748,N_6685,N_6702);
xor U6749 (N_6749,N_6583,N_6591);
or U6750 (N_6750,N_6611,N_6665);
or U6751 (N_6751,N_6578,N_6662);
nand U6752 (N_6752,N_6672,N_6603);
or U6753 (N_6753,N_6642,N_6686);
nor U6754 (N_6754,N_6569,N_6590);
and U6755 (N_6755,N_6692,N_6673);
and U6756 (N_6756,N_6634,N_6658);
or U6757 (N_6757,N_6623,N_6601);
and U6758 (N_6758,N_6628,N_6605);
nand U6759 (N_6759,N_6667,N_6584);
nor U6760 (N_6760,N_6666,N_6597);
nor U6761 (N_6761,N_6608,N_6618);
and U6762 (N_6762,N_6627,N_6630);
nand U6763 (N_6763,N_6704,N_6661);
or U6764 (N_6764,N_6700,N_6604);
xor U6765 (N_6765,N_6576,N_6697);
xor U6766 (N_6766,N_6600,N_6585);
nand U6767 (N_6767,N_6577,N_6664);
and U6768 (N_6768,N_6696,N_6688);
nand U6769 (N_6769,N_6645,N_6596);
and U6770 (N_6770,N_6713,N_6615);
nand U6771 (N_6771,N_6641,N_6565);
nor U6772 (N_6772,N_6587,N_6695);
xor U6773 (N_6773,N_6575,N_6714);
nor U6774 (N_6774,N_6586,N_6561);
xor U6775 (N_6775,N_6671,N_6656);
or U6776 (N_6776,N_6566,N_6717);
nor U6777 (N_6777,N_6613,N_6602);
or U6778 (N_6778,N_6635,N_6716);
nor U6779 (N_6779,N_6678,N_6706);
or U6780 (N_6780,N_6670,N_6625);
xor U6781 (N_6781,N_6567,N_6581);
nand U6782 (N_6782,N_6650,N_6588);
nand U6783 (N_6783,N_6698,N_6699);
nand U6784 (N_6784,N_6594,N_6571);
and U6785 (N_6785,N_6595,N_6640);
nand U6786 (N_6786,N_6647,N_6593);
nor U6787 (N_6787,N_6574,N_6599);
nand U6788 (N_6788,N_6638,N_6653);
nor U6789 (N_6789,N_6649,N_6718);
or U6790 (N_6790,N_6683,N_6564);
nor U6791 (N_6791,N_6572,N_6677);
xnor U6792 (N_6792,N_6573,N_6614);
nand U6793 (N_6793,N_6719,N_6663);
nor U6794 (N_6794,N_6609,N_6668);
and U6795 (N_6795,N_6616,N_6712);
nand U6796 (N_6796,N_6629,N_6579);
nor U6797 (N_6797,N_6632,N_6691);
nand U6798 (N_6798,N_6636,N_6703);
nand U6799 (N_6799,N_6687,N_6626);
nor U6800 (N_6800,N_6680,N_6575);
nand U6801 (N_6801,N_6589,N_6660);
nor U6802 (N_6802,N_6662,N_6708);
and U6803 (N_6803,N_6610,N_6647);
or U6804 (N_6804,N_6708,N_6606);
nand U6805 (N_6805,N_6632,N_6716);
nor U6806 (N_6806,N_6658,N_6644);
or U6807 (N_6807,N_6647,N_6561);
xnor U6808 (N_6808,N_6609,N_6638);
nand U6809 (N_6809,N_6703,N_6604);
nor U6810 (N_6810,N_6650,N_6597);
nor U6811 (N_6811,N_6710,N_6650);
or U6812 (N_6812,N_6689,N_6696);
and U6813 (N_6813,N_6701,N_6718);
nand U6814 (N_6814,N_6641,N_6657);
nor U6815 (N_6815,N_6684,N_6705);
nor U6816 (N_6816,N_6582,N_6686);
or U6817 (N_6817,N_6585,N_6664);
or U6818 (N_6818,N_6572,N_6606);
nand U6819 (N_6819,N_6615,N_6569);
nand U6820 (N_6820,N_6652,N_6644);
and U6821 (N_6821,N_6570,N_6631);
nand U6822 (N_6822,N_6592,N_6606);
or U6823 (N_6823,N_6630,N_6684);
xnor U6824 (N_6824,N_6582,N_6588);
xnor U6825 (N_6825,N_6594,N_6634);
nand U6826 (N_6826,N_6570,N_6615);
or U6827 (N_6827,N_6704,N_6678);
nand U6828 (N_6828,N_6706,N_6663);
nand U6829 (N_6829,N_6629,N_6709);
and U6830 (N_6830,N_6673,N_6710);
nand U6831 (N_6831,N_6662,N_6594);
xor U6832 (N_6832,N_6600,N_6706);
nand U6833 (N_6833,N_6640,N_6700);
and U6834 (N_6834,N_6629,N_6580);
and U6835 (N_6835,N_6681,N_6587);
xor U6836 (N_6836,N_6657,N_6594);
nor U6837 (N_6837,N_6622,N_6615);
nor U6838 (N_6838,N_6654,N_6685);
nor U6839 (N_6839,N_6580,N_6593);
or U6840 (N_6840,N_6625,N_6687);
nand U6841 (N_6841,N_6607,N_6663);
nor U6842 (N_6842,N_6631,N_6692);
and U6843 (N_6843,N_6627,N_6602);
and U6844 (N_6844,N_6580,N_6678);
or U6845 (N_6845,N_6679,N_6637);
xor U6846 (N_6846,N_6678,N_6671);
or U6847 (N_6847,N_6691,N_6598);
xnor U6848 (N_6848,N_6657,N_6611);
and U6849 (N_6849,N_6566,N_6715);
nand U6850 (N_6850,N_6632,N_6708);
nor U6851 (N_6851,N_6672,N_6591);
or U6852 (N_6852,N_6561,N_6655);
and U6853 (N_6853,N_6699,N_6642);
or U6854 (N_6854,N_6674,N_6717);
nor U6855 (N_6855,N_6675,N_6655);
nor U6856 (N_6856,N_6661,N_6601);
or U6857 (N_6857,N_6713,N_6574);
xnor U6858 (N_6858,N_6680,N_6698);
nand U6859 (N_6859,N_6670,N_6659);
nand U6860 (N_6860,N_6660,N_6711);
xor U6861 (N_6861,N_6592,N_6593);
or U6862 (N_6862,N_6621,N_6606);
nand U6863 (N_6863,N_6637,N_6648);
and U6864 (N_6864,N_6714,N_6662);
nor U6865 (N_6865,N_6708,N_6690);
or U6866 (N_6866,N_6640,N_6633);
and U6867 (N_6867,N_6608,N_6706);
and U6868 (N_6868,N_6577,N_6605);
xor U6869 (N_6869,N_6639,N_6654);
xnor U6870 (N_6870,N_6578,N_6595);
nor U6871 (N_6871,N_6712,N_6562);
nor U6872 (N_6872,N_6707,N_6693);
and U6873 (N_6873,N_6663,N_6701);
nand U6874 (N_6874,N_6623,N_6616);
and U6875 (N_6875,N_6719,N_6681);
xor U6876 (N_6876,N_6638,N_6642);
and U6877 (N_6877,N_6566,N_6697);
nand U6878 (N_6878,N_6650,N_6594);
and U6879 (N_6879,N_6687,N_6649);
xnor U6880 (N_6880,N_6793,N_6786);
nand U6881 (N_6881,N_6745,N_6775);
nand U6882 (N_6882,N_6773,N_6762);
xor U6883 (N_6883,N_6750,N_6870);
and U6884 (N_6884,N_6831,N_6777);
or U6885 (N_6885,N_6869,N_6739);
or U6886 (N_6886,N_6760,N_6801);
xor U6887 (N_6887,N_6725,N_6764);
or U6888 (N_6888,N_6744,N_6733);
nand U6889 (N_6889,N_6763,N_6844);
nor U6890 (N_6890,N_6868,N_6726);
or U6891 (N_6891,N_6852,N_6808);
nor U6892 (N_6892,N_6840,N_6874);
nand U6893 (N_6893,N_6792,N_6730);
nand U6894 (N_6894,N_6779,N_6778);
nand U6895 (N_6895,N_6794,N_6729);
and U6896 (N_6896,N_6836,N_6823);
xor U6897 (N_6897,N_6765,N_6867);
nand U6898 (N_6898,N_6788,N_6858);
xnor U6899 (N_6899,N_6757,N_6811);
or U6900 (N_6900,N_6720,N_6766);
nor U6901 (N_6901,N_6740,N_6724);
xor U6902 (N_6902,N_6846,N_6842);
xor U6903 (N_6903,N_6721,N_6857);
or U6904 (N_6904,N_6828,N_6803);
nor U6905 (N_6905,N_6837,N_6806);
xnor U6906 (N_6906,N_6848,N_6850);
or U6907 (N_6907,N_6754,N_6865);
or U6908 (N_6908,N_6772,N_6748);
nand U6909 (N_6909,N_6816,N_6818);
or U6910 (N_6910,N_6738,N_6789);
xnor U6911 (N_6911,N_6854,N_6727);
or U6912 (N_6912,N_6761,N_6791);
nand U6913 (N_6913,N_6785,N_6807);
xor U6914 (N_6914,N_6787,N_6735);
nor U6915 (N_6915,N_6847,N_6878);
nor U6916 (N_6916,N_6810,N_6824);
or U6917 (N_6917,N_6841,N_6722);
and U6918 (N_6918,N_6776,N_6835);
or U6919 (N_6919,N_6774,N_6845);
and U6920 (N_6920,N_6876,N_6820);
nor U6921 (N_6921,N_6755,N_6770);
and U6922 (N_6922,N_6822,N_6859);
nor U6923 (N_6923,N_6747,N_6839);
or U6924 (N_6924,N_6734,N_6826);
nand U6925 (N_6925,N_6804,N_6853);
xnor U6926 (N_6926,N_6838,N_6809);
nor U6927 (N_6927,N_6812,N_6814);
nand U6928 (N_6928,N_6872,N_6782);
xor U6929 (N_6929,N_6856,N_6796);
nand U6930 (N_6930,N_6805,N_6742);
nand U6931 (N_6931,N_6759,N_6758);
nand U6932 (N_6932,N_6731,N_6834);
nor U6933 (N_6933,N_6877,N_6784);
or U6934 (N_6934,N_6833,N_6821);
and U6935 (N_6935,N_6795,N_6855);
and U6936 (N_6936,N_6781,N_6780);
or U6937 (N_6937,N_6732,N_6736);
nand U6938 (N_6938,N_6771,N_6843);
or U6939 (N_6939,N_6753,N_6790);
nor U6940 (N_6940,N_6862,N_6863);
and U6941 (N_6941,N_6800,N_6751);
or U6942 (N_6942,N_6827,N_6851);
nor U6943 (N_6943,N_6864,N_6798);
and U6944 (N_6944,N_6866,N_6749);
and U6945 (N_6945,N_6849,N_6873);
xnor U6946 (N_6946,N_6783,N_6768);
nand U6947 (N_6947,N_6832,N_6875);
nor U6948 (N_6948,N_6799,N_6830);
xnor U6949 (N_6949,N_6879,N_6860);
and U6950 (N_6950,N_6825,N_6737);
and U6951 (N_6951,N_6767,N_6819);
or U6952 (N_6952,N_6741,N_6746);
nand U6953 (N_6953,N_6802,N_6817);
and U6954 (N_6954,N_6861,N_6829);
nand U6955 (N_6955,N_6813,N_6797);
nor U6956 (N_6956,N_6728,N_6815);
nor U6957 (N_6957,N_6871,N_6756);
nor U6958 (N_6958,N_6743,N_6752);
nand U6959 (N_6959,N_6723,N_6769);
nor U6960 (N_6960,N_6848,N_6726);
xor U6961 (N_6961,N_6869,N_6853);
nand U6962 (N_6962,N_6834,N_6849);
xor U6963 (N_6963,N_6737,N_6879);
or U6964 (N_6964,N_6782,N_6850);
or U6965 (N_6965,N_6826,N_6755);
or U6966 (N_6966,N_6875,N_6806);
nand U6967 (N_6967,N_6722,N_6856);
xnor U6968 (N_6968,N_6750,N_6751);
nor U6969 (N_6969,N_6862,N_6784);
xor U6970 (N_6970,N_6853,N_6733);
and U6971 (N_6971,N_6785,N_6818);
xor U6972 (N_6972,N_6736,N_6768);
and U6973 (N_6973,N_6748,N_6744);
nand U6974 (N_6974,N_6856,N_6850);
and U6975 (N_6975,N_6854,N_6799);
xnor U6976 (N_6976,N_6834,N_6840);
xnor U6977 (N_6977,N_6804,N_6831);
nand U6978 (N_6978,N_6819,N_6830);
or U6979 (N_6979,N_6845,N_6837);
xnor U6980 (N_6980,N_6876,N_6864);
nand U6981 (N_6981,N_6812,N_6819);
xor U6982 (N_6982,N_6794,N_6745);
xor U6983 (N_6983,N_6851,N_6814);
or U6984 (N_6984,N_6747,N_6745);
and U6985 (N_6985,N_6746,N_6754);
xor U6986 (N_6986,N_6857,N_6807);
nor U6987 (N_6987,N_6798,N_6748);
xor U6988 (N_6988,N_6811,N_6829);
or U6989 (N_6989,N_6862,N_6851);
xnor U6990 (N_6990,N_6725,N_6777);
nor U6991 (N_6991,N_6876,N_6761);
xor U6992 (N_6992,N_6787,N_6866);
xor U6993 (N_6993,N_6856,N_6847);
or U6994 (N_6994,N_6763,N_6732);
nand U6995 (N_6995,N_6785,N_6747);
or U6996 (N_6996,N_6752,N_6770);
xor U6997 (N_6997,N_6834,N_6816);
xnor U6998 (N_6998,N_6776,N_6797);
nand U6999 (N_6999,N_6740,N_6776);
or U7000 (N_7000,N_6781,N_6805);
and U7001 (N_7001,N_6812,N_6740);
or U7002 (N_7002,N_6765,N_6852);
xnor U7003 (N_7003,N_6740,N_6742);
and U7004 (N_7004,N_6767,N_6772);
nor U7005 (N_7005,N_6772,N_6804);
and U7006 (N_7006,N_6819,N_6727);
nand U7007 (N_7007,N_6825,N_6742);
and U7008 (N_7008,N_6802,N_6748);
xnor U7009 (N_7009,N_6860,N_6846);
or U7010 (N_7010,N_6829,N_6826);
nand U7011 (N_7011,N_6841,N_6803);
nor U7012 (N_7012,N_6870,N_6794);
nor U7013 (N_7013,N_6830,N_6796);
nand U7014 (N_7014,N_6811,N_6850);
xor U7015 (N_7015,N_6788,N_6733);
xnor U7016 (N_7016,N_6826,N_6827);
nor U7017 (N_7017,N_6791,N_6834);
xnor U7018 (N_7018,N_6815,N_6851);
xor U7019 (N_7019,N_6788,N_6853);
or U7020 (N_7020,N_6871,N_6831);
nand U7021 (N_7021,N_6809,N_6748);
nand U7022 (N_7022,N_6842,N_6744);
or U7023 (N_7023,N_6723,N_6740);
nand U7024 (N_7024,N_6725,N_6774);
nand U7025 (N_7025,N_6838,N_6759);
or U7026 (N_7026,N_6850,N_6853);
xnor U7027 (N_7027,N_6845,N_6734);
xor U7028 (N_7028,N_6870,N_6843);
and U7029 (N_7029,N_6787,N_6836);
nor U7030 (N_7030,N_6806,N_6734);
xor U7031 (N_7031,N_6733,N_6786);
or U7032 (N_7032,N_6808,N_6749);
or U7033 (N_7033,N_6868,N_6806);
and U7034 (N_7034,N_6875,N_6779);
or U7035 (N_7035,N_6735,N_6726);
nor U7036 (N_7036,N_6780,N_6765);
or U7037 (N_7037,N_6752,N_6814);
xor U7038 (N_7038,N_6866,N_6768);
or U7039 (N_7039,N_6826,N_6819);
or U7040 (N_7040,N_7003,N_6908);
nor U7041 (N_7041,N_6937,N_6980);
and U7042 (N_7042,N_6942,N_6890);
xor U7043 (N_7043,N_6968,N_6921);
or U7044 (N_7044,N_7032,N_6901);
or U7045 (N_7045,N_7025,N_6880);
xnor U7046 (N_7046,N_6907,N_7009);
or U7047 (N_7047,N_6960,N_6931);
or U7048 (N_7048,N_6945,N_7012);
nor U7049 (N_7049,N_6902,N_7002);
nand U7050 (N_7050,N_6930,N_6952);
xor U7051 (N_7051,N_6881,N_7034);
xnor U7052 (N_7052,N_6899,N_7019);
nand U7053 (N_7053,N_7027,N_6894);
and U7054 (N_7054,N_7022,N_6918);
and U7055 (N_7055,N_7004,N_6947);
xor U7056 (N_7056,N_7030,N_7029);
xor U7057 (N_7057,N_7021,N_6974);
and U7058 (N_7058,N_6933,N_7000);
and U7059 (N_7059,N_6976,N_6936);
xnor U7060 (N_7060,N_6944,N_6941);
nor U7061 (N_7061,N_6983,N_6935);
nor U7062 (N_7062,N_6929,N_6950);
or U7063 (N_7063,N_6892,N_7033);
and U7064 (N_7064,N_6926,N_6896);
and U7065 (N_7065,N_6905,N_6897);
nor U7066 (N_7066,N_6955,N_6906);
and U7067 (N_7067,N_6953,N_6991);
or U7068 (N_7068,N_6882,N_7010);
nor U7069 (N_7069,N_6981,N_6964);
xnor U7070 (N_7070,N_6939,N_6971);
nor U7071 (N_7071,N_7011,N_6979);
nand U7072 (N_7072,N_6938,N_6949);
xnor U7073 (N_7073,N_6884,N_6956);
nand U7074 (N_7074,N_6966,N_6987);
or U7075 (N_7075,N_7026,N_6995);
nand U7076 (N_7076,N_6977,N_7039);
nand U7077 (N_7077,N_6969,N_6927);
nand U7078 (N_7078,N_6993,N_7013);
nor U7079 (N_7079,N_6963,N_6948);
nor U7080 (N_7080,N_6885,N_6975);
nand U7081 (N_7081,N_6900,N_6973);
nor U7082 (N_7082,N_6911,N_6920);
or U7083 (N_7083,N_7035,N_6889);
and U7084 (N_7084,N_6916,N_6910);
or U7085 (N_7085,N_6893,N_7017);
or U7086 (N_7086,N_6912,N_6922);
and U7087 (N_7087,N_6886,N_6996);
nor U7088 (N_7088,N_7023,N_6932);
nor U7089 (N_7089,N_6997,N_7007);
or U7090 (N_7090,N_7031,N_6998);
nor U7091 (N_7091,N_6958,N_6957);
and U7092 (N_7092,N_6984,N_6913);
or U7093 (N_7093,N_7024,N_6961);
nor U7094 (N_7094,N_7014,N_7006);
nor U7095 (N_7095,N_6883,N_7038);
and U7096 (N_7096,N_7008,N_6999);
and U7097 (N_7097,N_7020,N_6951);
xor U7098 (N_7098,N_7001,N_6965);
or U7099 (N_7099,N_6986,N_6989);
nand U7100 (N_7100,N_6915,N_7016);
nor U7101 (N_7101,N_6909,N_6954);
and U7102 (N_7102,N_6982,N_6994);
xnor U7103 (N_7103,N_6972,N_6990);
nand U7104 (N_7104,N_6923,N_6940);
nand U7105 (N_7105,N_6891,N_7028);
nor U7106 (N_7106,N_6928,N_6904);
or U7107 (N_7107,N_6925,N_7015);
nor U7108 (N_7108,N_6903,N_6967);
xnor U7109 (N_7109,N_7005,N_6970);
nand U7110 (N_7110,N_6985,N_6959);
nor U7111 (N_7111,N_6962,N_6898);
nor U7112 (N_7112,N_6978,N_6917);
or U7113 (N_7113,N_6919,N_6914);
nand U7114 (N_7114,N_6895,N_6934);
nand U7115 (N_7115,N_7018,N_6992);
nor U7116 (N_7116,N_6887,N_7036);
xor U7117 (N_7117,N_6924,N_6946);
nand U7118 (N_7118,N_7037,N_6943);
xor U7119 (N_7119,N_6888,N_6988);
nand U7120 (N_7120,N_6915,N_6993);
nand U7121 (N_7121,N_6987,N_6898);
nand U7122 (N_7122,N_6955,N_6978);
xnor U7123 (N_7123,N_6967,N_6984);
or U7124 (N_7124,N_6907,N_6990);
xnor U7125 (N_7125,N_6899,N_6914);
xnor U7126 (N_7126,N_7034,N_7009);
nor U7127 (N_7127,N_7020,N_6905);
and U7128 (N_7128,N_6976,N_6985);
xor U7129 (N_7129,N_6882,N_6889);
and U7130 (N_7130,N_6904,N_6906);
and U7131 (N_7131,N_6950,N_6888);
xor U7132 (N_7132,N_6990,N_6889);
nor U7133 (N_7133,N_6926,N_6882);
and U7134 (N_7134,N_6943,N_6995);
nand U7135 (N_7135,N_6934,N_6933);
or U7136 (N_7136,N_6961,N_6890);
nand U7137 (N_7137,N_6956,N_6930);
xnor U7138 (N_7138,N_6928,N_6958);
and U7139 (N_7139,N_7030,N_6957);
nor U7140 (N_7140,N_6950,N_6967);
nand U7141 (N_7141,N_7003,N_7013);
or U7142 (N_7142,N_7001,N_6939);
nor U7143 (N_7143,N_6942,N_6917);
xor U7144 (N_7144,N_6924,N_6966);
nand U7145 (N_7145,N_6925,N_7011);
nand U7146 (N_7146,N_7018,N_6945);
and U7147 (N_7147,N_7033,N_7005);
and U7148 (N_7148,N_6908,N_6900);
nor U7149 (N_7149,N_6972,N_6970);
nand U7150 (N_7150,N_6894,N_6952);
and U7151 (N_7151,N_6939,N_6927);
and U7152 (N_7152,N_6969,N_6967);
xor U7153 (N_7153,N_7032,N_7031);
and U7154 (N_7154,N_6912,N_7007);
and U7155 (N_7155,N_6991,N_6936);
xnor U7156 (N_7156,N_7023,N_7005);
and U7157 (N_7157,N_7034,N_6979);
or U7158 (N_7158,N_6885,N_7015);
or U7159 (N_7159,N_6896,N_6912);
or U7160 (N_7160,N_6960,N_6979);
and U7161 (N_7161,N_6914,N_6944);
and U7162 (N_7162,N_7027,N_6944);
and U7163 (N_7163,N_6987,N_6884);
nand U7164 (N_7164,N_6955,N_6884);
nor U7165 (N_7165,N_6903,N_6891);
and U7166 (N_7166,N_6911,N_6965);
xnor U7167 (N_7167,N_7028,N_6915);
and U7168 (N_7168,N_7011,N_6943);
nor U7169 (N_7169,N_6912,N_6916);
and U7170 (N_7170,N_7007,N_6926);
or U7171 (N_7171,N_6991,N_6886);
nor U7172 (N_7172,N_6950,N_6961);
or U7173 (N_7173,N_6980,N_6963);
or U7174 (N_7174,N_6987,N_6926);
nand U7175 (N_7175,N_7011,N_7005);
and U7176 (N_7176,N_6894,N_6993);
nand U7177 (N_7177,N_6985,N_6978);
nand U7178 (N_7178,N_6943,N_6960);
nor U7179 (N_7179,N_6983,N_6916);
or U7180 (N_7180,N_6892,N_6924);
nor U7181 (N_7181,N_7037,N_6979);
nor U7182 (N_7182,N_6973,N_7010);
and U7183 (N_7183,N_6964,N_7023);
and U7184 (N_7184,N_6915,N_6955);
or U7185 (N_7185,N_6957,N_7026);
nor U7186 (N_7186,N_6958,N_6954);
xnor U7187 (N_7187,N_6946,N_6972);
and U7188 (N_7188,N_6988,N_7013);
nor U7189 (N_7189,N_6962,N_7036);
and U7190 (N_7190,N_6957,N_7020);
and U7191 (N_7191,N_6939,N_6883);
nor U7192 (N_7192,N_6951,N_6979);
xnor U7193 (N_7193,N_6991,N_6961);
and U7194 (N_7194,N_6881,N_7007);
or U7195 (N_7195,N_7018,N_6959);
nor U7196 (N_7196,N_7024,N_6962);
or U7197 (N_7197,N_6941,N_6982);
or U7198 (N_7198,N_6976,N_6961);
nand U7199 (N_7199,N_7016,N_7019);
nor U7200 (N_7200,N_7122,N_7055);
and U7201 (N_7201,N_7194,N_7123);
nor U7202 (N_7202,N_7114,N_7131);
or U7203 (N_7203,N_7191,N_7116);
xor U7204 (N_7204,N_7048,N_7109);
and U7205 (N_7205,N_7184,N_7059);
nand U7206 (N_7206,N_7119,N_7105);
nor U7207 (N_7207,N_7172,N_7046);
nor U7208 (N_7208,N_7087,N_7101);
nor U7209 (N_7209,N_7064,N_7052);
xnor U7210 (N_7210,N_7077,N_7042);
nand U7211 (N_7211,N_7189,N_7082);
nand U7212 (N_7212,N_7186,N_7090);
and U7213 (N_7213,N_7112,N_7089);
xor U7214 (N_7214,N_7060,N_7148);
xnor U7215 (N_7215,N_7085,N_7056);
and U7216 (N_7216,N_7076,N_7110);
nor U7217 (N_7217,N_7185,N_7115);
nor U7218 (N_7218,N_7104,N_7153);
or U7219 (N_7219,N_7138,N_7049);
nand U7220 (N_7220,N_7080,N_7107);
nor U7221 (N_7221,N_7066,N_7074);
and U7222 (N_7222,N_7111,N_7069);
or U7223 (N_7223,N_7192,N_7041);
or U7224 (N_7224,N_7062,N_7158);
or U7225 (N_7225,N_7054,N_7171);
nand U7226 (N_7226,N_7176,N_7100);
nor U7227 (N_7227,N_7043,N_7120);
nor U7228 (N_7228,N_7108,N_7098);
or U7229 (N_7229,N_7146,N_7167);
nand U7230 (N_7230,N_7198,N_7195);
nor U7231 (N_7231,N_7163,N_7168);
xor U7232 (N_7232,N_7129,N_7099);
nand U7233 (N_7233,N_7175,N_7177);
xnor U7234 (N_7234,N_7067,N_7045);
xor U7235 (N_7235,N_7174,N_7065);
xnor U7236 (N_7236,N_7150,N_7161);
nand U7237 (N_7237,N_7199,N_7160);
nand U7238 (N_7238,N_7050,N_7144);
nor U7239 (N_7239,N_7078,N_7196);
xor U7240 (N_7240,N_7127,N_7187);
xor U7241 (N_7241,N_7061,N_7128);
xnor U7242 (N_7242,N_7140,N_7121);
xor U7243 (N_7243,N_7102,N_7134);
nand U7244 (N_7244,N_7135,N_7094);
xnor U7245 (N_7245,N_7143,N_7070);
xnor U7246 (N_7246,N_7159,N_7132);
xnor U7247 (N_7247,N_7149,N_7040);
nand U7248 (N_7248,N_7145,N_7180);
nor U7249 (N_7249,N_7178,N_7051);
xnor U7250 (N_7250,N_7133,N_7157);
nand U7251 (N_7251,N_7079,N_7124);
and U7252 (N_7252,N_7139,N_7164);
and U7253 (N_7253,N_7165,N_7068);
or U7254 (N_7254,N_7063,N_7097);
xor U7255 (N_7255,N_7142,N_7173);
and U7256 (N_7256,N_7117,N_7181);
and U7257 (N_7257,N_7147,N_7183);
and U7258 (N_7258,N_7091,N_7095);
xor U7259 (N_7259,N_7169,N_7086);
xnor U7260 (N_7260,N_7081,N_7058);
nor U7261 (N_7261,N_7096,N_7125);
nor U7262 (N_7262,N_7103,N_7136);
or U7263 (N_7263,N_7152,N_7044);
or U7264 (N_7264,N_7154,N_7071);
or U7265 (N_7265,N_7151,N_7156);
nand U7266 (N_7266,N_7126,N_7083);
nor U7267 (N_7267,N_7106,N_7162);
nor U7268 (N_7268,N_7084,N_7088);
nand U7269 (N_7269,N_7130,N_7047);
or U7270 (N_7270,N_7118,N_7137);
nor U7271 (N_7271,N_7188,N_7093);
xnor U7272 (N_7272,N_7141,N_7053);
xor U7273 (N_7273,N_7155,N_7073);
nand U7274 (N_7274,N_7072,N_7092);
or U7275 (N_7275,N_7113,N_7190);
xnor U7276 (N_7276,N_7193,N_7179);
or U7277 (N_7277,N_7057,N_7182);
xnor U7278 (N_7278,N_7197,N_7075);
nor U7279 (N_7279,N_7166,N_7170);
or U7280 (N_7280,N_7120,N_7119);
and U7281 (N_7281,N_7174,N_7194);
and U7282 (N_7282,N_7059,N_7139);
nand U7283 (N_7283,N_7151,N_7159);
or U7284 (N_7284,N_7071,N_7174);
nand U7285 (N_7285,N_7076,N_7147);
nor U7286 (N_7286,N_7124,N_7108);
and U7287 (N_7287,N_7174,N_7045);
and U7288 (N_7288,N_7055,N_7051);
and U7289 (N_7289,N_7051,N_7058);
or U7290 (N_7290,N_7048,N_7150);
nor U7291 (N_7291,N_7072,N_7051);
nor U7292 (N_7292,N_7092,N_7145);
nor U7293 (N_7293,N_7173,N_7082);
nand U7294 (N_7294,N_7106,N_7152);
nor U7295 (N_7295,N_7153,N_7140);
or U7296 (N_7296,N_7095,N_7074);
or U7297 (N_7297,N_7111,N_7044);
nand U7298 (N_7298,N_7110,N_7119);
xor U7299 (N_7299,N_7075,N_7094);
nor U7300 (N_7300,N_7130,N_7132);
or U7301 (N_7301,N_7170,N_7103);
nand U7302 (N_7302,N_7178,N_7055);
xnor U7303 (N_7303,N_7146,N_7124);
xnor U7304 (N_7304,N_7078,N_7136);
nand U7305 (N_7305,N_7098,N_7141);
xor U7306 (N_7306,N_7100,N_7131);
or U7307 (N_7307,N_7108,N_7139);
and U7308 (N_7308,N_7105,N_7133);
xor U7309 (N_7309,N_7143,N_7087);
and U7310 (N_7310,N_7179,N_7199);
nor U7311 (N_7311,N_7078,N_7055);
nor U7312 (N_7312,N_7186,N_7068);
nor U7313 (N_7313,N_7114,N_7090);
or U7314 (N_7314,N_7053,N_7066);
nor U7315 (N_7315,N_7106,N_7177);
and U7316 (N_7316,N_7108,N_7114);
nor U7317 (N_7317,N_7089,N_7059);
or U7318 (N_7318,N_7174,N_7048);
xnor U7319 (N_7319,N_7092,N_7077);
xnor U7320 (N_7320,N_7137,N_7074);
nand U7321 (N_7321,N_7148,N_7053);
and U7322 (N_7322,N_7076,N_7193);
nand U7323 (N_7323,N_7057,N_7124);
nand U7324 (N_7324,N_7149,N_7176);
and U7325 (N_7325,N_7071,N_7088);
nand U7326 (N_7326,N_7181,N_7199);
nand U7327 (N_7327,N_7082,N_7073);
xor U7328 (N_7328,N_7117,N_7092);
and U7329 (N_7329,N_7186,N_7081);
nand U7330 (N_7330,N_7106,N_7076);
and U7331 (N_7331,N_7089,N_7049);
nand U7332 (N_7332,N_7194,N_7095);
and U7333 (N_7333,N_7122,N_7125);
xnor U7334 (N_7334,N_7194,N_7157);
nand U7335 (N_7335,N_7172,N_7049);
or U7336 (N_7336,N_7088,N_7074);
nor U7337 (N_7337,N_7149,N_7066);
and U7338 (N_7338,N_7119,N_7040);
xnor U7339 (N_7339,N_7192,N_7098);
xnor U7340 (N_7340,N_7070,N_7074);
xnor U7341 (N_7341,N_7193,N_7128);
or U7342 (N_7342,N_7074,N_7082);
xor U7343 (N_7343,N_7134,N_7116);
and U7344 (N_7344,N_7088,N_7123);
and U7345 (N_7345,N_7159,N_7121);
nand U7346 (N_7346,N_7106,N_7073);
or U7347 (N_7347,N_7057,N_7127);
and U7348 (N_7348,N_7174,N_7120);
xnor U7349 (N_7349,N_7058,N_7066);
xor U7350 (N_7350,N_7132,N_7114);
and U7351 (N_7351,N_7134,N_7155);
and U7352 (N_7352,N_7168,N_7106);
nor U7353 (N_7353,N_7186,N_7099);
nor U7354 (N_7354,N_7045,N_7079);
and U7355 (N_7355,N_7084,N_7198);
nor U7356 (N_7356,N_7081,N_7181);
nand U7357 (N_7357,N_7182,N_7195);
nand U7358 (N_7358,N_7105,N_7076);
and U7359 (N_7359,N_7158,N_7135);
nand U7360 (N_7360,N_7244,N_7337);
nor U7361 (N_7361,N_7330,N_7271);
and U7362 (N_7362,N_7237,N_7257);
xor U7363 (N_7363,N_7218,N_7333);
or U7364 (N_7364,N_7304,N_7207);
xnor U7365 (N_7365,N_7281,N_7262);
xnor U7366 (N_7366,N_7354,N_7352);
nor U7367 (N_7367,N_7270,N_7239);
or U7368 (N_7368,N_7228,N_7291);
xor U7369 (N_7369,N_7280,N_7320);
nand U7370 (N_7370,N_7314,N_7263);
nand U7371 (N_7371,N_7276,N_7305);
or U7372 (N_7372,N_7356,N_7222);
nor U7373 (N_7373,N_7254,N_7290);
or U7374 (N_7374,N_7203,N_7250);
xnor U7375 (N_7375,N_7231,N_7349);
nand U7376 (N_7376,N_7308,N_7296);
nand U7377 (N_7377,N_7329,N_7358);
and U7378 (N_7378,N_7325,N_7359);
nor U7379 (N_7379,N_7230,N_7242);
or U7380 (N_7380,N_7260,N_7233);
xor U7381 (N_7381,N_7248,N_7241);
nand U7382 (N_7382,N_7220,N_7215);
nand U7383 (N_7383,N_7286,N_7229);
nand U7384 (N_7384,N_7326,N_7216);
or U7385 (N_7385,N_7210,N_7315);
nor U7386 (N_7386,N_7346,N_7264);
xor U7387 (N_7387,N_7219,N_7297);
or U7388 (N_7388,N_7341,N_7251);
nand U7389 (N_7389,N_7221,N_7313);
nand U7390 (N_7390,N_7284,N_7268);
nand U7391 (N_7391,N_7336,N_7294);
xnor U7392 (N_7392,N_7345,N_7278);
nand U7393 (N_7393,N_7307,N_7225);
nand U7394 (N_7394,N_7328,N_7211);
and U7395 (N_7395,N_7288,N_7299);
nor U7396 (N_7396,N_7316,N_7338);
nand U7397 (N_7397,N_7240,N_7351);
or U7398 (N_7398,N_7298,N_7217);
or U7399 (N_7399,N_7253,N_7277);
xnor U7400 (N_7400,N_7234,N_7310);
xnor U7401 (N_7401,N_7283,N_7223);
or U7402 (N_7402,N_7355,N_7292);
nor U7403 (N_7403,N_7334,N_7312);
nand U7404 (N_7404,N_7332,N_7342);
or U7405 (N_7405,N_7272,N_7266);
or U7406 (N_7406,N_7212,N_7256);
and U7407 (N_7407,N_7214,N_7347);
or U7408 (N_7408,N_7335,N_7331);
nand U7409 (N_7409,N_7300,N_7340);
nand U7410 (N_7410,N_7285,N_7238);
nor U7411 (N_7411,N_7261,N_7255);
nor U7412 (N_7412,N_7321,N_7259);
and U7413 (N_7413,N_7279,N_7323);
nor U7414 (N_7414,N_7311,N_7213);
nor U7415 (N_7415,N_7350,N_7243);
or U7416 (N_7416,N_7227,N_7327);
or U7417 (N_7417,N_7324,N_7204);
nand U7418 (N_7418,N_7319,N_7232);
nand U7419 (N_7419,N_7202,N_7200);
or U7420 (N_7420,N_7209,N_7309);
or U7421 (N_7421,N_7306,N_7275);
nor U7422 (N_7422,N_7293,N_7303);
nor U7423 (N_7423,N_7201,N_7357);
and U7424 (N_7424,N_7205,N_7282);
nor U7425 (N_7425,N_7226,N_7317);
nand U7426 (N_7426,N_7235,N_7343);
nand U7427 (N_7427,N_7249,N_7274);
and U7428 (N_7428,N_7295,N_7247);
nand U7429 (N_7429,N_7267,N_7302);
nor U7430 (N_7430,N_7289,N_7344);
nand U7431 (N_7431,N_7252,N_7206);
xnor U7432 (N_7432,N_7287,N_7208);
or U7433 (N_7433,N_7258,N_7236);
nand U7434 (N_7434,N_7246,N_7339);
nor U7435 (N_7435,N_7265,N_7348);
and U7436 (N_7436,N_7245,N_7353);
or U7437 (N_7437,N_7318,N_7269);
nor U7438 (N_7438,N_7224,N_7301);
nand U7439 (N_7439,N_7322,N_7273);
or U7440 (N_7440,N_7339,N_7304);
or U7441 (N_7441,N_7303,N_7240);
and U7442 (N_7442,N_7203,N_7205);
or U7443 (N_7443,N_7222,N_7232);
and U7444 (N_7444,N_7253,N_7288);
or U7445 (N_7445,N_7297,N_7238);
or U7446 (N_7446,N_7220,N_7228);
or U7447 (N_7447,N_7306,N_7331);
nor U7448 (N_7448,N_7291,N_7284);
and U7449 (N_7449,N_7287,N_7315);
or U7450 (N_7450,N_7275,N_7270);
or U7451 (N_7451,N_7207,N_7335);
or U7452 (N_7452,N_7217,N_7358);
and U7453 (N_7453,N_7246,N_7232);
nand U7454 (N_7454,N_7327,N_7204);
or U7455 (N_7455,N_7271,N_7287);
and U7456 (N_7456,N_7212,N_7341);
or U7457 (N_7457,N_7309,N_7271);
or U7458 (N_7458,N_7222,N_7332);
or U7459 (N_7459,N_7342,N_7274);
or U7460 (N_7460,N_7335,N_7200);
nor U7461 (N_7461,N_7256,N_7219);
and U7462 (N_7462,N_7309,N_7202);
nor U7463 (N_7463,N_7323,N_7247);
and U7464 (N_7464,N_7322,N_7336);
nand U7465 (N_7465,N_7206,N_7319);
xor U7466 (N_7466,N_7266,N_7323);
and U7467 (N_7467,N_7297,N_7338);
nor U7468 (N_7468,N_7296,N_7289);
xnor U7469 (N_7469,N_7358,N_7234);
and U7470 (N_7470,N_7204,N_7209);
and U7471 (N_7471,N_7231,N_7303);
xnor U7472 (N_7472,N_7272,N_7284);
nor U7473 (N_7473,N_7303,N_7346);
and U7474 (N_7474,N_7333,N_7287);
xor U7475 (N_7475,N_7242,N_7337);
nand U7476 (N_7476,N_7228,N_7354);
nand U7477 (N_7477,N_7254,N_7312);
and U7478 (N_7478,N_7262,N_7220);
and U7479 (N_7479,N_7227,N_7237);
nand U7480 (N_7480,N_7320,N_7249);
and U7481 (N_7481,N_7295,N_7339);
or U7482 (N_7482,N_7358,N_7281);
xnor U7483 (N_7483,N_7238,N_7314);
nand U7484 (N_7484,N_7334,N_7343);
nor U7485 (N_7485,N_7269,N_7228);
xor U7486 (N_7486,N_7346,N_7251);
xnor U7487 (N_7487,N_7265,N_7275);
or U7488 (N_7488,N_7237,N_7236);
or U7489 (N_7489,N_7255,N_7301);
or U7490 (N_7490,N_7266,N_7203);
nor U7491 (N_7491,N_7259,N_7350);
nand U7492 (N_7492,N_7307,N_7322);
nand U7493 (N_7493,N_7263,N_7306);
xnor U7494 (N_7494,N_7339,N_7356);
xor U7495 (N_7495,N_7301,N_7240);
or U7496 (N_7496,N_7293,N_7227);
and U7497 (N_7497,N_7329,N_7317);
nand U7498 (N_7498,N_7348,N_7333);
nor U7499 (N_7499,N_7269,N_7328);
xnor U7500 (N_7500,N_7302,N_7321);
and U7501 (N_7501,N_7270,N_7204);
or U7502 (N_7502,N_7226,N_7316);
xor U7503 (N_7503,N_7228,N_7329);
and U7504 (N_7504,N_7235,N_7304);
or U7505 (N_7505,N_7345,N_7348);
nor U7506 (N_7506,N_7330,N_7334);
and U7507 (N_7507,N_7302,N_7210);
nor U7508 (N_7508,N_7299,N_7258);
xor U7509 (N_7509,N_7290,N_7344);
nor U7510 (N_7510,N_7267,N_7261);
nand U7511 (N_7511,N_7206,N_7239);
or U7512 (N_7512,N_7300,N_7332);
and U7513 (N_7513,N_7325,N_7241);
and U7514 (N_7514,N_7211,N_7264);
and U7515 (N_7515,N_7205,N_7290);
xnor U7516 (N_7516,N_7337,N_7319);
and U7517 (N_7517,N_7295,N_7304);
xnor U7518 (N_7518,N_7208,N_7207);
nand U7519 (N_7519,N_7300,N_7270);
xor U7520 (N_7520,N_7377,N_7493);
nor U7521 (N_7521,N_7458,N_7488);
nand U7522 (N_7522,N_7470,N_7403);
and U7523 (N_7523,N_7506,N_7468);
xor U7524 (N_7524,N_7417,N_7497);
nor U7525 (N_7525,N_7504,N_7391);
nor U7526 (N_7526,N_7370,N_7467);
and U7527 (N_7527,N_7379,N_7412);
and U7528 (N_7528,N_7371,N_7369);
nand U7529 (N_7529,N_7519,N_7374);
and U7530 (N_7530,N_7446,N_7515);
nor U7531 (N_7531,N_7409,N_7388);
and U7532 (N_7532,N_7384,N_7436);
xnor U7533 (N_7533,N_7413,N_7380);
or U7534 (N_7534,N_7435,N_7418);
xor U7535 (N_7535,N_7411,N_7381);
and U7536 (N_7536,N_7494,N_7364);
nor U7537 (N_7537,N_7396,N_7472);
and U7538 (N_7538,N_7410,N_7429);
and U7539 (N_7539,N_7444,N_7518);
and U7540 (N_7540,N_7441,N_7485);
nand U7541 (N_7541,N_7492,N_7390);
or U7542 (N_7542,N_7462,N_7438);
xnor U7543 (N_7543,N_7376,N_7400);
nor U7544 (N_7544,N_7496,N_7419);
xnor U7545 (N_7545,N_7430,N_7471);
nor U7546 (N_7546,N_7510,N_7466);
xor U7547 (N_7547,N_7461,N_7484);
nor U7548 (N_7548,N_7363,N_7407);
nor U7549 (N_7549,N_7425,N_7427);
and U7550 (N_7550,N_7439,N_7476);
xor U7551 (N_7551,N_7431,N_7422);
nor U7552 (N_7552,N_7480,N_7426);
xnor U7553 (N_7553,N_7455,N_7509);
nor U7554 (N_7554,N_7420,N_7508);
or U7555 (N_7555,N_7464,N_7399);
nand U7556 (N_7556,N_7449,N_7448);
or U7557 (N_7557,N_7360,N_7482);
nor U7558 (N_7558,N_7502,N_7372);
nor U7559 (N_7559,N_7428,N_7490);
nor U7560 (N_7560,N_7405,N_7454);
nor U7561 (N_7561,N_7404,N_7451);
or U7562 (N_7562,N_7511,N_7406);
nand U7563 (N_7563,N_7491,N_7478);
nor U7564 (N_7564,N_7362,N_7477);
nor U7565 (N_7565,N_7495,N_7456);
xor U7566 (N_7566,N_7487,N_7463);
nor U7567 (N_7567,N_7445,N_7474);
xor U7568 (N_7568,N_7483,N_7366);
xor U7569 (N_7569,N_7473,N_7397);
nor U7570 (N_7570,N_7516,N_7416);
nor U7571 (N_7571,N_7513,N_7424);
or U7572 (N_7572,N_7401,N_7378);
nor U7573 (N_7573,N_7465,N_7368);
xor U7574 (N_7574,N_7434,N_7361);
and U7575 (N_7575,N_7386,N_7500);
and U7576 (N_7576,N_7489,N_7389);
nor U7577 (N_7577,N_7442,N_7393);
xnor U7578 (N_7578,N_7382,N_7453);
nand U7579 (N_7579,N_7479,N_7395);
and U7580 (N_7580,N_7501,N_7433);
xor U7581 (N_7581,N_7392,N_7459);
and U7582 (N_7582,N_7514,N_7437);
nor U7583 (N_7583,N_7503,N_7394);
nand U7584 (N_7584,N_7517,N_7408);
nand U7585 (N_7585,N_7365,N_7443);
nor U7586 (N_7586,N_7414,N_7447);
or U7587 (N_7587,N_7452,N_7421);
or U7588 (N_7588,N_7373,N_7383);
nor U7589 (N_7589,N_7398,N_7415);
nor U7590 (N_7590,N_7423,N_7460);
or U7591 (N_7591,N_7507,N_7450);
nor U7592 (N_7592,N_7469,N_7457);
xnor U7593 (N_7593,N_7498,N_7481);
xor U7594 (N_7594,N_7367,N_7486);
nand U7595 (N_7595,N_7432,N_7499);
and U7596 (N_7596,N_7385,N_7505);
nand U7597 (N_7597,N_7387,N_7440);
or U7598 (N_7598,N_7475,N_7512);
xor U7599 (N_7599,N_7375,N_7402);
nor U7600 (N_7600,N_7424,N_7372);
or U7601 (N_7601,N_7519,N_7422);
or U7602 (N_7602,N_7511,N_7438);
xnor U7603 (N_7603,N_7512,N_7435);
or U7604 (N_7604,N_7373,N_7403);
or U7605 (N_7605,N_7421,N_7469);
and U7606 (N_7606,N_7365,N_7491);
nor U7607 (N_7607,N_7407,N_7469);
nand U7608 (N_7608,N_7435,N_7374);
nor U7609 (N_7609,N_7369,N_7384);
xor U7610 (N_7610,N_7489,N_7372);
xnor U7611 (N_7611,N_7373,N_7513);
nand U7612 (N_7612,N_7475,N_7503);
or U7613 (N_7613,N_7445,N_7467);
and U7614 (N_7614,N_7363,N_7483);
nor U7615 (N_7615,N_7455,N_7501);
nand U7616 (N_7616,N_7388,N_7458);
nand U7617 (N_7617,N_7416,N_7485);
nor U7618 (N_7618,N_7392,N_7442);
xor U7619 (N_7619,N_7447,N_7422);
nand U7620 (N_7620,N_7479,N_7370);
nor U7621 (N_7621,N_7414,N_7361);
xnor U7622 (N_7622,N_7432,N_7469);
xnor U7623 (N_7623,N_7496,N_7460);
nand U7624 (N_7624,N_7461,N_7512);
xor U7625 (N_7625,N_7495,N_7388);
nand U7626 (N_7626,N_7512,N_7400);
or U7627 (N_7627,N_7383,N_7396);
and U7628 (N_7628,N_7473,N_7429);
xor U7629 (N_7629,N_7474,N_7498);
nand U7630 (N_7630,N_7446,N_7364);
nor U7631 (N_7631,N_7405,N_7513);
nand U7632 (N_7632,N_7446,N_7403);
xor U7633 (N_7633,N_7505,N_7481);
xor U7634 (N_7634,N_7373,N_7406);
nor U7635 (N_7635,N_7475,N_7386);
or U7636 (N_7636,N_7387,N_7507);
or U7637 (N_7637,N_7374,N_7379);
nor U7638 (N_7638,N_7465,N_7401);
and U7639 (N_7639,N_7457,N_7478);
nand U7640 (N_7640,N_7423,N_7361);
or U7641 (N_7641,N_7495,N_7382);
and U7642 (N_7642,N_7497,N_7426);
or U7643 (N_7643,N_7362,N_7394);
nor U7644 (N_7644,N_7363,N_7486);
nand U7645 (N_7645,N_7374,N_7471);
nand U7646 (N_7646,N_7447,N_7437);
or U7647 (N_7647,N_7483,N_7447);
and U7648 (N_7648,N_7502,N_7475);
nand U7649 (N_7649,N_7476,N_7515);
xnor U7650 (N_7650,N_7415,N_7422);
nand U7651 (N_7651,N_7457,N_7391);
and U7652 (N_7652,N_7420,N_7498);
nand U7653 (N_7653,N_7432,N_7380);
or U7654 (N_7654,N_7410,N_7445);
nor U7655 (N_7655,N_7413,N_7360);
or U7656 (N_7656,N_7429,N_7412);
or U7657 (N_7657,N_7397,N_7385);
or U7658 (N_7658,N_7465,N_7381);
or U7659 (N_7659,N_7365,N_7479);
nand U7660 (N_7660,N_7519,N_7477);
and U7661 (N_7661,N_7409,N_7479);
xnor U7662 (N_7662,N_7458,N_7402);
nor U7663 (N_7663,N_7489,N_7371);
xnor U7664 (N_7664,N_7389,N_7383);
or U7665 (N_7665,N_7361,N_7374);
or U7666 (N_7666,N_7434,N_7478);
xnor U7667 (N_7667,N_7440,N_7512);
xnor U7668 (N_7668,N_7502,N_7388);
nor U7669 (N_7669,N_7381,N_7478);
nand U7670 (N_7670,N_7383,N_7497);
or U7671 (N_7671,N_7387,N_7457);
or U7672 (N_7672,N_7430,N_7437);
xnor U7673 (N_7673,N_7483,N_7401);
nand U7674 (N_7674,N_7431,N_7437);
or U7675 (N_7675,N_7388,N_7459);
xor U7676 (N_7676,N_7417,N_7376);
or U7677 (N_7677,N_7465,N_7469);
and U7678 (N_7678,N_7439,N_7432);
or U7679 (N_7679,N_7402,N_7489);
and U7680 (N_7680,N_7626,N_7667);
or U7681 (N_7681,N_7602,N_7629);
xor U7682 (N_7682,N_7616,N_7644);
nor U7683 (N_7683,N_7621,N_7587);
or U7684 (N_7684,N_7523,N_7531);
nor U7685 (N_7685,N_7663,N_7595);
nand U7686 (N_7686,N_7532,N_7664);
nor U7687 (N_7687,N_7655,N_7588);
nor U7688 (N_7688,N_7677,N_7582);
or U7689 (N_7689,N_7615,N_7635);
nor U7690 (N_7690,N_7631,N_7641);
nor U7691 (N_7691,N_7653,N_7560);
nand U7692 (N_7692,N_7646,N_7648);
xnor U7693 (N_7693,N_7565,N_7527);
and U7694 (N_7694,N_7557,N_7666);
xnor U7695 (N_7695,N_7617,N_7575);
xor U7696 (N_7696,N_7542,N_7541);
xor U7697 (N_7697,N_7606,N_7651);
or U7698 (N_7698,N_7567,N_7547);
and U7699 (N_7699,N_7630,N_7611);
nor U7700 (N_7700,N_7570,N_7605);
nor U7701 (N_7701,N_7622,N_7632);
xnor U7702 (N_7702,N_7573,N_7571);
or U7703 (N_7703,N_7544,N_7533);
and U7704 (N_7704,N_7665,N_7566);
nor U7705 (N_7705,N_7551,N_7619);
xnor U7706 (N_7706,N_7555,N_7579);
and U7707 (N_7707,N_7558,N_7581);
nor U7708 (N_7708,N_7604,N_7559);
nand U7709 (N_7709,N_7623,N_7613);
nor U7710 (N_7710,N_7625,N_7548);
nor U7711 (N_7711,N_7652,N_7563);
and U7712 (N_7712,N_7539,N_7601);
nand U7713 (N_7713,N_7549,N_7536);
and U7714 (N_7714,N_7524,N_7660);
and U7715 (N_7715,N_7657,N_7642);
nand U7716 (N_7716,N_7650,N_7538);
nor U7717 (N_7717,N_7574,N_7529);
and U7718 (N_7718,N_7535,N_7578);
and U7719 (N_7719,N_7636,N_7675);
xnor U7720 (N_7720,N_7676,N_7645);
and U7721 (N_7721,N_7564,N_7678);
nor U7722 (N_7722,N_7598,N_7600);
xor U7723 (N_7723,N_7639,N_7594);
nor U7724 (N_7724,N_7552,N_7568);
xnor U7725 (N_7725,N_7543,N_7671);
nand U7726 (N_7726,N_7674,N_7597);
nor U7727 (N_7727,N_7537,N_7596);
nand U7728 (N_7728,N_7599,N_7521);
nand U7729 (N_7729,N_7608,N_7591);
and U7730 (N_7730,N_7624,N_7638);
nand U7731 (N_7731,N_7633,N_7586);
or U7732 (N_7732,N_7669,N_7577);
or U7733 (N_7733,N_7620,N_7528);
nand U7734 (N_7734,N_7670,N_7534);
nand U7735 (N_7735,N_7662,N_7576);
or U7736 (N_7736,N_7659,N_7672);
xor U7737 (N_7737,N_7584,N_7592);
nor U7738 (N_7738,N_7612,N_7603);
xnor U7739 (N_7739,N_7580,N_7637);
or U7740 (N_7740,N_7679,N_7583);
nor U7741 (N_7741,N_7561,N_7614);
nand U7742 (N_7742,N_7634,N_7658);
and U7743 (N_7743,N_7618,N_7545);
nand U7744 (N_7744,N_7668,N_7553);
or U7745 (N_7745,N_7520,N_7609);
nand U7746 (N_7746,N_7546,N_7526);
and U7747 (N_7747,N_7661,N_7556);
nand U7748 (N_7748,N_7627,N_7522);
xor U7749 (N_7749,N_7640,N_7593);
or U7750 (N_7750,N_7562,N_7673);
xor U7751 (N_7751,N_7654,N_7590);
nand U7752 (N_7752,N_7589,N_7610);
xnor U7753 (N_7753,N_7647,N_7525);
and U7754 (N_7754,N_7656,N_7649);
and U7755 (N_7755,N_7585,N_7540);
xor U7756 (N_7756,N_7550,N_7607);
xor U7757 (N_7757,N_7628,N_7554);
nand U7758 (N_7758,N_7530,N_7643);
xnor U7759 (N_7759,N_7569,N_7572);
and U7760 (N_7760,N_7670,N_7543);
nand U7761 (N_7761,N_7594,N_7571);
nor U7762 (N_7762,N_7592,N_7635);
or U7763 (N_7763,N_7552,N_7668);
and U7764 (N_7764,N_7657,N_7673);
and U7765 (N_7765,N_7587,N_7539);
or U7766 (N_7766,N_7663,N_7527);
xnor U7767 (N_7767,N_7642,N_7542);
nand U7768 (N_7768,N_7576,N_7563);
and U7769 (N_7769,N_7565,N_7593);
and U7770 (N_7770,N_7555,N_7571);
nor U7771 (N_7771,N_7662,N_7571);
and U7772 (N_7772,N_7658,N_7666);
nand U7773 (N_7773,N_7663,N_7569);
or U7774 (N_7774,N_7618,N_7555);
nor U7775 (N_7775,N_7660,N_7609);
nor U7776 (N_7776,N_7636,N_7560);
nor U7777 (N_7777,N_7526,N_7522);
or U7778 (N_7778,N_7665,N_7568);
xnor U7779 (N_7779,N_7612,N_7568);
xnor U7780 (N_7780,N_7618,N_7634);
and U7781 (N_7781,N_7576,N_7572);
xor U7782 (N_7782,N_7621,N_7652);
and U7783 (N_7783,N_7549,N_7623);
nand U7784 (N_7784,N_7533,N_7642);
xor U7785 (N_7785,N_7585,N_7613);
and U7786 (N_7786,N_7599,N_7573);
and U7787 (N_7787,N_7588,N_7607);
or U7788 (N_7788,N_7532,N_7594);
xor U7789 (N_7789,N_7655,N_7658);
or U7790 (N_7790,N_7657,N_7557);
and U7791 (N_7791,N_7527,N_7621);
nand U7792 (N_7792,N_7554,N_7637);
xor U7793 (N_7793,N_7561,N_7603);
xor U7794 (N_7794,N_7575,N_7625);
nor U7795 (N_7795,N_7570,N_7591);
nand U7796 (N_7796,N_7523,N_7600);
xnor U7797 (N_7797,N_7606,N_7573);
nor U7798 (N_7798,N_7585,N_7639);
xnor U7799 (N_7799,N_7563,N_7579);
nor U7800 (N_7800,N_7551,N_7547);
xor U7801 (N_7801,N_7678,N_7529);
nand U7802 (N_7802,N_7598,N_7539);
and U7803 (N_7803,N_7589,N_7658);
nand U7804 (N_7804,N_7679,N_7571);
nand U7805 (N_7805,N_7577,N_7650);
xor U7806 (N_7806,N_7625,N_7675);
and U7807 (N_7807,N_7625,N_7673);
or U7808 (N_7808,N_7573,N_7590);
or U7809 (N_7809,N_7609,N_7625);
nor U7810 (N_7810,N_7594,N_7614);
or U7811 (N_7811,N_7572,N_7615);
and U7812 (N_7812,N_7631,N_7605);
and U7813 (N_7813,N_7677,N_7597);
or U7814 (N_7814,N_7636,N_7674);
nand U7815 (N_7815,N_7604,N_7611);
or U7816 (N_7816,N_7647,N_7556);
or U7817 (N_7817,N_7635,N_7629);
and U7818 (N_7818,N_7570,N_7559);
nor U7819 (N_7819,N_7542,N_7653);
and U7820 (N_7820,N_7565,N_7553);
or U7821 (N_7821,N_7641,N_7559);
nor U7822 (N_7822,N_7629,N_7582);
or U7823 (N_7823,N_7522,N_7657);
or U7824 (N_7824,N_7535,N_7591);
nand U7825 (N_7825,N_7621,N_7639);
nand U7826 (N_7826,N_7619,N_7565);
xor U7827 (N_7827,N_7585,N_7538);
xor U7828 (N_7828,N_7679,N_7660);
xor U7829 (N_7829,N_7664,N_7562);
or U7830 (N_7830,N_7651,N_7614);
or U7831 (N_7831,N_7577,N_7629);
and U7832 (N_7832,N_7618,N_7554);
xor U7833 (N_7833,N_7601,N_7549);
nand U7834 (N_7834,N_7621,N_7656);
xor U7835 (N_7835,N_7641,N_7592);
nand U7836 (N_7836,N_7576,N_7650);
and U7837 (N_7837,N_7567,N_7606);
xnor U7838 (N_7838,N_7586,N_7659);
nor U7839 (N_7839,N_7547,N_7616);
and U7840 (N_7840,N_7706,N_7718);
xnor U7841 (N_7841,N_7764,N_7741);
or U7842 (N_7842,N_7698,N_7696);
or U7843 (N_7843,N_7795,N_7762);
and U7844 (N_7844,N_7729,N_7783);
nand U7845 (N_7845,N_7827,N_7799);
or U7846 (N_7846,N_7801,N_7756);
nand U7847 (N_7847,N_7808,N_7763);
and U7848 (N_7848,N_7750,N_7720);
nand U7849 (N_7849,N_7812,N_7839);
or U7850 (N_7850,N_7734,N_7733);
nor U7851 (N_7851,N_7830,N_7722);
or U7852 (N_7852,N_7794,N_7784);
nand U7853 (N_7853,N_7754,N_7715);
xnor U7854 (N_7854,N_7702,N_7802);
nand U7855 (N_7855,N_7695,N_7781);
nand U7856 (N_7856,N_7811,N_7758);
nand U7857 (N_7857,N_7690,N_7787);
and U7858 (N_7858,N_7680,N_7692);
or U7859 (N_7859,N_7831,N_7752);
nor U7860 (N_7860,N_7791,N_7719);
nand U7861 (N_7861,N_7714,N_7745);
nor U7862 (N_7862,N_7828,N_7689);
xnor U7863 (N_7863,N_7742,N_7759);
or U7864 (N_7864,N_7682,N_7738);
or U7865 (N_7865,N_7814,N_7786);
xnor U7866 (N_7866,N_7780,N_7751);
and U7867 (N_7867,N_7772,N_7815);
nand U7868 (N_7868,N_7761,N_7757);
xnor U7869 (N_7869,N_7701,N_7712);
nor U7870 (N_7870,N_7825,N_7697);
nand U7871 (N_7871,N_7768,N_7806);
xnor U7872 (N_7872,N_7837,N_7823);
xnor U7873 (N_7873,N_7708,N_7833);
nand U7874 (N_7874,N_7797,N_7707);
nand U7875 (N_7875,N_7703,N_7727);
xor U7876 (N_7876,N_7832,N_7771);
and U7877 (N_7877,N_7728,N_7743);
nand U7878 (N_7878,N_7782,N_7735);
nand U7879 (N_7879,N_7793,N_7760);
nor U7880 (N_7880,N_7813,N_7717);
or U7881 (N_7881,N_7713,N_7681);
and U7882 (N_7882,N_7809,N_7816);
nor U7883 (N_7883,N_7822,N_7687);
xor U7884 (N_7884,N_7705,N_7800);
nand U7885 (N_7885,N_7834,N_7723);
or U7886 (N_7886,N_7753,N_7818);
and U7887 (N_7887,N_7798,N_7805);
or U7888 (N_7888,N_7765,N_7688);
and U7889 (N_7889,N_7835,N_7699);
or U7890 (N_7890,N_7819,N_7776);
xor U7891 (N_7891,N_7724,N_7691);
or U7892 (N_7892,N_7836,N_7792);
nor U7893 (N_7893,N_7767,N_7803);
nand U7894 (N_7894,N_7769,N_7770);
nor U7895 (N_7895,N_7748,N_7704);
xor U7896 (N_7896,N_7777,N_7725);
nand U7897 (N_7897,N_7684,N_7726);
xnor U7898 (N_7898,N_7755,N_7820);
or U7899 (N_7899,N_7746,N_7826);
or U7900 (N_7900,N_7773,N_7693);
nand U7901 (N_7901,N_7747,N_7817);
or U7902 (N_7902,N_7779,N_7778);
xnor U7903 (N_7903,N_7694,N_7774);
or U7904 (N_7904,N_7744,N_7824);
nor U7905 (N_7905,N_7710,N_7821);
xor U7906 (N_7906,N_7685,N_7711);
nor U7907 (N_7907,N_7789,N_7730);
or U7908 (N_7908,N_7683,N_7829);
or U7909 (N_7909,N_7766,N_7807);
xnor U7910 (N_7910,N_7732,N_7788);
nand U7911 (N_7911,N_7737,N_7790);
xnor U7912 (N_7912,N_7804,N_7709);
nand U7913 (N_7913,N_7838,N_7749);
xnor U7914 (N_7914,N_7785,N_7739);
or U7915 (N_7915,N_7716,N_7700);
and U7916 (N_7916,N_7796,N_7736);
xor U7917 (N_7917,N_7731,N_7721);
xor U7918 (N_7918,N_7810,N_7775);
nor U7919 (N_7919,N_7740,N_7686);
nand U7920 (N_7920,N_7739,N_7745);
and U7921 (N_7921,N_7815,N_7720);
nand U7922 (N_7922,N_7716,N_7730);
xnor U7923 (N_7923,N_7731,N_7735);
xnor U7924 (N_7924,N_7772,N_7746);
xor U7925 (N_7925,N_7697,N_7684);
nand U7926 (N_7926,N_7828,N_7684);
nand U7927 (N_7927,N_7821,N_7801);
and U7928 (N_7928,N_7730,N_7782);
or U7929 (N_7929,N_7825,N_7834);
or U7930 (N_7930,N_7711,N_7833);
nor U7931 (N_7931,N_7819,N_7693);
nor U7932 (N_7932,N_7720,N_7790);
xor U7933 (N_7933,N_7742,N_7756);
and U7934 (N_7934,N_7799,N_7834);
and U7935 (N_7935,N_7752,N_7745);
and U7936 (N_7936,N_7772,N_7687);
nor U7937 (N_7937,N_7726,N_7825);
and U7938 (N_7938,N_7793,N_7766);
and U7939 (N_7939,N_7755,N_7772);
xor U7940 (N_7940,N_7712,N_7700);
and U7941 (N_7941,N_7832,N_7708);
nor U7942 (N_7942,N_7822,N_7754);
or U7943 (N_7943,N_7826,N_7686);
nor U7944 (N_7944,N_7751,N_7723);
and U7945 (N_7945,N_7832,N_7778);
and U7946 (N_7946,N_7749,N_7696);
nand U7947 (N_7947,N_7697,N_7695);
and U7948 (N_7948,N_7824,N_7798);
or U7949 (N_7949,N_7795,N_7690);
nand U7950 (N_7950,N_7823,N_7680);
xor U7951 (N_7951,N_7694,N_7729);
nand U7952 (N_7952,N_7781,N_7718);
nor U7953 (N_7953,N_7699,N_7838);
xor U7954 (N_7954,N_7738,N_7797);
or U7955 (N_7955,N_7783,N_7706);
and U7956 (N_7956,N_7753,N_7835);
nor U7957 (N_7957,N_7732,N_7793);
nand U7958 (N_7958,N_7809,N_7771);
or U7959 (N_7959,N_7706,N_7832);
nand U7960 (N_7960,N_7694,N_7773);
nand U7961 (N_7961,N_7789,N_7806);
or U7962 (N_7962,N_7726,N_7828);
xor U7963 (N_7963,N_7813,N_7746);
and U7964 (N_7964,N_7774,N_7826);
nor U7965 (N_7965,N_7703,N_7801);
or U7966 (N_7966,N_7834,N_7704);
nand U7967 (N_7967,N_7724,N_7738);
nand U7968 (N_7968,N_7831,N_7706);
nor U7969 (N_7969,N_7783,N_7697);
xor U7970 (N_7970,N_7809,N_7737);
xor U7971 (N_7971,N_7833,N_7683);
or U7972 (N_7972,N_7706,N_7756);
xnor U7973 (N_7973,N_7809,N_7786);
or U7974 (N_7974,N_7836,N_7763);
or U7975 (N_7975,N_7811,N_7835);
or U7976 (N_7976,N_7794,N_7701);
nand U7977 (N_7977,N_7742,N_7769);
and U7978 (N_7978,N_7681,N_7692);
nor U7979 (N_7979,N_7722,N_7750);
nor U7980 (N_7980,N_7743,N_7781);
and U7981 (N_7981,N_7747,N_7826);
nand U7982 (N_7982,N_7747,N_7779);
and U7983 (N_7983,N_7821,N_7691);
nor U7984 (N_7984,N_7822,N_7800);
and U7985 (N_7985,N_7720,N_7769);
nand U7986 (N_7986,N_7825,N_7805);
nor U7987 (N_7987,N_7697,N_7752);
xor U7988 (N_7988,N_7810,N_7727);
xor U7989 (N_7989,N_7725,N_7707);
nand U7990 (N_7990,N_7826,N_7813);
nand U7991 (N_7991,N_7747,N_7694);
or U7992 (N_7992,N_7773,N_7807);
and U7993 (N_7993,N_7780,N_7825);
nor U7994 (N_7994,N_7764,N_7687);
xnor U7995 (N_7995,N_7792,N_7798);
xor U7996 (N_7996,N_7758,N_7786);
and U7997 (N_7997,N_7773,N_7703);
nand U7998 (N_7998,N_7696,N_7746);
or U7999 (N_7999,N_7813,N_7699);
and U8000 (N_8000,N_7935,N_7945);
or U8001 (N_8001,N_7856,N_7874);
nand U8002 (N_8002,N_7992,N_7900);
and U8003 (N_8003,N_7887,N_7854);
xor U8004 (N_8004,N_7853,N_7847);
nor U8005 (N_8005,N_7988,N_7848);
or U8006 (N_8006,N_7923,N_7949);
nand U8007 (N_8007,N_7989,N_7991);
or U8008 (N_8008,N_7963,N_7946);
nor U8009 (N_8009,N_7855,N_7908);
xor U8010 (N_8010,N_7893,N_7926);
xnor U8011 (N_8011,N_7944,N_7960);
or U8012 (N_8012,N_7934,N_7849);
xor U8013 (N_8013,N_7857,N_7880);
and U8014 (N_8014,N_7879,N_7948);
nor U8015 (N_8015,N_7843,N_7890);
nor U8016 (N_8016,N_7902,N_7881);
and U8017 (N_8017,N_7999,N_7928);
xnor U8018 (N_8018,N_7937,N_7905);
nand U8019 (N_8019,N_7886,N_7955);
and U8020 (N_8020,N_7921,N_7965);
or U8021 (N_8021,N_7968,N_7967);
and U8022 (N_8022,N_7850,N_7914);
xnor U8023 (N_8023,N_7891,N_7922);
nor U8024 (N_8024,N_7933,N_7942);
or U8025 (N_8025,N_7950,N_7977);
and U8026 (N_8026,N_7998,N_7938);
nand U8027 (N_8027,N_7846,N_7986);
nor U8028 (N_8028,N_7978,N_7969);
nand U8029 (N_8029,N_7985,N_7917);
xor U8030 (N_8030,N_7918,N_7876);
nand U8031 (N_8031,N_7872,N_7907);
and U8032 (N_8032,N_7841,N_7929);
xor U8033 (N_8033,N_7971,N_7994);
nor U8034 (N_8034,N_7973,N_7844);
and U8035 (N_8035,N_7924,N_7885);
and U8036 (N_8036,N_7952,N_7901);
xnor U8037 (N_8037,N_7882,N_7959);
or U8038 (N_8038,N_7927,N_7883);
or U8039 (N_8039,N_7852,N_7851);
or U8040 (N_8040,N_7983,N_7972);
nor U8041 (N_8041,N_7873,N_7966);
nor U8042 (N_8042,N_7916,N_7982);
and U8043 (N_8043,N_7884,N_7892);
or U8044 (N_8044,N_7863,N_7899);
and U8045 (N_8045,N_7995,N_7906);
xor U8046 (N_8046,N_7984,N_7996);
and U8047 (N_8047,N_7990,N_7909);
nor U8048 (N_8048,N_7866,N_7889);
nor U8049 (N_8049,N_7870,N_7930);
nor U8050 (N_8050,N_7915,N_7862);
or U8051 (N_8051,N_7957,N_7940);
nand U8052 (N_8052,N_7859,N_7869);
nor U8053 (N_8053,N_7910,N_7840);
and U8054 (N_8054,N_7931,N_7919);
or U8055 (N_8055,N_7964,N_7941);
nand U8056 (N_8056,N_7913,N_7936);
xor U8057 (N_8057,N_7947,N_7970);
or U8058 (N_8058,N_7904,N_7962);
xor U8059 (N_8059,N_7865,N_7932);
and U8060 (N_8060,N_7980,N_7867);
nand U8061 (N_8061,N_7981,N_7911);
and U8062 (N_8062,N_7895,N_7976);
nand U8063 (N_8063,N_7888,N_7896);
and U8064 (N_8064,N_7997,N_7958);
xor U8065 (N_8065,N_7974,N_7858);
xnor U8066 (N_8066,N_7860,N_7868);
or U8067 (N_8067,N_7956,N_7975);
nand U8068 (N_8068,N_7897,N_7993);
nand U8069 (N_8069,N_7939,N_7878);
and U8070 (N_8070,N_7954,N_7845);
or U8071 (N_8071,N_7920,N_7875);
nor U8072 (N_8072,N_7987,N_7871);
nand U8073 (N_8073,N_7953,N_7925);
and U8074 (N_8074,N_7979,N_7877);
and U8075 (N_8075,N_7961,N_7951);
xnor U8076 (N_8076,N_7894,N_7864);
nor U8077 (N_8077,N_7898,N_7861);
xor U8078 (N_8078,N_7903,N_7842);
and U8079 (N_8079,N_7912,N_7943);
or U8080 (N_8080,N_7878,N_7971);
and U8081 (N_8081,N_7893,N_7918);
or U8082 (N_8082,N_7956,N_7923);
nand U8083 (N_8083,N_7878,N_7993);
and U8084 (N_8084,N_7944,N_7865);
nand U8085 (N_8085,N_7872,N_7945);
xor U8086 (N_8086,N_7887,N_7855);
nor U8087 (N_8087,N_7917,N_7998);
nand U8088 (N_8088,N_7881,N_7893);
and U8089 (N_8089,N_7967,N_7927);
nor U8090 (N_8090,N_7995,N_7847);
nand U8091 (N_8091,N_7858,N_7894);
xor U8092 (N_8092,N_7938,N_7982);
nor U8093 (N_8093,N_7875,N_7982);
nand U8094 (N_8094,N_7855,N_7973);
xor U8095 (N_8095,N_7979,N_7918);
or U8096 (N_8096,N_7899,N_7961);
nor U8097 (N_8097,N_7918,N_7946);
nand U8098 (N_8098,N_7871,N_7959);
nand U8099 (N_8099,N_7856,N_7932);
nand U8100 (N_8100,N_7886,N_7889);
and U8101 (N_8101,N_7938,N_7948);
nor U8102 (N_8102,N_7922,N_7997);
and U8103 (N_8103,N_7864,N_7842);
nor U8104 (N_8104,N_7888,N_7866);
xor U8105 (N_8105,N_7870,N_7907);
xnor U8106 (N_8106,N_7892,N_7851);
or U8107 (N_8107,N_7909,N_7906);
xnor U8108 (N_8108,N_7984,N_7873);
or U8109 (N_8109,N_7868,N_7993);
nor U8110 (N_8110,N_7891,N_7882);
nor U8111 (N_8111,N_7874,N_7938);
xnor U8112 (N_8112,N_7889,N_7861);
or U8113 (N_8113,N_7861,N_7963);
nor U8114 (N_8114,N_7883,N_7856);
nand U8115 (N_8115,N_7857,N_7894);
and U8116 (N_8116,N_7915,N_7996);
or U8117 (N_8117,N_7946,N_7861);
xnor U8118 (N_8118,N_7902,N_7954);
xor U8119 (N_8119,N_7873,N_7919);
nand U8120 (N_8120,N_7869,N_7945);
nor U8121 (N_8121,N_7906,N_7911);
nand U8122 (N_8122,N_7918,N_7915);
and U8123 (N_8123,N_7893,N_7847);
nor U8124 (N_8124,N_7873,N_7861);
or U8125 (N_8125,N_7898,N_7930);
nand U8126 (N_8126,N_7917,N_7899);
and U8127 (N_8127,N_7948,N_7842);
or U8128 (N_8128,N_7923,N_7928);
xnor U8129 (N_8129,N_7968,N_7864);
or U8130 (N_8130,N_7950,N_7899);
xor U8131 (N_8131,N_7893,N_7998);
xor U8132 (N_8132,N_7901,N_7977);
xor U8133 (N_8133,N_7912,N_7923);
nand U8134 (N_8134,N_7845,N_7862);
nand U8135 (N_8135,N_7973,N_7908);
xor U8136 (N_8136,N_7982,N_7879);
xnor U8137 (N_8137,N_7956,N_7862);
xor U8138 (N_8138,N_7870,N_7901);
nor U8139 (N_8139,N_7848,N_7853);
xor U8140 (N_8140,N_7886,N_7944);
xor U8141 (N_8141,N_7898,N_7995);
and U8142 (N_8142,N_7971,N_7973);
and U8143 (N_8143,N_7978,N_7914);
nor U8144 (N_8144,N_7900,N_7994);
xor U8145 (N_8145,N_7910,N_7887);
nor U8146 (N_8146,N_7973,N_7868);
nand U8147 (N_8147,N_7861,N_7854);
xor U8148 (N_8148,N_7970,N_7880);
nor U8149 (N_8149,N_7882,N_7953);
nand U8150 (N_8150,N_7874,N_7870);
nand U8151 (N_8151,N_7883,N_7863);
and U8152 (N_8152,N_7910,N_7898);
nand U8153 (N_8153,N_7869,N_7881);
or U8154 (N_8154,N_7953,N_7923);
nor U8155 (N_8155,N_7849,N_7887);
xnor U8156 (N_8156,N_7991,N_7843);
and U8157 (N_8157,N_7910,N_7903);
nor U8158 (N_8158,N_7906,N_7968);
nand U8159 (N_8159,N_7902,N_7973);
and U8160 (N_8160,N_8094,N_8100);
nor U8161 (N_8161,N_8014,N_8134);
nor U8162 (N_8162,N_8101,N_8062);
xnor U8163 (N_8163,N_8002,N_8072);
or U8164 (N_8164,N_8027,N_8077);
nor U8165 (N_8165,N_8079,N_8128);
xor U8166 (N_8166,N_8105,N_8143);
nor U8167 (N_8167,N_8037,N_8082);
xnor U8168 (N_8168,N_8000,N_8118);
or U8169 (N_8169,N_8106,N_8123);
or U8170 (N_8170,N_8113,N_8036);
nor U8171 (N_8171,N_8125,N_8075);
xnor U8172 (N_8172,N_8110,N_8074);
and U8173 (N_8173,N_8119,N_8097);
or U8174 (N_8174,N_8147,N_8108);
and U8175 (N_8175,N_8070,N_8006);
nor U8176 (N_8176,N_8124,N_8022);
nand U8177 (N_8177,N_8035,N_8059);
nand U8178 (N_8178,N_8144,N_8088);
nor U8179 (N_8179,N_8126,N_8137);
xor U8180 (N_8180,N_8056,N_8052);
nor U8181 (N_8181,N_8115,N_8007);
and U8182 (N_8182,N_8004,N_8151);
nor U8183 (N_8183,N_8005,N_8020);
nand U8184 (N_8184,N_8089,N_8140);
and U8185 (N_8185,N_8114,N_8139);
or U8186 (N_8186,N_8107,N_8026);
or U8187 (N_8187,N_8154,N_8029);
xnor U8188 (N_8188,N_8068,N_8085);
nor U8189 (N_8189,N_8017,N_8092);
or U8190 (N_8190,N_8042,N_8055);
and U8191 (N_8191,N_8048,N_8112);
or U8192 (N_8192,N_8011,N_8127);
and U8193 (N_8193,N_8087,N_8116);
nor U8194 (N_8194,N_8096,N_8031);
and U8195 (N_8195,N_8155,N_8086);
nand U8196 (N_8196,N_8095,N_8003);
nand U8197 (N_8197,N_8044,N_8083);
nand U8198 (N_8198,N_8061,N_8084);
nor U8199 (N_8199,N_8013,N_8030);
or U8200 (N_8200,N_8152,N_8051);
or U8201 (N_8201,N_8148,N_8111);
and U8202 (N_8202,N_8023,N_8104);
nand U8203 (N_8203,N_8025,N_8135);
nand U8204 (N_8204,N_8131,N_8133);
xnor U8205 (N_8205,N_8149,N_8129);
xnor U8206 (N_8206,N_8136,N_8159);
nor U8207 (N_8207,N_8039,N_8049);
nand U8208 (N_8208,N_8099,N_8073);
or U8209 (N_8209,N_8078,N_8040);
xnor U8210 (N_8210,N_8080,N_8019);
and U8211 (N_8211,N_8033,N_8142);
and U8212 (N_8212,N_8141,N_8153);
nor U8213 (N_8213,N_8021,N_8145);
nand U8214 (N_8214,N_8066,N_8008);
or U8215 (N_8215,N_8121,N_8117);
nor U8216 (N_8216,N_8045,N_8001);
xor U8217 (N_8217,N_8067,N_8034);
nor U8218 (N_8218,N_8157,N_8053);
nand U8219 (N_8219,N_8057,N_8063);
nand U8220 (N_8220,N_8109,N_8046);
nand U8221 (N_8221,N_8050,N_8024);
or U8222 (N_8222,N_8138,N_8076);
xnor U8223 (N_8223,N_8060,N_8058);
and U8224 (N_8224,N_8043,N_8122);
nor U8225 (N_8225,N_8156,N_8047);
and U8226 (N_8226,N_8010,N_8069);
xnor U8227 (N_8227,N_8012,N_8158);
nor U8228 (N_8228,N_8038,N_8064);
and U8229 (N_8229,N_8028,N_8032);
or U8230 (N_8230,N_8016,N_8098);
and U8231 (N_8231,N_8120,N_8103);
or U8232 (N_8232,N_8054,N_8150);
xnor U8233 (N_8233,N_8009,N_8071);
and U8234 (N_8234,N_8081,N_8091);
xor U8235 (N_8235,N_8090,N_8041);
nor U8236 (N_8236,N_8093,N_8065);
nand U8237 (N_8237,N_8018,N_8146);
and U8238 (N_8238,N_8132,N_8102);
or U8239 (N_8239,N_8015,N_8130);
and U8240 (N_8240,N_8138,N_8063);
and U8241 (N_8241,N_8120,N_8027);
nand U8242 (N_8242,N_8054,N_8013);
and U8243 (N_8243,N_8043,N_8145);
and U8244 (N_8244,N_8002,N_8088);
nor U8245 (N_8245,N_8010,N_8145);
nor U8246 (N_8246,N_8116,N_8106);
nand U8247 (N_8247,N_8065,N_8108);
nor U8248 (N_8248,N_8091,N_8113);
and U8249 (N_8249,N_8033,N_8090);
nor U8250 (N_8250,N_8006,N_8038);
or U8251 (N_8251,N_8141,N_8126);
or U8252 (N_8252,N_8103,N_8135);
or U8253 (N_8253,N_8055,N_8156);
nor U8254 (N_8254,N_8040,N_8013);
xor U8255 (N_8255,N_8069,N_8120);
nor U8256 (N_8256,N_8102,N_8134);
nor U8257 (N_8257,N_8000,N_8080);
or U8258 (N_8258,N_8094,N_8007);
or U8259 (N_8259,N_8153,N_8045);
and U8260 (N_8260,N_8121,N_8047);
or U8261 (N_8261,N_8115,N_8075);
nor U8262 (N_8262,N_8081,N_8026);
nand U8263 (N_8263,N_8104,N_8156);
xor U8264 (N_8264,N_8095,N_8017);
xor U8265 (N_8265,N_8026,N_8100);
xnor U8266 (N_8266,N_8064,N_8075);
and U8267 (N_8267,N_8069,N_8031);
xnor U8268 (N_8268,N_8145,N_8022);
or U8269 (N_8269,N_8060,N_8074);
xor U8270 (N_8270,N_8027,N_8110);
and U8271 (N_8271,N_8000,N_8076);
nand U8272 (N_8272,N_8088,N_8147);
xnor U8273 (N_8273,N_8043,N_8139);
xor U8274 (N_8274,N_8092,N_8087);
and U8275 (N_8275,N_8048,N_8141);
nor U8276 (N_8276,N_8108,N_8058);
xor U8277 (N_8277,N_8105,N_8001);
nand U8278 (N_8278,N_8088,N_8062);
xor U8279 (N_8279,N_8034,N_8020);
xnor U8280 (N_8280,N_8076,N_8084);
and U8281 (N_8281,N_8055,N_8020);
and U8282 (N_8282,N_8045,N_8084);
xnor U8283 (N_8283,N_8023,N_8154);
xor U8284 (N_8284,N_8059,N_8093);
and U8285 (N_8285,N_8150,N_8113);
or U8286 (N_8286,N_8113,N_8032);
xnor U8287 (N_8287,N_8072,N_8052);
nor U8288 (N_8288,N_8132,N_8028);
nand U8289 (N_8289,N_8157,N_8116);
and U8290 (N_8290,N_8116,N_8092);
nand U8291 (N_8291,N_8130,N_8018);
or U8292 (N_8292,N_8098,N_8110);
nor U8293 (N_8293,N_8013,N_8149);
nor U8294 (N_8294,N_8065,N_8049);
or U8295 (N_8295,N_8068,N_8153);
or U8296 (N_8296,N_8109,N_8076);
or U8297 (N_8297,N_8038,N_8033);
nor U8298 (N_8298,N_8016,N_8104);
nand U8299 (N_8299,N_8099,N_8000);
or U8300 (N_8300,N_8078,N_8044);
nand U8301 (N_8301,N_8106,N_8146);
nand U8302 (N_8302,N_8002,N_8032);
or U8303 (N_8303,N_8104,N_8032);
xnor U8304 (N_8304,N_8062,N_8043);
and U8305 (N_8305,N_8039,N_8034);
xnor U8306 (N_8306,N_8022,N_8068);
and U8307 (N_8307,N_8084,N_8012);
nand U8308 (N_8308,N_8053,N_8122);
nand U8309 (N_8309,N_8115,N_8079);
nand U8310 (N_8310,N_8123,N_8105);
nor U8311 (N_8311,N_8126,N_8013);
or U8312 (N_8312,N_8015,N_8059);
and U8313 (N_8313,N_8076,N_8052);
xor U8314 (N_8314,N_8001,N_8020);
nor U8315 (N_8315,N_8138,N_8150);
nor U8316 (N_8316,N_8085,N_8012);
nor U8317 (N_8317,N_8088,N_8152);
nor U8318 (N_8318,N_8088,N_8029);
nand U8319 (N_8319,N_8027,N_8108);
nand U8320 (N_8320,N_8218,N_8161);
nand U8321 (N_8321,N_8205,N_8303);
and U8322 (N_8322,N_8209,N_8263);
xor U8323 (N_8323,N_8227,N_8253);
nand U8324 (N_8324,N_8222,N_8273);
nand U8325 (N_8325,N_8245,N_8219);
xor U8326 (N_8326,N_8224,N_8292);
nand U8327 (N_8327,N_8255,N_8283);
or U8328 (N_8328,N_8233,N_8295);
xor U8329 (N_8329,N_8201,N_8204);
and U8330 (N_8330,N_8257,N_8185);
nand U8331 (N_8331,N_8293,N_8314);
and U8332 (N_8332,N_8168,N_8199);
nand U8333 (N_8333,N_8179,N_8306);
nor U8334 (N_8334,N_8296,N_8301);
nand U8335 (N_8335,N_8281,N_8284);
or U8336 (N_8336,N_8318,N_8234);
nand U8337 (N_8337,N_8210,N_8177);
nand U8338 (N_8338,N_8265,N_8237);
xnor U8339 (N_8339,N_8180,N_8243);
and U8340 (N_8340,N_8195,N_8280);
nor U8341 (N_8341,N_8276,N_8275);
and U8342 (N_8342,N_8184,N_8240);
nand U8343 (N_8343,N_8178,N_8191);
nor U8344 (N_8344,N_8260,N_8213);
or U8345 (N_8345,N_8236,N_8262);
nor U8346 (N_8346,N_8172,N_8194);
nor U8347 (N_8347,N_8193,N_8174);
nor U8348 (N_8348,N_8220,N_8216);
xor U8349 (N_8349,N_8206,N_8305);
xnor U8350 (N_8350,N_8186,N_8256);
nand U8351 (N_8351,N_8182,N_8183);
and U8352 (N_8352,N_8162,N_8259);
and U8353 (N_8353,N_8287,N_8315);
nor U8354 (N_8354,N_8254,N_8304);
or U8355 (N_8355,N_8181,N_8268);
and U8356 (N_8356,N_8290,N_8228);
nand U8357 (N_8357,N_8238,N_8249);
xor U8358 (N_8358,N_8308,N_8307);
nor U8359 (N_8359,N_8267,N_8163);
or U8360 (N_8360,N_8312,N_8248);
nand U8361 (N_8361,N_8202,N_8317);
or U8362 (N_8362,N_8198,N_8190);
xnor U8363 (N_8363,N_8300,N_8244);
and U8364 (N_8364,N_8231,N_8250);
or U8365 (N_8365,N_8241,N_8196);
nand U8366 (N_8366,N_8282,N_8242);
nand U8367 (N_8367,N_8203,N_8160);
xnor U8368 (N_8368,N_8310,N_8247);
nor U8369 (N_8369,N_8211,N_8167);
nor U8370 (N_8370,N_8298,N_8229);
nand U8371 (N_8371,N_8169,N_8272);
nand U8372 (N_8372,N_8309,N_8217);
and U8373 (N_8373,N_8264,N_8269);
or U8374 (N_8374,N_8289,N_8230);
nand U8375 (N_8375,N_8246,N_8302);
nor U8376 (N_8376,N_8207,N_8166);
nand U8377 (N_8377,N_8286,N_8258);
xnor U8378 (N_8378,N_8274,N_8212);
nor U8379 (N_8379,N_8200,N_8173);
and U8380 (N_8380,N_8266,N_8313);
xor U8381 (N_8381,N_8188,N_8165);
nor U8382 (N_8382,N_8225,N_8171);
nor U8383 (N_8383,N_8294,N_8271);
nand U8384 (N_8384,N_8175,N_8299);
and U8385 (N_8385,N_8197,N_8311);
nor U8386 (N_8386,N_8297,N_8221);
nand U8387 (N_8387,N_8319,N_8164);
nor U8388 (N_8388,N_8176,N_8291);
or U8389 (N_8389,N_8278,N_8279);
and U8390 (N_8390,N_8261,N_8239);
xnor U8391 (N_8391,N_8170,N_8189);
and U8392 (N_8392,N_8251,N_8285);
xnor U8393 (N_8393,N_8277,N_8252);
nor U8394 (N_8394,N_8208,N_8215);
xor U8395 (N_8395,N_8214,N_8288);
or U8396 (N_8396,N_8316,N_8187);
nor U8397 (N_8397,N_8270,N_8226);
nand U8398 (N_8398,N_8235,N_8223);
nor U8399 (N_8399,N_8232,N_8192);
xnor U8400 (N_8400,N_8193,N_8179);
and U8401 (N_8401,N_8199,N_8242);
or U8402 (N_8402,N_8286,N_8162);
and U8403 (N_8403,N_8213,N_8276);
and U8404 (N_8404,N_8271,N_8313);
nor U8405 (N_8405,N_8166,N_8268);
and U8406 (N_8406,N_8198,N_8222);
xnor U8407 (N_8407,N_8228,N_8279);
nor U8408 (N_8408,N_8311,N_8223);
and U8409 (N_8409,N_8292,N_8214);
xnor U8410 (N_8410,N_8165,N_8198);
xnor U8411 (N_8411,N_8164,N_8278);
xor U8412 (N_8412,N_8272,N_8312);
nand U8413 (N_8413,N_8294,N_8295);
nor U8414 (N_8414,N_8190,N_8176);
nor U8415 (N_8415,N_8297,N_8303);
and U8416 (N_8416,N_8200,N_8301);
or U8417 (N_8417,N_8208,N_8296);
or U8418 (N_8418,N_8257,N_8313);
or U8419 (N_8419,N_8218,N_8305);
xnor U8420 (N_8420,N_8319,N_8274);
and U8421 (N_8421,N_8183,N_8317);
or U8422 (N_8422,N_8243,N_8301);
or U8423 (N_8423,N_8238,N_8189);
nor U8424 (N_8424,N_8201,N_8271);
or U8425 (N_8425,N_8186,N_8285);
nor U8426 (N_8426,N_8228,N_8194);
nand U8427 (N_8427,N_8285,N_8209);
or U8428 (N_8428,N_8220,N_8215);
and U8429 (N_8429,N_8217,N_8226);
or U8430 (N_8430,N_8174,N_8175);
and U8431 (N_8431,N_8189,N_8299);
nor U8432 (N_8432,N_8181,N_8173);
or U8433 (N_8433,N_8292,N_8245);
or U8434 (N_8434,N_8257,N_8192);
xnor U8435 (N_8435,N_8270,N_8283);
nand U8436 (N_8436,N_8219,N_8311);
nand U8437 (N_8437,N_8241,N_8213);
and U8438 (N_8438,N_8167,N_8239);
nor U8439 (N_8439,N_8208,N_8210);
or U8440 (N_8440,N_8179,N_8304);
nor U8441 (N_8441,N_8237,N_8292);
or U8442 (N_8442,N_8216,N_8256);
xor U8443 (N_8443,N_8271,N_8245);
nand U8444 (N_8444,N_8205,N_8314);
nor U8445 (N_8445,N_8230,N_8192);
nor U8446 (N_8446,N_8315,N_8306);
or U8447 (N_8447,N_8243,N_8234);
and U8448 (N_8448,N_8302,N_8198);
nor U8449 (N_8449,N_8313,N_8184);
or U8450 (N_8450,N_8205,N_8164);
nand U8451 (N_8451,N_8289,N_8300);
and U8452 (N_8452,N_8220,N_8198);
and U8453 (N_8453,N_8254,N_8223);
xnor U8454 (N_8454,N_8277,N_8199);
or U8455 (N_8455,N_8203,N_8266);
and U8456 (N_8456,N_8186,N_8316);
or U8457 (N_8457,N_8314,N_8237);
xor U8458 (N_8458,N_8247,N_8312);
or U8459 (N_8459,N_8225,N_8168);
nand U8460 (N_8460,N_8274,N_8249);
xnor U8461 (N_8461,N_8237,N_8234);
nand U8462 (N_8462,N_8301,N_8180);
nand U8463 (N_8463,N_8204,N_8309);
or U8464 (N_8464,N_8234,N_8285);
nand U8465 (N_8465,N_8181,N_8222);
and U8466 (N_8466,N_8225,N_8221);
nand U8467 (N_8467,N_8254,N_8318);
or U8468 (N_8468,N_8234,N_8182);
and U8469 (N_8469,N_8279,N_8275);
nand U8470 (N_8470,N_8179,N_8295);
or U8471 (N_8471,N_8231,N_8236);
nand U8472 (N_8472,N_8268,N_8298);
nand U8473 (N_8473,N_8164,N_8165);
nand U8474 (N_8474,N_8221,N_8275);
nor U8475 (N_8475,N_8194,N_8290);
and U8476 (N_8476,N_8299,N_8290);
or U8477 (N_8477,N_8181,N_8185);
or U8478 (N_8478,N_8170,N_8276);
nand U8479 (N_8479,N_8185,N_8199);
nor U8480 (N_8480,N_8339,N_8379);
and U8481 (N_8481,N_8423,N_8447);
and U8482 (N_8482,N_8371,N_8393);
xor U8483 (N_8483,N_8475,N_8430);
nor U8484 (N_8484,N_8449,N_8378);
xnor U8485 (N_8485,N_8408,N_8452);
xor U8486 (N_8486,N_8437,N_8350);
nor U8487 (N_8487,N_8338,N_8381);
and U8488 (N_8488,N_8348,N_8477);
or U8489 (N_8489,N_8400,N_8335);
nor U8490 (N_8490,N_8441,N_8330);
or U8491 (N_8491,N_8389,N_8443);
nor U8492 (N_8492,N_8431,N_8427);
nor U8493 (N_8493,N_8363,N_8445);
xnor U8494 (N_8494,N_8388,N_8444);
or U8495 (N_8495,N_8356,N_8438);
nor U8496 (N_8496,N_8417,N_8352);
nand U8497 (N_8497,N_8420,N_8413);
and U8498 (N_8498,N_8377,N_8354);
or U8499 (N_8499,N_8424,N_8333);
or U8500 (N_8500,N_8332,N_8422);
nor U8501 (N_8501,N_8344,N_8395);
xor U8502 (N_8502,N_8385,N_8364);
nand U8503 (N_8503,N_8349,N_8478);
and U8504 (N_8504,N_8373,N_8347);
or U8505 (N_8505,N_8465,N_8382);
or U8506 (N_8506,N_8326,N_8345);
nand U8507 (N_8507,N_8342,N_8359);
and U8508 (N_8508,N_8426,N_8453);
nand U8509 (N_8509,N_8468,N_8450);
nand U8510 (N_8510,N_8479,N_8463);
nor U8511 (N_8511,N_8457,N_8384);
nor U8512 (N_8512,N_8451,N_8394);
nand U8513 (N_8513,N_8372,N_8414);
xor U8514 (N_8514,N_8402,N_8473);
or U8515 (N_8515,N_8460,N_8432);
or U8516 (N_8516,N_8440,N_8472);
and U8517 (N_8517,N_8397,N_8376);
nor U8518 (N_8518,N_8328,N_8458);
xnor U8519 (N_8519,N_8464,N_8419);
or U8520 (N_8520,N_8321,N_8446);
xnor U8521 (N_8521,N_8462,N_8398);
and U8522 (N_8522,N_8396,N_8329);
xnor U8523 (N_8523,N_8365,N_8405);
or U8524 (N_8524,N_8401,N_8410);
and U8525 (N_8525,N_8340,N_8366);
and U8526 (N_8526,N_8375,N_8399);
or U8527 (N_8527,N_8324,N_8411);
xor U8528 (N_8528,N_8322,N_8415);
and U8529 (N_8529,N_8407,N_8341);
and U8530 (N_8530,N_8436,N_8323);
and U8531 (N_8531,N_8362,N_8428);
and U8532 (N_8532,N_8474,N_8467);
xnor U8533 (N_8533,N_8383,N_8368);
or U8534 (N_8534,N_8421,N_8390);
xor U8535 (N_8535,N_8403,N_8331);
and U8536 (N_8536,N_8374,N_8351);
and U8537 (N_8537,N_8353,N_8459);
nand U8538 (N_8538,N_8433,N_8429);
or U8539 (N_8539,N_8392,N_8412);
or U8540 (N_8540,N_8391,N_8425);
nand U8541 (N_8541,N_8439,N_8367);
xor U8542 (N_8542,N_8325,N_8466);
xor U8543 (N_8543,N_8406,N_8469);
nand U8544 (N_8544,N_8358,N_8418);
or U8545 (N_8545,N_8386,N_8434);
and U8546 (N_8546,N_8380,N_8454);
and U8547 (N_8547,N_8387,N_8476);
and U8548 (N_8548,N_8360,N_8336);
and U8549 (N_8549,N_8320,N_8435);
or U8550 (N_8550,N_8448,N_8409);
and U8551 (N_8551,N_8346,N_8357);
nor U8552 (N_8552,N_8456,N_8361);
nand U8553 (N_8553,N_8471,N_8442);
nand U8554 (N_8554,N_8337,N_8369);
nand U8555 (N_8555,N_8370,N_8455);
nand U8556 (N_8556,N_8334,N_8470);
and U8557 (N_8557,N_8355,N_8404);
xnor U8558 (N_8558,N_8343,N_8416);
nand U8559 (N_8559,N_8461,N_8327);
xnor U8560 (N_8560,N_8331,N_8443);
or U8561 (N_8561,N_8454,N_8334);
nor U8562 (N_8562,N_8404,N_8469);
or U8563 (N_8563,N_8475,N_8382);
xor U8564 (N_8564,N_8379,N_8354);
nand U8565 (N_8565,N_8437,N_8341);
nand U8566 (N_8566,N_8321,N_8404);
or U8567 (N_8567,N_8378,N_8369);
xor U8568 (N_8568,N_8339,N_8463);
and U8569 (N_8569,N_8412,N_8433);
and U8570 (N_8570,N_8441,N_8344);
and U8571 (N_8571,N_8332,N_8348);
nor U8572 (N_8572,N_8320,N_8348);
nor U8573 (N_8573,N_8355,N_8476);
or U8574 (N_8574,N_8468,N_8365);
nand U8575 (N_8575,N_8365,N_8366);
nand U8576 (N_8576,N_8402,N_8331);
and U8577 (N_8577,N_8416,N_8407);
nor U8578 (N_8578,N_8460,N_8323);
nor U8579 (N_8579,N_8463,N_8367);
xnor U8580 (N_8580,N_8340,N_8376);
nand U8581 (N_8581,N_8403,N_8461);
or U8582 (N_8582,N_8321,N_8343);
xor U8583 (N_8583,N_8428,N_8379);
and U8584 (N_8584,N_8477,N_8440);
nand U8585 (N_8585,N_8330,N_8353);
nor U8586 (N_8586,N_8452,N_8438);
and U8587 (N_8587,N_8357,N_8409);
nor U8588 (N_8588,N_8421,N_8392);
or U8589 (N_8589,N_8424,N_8423);
xor U8590 (N_8590,N_8345,N_8426);
xor U8591 (N_8591,N_8413,N_8449);
and U8592 (N_8592,N_8460,N_8385);
xor U8593 (N_8593,N_8419,N_8411);
or U8594 (N_8594,N_8395,N_8417);
nand U8595 (N_8595,N_8467,N_8436);
nand U8596 (N_8596,N_8336,N_8386);
nand U8597 (N_8597,N_8371,N_8395);
or U8598 (N_8598,N_8471,N_8469);
and U8599 (N_8599,N_8410,N_8444);
or U8600 (N_8600,N_8401,N_8383);
nand U8601 (N_8601,N_8461,N_8348);
nor U8602 (N_8602,N_8346,N_8479);
nor U8603 (N_8603,N_8347,N_8342);
nor U8604 (N_8604,N_8352,N_8398);
nand U8605 (N_8605,N_8396,N_8386);
nand U8606 (N_8606,N_8467,N_8325);
xnor U8607 (N_8607,N_8432,N_8424);
and U8608 (N_8608,N_8381,N_8416);
nor U8609 (N_8609,N_8349,N_8325);
xnor U8610 (N_8610,N_8335,N_8449);
nor U8611 (N_8611,N_8382,N_8368);
nand U8612 (N_8612,N_8331,N_8440);
nand U8613 (N_8613,N_8417,N_8430);
xor U8614 (N_8614,N_8437,N_8337);
or U8615 (N_8615,N_8420,N_8388);
xor U8616 (N_8616,N_8394,N_8433);
nor U8617 (N_8617,N_8339,N_8455);
nand U8618 (N_8618,N_8423,N_8374);
or U8619 (N_8619,N_8428,N_8456);
nor U8620 (N_8620,N_8365,N_8453);
nor U8621 (N_8621,N_8330,N_8458);
or U8622 (N_8622,N_8478,N_8369);
or U8623 (N_8623,N_8372,N_8432);
and U8624 (N_8624,N_8450,N_8339);
or U8625 (N_8625,N_8380,N_8375);
or U8626 (N_8626,N_8424,N_8431);
nand U8627 (N_8627,N_8329,N_8478);
and U8628 (N_8628,N_8398,N_8443);
nand U8629 (N_8629,N_8422,N_8434);
or U8630 (N_8630,N_8421,N_8438);
xnor U8631 (N_8631,N_8384,N_8411);
nor U8632 (N_8632,N_8421,N_8335);
nor U8633 (N_8633,N_8397,N_8462);
and U8634 (N_8634,N_8347,N_8320);
and U8635 (N_8635,N_8474,N_8438);
and U8636 (N_8636,N_8377,N_8359);
nand U8637 (N_8637,N_8377,N_8382);
and U8638 (N_8638,N_8362,N_8475);
xor U8639 (N_8639,N_8362,N_8333);
nand U8640 (N_8640,N_8568,N_8520);
nor U8641 (N_8641,N_8517,N_8519);
xor U8642 (N_8642,N_8622,N_8589);
and U8643 (N_8643,N_8518,N_8480);
or U8644 (N_8644,N_8535,N_8626);
and U8645 (N_8645,N_8513,N_8567);
or U8646 (N_8646,N_8625,N_8538);
or U8647 (N_8647,N_8597,N_8552);
and U8648 (N_8648,N_8631,N_8491);
nor U8649 (N_8649,N_8607,N_8492);
nand U8650 (N_8650,N_8566,N_8493);
nor U8651 (N_8651,N_8541,N_8588);
nor U8652 (N_8652,N_8526,N_8634);
nor U8653 (N_8653,N_8485,N_8522);
xnor U8654 (N_8654,N_8553,N_8515);
or U8655 (N_8655,N_8636,N_8505);
or U8656 (N_8656,N_8612,N_8594);
nand U8657 (N_8657,N_8577,N_8592);
xor U8658 (N_8658,N_8586,N_8604);
and U8659 (N_8659,N_8570,N_8495);
or U8660 (N_8660,N_8621,N_8565);
or U8661 (N_8661,N_8619,N_8628);
and U8662 (N_8662,N_8534,N_8521);
and U8663 (N_8663,N_8501,N_8532);
xor U8664 (N_8664,N_8523,N_8635);
xor U8665 (N_8665,N_8638,N_8593);
nand U8666 (N_8666,N_8598,N_8563);
nand U8667 (N_8667,N_8569,N_8602);
xnor U8668 (N_8668,N_8595,N_8571);
and U8669 (N_8669,N_8527,N_8591);
nor U8670 (N_8670,N_8632,N_8606);
or U8671 (N_8671,N_8556,N_8600);
nand U8672 (N_8672,N_8536,N_8550);
and U8673 (N_8673,N_8525,N_8512);
or U8674 (N_8674,N_8530,N_8561);
xor U8675 (N_8675,N_8555,N_8544);
nand U8676 (N_8676,N_8585,N_8630);
and U8677 (N_8677,N_8564,N_8503);
and U8678 (N_8678,N_8543,N_8587);
and U8679 (N_8679,N_8610,N_8494);
and U8680 (N_8680,N_8484,N_8508);
or U8681 (N_8681,N_8509,N_8616);
nor U8682 (N_8682,N_8599,N_8539);
nor U8683 (N_8683,N_8497,N_8615);
nand U8684 (N_8684,N_8580,N_8540);
and U8685 (N_8685,N_8504,N_8579);
xnor U8686 (N_8686,N_8611,N_8605);
nand U8687 (N_8687,N_8576,N_8581);
or U8688 (N_8688,N_8537,N_8528);
xnor U8689 (N_8689,N_8608,N_8629);
nand U8690 (N_8690,N_8558,N_8637);
and U8691 (N_8691,N_8510,N_8562);
or U8692 (N_8692,N_8551,N_8627);
and U8693 (N_8693,N_8533,N_8590);
nand U8694 (N_8694,N_8488,N_8511);
and U8695 (N_8695,N_8483,N_8603);
nor U8696 (N_8696,N_8623,N_8609);
nor U8697 (N_8697,N_8531,N_8557);
and U8698 (N_8698,N_8542,N_8601);
nand U8699 (N_8699,N_8618,N_8490);
and U8700 (N_8700,N_8554,N_8506);
or U8701 (N_8701,N_8529,N_8559);
nor U8702 (N_8702,N_8547,N_8583);
xnor U8703 (N_8703,N_8507,N_8624);
nand U8704 (N_8704,N_8496,N_8524);
nand U8705 (N_8705,N_8633,N_8500);
nor U8706 (N_8706,N_8575,N_8481);
xor U8707 (N_8707,N_8578,N_8486);
xnor U8708 (N_8708,N_8514,N_8614);
nand U8709 (N_8709,N_8498,N_8499);
xnor U8710 (N_8710,N_8573,N_8584);
xnor U8711 (N_8711,N_8482,N_8582);
xor U8712 (N_8712,N_8613,N_8548);
nand U8713 (N_8713,N_8489,N_8560);
and U8714 (N_8714,N_8549,N_8620);
and U8715 (N_8715,N_8487,N_8502);
nand U8716 (N_8716,N_8639,N_8617);
nor U8717 (N_8717,N_8516,N_8572);
nand U8718 (N_8718,N_8545,N_8596);
nand U8719 (N_8719,N_8546,N_8574);
nor U8720 (N_8720,N_8545,N_8581);
nor U8721 (N_8721,N_8606,N_8626);
and U8722 (N_8722,N_8550,N_8633);
xor U8723 (N_8723,N_8637,N_8587);
and U8724 (N_8724,N_8628,N_8584);
or U8725 (N_8725,N_8563,N_8574);
or U8726 (N_8726,N_8622,N_8566);
nor U8727 (N_8727,N_8606,N_8554);
nand U8728 (N_8728,N_8630,N_8577);
xnor U8729 (N_8729,N_8542,N_8524);
and U8730 (N_8730,N_8562,N_8635);
nand U8731 (N_8731,N_8524,N_8538);
nor U8732 (N_8732,N_8493,N_8508);
xor U8733 (N_8733,N_8567,N_8629);
nor U8734 (N_8734,N_8586,N_8498);
nor U8735 (N_8735,N_8611,N_8516);
or U8736 (N_8736,N_8521,N_8597);
nand U8737 (N_8737,N_8576,N_8512);
xor U8738 (N_8738,N_8589,N_8545);
nand U8739 (N_8739,N_8501,N_8549);
and U8740 (N_8740,N_8636,N_8525);
and U8741 (N_8741,N_8541,N_8558);
nand U8742 (N_8742,N_8525,N_8571);
and U8743 (N_8743,N_8593,N_8486);
nand U8744 (N_8744,N_8639,N_8514);
xnor U8745 (N_8745,N_8558,N_8622);
nor U8746 (N_8746,N_8584,N_8572);
or U8747 (N_8747,N_8562,N_8594);
nor U8748 (N_8748,N_8499,N_8626);
or U8749 (N_8749,N_8586,N_8482);
and U8750 (N_8750,N_8595,N_8628);
xor U8751 (N_8751,N_8594,N_8544);
or U8752 (N_8752,N_8549,N_8584);
or U8753 (N_8753,N_8505,N_8491);
nand U8754 (N_8754,N_8577,N_8600);
nand U8755 (N_8755,N_8577,N_8586);
nand U8756 (N_8756,N_8580,N_8511);
xor U8757 (N_8757,N_8595,N_8489);
nand U8758 (N_8758,N_8584,N_8638);
nor U8759 (N_8759,N_8639,N_8611);
or U8760 (N_8760,N_8534,N_8582);
or U8761 (N_8761,N_8626,N_8608);
xor U8762 (N_8762,N_8587,N_8626);
xnor U8763 (N_8763,N_8617,N_8586);
and U8764 (N_8764,N_8558,N_8539);
xnor U8765 (N_8765,N_8488,N_8515);
nand U8766 (N_8766,N_8497,N_8617);
nor U8767 (N_8767,N_8548,N_8606);
and U8768 (N_8768,N_8585,N_8597);
xor U8769 (N_8769,N_8639,N_8561);
xnor U8770 (N_8770,N_8504,N_8632);
or U8771 (N_8771,N_8506,N_8556);
and U8772 (N_8772,N_8636,N_8582);
and U8773 (N_8773,N_8536,N_8579);
or U8774 (N_8774,N_8514,N_8593);
nor U8775 (N_8775,N_8617,N_8567);
nor U8776 (N_8776,N_8504,N_8558);
and U8777 (N_8777,N_8621,N_8507);
and U8778 (N_8778,N_8525,N_8608);
nor U8779 (N_8779,N_8507,N_8582);
nor U8780 (N_8780,N_8606,N_8498);
nor U8781 (N_8781,N_8577,N_8559);
or U8782 (N_8782,N_8518,N_8571);
nand U8783 (N_8783,N_8545,N_8483);
nor U8784 (N_8784,N_8592,N_8636);
nor U8785 (N_8785,N_8560,N_8483);
xor U8786 (N_8786,N_8489,N_8626);
or U8787 (N_8787,N_8633,N_8510);
or U8788 (N_8788,N_8542,N_8551);
nand U8789 (N_8789,N_8535,N_8604);
and U8790 (N_8790,N_8627,N_8542);
and U8791 (N_8791,N_8565,N_8505);
nor U8792 (N_8792,N_8575,N_8518);
xnor U8793 (N_8793,N_8554,N_8588);
or U8794 (N_8794,N_8628,N_8583);
xnor U8795 (N_8795,N_8546,N_8501);
nor U8796 (N_8796,N_8583,N_8585);
or U8797 (N_8797,N_8513,N_8580);
xnor U8798 (N_8798,N_8499,N_8514);
nor U8799 (N_8799,N_8558,N_8510);
or U8800 (N_8800,N_8643,N_8673);
xnor U8801 (N_8801,N_8739,N_8709);
xor U8802 (N_8802,N_8688,N_8648);
nor U8803 (N_8803,N_8789,N_8654);
nor U8804 (N_8804,N_8747,N_8730);
or U8805 (N_8805,N_8665,N_8794);
nor U8806 (N_8806,N_8725,N_8722);
or U8807 (N_8807,N_8732,N_8710);
nand U8808 (N_8808,N_8651,N_8678);
nand U8809 (N_8809,N_8670,N_8757);
or U8810 (N_8810,N_8715,N_8644);
nor U8811 (N_8811,N_8771,N_8679);
or U8812 (N_8812,N_8795,N_8690);
nand U8813 (N_8813,N_8772,N_8748);
nor U8814 (N_8814,N_8759,N_8787);
xnor U8815 (N_8815,N_8706,N_8749);
nand U8816 (N_8816,N_8752,N_8735);
nor U8817 (N_8817,N_8685,N_8782);
or U8818 (N_8818,N_8788,N_8741);
and U8819 (N_8819,N_8712,N_8780);
xor U8820 (N_8820,N_8658,N_8770);
or U8821 (N_8821,N_8705,N_8768);
nand U8822 (N_8822,N_8737,N_8773);
nor U8823 (N_8823,N_8761,N_8674);
nand U8824 (N_8824,N_8698,N_8704);
and U8825 (N_8825,N_8797,N_8784);
or U8826 (N_8826,N_8786,N_8720);
or U8827 (N_8827,N_8677,N_8764);
or U8828 (N_8828,N_8781,N_8796);
or U8829 (N_8829,N_8672,N_8765);
nand U8830 (N_8830,N_8776,N_8726);
or U8831 (N_8831,N_8645,N_8684);
xor U8832 (N_8832,N_8662,N_8708);
nand U8833 (N_8833,N_8640,N_8680);
or U8834 (N_8834,N_8791,N_8790);
nand U8835 (N_8835,N_8667,N_8754);
xnor U8836 (N_8836,N_8642,N_8681);
nand U8837 (N_8837,N_8655,N_8641);
and U8838 (N_8838,N_8671,N_8779);
nor U8839 (N_8839,N_8700,N_8650);
and U8840 (N_8840,N_8711,N_8734);
xor U8841 (N_8841,N_8716,N_8693);
nand U8842 (N_8842,N_8743,N_8659);
and U8843 (N_8843,N_8753,N_8703);
nor U8844 (N_8844,N_8663,N_8664);
or U8845 (N_8845,N_8668,N_8646);
and U8846 (N_8846,N_8755,N_8660);
nand U8847 (N_8847,N_8694,N_8758);
nor U8848 (N_8848,N_8717,N_8689);
nand U8849 (N_8849,N_8683,N_8652);
or U8850 (N_8850,N_8657,N_8740);
nor U8851 (N_8851,N_8774,N_8799);
nor U8852 (N_8852,N_8727,N_8778);
or U8853 (N_8853,N_8738,N_8713);
and U8854 (N_8854,N_8762,N_8783);
nor U8855 (N_8855,N_8767,N_8736);
nand U8856 (N_8856,N_8697,N_8707);
nand U8857 (N_8857,N_8675,N_8723);
or U8858 (N_8858,N_8691,N_8729);
nand U8859 (N_8859,N_8751,N_8744);
nor U8860 (N_8860,N_8721,N_8793);
nor U8861 (N_8861,N_8692,N_8647);
nand U8862 (N_8862,N_8669,N_8766);
and U8863 (N_8863,N_8745,N_8756);
xor U8864 (N_8864,N_8696,N_8719);
nor U8865 (N_8865,N_8702,N_8769);
nor U8866 (N_8866,N_8682,N_8699);
and U8867 (N_8867,N_8760,N_8656);
or U8868 (N_8868,N_8661,N_8742);
nand U8869 (N_8869,N_8763,N_8792);
nand U8870 (N_8870,N_8666,N_8777);
and U8871 (N_8871,N_8687,N_8728);
and U8872 (N_8872,N_8785,N_8686);
or U8873 (N_8873,N_8676,N_8649);
and U8874 (N_8874,N_8731,N_8746);
nor U8875 (N_8875,N_8733,N_8798);
xnor U8876 (N_8876,N_8695,N_8653);
or U8877 (N_8877,N_8724,N_8718);
nor U8878 (N_8878,N_8701,N_8775);
xor U8879 (N_8879,N_8714,N_8750);
nor U8880 (N_8880,N_8705,N_8747);
and U8881 (N_8881,N_8740,N_8729);
xor U8882 (N_8882,N_8682,N_8642);
and U8883 (N_8883,N_8640,N_8681);
and U8884 (N_8884,N_8720,N_8789);
or U8885 (N_8885,N_8740,N_8786);
and U8886 (N_8886,N_8775,N_8679);
xor U8887 (N_8887,N_8728,N_8699);
nor U8888 (N_8888,N_8740,N_8767);
nand U8889 (N_8889,N_8721,N_8677);
and U8890 (N_8890,N_8753,N_8771);
nor U8891 (N_8891,N_8703,N_8718);
xor U8892 (N_8892,N_8751,N_8731);
nor U8893 (N_8893,N_8751,N_8661);
or U8894 (N_8894,N_8678,N_8774);
nor U8895 (N_8895,N_8730,N_8714);
nor U8896 (N_8896,N_8788,N_8686);
nor U8897 (N_8897,N_8782,N_8789);
and U8898 (N_8898,N_8738,N_8675);
nor U8899 (N_8899,N_8679,N_8758);
or U8900 (N_8900,N_8708,N_8742);
and U8901 (N_8901,N_8764,N_8650);
xnor U8902 (N_8902,N_8695,N_8715);
nor U8903 (N_8903,N_8683,N_8709);
xnor U8904 (N_8904,N_8699,N_8730);
xnor U8905 (N_8905,N_8694,N_8677);
or U8906 (N_8906,N_8646,N_8643);
nor U8907 (N_8907,N_8743,N_8752);
or U8908 (N_8908,N_8788,N_8702);
and U8909 (N_8909,N_8706,N_8733);
and U8910 (N_8910,N_8696,N_8756);
or U8911 (N_8911,N_8689,N_8735);
or U8912 (N_8912,N_8798,N_8693);
nand U8913 (N_8913,N_8690,N_8659);
nor U8914 (N_8914,N_8781,N_8765);
and U8915 (N_8915,N_8657,N_8789);
nand U8916 (N_8916,N_8769,N_8663);
xnor U8917 (N_8917,N_8758,N_8790);
or U8918 (N_8918,N_8705,N_8689);
nand U8919 (N_8919,N_8709,N_8742);
nand U8920 (N_8920,N_8703,N_8735);
nand U8921 (N_8921,N_8751,N_8735);
or U8922 (N_8922,N_8646,N_8736);
and U8923 (N_8923,N_8678,N_8740);
nor U8924 (N_8924,N_8698,N_8746);
and U8925 (N_8925,N_8744,N_8677);
nor U8926 (N_8926,N_8744,N_8781);
xor U8927 (N_8927,N_8661,N_8687);
xor U8928 (N_8928,N_8764,N_8673);
nand U8929 (N_8929,N_8716,N_8744);
or U8930 (N_8930,N_8699,N_8674);
or U8931 (N_8931,N_8753,N_8724);
xnor U8932 (N_8932,N_8643,N_8765);
and U8933 (N_8933,N_8716,N_8752);
xor U8934 (N_8934,N_8784,N_8751);
and U8935 (N_8935,N_8684,N_8705);
or U8936 (N_8936,N_8698,N_8691);
xor U8937 (N_8937,N_8786,N_8657);
nand U8938 (N_8938,N_8670,N_8766);
nand U8939 (N_8939,N_8760,N_8726);
or U8940 (N_8940,N_8749,N_8686);
and U8941 (N_8941,N_8670,N_8688);
nand U8942 (N_8942,N_8724,N_8653);
or U8943 (N_8943,N_8700,N_8688);
nand U8944 (N_8944,N_8784,N_8768);
xnor U8945 (N_8945,N_8791,N_8733);
xor U8946 (N_8946,N_8672,N_8788);
xnor U8947 (N_8947,N_8758,N_8798);
and U8948 (N_8948,N_8719,N_8720);
nor U8949 (N_8949,N_8712,N_8701);
or U8950 (N_8950,N_8773,N_8724);
or U8951 (N_8951,N_8765,N_8746);
and U8952 (N_8952,N_8699,N_8676);
or U8953 (N_8953,N_8790,N_8667);
and U8954 (N_8954,N_8720,N_8740);
or U8955 (N_8955,N_8721,N_8709);
or U8956 (N_8956,N_8727,N_8687);
or U8957 (N_8957,N_8727,N_8690);
and U8958 (N_8958,N_8787,N_8714);
nor U8959 (N_8959,N_8778,N_8669);
xor U8960 (N_8960,N_8914,N_8806);
xnor U8961 (N_8961,N_8803,N_8910);
or U8962 (N_8962,N_8928,N_8872);
or U8963 (N_8963,N_8802,N_8925);
xnor U8964 (N_8964,N_8952,N_8901);
xor U8965 (N_8965,N_8862,N_8844);
nand U8966 (N_8966,N_8883,N_8935);
or U8967 (N_8967,N_8851,N_8959);
and U8968 (N_8968,N_8827,N_8801);
or U8969 (N_8969,N_8907,N_8825);
or U8970 (N_8970,N_8930,N_8813);
nand U8971 (N_8971,N_8889,N_8831);
nand U8972 (N_8972,N_8919,N_8846);
nand U8973 (N_8973,N_8835,N_8882);
xor U8974 (N_8974,N_8954,N_8957);
or U8975 (N_8975,N_8843,N_8874);
or U8976 (N_8976,N_8847,N_8824);
nand U8977 (N_8977,N_8865,N_8921);
and U8978 (N_8978,N_8892,N_8854);
and U8979 (N_8979,N_8924,N_8871);
xnor U8980 (N_8980,N_8936,N_8842);
and U8981 (N_8981,N_8927,N_8819);
xor U8982 (N_8982,N_8867,N_8911);
xnor U8983 (N_8983,N_8884,N_8855);
xor U8984 (N_8984,N_8894,N_8948);
or U8985 (N_8985,N_8893,N_8931);
nor U8986 (N_8986,N_8941,N_8933);
and U8987 (N_8987,N_8923,N_8800);
and U8988 (N_8988,N_8953,N_8908);
nand U8989 (N_8989,N_8885,N_8869);
nand U8990 (N_8990,N_8856,N_8913);
nor U8991 (N_8991,N_8958,N_8860);
xnor U8992 (N_8992,N_8906,N_8934);
and U8993 (N_8993,N_8840,N_8942);
nor U8994 (N_8994,N_8956,N_8838);
nor U8995 (N_8995,N_8810,N_8861);
nand U8996 (N_8996,N_8903,N_8822);
xor U8997 (N_8997,N_8818,N_8805);
and U8998 (N_8998,N_8951,N_8809);
nor U8999 (N_8999,N_8826,N_8937);
and U9000 (N_9000,N_8857,N_8904);
nor U9001 (N_9001,N_8900,N_8898);
nor U9002 (N_9002,N_8859,N_8940);
nor U9003 (N_9003,N_8881,N_8852);
nor U9004 (N_9004,N_8929,N_8814);
nand U9005 (N_9005,N_8864,N_8938);
xor U9006 (N_9006,N_8834,N_8946);
nor U9007 (N_9007,N_8915,N_8902);
and U9008 (N_9008,N_8916,N_8823);
xor U9009 (N_9009,N_8876,N_8870);
and U9010 (N_9010,N_8899,N_8815);
xor U9011 (N_9011,N_8841,N_8812);
and U9012 (N_9012,N_8879,N_8897);
xnor U9013 (N_9013,N_8820,N_8947);
nand U9014 (N_9014,N_8829,N_8895);
or U9015 (N_9015,N_8804,N_8890);
nor U9016 (N_9016,N_8886,N_8853);
and U9017 (N_9017,N_8950,N_8873);
or U9018 (N_9018,N_8909,N_8830);
or U9019 (N_9019,N_8807,N_8922);
nor U9020 (N_9020,N_8905,N_8808);
or U9021 (N_9021,N_8868,N_8863);
nor U9022 (N_9022,N_8888,N_8949);
or U9023 (N_9023,N_8817,N_8821);
or U9024 (N_9024,N_8891,N_8836);
nor U9025 (N_9025,N_8832,N_8887);
xor U9026 (N_9026,N_8858,N_8926);
and U9027 (N_9027,N_8816,N_8918);
or U9028 (N_9028,N_8880,N_8943);
nor U9029 (N_9029,N_8811,N_8837);
and U9030 (N_9030,N_8920,N_8875);
xnor U9031 (N_9031,N_8917,N_8944);
or U9032 (N_9032,N_8848,N_8877);
nand U9033 (N_9033,N_8850,N_8945);
and U9034 (N_9034,N_8912,N_8896);
nand U9035 (N_9035,N_8878,N_8839);
xnor U9036 (N_9036,N_8932,N_8955);
or U9037 (N_9037,N_8939,N_8866);
nand U9038 (N_9038,N_8849,N_8845);
nor U9039 (N_9039,N_8833,N_8828);
nor U9040 (N_9040,N_8864,N_8942);
or U9041 (N_9041,N_8936,N_8901);
nand U9042 (N_9042,N_8916,N_8818);
nand U9043 (N_9043,N_8958,N_8807);
xor U9044 (N_9044,N_8876,N_8889);
nand U9045 (N_9045,N_8889,N_8919);
or U9046 (N_9046,N_8837,N_8805);
or U9047 (N_9047,N_8890,N_8854);
or U9048 (N_9048,N_8881,N_8903);
nand U9049 (N_9049,N_8947,N_8802);
xnor U9050 (N_9050,N_8809,N_8835);
nor U9051 (N_9051,N_8943,N_8848);
nor U9052 (N_9052,N_8904,N_8894);
xnor U9053 (N_9053,N_8945,N_8946);
xor U9054 (N_9054,N_8819,N_8863);
nor U9055 (N_9055,N_8911,N_8944);
nor U9056 (N_9056,N_8804,N_8874);
xnor U9057 (N_9057,N_8918,N_8837);
xnor U9058 (N_9058,N_8848,N_8827);
and U9059 (N_9059,N_8837,N_8928);
xnor U9060 (N_9060,N_8857,N_8861);
or U9061 (N_9061,N_8810,N_8883);
nor U9062 (N_9062,N_8893,N_8891);
and U9063 (N_9063,N_8801,N_8814);
nand U9064 (N_9064,N_8933,N_8813);
and U9065 (N_9065,N_8885,N_8917);
or U9066 (N_9066,N_8935,N_8810);
nor U9067 (N_9067,N_8884,N_8836);
xor U9068 (N_9068,N_8847,N_8901);
nor U9069 (N_9069,N_8928,N_8932);
xor U9070 (N_9070,N_8809,N_8813);
nor U9071 (N_9071,N_8822,N_8843);
and U9072 (N_9072,N_8814,N_8940);
nor U9073 (N_9073,N_8958,N_8853);
nor U9074 (N_9074,N_8813,N_8871);
nand U9075 (N_9075,N_8933,N_8854);
and U9076 (N_9076,N_8904,N_8919);
xor U9077 (N_9077,N_8832,N_8958);
or U9078 (N_9078,N_8957,N_8883);
nor U9079 (N_9079,N_8900,N_8840);
nor U9080 (N_9080,N_8947,N_8844);
or U9081 (N_9081,N_8806,N_8916);
or U9082 (N_9082,N_8858,N_8819);
and U9083 (N_9083,N_8863,N_8878);
nor U9084 (N_9084,N_8927,N_8836);
nand U9085 (N_9085,N_8856,N_8904);
nor U9086 (N_9086,N_8958,N_8884);
nor U9087 (N_9087,N_8844,N_8875);
nor U9088 (N_9088,N_8848,N_8950);
nor U9089 (N_9089,N_8882,N_8934);
nor U9090 (N_9090,N_8876,N_8820);
nand U9091 (N_9091,N_8835,N_8808);
or U9092 (N_9092,N_8902,N_8943);
nand U9093 (N_9093,N_8816,N_8934);
xnor U9094 (N_9094,N_8841,N_8843);
and U9095 (N_9095,N_8931,N_8896);
nand U9096 (N_9096,N_8881,N_8814);
xor U9097 (N_9097,N_8956,N_8850);
and U9098 (N_9098,N_8812,N_8851);
and U9099 (N_9099,N_8935,N_8899);
xnor U9100 (N_9100,N_8894,N_8839);
nor U9101 (N_9101,N_8861,N_8905);
nor U9102 (N_9102,N_8813,N_8957);
xor U9103 (N_9103,N_8890,N_8871);
or U9104 (N_9104,N_8882,N_8838);
nand U9105 (N_9105,N_8942,N_8911);
nand U9106 (N_9106,N_8817,N_8935);
nand U9107 (N_9107,N_8834,N_8890);
nor U9108 (N_9108,N_8852,N_8885);
and U9109 (N_9109,N_8843,N_8913);
or U9110 (N_9110,N_8896,N_8858);
nand U9111 (N_9111,N_8803,N_8959);
or U9112 (N_9112,N_8889,N_8950);
or U9113 (N_9113,N_8947,N_8849);
nand U9114 (N_9114,N_8926,N_8949);
nand U9115 (N_9115,N_8820,N_8918);
or U9116 (N_9116,N_8900,N_8885);
or U9117 (N_9117,N_8945,N_8930);
and U9118 (N_9118,N_8869,N_8835);
xor U9119 (N_9119,N_8931,N_8885);
or U9120 (N_9120,N_9045,N_9030);
and U9121 (N_9121,N_9068,N_9050);
nand U9122 (N_9122,N_9061,N_9076);
and U9123 (N_9123,N_9115,N_9042);
xnor U9124 (N_9124,N_9102,N_9022);
and U9125 (N_9125,N_9037,N_9017);
or U9126 (N_9126,N_9097,N_9053);
xor U9127 (N_9127,N_9048,N_9019);
or U9128 (N_9128,N_8975,N_9101);
nand U9129 (N_9129,N_8996,N_9106);
and U9130 (N_9130,N_9078,N_9012);
or U9131 (N_9131,N_8967,N_9031);
and U9132 (N_9132,N_9040,N_8984);
and U9133 (N_9133,N_9103,N_9059);
nor U9134 (N_9134,N_8974,N_8982);
nor U9135 (N_9135,N_8976,N_9085);
nor U9136 (N_9136,N_9046,N_9054);
and U9137 (N_9137,N_9036,N_9070);
nor U9138 (N_9138,N_9077,N_8962);
and U9139 (N_9139,N_8973,N_9038);
and U9140 (N_9140,N_9075,N_9058);
nor U9141 (N_9141,N_8979,N_9113);
nor U9142 (N_9142,N_9000,N_8970);
or U9143 (N_9143,N_9009,N_9079);
xor U9144 (N_9144,N_8988,N_9082);
nor U9145 (N_9145,N_9024,N_9013);
xnor U9146 (N_9146,N_8999,N_9107);
nand U9147 (N_9147,N_8990,N_9057);
and U9148 (N_9148,N_9092,N_9096);
xnor U9149 (N_9149,N_9032,N_9065);
nor U9150 (N_9150,N_9015,N_9035);
nor U9151 (N_9151,N_9091,N_9027);
or U9152 (N_9152,N_9008,N_9081);
xnor U9153 (N_9153,N_8977,N_9087);
nor U9154 (N_9154,N_8992,N_9062);
and U9155 (N_9155,N_9117,N_9071);
nor U9156 (N_9156,N_8994,N_9016);
nor U9157 (N_9157,N_9086,N_9014);
nor U9158 (N_9158,N_9100,N_9025);
xor U9159 (N_9159,N_9110,N_9011);
or U9160 (N_9160,N_8991,N_9029);
or U9161 (N_9161,N_9063,N_9119);
xnor U9162 (N_9162,N_8972,N_9010);
nand U9163 (N_9163,N_8985,N_8987);
xnor U9164 (N_9164,N_8995,N_9033);
nand U9165 (N_9165,N_9051,N_8983);
nor U9166 (N_9166,N_9023,N_9034);
or U9167 (N_9167,N_9114,N_9064);
xnor U9168 (N_9168,N_8998,N_9018);
and U9169 (N_9169,N_9111,N_9060);
and U9170 (N_9170,N_9002,N_8960);
or U9171 (N_9171,N_9007,N_9108);
xor U9172 (N_9172,N_8971,N_9044);
nor U9173 (N_9173,N_8969,N_9028);
or U9174 (N_9174,N_9093,N_9067);
xnor U9175 (N_9175,N_9026,N_9047);
or U9176 (N_9176,N_9083,N_9005);
nor U9177 (N_9177,N_9041,N_8993);
nor U9178 (N_9178,N_9069,N_9074);
nand U9179 (N_9179,N_9020,N_9109);
or U9180 (N_9180,N_9056,N_8981);
nor U9181 (N_9181,N_9049,N_9094);
or U9182 (N_9182,N_8997,N_9089);
xnor U9183 (N_9183,N_9099,N_9001);
or U9184 (N_9184,N_8961,N_9043);
nand U9185 (N_9185,N_9080,N_9055);
xor U9186 (N_9186,N_9104,N_8965);
or U9187 (N_9187,N_9116,N_8968);
or U9188 (N_9188,N_9090,N_8989);
xnor U9189 (N_9189,N_9006,N_9021);
nor U9190 (N_9190,N_9039,N_9084);
and U9191 (N_9191,N_8978,N_9105);
xor U9192 (N_9192,N_8980,N_9066);
nor U9193 (N_9193,N_8966,N_8964);
and U9194 (N_9194,N_9052,N_8963);
or U9195 (N_9195,N_9088,N_9072);
nand U9196 (N_9196,N_9004,N_9095);
xnor U9197 (N_9197,N_9073,N_9118);
and U9198 (N_9198,N_9003,N_8986);
nor U9199 (N_9199,N_9112,N_9098);
and U9200 (N_9200,N_9058,N_8985);
nor U9201 (N_9201,N_9107,N_9077);
nand U9202 (N_9202,N_9113,N_9017);
xnor U9203 (N_9203,N_9077,N_8967);
or U9204 (N_9204,N_8998,N_8960);
xor U9205 (N_9205,N_9111,N_9092);
or U9206 (N_9206,N_9051,N_9008);
nand U9207 (N_9207,N_9011,N_9067);
xnor U9208 (N_9208,N_9004,N_8979);
nor U9209 (N_9209,N_8976,N_9003);
nor U9210 (N_9210,N_9028,N_9064);
nand U9211 (N_9211,N_8992,N_8981);
nand U9212 (N_9212,N_9027,N_9083);
xor U9213 (N_9213,N_8983,N_9020);
or U9214 (N_9214,N_9111,N_9059);
nor U9215 (N_9215,N_9025,N_8981);
nand U9216 (N_9216,N_9115,N_9060);
or U9217 (N_9217,N_9009,N_9005);
or U9218 (N_9218,N_9029,N_9075);
and U9219 (N_9219,N_8967,N_9013);
or U9220 (N_9220,N_8964,N_9030);
xor U9221 (N_9221,N_9010,N_9103);
nand U9222 (N_9222,N_9071,N_9115);
nand U9223 (N_9223,N_9035,N_9077);
nor U9224 (N_9224,N_9052,N_8985);
and U9225 (N_9225,N_9088,N_9001);
and U9226 (N_9226,N_9071,N_9066);
nand U9227 (N_9227,N_8997,N_9026);
or U9228 (N_9228,N_9020,N_9054);
nor U9229 (N_9229,N_8983,N_9047);
or U9230 (N_9230,N_9108,N_8965);
or U9231 (N_9231,N_9018,N_9000);
nor U9232 (N_9232,N_9009,N_9002);
and U9233 (N_9233,N_9114,N_9075);
xor U9234 (N_9234,N_8993,N_8983);
nor U9235 (N_9235,N_9117,N_8983);
nand U9236 (N_9236,N_9035,N_8996);
nor U9237 (N_9237,N_9061,N_9046);
nand U9238 (N_9238,N_8969,N_9118);
or U9239 (N_9239,N_9063,N_9057);
nor U9240 (N_9240,N_9009,N_9044);
nor U9241 (N_9241,N_9073,N_8977);
or U9242 (N_9242,N_9092,N_8984);
nor U9243 (N_9243,N_9059,N_9113);
nor U9244 (N_9244,N_9095,N_8969);
or U9245 (N_9245,N_9048,N_8980);
xnor U9246 (N_9246,N_9004,N_9093);
xor U9247 (N_9247,N_9012,N_8999);
nor U9248 (N_9248,N_8985,N_9014);
nor U9249 (N_9249,N_9077,N_9117);
and U9250 (N_9250,N_8996,N_9094);
or U9251 (N_9251,N_9089,N_9063);
or U9252 (N_9252,N_9055,N_8970);
nand U9253 (N_9253,N_9088,N_8984);
or U9254 (N_9254,N_9090,N_9017);
nand U9255 (N_9255,N_9074,N_8961);
nand U9256 (N_9256,N_9076,N_9018);
and U9257 (N_9257,N_9019,N_9068);
nand U9258 (N_9258,N_9039,N_8973);
and U9259 (N_9259,N_8992,N_9093);
xnor U9260 (N_9260,N_9008,N_9113);
nor U9261 (N_9261,N_9019,N_9009);
nor U9262 (N_9262,N_9065,N_8973);
and U9263 (N_9263,N_9032,N_9106);
and U9264 (N_9264,N_9098,N_8972);
nor U9265 (N_9265,N_9072,N_8968);
nor U9266 (N_9266,N_9011,N_9094);
xor U9267 (N_9267,N_9011,N_9033);
nor U9268 (N_9268,N_9019,N_9101);
or U9269 (N_9269,N_9078,N_8972);
xnor U9270 (N_9270,N_9094,N_9009);
or U9271 (N_9271,N_8984,N_9107);
nand U9272 (N_9272,N_9032,N_9080);
nor U9273 (N_9273,N_9024,N_9111);
or U9274 (N_9274,N_8992,N_9102);
and U9275 (N_9275,N_9046,N_9119);
or U9276 (N_9276,N_9100,N_9059);
nand U9277 (N_9277,N_9066,N_9025);
nor U9278 (N_9278,N_9114,N_9023);
nand U9279 (N_9279,N_9067,N_9051);
or U9280 (N_9280,N_9221,N_9148);
or U9281 (N_9281,N_9263,N_9219);
xnor U9282 (N_9282,N_9246,N_9279);
and U9283 (N_9283,N_9211,N_9226);
xnor U9284 (N_9284,N_9169,N_9201);
xor U9285 (N_9285,N_9171,N_9196);
or U9286 (N_9286,N_9218,N_9165);
nor U9287 (N_9287,N_9262,N_9124);
and U9288 (N_9288,N_9158,N_9257);
xor U9289 (N_9289,N_9247,N_9276);
or U9290 (N_9290,N_9224,N_9238);
xnor U9291 (N_9291,N_9248,N_9233);
xnor U9292 (N_9292,N_9156,N_9144);
xor U9293 (N_9293,N_9191,N_9130);
or U9294 (N_9294,N_9265,N_9155);
nor U9295 (N_9295,N_9222,N_9195);
nand U9296 (N_9296,N_9188,N_9183);
or U9297 (N_9297,N_9208,N_9261);
nor U9298 (N_9298,N_9167,N_9234);
xor U9299 (N_9299,N_9204,N_9227);
or U9300 (N_9300,N_9128,N_9239);
nor U9301 (N_9301,N_9244,N_9176);
nand U9302 (N_9302,N_9228,N_9223);
and U9303 (N_9303,N_9185,N_9152);
or U9304 (N_9304,N_9267,N_9189);
and U9305 (N_9305,N_9172,N_9162);
or U9306 (N_9306,N_9166,N_9243);
nor U9307 (N_9307,N_9139,N_9136);
nand U9308 (N_9308,N_9255,N_9236);
xor U9309 (N_9309,N_9142,N_9134);
nor U9310 (N_9310,N_9123,N_9121);
xor U9311 (N_9311,N_9249,N_9140);
nor U9312 (N_9312,N_9174,N_9251);
nor U9313 (N_9313,N_9203,N_9151);
or U9314 (N_9314,N_9120,N_9275);
nor U9315 (N_9315,N_9192,N_9154);
nand U9316 (N_9316,N_9153,N_9206);
xnor U9317 (N_9317,N_9256,N_9168);
and U9318 (N_9318,N_9181,N_9150);
xor U9319 (N_9319,N_9202,N_9160);
and U9320 (N_9320,N_9235,N_9197);
nor U9321 (N_9321,N_9273,N_9159);
and U9322 (N_9322,N_9164,N_9253);
or U9323 (N_9323,N_9241,N_9180);
nor U9324 (N_9324,N_9259,N_9175);
nor U9325 (N_9325,N_9250,N_9271);
xor U9326 (N_9326,N_9240,N_9252);
xnor U9327 (N_9327,N_9210,N_9245);
xor U9328 (N_9328,N_9200,N_9272);
nor U9329 (N_9329,N_9135,N_9264);
nor U9330 (N_9330,N_9242,N_9141);
or U9331 (N_9331,N_9237,N_9230);
and U9332 (N_9332,N_9173,N_9170);
xor U9333 (N_9333,N_9122,N_9187);
or U9334 (N_9334,N_9198,N_9199);
xnor U9335 (N_9335,N_9186,N_9231);
and U9336 (N_9336,N_9277,N_9138);
nand U9337 (N_9337,N_9129,N_9225);
nand U9338 (N_9338,N_9149,N_9214);
xor U9339 (N_9339,N_9145,N_9126);
nor U9340 (N_9340,N_9179,N_9207);
xor U9341 (N_9341,N_9157,N_9127);
nand U9342 (N_9342,N_9270,N_9209);
or U9343 (N_9343,N_9274,N_9163);
nand U9344 (N_9344,N_9215,N_9133);
xor U9345 (N_9345,N_9177,N_9132);
nand U9346 (N_9346,N_9178,N_9125);
xor U9347 (N_9347,N_9278,N_9190);
and U9348 (N_9348,N_9182,N_9212);
xnor U9349 (N_9349,N_9131,N_9232);
xor U9350 (N_9350,N_9258,N_9147);
nand U9351 (N_9351,N_9229,N_9194);
nand U9352 (N_9352,N_9266,N_9184);
and U9353 (N_9353,N_9143,N_9268);
or U9354 (N_9354,N_9193,N_9213);
nor U9355 (N_9355,N_9161,N_9216);
or U9356 (N_9356,N_9254,N_9205);
xnor U9357 (N_9357,N_9260,N_9220);
and U9358 (N_9358,N_9137,N_9217);
xnor U9359 (N_9359,N_9269,N_9146);
nor U9360 (N_9360,N_9134,N_9158);
or U9361 (N_9361,N_9165,N_9259);
xor U9362 (N_9362,N_9207,N_9180);
nor U9363 (N_9363,N_9232,N_9165);
nor U9364 (N_9364,N_9254,N_9195);
or U9365 (N_9365,N_9141,N_9213);
xor U9366 (N_9366,N_9240,N_9243);
xor U9367 (N_9367,N_9256,N_9156);
or U9368 (N_9368,N_9210,N_9257);
or U9369 (N_9369,N_9218,N_9278);
nor U9370 (N_9370,N_9120,N_9277);
and U9371 (N_9371,N_9262,N_9223);
or U9372 (N_9372,N_9265,N_9223);
and U9373 (N_9373,N_9189,N_9152);
nor U9374 (N_9374,N_9222,N_9146);
and U9375 (N_9375,N_9237,N_9204);
or U9376 (N_9376,N_9195,N_9152);
xor U9377 (N_9377,N_9191,N_9277);
xor U9378 (N_9378,N_9211,N_9215);
nor U9379 (N_9379,N_9141,N_9134);
and U9380 (N_9380,N_9247,N_9218);
xor U9381 (N_9381,N_9183,N_9185);
and U9382 (N_9382,N_9143,N_9180);
nand U9383 (N_9383,N_9255,N_9140);
and U9384 (N_9384,N_9259,N_9219);
nand U9385 (N_9385,N_9251,N_9209);
nor U9386 (N_9386,N_9199,N_9219);
or U9387 (N_9387,N_9156,N_9236);
or U9388 (N_9388,N_9248,N_9270);
nor U9389 (N_9389,N_9192,N_9221);
and U9390 (N_9390,N_9212,N_9259);
nand U9391 (N_9391,N_9273,N_9160);
nor U9392 (N_9392,N_9159,N_9123);
or U9393 (N_9393,N_9147,N_9202);
nand U9394 (N_9394,N_9133,N_9176);
xor U9395 (N_9395,N_9200,N_9223);
nand U9396 (N_9396,N_9216,N_9179);
and U9397 (N_9397,N_9147,N_9236);
or U9398 (N_9398,N_9245,N_9223);
nand U9399 (N_9399,N_9217,N_9232);
nand U9400 (N_9400,N_9235,N_9160);
and U9401 (N_9401,N_9192,N_9273);
or U9402 (N_9402,N_9217,N_9188);
and U9403 (N_9403,N_9186,N_9160);
nor U9404 (N_9404,N_9241,N_9246);
xnor U9405 (N_9405,N_9149,N_9145);
and U9406 (N_9406,N_9211,N_9212);
xor U9407 (N_9407,N_9184,N_9176);
xnor U9408 (N_9408,N_9232,N_9230);
nor U9409 (N_9409,N_9270,N_9259);
or U9410 (N_9410,N_9140,N_9243);
and U9411 (N_9411,N_9192,N_9257);
xnor U9412 (N_9412,N_9124,N_9213);
xnor U9413 (N_9413,N_9175,N_9215);
and U9414 (N_9414,N_9123,N_9170);
and U9415 (N_9415,N_9153,N_9185);
nor U9416 (N_9416,N_9181,N_9205);
nor U9417 (N_9417,N_9179,N_9213);
nand U9418 (N_9418,N_9212,N_9276);
nor U9419 (N_9419,N_9169,N_9218);
or U9420 (N_9420,N_9218,N_9152);
and U9421 (N_9421,N_9245,N_9179);
nand U9422 (N_9422,N_9159,N_9232);
xnor U9423 (N_9423,N_9199,N_9277);
xor U9424 (N_9424,N_9155,N_9159);
nor U9425 (N_9425,N_9184,N_9211);
nand U9426 (N_9426,N_9152,N_9233);
nor U9427 (N_9427,N_9212,N_9181);
nand U9428 (N_9428,N_9146,N_9155);
nand U9429 (N_9429,N_9186,N_9168);
and U9430 (N_9430,N_9160,N_9278);
nand U9431 (N_9431,N_9122,N_9169);
and U9432 (N_9432,N_9203,N_9243);
and U9433 (N_9433,N_9191,N_9178);
xor U9434 (N_9434,N_9255,N_9273);
nand U9435 (N_9435,N_9146,N_9262);
or U9436 (N_9436,N_9123,N_9133);
xnor U9437 (N_9437,N_9232,N_9129);
nor U9438 (N_9438,N_9130,N_9202);
nand U9439 (N_9439,N_9138,N_9249);
and U9440 (N_9440,N_9324,N_9430);
nor U9441 (N_9441,N_9365,N_9347);
or U9442 (N_9442,N_9287,N_9286);
nor U9443 (N_9443,N_9431,N_9320);
nor U9444 (N_9444,N_9295,N_9400);
nand U9445 (N_9445,N_9407,N_9392);
nand U9446 (N_9446,N_9304,N_9396);
nand U9447 (N_9447,N_9360,N_9427);
xnor U9448 (N_9448,N_9391,N_9294);
and U9449 (N_9449,N_9351,N_9372);
nand U9450 (N_9450,N_9305,N_9301);
nand U9451 (N_9451,N_9422,N_9423);
and U9452 (N_9452,N_9327,N_9373);
and U9453 (N_9453,N_9385,N_9388);
nor U9454 (N_9454,N_9299,N_9376);
nand U9455 (N_9455,N_9420,N_9429);
and U9456 (N_9456,N_9436,N_9367);
and U9457 (N_9457,N_9408,N_9426);
nand U9458 (N_9458,N_9318,N_9352);
and U9459 (N_9459,N_9290,N_9355);
or U9460 (N_9460,N_9433,N_9383);
and U9461 (N_9461,N_9283,N_9411);
nand U9462 (N_9462,N_9316,N_9415);
nor U9463 (N_9463,N_9343,N_9369);
or U9464 (N_9464,N_9394,N_9379);
and U9465 (N_9465,N_9371,N_9425);
xnor U9466 (N_9466,N_9358,N_9406);
and U9467 (N_9467,N_9311,N_9280);
or U9468 (N_9468,N_9418,N_9409);
nor U9469 (N_9469,N_9310,N_9337);
or U9470 (N_9470,N_9300,N_9325);
xor U9471 (N_9471,N_9346,N_9378);
xor U9472 (N_9472,N_9281,N_9289);
xor U9473 (N_9473,N_9306,N_9307);
or U9474 (N_9474,N_9326,N_9417);
or U9475 (N_9475,N_9357,N_9313);
nor U9476 (N_9476,N_9363,N_9416);
and U9477 (N_9477,N_9292,N_9303);
nand U9478 (N_9478,N_9332,N_9368);
or U9479 (N_9479,N_9359,N_9366);
and U9480 (N_9480,N_9288,N_9317);
nor U9481 (N_9481,N_9386,N_9336);
and U9482 (N_9482,N_9323,N_9319);
and U9483 (N_9483,N_9342,N_9398);
or U9484 (N_9484,N_9393,N_9348);
xnor U9485 (N_9485,N_9395,N_9381);
or U9486 (N_9486,N_9302,N_9361);
or U9487 (N_9487,N_9329,N_9282);
nand U9488 (N_9488,N_9437,N_9345);
nor U9489 (N_9489,N_9382,N_9374);
and U9490 (N_9490,N_9370,N_9315);
or U9491 (N_9491,N_9375,N_9403);
nor U9492 (N_9492,N_9434,N_9405);
or U9493 (N_9493,N_9341,N_9297);
or U9494 (N_9494,N_9414,N_9291);
and U9495 (N_9495,N_9404,N_9389);
and U9496 (N_9496,N_9384,N_9293);
nand U9497 (N_9497,N_9328,N_9333);
nor U9498 (N_9498,N_9312,N_9432);
nor U9499 (N_9499,N_9338,N_9334);
xnor U9500 (N_9500,N_9339,N_9439);
or U9501 (N_9501,N_9410,N_9335);
xnor U9502 (N_9502,N_9331,N_9438);
nand U9503 (N_9503,N_9309,N_9421);
nand U9504 (N_9504,N_9321,N_9399);
nand U9505 (N_9505,N_9364,N_9284);
nand U9506 (N_9506,N_9377,N_9296);
nand U9507 (N_9507,N_9314,N_9387);
or U9508 (N_9508,N_9344,N_9308);
xnor U9509 (N_9509,N_9397,N_9380);
and U9510 (N_9510,N_9356,N_9330);
or U9511 (N_9511,N_9285,N_9322);
and U9512 (N_9512,N_9362,N_9340);
and U9513 (N_9513,N_9412,N_9350);
nand U9514 (N_9514,N_9349,N_9401);
and U9515 (N_9515,N_9435,N_9354);
nor U9516 (N_9516,N_9424,N_9402);
nor U9517 (N_9517,N_9413,N_9419);
nand U9518 (N_9518,N_9353,N_9428);
nand U9519 (N_9519,N_9298,N_9390);
or U9520 (N_9520,N_9307,N_9350);
and U9521 (N_9521,N_9315,N_9355);
nor U9522 (N_9522,N_9349,N_9302);
and U9523 (N_9523,N_9301,N_9431);
or U9524 (N_9524,N_9373,N_9387);
and U9525 (N_9525,N_9356,N_9296);
xnor U9526 (N_9526,N_9420,N_9377);
and U9527 (N_9527,N_9439,N_9300);
or U9528 (N_9528,N_9284,N_9351);
and U9529 (N_9529,N_9327,N_9314);
or U9530 (N_9530,N_9398,N_9344);
nor U9531 (N_9531,N_9388,N_9353);
nand U9532 (N_9532,N_9432,N_9346);
and U9533 (N_9533,N_9392,N_9314);
xnor U9534 (N_9534,N_9295,N_9365);
or U9535 (N_9535,N_9423,N_9376);
and U9536 (N_9536,N_9428,N_9378);
nor U9537 (N_9537,N_9343,N_9335);
or U9538 (N_9538,N_9350,N_9389);
and U9539 (N_9539,N_9381,N_9424);
nor U9540 (N_9540,N_9401,N_9296);
nor U9541 (N_9541,N_9378,N_9411);
xnor U9542 (N_9542,N_9415,N_9356);
xor U9543 (N_9543,N_9379,N_9407);
nand U9544 (N_9544,N_9385,N_9429);
or U9545 (N_9545,N_9382,N_9328);
nand U9546 (N_9546,N_9439,N_9348);
xnor U9547 (N_9547,N_9398,N_9368);
and U9548 (N_9548,N_9392,N_9287);
nand U9549 (N_9549,N_9343,N_9381);
xnor U9550 (N_9550,N_9336,N_9430);
nand U9551 (N_9551,N_9417,N_9401);
nor U9552 (N_9552,N_9352,N_9370);
nand U9553 (N_9553,N_9328,N_9378);
xor U9554 (N_9554,N_9347,N_9371);
or U9555 (N_9555,N_9338,N_9415);
nor U9556 (N_9556,N_9352,N_9359);
or U9557 (N_9557,N_9330,N_9360);
xor U9558 (N_9558,N_9372,N_9347);
nor U9559 (N_9559,N_9409,N_9401);
or U9560 (N_9560,N_9310,N_9334);
nand U9561 (N_9561,N_9307,N_9392);
or U9562 (N_9562,N_9394,N_9340);
nand U9563 (N_9563,N_9325,N_9376);
xnor U9564 (N_9564,N_9390,N_9339);
nor U9565 (N_9565,N_9318,N_9283);
xor U9566 (N_9566,N_9423,N_9314);
nor U9567 (N_9567,N_9327,N_9298);
and U9568 (N_9568,N_9379,N_9395);
nor U9569 (N_9569,N_9431,N_9351);
and U9570 (N_9570,N_9402,N_9360);
or U9571 (N_9571,N_9344,N_9330);
nand U9572 (N_9572,N_9396,N_9433);
or U9573 (N_9573,N_9359,N_9283);
nor U9574 (N_9574,N_9317,N_9434);
or U9575 (N_9575,N_9387,N_9410);
and U9576 (N_9576,N_9402,N_9410);
xnor U9577 (N_9577,N_9383,N_9321);
and U9578 (N_9578,N_9295,N_9293);
and U9579 (N_9579,N_9438,N_9376);
xor U9580 (N_9580,N_9337,N_9421);
nand U9581 (N_9581,N_9381,N_9417);
or U9582 (N_9582,N_9317,N_9312);
or U9583 (N_9583,N_9425,N_9367);
nor U9584 (N_9584,N_9310,N_9420);
nand U9585 (N_9585,N_9323,N_9314);
xor U9586 (N_9586,N_9361,N_9300);
and U9587 (N_9587,N_9309,N_9378);
nor U9588 (N_9588,N_9307,N_9364);
or U9589 (N_9589,N_9418,N_9360);
or U9590 (N_9590,N_9433,N_9361);
or U9591 (N_9591,N_9339,N_9337);
and U9592 (N_9592,N_9389,N_9281);
nor U9593 (N_9593,N_9411,N_9307);
and U9594 (N_9594,N_9368,N_9439);
and U9595 (N_9595,N_9369,N_9337);
nor U9596 (N_9596,N_9339,N_9414);
xnor U9597 (N_9597,N_9335,N_9320);
and U9598 (N_9598,N_9345,N_9417);
or U9599 (N_9599,N_9299,N_9389);
and U9600 (N_9600,N_9485,N_9445);
nor U9601 (N_9601,N_9470,N_9441);
or U9602 (N_9602,N_9452,N_9527);
nand U9603 (N_9603,N_9538,N_9454);
xor U9604 (N_9604,N_9534,N_9461);
nand U9605 (N_9605,N_9559,N_9489);
and U9606 (N_9606,N_9487,N_9543);
xnor U9607 (N_9607,N_9569,N_9572);
or U9608 (N_9608,N_9440,N_9563);
nand U9609 (N_9609,N_9451,N_9583);
and U9610 (N_9610,N_9468,N_9592);
xnor U9611 (N_9611,N_9514,N_9593);
nand U9612 (N_9612,N_9504,N_9587);
nand U9613 (N_9613,N_9455,N_9530);
and U9614 (N_9614,N_9523,N_9469);
or U9615 (N_9615,N_9542,N_9540);
xor U9616 (N_9616,N_9558,N_9575);
nand U9617 (N_9617,N_9573,N_9532);
and U9618 (N_9618,N_9535,N_9537);
xnor U9619 (N_9619,N_9599,N_9566);
xor U9620 (N_9620,N_9588,N_9528);
nand U9621 (N_9621,N_9525,N_9449);
nand U9622 (N_9622,N_9529,N_9505);
nor U9623 (N_9623,N_9510,N_9536);
nor U9624 (N_9624,N_9479,N_9478);
and U9625 (N_9625,N_9442,N_9581);
nor U9626 (N_9626,N_9477,N_9458);
nand U9627 (N_9627,N_9544,N_9522);
or U9628 (N_9628,N_9517,N_9476);
and U9629 (N_9629,N_9494,N_9554);
xor U9630 (N_9630,N_9590,N_9561);
nand U9631 (N_9631,N_9594,N_9481);
nor U9632 (N_9632,N_9516,N_9511);
nand U9633 (N_9633,N_9465,N_9490);
nor U9634 (N_9634,N_9589,N_9556);
and U9635 (N_9635,N_9598,N_9456);
nor U9636 (N_9636,N_9576,N_9515);
nor U9637 (N_9637,N_9521,N_9518);
nand U9638 (N_9638,N_9578,N_9482);
nand U9639 (N_9639,N_9472,N_9552);
xor U9640 (N_9640,N_9462,N_9507);
nand U9641 (N_9641,N_9553,N_9565);
or U9642 (N_9642,N_9501,N_9500);
nand U9643 (N_9643,N_9577,N_9548);
and U9644 (N_9644,N_9595,N_9550);
and U9645 (N_9645,N_9513,N_9460);
nand U9646 (N_9646,N_9493,N_9498);
nor U9647 (N_9647,N_9509,N_9547);
and U9648 (N_9648,N_9564,N_9475);
xor U9649 (N_9649,N_9560,N_9503);
nand U9650 (N_9650,N_9463,N_9471);
or U9651 (N_9651,N_9488,N_9539);
or U9652 (N_9652,N_9571,N_9484);
nor U9653 (N_9653,N_9519,N_9467);
xnor U9654 (N_9654,N_9585,N_9562);
nand U9655 (N_9655,N_9551,N_9555);
nand U9656 (N_9656,N_9582,N_9492);
nand U9657 (N_9657,N_9597,N_9584);
nand U9658 (N_9658,N_9533,N_9443);
and U9659 (N_9659,N_9591,N_9586);
nor U9660 (N_9660,N_9464,N_9448);
nor U9661 (N_9661,N_9508,N_9457);
nor U9662 (N_9662,N_9526,N_9495);
xor U9663 (N_9663,N_9520,N_9459);
and U9664 (N_9664,N_9502,N_9473);
or U9665 (N_9665,N_9574,N_9506);
and U9666 (N_9666,N_9549,N_9483);
xor U9667 (N_9667,N_9444,N_9446);
xnor U9668 (N_9668,N_9447,N_9570);
nand U9669 (N_9669,N_9596,N_9499);
xnor U9670 (N_9670,N_9497,N_9453);
nor U9671 (N_9671,N_9466,N_9480);
xnor U9672 (N_9672,N_9557,N_9541);
and U9673 (N_9673,N_9580,N_9567);
nor U9674 (N_9674,N_9579,N_9568);
and U9675 (N_9675,N_9546,N_9512);
xor U9676 (N_9676,N_9486,N_9531);
and U9677 (N_9677,N_9491,N_9524);
xnor U9678 (N_9678,N_9496,N_9545);
nand U9679 (N_9679,N_9474,N_9450);
nand U9680 (N_9680,N_9527,N_9537);
or U9681 (N_9681,N_9589,N_9464);
nand U9682 (N_9682,N_9457,N_9470);
nor U9683 (N_9683,N_9592,N_9585);
or U9684 (N_9684,N_9524,N_9594);
or U9685 (N_9685,N_9565,N_9469);
xor U9686 (N_9686,N_9560,N_9543);
and U9687 (N_9687,N_9579,N_9511);
nor U9688 (N_9688,N_9452,N_9519);
xor U9689 (N_9689,N_9475,N_9559);
nand U9690 (N_9690,N_9544,N_9590);
nor U9691 (N_9691,N_9514,N_9518);
xnor U9692 (N_9692,N_9474,N_9477);
xor U9693 (N_9693,N_9511,N_9545);
and U9694 (N_9694,N_9541,N_9551);
or U9695 (N_9695,N_9449,N_9563);
xor U9696 (N_9696,N_9469,N_9510);
nand U9697 (N_9697,N_9452,N_9539);
xor U9698 (N_9698,N_9484,N_9550);
and U9699 (N_9699,N_9591,N_9560);
and U9700 (N_9700,N_9592,N_9574);
nor U9701 (N_9701,N_9547,N_9595);
xnor U9702 (N_9702,N_9538,N_9526);
xnor U9703 (N_9703,N_9462,N_9487);
nor U9704 (N_9704,N_9446,N_9490);
nand U9705 (N_9705,N_9539,N_9541);
nor U9706 (N_9706,N_9446,N_9547);
nor U9707 (N_9707,N_9587,N_9559);
or U9708 (N_9708,N_9475,N_9580);
nor U9709 (N_9709,N_9572,N_9584);
nor U9710 (N_9710,N_9585,N_9465);
or U9711 (N_9711,N_9473,N_9531);
nand U9712 (N_9712,N_9542,N_9485);
or U9713 (N_9713,N_9585,N_9512);
xor U9714 (N_9714,N_9516,N_9599);
and U9715 (N_9715,N_9500,N_9547);
xnor U9716 (N_9716,N_9574,N_9448);
and U9717 (N_9717,N_9461,N_9554);
xnor U9718 (N_9718,N_9567,N_9503);
and U9719 (N_9719,N_9511,N_9539);
nor U9720 (N_9720,N_9559,N_9524);
xor U9721 (N_9721,N_9554,N_9586);
xor U9722 (N_9722,N_9500,N_9462);
nand U9723 (N_9723,N_9446,N_9491);
and U9724 (N_9724,N_9499,N_9535);
xnor U9725 (N_9725,N_9468,N_9480);
xnor U9726 (N_9726,N_9441,N_9572);
nand U9727 (N_9727,N_9498,N_9442);
and U9728 (N_9728,N_9549,N_9537);
xor U9729 (N_9729,N_9567,N_9588);
nor U9730 (N_9730,N_9554,N_9581);
nor U9731 (N_9731,N_9558,N_9541);
nor U9732 (N_9732,N_9563,N_9541);
nand U9733 (N_9733,N_9512,N_9503);
nand U9734 (N_9734,N_9517,N_9579);
and U9735 (N_9735,N_9526,N_9536);
and U9736 (N_9736,N_9479,N_9496);
or U9737 (N_9737,N_9448,N_9465);
xor U9738 (N_9738,N_9565,N_9554);
nand U9739 (N_9739,N_9493,N_9463);
nand U9740 (N_9740,N_9478,N_9448);
nand U9741 (N_9741,N_9483,N_9531);
or U9742 (N_9742,N_9508,N_9531);
nor U9743 (N_9743,N_9576,N_9508);
nor U9744 (N_9744,N_9471,N_9593);
or U9745 (N_9745,N_9472,N_9570);
xnor U9746 (N_9746,N_9483,N_9471);
and U9747 (N_9747,N_9589,N_9471);
and U9748 (N_9748,N_9454,N_9473);
or U9749 (N_9749,N_9495,N_9570);
nor U9750 (N_9750,N_9550,N_9523);
and U9751 (N_9751,N_9465,N_9544);
xor U9752 (N_9752,N_9517,N_9486);
or U9753 (N_9753,N_9467,N_9573);
or U9754 (N_9754,N_9588,N_9480);
xnor U9755 (N_9755,N_9577,N_9564);
nor U9756 (N_9756,N_9588,N_9521);
or U9757 (N_9757,N_9543,N_9582);
and U9758 (N_9758,N_9560,N_9535);
nand U9759 (N_9759,N_9568,N_9490);
nand U9760 (N_9760,N_9667,N_9697);
nand U9761 (N_9761,N_9625,N_9619);
xnor U9762 (N_9762,N_9611,N_9746);
or U9763 (N_9763,N_9684,N_9606);
or U9764 (N_9764,N_9680,N_9695);
nor U9765 (N_9765,N_9636,N_9617);
nand U9766 (N_9766,N_9649,N_9759);
and U9767 (N_9767,N_9681,N_9605);
or U9768 (N_9768,N_9732,N_9730);
or U9769 (N_9769,N_9635,N_9712);
and U9770 (N_9770,N_9700,N_9683);
or U9771 (N_9771,N_9647,N_9656);
xnor U9772 (N_9772,N_9716,N_9705);
or U9773 (N_9773,N_9729,N_9754);
nand U9774 (N_9774,N_9715,N_9628);
nor U9775 (N_9775,N_9604,N_9740);
xor U9776 (N_9776,N_9634,N_9672);
nor U9777 (N_9777,N_9663,N_9731);
or U9778 (N_9778,N_9723,N_9629);
nand U9779 (N_9779,N_9748,N_9721);
xor U9780 (N_9780,N_9758,N_9670);
xnor U9781 (N_9781,N_9643,N_9718);
and U9782 (N_9782,N_9600,N_9620);
xor U9783 (N_9783,N_9638,N_9659);
nor U9784 (N_9784,N_9607,N_9690);
and U9785 (N_9785,N_9756,N_9713);
and U9786 (N_9786,N_9671,N_9645);
xnor U9787 (N_9787,N_9693,N_9698);
xnor U9788 (N_9788,N_9673,N_9678);
or U9789 (N_9789,N_9660,N_9624);
or U9790 (N_9790,N_9743,N_9736);
nor U9791 (N_9791,N_9669,N_9750);
nor U9792 (N_9792,N_9733,N_9666);
nor U9793 (N_9793,N_9696,N_9685);
nand U9794 (N_9794,N_9612,N_9626);
xnor U9795 (N_9795,N_9714,N_9602);
and U9796 (N_9796,N_9675,N_9637);
nor U9797 (N_9797,N_9615,N_9664);
or U9798 (N_9798,N_9662,N_9711);
or U9799 (N_9799,N_9622,N_9744);
nand U9800 (N_9800,N_9654,N_9701);
or U9801 (N_9801,N_9734,N_9603);
or U9802 (N_9802,N_9727,N_9640);
nor U9803 (N_9803,N_9631,N_9728);
or U9804 (N_9804,N_9601,N_9609);
xnor U9805 (N_9805,N_9742,N_9652);
or U9806 (N_9806,N_9689,N_9738);
nand U9807 (N_9807,N_9676,N_9632);
or U9808 (N_9808,N_9655,N_9614);
xor U9809 (N_9809,N_9692,N_9749);
xnor U9810 (N_9810,N_9665,N_9737);
and U9811 (N_9811,N_9610,N_9691);
nor U9812 (N_9812,N_9707,N_9613);
nand U9813 (N_9813,N_9630,N_9703);
or U9814 (N_9814,N_9752,N_9639);
xnor U9815 (N_9815,N_9687,N_9642);
or U9816 (N_9816,N_9674,N_9694);
nor U9817 (N_9817,N_9717,N_9621);
and U9818 (N_9818,N_9616,N_9755);
xnor U9819 (N_9819,N_9757,N_9725);
xor U9820 (N_9820,N_9646,N_9657);
xnor U9821 (N_9821,N_9709,N_9747);
and U9822 (N_9822,N_9739,N_9702);
xnor U9823 (N_9823,N_9741,N_9608);
nand U9824 (N_9824,N_9648,N_9688);
or U9825 (N_9825,N_9623,N_9745);
xor U9826 (N_9826,N_9720,N_9753);
xnor U9827 (N_9827,N_9627,N_9661);
xnor U9828 (N_9828,N_9686,N_9658);
nor U9829 (N_9829,N_9653,N_9735);
or U9830 (N_9830,N_9710,N_9679);
or U9831 (N_9831,N_9724,N_9651);
and U9832 (N_9832,N_9708,N_9682);
nand U9833 (N_9833,N_9751,N_9641);
nand U9834 (N_9834,N_9633,N_9668);
nor U9835 (N_9835,N_9719,N_9650);
nor U9836 (N_9836,N_9644,N_9722);
nor U9837 (N_9837,N_9699,N_9618);
and U9838 (N_9838,N_9706,N_9677);
and U9839 (N_9839,N_9704,N_9726);
nand U9840 (N_9840,N_9652,N_9616);
or U9841 (N_9841,N_9706,N_9727);
or U9842 (N_9842,N_9652,N_9682);
nor U9843 (N_9843,N_9644,N_9602);
nor U9844 (N_9844,N_9696,N_9747);
nor U9845 (N_9845,N_9739,N_9648);
nand U9846 (N_9846,N_9669,N_9602);
nor U9847 (N_9847,N_9747,N_9674);
or U9848 (N_9848,N_9731,N_9607);
and U9849 (N_9849,N_9693,N_9639);
nor U9850 (N_9850,N_9759,N_9706);
xor U9851 (N_9851,N_9608,N_9610);
nand U9852 (N_9852,N_9600,N_9666);
or U9853 (N_9853,N_9735,N_9708);
and U9854 (N_9854,N_9749,N_9719);
and U9855 (N_9855,N_9607,N_9696);
nor U9856 (N_9856,N_9605,N_9733);
nor U9857 (N_9857,N_9741,N_9747);
and U9858 (N_9858,N_9621,N_9625);
nand U9859 (N_9859,N_9704,N_9660);
and U9860 (N_9860,N_9722,N_9672);
xnor U9861 (N_9861,N_9691,N_9742);
and U9862 (N_9862,N_9612,N_9661);
and U9863 (N_9863,N_9705,N_9671);
xor U9864 (N_9864,N_9618,N_9604);
xnor U9865 (N_9865,N_9703,N_9628);
and U9866 (N_9866,N_9636,N_9727);
nor U9867 (N_9867,N_9714,N_9662);
or U9868 (N_9868,N_9722,N_9692);
xor U9869 (N_9869,N_9725,N_9715);
and U9870 (N_9870,N_9655,N_9749);
xor U9871 (N_9871,N_9687,N_9688);
or U9872 (N_9872,N_9744,N_9620);
and U9873 (N_9873,N_9698,N_9737);
and U9874 (N_9874,N_9757,N_9730);
nand U9875 (N_9875,N_9621,N_9744);
xnor U9876 (N_9876,N_9745,N_9606);
nand U9877 (N_9877,N_9748,N_9605);
and U9878 (N_9878,N_9705,N_9718);
nor U9879 (N_9879,N_9680,N_9638);
nor U9880 (N_9880,N_9677,N_9636);
and U9881 (N_9881,N_9730,N_9684);
nand U9882 (N_9882,N_9615,N_9626);
and U9883 (N_9883,N_9648,N_9719);
or U9884 (N_9884,N_9612,N_9663);
or U9885 (N_9885,N_9634,N_9750);
and U9886 (N_9886,N_9745,N_9753);
nor U9887 (N_9887,N_9698,N_9738);
nand U9888 (N_9888,N_9603,N_9738);
or U9889 (N_9889,N_9698,N_9642);
xnor U9890 (N_9890,N_9627,N_9729);
xnor U9891 (N_9891,N_9740,N_9734);
xor U9892 (N_9892,N_9627,N_9635);
xor U9893 (N_9893,N_9691,N_9640);
and U9894 (N_9894,N_9677,N_9685);
or U9895 (N_9895,N_9720,N_9684);
or U9896 (N_9896,N_9690,N_9605);
nand U9897 (N_9897,N_9750,N_9725);
and U9898 (N_9898,N_9633,N_9621);
nand U9899 (N_9899,N_9725,N_9680);
nor U9900 (N_9900,N_9623,N_9665);
nor U9901 (N_9901,N_9658,N_9738);
or U9902 (N_9902,N_9623,N_9637);
xnor U9903 (N_9903,N_9603,N_9684);
nor U9904 (N_9904,N_9603,N_9710);
nand U9905 (N_9905,N_9624,N_9736);
xor U9906 (N_9906,N_9642,N_9679);
or U9907 (N_9907,N_9717,N_9602);
xnor U9908 (N_9908,N_9705,N_9695);
nand U9909 (N_9909,N_9707,N_9651);
nand U9910 (N_9910,N_9717,N_9649);
xor U9911 (N_9911,N_9752,N_9670);
nor U9912 (N_9912,N_9659,N_9732);
xor U9913 (N_9913,N_9756,N_9629);
or U9914 (N_9914,N_9728,N_9617);
xnor U9915 (N_9915,N_9652,N_9732);
nand U9916 (N_9916,N_9740,N_9695);
nor U9917 (N_9917,N_9717,N_9667);
nor U9918 (N_9918,N_9717,N_9707);
nor U9919 (N_9919,N_9627,N_9744);
or U9920 (N_9920,N_9805,N_9761);
nor U9921 (N_9921,N_9766,N_9855);
or U9922 (N_9922,N_9814,N_9886);
and U9923 (N_9923,N_9793,N_9810);
nand U9924 (N_9924,N_9765,N_9880);
and U9925 (N_9925,N_9853,N_9887);
xnor U9926 (N_9926,N_9790,N_9822);
and U9927 (N_9927,N_9840,N_9797);
nor U9928 (N_9928,N_9884,N_9770);
xnor U9929 (N_9929,N_9857,N_9895);
nand U9930 (N_9930,N_9777,N_9901);
xor U9931 (N_9931,N_9815,N_9772);
nand U9932 (N_9932,N_9760,N_9803);
and U9933 (N_9933,N_9919,N_9866);
and U9934 (N_9934,N_9899,N_9861);
nor U9935 (N_9935,N_9826,N_9883);
nand U9936 (N_9936,N_9812,N_9903);
nor U9937 (N_9937,N_9786,N_9780);
nand U9938 (N_9938,N_9896,N_9862);
nor U9939 (N_9939,N_9858,N_9906);
xor U9940 (N_9940,N_9823,N_9769);
nor U9941 (N_9941,N_9912,N_9849);
nor U9942 (N_9942,N_9848,N_9825);
or U9943 (N_9943,N_9764,N_9854);
nand U9944 (N_9944,N_9802,N_9834);
and U9945 (N_9945,N_9804,N_9794);
xor U9946 (N_9946,N_9821,N_9787);
nand U9947 (N_9947,N_9763,N_9776);
and U9948 (N_9948,N_9845,N_9791);
nand U9949 (N_9949,N_9808,N_9865);
xor U9950 (N_9950,N_9875,N_9867);
nand U9951 (N_9951,N_9820,N_9859);
or U9952 (N_9952,N_9762,N_9842);
or U9953 (N_9953,N_9836,N_9773);
xnor U9954 (N_9954,N_9789,N_9900);
nor U9955 (N_9955,N_9908,N_9910);
nand U9956 (N_9956,N_9796,N_9778);
or U9957 (N_9957,N_9891,N_9851);
nor U9958 (N_9958,N_9915,N_9843);
nor U9959 (N_9959,N_9811,N_9824);
and U9960 (N_9960,N_9782,N_9835);
nor U9961 (N_9961,N_9874,N_9800);
nand U9962 (N_9962,N_9828,N_9841);
nor U9963 (N_9963,N_9829,N_9898);
xnor U9964 (N_9964,N_9864,N_9827);
or U9965 (N_9965,N_9831,N_9885);
or U9966 (N_9966,N_9871,N_9894);
xor U9967 (N_9967,N_9819,N_9846);
nand U9968 (N_9968,N_9767,N_9888);
nor U9969 (N_9969,N_9881,N_9784);
xnor U9970 (N_9970,N_9783,N_9918);
nor U9971 (N_9971,N_9774,N_9809);
nand U9972 (N_9972,N_9889,N_9914);
and U9973 (N_9973,N_9817,N_9795);
and U9974 (N_9974,N_9856,N_9905);
or U9975 (N_9975,N_9779,N_9832);
and U9976 (N_9976,N_9837,N_9813);
and U9977 (N_9977,N_9913,N_9882);
nor U9978 (N_9978,N_9768,N_9830);
xnor U9979 (N_9979,N_9792,N_9788);
or U9980 (N_9980,N_9801,N_9904);
and U9981 (N_9981,N_9775,N_9799);
xnor U9982 (N_9982,N_9847,N_9873);
nand U9983 (N_9983,N_9876,N_9868);
or U9984 (N_9984,N_9863,N_9771);
nor U9985 (N_9985,N_9911,N_9917);
nor U9986 (N_9986,N_9850,N_9785);
nor U9987 (N_9987,N_9872,N_9879);
or U9988 (N_9988,N_9877,N_9878);
xnor U9989 (N_9989,N_9844,N_9892);
and U9990 (N_9990,N_9806,N_9807);
or U9991 (N_9991,N_9869,N_9897);
nand U9992 (N_9992,N_9839,N_9890);
nor U9993 (N_9993,N_9838,N_9833);
and U9994 (N_9994,N_9860,N_9902);
or U9995 (N_9995,N_9916,N_9893);
xor U9996 (N_9996,N_9816,N_9909);
nor U9997 (N_9997,N_9852,N_9907);
nor U9998 (N_9998,N_9781,N_9798);
xnor U9999 (N_9999,N_9818,N_9870);
and U10000 (N_10000,N_9890,N_9799);
or U10001 (N_10001,N_9773,N_9889);
nand U10002 (N_10002,N_9768,N_9821);
nand U10003 (N_10003,N_9798,N_9810);
or U10004 (N_10004,N_9893,N_9826);
nor U10005 (N_10005,N_9822,N_9883);
and U10006 (N_10006,N_9816,N_9866);
xor U10007 (N_10007,N_9881,N_9847);
nor U10008 (N_10008,N_9789,N_9829);
or U10009 (N_10009,N_9914,N_9779);
or U10010 (N_10010,N_9911,N_9888);
nand U10011 (N_10011,N_9824,N_9771);
or U10012 (N_10012,N_9837,N_9851);
xnor U10013 (N_10013,N_9869,N_9782);
nor U10014 (N_10014,N_9857,N_9828);
nor U10015 (N_10015,N_9774,N_9801);
and U10016 (N_10016,N_9772,N_9862);
nand U10017 (N_10017,N_9821,N_9856);
nand U10018 (N_10018,N_9764,N_9887);
or U10019 (N_10019,N_9777,N_9842);
or U10020 (N_10020,N_9910,N_9794);
nor U10021 (N_10021,N_9800,N_9914);
xnor U10022 (N_10022,N_9794,N_9856);
or U10023 (N_10023,N_9837,N_9791);
or U10024 (N_10024,N_9837,N_9860);
nor U10025 (N_10025,N_9783,N_9832);
nor U10026 (N_10026,N_9784,N_9918);
nand U10027 (N_10027,N_9778,N_9765);
xor U10028 (N_10028,N_9783,N_9812);
or U10029 (N_10029,N_9837,N_9817);
or U10030 (N_10030,N_9840,N_9889);
nand U10031 (N_10031,N_9801,N_9856);
nand U10032 (N_10032,N_9794,N_9774);
xor U10033 (N_10033,N_9812,N_9789);
xor U10034 (N_10034,N_9840,N_9808);
or U10035 (N_10035,N_9830,N_9917);
nand U10036 (N_10036,N_9849,N_9774);
nor U10037 (N_10037,N_9850,N_9833);
and U10038 (N_10038,N_9912,N_9799);
nand U10039 (N_10039,N_9907,N_9881);
and U10040 (N_10040,N_9829,N_9779);
nand U10041 (N_10041,N_9845,N_9806);
and U10042 (N_10042,N_9919,N_9813);
or U10043 (N_10043,N_9837,N_9917);
nand U10044 (N_10044,N_9784,N_9814);
and U10045 (N_10045,N_9901,N_9851);
xor U10046 (N_10046,N_9896,N_9766);
and U10047 (N_10047,N_9810,N_9781);
nand U10048 (N_10048,N_9877,N_9835);
or U10049 (N_10049,N_9805,N_9830);
nor U10050 (N_10050,N_9783,N_9818);
xnor U10051 (N_10051,N_9905,N_9818);
or U10052 (N_10052,N_9913,N_9863);
or U10053 (N_10053,N_9777,N_9812);
nor U10054 (N_10054,N_9813,N_9887);
and U10055 (N_10055,N_9825,N_9806);
xor U10056 (N_10056,N_9847,N_9843);
or U10057 (N_10057,N_9890,N_9773);
and U10058 (N_10058,N_9844,N_9916);
nand U10059 (N_10059,N_9769,N_9914);
nor U10060 (N_10060,N_9883,N_9908);
or U10061 (N_10061,N_9873,N_9812);
nor U10062 (N_10062,N_9777,N_9850);
nor U10063 (N_10063,N_9834,N_9839);
and U10064 (N_10064,N_9786,N_9853);
nand U10065 (N_10065,N_9818,N_9898);
or U10066 (N_10066,N_9826,N_9815);
and U10067 (N_10067,N_9863,N_9779);
or U10068 (N_10068,N_9881,N_9793);
nor U10069 (N_10069,N_9764,N_9895);
or U10070 (N_10070,N_9793,N_9876);
and U10071 (N_10071,N_9855,N_9795);
nor U10072 (N_10072,N_9806,N_9843);
or U10073 (N_10073,N_9831,N_9824);
and U10074 (N_10074,N_9854,N_9882);
and U10075 (N_10075,N_9875,N_9809);
nor U10076 (N_10076,N_9786,N_9826);
and U10077 (N_10077,N_9862,N_9864);
nor U10078 (N_10078,N_9902,N_9774);
or U10079 (N_10079,N_9861,N_9788);
and U10080 (N_10080,N_10019,N_10078);
nand U10081 (N_10081,N_9962,N_9934);
xnor U10082 (N_10082,N_9946,N_9940);
or U10083 (N_10083,N_9926,N_9964);
nor U10084 (N_10084,N_9945,N_9941);
xor U10085 (N_10085,N_10014,N_10060);
nor U10086 (N_10086,N_10021,N_10006);
nand U10087 (N_10087,N_10056,N_9986);
and U10088 (N_10088,N_10018,N_9990);
nand U10089 (N_10089,N_9938,N_10031);
xor U10090 (N_10090,N_9923,N_10012);
and U10091 (N_10091,N_10049,N_10023);
and U10092 (N_10092,N_9953,N_9965);
nor U10093 (N_10093,N_10068,N_9979);
nand U10094 (N_10094,N_9925,N_9996);
or U10095 (N_10095,N_10042,N_10002);
and U10096 (N_10096,N_10036,N_10069);
or U10097 (N_10097,N_9935,N_9967);
nand U10098 (N_10098,N_10079,N_9955);
xnor U10099 (N_10099,N_9943,N_9949);
xor U10100 (N_10100,N_9961,N_10070);
nor U10101 (N_10101,N_9936,N_10030);
nor U10102 (N_10102,N_9997,N_9969);
nand U10103 (N_10103,N_10028,N_9952);
and U10104 (N_10104,N_10003,N_9947);
and U10105 (N_10105,N_9981,N_10041);
nand U10106 (N_10106,N_10046,N_10071);
nand U10107 (N_10107,N_10048,N_9924);
nand U10108 (N_10108,N_10017,N_9994);
and U10109 (N_10109,N_9931,N_10052);
and U10110 (N_10110,N_9929,N_10067);
nand U10111 (N_10111,N_9937,N_9999);
nand U10112 (N_10112,N_9972,N_10050);
and U10113 (N_10113,N_9974,N_10038);
nand U10114 (N_10114,N_10008,N_9958);
or U10115 (N_10115,N_10065,N_10055);
xnor U10116 (N_10116,N_9993,N_10001);
xnor U10117 (N_10117,N_10000,N_10061);
nand U10118 (N_10118,N_9978,N_9968);
or U10119 (N_10119,N_9980,N_10010);
nand U10120 (N_10120,N_10045,N_10073);
xnor U10121 (N_10121,N_10044,N_10057);
nor U10122 (N_10122,N_9950,N_9984);
and U10123 (N_10123,N_9944,N_9977);
nand U10124 (N_10124,N_10039,N_9971);
xor U10125 (N_10125,N_10035,N_10051);
nor U10126 (N_10126,N_9989,N_10004);
and U10127 (N_10127,N_9942,N_10007);
nor U10128 (N_10128,N_10032,N_9956);
nor U10129 (N_10129,N_9975,N_10062);
nand U10130 (N_10130,N_9933,N_10037);
and U10131 (N_10131,N_9983,N_9991);
nand U10132 (N_10132,N_9966,N_9976);
xor U10133 (N_10133,N_10016,N_10059);
or U10134 (N_10134,N_9954,N_9982);
and U10135 (N_10135,N_9951,N_9987);
nor U10136 (N_10136,N_10009,N_10020);
xnor U10137 (N_10137,N_9932,N_10054);
nor U10138 (N_10138,N_9960,N_10063);
or U10139 (N_10139,N_9992,N_10011);
nor U10140 (N_10140,N_10076,N_10053);
or U10141 (N_10141,N_10077,N_9963);
and U10142 (N_10142,N_9922,N_9928);
xor U10143 (N_10143,N_10027,N_9921);
or U10144 (N_10144,N_9920,N_9995);
xnor U10145 (N_10145,N_10033,N_9939);
nor U10146 (N_10146,N_10025,N_10026);
and U10147 (N_10147,N_10034,N_10064);
or U10148 (N_10148,N_10040,N_9985);
or U10149 (N_10149,N_9927,N_10043);
nand U10150 (N_10150,N_10022,N_9970);
xnor U10151 (N_10151,N_10029,N_10066);
or U10152 (N_10152,N_9930,N_10005);
xnor U10153 (N_10153,N_10047,N_10075);
xnor U10154 (N_10154,N_10024,N_9988);
or U10155 (N_10155,N_10058,N_10074);
nor U10156 (N_10156,N_10013,N_9948);
nand U10157 (N_10157,N_9957,N_9973);
nor U10158 (N_10158,N_10015,N_9998);
nand U10159 (N_10159,N_9959,N_10072);
nor U10160 (N_10160,N_9966,N_10039);
nor U10161 (N_10161,N_10035,N_9941);
or U10162 (N_10162,N_10062,N_9966);
xor U10163 (N_10163,N_10077,N_10063);
xor U10164 (N_10164,N_10052,N_9958);
and U10165 (N_10165,N_9991,N_9925);
and U10166 (N_10166,N_10027,N_9923);
or U10167 (N_10167,N_10061,N_9942);
nand U10168 (N_10168,N_9999,N_10043);
xor U10169 (N_10169,N_9999,N_9988);
nand U10170 (N_10170,N_9939,N_9969);
or U10171 (N_10171,N_9938,N_10004);
xnor U10172 (N_10172,N_9928,N_9967);
or U10173 (N_10173,N_9995,N_9925);
and U10174 (N_10174,N_10018,N_10059);
nor U10175 (N_10175,N_10010,N_10061);
or U10176 (N_10176,N_9964,N_9989);
xor U10177 (N_10177,N_10061,N_10021);
nand U10178 (N_10178,N_9971,N_10070);
nor U10179 (N_10179,N_9932,N_10079);
and U10180 (N_10180,N_9972,N_10079);
nand U10181 (N_10181,N_10001,N_10004);
xnor U10182 (N_10182,N_10011,N_10070);
xor U10183 (N_10183,N_10029,N_9999);
and U10184 (N_10184,N_10014,N_10017);
nor U10185 (N_10185,N_10008,N_9950);
xor U10186 (N_10186,N_10023,N_10033);
or U10187 (N_10187,N_9951,N_10068);
and U10188 (N_10188,N_10042,N_10022);
nand U10189 (N_10189,N_10037,N_9943);
or U10190 (N_10190,N_9981,N_9923);
and U10191 (N_10191,N_9985,N_9972);
xnor U10192 (N_10192,N_10036,N_10029);
or U10193 (N_10193,N_9973,N_9932);
xor U10194 (N_10194,N_9977,N_9935);
xor U10195 (N_10195,N_9973,N_9940);
and U10196 (N_10196,N_10016,N_10053);
or U10197 (N_10197,N_10022,N_9952);
and U10198 (N_10198,N_10000,N_9986);
and U10199 (N_10199,N_10040,N_9969);
and U10200 (N_10200,N_10026,N_10040);
nand U10201 (N_10201,N_10004,N_10032);
and U10202 (N_10202,N_10005,N_9938);
and U10203 (N_10203,N_9995,N_9981);
nor U10204 (N_10204,N_10026,N_9970);
nor U10205 (N_10205,N_10053,N_10027);
or U10206 (N_10206,N_10010,N_10076);
xor U10207 (N_10207,N_10079,N_9983);
or U10208 (N_10208,N_10025,N_9924);
nor U10209 (N_10209,N_10054,N_10064);
xor U10210 (N_10210,N_9933,N_10012);
nand U10211 (N_10211,N_9990,N_10071);
or U10212 (N_10212,N_9964,N_9968);
nor U10213 (N_10213,N_10070,N_9969);
nor U10214 (N_10214,N_10020,N_10043);
nor U10215 (N_10215,N_9941,N_10010);
or U10216 (N_10216,N_9952,N_10066);
and U10217 (N_10217,N_9993,N_9947);
and U10218 (N_10218,N_9971,N_10033);
nand U10219 (N_10219,N_10033,N_10068);
nor U10220 (N_10220,N_9981,N_9994);
nand U10221 (N_10221,N_10077,N_10046);
or U10222 (N_10222,N_9950,N_10043);
nor U10223 (N_10223,N_10016,N_10079);
nand U10224 (N_10224,N_10040,N_9928);
xnor U10225 (N_10225,N_9990,N_9939);
or U10226 (N_10226,N_10048,N_10022);
nor U10227 (N_10227,N_9963,N_10078);
or U10228 (N_10228,N_9940,N_9943);
xnor U10229 (N_10229,N_10060,N_9933);
nand U10230 (N_10230,N_9938,N_10048);
xnor U10231 (N_10231,N_9936,N_9935);
and U10232 (N_10232,N_10030,N_9979);
and U10233 (N_10233,N_10055,N_10057);
or U10234 (N_10234,N_10028,N_9976);
and U10235 (N_10235,N_10019,N_10028);
nor U10236 (N_10236,N_10058,N_9933);
and U10237 (N_10237,N_10025,N_10023);
nand U10238 (N_10238,N_10079,N_9964);
xor U10239 (N_10239,N_10077,N_9937);
nand U10240 (N_10240,N_10217,N_10183);
xnor U10241 (N_10241,N_10237,N_10198);
nand U10242 (N_10242,N_10109,N_10223);
or U10243 (N_10243,N_10186,N_10197);
and U10244 (N_10244,N_10165,N_10104);
xnor U10245 (N_10245,N_10224,N_10094);
nor U10246 (N_10246,N_10154,N_10081);
or U10247 (N_10247,N_10150,N_10175);
and U10248 (N_10248,N_10185,N_10236);
xor U10249 (N_10249,N_10204,N_10188);
nor U10250 (N_10250,N_10173,N_10116);
xor U10251 (N_10251,N_10147,N_10202);
and U10252 (N_10252,N_10130,N_10097);
nor U10253 (N_10253,N_10152,N_10235);
and U10254 (N_10254,N_10201,N_10122);
and U10255 (N_10255,N_10196,N_10099);
nand U10256 (N_10256,N_10164,N_10146);
and U10257 (N_10257,N_10213,N_10091);
and U10258 (N_10258,N_10163,N_10149);
nor U10259 (N_10259,N_10086,N_10229);
nor U10260 (N_10260,N_10108,N_10231);
and U10261 (N_10261,N_10189,N_10101);
nand U10262 (N_10262,N_10082,N_10093);
nand U10263 (N_10263,N_10187,N_10098);
nand U10264 (N_10264,N_10092,N_10143);
xor U10265 (N_10265,N_10100,N_10083);
nand U10266 (N_10266,N_10084,N_10238);
nand U10267 (N_10267,N_10141,N_10102);
and U10268 (N_10268,N_10191,N_10095);
or U10269 (N_10269,N_10111,N_10087);
nor U10270 (N_10270,N_10182,N_10123);
or U10271 (N_10271,N_10127,N_10157);
or U10272 (N_10272,N_10113,N_10106);
nand U10273 (N_10273,N_10153,N_10207);
xnor U10274 (N_10274,N_10214,N_10105);
xor U10275 (N_10275,N_10115,N_10221);
and U10276 (N_10276,N_10103,N_10218);
nand U10277 (N_10277,N_10232,N_10118);
or U10278 (N_10278,N_10225,N_10222);
nand U10279 (N_10279,N_10233,N_10228);
xnor U10280 (N_10280,N_10166,N_10205);
xnor U10281 (N_10281,N_10126,N_10220);
xor U10282 (N_10282,N_10124,N_10226);
and U10283 (N_10283,N_10090,N_10190);
or U10284 (N_10284,N_10216,N_10178);
nand U10285 (N_10285,N_10134,N_10156);
nand U10286 (N_10286,N_10227,N_10159);
nor U10287 (N_10287,N_10206,N_10212);
nor U10288 (N_10288,N_10107,N_10133);
nor U10289 (N_10289,N_10096,N_10209);
nor U10290 (N_10290,N_10171,N_10121);
nor U10291 (N_10291,N_10158,N_10120);
and U10292 (N_10292,N_10219,N_10174);
and U10293 (N_10293,N_10089,N_10162);
nand U10294 (N_10294,N_10144,N_10131);
nand U10295 (N_10295,N_10210,N_10138);
and U10296 (N_10296,N_10195,N_10192);
nor U10297 (N_10297,N_10234,N_10177);
and U10298 (N_10298,N_10117,N_10211);
and U10299 (N_10299,N_10208,N_10170);
nand U10300 (N_10300,N_10112,N_10136);
xnor U10301 (N_10301,N_10145,N_10139);
nor U10302 (N_10302,N_10129,N_10161);
nor U10303 (N_10303,N_10230,N_10125);
xnor U10304 (N_10304,N_10169,N_10203);
nor U10305 (N_10305,N_10199,N_10179);
nand U10306 (N_10306,N_10176,N_10085);
nand U10307 (N_10307,N_10200,N_10180);
or U10308 (N_10308,N_10215,N_10142);
xnor U10309 (N_10309,N_10132,N_10137);
and U10310 (N_10310,N_10119,N_10194);
nand U10311 (N_10311,N_10110,N_10239);
and U10312 (N_10312,N_10114,N_10172);
and U10313 (N_10313,N_10088,N_10148);
xnor U10314 (N_10314,N_10155,N_10184);
or U10315 (N_10315,N_10135,N_10140);
nand U10316 (N_10316,N_10167,N_10193);
and U10317 (N_10317,N_10080,N_10160);
nor U10318 (N_10318,N_10151,N_10128);
xnor U10319 (N_10319,N_10168,N_10181);
xnor U10320 (N_10320,N_10209,N_10145);
or U10321 (N_10321,N_10111,N_10146);
nor U10322 (N_10322,N_10227,N_10107);
nor U10323 (N_10323,N_10235,N_10167);
and U10324 (N_10324,N_10154,N_10093);
nor U10325 (N_10325,N_10128,N_10140);
or U10326 (N_10326,N_10154,N_10085);
nand U10327 (N_10327,N_10187,N_10213);
nor U10328 (N_10328,N_10178,N_10180);
and U10329 (N_10329,N_10116,N_10148);
and U10330 (N_10330,N_10236,N_10087);
xor U10331 (N_10331,N_10119,N_10177);
and U10332 (N_10332,N_10234,N_10118);
xnor U10333 (N_10333,N_10196,N_10095);
and U10334 (N_10334,N_10180,N_10098);
or U10335 (N_10335,N_10124,N_10147);
and U10336 (N_10336,N_10132,N_10139);
xnor U10337 (N_10337,N_10148,N_10122);
nand U10338 (N_10338,N_10196,N_10185);
nor U10339 (N_10339,N_10110,N_10095);
xnor U10340 (N_10340,N_10184,N_10156);
nor U10341 (N_10341,N_10145,N_10158);
nand U10342 (N_10342,N_10217,N_10120);
xnor U10343 (N_10343,N_10206,N_10186);
nand U10344 (N_10344,N_10129,N_10136);
nor U10345 (N_10345,N_10208,N_10147);
nand U10346 (N_10346,N_10225,N_10107);
nand U10347 (N_10347,N_10185,N_10105);
xor U10348 (N_10348,N_10121,N_10153);
xor U10349 (N_10349,N_10225,N_10197);
and U10350 (N_10350,N_10195,N_10164);
nand U10351 (N_10351,N_10099,N_10192);
and U10352 (N_10352,N_10086,N_10237);
or U10353 (N_10353,N_10236,N_10101);
nor U10354 (N_10354,N_10083,N_10181);
nand U10355 (N_10355,N_10226,N_10111);
xnor U10356 (N_10356,N_10198,N_10193);
or U10357 (N_10357,N_10197,N_10144);
xor U10358 (N_10358,N_10223,N_10111);
xnor U10359 (N_10359,N_10161,N_10150);
xnor U10360 (N_10360,N_10086,N_10222);
nor U10361 (N_10361,N_10120,N_10216);
and U10362 (N_10362,N_10085,N_10125);
xnor U10363 (N_10363,N_10080,N_10226);
nor U10364 (N_10364,N_10137,N_10231);
xor U10365 (N_10365,N_10182,N_10132);
and U10366 (N_10366,N_10106,N_10217);
or U10367 (N_10367,N_10168,N_10189);
nor U10368 (N_10368,N_10100,N_10186);
xnor U10369 (N_10369,N_10146,N_10096);
nand U10370 (N_10370,N_10214,N_10114);
nand U10371 (N_10371,N_10182,N_10229);
and U10372 (N_10372,N_10208,N_10193);
or U10373 (N_10373,N_10172,N_10196);
nand U10374 (N_10374,N_10194,N_10108);
nand U10375 (N_10375,N_10098,N_10194);
nor U10376 (N_10376,N_10137,N_10091);
nand U10377 (N_10377,N_10108,N_10196);
xnor U10378 (N_10378,N_10193,N_10137);
nor U10379 (N_10379,N_10171,N_10100);
and U10380 (N_10380,N_10163,N_10176);
nand U10381 (N_10381,N_10148,N_10143);
nand U10382 (N_10382,N_10228,N_10181);
nand U10383 (N_10383,N_10165,N_10166);
xnor U10384 (N_10384,N_10226,N_10200);
or U10385 (N_10385,N_10166,N_10086);
nand U10386 (N_10386,N_10186,N_10192);
nand U10387 (N_10387,N_10144,N_10125);
xor U10388 (N_10388,N_10170,N_10190);
nand U10389 (N_10389,N_10137,N_10144);
or U10390 (N_10390,N_10138,N_10149);
nand U10391 (N_10391,N_10192,N_10238);
nor U10392 (N_10392,N_10171,N_10192);
xnor U10393 (N_10393,N_10200,N_10165);
xnor U10394 (N_10394,N_10149,N_10129);
nor U10395 (N_10395,N_10083,N_10189);
or U10396 (N_10396,N_10136,N_10108);
nand U10397 (N_10397,N_10108,N_10193);
nor U10398 (N_10398,N_10167,N_10185);
nor U10399 (N_10399,N_10188,N_10096);
and U10400 (N_10400,N_10341,N_10304);
and U10401 (N_10401,N_10241,N_10336);
xor U10402 (N_10402,N_10376,N_10396);
and U10403 (N_10403,N_10386,N_10328);
or U10404 (N_10404,N_10276,N_10302);
or U10405 (N_10405,N_10279,N_10398);
or U10406 (N_10406,N_10368,N_10322);
nor U10407 (N_10407,N_10282,N_10323);
and U10408 (N_10408,N_10289,N_10327);
nor U10409 (N_10409,N_10337,N_10308);
or U10410 (N_10410,N_10300,N_10278);
xnor U10411 (N_10411,N_10256,N_10360);
and U10412 (N_10412,N_10292,N_10370);
nand U10413 (N_10413,N_10391,N_10262);
nor U10414 (N_10414,N_10394,N_10258);
nor U10415 (N_10415,N_10268,N_10266);
nor U10416 (N_10416,N_10363,N_10293);
or U10417 (N_10417,N_10338,N_10381);
or U10418 (N_10418,N_10367,N_10250);
nor U10419 (N_10419,N_10343,N_10379);
nand U10420 (N_10420,N_10371,N_10257);
xor U10421 (N_10421,N_10362,N_10320);
and U10422 (N_10422,N_10314,N_10380);
nand U10423 (N_10423,N_10387,N_10309);
xnor U10424 (N_10424,N_10244,N_10388);
and U10425 (N_10425,N_10374,N_10330);
and U10426 (N_10426,N_10285,N_10348);
nor U10427 (N_10427,N_10283,N_10267);
or U10428 (N_10428,N_10366,N_10357);
nor U10429 (N_10429,N_10354,N_10253);
and U10430 (N_10430,N_10325,N_10392);
nand U10431 (N_10431,N_10318,N_10312);
xnor U10432 (N_10432,N_10275,N_10333);
nor U10433 (N_10433,N_10332,N_10247);
and U10434 (N_10434,N_10378,N_10271);
and U10435 (N_10435,N_10383,N_10375);
and U10436 (N_10436,N_10390,N_10321);
xor U10437 (N_10437,N_10353,N_10242);
and U10438 (N_10438,N_10310,N_10399);
nor U10439 (N_10439,N_10260,N_10284);
and U10440 (N_10440,N_10270,N_10305);
nand U10441 (N_10441,N_10265,N_10299);
nor U10442 (N_10442,N_10372,N_10254);
or U10443 (N_10443,N_10356,N_10349);
nand U10444 (N_10444,N_10251,N_10280);
nand U10445 (N_10445,N_10334,N_10384);
or U10446 (N_10446,N_10355,N_10246);
or U10447 (N_10447,N_10307,N_10306);
and U10448 (N_10448,N_10373,N_10339);
nand U10449 (N_10449,N_10311,N_10365);
or U10450 (N_10450,N_10364,N_10358);
or U10451 (N_10451,N_10288,N_10303);
or U10452 (N_10452,N_10351,N_10345);
xor U10453 (N_10453,N_10261,N_10240);
and U10454 (N_10454,N_10393,N_10259);
or U10455 (N_10455,N_10255,N_10248);
nand U10456 (N_10456,N_10340,N_10290);
or U10457 (N_10457,N_10273,N_10286);
nand U10458 (N_10458,N_10316,N_10269);
nand U10459 (N_10459,N_10317,N_10264);
nor U10460 (N_10460,N_10287,N_10324);
or U10461 (N_10461,N_10291,N_10397);
xor U10462 (N_10462,N_10346,N_10295);
nor U10463 (N_10463,N_10331,N_10263);
or U10464 (N_10464,N_10252,N_10389);
and U10465 (N_10465,N_10352,N_10298);
nand U10466 (N_10466,N_10395,N_10344);
or U10467 (N_10467,N_10296,N_10313);
and U10468 (N_10468,N_10369,N_10245);
xor U10469 (N_10469,N_10326,N_10359);
nor U10470 (N_10470,N_10319,N_10297);
nor U10471 (N_10471,N_10361,N_10382);
and U10472 (N_10472,N_10385,N_10342);
and U10473 (N_10473,N_10272,N_10377);
and U10474 (N_10474,N_10249,N_10335);
xnor U10475 (N_10475,N_10281,N_10243);
nor U10476 (N_10476,N_10347,N_10329);
nor U10477 (N_10477,N_10277,N_10350);
nor U10478 (N_10478,N_10301,N_10294);
or U10479 (N_10479,N_10315,N_10274);
or U10480 (N_10480,N_10279,N_10318);
and U10481 (N_10481,N_10282,N_10387);
nand U10482 (N_10482,N_10392,N_10341);
xnor U10483 (N_10483,N_10347,N_10296);
nand U10484 (N_10484,N_10313,N_10270);
nor U10485 (N_10485,N_10365,N_10242);
xnor U10486 (N_10486,N_10296,N_10251);
xor U10487 (N_10487,N_10382,N_10354);
or U10488 (N_10488,N_10271,N_10290);
xor U10489 (N_10489,N_10362,N_10369);
nand U10490 (N_10490,N_10256,N_10393);
and U10491 (N_10491,N_10293,N_10376);
nand U10492 (N_10492,N_10323,N_10371);
and U10493 (N_10493,N_10277,N_10344);
nand U10494 (N_10494,N_10244,N_10278);
nand U10495 (N_10495,N_10306,N_10392);
and U10496 (N_10496,N_10373,N_10309);
nand U10497 (N_10497,N_10393,N_10332);
or U10498 (N_10498,N_10352,N_10328);
and U10499 (N_10499,N_10242,N_10378);
nand U10500 (N_10500,N_10243,N_10300);
and U10501 (N_10501,N_10331,N_10394);
and U10502 (N_10502,N_10312,N_10285);
xnor U10503 (N_10503,N_10252,N_10278);
and U10504 (N_10504,N_10298,N_10322);
and U10505 (N_10505,N_10343,N_10354);
or U10506 (N_10506,N_10311,N_10325);
and U10507 (N_10507,N_10267,N_10348);
and U10508 (N_10508,N_10254,N_10330);
nand U10509 (N_10509,N_10320,N_10345);
nand U10510 (N_10510,N_10395,N_10304);
and U10511 (N_10511,N_10264,N_10369);
nor U10512 (N_10512,N_10296,N_10392);
nand U10513 (N_10513,N_10379,N_10293);
nand U10514 (N_10514,N_10264,N_10391);
nor U10515 (N_10515,N_10338,N_10358);
nand U10516 (N_10516,N_10278,N_10284);
and U10517 (N_10517,N_10281,N_10263);
nand U10518 (N_10518,N_10304,N_10249);
nand U10519 (N_10519,N_10372,N_10312);
and U10520 (N_10520,N_10317,N_10296);
xor U10521 (N_10521,N_10257,N_10333);
and U10522 (N_10522,N_10305,N_10300);
nand U10523 (N_10523,N_10397,N_10353);
xor U10524 (N_10524,N_10249,N_10284);
nor U10525 (N_10525,N_10310,N_10363);
and U10526 (N_10526,N_10284,N_10298);
xnor U10527 (N_10527,N_10274,N_10369);
xor U10528 (N_10528,N_10260,N_10281);
nand U10529 (N_10529,N_10387,N_10254);
xnor U10530 (N_10530,N_10323,N_10255);
nand U10531 (N_10531,N_10365,N_10378);
nand U10532 (N_10532,N_10343,N_10326);
nand U10533 (N_10533,N_10344,N_10260);
or U10534 (N_10534,N_10249,N_10287);
or U10535 (N_10535,N_10250,N_10376);
xnor U10536 (N_10536,N_10391,N_10382);
xor U10537 (N_10537,N_10248,N_10292);
nand U10538 (N_10538,N_10333,N_10342);
or U10539 (N_10539,N_10316,N_10303);
or U10540 (N_10540,N_10300,N_10320);
xnor U10541 (N_10541,N_10260,N_10272);
nand U10542 (N_10542,N_10324,N_10348);
nor U10543 (N_10543,N_10256,N_10269);
and U10544 (N_10544,N_10335,N_10318);
and U10545 (N_10545,N_10334,N_10332);
or U10546 (N_10546,N_10269,N_10347);
or U10547 (N_10547,N_10307,N_10277);
nor U10548 (N_10548,N_10275,N_10392);
nand U10549 (N_10549,N_10341,N_10308);
nor U10550 (N_10550,N_10275,N_10321);
nor U10551 (N_10551,N_10340,N_10366);
or U10552 (N_10552,N_10299,N_10286);
xor U10553 (N_10553,N_10351,N_10368);
xor U10554 (N_10554,N_10350,N_10397);
nand U10555 (N_10555,N_10366,N_10256);
or U10556 (N_10556,N_10317,N_10310);
or U10557 (N_10557,N_10395,N_10283);
xnor U10558 (N_10558,N_10327,N_10286);
nor U10559 (N_10559,N_10263,N_10351);
nor U10560 (N_10560,N_10441,N_10500);
nand U10561 (N_10561,N_10532,N_10417);
nor U10562 (N_10562,N_10524,N_10480);
nand U10563 (N_10563,N_10422,N_10424);
and U10564 (N_10564,N_10485,N_10423);
or U10565 (N_10565,N_10452,N_10559);
nand U10566 (N_10566,N_10547,N_10482);
or U10567 (N_10567,N_10510,N_10474);
nand U10568 (N_10568,N_10428,N_10479);
and U10569 (N_10569,N_10418,N_10539);
nor U10570 (N_10570,N_10543,N_10463);
and U10571 (N_10571,N_10407,N_10549);
or U10572 (N_10572,N_10436,N_10409);
nand U10573 (N_10573,N_10408,N_10427);
nor U10574 (N_10574,N_10536,N_10451);
and U10575 (N_10575,N_10552,N_10495);
nor U10576 (N_10576,N_10459,N_10433);
nor U10577 (N_10577,N_10553,N_10509);
and U10578 (N_10578,N_10429,N_10513);
nand U10579 (N_10579,N_10499,N_10456);
xor U10580 (N_10580,N_10481,N_10530);
nand U10581 (N_10581,N_10516,N_10534);
nand U10582 (N_10582,N_10440,N_10420);
or U10583 (N_10583,N_10557,N_10448);
and U10584 (N_10584,N_10522,N_10467);
xnor U10585 (N_10585,N_10434,N_10492);
nand U10586 (N_10586,N_10455,N_10556);
nor U10587 (N_10587,N_10437,N_10506);
or U10588 (N_10588,N_10526,N_10486);
nor U10589 (N_10589,N_10465,N_10478);
xnor U10590 (N_10590,N_10405,N_10512);
nor U10591 (N_10591,N_10507,N_10454);
and U10592 (N_10592,N_10403,N_10489);
xnor U10593 (N_10593,N_10501,N_10477);
nor U10594 (N_10594,N_10401,N_10523);
nor U10595 (N_10595,N_10439,N_10446);
nor U10596 (N_10596,N_10431,N_10551);
and U10597 (N_10597,N_10515,N_10538);
xor U10598 (N_10598,N_10484,N_10504);
nor U10599 (N_10599,N_10466,N_10410);
or U10600 (N_10600,N_10430,N_10545);
and U10601 (N_10601,N_10502,N_10473);
nand U10602 (N_10602,N_10494,N_10476);
nor U10603 (N_10603,N_10444,N_10442);
or U10604 (N_10604,N_10520,N_10491);
nor U10605 (N_10605,N_10531,N_10497);
and U10606 (N_10606,N_10464,N_10508);
xor U10607 (N_10607,N_10450,N_10488);
nor U10608 (N_10608,N_10402,N_10438);
and U10609 (N_10609,N_10498,N_10535);
nor U10610 (N_10610,N_10413,N_10449);
and U10611 (N_10611,N_10550,N_10518);
nor U10612 (N_10612,N_10404,N_10548);
xor U10613 (N_10613,N_10469,N_10490);
nand U10614 (N_10614,N_10443,N_10453);
or U10615 (N_10615,N_10493,N_10457);
nor U10616 (N_10616,N_10517,N_10525);
or U10617 (N_10617,N_10527,N_10546);
or U10618 (N_10618,N_10445,N_10511);
nor U10619 (N_10619,N_10519,N_10528);
nand U10620 (N_10620,N_10458,N_10521);
nand U10621 (N_10621,N_10461,N_10421);
or U10622 (N_10622,N_10487,N_10406);
xnor U10623 (N_10623,N_10470,N_10415);
xnor U10624 (N_10624,N_10472,N_10537);
xnor U10625 (N_10625,N_10471,N_10540);
nor U10626 (N_10626,N_10514,N_10462);
and U10627 (N_10627,N_10426,N_10400);
xor U10628 (N_10628,N_10533,N_10542);
and U10629 (N_10629,N_10483,N_10544);
or U10630 (N_10630,N_10419,N_10460);
xnor U10631 (N_10631,N_10529,N_10503);
or U10632 (N_10632,N_10411,N_10554);
and U10633 (N_10633,N_10475,N_10412);
or U10634 (N_10634,N_10496,N_10414);
or U10635 (N_10635,N_10468,N_10505);
nor U10636 (N_10636,N_10425,N_10416);
and U10637 (N_10637,N_10435,N_10555);
or U10638 (N_10638,N_10432,N_10541);
or U10639 (N_10639,N_10447,N_10558);
and U10640 (N_10640,N_10529,N_10526);
nand U10641 (N_10641,N_10551,N_10404);
or U10642 (N_10642,N_10559,N_10404);
and U10643 (N_10643,N_10420,N_10463);
nand U10644 (N_10644,N_10477,N_10441);
xnor U10645 (N_10645,N_10530,N_10538);
xor U10646 (N_10646,N_10508,N_10450);
nand U10647 (N_10647,N_10446,N_10481);
nor U10648 (N_10648,N_10448,N_10444);
xor U10649 (N_10649,N_10558,N_10507);
nor U10650 (N_10650,N_10429,N_10441);
xor U10651 (N_10651,N_10525,N_10414);
nand U10652 (N_10652,N_10531,N_10453);
nand U10653 (N_10653,N_10542,N_10430);
or U10654 (N_10654,N_10537,N_10526);
or U10655 (N_10655,N_10559,N_10446);
or U10656 (N_10656,N_10457,N_10488);
or U10657 (N_10657,N_10419,N_10471);
and U10658 (N_10658,N_10558,N_10496);
or U10659 (N_10659,N_10451,N_10464);
xnor U10660 (N_10660,N_10521,N_10520);
xnor U10661 (N_10661,N_10417,N_10437);
nand U10662 (N_10662,N_10483,N_10551);
xnor U10663 (N_10663,N_10544,N_10555);
nand U10664 (N_10664,N_10423,N_10413);
nor U10665 (N_10665,N_10528,N_10496);
and U10666 (N_10666,N_10559,N_10451);
and U10667 (N_10667,N_10533,N_10551);
xor U10668 (N_10668,N_10405,N_10401);
nor U10669 (N_10669,N_10454,N_10460);
nand U10670 (N_10670,N_10447,N_10488);
and U10671 (N_10671,N_10543,N_10413);
nor U10672 (N_10672,N_10519,N_10406);
nor U10673 (N_10673,N_10427,N_10502);
or U10674 (N_10674,N_10525,N_10546);
or U10675 (N_10675,N_10506,N_10409);
nor U10676 (N_10676,N_10513,N_10484);
nor U10677 (N_10677,N_10470,N_10442);
and U10678 (N_10678,N_10491,N_10426);
nand U10679 (N_10679,N_10439,N_10471);
xnor U10680 (N_10680,N_10449,N_10432);
nor U10681 (N_10681,N_10509,N_10506);
or U10682 (N_10682,N_10440,N_10425);
xnor U10683 (N_10683,N_10551,N_10487);
and U10684 (N_10684,N_10437,N_10422);
or U10685 (N_10685,N_10426,N_10469);
or U10686 (N_10686,N_10493,N_10452);
or U10687 (N_10687,N_10450,N_10559);
nor U10688 (N_10688,N_10440,N_10543);
or U10689 (N_10689,N_10470,N_10552);
nor U10690 (N_10690,N_10537,N_10425);
or U10691 (N_10691,N_10533,N_10485);
xor U10692 (N_10692,N_10467,N_10525);
or U10693 (N_10693,N_10497,N_10541);
and U10694 (N_10694,N_10434,N_10506);
nand U10695 (N_10695,N_10491,N_10446);
nand U10696 (N_10696,N_10546,N_10544);
and U10697 (N_10697,N_10415,N_10430);
or U10698 (N_10698,N_10510,N_10531);
nor U10699 (N_10699,N_10427,N_10512);
nor U10700 (N_10700,N_10401,N_10437);
nand U10701 (N_10701,N_10403,N_10447);
nor U10702 (N_10702,N_10539,N_10500);
or U10703 (N_10703,N_10406,N_10555);
nor U10704 (N_10704,N_10488,N_10548);
nand U10705 (N_10705,N_10450,N_10539);
nand U10706 (N_10706,N_10454,N_10537);
and U10707 (N_10707,N_10486,N_10558);
and U10708 (N_10708,N_10535,N_10516);
and U10709 (N_10709,N_10458,N_10523);
nor U10710 (N_10710,N_10482,N_10491);
xor U10711 (N_10711,N_10502,N_10512);
nor U10712 (N_10712,N_10470,N_10406);
and U10713 (N_10713,N_10444,N_10521);
nor U10714 (N_10714,N_10461,N_10435);
nand U10715 (N_10715,N_10473,N_10534);
and U10716 (N_10716,N_10559,N_10489);
nand U10717 (N_10717,N_10434,N_10425);
nor U10718 (N_10718,N_10535,N_10406);
or U10719 (N_10719,N_10463,N_10419);
nor U10720 (N_10720,N_10563,N_10666);
nand U10721 (N_10721,N_10592,N_10694);
or U10722 (N_10722,N_10618,N_10639);
or U10723 (N_10723,N_10638,N_10613);
xor U10724 (N_10724,N_10573,N_10669);
xnor U10725 (N_10725,N_10603,N_10675);
or U10726 (N_10726,N_10568,N_10567);
or U10727 (N_10727,N_10649,N_10579);
nand U10728 (N_10728,N_10598,N_10619);
or U10729 (N_10729,N_10577,N_10702);
or U10730 (N_10730,N_10691,N_10647);
and U10731 (N_10731,N_10695,N_10692);
and U10732 (N_10732,N_10597,N_10687);
nor U10733 (N_10733,N_10654,N_10585);
or U10734 (N_10734,N_10688,N_10587);
or U10735 (N_10735,N_10630,N_10662);
or U10736 (N_10736,N_10710,N_10718);
xor U10737 (N_10737,N_10594,N_10571);
xnor U10738 (N_10738,N_10665,N_10679);
nor U10739 (N_10739,N_10623,N_10609);
xor U10740 (N_10740,N_10570,N_10709);
xor U10741 (N_10741,N_10670,N_10705);
xnor U10742 (N_10742,N_10651,N_10655);
nand U10743 (N_10743,N_10605,N_10578);
or U10744 (N_10744,N_10667,N_10606);
and U10745 (N_10745,N_10624,N_10690);
and U10746 (N_10746,N_10706,N_10676);
nor U10747 (N_10747,N_10633,N_10627);
xnor U10748 (N_10748,N_10696,N_10574);
nand U10749 (N_10749,N_10614,N_10652);
or U10750 (N_10750,N_10715,N_10714);
and U10751 (N_10751,N_10678,N_10712);
and U10752 (N_10752,N_10707,N_10608);
or U10753 (N_10753,N_10693,N_10634);
or U10754 (N_10754,N_10615,N_10560);
nor U10755 (N_10755,N_10628,N_10663);
nand U10756 (N_10756,N_10717,N_10644);
xor U10757 (N_10757,N_10704,N_10565);
nor U10758 (N_10758,N_10575,N_10607);
nand U10759 (N_10759,N_10599,N_10672);
xor U10760 (N_10760,N_10617,N_10631);
and U10761 (N_10761,N_10686,N_10586);
and U10762 (N_10762,N_10700,N_10610);
nand U10763 (N_10763,N_10659,N_10641);
nor U10764 (N_10764,N_10581,N_10648);
and U10765 (N_10765,N_10658,N_10602);
nor U10766 (N_10766,N_10682,N_10632);
xnor U10767 (N_10767,N_10650,N_10697);
nor U10768 (N_10768,N_10640,N_10699);
nor U10769 (N_10769,N_10681,N_10561);
xnor U10770 (N_10770,N_10626,N_10685);
and U10771 (N_10771,N_10572,N_10595);
xor U10772 (N_10772,N_10645,N_10677);
xnor U10773 (N_10773,N_10698,N_10564);
or U10774 (N_10774,N_10620,N_10569);
or U10775 (N_10775,N_10566,N_10683);
and U10776 (N_10776,N_10576,N_10593);
nand U10777 (N_10777,N_10590,N_10562);
nand U10778 (N_10778,N_10680,N_10622);
and U10779 (N_10779,N_10674,N_10635);
and U10780 (N_10780,N_10661,N_10642);
and U10781 (N_10781,N_10583,N_10604);
nand U10782 (N_10782,N_10657,N_10591);
nor U10783 (N_10783,N_10684,N_10671);
xor U10784 (N_10784,N_10582,N_10637);
and U10785 (N_10785,N_10673,N_10708);
xnor U10786 (N_10786,N_10713,N_10646);
nand U10787 (N_10787,N_10664,N_10703);
and U10788 (N_10788,N_10711,N_10716);
or U10789 (N_10789,N_10611,N_10689);
xor U10790 (N_10790,N_10616,N_10653);
nor U10791 (N_10791,N_10656,N_10621);
and U10792 (N_10792,N_10600,N_10636);
xnor U10793 (N_10793,N_10601,N_10580);
nor U10794 (N_10794,N_10643,N_10588);
or U10795 (N_10795,N_10660,N_10625);
nor U10796 (N_10796,N_10719,N_10612);
nor U10797 (N_10797,N_10589,N_10668);
or U10798 (N_10798,N_10629,N_10701);
and U10799 (N_10799,N_10584,N_10596);
or U10800 (N_10800,N_10662,N_10635);
xnor U10801 (N_10801,N_10588,N_10666);
and U10802 (N_10802,N_10708,N_10610);
or U10803 (N_10803,N_10705,N_10601);
and U10804 (N_10804,N_10693,N_10701);
nand U10805 (N_10805,N_10709,N_10688);
xnor U10806 (N_10806,N_10658,N_10674);
and U10807 (N_10807,N_10701,N_10643);
nand U10808 (N_10808,N_10712,N_10569);
nand U10809 (N_10809,N_10646,N_10647);
nor U10810 (N_10810,N_10718,N_10614);
and U10811 (N_10811,N_10602,N_10661);
or U10812 (N_10812,N_10576,N_10603);
nor U10813 (N_10813,N_10637,N_10719);
nand U10814 (N_10814,N_10593,N_10660);
nor U10815 (N_10815,N_10598,N_10577);
or U10816 (N_10816,N_10664,N_10679);
and U10817 (N_10817,N_10692,N_10630);
nor U10818 (N_10818,N_10705,N_10591);
nand U10819 (N_10819,N_10574,N_10589);
and U10820 (N_10820,N_10639,N_10591);
or U10821 (N_10821,N_10689,N_10613);
nand U10822 (N_10822,N_10583,N_10601);
nor U10823 (N_10823,N_10684,N_10615);
nor U10824 (N_10824,N_10641,N_10709);
and U10825 (N_10825,N_10661,N_10698);
or U10826 (N_10826,N_10674,N_10564);
xor U10827 (N_10827,N_10595,N_10619);
nand U10828 (N_10828,N_10627,N_10638);
nand U10829 (N_10829,N_10715,N_10648);
nand U10830 (N_10830,N_10611,N_10596);
and U10831 (N_10831,N_10691,N_10611);
nand U10832 (N_10832,N_10604,N_10571);
and U10833 (N_10833,N_10698,N_10560);
nor U10834 (N_10834,N_10591,N_10674);
nor U10835 (N_10835,N_10564,N_10654);
nor U10836 (N_10836,N_10660,N_10697);
nand U10837 (N_10837,N_10694,N_10688);
nor U10838 (N_10838,N_10675,N_10563);
or U10839 (N_10839,N_10567,N_10573);
xor U10840 (N_10840,N_10669,N_10701);
nor U10841 (N_10841,N_10639,N_10640);
and U10842 (N_10842,N_10595,N_10691);
nor U10843 (N_10843,N_10590,N_10583);
nor U10844 (N_10844,N_10628,N_10688);
nor U10845 (N_10845,N_10632,N_10578);
and U10846 (N_10846,N_10567,N_10560);
nand U10847 (N_10847,N_10647,N_10686);
or U10848 (N_10848,N_10646,N_10660);
nor U10849 (N_10849,N_10610,N_10661);
and U10850 (N_10850,N_10679,N_10632);
xnor U10851 (N_10851,N_10681,N_10674);
nor U10852 (N_10852,N_10649,N_10638);
xnor U10853 (N_10853,N_10630,N_10578);
or U10854 (N_10854,N_10675,N_10717);
nand U10855 (N_10855,N_10621,N_10674);
or U10856 (N_10856,N_10698,N_10691);
and U10857 (N_10857,N_10705,N_10565);
and U10858 (N_10858,N_10674,N_10714);
or U10859 (N_10859,N_10568,N_10704);
nor U10860 (N_10860,N_10621,N_10709);
and U10861 (N_10861,N_10617,N_10702);
nand U10862 (N_10862,N_10592,N_10641);
nor U10863 (N_10863,N_10569,N_10644);
and U10864 (N_10864,N_10647,N_10656);
nor U10865 (N_10865,N_10686,N_10652);
or U10866 (N_10866,N_10606,N_10697);
nor U10867 (N_10867,N_10578,N_10624);
nor U10868 (N_10868,N_10627,N_10696);
or U10869 (N_10869,N_10634,N_10711);
and U10870 (N_10870,N_10598,N_10581);
xor U10871 (N_10871,N_10625,N_10659);
xnor U10872 (N_10872,N_10577,N_10603);
xor U10873 (N_10873,N_10565,N_10702);
xnor U10874 (N_10874,N_10711,N_10561);
xor U10875 (N_10875,N_10614,N_10688);
nor U10876 (N_10876,N_10619,N_10646);
nand U10877 (N_10877,N_10688,N_10643);
or U10878 (N_10878,N_10597,N_10569);
and U10879 (N_10879,N_10647,N_10632);
nand U10880 (N_10880,N_10866,N_10733);
xnor U10881 (N_10881,N_10849,N_10778);
nor U10882 (N_10882,N_10731,N_10856);
nand U10883 (N_10883,N_10785,N_10762);
or U10884 (N_10884,N_10875,N_10831);
nand U10885 (N_10885,N_10734,N_10729);
or U10886 (N_10886,N_10868,N_10863);
nand U10887 (N_10887,N_10823,N_10828);
nor U10888 (N_10888,N_10877,N_10844);
or U10889 (N_10889,N_10801,N_10737);
or U10890 (N_10890,N_10857,N_10878);
and U10891 (N_10891,N_10821,N_10783);
nand U10892 (N_10892,N_10841,N_10855);
nand U10893 (N_10893,N_10832,N_10755);
nor U10894 (N_10894,N_10790,N_10776);
xnor U10895 (N_10895,N_10772,N_10787);
and U10896 (N_10896,N_10767,N_10822);
xor U10897 (N_10897,N_10846,N_10759);
xor U10898 (N_10898,N_10774,N_10869);
xnor U10899 (N_10899,N_10725,N_10824);
xor U10900 (N_10900,N_10751,N_10839);
or U10901 (N_10901,N_10808,N_10728);
and U10902 (N_10902,N_10835,N_10840);
and U10903 (N_10903,N_10813,N_10848);
or U10904 (N_10904,N_10852,N_10757);
nor U10905 (N_10905,N_10815,N_10872);
nor U10906 (N_10906,N_10876,N_10853);
xnor U10907 (N_10907,N_10739,N_10789);
and U10908 (N_10908,N_10804,N_10825);
nand U10909 (N_10909,N_10740,N_10721);
nor U10910 (N_10910,N_10727,N_10742);
nor U10911 (N_10911,N_10837,N_10793);
nor U10912 (N_10912,N_10847,N_10761);
xor U10913 (N_10913,N_10756,N_10810);
xor U10914 (N_10914,N_10879,N_10748);
nor U10915 (N_10915,N_10747,N_10765);
nor U10916 (N_10916,N_10838,N_10780);
xnor U10917 (N_10917,N_10809,N_10760);
nand U10918 (N_10918,N_10792,N_10750);
or U10919 (N_10919,N_10854,N_10842);
nor U10920 (N_10920,N_10732,N_10766);
and U10921 (N_10921,N_10830,N_10867);
or U10922 (N_10922,N_10749,N_10743);
xor U10923 (N_10923,N_10850,N_10771);
and U10924 (N_10924,N_10738,N_10769);
xor U10925 (N_10925,N_10795,N_10741);
nand U10926 (N_10926,N_10812,N_10758);
nand U10927 (N_10927,N_10799,N_10768);
nor U10928 (N_10928,N_10827,N_10735);
or U10929 (N_10929,N_10797,N_10820);
and U10930 (N_10930,N_10843,N_10826);
nor U10931 (N_10931,N_10802,N_10816);
and U10932 (N_10932,N_10775,N_10818);
and U10933 (N_10933,N_10752,N_10720);
xnor U10934 (N_10934,N_10834,N_10745);
nor U10935 (N_10935,N_10798,N_10833);
and U10936 (N_10936,N_10858,N_10817);
nor U10937 (N_10937,N_10754,N_10746);
nand U10938 (N_10938,N_10773,N_10811);
nor U10939 (N_10939,N_10806,N_10845);
or U10940 (N_10940,N_10814,N_10861);
and U10941 (N_10941,N_10851,N_10794);
or U10942 (N_10942,N_10803,N_10836);
or U10943 (N_10943,N_10796,N_10807);
nor U10944 (N_10944,N_10784,N_10873);
or U10945 (N_10945,N_10744,N_10724);
nor U10946 (N_10946,N_10859,N_10753);
nor U10947 (N_10947,N_10730,N_10781);
or U10948 (N_10948,N_10722,N_10865);
xor U10949 (N_10949,N_10763,N_10726);
nand U10950 (N_10950,N_10779,N_10819);
xnor U10951 (N_10951,N_10770,N_10864);
nor U10952 (N_10952,N_10788,N_10764);
or U10953 (N_10953,N_10860,N_10791);
xor U10954 (N_10954,N_10723,N_10800);
xor U10955 (N_10955,N_10777,N_10871);
nor U10956 (N_10956,N_10874,N_10805);
or U10957 (N_10957,N_10736,N_10870);
nand U10958 (N_10958,N_10862,N_10829);
nor U10959 (N_10959,N_10782,N_10786);
nor U10960 (N_10960,N_10779,N_10822);
xnor U10961 (N_10961,N_10851,N_10874);
or U10962 (N_10962,N_10795,N_10866);
or U10963 (N_10963,N_10723,N_10721);
or U10964 (N_10964,N_10727,N_10786);
nor U10965 (N_10965,N_10792,N_10808);
xor U10966 (N_10966,N_10822,N_10745);
nor U10967 (N_10967,N_10859,N_10798);
nand U10968 (N_10968,N_10811,N_10797);
or U10969 (N_10969,N_10798,N_10721);
and U10970 (N_10970,N_10804,N_10733);
xnor U10971 (N_10971,N_10763,N_10757);
nor U10972 (N_10972,N_10770,N_10720);
xor U10973 (N_10973,N_10760,N_10845);
or U10974 (N_10974,N_10793,N_10832);
nor U10975 (N_10975,N_10843,N_10758);
or U10976 (N_10976,N_10784,N_10810);
nand U10977 (N_10977,N_10745,N_10809);
nor U10978 (N_10978,N_10854,N_10723);
and U10979 (N_10979,N_10733,N_10756);
and U10980 (N_10980,N_10728,N_10748);
nand U10981 (N_10981,N_10783,N_10867);
xnor U10982 (N_10982,N_10734,N_10874);
nand U10983 (N_10983,N_10781,N_10838);
xnor U10984 (N_10984,N_10813,N_10835);
nor U10985 (N_10985,N_10853,N_10750);
nand U10986 (N_10986,N_10843,N_10762);
nor U10987 (N_10987,N_10815,N_10749);
and U10988 (N_10988,N_10795,N_10734);
or U10989 (N_10989,N_10868,N_10764);
and U10990 (N_10990,N_10799,N_10766);
nor U10991 (N_10991,N_10832,N_10760);
xnor U10992 (N_10992,N_10813,N_10740);
and U10993 (N_10993,N_10743,N_10766);
and U10994 (N_10994,N_10758,N_10779);
or U10995 (N_10995,N_10754,N_10812);
nand U10996 (N_10996,N_10764,N_10879);
nor U10997 (N_10997,N_10864,N_10780);
nand U10998 (N_10998,N_10852,N_10721);
and U10999 (N_10999,N_10809,N_10807);
xnor U11000 (N_11000,N_10795,N_10761);
or U11001 (N_11001,N_10850,N_10745);
xor U11002 (N_11002,N_10729,N_10764);
and U11003 (N_11003,N_10793,N_10772);
xnor U11004 (N_11004,N_10857,N_10842);
xnor U11005 (N_11005,N_10850,N_10775);
and U11006 (N_11006,N_10844,N_10724);
or U11007 (N_11007,N_10773,N_10755);
and U11008 (N_11008,N_10802,N_10778);
xnor U11009 (N_11009,N_10829,N_10749);
nand U11010 (N_11010,N_10766,N_10844);
xor U11011 (N_11011,N_10837,N_10818);
nand U11012 (N_11012,N_10846,N_10821);
or U11013 (N_11013,N_10756,N_10845);
nand U11014 (N_11014,N_10860,N_10748);
or U11015 (N_11015,N_10786,N_10734);
nand U11016 (N_11016,N_10835,N_10785);
or U11017 (N_11017,N_10766,N_10875);
nand U11018 (N_11018,N_10850,N_10746);
xor U11019 (N_11019,N_10814,N_10782);
nor U11020 (N_11020,N_10751,N_10831);
or U11021 (N_11021,N_10874,N_10803);
xnor U11022 (N_11022,N_10838,N_10728);
and U11023 (N_11023,N_10813,N_10730);
or U11024 (N_11024,N_10818,N_10823);
and U11025 (N_11025,N_10790,N_10866);
nor U11026 (N_11026,N_10767,N_10819);
nor U11027 (N_11027,N_10828,N_10824);
nor U11028 (N_11028,N_10794,N_10754);
xnor U11029 (N_11029,N_10724,N_10839);
and U11030 (N_11030,N_10791,N_10789);
xor U11031 (N_11031,N_10873,N_10731);
and U11032 (N_11032,N_10843,N_10787);
or U11033 (N_11033,N_10729,N_10841);
nor U11034 (N_11034,N_10854,N_10872);
and U11035 (N_11035,N_10836,N_10826);
nor U11036 (N_11036,N_10862,N_10866);
xnor U11037 (N_11037,N_10843,N_10806);
nor U11038 (N_11038,N_10820,N_10851);
nand U11039 (N_11039,N_10730,N_10842);
xnor U11040 (N_11040,N_11032,N_10974);
xor U11041 (N_11041,N_10933,N_11018);
nor U11042 (N_11042,N_10915,N_10952);
or U11043 (N_11043,N_10927,N_10993);
xor U11044 (N_11044,N_10978,N_10890);
nand U11045 (N_11045,N_10953,N_10912);
or U11046 (N_11046,N_10976,N_10884);
nor U11047 (N_11047,N_10997,N_10958);
nand U11048 (N_11048,N_10956,N_11012);
nand U11049 (N_11049,N_10977,N_10896);
nand U11050 (N_11050,N_11011,N_10911);
nand U11051 (N_11051,N_11010,N_10969);
nand U11052 (N_11052,N_10960,N_10889);
and U11053 (N_11053,N_10981,N_10972);
or U11054 (N_11054,N_11008,N_10880);
and U11055 (N_11055,N_10948,N_10916);
nand U11056 (N_11056,N_10973,N_10982);
and U11057 (N_11057,N_11000,N_11013);
and U11058 (N_11058,N_10954,N_11037);
nand U11059 (N_11059,N_10907,N_10934);
xnor U11060 (N_11060,N_10910,N_10996);
xnor U11061 (N_11061,N_10900,N_10888);
and U11062 (N_11062,N_10945,N_10897);
or U11063 (N_11063,N_10968,N_10930);
or U11064 (N_11064,N_11034,N_10929);
nand U11065 (N_11065,N_10965,N_10946);
nand U11066 (N_11066,N_10939,N_10931);
or U11067 (N_11067,N_10938,N_10892);
and U11068 (N_11068,N_10923,N_10921);
and U11069 (N_11069,N_11038,N_10963);
nor U11070 (N_11070,N_10999,N_10899);
or U11071 (N_11071,N_10898,N_11014);
nand U11072 (N_11072,N_10883,N_10971);
or U11073 (N_11073,N_10951,N_10904);
nor U11074 (N_11074,N_11026,N_10935);
xnor U11075 (N_11075,N_10881,N_10885);
nor U11076 (N_11076,N_10909,N_10949);
xor U11077 (N_11077,N_10959,N_11022);
nor U11078 (N_11078,N_10895,N_11015);
nand U11079 (N_11079,N_11004,N_11035);
nor U11080 (N_11080,N_10922,N_10924);
nand U11081 (N_11081,N_10962,N_10919);
xor U11082 (N_11082,N_10928,N_10955);
and U11083 (N_11083,N_10998,N_10992);
nand U11084 (N_11084,N_10925,N_11023);
xnor U11085 (N_11085,N_11017,N_10942);
and U11086 (N_11086,N_10891,N_11021);
nand U11087 (N_11087,N_10970,N_11025);
xor U11088 (N_11088,N_10991,N_10914);
and U11089 (N_11089,N_10920,N_10882);
nor U11090 (N_11090,N_10943,N_10966);
nand U11091 (N_11091,N_11009,N_11006);
xor U11092 (N_11092,N_11007,N_11028);
and U11093 (N_11093,N_11005,N_10988);
xor U11094 (N_11094,N_10918,N_10886);
and U11095 (N_11095,N_10980,N_11029);
or U11096 (N_11096,N_10979,N_11002);
nor U11097 (N_11097,N_10936,N_10903);
or U11098 (N_11098,N_11030,N_10961);
and U11099 (N_11099,N_10901,N_11039);
xor U11100 (N_11100,N_10950,N_10893);
and U11101 (N_11101,N_10987,N_11024);
or U11102 (N_11102,N_11001,N_10905);
or U11103 (N_11103,N_10941,N_10964);
or U11104 (N_11104,N_10887,N_10926);
nand U11105 (N_11105,N_10989,N_10986);
xnor U11106 (N_11106,N_10894,N_11033);
nand U11107 (N_11107,N_10994,N_10913);
nor U11108 (N_11108,N_10902,N_10984);
and U11109 (N_11109,N_10967,N_11036);
nand U11110 (N_11110,N_10937,N_11016);
nor U11111 (N_11111,N_10917,N_10995);
nand U11112 (N_11112,N_10957,N_10990);
and U11113 (N_11113,N_11027,N_10985);
or U11114 (N_11114,N_10975,N_11020);
and U11115 (N_11115,N_10932,N_11003);
nor U11116 (N_11116,N_11031,N_10906);
nor U11117 (N_11117,N_10940,N_10983);
xnor U11118 (N_11118,N_10947,N_10944);
nand U11119 (N_11119,N_11019,N_10908);
nor U11120 (N_11120,N_11016,N_11029);
or U11121 (N_11121,N_10914,N_10953);
nor U11122 (N_11122,N_11007,N_10982);
nand U11123 (N_11123,N_10934,N_11003);
nor U11124 (N_11124,N_10951,N_10912);
xor U11125 (N_11125,N_10896,N_11036);
nor U11126 (N_11126,N_10895,N_10931);
nor U11127 (N_11127,N_10991,N_10882);
and U11128 (N_11128,N_10991,N_10888);
or U11129 (N_11129,N_10957,N_10907);
or U11130 (N_11130,N_11013,N_10940);
and U11131 (N_11131,N_10979,N_10890);
or U11132 (N_11132,N_10915,N_10916);
nand U11133 (N_11133,N_10984,N_10945);
and U11134 (N_11134,N_10954,N_10904);
xnor U11135 (N_11135,N_10896,N_11007);
nand U11136 (N_11136,N_11009,N_10893);
and U11137 (N_11137,N_11010,N_10955);
nor U11138 (N_11138,N_10902,N_11018);
nor U11139 (N_11139,N_10947,N_11037);
nand U11140 (N_11140,N_10885,N_10937);
nor U11141 (N_11141,N_10966,N_10956);
or U11142 (N_11142,N_10930,N_10984);
xor U11143 (N_11143,N_10941,N_10916);
and U11144 (N_11144,N_10887,N_10935);
xnor U11145 (N_11145,N_10938,N_10936);
xnor U11146 (N_11146,N_10956,N_10893);
nor U11147 (N_11147,N_11019,N_11006);
and U11148 (N_11148,N_10915,N_10950);
nand U11149 (N_11149,N_10924,N_10945);
and U11150 (N_11150,N_10958,N_10978);
or U11151 (N_11151,N_10934,N_10951);
xnor U11152 (N_11152,N_11039,N_10980);
or U11153 (N_11153,N_10961,N_10927);
nor U11154 (N_11154,N_10906,N_11030);
and U11155 (N_11155,N_10883,N_11038);
and U11156 (N_11156,N_10948,N_10880);
xor U11157 (N_11157,N_10933,N_11015);
xor U11158 (N_11158,N_10994,N_10910);
and U11159 (N_11159,N_10973,N_10909);
xnor U11160 (N_11160,N_11026,N_10984);
nor U11161 (N_11161,N_10994,N_10970);
xnor U11162 (N_11162,N_10996,N_11023);
nand U11163 (N_11163,N_10981,N_10991);
nor U11164 (N_11164,N_11018,N_11016);
and U11165 (N_11165,N_11030,N_10956);
and U11166 (N_11166,N_10888,N_10979);
or U11167 (N_11167,N_11034,N_11003);
xnor U11168 (N_11168,N_10983,N_10888);
and U11169 (N_11169,N_10891,N_10884);
xnor U11170 (N_11170,N_10952,N_10951);
xor U11171 (N_11171,N_10988,N_10995);
nor U11172 (N_11172,N_10939,N_10948);
and U11173 (N_11173,N_11025,N_10953);
or U11174 (N_11174,N_11029,N_10921);
and U11175 (N_11175,N_10990,N_10953);
and U11176 (N_11176,N_10980,N_10933);
nand U11177 (N_11177,N_10964,N_10999);
and U11178 (N_11178,N_10960,N_10888);
nor U11179 (N_11179,N_10953,N_10963);
or U11180 (N_11180,N_10944,N_10892);
or U11181 (N_11181,N_11007,N_10997);
xnor U11182 (N_11182,N_10895,N_10949);
and U11183 (N_11183,N_10893,N_10912);
and U11184 (N_11184,N_10882,N_10942);
nor U11185 (N_11185,N_10980,N_11016);
or U11186 (N_11186,N_10965,N_10910);
nand U11187 (N_11187,N_11016,N_11004);
nor U11188 (N_11188,N_10986,N_10920);
or U11189 (N_11189,N_10895,N_11031);
and U11190 (N_11190,N_10980,N_10936);
nor U11191 (N_11191,N_10999,N_10959);
or U11192 (N_11192,N_10911,N_10999);
xnor U11193 (N_11193,N_10986,N_11031);
and U11194 (N_11194,N_10905,N_10961);
xnor U11195 (N_11195,N_10968,N_11032);
xnor U11196 (N_11196,N_10929,N_10887);
and U11197 (N_11197,N_10960,N_10919);
and U11198 (N_11198,N_11008,N_10912);
and U11199 (N_11199,N_10906,N_11020);
or U11200 (N_11200,N_11077,N_11195);
or U11201 (N_11201,N_11151,N_11090);
xor U11202 (N_11202,N_11115,N_11066);
or U11203 (N_11203,N_11169,N_11104);
nor U11204 (N_11204,N_11172,N_11101);
and U11205 (N_11205,N_11046,N_11041);
or U11206 (N_11206,N_11106,N_11160);
or U11207 (N_11207,N_11196,N_11154);
nand U11208 (N_11208,N_11109,N_11052);
or U11209 (N_11209,N_11087,N_11163);
and U11210 (N_11210,N_11111,N_11059);
xor U11211 (N_11211,N_11141,N_11187);
nand U11212 (N_11212,N_11194,N_11110);
or U11213 (N_11213,N_11074,N_11085);
xnor U11214 (N_11214,N_11197,N_11124);
and U11215 (N_11215,N_11153,N_11050);
nand U11216 (N_11216,N_11045,N_11072);
and U11217 (N_11217,N_11136,N_11135);
or U11218 (N_11218,N_11152,N_11150);
xnor U11219 (N_11219,N_11155,N_11058);
nor U11220 (N_11220,N_11182,N_11061);
nand U11221 (N_11221,N_11047,N_11137);
nand U11222 (N_11222,N_11100,N_11130);
nor U11223 (N_11223,N_11145,N_11185);
and U11224 (N_11224,N_11198,N_11044);
xnor U11225 (N_11225,N_11177,N_11147);
and U11226 (N_11226,N_11113,N_11120);
xnor U11227 (N_11227,N_11125,N_11088);
xor U11228 (N_11228,N_11099,N_11096);
nand U11229 (N_11229,N_11092,N_11083);
nor U11230 (N_11230,N_11138,N_11078);
or U11231 (N_11231,N_11091,N_11123);
and U11232 (N_11232,N_11127,N_11089);
xor U11233 (N_11233,N_11054,N_11057);
and U11234 (N_11234,N_11042,N_11128);
or U11235 (N_11235,N_11093,N_11076);
and U11236 (N_11236,N_11180,N_11073);
nand U11237 (N_11237,N_11188,N_11064);
nor U11238 (N_11238,N_11112,N_11049);
xor U11239 (N_11239,N_11065,N_11134);
xnor U11240 (N_11240,N_11040,N_11149);
xnor U11241 (N_11241,N_11055,N_11114);
or U11242 (N_11242,N_11159,N_11157);
and U11243 (N_11243,N_11139,N_11082);
nor U11244 (N_11244,N_11133,N_11164);
nor U11245 (N_11245,N_11166,N_11170);
and U11246 (N_11246,N_11080,N_11118);
nor U11247 (N_11247,N_11097,N_11146);
nor U11248 (N_11248,N_11084,N_11189);
nand U11249 (N_11249,N_11165,N_11167);
or U11250 (N_11250,N_11119,N_11094);
and U11251 (N_11251,N_11131,N_11086);
and U11252 (N_11252,N_11148,N_11043);
nor U11253 (N_11253,N_11105,N_11116);
nor U11254 (N_11254,N_11081,N_11122);
and U11255 (N_11255,N_11174,N_11102);
nor U11256 (N_11256,N_11095,N_11068);
and U11257 (N_11257,N_11190,N_11056);
nand U11258 (N_11258,N_11142,N_11184);
and U11259 (N_11259,N_11140,N_11062);
or U11260 (N_11260,N_11179,N_11098);
or U11261 (N_11261,N_11144,N_11191);
and U11262 (N_11262,N_11143,N_11156);
nand U11263 (N_11263,N_11126,N_11075);
and U11264 (N_11264,N_11199,N_11186);
and U11265 (N_11265,N_11070,N_11168);
nand U11266 (N_11266,N_11067,N_11053);
xnor U11267 (N_11267,N_11060,N_11051);
xor U11268 (N_11268,N_11158,N_11181);
and U11269 (N_11269,N_11117,N_11132);
and U11270 (N_11270,N_11063,N_11178);
xnor U11271 (N_11271,N_11162,N_11193);
nor U11272 (N_11272,N_11183,N_11107);
nand U11273 (N_11273,N_11192,N_11103);
nor U11274 (N_11274,N_11108,N_11173);
xor U11275 (N_11275,N_11079,N_11176);
nor U11276 (N_11276,N_11175,N_11048);
nor U11277 (N_11277,N_11069,N_11171);
nand U11278 (N_11278,N_11161,N_11121);
and U11279 (N_11279,N_11071,N_11129);
nand U11280 (N_11280,N_11041,N_11186);
nor U11281 (N_11281,N_11068,N_11041);
xor U11282 (N_11282,N_11175,N_11093);
xor U11283 (N_11283,N_11184,N_11180);
and U11284 (N_11284,N_11072,N_11075);
nand U11285 (N_11285,N_11155,N_11078);
nor U11286 (N_11286,N_11071,N_11159);
nand U11287 (N_11287,N_11132,N_11169);
or U11288 (N_11288,N_11189,N_11055);
or U11289 (N_11289,N_11150,N_11178);
or U11290 (N_11290,N_11070,N_11069);
nor U11291 (N_11291,N_11175,N_11160);
nor U11292 (N_11292,N_11079,N_11086);
nor U11293 (N_11293,N_11175,N_11080);
nand U11294 (N_11294,N_11088,N_11072);
and U11295 (N_11295,N_11054,N_11184);
xnor U11296 (N_11296,N_11144,N_11178);
nor U11297 (N_11297,N_11050,N_11065);
nand U11298 (N_11298,N_11105,N_11138);
nand U11299 (N_11299,N_11177,N_11056);
nor U11300 (N_11300,N_11160,N_11050);
xnor U11301 (N_11301,N_11051,N_11159);
and U11302 (N_11302,N_11126,N_11141);
and U11303 (N_11303,N_11066,N_11190);
and U11304 (N_11304,N_11174,N_11092);
or U11305 (N_11305,N_11097,N_11133);
or U11306 (N_11306,N_11173,N_11049);
nand U11307 (N_11307,N_11121,N_11062);
nand U11308 (N_11308,N_11045,N_11172);
xnor U11309 (N_11309,N_11062,N_11175);
or U11310 (N_11310,N_11174,N_11172);
nor U11311 (N_11311,N_11154,N_11179);
and U11312 (N_11312,N_11084,N_11149);
nor U11313 (N_11313,N_11043,N_11186);
and U11314 (N_11314,N_11132,N_11145);
nand U11315 (N_11315,N_11161,N_11069);
or U11316 (N_11316,N_11154,N_11124);
and U11317 (N_11317,N_11059,N_11075);
or U11318 (N_11318,N_11175,N_11115);
nand U11319 (N_11319,N_11065,N_11042);
nand U11320 (N_11320,N_11131,N_11059);
nor U11321 (N_11321,N_11048,N_11061);
nor U11322 (N_11322,N_11076,N_11177);
nor U11323 (N_11323,N_11154,N_11158);
nor U11324 (N_11324,N_11113,N_11088);
nor U11325 (N_11325,N_11112,N_11106);
xor U11326 (N_11326,N_11189,N_11192);
and U11327 (N_11327,N_11151,N_11071);
nor U11328 (N_11328,N_11104,N_11046);
nand U11329 (N_11329,N_11145,N_11134);
xor U11330 (N_11330,N_11158,N_11086);
nand U11331 (N_11331,N_11126,N_11152);
xnor U11332 (N_11332,N_11116,N_11152);
nand U11333 (N_11333,N_11146,N_11128);
nand U11334 (N_11334,N_11119,N_11199);
or U11335 (N_11335,N_11143,N_11168);
nand U11336 (N_11336,N_11188,N_11050);
xor U11337 (N_11337,N_11053,N_11079);
nand U11338 (N_11338,N_11186,N_11144);
nand U11339 (N_11339,N_11050,N_11135);
xor U11340 (N_11340,N_11176,N_11121);
nand U11341 (N_11341,N_11184,N_11168);
nand U11342 (N_11342,N_11041,N_11069);
nand U11343 (N_11343,N_11112,N_11124);
xor U11344 (N_11344,N_11054,N_11040);
xor U11345 (N_11345,N_11089,N_11072);
or U11346 (N_11346,N_11079,N_11188);
nor U11347 (N_11347,N_11183,N_11097);
or U11348 (N_11348,N_11101,N_11130);
nand U11349 (N_11349,N_11086,N_11045);
xor U11350 (N_11350,N_11040,N_11136);
and U11351 (N_11351,N_11139,N_11155);
nand U11352 (N_11352,N_11047,N_11177);
or U11353 (N_11353,N_11131,N_11119);
xor U11354 (N_11354,N_11070,N_11090);
and U11355 (N_11355,N_11107,N_11080);
nand U11356 (N_11356,N_11077,N_11128);
nor U11357 (N_11357,N_11057,N_11151);
and U11358 (N_11358,N_11119,N_11076);
and U11359 (N_11359,N_11166,N_11172);
or U11360 (N_11360,N_11249,N_11230);
xor U11361 (N_11361,N_11241,N_11272);
or U11362 (N_11362,N_11352,N_11353);
xor U11363 (N_11363,N_11255,N_11315);
or U11364 (N_11364,N_11227,N_11330);
xnor U11365 (N_11365,N_11348,N_11321);
xor U11366 (N_11366,N_11277,N_11294);
or U11367 (N_11367,N_11295,N_11316);
or U11368 (N_11368,N_11349,N_11209);
nand U11369 (N_11369,N_11200,N_11237);
nand U11370 (N_11370,N_11344,N_11350);
nor U11371 (N_11371,N_11259,N_11318);
or U11372 (N_11372,N_11319,N_11359);
nand U11373 (N_11373,N_11236,N_11287);
nand U11374 (N_11374,N_11280,N_11358);
and U11375 (N_11375,N_11341,N_11256);
or U11376 (N_11376,N_11284,N_11307);
nor U11377 (N_11377,N_11216,N_11302);
and U11378 (N_11378,N_11323,N_11310);
nand U11379 (N_11379,N_11224,N_11311);
nor U11380 (N_11380,N_11252,N_11235);
nand U11381 (N_11381,N_11313,N_11234);
nand U11382 (N_11382,N_11312,N_11248);
and U11383 (N_11383,N_11221,N_11212);
and U11384 (N_11384,N_11297,N_11265);
or U11385 (N_11385,N_11210,N_11223);
xor U11386 (N_11386,N_11240,N_11329);
nor U11387 (N_11387,N_11276,N_11334);
and U11388 (N_11388,N_11304,N_11268);
xor U11389 (N_11389,N_11225,N_11232);
nor U11390 (N_11390,N_11260,N_11203);
and U11391 (N_11391,N_11205,N_11288);
nand U11392 (N_11392,N_11322,N_11266);
and U11393 (N_11393,N_11290,N_11245);
xor U11394 (N_11394,N_11250,N_11273);
and U11395 (N_11395,N_11242,N_11337);
or U11396 (N_11396,N_11356,N_11253);
or U11397 (N_11397,N_11305,N_11338);
nor U11398 (N_11398,N_11347,N_11296);
and U11399 (N_11399,N_11231,N_11309);
and U11400 (N_11400,N_11303,N_11326);
nor U11401 (N_11401,N_11261,N_11293);
or U11402 (N_11402,N_11208,N_11340);
nand U11403 (N_11403,N_11342,N_11264);
xor U11404 (N_11404,N_11233,N_11283);
or U11405 (N_11405,N_11324,N_11299);
nand U11406 (N_11406,N_11317,N_11239);
nand U11407 (N_11407,N_11282,N_11332);
and U11408 (N_11408,N_11269,N_11238);
and U11409 (N_11409,N_11211,N_11289);
and U11410 (N_11410,N_11247,N_11263);
or U11411 (N_11411,N_11325,N_11333);
and U11412 (N_11412,N_11251,N_11335);
xnor U11413 (N_11413,N_11343,N_11219);
and U11414 (N_11414,N_11270,N_11246);
nand U11415 (N_11415,N_11274,N_11206);
xor U11416 (N_11416,N_11327,N_11262);
xnor U11417 (N_11417,N_11218,N_11229);
or U11418 (N_11418,N_11320,N_11278);
xor U11419 (N_11419,N_11281,N_11201);
xnor U11420 (N_11420,N_11228,N_11220);
nor U11421 (N_11421,N_11254,N_11279);
and U11422 (N_11422,N_11346,N_11292);
nor U11423 (N_11423,N_11306,N_11291);
or U11424 (N_11424,N_11336,N_11213);
nor U11425 (N_11425,N_11357,N_11202);
and U11426 (N_11426,N_11300,N_11215);
nand U11427 (N_11427,N_11275,N_11257);
xor U11428 (N_11428,N_11355,N_11207);
or U11429 (N_11429,N_11226,N_11267);
nand U11430 (N_11430,N_11286,N_11258);
nor U11431 (N_11431,N_11217,N_11339);
and U11432 (N_11432,N_11222,N_11243);
xnor U11433 (N_11433,N_11271,N_11244);
xor U11434 (N_11434,N_11204,N_11285);
and U11435 (N_11435,N_11298,N_11351);
nand U11436 (N_11436,N_11331,N_11345);
xnor U11437 (N_11437,N_11314,N_11214);
nor U11438 (N_11438,N_11354,N_11328);
and U11439 (N_11439,N_11308,N_11301);
nor U11440 (N_11440,N_11300,N_11243);
nor U11441 (N_11441,N_11274,N_11310);
nor U11442 (N_11442,N_11287,N_11299);
and U11443 (N_11443,N_11207,N_11285);
nor U11444 (N_11444,N_11214,N_11247);
nand U11445 (N_11445,N_11272,N_11325);
nor U11446 (N_11446,N_11211,N_11275);
or U11447 (N_11447,N_11222,N_11247);
or U11448 (N_11448,N_11254,N_11297);
and U11449 (N_11449,N_11260,N_11251);
xnor U11450 (N_11450,N_11231,N_11306);
xnor U11451 (N_11451,N_11328,N_11357);
xnor U11452 (N_11452,N_11251,N_11283);
nand U11453 (N_11453,N_11262,N_11251);
nand U11454 (N_11454,N_11311,N_11310);
nand U11455 (N_11455,N_11256,N_11351);
xor U11456 (N_11456,N_11234,N_11246);
and U11457 (N_11457,N_11251,N_11269);
nand U11458 (N_11458,N_11317,N_11355);
nor U11459 (N_11459,N_11225,N_11221);
nor U11460 (N_11460,N_11339,N_11233);
nand U11461 (N_11461,N_11325,N_11356);
nand U11462 (N_11462,N_11338,N_11297);
or U11463 (N_11463,N_11337,N_11343);
nand U11464 (N_11464,N_11254,N_11222);
or U11465 (N_11465,N_11241,N_11206);
and U11466 (N_11466,N_11225,N_11355);
or U11467 (N_11467,N_11249,N_11210);
and U11468 (N_11468,N_11227,N_11303);
and U11469 (N_11469,N_11236,N_11329);
xnor U11470 (N_11470,N_11353,N_11324);
or U11471 (N_11471,N_11318,N_11323);
and U11472 (N_11472,N_11324,N_11316);
nand U11473 (N_11473,N_11202,N_11248);
and U11474 (N_11474,N_11312,N_11355);
xnor U11475 (N_11475,N_11346,N_11246);
nor U11476 (N_11476,N_11329,N_11249);
or U11477 (N_11477,N_11240,N_11204);
nor U11478 (N_11478,N_11291,N_11319);
xor U11479 (N_11479,N_11283,N_11294);
or U11480 (N_11480,N_11267,N_11257);
nand U11481 (N_11481,N_11347,N_11278);
xor U11482 (N_11482,N_11229,N_11305);
nand U11483 (N_11483,N_11243,N_11210);
nor U11484 (N_11484,N_11351,N_11334);
or U11485 (N_11485,N_11218,N_11316);
nand U11486 (N_11486,N_11311,N_11223);
nand U11487 (N_11487,N_11253,N_11320);
and U11488 (N_11488,N_11212,N_11339);
nor U11489 (N_11489,N_11329,N_11306);
nand U11490 (N_11490,N_11270,N_11212);
and U11491 (N_11491,N_11219,N_11274);
and U11492 (N_11492,N_11290,N_11317);
or U11493 (N_11493,N_11222,N_11345);
nand U11494 (N_11494,N_11295,N_11247);
or U11495 (N_11495,N_11234,N_11301);
nand U11496 (N_11496,N_11338,N_11251);
xor U11497 (N_11497,N_11266,N_11318);
xnor U11498 (N_11498,N_11321,N_11220);
xnor U11499 (N_11499,N_11350,N_11282);
or U11500 (N_11500,N_11235,N_11311);
nor U11501 (N_11501,N_11353,N_11337);
or U11502 (N_11502,N_11341,N_11246);
xnor U11503 (N_11503,N_11292,N_11220);
xor U11504 (N_11504,N_11218,N_11274);
nand U11505 (N_11505,N_11317,N_11222);
nor U11506 (N_11506,N_11330,N_11200);
nand U11507 (N_11507,N_11226,N_11283);
xor U11508 (N_11508,N_11207,N_11244);
nand U11509 (N_11509,N_11357,N_11222);
and U11510 (N_11510,N_11286,N_11343);
or U11511 (N_11511,N_11211,N_11213);
xnor U11512 (N_11512,N_11292,N_11203);
nand U11513 (N_11513,N_11237,N_11296);
or U11514 (N_11514,N_11238,N_11223);
xor U11515 (N_11515,N_11356,N_11298);
xnor U11516 (N_11516,N_11335,N_11228);
nor U11517 (N_11517,N_11245,N_11329);
or U11518 (N_11518,N_11209,N_11260);
or U11519 (N_11519,N_11310,N_11251);
nor U11520 (N_11520,N_11384,N_11427);
or U11521 (N_11521,N_11440,N_11387);
nor U11522 (N_11522,N_11409,N_11395);
nand U11523 (N_11523,N_11450,N_11471);
or U11524 (N_11524,N_11415,N_11375);
xnor U11525 (N_11525,N_11424,N_11422);
nand U11526 (N_11526,N_11438,N_11499);
nand U11527 (N_11527,N_11369,N_11442);
nand U11528 (N_11528,N_11452,N_11372);
or U11529 (N_11529,N_11413,N_11462);
and U11530 (N_11530,N_11461,N_11429);
nand U11531 (N_11531,N_11366,N_11410);
nand U11532 (N_11532,N_11490,N_11463);
xnor U11533 (N_11533,N_11514,N_11420);
or U11534 (N_11534,N_11382,N_11404);
xor U11535 (N_11535,N_11444,N_11393);
and U11536 (N_11536,N_11511,N_11367);
nor U11537 (N_11537,N_11371,N_11465);
or U11538 (N_11538,N_11446,N_11360);
or U11539 (N_11539,N_11458,N_11492);
nor U11540 (N_11540,N_11378,N_11428);
and U11541 (N_11541,N_11421,N_11425);
or U11542 (N_11542,N_11419,N_11518);
xor U11543 (N_11543,N_11370,N_11368);
xor U11544 (N_11544,N_11362,N_11361);
and U11545 (N_11545,N_11436,N_11397);
or U11546 (N_11546,N_11475,N_11416);
or U11547 (N_11547,N_11430,N_11487);
xnor U11548 (N_11548,N_11474,N_11480);
and U11549 (N_11549,N_11488,N_11503);
and U11550 (N_11550,N_11402,N_11407);
or U11551 (N_11551,N_11379,N_11403);
nand U11552 (N_11552,N_11512,N_11516);
and U11553 (N_11553,N_11373,N_11501);
and U11554 (N_11554,N_11449,N_11437);
and U11555 (N_11555,N_11390,N_11432);
nor U11556 (N_11556,N_11472,N_11392);
or U11557 (N_11557,N_11464,N_11401);
xor U11558 (N_11558,N_11500,N_11447);
xor U11559 (N_11559,N_11426,N_11502);
nor U11560 (N_11560,N_11376,N_11453);
nor U11561 (N_11561,N_11493,N_11494);
nand U11562 (N_11562,N_11377,N_11506);
and U11563 (N_11563,N_11431,N_11417);
xor U11564 (N_11564,N_11385,N_11510);
nand U11565 (N_11565,N_11495,N_11473);
nand U11566 (N_11566,N_11466,N_11457);
nand U11567 (N_11567,N_11505,N_11485);
nand U11568 (N_11568,N_11405,N_11406);
and U11569 (N_11569,N_11381,N_11477);
or U11570 (N_11570,N_11504,N_11414);
or U11571 (N_11571,N_11399,N_11433);
xor U11572 (N_11572,N_11398,N_11408);
nor U11573 (N_11573,N_11363,N_11411);
xnor U11574 (N_11574,N_11389,N_11445);
and U11575 (N_11575,N_11386,N_11481);
nor U11576 (N_11576,N_11455,N_11439);
or U11577 (N_11577,N_11478,N_11391);
nor U11578 (N_11578,N_11400,N_11515);
and U11579 (N_11579,N_11364,N_11508);
and U11580 (N_11580,N_11434,N_11435);
nand U11581 (N_11581,N_11470,N_11412);
nand U11582 (N_11582,N_11519,N_11467);
or U11583 (N_11583,N_11496,N_11383);
and U11584 (N_11584,N_11454,N_11468);
and U11585 (N_11585,N_11489,N_11396);
nor U11586 (N_11586,N_11476,N_11388);
and U11587 (N_11587,N_11460,N_11451);
xor U11588 (N_11588,N_11448,N_11507);
nand U11589 (N_11589,N_11497,N_11483);
nor U11590 (N_11590,N_11482,N_11459);
and U11591 (N_11591,N_11509,N_11456);
and U11592 (N_11592,N_11418,N_11394);
nand U11593 (N_11593,N_11479,N_11491);
nor U11594 (N_11594,N_11469,N_11443);
or U11595 (N_11595,N_11441,N_11498);
xor U11596 (N_11596,N_11365,N_11380);
or U11597 (N_11597,N_11374,N_11423);
nor U11598 (N_11598,N_11513,N_11484);
nor U11599 (N_11599,N_11486,N_11517);
nand U11600 (N_11600,N_11405,N_11512);
nand U11601 (N_11601,N_11372,N_11397);
xnor U11602 (N_11602,N_11438,N_11423);
xor U11603 (N_11603,N_11486,N_11483);
nand U11604 (N_11604,N_11492,N_11479);
nand U11605 (N_11605,N_11454,N_11464);
nand U11606 (N_11606,N_11414,N_11482);
xor U11607 (N_11607,N_11473,N_11366);
and U11608 (N_11608,N_11470,N_11425);
and U11609 (N_11609,N_11518,N_11380);
xnor U11610 (N_11610,N_11452,N_11485);
nor U11611 (N_11611,N_11448,N_11412);
xor U11612 (N_11612,N_11507,N_11450);
and U11613 (N_11613,N_11377,N_11446);
or U11614 (N_11614,N_11501,N_11399);
nor U11615 (N_11615,N_11421,N_11409);
and U11616 (N_11616,N_11383,N_11456);
xor U11617 (N_11617,N_11374,N_11445);
and U11618 (N_11618,N_11514,N_11438);
nor U11619 (N_11619,N_11372,N_11373);
nand U11620 (N_11620,N_11383,N_11364);
xnor U11621 (N_11621,N_11419,N_11470);
or U11622 (N_11622,N_11448,N_11427);
or U11623 (N_11623,N_11473,N_11442);
xnor U11624 (N_11624,N_11492,N_11384);
nand U11625 (N_11625,N_11454,N_11456);
nor U11626 (N_11626,N_11499,N_11444);
and U11627 (N_11627,N_11448,N_11447);
xnor U11628 (N_11628,N_11504,N_11391);
nand U11629 (N_11629,N_11500,N_11440);
or U11630 (N_11630,N_11367,N_11503);
or U11631 (N_11631,N_11424,N_11403);
nand U11632 (N_11632,N_11430,N_11433);
nand U11633 (N_11633,N_11426,N_11506);
xnor U11634 (N_11634,N_11385,N_11426);
nand U11635 (N_11635,N_11392,N_11517);
or U11636 (N_11636,N_11513,N_11500);
or U11637 (N_11637,N_11371,N_11495);
nand U11638 (N_11638,N_11510,N_11473);
xnor U11639 (N_11639,N_11509,N_11399);
nor U11640 (N_11640,N_11450,N_11382);
or U11641 (N_11641,N_11425,N_11482);
or U11642 (N_11642,N_11455,N_11511);
nand U11643 (N_11643,N_11508,N_11445);
and U11644 (N_11644,N_11459,N_11483);
nor U11645 (N_11645,N_11517,N_11363);
or U11646 (N_11646,N_11361,N_11360);
and U11647 (N_11647,N_11400,N_11506);
nor U11648 (N_11648,N_11462,N_11370);
and U11649 (N_11649,N_11504,N_11424);
nand U11650 (N_11650,N_11503,N_11397);
or U11651 (N_11651,N_11459,N_11497);
nor U11652 (N_11652,N_11466,N_11370);
and U11653 (N_11653,N_11498,N_11487);
nand U11654 (N_11654,N_11378,N_11365);
nand U11655 (N_11655,N_11417,N_11496);
and U11656 (N_11656,N_11436,N_11406);
xnor U11657 (N_11657,N_11411,N_11513);
or U11658 (N_11658,N_11393,N_11501);
xnor U11659 (N_11659,N_11366,N_11419);
xnor U11660 (N_11660,N_11437,N_11492);
or U11661 (N_11661,N_11371,N_11414);
nor U11662 (N_11662,N_11442,N_11462);
and U11663 (N_11663,N_11376,N_11463);
xor U11664 (N_11664,N_11369,N_11455);
nor U11665 (N_11665,N_11453,N_11414);
nand U11666 (N_11666,N_11380,N_11401);
xor U11667 (N_11667,N_11500,N_11417);
nand U11668 (N_11668,N_11469,N_11452);
or U11669 (N_11669,N_11511,N_11381);
or U11670 (N_11670,N_11490,N_11446);
and U11671 (N_11671,N_11401,N_11447);
or U11672 (N_11672,N_11438,N_11426);
xnor U11673 (N_11673,N_11463,N_11457);
or U11674 (N_11674,N_11397,N_11440);
and U11675 (N_11675,N_11508,N_11516);
or U11676 (N_11676,N_11361,N_11503);
nor U11677 (N_11677,N_11444,N_11493);
and U11678 (N_11678,N_11393,N_11475);
xor U11679 (N_11679,N_11449,N_11419);
or U11680 (N_11680,N_11574,N_11611);
nand U11681 (N_11681,N_11580,N_11598);
or U11682 (N_11682,N_11656,N_11567);
nor U11683 (N_11683,N_11561,N_11654);
xor U11684 (N_11684,N_11628,N_11608);
and U11685 (N_11685,N_11658,N_11660);
nor U11686 (N_11686,N_11582,N_11621);
nand U11687 (N_11687,N_11665,N_11586);
nand U11688 (N_11688,N_11570,N_11559);
xor U11689 (N_11689,N_11653,N_11637);
xor U11690 (N_11690,N_11644,N_11542);
nand U11691 (N_11691,N_11547,N_11618);
xor U11692 (N_11692,N_11594,N_11600);
or U11693 (N_11693,N_11626,N_11669);
nor U11694 (N_11694,N_11620,N_11529);
or U11695 (N_11695,N_11573,N_11655);
nand U11696 (N_11696,N_11630,N_11615);
and U11697 (N_11697,N_11604,N_11591);
and U11698 (N_11698,N_11564,N_11575);
nand U11699 (N_11699,N_11617,N_11577);
and U11700 (N_11700,N_11593,N_11581);
and U11701 (N_11701,N_11526,N_11633);
nand U11702 (N_11702,N_11651,N_11613);
nand U11703 (N_11703,N_11652,N_11554);
and U11704 (N_11704,N_11595,N_11558);
nor U11705 (N_11705,N_11556,N_11589);
nor U11706 (N_11706,N_11545,N_11670);
nor U11707 (N_11707,N_11642,N_11602);
xnor U11708 (N_11708,N_11601,N_11674);
or U11709 (N_11709,N_11555,N_11640);
nand U11710 (N_11710,N_11534,N_11678);
nor U11711 (N_11711,N_11647,N_11629);
nand U11712 (N_11712,N_11579,N_11522);
nand U11713 (N_11713,N_11540,N_11537);
or U11714 (N_11714,N_11548,N_11624);
nor U11715 (N_11715,N_11648,N_11675);
nand U11716 (N_11716,N_11557,N_11596);
or U11717 (N_11717,N_11673,N_11677);
and U11718 (N_11718,N_11523,N_11571);
and U11719 (N_11719,N_11623,N_11610);
and U11720 (N_11720,N_11532,N_11551);
xor U11721 (N_11721,N_11597,N_11657);
xnor U11722 (N_11722,N_11520,N_11546);
and U11723 (N_11723,N_11659,N_11566);
nor U11724 (N_11724,N_11576,N_11625);
nor U11725 (N_11725,N_11664,N_11614);
and U11726 (N_11726,N_11607,N_11643);
nand U11727 (N_11727,N_11544,N_11616);
xor U11728 (N_11728,N_11584,N_11627);
and U11729 (N_11729,N_11612,N_11524);
nand U11730 (N_11730,N_11638,N_11622);
nand U11731 (N_11731,N_11527,N_11631);
nand U11732 (N_11732,N_11635,N_11599);
xor U11733 (N_11733,N_11583,N_11560);
xnor U11734 (N_11734,N_11605,N_11671);
nand U11735 (N_11735,N_11578,N_11565);
xnor U11736 (N_11736,N_11645,N_11552);
xor U11737 (N_11737,N_11563,N_11585);
nand U11738 (N_11738,N_11662,N_11636);
and U11739 (N_11739,N_11592,N_11590);
xor U11740 (N_11740,N_11666,N_11533);
nand U11741 (N_11741,N_11619,N_11639);
nand U11742 (N_11742,N_11676,N_11530);
nand U11743 (N_11743,N_11606,N_11587);
nor U11744 (N_11744,N_11538,N_11641);
nand U11745 (N_11745,N_11568,N_11531);
or U11746 (N_11746,N_11528,N_11672);
nor U11747 (N_11747,N_11667,N_11541);
or U11748 (N_11748,N_11663,N_11553);
nand U11749 (N_11749,N_11634,N_11562);
and U11750 (N_11750,N_11535,N_11650);
and U11751 (N_11751,N_11543,N_11550);
and U11752 (N_11752,N_11521,N_11525);
nand U11753 (N_11753,N_11549,N_11603);
and U11754 (N_11754,N_11679,N_11661);
or U11755 (N_11755,N_11536,N_11588);
or U11756 (N_11756,N_11539,N_11646);
xnor U11757 (N_11757,N_11668,N_11572);
nor U11758 (N_11758,N_11632,N_11609);
xnor U11759 (N_11759,N_11649,N_11569);
nor U11760 (N_11760,N_11587,N_11552);
or U11761 (N_11761,N_11640,N_11666);
nand U11762 (N_11762,N_11536,N_11662);
nand U11763 (N_11763,N_11671,N_11669);
and U11764 (N_11764,N_11555,N_11625);
and U11765 (N_11765,N_11664,N_11671);
nand U11766 (N_11766,N_11597,N_11631);
nor U11767 (N_11767,N_11671,N_11557);
nor U11768 (N_11768,N_11589,N_11598);
nand U11769 (N_11769,N_11567,N_11662);
and U11770 (N_11770,N_11662,N_11583);
nand U11771 (N_11771,N_11672,N_11629);
and U11772 (N_11772,N_11571,N_11537);
nand U11773 (N_11773,N_11556,N_11616);
and U11774 (N_11774,N_11586,N_11570);
xnor U11775 (N_11775,N_11564,N_11536);
or U11776 (N_11776,N_11614,N_11567);
nor U11777 (N_11777,N_11574,N_11667);
or U11778 (N_11778,N_11563,N_11580);
xor U11779 (N_11779,N_11586,N_11649);
or U11780 (N_11780,N_11654,N_11523);
nor U11781 (N_11781,N_11560,N_11584);
and U11782 (N_11782,N_11571,N_11579);
nand U11783 (N_11783,N_11618,N_11568);
and U11784 (N_11784,N_11524,N_11630);
nand U11785 (N_11785,N_11531,N_11553);
nand U11786 (N_11786,N_11554,N_11597);
xnor U11787 (N_11787,N_11568,N_11588);
nand U11788 (N_11788,N_11606,N_11624);
xnor U11789 (N_11789,N_11566,N_11611);
nor U11790 (N_11790,N_11622,N_11582);
or U11791 (N_11791,N_11552,N_11658);
nand U11792 (N_11792,N_11541,N_11664);
nor U11793 (N_11793,N_11624,N_11546);
nand U11794 (N_11794,N_11588,N_11663);
and U11795 (N_11795,N_11606,N_11664);
and U11796 (N_11796,N_11653,N_11622);
and U11797 (N_11797,N_11650,N_11572);
nor U11798 (N_11798,N_11589,N_11539);
and U11799 (N_11799,N_11533,N_11621);
or U11800 (N_11800,N_11547,N_11552);
and U11801 (N_11801,N_11564,N_11525);
or U11802 (N_11802,N_11560,N_11576);
or U11803 (N_11803,N_11654,N_11665);
nand U11804 (N_11804,N_11595,N_11562);
and U11805 (N_11805,N_11533,N_11655);
nand U11806 (N_11806,N_11649,N_11578);
nor U11807 (N_11807,N_11635,N_11651);
xor U11808 (N_11808,N_11585,N_11612);
and U11809 (N_11809,N_11630,N_11554);
nand U11810 (N_11810,N_11612,N_11594);
and U11811 (N_11811,N_11641,N_11643);
and U11812 (N_11812,N_11594,N_11653);
nand U11813 (N_11813,N_11555,N_11599);
nand U11814 (N_11814,N_11550,N_11622);
or U11815 (N_11815,N_11623,N_11541);
xnor U11816 (N_11816,N_11563,N_11665);
and U11817 (N_11817,N_11548,N_11638);
and U11818 (N_11818,N_11648,N_11610);
nor U11819 (N_11819,N_11578,N_11610);
nor U11820 (N_11820,N_11536,N_11524);
nand U11821 (N_11821,N_11611,N_11663);
or U11822 (N_11822,N_11583,N_11552);
xor U11823 (N_11823,N_11560,N_11621);
and U11824 (N_11824,N_11619,N_11650);
and U11825 (N_11825,N_11582,N_11641);
and U11826 (N_11826,N_11594,N_11593);
or U11827 (N_11827,N_11546,N_11548);
and U11828 (N_11828,N_11581,N_11607);
nand U11829 (N_11829,N_11562,N_11643);
nor U11830 (N_11830,N_11598,N_11530);
or U11831 (N_11831,N_11595,N_11615);
xor U11832 (N_11832,N_11677,N_11668);
or U11833 (N_11833,N_11629,N_11637);
or U11834 (N_11834,N_11679,N_11667);
or U11835 (N_11835,N_11611,N_11601);
nand U11836 (N_11836,N_11611,N_11647);
or U11837 (N_11837,N_11641,N_11622);
nand U11838 (N_11838,N_11646,N_11582);
or U11839 (N_11839,N_11659,N_11648);
nand U11840 (N_11840,N_11818,N_11691);
xor U11841 (N_11841,N_11697,N_11751);
and U11842 (N_11842,N_11696,N_11733);
and U11843 (N_11843,N_11698,N_11769);
xor U11844 (N_11844,N_11794,N_11776);
nand U11845 (N_11845,N_11713,N_11762);
and U11846 (N_11846,N_11786,N_11711);
nor U11847 (N_11847,N_11832,N_11837);
nor U11848 (N_11848,N_11771,N_11739);
and U11849 (N_11849,N_11716,N_11808);
nor U11850 (N_11850,N_11759,N_11732);
or U11851 (N_11851,N_11811,N_11750);
nor U11852 (N_11852,N_11805,N_11684);
nor U11853 (N_11853,N_11815,N_11755);
xor U11854 (N_11854,N_11726,N_11825);
nand U11855 (N_11855,N_11827,N_11809);
and U11856 (N_11856,N_11694,N_11826);
xor U11857 (N_11857,N_11719,N_11753);
or U11858 (N_11858,N_11788,N_11728);
nor U11859 (N_11859,N_11816,N_11704);
and U11860 (N_11860,N_11774,N_11708);
nor U11861 (N_11861,N_11775,N_11839);
and U11862 (N_11862,N_11783,N_11767);
nand U11863 (N_11863,N_11787,N_11830);
xnor U11864 (N_11864,N_11712,N_11686);
and U11865 (N_11865,N_11798,N_11799);
xor U11866 (N_11866,N_11792,N_11810);
nand U11867 (N_11867,N_11784,N_11770);
xor U11868 (N_11868,N_11718,N_11724);
nor U11869 (N_11869,N_11829,N_11763);
and U11870 (N_11870,N_11789,N_11741);
nand U11871 (N_11871,N_11781,N_11800);
or U11872 (N_11872,N_11692,N_11779);
or U11873 (N_11873,N_11836,N_11793);
nand U11874 (N_11874,N_11831,N_11764);
and U11875 (N_11875,N_11703,N_11778);
nor U11876 (N_11876,N_11821,N_11761);
and U11877 (N_11877,N_11782,N_11828);
nor U11878 (N_11878,N_11777,N_11746);
or U11879 (N_11879,N_11700,N_11817);
nand U11880 (N_11880,N_11747,N_11699);
or U11881 (N_11881,N_11780,N_11772);
nand U11882 (N_11882,N_11785,N_11721);
nand U11883 (N_11883,N_11695,N_11680);
xor U11884 (N_11884,N_11707,N_11714);
xnor U11885 (N_11885,N_11819,N_11738);
nor U11886 (N_11886,N_11824,N_11731);
nand U11887 (N_11887,N_11814,N_11754);
nor U11888 (N_11888,N_11757,N_11802);
xor U11889 (N_11889,N_11737,N_11835);
and U11890 (N_11890,N_11822,N_11801);
and U11891 (N_11891,N_11796,N_11717);
and U11892 (N_11892,N_11742,N_11729);
and U11893 (N_11893,N_11734,N_11693);
nand U11894 (N_11894,N_11807,N_11806);
nand U11895 (N_11895,N_11790,N_11758);
nor U11896 (N_11896,N_11834,N_11683);
xnor U11897 (N_11897,N_11702,N_11773);
nor U11898 (N_11898,N_11690,N_11722);
xnor U11899 (N_11899,N_11752,N_11749);
xnor U11900 (N_11900,N_11804,N_11688);
nand U11901 (N_11901,N_11797,N_11748);
xor U11902 (N_11902,N_11820,N_11743);
nand U11903 (N_11903,N_11812,N_11689);
nand U11904 (N_11904,N_11765,N_11685);
xnor U11905 (N_11905,N_11705,N_11795);
or U11906 (N_11906,N_11720,N_11706);
nand U11907 (N_11907,N_11744,N_11681);
and U11908 (N_11908,N_11735,N_11730);
or U11909 (N_11909,N_11715,N_11803);
nand U11910 (N_11910,N_11791,N_11745);
xnor U11911 (N_11911,N_11723,N_11813);
nor U11912 (N_11912,N_11736,N_11687);
and U11913 (N_11913,N_11682,N_11823);
nor U11914 (N_11914,N_11760,N_11838);
or U11915 (N_11915,N_11768,N_11701);
xor U11916 (N_11916,N_11727,N_11766);
and U11917 (N_11917,N_11710,N_11740);
nor U11918 (N_11918,N_11833,N_11709);
or U11919 (N_11919,N_11725,N_11756);
or U11920 (N_11920,N_11726,N_11816);
xor U11921 (N_11921,N_11700,N_11720);
nor U11922 (N_11922,N_11764,N_11796);
xnor U11923 (N_11923,N_11782,N_11719);
nor U11924 (N_11924,N_11797,N_11746);
nor U11925 (N_11925,N_11834,N_11767);
xnor U11926 (N_11926,N_11795,N_11807);
nor U11927 (N_11927,N_11717,N_11708);
xor U11928 (N_11928,N_11759,N_11822);
or U11929 (N_11929,N_11754,N_11726);
nand U11930 (N_11930,N_11806,N_11737);
nor U11931 (N_11931,N_11762,N_11835);
nor U11932 (N_11932,N_11743,N_11764);
or U11933 (N_11933,N_11740,N_11777);
and U11934 (N_11934,N_11727,N_11701);
and U11935 (N_11935,N_11817,N_11766);
nor U11936 (N_11936,N_11682,N_11747);
xnor U11937 (N_11937,N_11749,N_11727);
or U11938 (N_11938,N_11704,N_11693);
xor U11939 (N_11939,N_11791,N_11714);
nand U11940 (N_11940,N_11699,N_11731);
nor U11941 (N_11941,N_11783,N_11684);
or U11942 (N_11942,N_11787,N_11740);
nand U11943 (N_11943,N_11739,N_11784);
nor U11944 (N_11944,N_11737,N_11699);
and U11945 (N_11945,N_11832,N_11690);
and U11946 (N_11946,N_11727,N_11716);
nor U11947 (N_11947,N_11701,N_11741);
xor U11948 (N_11948,N_11728,N_11755);
xnor U11949 (N_11949,N_11680,N_11813);
nor U11950 (N_11950,N_11818,N_11695);
or U11951 (N_11951,N_11812,N_11754);
nand U11952 (N_11952,N_11839,N_11706);
and U11953 (N_11953,N_11831,N_11688);
nand U11954 (N_11954,N_11729,N_11782);
nand U11955 (N_11955,N_11725,N_11766);
xor U11956 (N_11956,N_11741,N_11828);
or U11957 (N_11957,N_11705,N_11688);
nor U11958 (N_11958,N_11758,N_11743);
nand U11959 (N_11959,N_11720,N_11766);
and U11960 (N_11960,N_11755,N_11686);
nand U11961 (N_11961,N_11826,N_11707);
nand U11962 (N_11962,N_11779,N_11757);
or U11963 (N_11963,N_11724,N_11709);
nand U11964 (N_11964,N_11834,N_11786);
and U11965 (N_11965,N_11731,N_11746);
or U11966 (N_11966,N_11792,N_11683);
or U11967 (N_11967,N_11808,N_11805);
and U11968 (N_11968,N_11811,N_11743);
or U11969 (N_11969,N_11699,N_11828);
and U11970 (N_11970,N_11789,N_11733);
nor U11971 (N_11971,N_11682,N_11685);
xnor U11972 (N_11972,N_11771,N_11702);
or U11973 (N_11973,N_11771,N_11716);
nor U11974 (N_11974,N_11699,N_11709);
or U11975 (N_11975,N_11758,N_11682);
nor U11976 (N_11976,N_11756,N_11687);
nor U11977 (N_11977,N_11716,N_11820);
or U11978 (N_11978,N_11807,N_11710);
nor U11979 (N_11979,N_11771,N_11795);
or U11980 (N_11980,N_11692,N_11739);
or U11981 (N_11981,N_11780,N_11826);
xor U11982 (N_11982,N_11682,N_11733);
or U11983 (N_11983,N_11812,N_11803);
nand U11984 (N_11984,N_11758,N_11781);
or U11985 (N_11985,N_11831,N_11814);
nand U11986 (N_11986,N_11716,N_11699);
nand U11987 (N_11987,N_11767,N_11718);
nand U11988 (N_11988,N_11776,N_11816);
or U11989 (N_11989,N_11712,N_11795);
nor U11990 (N_11990,N_11719,N_11780);
or U11991 (N_11991,N_11774,N_11728);
xnor U11992 (N_11992,N_11804,N_11810);
and U11993 (N_11993,N_11798,N_11813);
nor U11994 (N_11994,N_11778,N_11742);
xnor U11995 (N_11995,N_11775,N_11736);
nor U11996 (N_11996,N_11803,N_11725);
nand U11997 (N_11997,N_11830,N_11733);
and U11998 (N_11998,N_11751,N_11762);
xnor U11999 (N_11999,N_11787,N_11692);
nor U12000 (N_12000,N_11992,N_11991);
nor U12001 (N_12001,N_11954,N_11841);
xor U12002 (N_12002,N_11950,N_11902);
and U12003 (N_12003,N_11868,N_11901);
and U12004 (N_12004,N_11871,N_11978);
nor U12005 (N_12005,N_11996,N_11908);
nand U12006 (N_12006,N_11988,N_11851);
xnor U12007 (N_12007,N_11937,N_11930);
nor U12008 (N_12008,N_11966,N_11926);
and U12009 (N_12009,N_11971,N_11927);
nand U12010 (N_12010,N_11845,N_11892);
nand U12011 (N_12011,N_11975,N_11893);
or U12012 (N_12012,N_11906,N_11934);
nand U12013 (N_12013,N_11920,N_11890);
and U12014 (N_12014,N_11874,N_11929);
nand U12015 (N_12015,N_11899,N_11863);
xor U12016 (N_12016,N_11942,N_11945);
nor U12017 (N_12017,N_11947,N_11907);
nor U12018 (N_12018,N_11867,N_11982);
nor U12019 (N_12019,N_11921,N_11858);
and U12020 (N_12020,N_11925,N_11849);
nand U12021 (N_12021,N_11919,N_11963);
nor U12022 (N_12022,N_11923,N_11913);
nor U12023 (N_12023,N_11957,N_11969);
nor U12024 (N_12024,N_11887,N_11897);
nor U12025 (N_12025,N_11968,N_11864);
xor U12026 (N_12026,N_11846,N_11854);
xor U12027 (N_12027,N_11914,N_11941);
nor U12028 (N_12028,N_11997,N_11967);
nor U12029 (N_12029,N_11974,N_11844);
nor U12030 (N_12030,N_11928,N_11904);
xnor U12031 (N_12031,N_11961,N_11884);
nand U12032 (N_12032,N_11980,N_11873);
xor U12033 (N_12033,N_11935,N_11903);
and U12034 (N_12034,N_11933,N_11883);
nor U12035 (N_12035,N_11865,N_11847);
and U12036 (N_12036,N_11960,N_11981);
or U12037 (N_12037,N_11886,N_11993);
nand U12038 (N_12038,N_11965,N_11924);
nor U12039 (N_12039,N_11877,N_11880);
and U12040 (N_12040,N_11972,N_11931);
nand U12041 (N_12041,N_11852,N_11912);
or U12042 (N_12042,N_11916,N_11885);
nor U12043 (N_12043,N_11848,N_11973);
nor U12044 (N_12044,N_11895,N_11918);
nor U12045 (N_12045,N_11987,N_11940);
or U12046 (N_12046,N_11939,N_11917);
and U12047 (N_12047,N_11900,N_11952);
xor U12048 (N_12048,N_11909,N_11976);
nor U12049 (N_12049,N_11956,N_11989);
nand U12050 (N_12050,N_11985,N_11882);
xnor U12051 (N_12051,N_11898,N_11958);
xnor U12052 (N_12052,N_11944,N_11911);
xnor U12053 (N_12053,N_11955,N_11995);
or U12054 (N_12054,N_11872,N_11959);
or U12055 (N_12055,N_11994,N_11861);
or U12056 (N_12056,N_11979,N_11905);
nor U12057 (N_12057,N_11855,N_11889);
nor U12058 (N_12058,N_11875,N_11922);
or U12059 (N_12059,N_11910,N_11843);
xnor U12060 (N_12060,N_11938,N_11842);
and U12061 (N_12061,N_11881,N_11857);
xnor U12062 (N_12062,N_11949,N_11953);
or U12063 (N_12063,N_11946,N_11856);
or U12064 (N_12064,N_11970,N_11870);
or U12065 (N_12065,N_11964,N_11999);
nor U12066 (N_12066,N_11951,N_11859);
or U12067 (N_12067,N_11986,N_11840);
and U12068 (N_12068,N_11850,N_11983);
or U12069 (N_12069,N_11896,N_11998);
or U12070 (N_12070,N_11891,N_11853);
nor U12071 (N_12071,N_11977,N_11984);
nand U12072 (N_12072,N_11932,N_11878);
xnor U12073 (N_12073,N_11915,N_11860);
nor U12074 (N_12074,N_11869,N_11894);
nor U12075 (N_12075,N_11962,N_11943);
nor U12076 (N_12076,N_11888,N_11866);
nor U12077 (N_12077,N_11876,N_11948);
or U12078 (N_12078,N_11862,N_11990);
and U12079 (N_12079,N_11879,N_11936);
or U12080 (N_12080,N_11856,N_11853);
xor U12081 (N_12081,N_11879,N_11954);
and U12082 (N_12082,N_11905,N_11909);
and U12083 (N_12083,N_11922,N_11913);
nor U12084 (N_12084,N_11951,N_11899);
nor U12085 (N_12085,N_11883,N_11904);
and U12086 (N_12086,N_11879,N_11850);
nor U12087 (N_12087,N_11874,N_11983);
nand U12088 (N_12088,N_11934,N_11901);
nor U12089 (N_12089,N_11897,N_11900);
nand U12090 (N_12090,N_11907,N_11923);
or U12091 (N_12091,N_11898,N_11896);
and U12092 (N_12092,N_11902,N_11995);
or U12093 (N_12093,N_11922,N_11884);
xnor U12094 (N_12094,N_11951,N_11954);
nor U12095 (N_12095,N_11999,N_11996);
nor U12096 (N_12096,N_11853,N_11889);
xor U12097 (N_12097,N_11958,N_11995);
nand U12098 (N_12098,N_11947,N_11948);
or U12099 (N_12099,N_11867,N_11921);
nor U12100 (N_12100,N_11892,N_11934);
nor U12101 (N_12101,N_11861,N_11936);
nor U12102 (N_12102,N_11983,N_11897);
or U12103 (N_12103,N_11936,N_11907);
nor U12104 (N_12104,N_11973,N_11850);
nand U12105 (N_12105,N_11897,N_11863);
or U12106 (N_12106,N_11845,N_11951);
nand U12107 (N_12107,N_11955,N_11942);
xnor U12108 (N_12108,N_11847,N_11945);
nor U12109 (N_12109,N_11890,N_11919);
xnor U12110 (N_12110,N_11912,N_11999);
nor U12111 (N_12111,N_11995,N_11873);
nand U12112 (N_12112,N_11862,N_11998);
nor U12113 (N_12113,N_11979,N_11904);
nor U12114 (N_12114,N_11952,N_11886);
xor U12115 (N_12115,N_11972,N_11980);
nor U12116 (N_12116,N_11982,N_11977);
and U12117 (N_12117,N_11907,N_11968);
and U12118 (N_12118,N_11976,N_11962);
xnor U12119 (N_12119,N_11986,N_11966);
or U12120 (N_12120,N_11910,N_11886);
nor U12121 (N_12121,N_11998,N_11876);
nor U12122 (N_12122,N_11993,N_11981);
nor U12123 (N_12123,N_11921,N_11998);
nand U12124 (N_12124,N_11874,N_11986);
or U12125 (N_12125,N_11911,N_11953);
nand U12126 (N_12126,N_11919,N_11920);
and U12127 (N_12127,N_11905,N_11879);
and U12128 (N_12128,N_11919,N_11908);
xor U12129 (N_12129,N_11904,N_11998);
nor U12130 (N_12130,N_11891,N_11930);
xor U12131 (N_12131,N_11937,N_11867);
or U12132 (N_12132,N_11905,N_11941);
nor U12133 (N_12133,N_11848,N_11922);
nor U12134 (N_12134,N_11979,N_11866);
xor U12135 (N_12135,N_11934,N_11897);
xor U12136 (N_12136,N_11984,N_11890);
nand U12137 (N_12137,N_11909,N_11927);
or U12138 (N_12138,N_11942,N_11856);
nand U12139 (N_12139,N_11953,N_11849);
nand U12140 (N_12140,N_11968,N_11985);
or U12141 (N_12141,N_11865,N_11980);
nor U12142 (N_12142,N_11947,N_11954);
nor U12143 (N_12143,N_11888,N_11903);
nand U12144 (N_12144,N_11901,N_11982);
nor U12145 (N_12145,N_11854,N_11881);
xor U12146 (N_12146,N_11928,N_11946);
xnor U12147 (N_12147,N_11998,N_11939);
nor U12148 (N_12148,N_11999,N_11872);
xnor U12149 (N_12149,N_11923,N_11924);
nand U12150 (N_12150,N_11887,N_11860);
nand U12151 (N_12151,N_11843,N_11867);
or U12152 (N_12152,N_11850,N_11887);
nor U12153 (N_12153,N_11879,N_11890);
xnor U12154 (N_12154,N_11999,N_11875);
nor U12155 (N_12155,N_11938,N_11920);
nor U12156 (N_12156,N_11939,N_11875);
xor U12157 (N_12157,N_11857,N_11871);
xor U12158 (N_12158,N_11936,N_11844);
nor U12159 (N_12159,N_11981,N_11916);
and U12160 (N_12160,N_12019,N_12082);
nand U12161 (N_12161,N_12097,N_12047);
and U12162 (N_12162,N_12098,N_12042);
xor U12163 (N_12163,N_12158,N_12037);
or U12164 (N_12164,N_12015,N_12014);
xnor U12165 (N_12165,N_12030,N_12106);
nand U12166 (N_12166,N_12068,N_12058);
and U12167 (N_12167,N_12117,N_12100);
or U12168 (N_12168,N_12149,N_12033);
nor U12169 (N_12169,N_12133,N_12079);
nand U12170 (N_12170,N_12006,N_12043);
and U12171 (N_12171,N_12074,N_12104);
and U12172 (N_12172,N_12076,N_12157);
or U12173 (N_12173,N_12084,N_12114);
nand U12174 (N_12174,N_12034,N_12110);
and U12175 (N_12175,N_12062,N_12108);
nand U12176 (N_12176,N_12025,N_12101);
nand U12177 (N_12177,N_12077,N_12010);
xnor U12178 (N_12178,N_12064,N_12136);
xor U12179 (N_12179,N_12009,N_12142);
nand U12180 (N_12180,N_12003,N_12138);
or U12181 (N_12181,N_12028,N_12128);
nand U12182 (N_12182,N_12150,N_12032);
and U12183 (N_12183,N_12054,N_12130);
and U12184 (N_12184,N_12039,N_12027);
nand U12185 (N_12185,N_12029,N_12125);
nor U12186 (N_12186,N_12159,N_12073);
and U12187 (N_12187,N_12078,N_12144);
and U12188 (N_12188,N_12135,N_12035);
xnor U12189 (N_12189,N_12066,N_12080);
and U12190 (N_12190,N_12123,N_12140);
nor U12191 (N_12191,N_12105,N_12118);
nand U12192 (N_12192,N_12056,N_12057);
xnor U12193 (N_12193,N_12093,N_12008);
and U12194 (N_12194,N_12070,N_12086);
or U12195 (N_12195,N_12132,N_12102);
xnor U12196 (N_12196,N_12038,N_12156);
or U12197 (N_12197,N_12022,N_12036);
xnor U12198 (N_12198,N_12088,N_12116);
and U12199 (N_12199,N_12099,N_12012);
and U12200 (N_12200,N_12134,N_12083);
xnor U12201 (N_12201,N_12063,N_12126);
xnor U12202 (N_12202,N_12155,N_12005);
nand U12203 (N_12203,N_12154,N_12148);
or U12204 (N_12204,N_12040,N_12115);
or U12205 (N_12205,N_12041,N_12020);
nand U12206 (N_12206,N_12146,N_12002);
nand U12207 (N_12207,N_12004,N_12051);
nor U12208 (N_12208,N_12026,N_12087);
xor U12209 (N_12209,N_12153,N_12075);
and U12210 (N_12210,N_12122,N_12145);
nor U12211 (N_12211,N_12061,N_12120);
nand U12212 (N_12212,N_12001,N_12007);
and U12213 (N_12213,N_12024,N_12092);
nand U12214 (N_12214,N_12072,N_12055);
and U12215 (N_12215,N_12143,N_12000);
or U12216 (N_12216,N_12141,N_12147);
xnor U12217 (N_12217,N_12018,N_12021);
nor U12218 (N_12218,N_12121,N_12113);
xnor U12219 (N_12219,N_12107,N_12045);
or U12220 (N_12220,N_12119,N_12053);
nand U12221 (N_12221,N_12112,N_12089);
nor U12222 (N_12222,N_12048,N_12052);
xor U12223 (N_12223,N_12049,N_12050);
nand U12224 (N_12224,N_12094,N_12111);
or U12225 (N_12225,N_12071,N_12059);
xor U12226 (N_12226,N_12085,N_12131);
xor U12227 (N_12227,N_12091,N_12046);
nand U12228 (N_12228,N_12109,N_12067);
xnor U12229 (N_12229,N_12031,N_12081);
and U12230 (N_12230,N_12069,N_12013);
or U12231 (N_12231,N_12017,N_12124);
xor U12232 (N_12232,N_12065,N_12152);
nor U12233 (N_12233,N_12151,N_12044);
xnor U12234 (N_12234,N_12016,N_12060);
or U12235 (N_12235,N_12137,N_12127);
and U12236 (N_12236,N_12023,N_12096);
xnor U12237 (N_12237,N_12129,N_12090);
and U12238 (N_12238,N_12095,N_12139);
and U12239 (N_12239,N_12011,N_12103);
nor U12240 (N_12240,N_12125,N_12041);
or U12241 (N_12241,N_12118,N_12043);
and U12242 (N_12242,N_12071,N_12103);
xor U12243 (N_12243,N_12095,N_12147);
or U12244 (N_12244,N_12071,N_12057);
nand U12245 (N_12245,N_12065,N_12146);
and U12246 (N_12246,N_12115,N_12004);
and U12247 (N_12247,N_12002,N_12091);
and U12248 (N_12248,N_12069,N_12029);
or U12249 (N_12249,N_12057,N_12112);
nand U12250 (N_12250,N_12001,N_12073);
or U12251 (N_12251,N_12102,N_12085);
nor U12252 (N_12252,N_12029,N_12122);
nand U12253 (N_12253,N_12091,N_12059);
and U12254 (N_12254,N_12054,N_12045);
xor U12255 (N_12255,N_12147,N_12115);
nor U12256 (N_12256,N_12071,N_12148);
xnor U12257 (N_12257,N_12059,N_12125);
nand U12258 (N_12258,N_12138,N_12058);
and U12259 (N_12259,N_12130,N_12028);
nor U12260 (N_12260,N_12079,N_12123);
xor U12261 (N_12261,N_12111,N_12058);
and U12262 (N_12262,N_12021,N_12022);
and U12263 (N_12263,N_12075,N_12032);
and U12264 (N_12264,N_12097,N_12002);
or U12265 (N_12265,N_12032,N_12040);
nand U12266 (N_12266,N_12096,N_12021);
or U12267 (N_12267,N_12066,N_12068);
xor U12268 (N_12268,N_12022,N_12032);
xor U12269 (N_12269,N_12135,N_12005);
nor U12270 (N_12270,N_12069,N_12116);
nor U12271 (N_12271,N_12023,N_12106);
nand U12272 (N_12272,N_12054,N_12016);
nand U12273 (N_12273,N_12029,N_12028);
or U12274 (N_12274,N_12158,N_12084);
nor U12275 (N_12275,N_12054,N_12089);
or U12276 (N_12276,N_12023,N_12159);
and U12277 (N_12277,N_12005,N_12069);
nand U12278 (N_12278,N_12018,N_12146);
nor U12279 (N_12279,N_12013,N_12040);
nor U12280 (N_12280,N_12040,N_12026);
nand U12281 (N_12281,N_12010,N_12122);
nor U12282 (N_12282,N_12101,N_12073);
and U12283 (N_12283,N_12056,N_12045);
nor U12284 (N_12284,N_12133,N_12140);
or U12285 (N_12285,N_12110,N_12138);
nor U12286 (N_12286,N_12082,N_12087);
xnor U12287 (N_12287,N_12083,N_12139);
nor U12288 (N_12288,N_12117,N_12017);
xnor U12289 (N_12289,N_12097,N_12034);
nand U12290 (N_12290,N_12089,N_12061);
xnor U12291 (N_12291,N_12148,N_12144);
and U12292 (N_12292,N_12156,N_12042);
nor U12293 (N_12293,N_12154,N_12037);
nor U12294 (N_12294,N_12116,N_12025);
and U12295 (N_12295,N_12006,N_12137);
and U12296 (N_12296,N_12124,N_12086);
or U12297 (N_12297,N_12078,N_12053);
nor U12298 (N_12298,N_12106,N_12152);
and U12299 (N_12299,N_12011,N_12000);
nand U12300 (N_12300,N_12087,N_12074);
and U12301 (N_12301,N_12115,N_12022);
xnor U12302 (N_12302,N_12149,N_12089);
xnor U12303 (N_12303,N_12137,N_12100);
or U12304 (N_12304,N_12077,N_12155);
nor U12305 (N_12305,N_12138,N_12145);
nor U12306 (N_12306,N_12105,N_12108);
and U12307 (N_12307,N_12158,N_12048);
and U12308 (N_12308,N_12106,N_12084);
and U12309 (N_12309,N_12100,N_12065);
or U12310 (N_12310,N_12117,N_12126);
nor U12311 (N_12311,N_12045,N_12092);
or U12312 (N_12312,N_12017,N_12093);
nand U12313 (N_12313,N_12067,N_12153);
nand U12314 (N_12314,N_12053,N_12147);
and U12315 (N_12315,N_12152,N_12028);
and U12316 (N_12316,N_12080,N_12052);
and U12317 (N_12317,N_12006,N_12076);
and U12318 (N_12318,N_12017,N_12076);
and U12319 (N_12319,N_12016,N_12070);
or U12320 (N_12320,N_12313,N_12211);
xor U12321 (N_12321,N_12256,N_12178);
nor U12322 (N_12322,N_12215,N_12306);
and U12323 (N_12323,N_12309,N_12168);
nor U12324 (N_12324,N_12225,N_12281);
or U12325 (N_12325,N_12175,N_12301);
and U12326 (N_12326,N_12199,N_12210);
and U12327 (N_12327,N_12254,N_12241);
and U12328 (N_12328,N_12314,N_12277);
or U12329 (N_12329,N_12180,N_12316);
or U12330 (N_12330,N_12247,N_12213);
nand U12331 (N_12331,N_12317,N_12297);
or U12332 (N_12332,N_12166,N_12228);
and U12333 (N_12333,N_12204,N_12183);
and U12334 (N_12334,N_12266,N_12289);
xor U12335 (N_12335,N_12226,N_12276);
nand U12336 (N_12336,N_12182,N_12235);
nor U12337 (N_12337,N_12236,N_12299);
or U12338 (N_12338,N_12305,N_12270);
and U12339 (N_12339,N_12217,N_12304);
or U12340 (N_12340,N_12188,N_12205);
xnor U12341 (N_12341,N_12238,N_12307);
nand U12342 (N_12342,N_12315,N_12233);
nand U12343 (N_12343,N_12222,N_12163);
and U12344 (N_12344,N_12230,N_12174);
and U12345 (N_12345,N_12169,N_12192);
xor U12346 (N_12346,N_12190,N_12224);
xnor U12347 (N_12347,N_12196,N_12223);
nor U12348 (N_12348,N_12308,N_12203);
and U12349 (N_12349,N_12264,N_12179);
nor U12350 (N_12350,N_12319,N_12285);
nand U12351 (N_12351,N_12227,N_12165);
nand U12352 (N_12352,N_12300,N_12257);
nand U12353 (N_12353,N_12310,N_12259);
nand U12354 (N_12354,N_12283,N_12253);
nor U12355 (N_12355,N_12292,N_12272);
nor U12356 (N_12356,N_12251,N_12275);
and U12357 (N_12357,N_12239,N_12186);
nand U12358 (N_12358,N_12209,N_12207);
xnor U12359 (N_12359,N_12185,N_12262);
or U12360 (N_12360,N_12258,N_12260);
and U12361 (N_12361,N_12242,N_12263);
and U12362 (N_12362,N_12231,N_12291);
or U12363 (N_12363,N_12206,N_12274);
nor U12364 (N_12364,N_12212,N_12279);
and U12365 (N_12365,N_12261,N_12244);
nand U12366 (N_12366,N_12245,N_12191);
or U12367 (N_12367,N_12255,N_12278);
xor U12368 (N_12368,N_12184,N_12271);
nand U12369 (N_12369,N_12214,N_12193);
nand U12370 (N_12370,N_12312,N_12219);
and U12371 (N_12371,N_12252,N_12160);
nand U12372 (N_12372,N_12218,N_12216);
xor U12373 (N_12373,N_12220,N_12290);
nand U12374 (N_12374,N_12197,N_12200);
nand U12375 (N_12375,N_12161,N_12298);
nor U12376 (N_12376,N_12237,N_12173);
nor U12377 (N_12377,N_12208,N_12195);
nand U12378 (N_12378,N_12229,N_12273);
or U12379 (N_12379,N_12243,N_12311);
nand U12380 (N_12380,N_12202,N_12286);
nor U12381 (N_12381,N_12201,N_12246);
nand U12382 (N_12382,N_12287,N_12198);
nor U12383 (N_12383,N_12234,N_12294);
and U12384 (N_12384,N_12296,N_12181);
nor U12385 (N_12385,N_12267,N_12284);
or U12386 (N_12386,N_12240,N_12302);
nor U12387 (N_12387,N_12176,N_12248);
and U12388 (N_12388,N_12268,N_12250);
and U12389 (N_12389,N_12318,N_12232);
nand U12390 (N_12390,N_12171,N_12288);
or U12391 (N_12391,N_12221,N_12269);
nor U12392 (N_12392,N_12164,N_12293);
and U12393 (N_12393,N_12167,N_12280);
nor U12394 (N_12394,N_12282,N_12303);
nand U12395 (N_12395,N_12162,N_12295);
and U12396 (N_12396,N_12249,N_12170);
xor U12397 (N_12397,N_12177,N_12187);
nand U12398 (N_12398,N_12194,N_12189);
nand U12399 (N_12399,N_12172,N_12265);
nor U12400 (N_12400,N_12247,N_12303);
and U12401 (N_12401,N_12291,N_12290);
nand U12402 (N_12402,N_12253,N_12201);
nor U12403 (N_12403,N_12271,N_12197);
nor U12404 (N_12404,N_12290,N_12266);
and U12405 (N_12405,N_12243,N_12266);
or U12406 (N_12406,N_12296,N_12309);
xnor U12407 (N_12407,N_12267,N_12176);
nor U12408 (N_12408,N_12218,N_12313);
and U12409 (N_12409,N_12200,N_12262);
xnor U12410 (N_12410,N_12170,N_12216);
and U12411 (N_12411,N_12162,N_12251);
nand U12412 (N_12412,N_12268,N_12215);
xnor U12413 (N_12413,N_12246,N_12282);
or U12414 (N_12414,N_12250,N_12225);
nor U12415 (N_12415,N_12308,N_12178);
and U12416 (N_12416,N_12255,N_12234);
nor U12417 (N_12417,N_12168,N_12273);
or U12418 (N_12418,N_12226,N_12230);
xor U12419 (N_12419,N_12210,N_12200);
xnor U12420 (N_12420,N_12245,N_12230);
xor U12421 (N_12421,N_12305,N_12218);
or U12422 (N_12422,N_12318,N_12248);
nor U12423 (N_12423,N_12315,N_12236);
nor U12424 (N_12424,N_12206,N_12254);
nand U12425 (N_12425,N_12310,N_12289);
xor U12426 (N_12426,N_12162,N_12317);
nand U12427 (N_12427,N_12309,N_12201);
xnor U12428 (N_12428,N_12296,N_12165);
nor U12429 (N_12429,N_12296,N_12286);
or U12430 (N_12430,N_12230,N_12235);
or U12431 (N_12431,N_12293,N_12176);
and U12432 (N_12432,N_12202,N_12232);
or U12433 (N_12433,N_12314,N_12200);
and U12434 (N_12434,N_12232,N_12297);
nand U12435 (N_12435,N_12302,N_12195);
nand U12436 (N_12436,N_12189,N_12315);
and U12437 (N_12437,N_12314,N_12170);
xor U12438 (N_12438,N_12270,N_12314);
nand U12439 (N_12439,N_12312,N_12166);
xor U12440 (N_12440,N_12271,N_12206);
or U12441 (N_12441,N_12192,N_12295);
nand U12442 (N_12442,N_12289,N_12177);
nor U12443 (N_12443,N_12279,N_12256);
nand U12444 (N_12444,N_12199,N_12295);
xnor U12445 (N_12445,N_12165,N_12313);
or U12446 (N_12446,N_12209,N_12275);
or U12447 (N_12447,N_12317,N_12199);
xor U12448 (N_12448,N_12223,N_12276);
and U12449 (N_12449,N_12211,N_12267);
nor U12450 (N_12450,N_12218,N_12165);
nor U12451 (N_12451,N_12183,N_12282);
xor U12452 (N_12452,N_12162,N_12254);
nor U12453 (N_12453,N_12244,N_12262);
xor U12454 (N_12454,N_12300,N_12301);
or U12455 (N_12455,N_12225,N_12160);
or U12456 (N_12456,N_12211,N_12212);
or U12457 (N_12457,N_12186,N_12222);
and U12458 (N_12458,N_12201,N_12162);
nand U12459 (N_12459,N_12314,N_12219);
and U12460 (N_12460,N_12189,N_12253);
xnor U12461 (N_12461,N_12291,N_12173);
nand U12462 (N_12462,N_12242,N_12266);
xnor U12463 (N_12463,N_12169,N_12283);
nor U12464 (N_12464,N_12282,N_12176);
or U12465 (N_12465,N_12309,N_12173);
or U12466 (N_12466,N_12223,N_12269);
xnor U12467 (N_12467,N_12243,N_12283);
xnor U12468 (N_12468,N_12236,N_12256);
xor U12469 (N_12469,N_12243,N_12265);
nor U12470 (N_12470,N_12183,N_12309);
nor U12471 (N_12471,N_12204,N_12193);
xor U12472 (N_12472,N_12266,N_12312);
nor U12473 (N_12473,N_12314,N_12208);
nand U12474 (N_12474,N_12225,N_12167);
nor U12475 (N_12475,N_12318,N_12167);
nor U12476 (N_12476,N_12180,N_12169);
or U12477 (N_12477,N_12268,N_12211);
nor U12478 (N_12478,N_12297,N_12262);
nor U12479 (N_12479,N_12246,N_12264);
or U12480 (N_12480,N_12331,N_12332);
xnor U12481 (N_12481,N_12432,N_12392);
or U12482 (N_12482,N_12391,N_12400);
nor U12483 (N_12483,N_12465,N_12404);
or U12484 (N_12484,N_12342,N_12455);
nor U12485 (N_12485,N_12386,N_12335);
nor U12486 (N_12486,N_12390,N_12394);
or U12487 (N_12487,N_12358,N_12377);
nand U12488 (N_12488,N_12410,N_12351);
nand U12489 (N_12489,N_12417,N_12461);
and U12490 (N_12490,N_12324,N_12396);
xor U12491 (N_12491,N_12424,N_12321);
and U12492 (N_12492,N_12338,N_12353);
or U12493 (N_12493,N_12464,N_12365);
nor U12494 (N_12494,N_12339,N_12333);
or U12495 (N_12495,N_12340,N_12395);
nor U12496 (N_12496,N_12433,N_12468);
nor U12497 (N_12497,N_12453,N_12393);
nor U12498 (N_12498,N_12344,N_12388);
or U12499 (N_12499,N_12323,N_12382);
and U12500 (N_12500,N_12438,N_12422);
nor U12501 (N_12501,N_12470,N_12457);
xnor U12502 (N_12502,N_12439,N_12372);
nor U12503 (N_12503,N_12431,N_12429);
and U12504 (N_12504,N_12381,N_12373);
nand U12505 (N_12505,N_12423,N_12345);
nand U12506 (N_12506,N_12436,N_12375);
nor U12507 (N_12507,N_12399,N_12369);
nor U12508 (N_12508,N_12419,N_12456);
xnor U12509 (N_12509,N_12346,N_12374);
nor U12510 (N_12510,N_12452,N_12364);
xnor U12511 (N_12511,N_12467,N_12343);
nor U12512 (N_12512,N_12367,N_12387);
or U12513 (N_12513,N_12444,N_12446);
nor U12514 (N_12514,N_12376,N_12421);
xnor U12515 (N_12515,N_12347,N_12384);
and U12516 (N_12516,N_12472,N_12334);
and U12517 (N_12517,N_12462,N_12426);
nand U12518 (N_12518,N_12360,N_12428);
nand U12519 (N_12519,N_12475,N_12418);
xnor U12520 (N_12520,N_12326,N_12328);
or U12521 (N_12521,N_12409,N_12448);
xor U12522 (N_12522,N_12469,N_12460);
xor U12523 (N_12523,N_12327,N_12477);
xor U12524 (N_12524,N_12336,N_12407);
nand U12525 (N_12525,N_12320,N_12449);
nor U12526 (N_12526,N_12348,N_12463);
or U12527 (N_12527,N_12385,N_12451);
nor U12528 (N_12528,N_12389,N_12441);
and U12529 (N_12529,N_12479,N_12378);
nor U12530 (N_12530,N_12383,N_12406);
or U12531 (N_12531,N_12450,N_12362);
nor U12532 (N_12532,N_12329,N_12380);
nand U12533 (N_12533,N_12445,N_12471);
nor U12534 (N_12534,N_12434,N_12357);
and U12535 (N_12535,N_12454,N_12459);
xnor U12536 (N_12536,N_12440,N_12371);
xor U12537 (N_12537,N_12361,N_12330);
nand U12538 (N_12538,N_12435,N_12447);
nor U12539 (N_12539,N_12416,N_12478);
or U12540 (N_12540,N_12354,N_12366);
or U12541 (N_12541,N_12322,N_12368);
nand U12542 (N_12542,N_12474,N_12341);
and U12543 (N_12543,N_12349,N_12398);
xor U12544 (N_12544,N_12427,N_12437);
and U12545 (N_12545,N_12408,N_12397);
nor U12546 (N_12546,N_12405,N_12413);
nand U12547 (N_12547,N_12420,N_12379);
xnor U12548 (N_12548,N_12425,N_12352);
nor U12549 (N_12549,N_12355,N_12403);
and U12550 (N_12550,N_12466,N_12359);
nand U12551 (N_12551,N_12442,N_12430);
nand U12552 (N_12552,N_12401,N_12476);
nand U12553 (N_12553,N_12356,N_12325);
xor U12554 (N_12554,N_12337,N_12414);
xnor U12555 (N_12555,N_12411,N_12370);
or U12556 (N_12556,N_12412,N_12443);
nand U12557 (N_12557,N_12363,N_12350);
nand U12558 (N_12558,N_12458,N_12415);
nor U12559 (N_12559,N_12402,N_12473);
or U12560 (N_12560,N_12442,N_12395);
nand U12561 (N_12561,N_12328,N_12454);
nand U12562 (N_12562,N_12340,N_12456);
nor U12563 (N_12563,N_12453,N_12479);
nor U12564 (N_12564,N_12361,N_12402);
and U12565 (N_12565,N_12461,N_12436);
or U12566 (N_12566,N_12378,N_12392);
or U12567 (N_12567,N_12436,N_12380);
or U12568 (N_12568,N_12391,N_12466);
xor U12569 (N_12569,N_12444,N_12371);
or U12570 (N_12570,N_12415,N_12457);
or U12571 (N_12571,N_12414,N_12411);
xor U12572 (N_12572,N_12454,N_12412);
xnor U12573 (N_12573,N_12426,N_12444);
nor U12574 (N_12574,N_12386,N_12461);
nor U12575 (N_12575,N_12449,N_12357);
and U12576 (N_12576,N_12370,N_12409);
and U12577 (N_12577,N_12428,N_12326);
xnor U12578 (N_12578,N_12366,N_12455);
nand U12579 (N_12579,N_12328,N_12334);
nor U12580 (N_12580,N_12376,N_12467);
or U12581 (N_12581,N_12440,N_12357);
nand U12582 (N_12582,N_12436,N_12425);
xor U12583 (N_12583,N_12419,N_12352);
nor U12584 (N_12584,N_12403,N_12397);
nor U12585 (N_12585,N_12386,N_12410);
nand U12586 (N_12586,N_12351,N_12399);
nor U12587 (N_12587,N_12343,N_12465);
or U12588 (N_12588,N_12343,N_12393);
xor U12589 (N_12589,N_12423,N_12331);
nand U12590 (N_12590,N_12432,N_12346);
xnor U12591 (N_12591,N_12332,N_12445);
or U12592 (N_12592,N_12455,N_12368);
or U12593 (N_12593,N_12331,N_12431);
and U12594 (N_12594,N_12343,N_12402);
nand U12595 (N_12595,N_12475,N_12463);
nand U12596 (N_12596,N_12425,N_12370);
nor U12597 (N_12597,N_12351,N_12381);
nor U12598 (N_12598,N_12329,N_12337);
xor U12599 (N_12599,N_12374,N_12385);
xor U12600 (N_12600,N_12451,N_12395);
nor U12601 (N_12601,N_12470,N_12326);
nor U12602 (N_12602,N_12438,N_12386);
nor U12603 (N_12603,N_12396,N_12401);
or U12604 (N_12604,N_12423,N_12454);
nand U12605 (N_12605,N_12408,N_12432);
or U12606 (N_12606,N_12425,N_12415);
xor U12607 (N_12607,N_12388,N_12457);
nor U12608 (N_12608,N_12338,N_12442);
nor U12609 (N_12609,N_12392,N_12472);
xnor U12610 (N_12610,N_12329,N_12421);
nand U12611 (N_12611,N_12468,N_12414);
and U12612 (N_12612,N_12478,N_12434);
nand U12613 (N_12613,N_12337,N_12429);
xor U12614 (N_12614,N_12389,N_12447);
nor U12615 (N_12615,N_12457,N_12421);
nand U12616 (N_12616,N_12441,N_12417);
nand U12617 (N_12617,N_12388,N_12347);
nor U12618 (N_12618,N_12356,N_12338);
and U12619 (N_12619,N_12456,N_12438);
and U12620 (N_12620,N_12327,N_12440);
xor U12621 (N_12621,N_12420,N_12460);
xor U12622 (N_12622,N_12443,N_12342);
xnor U12623 (N_12623,N_12412,N_12476);
nor U12624 (N_12624,N_12344,N_12347);
nand U12625 (N_12625,N_12350,N_12366);
nor U12626 (N_12626,N_12373,N_12352);
nor U12627 (N_12627,N_12359,N_12377);
xor U12628 (N_12628,N_12389,N_12360);
xnor U12629 (N_12629,N_12331,N_12479);
and U12630 (N_12630,N_12353,N_12379);
nand U12631 (N_12631,N_12475,N_12343);
or U12632 (N_12632,N_12455,N_12452);
nand U12633 (N_12633,N_12341,N_12418);
and U12634 (N_12634,N_12449,N_12348);
nand U12635 (N_12635,N_12454,N_12455);
xnor U12636 (N_12636,N_12403,N_12440);
xor U12637 (N_12637,N_12466,N_12369);
nor U12638 (N_12638,N_12435,N_12472);
nor U12639 (N_12639,N_12396,N_12344);
or U12640 (N_12640,N_12510,N_12501);
nor U12641 (N_12641,N_12592,N_12588);
nor U12642 (N_12642,N_12576,N_12532);
xor U12643 (N_12643,N_12531,N_12520);
or U12644 (N_12644,N_12546,N_12529);
nand U12645 (N_12645,N_12533,N_12563);
and U12646 (N_12646,N_12509,N_12575);
and U12647 (N_12647,N_12613,N_12630);
xnor U12648 (N_12648,N_12595,N_12511);
nor U12649 (N_12649,N_12550,N_12622);
or U12650 (N_12650,N_12549,N_12556);
nor U12651 (N_12651,N_12525,N_12499);
nand U12652 (N_12652,N_12616,N_12602);
nor U12653 (N_12653,N_12502,N_12605);
or U12654 (N_12654,N_12587,N_12559);
xor U12655 (N_12655,N_12580,N_12585);
xor U12656 (N_12656,N_12577,N_12600);
and U12657 (N_12657,N_12541,N_12631);
nand U12658 (N_12658,N_12625,N_12581);
or U12659 (N_12659,N_12483,N_12582);
and U12660 (N_12660,N_12621,N_12522);
and U12661 (N_12661,N_12539,N_12589);
nor U12662 (N_12662,N_12615,N_12491);
nand U12663 (N_12663,N_12552,N_12528);
xnor U12664 (N_12664,N_12495,N_12494);
or U12665 (N_12665,N_12612,N_12599);
and U12666 (N_12666,N_12598,N_12524);
or U12667 (N_12667,N_12526,N_12562);
xnor U12668 (N_12668,N_12516,N_12623);
and U12669 (N_12669,N_12540,N_12637);
and U12670 (N_12670,N_12633,N_12572);
nand U12671 (N_12671,N_12536,N_12503);
xor U12672 (N_12672,N_12597,N_12497);
nor U12673 (N_12673,N_12565,N_12610);
nor U12674 (N_12674,N_12618,N_12512);
and U12675 (N_12675,N_12578,N_12542);
nand U12676 (N_12676,N_12574,N_12628);
and U12677 (N_12677,N_12561,N_12627);
or U12678 (N_12678,N_12617,N_12603);
nor U12679 (N_12679,N_12496,N_12568);
xor U12680 (N_12680,N_12514,N_12564);
and U12681 (N_12681,N_12485,N_12634);
nand U12682 (N_12682,N_12596,N_12490);
nor U12683 (N_12683,N_12566,N_12569);
xor U12684 (N_12684,N_12489,N_12493);
nand U12685 (N_12685,N_12557,N_12498);
and U12686 (N_12686,N_12535,N_12638);
and U12687 (N_12687,N_12484,N_12636);
or U12688 (N_12688,N_12593,N_12586);
xnor U12689 (N_12689,N_12551,N_12591);
or U12690 (N_12690,N_12530,N_12521);
or U12691 (N_12691,N_12570,N_12500);
and U12692 (N_12692,N_12583,N_12547);
and U12693 (N_12693,N_12573,N_12534);
nor U12694 (N_12694,N_12619,N_12620);
or U12695 (N_12695,N_12555,N_12567);
nand U12696 (N_12696,N_12604,N_12505);
and U12697 (N_12697,N_12584,N_12554);
nor U12698 (N_12698,N_12639,N_12518);
nand U12699 (N_12699,N_12594,N_12519);
xor U12700 (N_12700,N_12527,N_12508);
or U12701 (N_12701,N_12506,N_12629);
nand U12702 (N_12702,N_12548,N_12611);
xor U12703 (N_12703,N_12553,N_12481);
nand U12704 (N_12704,N_12515,N_12608);
or U12705 (N_12705,N_12624,N_12487);
and U12706 (N_12706,N_12545,N_12537);
and U12707 (N_12707,N_12614,N_12544);
or U12708 (N_12708,N_12626,N_12517);
nor U12709 (N_12709,N_12606,N_12523);
or U12710 (N_12710,N_12558,N_12601);
nand U12711 (N_12711,N_12609,N_12635);
xnor U12712 (N_12712,N_12632,N_12482);
nor U12713 (N_12713,N_12488,N_12513);
or U12714 (N_12714,N_12543,N_12579);
xnor U12715 (N_12715,N_12571,N_12486);
nand U12716 (N_12716,N_12507,N_12560);
xor U12717 (N_12717,N_12607,N_12492);
nor U12718 (N_12718,N_12504,N_12480);
and U12719 (N_12719,N_12538,N_12590);
nor U12720 (N_12720,N_12557,N_12501);
nand U12721 (N_12721,N_12606,N_12569);
and U12722 (N_12722,N_12522,N_12488);
and U12723 (N_12723,N_12496,N_12574);
xnor U12724 (N_12724,N_12580,N_12630);
or U12725 (N_12725,N_12510,N_12500);
or U12726 (N_12726,N_12606,N_12583);
nand U12727 (N_12727,N_12552,N_12510);
nor U12728 (N_12728,N_12513,N_12615);
nand U12729 (N_12729,N_12551,N_12603);
nand U12730 (N_12730,N_12631,N_12555);
and U12731 (N_12731,N_12569,N_12577);
nor U12732 (N_12732,N_12596,N_12557);
and U12733 (N_12733,N_12570,N_12528);
nor U12734 (N_12734,N_12586,N_12507);
nand U12735 (N_12735,N_12544,N_12492);
nor U12736 (N_12736,N_12566,N_12602);
and U12737 (N_12737,N_12629,N_12584);
or U12738 (N_12738,N_12608,N_12509);
nand U12739 (N_12739,N_12485,N_12621);
xor U12740 (N_12740,N_12515,N_12618);
or U12741 (N_12741,N_12486,N_12496);
xor U12742 (N_12742,N_12574,N_12549);
nand U12743 (N_12743,N_12527,N_12544);
xnor U12744 (N_12744,N_12613,N_12592);
and U12745 (N_12745,N_12551,N_12546);
xor U12746 (N_12746,N_12511,N_12529);
xor U12747 (N_12747,N_12638,N_12624);
and U12748 (N_12748,N_12546,N_12505);
nand U12749 (N_12749,N_12557,N_12527);
nand U12750 (N_12750,N_12534,N_12582);
or U12751 (N_12751,N_12590,N_12634);
xor U12752 (N_12752,N_12588,N_12623);
nor U12753 (N_12753,N_12609,N_12517);
nor U12754 (N_12754,N_12526,N_12573);
and U12755 (N_12755,N_12516,N_12506);
nor U12756 (N_12756,N_12481,N_12531);
and U12757 (N_12757,N_12620,N_12508);
and U12758 (N_12758,N_12557,N_12537);
or U12759 (N_12759,N_12602,N_12543);
nand U12760 (N_12760,N_12493,N_12637);
nand U12761 (N_12761,N_12497,N_12569);
or U12762 (N_12762,N_12619,N_12487);
and U12763 (N_12763,N_12544,N_12557);
or U12764 (N_12764,N_12495,N_12574);
and U12765 (N_12765,N_12541,N_12505);
and U12766 (N_12766,N_12510,N_12605);
nor U12767 (N_12767,N_12577,N_12505);
and U12768 (N_12768,N_12493,N_12600);
nor U12769 (N_12769,N_12544,N_12589);
and U12770 (N_12770,N_12537,N_12632);
nand U12771 (N_12771,N_12480,N_12610);
or U12772 (N_12772,N_12578,N_12504);
nand U12773 (N_12773,N_12495,N_12560);
and U12774 (N_12774,N_12508,N_12553);
and U12775 (N_12775,N_12592,N_12597);
nor U12776 (N_12776,N_12545,N_12563);
nor U12777 (N_12777,N_12568,N_12556);
xnor U12778 (N_12778,N_12561,N_12527);
nor U12779 (N_12779,N_12488,N_12483);
nor U12780 (N_12780,N_12552,N_12586);
nor U12781 (N_12781,N_12611,N_12617);
nor U12782 (N_12782,N_12549,N_12484);
nor U12783 (N_12783,N_12516,N_12619);
nor U12784 (N_12784,N_12537,N_12578);
or U12785 (N_12785,N_12524,N_12542);
xnor U12786 (N_12786,N_12595,N_12509);
nand U12787 (N_12787,N_12611,N_12551);
xor U12788 (N_12788,N_12610,N_12512);
nor U12789 (N_12789,N_12585,N_12556);
nand U12790 (N_12790,N_12524,N_12494);
and U12791 (N_12791,N_12572,N_12549);
nor U12792 (N_12792,N_12542,N_12500);
xor U12793 (N_12793,N_12634,N_12504);
nand U12794 (N_12794,N_12580,N_12595);
nor U12795 (N_12795,N_12480,N_12564);
nor U12796 (N_12796,N_12551,N_12526);
and U12797 (N_12797,N_12554,N_12588);
and U12798 (N_12798,N_12539,N_12489);
or U12799 (N_12799,N_12542,N_12519);
xor U12800 (N_12800,N_12733,N_12669);
xor U12801 (N_12801,N_12747,N_12701);
nand U12802 (N_12802,N_12770,N_12736);
and U12803 (N_12803,N_12744,N_12727);
nor U12804 (N_12804,N_12791,N_12779);
xor U12805 (N_12805,N_12680,N_12725);
and U12806 (N_12806,N_12690,N_12702);
and U12807 (N_12807,N_12674,N_12652);
and U12808 (N_12808,N_12728,N_12651);
xnor U12809 (N_12809,N_12754,N_12792);
or U12810 (N_12810,N_12718,N_12668);
or U12811 (N_12811,N_12685,N_12769);
xnor U12812 (N_12812,N_12712,N_12784);
xor U12813 (N_12813,N_12675,N_12755);
or U12814 (N_12814,N_12714,N_12665);
xnor U12815 (N_12815,N_12798,N_12778);
and U12816 (N_12816,N_12726,N_12721);
and U12817 (N_12817,N_12793,N_12739);
or U12818 (N_12818,N_12737,N_12764);
nor U12819 (N_12819,N_12722,N_12772);
or U12820 (N_12820,N_12710,N_12765);
and U12821 (N_12821,N_12677,N_12662);
and U12822 (N_12822,N_12758,N_12750);
nand U12823 (N_12823,N_12654,N_12716);
nand U12824 (N_12824,N_12648,N_12761);
and U12825 (N_12825,N_12693,N_12655);
nor U12826 (N_12826,N_12653,N_12708);
or U12827 (N_12827,N_12647,N_12796);
nand U12828 (N_12828,N_12723,N_12717);
and U12829 (N_12829,N_12672,N_12641);
and U12830 (N_12830,N_12724,N_12650);
nand U12831 (N_12831,N_12745,N_12797);
or U12832 (N_12832,N_12679,N_12751);
or U12833 (N_12833,N_12698,N_12775);
xnor U12834 (N_12834,N_12704,N_12731);
nand U12835 (N_12835,N_12776,N_12743);
or U12836 (N_12836,N_12777,N_12729);
and U12837 (N_12837,N_12683,N_12794);
nand U12838 (N_12838,N_12645,N_12760);
xnor U12839 (N_12839,N_12782,N_12697);
nor U12840 (N_12840,N_12780,N_12789);
and U12841 (N_12841,N_12735,N_12766);
nand U12842 (N_12842,N_12676,N_12678);
and U12843 (N_12843,N_12783,N_12719);
nand U12844 (N_12844,N_12681,N_12699);
nor U12845 (N_12845,N_12670,N_12700);
and U12846 (N_12846,N_12642,N_12643);
nor U12847 (N_12847,N_12746,N_12711);
or U12848 (N_12848,N_12713,N_12742);
or U12849 (N_12849,N_12757,N_12646);
or U12850 (N_12850,N_12686,N_12738);
or U12851 (N_12851,N_12691,N_12640);
or U12852 (N_12852,N_12740,N_12656);
xor U12853 (N_12853,N_12694,N_12663);
and U12854 (N_12854,N_12785,N_12790);
xor U12855 (N_12855,N_12688,N_12787);
and U12856 (N_12856,N_12660,N_12734);
xor U12857 (N_12857,N_12795,N_12666);
xnor U12858 (N_12858,N_12774,N_12671);
xnor U12859 (N_12859,N_12799,N_12781);
xnor U12860 (N_12860,N_12657,N_12659);
xor U12861 (N_12861,N_12732,N_12673);
and U12862 (N_12862,N_12773,N_12759);
or U12863 (N_12863,N_12649,N_12664);
xor U12864 (N_12864,N_12771,N_12752);
and U12865 (N_12865,N_12705,N_12788);
or U12866 (N_12866,N_12644,N_12741);
nor U12867 (N_12867,N_12753,N_12762);
nand U12868 (N_12868,N_12749,N_12709);
nor U12869 (N_12869,N_12658,N_12763);
and U12870 (N_12870,N_12703,N_12682);
xor U12871 (N_12871,N_12695,N_12768);
xor U12872 (N_12872,N_12715,N_12689);
nand U12873 (N_12873,N_12720,N_12786);
and U12874 (N_12874,N_12707,N_12748);
nor U12875 (N_12875,N_12730,N_12684);
nand U12876 (N_12876,N_12767,N_12661);
nand U12877 (N_12877,N_12756,N_12706);
nand U12878 (N_12878,N_12696,N_12687);
xor U12879 (N_12879,N_12692,N_12667);
and U12880 (N_12880,N_12753,N_12665);
and U12881 (N_12881,N_12768,N_12715);
nand U12882 (N_12882,N_12667,N_12703);
or U12883 (N_12883,N_12688,N_12705);
nor U12884 (N_12884,N_12744,N_12662);
nor U12885 (N_12885,N_12684,N_12707);
xor U12886 (N_12886,N_12713,N_12725);
nor U12887 (N_12887,N_12642,N_12706);
and U12888 (N_12888,N_12666,N_12772);
nand U12889 (N_12889,N_12652,N_12732);
nor U12890 (N_12890,N_12763,N_12789);
nand U12891 (N_12891,N_12656,N_12780);
nand U12892 (N_12892,N_12722,N_12655);
or U12893 (N_12893,N_12690,N_12772);
nand U12894 (N_12894,N_12768,N_12781);
and U12895 (N_12895,N_12781,N_12749);
or U12896 (N_12896,N_12774,N_12700);
and U12897 (N_12897,N_12785,N_12701);
and U12898 (N_12898,N_12734,N_12647);
and U12899 (N_12899,N_12654,N_12669);
nor U12900 (N_12900,N_12663,N_12793);
or U12901 (N_12901,N_12763,N_12677);
nor U12902 (N_12902,N_12729,N_12660);
xnor U12903 (N_12903,N_12764,N_12776);
and U12904 (N_12904,N_12676,N_12739);
nand U12905 (N_12905,N_12772,N_12787);
and U12906 (N_12906,N_12668,N_12682);
and U12907 (N_12907,N_12704,N_12711);
nor U12908 (N_12908,N_12740,N_12799);
and U12909 (N_12909,N_12725,N_12705);
nor U12910 (N_12910,N_12654,N_12718);
and U12911 (N_12911,N_12640,N_12749);
xnor U12912 (N_12912,N_12792,N_12646);
xnor U12913 (N_12913,N_12675,N_12749);
or U12914 (N_12914,N_12676,N_12673);
nor U12915 (N_12915,N_12718,N_12730);
nand U12916 (N_12916,N_12739,N_12757);
nor U12917 (N_12917,N_12692,N_12668);
xor U12918 (N_12918,N_12648,N_12647);
nor U12919 (N_12919,N_12753,N_12663);
nand U12920 (N_12920,N_12751,N_12790);
xnor U12921 (N_12921,N_12682,N_12729);
nand U12922 (N_12922,N_12679,N_12680);
nand U12923 (N_12923,N_12787,N_12695);
nor U12924 (N_12924,N_12731,N_12761);
nor U12925 (N_12925,N_12767,N_12739);
nor U12926 (N_12926,N_12667,N_12711);
or U12927 (N_12927,N_12767,N_12667);
nor U12928 (N_12928,N_12746,N_12689);
nor U12929 (N_12929,N_12649,N_12747);
nand U12930 (N_12930,N_12723,N_12663);
nand U12931 (N_12931,N_12790,N_12693);
and U12932 (N_12932,N_12687,N_12760);
or U12933 (N_12933,N_12764,N_12677);
nor U12934 (N_12934,N_12646,N_12756);
nand U12935 (N_12935,N_12780,N_12705);
nand U12936 (N_12936,N_12771,N_12733);
nand U12937 (N_12937,N_12735,N_12691);
nor U12938 (N_12938,N_12688,N_12702);
nand U12939 (N_12939,N_12703,N_12660);
xnor U12940 (N_12940,N_12684,N_12744);
and U12941 (N_12941,N_12640,N_12729);
or U12942 (N_12942,N_12771,N_12722);
and U12943 (N_12943,N_12793,N_12756);
nand U12944 (N_12944,N_12749,N_12645);
and U12945 (N_12945,N_12695,N_12658);
and U12946 (N_12946,N_12678,N_12706);
or U12947 (N_12947,N_12729,N_12684);
nand U12948 (N_12948,N_12646,N_12772);
xnor U12949 (N_12949,N_12709,N_12767);
or U12950 (N_12950,N_12695,N_12646);
nor U12951 (N_12951,N_12764,N_12761);
or U12952 (N_12952,N_12650,N_12790);
xor U12953 (N_12953,N_12716,N_12707);
nand U12954 (N_12954,N_12701,N_12688);
nand U12955 (N_12955,N_12774,N_12667);
or U12956 (N_12956,N_12719,N_12781);
or U12957 (N_12957,N_12695,N_12741);
nand U12958 (N_12958,N_12799,N_12790);
nand U12959 (N_12959,N_12655,N_12695);
nor U12960 (N_12960,N_12953,N_12838);
xnor U12961 (N_12961,N_12872,N_12950);
xor U12962 (N_12962,N_12843,N_12952);
nor U12963 (N_12963,N_12893,N_12906);
nor U12964 (N_12964,N_12850,N_12949);
nand U12965 (N_12965,N_12932,N_12867);
or U12966 (N_12966,N_12920,N_12862);
nor U12967 (N_12967,N_12846,N_12842);
nand U12968 (N_12968,N_12848,N_12923);
xor U12969 (N_12969,N_12927,N_12802);
xor U12970 (N_12970,N_12814,N_12922);
or U12971 (N_12971,N_12878,N_12849);
or U12972 (N_12972,N_12921,N_12807);
xor U12973 (N_12973,N_12826,N_12855);
nand U12974 (N_12974,N_12942,N_12844);
or U12975 (N_12975,N_12874,N_12813);
nand U12976 (N_12976,N_12901,N_12957);
xor U12977 (N_12977,N_12888,N_12915);
or U12978 (N_12978,N_12903,N_12871);
nand U12979 (N_12979,N_12837,N_12944);
xor U12980 (N_12980,N_12860,N_12836);
nor U12981 (N_12981,N_12956,N_12830);
nand U12982 (N_12982,N_12812,N_12913);
and U12983 (N_12983,N_12821,N_12958);
xnor U12984 (N_12984,N_12820,N_12881);
nor U12985 (N_12985,N_12847,N_12909);
or U12986 (N_12986,N_12822,N_12869);
nand U12987 (N_12987,N_12818,N_12919);
and U12988 (N_12988,N_12943,N_12887);
nor U12989 (N_12989,N_12925,N_12839);
and U12990 (N_12990,N_12879,N_12800);
nand U12991 (N_12991,N_12833,N_12864);
and U12992 (N_12992,N_12866,N_12936);
and U12993 (N_12993,N_12870,N_12811);
xor U12994 (N_12994,N_12890,N_12828);
and U12995 (N_12995,N_12819,N_12889);
and U12996 (N_12996,N_12908,N_12829);
xnor U12997 (N_12997,N_12959,N_12857);
xor U12998 (N_12998,N_12840,N_12824);
xor U12999 (N_12999,N_12894,N_12801);
or U13000 (N_13000,N_12896,N_12933);
or U13001 (N_13001,N_12805,N_12907);
and U13002 (N_13002,N_12905,N_12954);
or U13003 (N_13003,N_12804,N_12930);
nand U13004 (N_13004,N_12924,N_12806);
or U13005 (N_13005,N_12876,N_12886);
and U13006 (N_13006,N_12823,N_12868);
and U13007 (N_13007,N_12934,N_12895);
or U13008 (N_13008,N_12834,N_12831);
nor U13009 (N_13009,N_12861,N_12841);
nor U13010 (N_13010,N_12947,N_12946);
and U13011 (N_13011,N_12825,N_12809);
nand U13012 (N_13012,N_12918,N_12882);
xnor U13013 (N_13013,N_12827,N_12935);
nor U13014 (N_13014,N_12945,N_12955);
and U13015 (N_13015,N_12897,N_12939);
and U13016 (N_13016,N_12928,N_12883);
nand U13017 (N_13017,N_12817,N_12938);
nor U13018 (N_13018,N_12931,N_12916);
nand U13019 (N_13019,N_12835,N_12852);
or U13020 (N_13020,N_12803,N_12912);
or U13021 (N_13021,N_12865,N_12951);
xor U13022 (N_13022,N_12832,N_12851);
xor U13023 (N_13023,N_12926,N_12911);
or U13024 (N_13024,N_12808,N_12904);
nand U13025 (N_13025,N_12875,N_12948);
and U13026 (N_13026,N_12900,N_12863);
and U13027 (N_13027,N_12884,N_12899);
xor U13028 (N_13028,N_12941,N_12816);
nand U13029 (N_13029,N_12810,N_12880);
or U13030 (N_13030,N_12856,N_12885);
and U13031 (N_13031,N_12902,N_12917);
or U13032 (N_13032,N_12891,N_12929);
xnor U13033 (N_13033,N_12853,N_12858);
nand U13034 (N_13034,N_12845,N_12854);
nand U13035 (N_13035,N_12898,N_12873);
nand U13036 (N_13036,N_12815,N_12892);
nand U13037 (N_13037,N_12940,N_12910);
nand U13038 (N_13038,N_12914,N_12859);
nand U13039 (N_13039,N_12937,N_12877);
nor U13040 (N_13040,N_12929,N_12802);
nand U13041 (N_13041,N_12914,N_12916);
and U13042 (N_13042,N_12842,N_12803);
nor U13043 (N_13043,N_12954,N_12858);
nand U13044 (N_13044,N_12843,N_12915);
nand U13045 (N_13045,N_12855,N_12927);
or U13046 (N_13046,N_12941,N_12841);
xnor U13047 (N_13047,N_12881,N_12946);
xnor U13048 (N_13048,N_12944,N_12854);
nor U13049 (N_13049,N_12838,N_12927);
or U13050 (N_13050,N_12883,N_12910);
xnor U13051 (N_13051,N_12888,N_12883);
nand U13052 (N_13052,N_12839,N_12945);
or U13053 (N_13053,N_12954,N_12832);
or U13054 (N_13054,N_12956,N_12916);
nand U13055 (N_13055,N_12808,N_12813);
and U13056 (N_13056,N_12913,N_12869);
nor U13057 (N_13057,N_12928,N_12814);
xnor U13058 (N_13058,N_12869,N_12956);
and U13059 (N_13059,N_12940,N_12926);
nor U13060 (N_13060,N_12849,N_12888);
nor U13061 (N_13061,N_12844,N_12893);
nand U13062 (N_13062,N_12810,N_12947);
or U13063 (N_13063,N_12931,N_12934);
xor U13064 (N_13064,N_12929,N_12875);
nand U13065 (N_13065,N_12918,N_12939);
nor U13066 (N_13066,N_12874,N_12913);
nand U13067 (N_13067,N_12930,N_12919);
nor U13068 (N_13068,N_12801,N_12852);
nand U13069 (N_13069,N_12915,N_12844);
nor U13070 (N_13070,N_12807,N_12877);
nor U13071 (N_13071,N_12868,N_12829);
xnor U13072 (N_13072,N_12898,N_12863);
nand U13073 (N_13073,N_12922,N_12860);
nand U13074 (N_13074,N_12895,N_12940);
or U13075 (N_13075,N_12847,N_12950);
nand U13076 (N_13076,N_12958,N_12940);
and U13077 (N_13077,N_12935,N_12808);
xor U13078 (N_13078,N_12956,N_12942);
and U13079 (N_13079,N_12871,N_12897);
nand U13080 (N_13080,N_12946,N_12850);
or U13081 (N_13081,N_12936,N_12948);
nor U13082 (N_13082,N_12947,N_12881);
and U13083 (N_13083,N_12874,N_12859);
and U13084 (N_13084,N_12903,N_12928);
or U13085 (N_13085,N_12809,N_12950);
xor U13086 (N_13086,N_12920,N_12848);
nand U13087 (N_13087,N_12937,N_12860);
xor U13088 (N_13088,N_12817,N_12959);
or U13089 (N_13089,N_12943,N_12894);
nor U13090 (N_13090,N_12849,N_12801);
or U13091 (N_13091,N_12861,N_12931);
nor U13092 (N_13092,N_12844,N_12865);
nor U13093 (N_13093,N_12886,N_12874);
nor U13094 (N_13094,N_12916,N_12871);
and U13095 (N_13095,N_12828,N_12853);
and U13096 (N_13096,N_12902,N_12956);
xor U13097 (N_13097,N_12924,N_12833);
nand U13098 (N_13098,N_12896,N_12905);
nand U13099 (N_13099,N_12917,N_12887);
nand U13100 (N_13100,N_12811,N_12884);
nor U13101 (N_13101,N_12804,N_12850);
and U13102 (N_13102,N_12908,N_12934);
nor U13103 (N_13103,N_12837,N_12909);
and U13104 (N_13104,N_12872,N_12938);
or U13105 (N_13105,N_12822,N_12835);
xor U13106 (N_13106,N_12800,N_12833);
and U13107 (N_13107,N_12831,N_12946);
and U13108 (N_13108,N_12843,N_12851);
xor U13109 (N_13109,N_12860,N_12825);
or U13110 (N_13110,N_12864,N_12848);
and U13111 (N_13111,N_12916,N_12864);
or U13112 (N_13112,N_12837,N_12890);
nor U13113 (N_13113,N_12933,N_12871);
or U13114 (N_13114,N_12882,N_12943);
nand U13115 (N_13115,N_12803,N_12917);
nor U13116 (N_13116,N_12946,N_12920);
and U13117 (N_13117,N_12881,N_12882);
xor U13118 (N_13118,N_12818,N_12901);
and U13119 (N_13119,N_12821,N_12807);
or U13120 (N_13120,N_13056,N_13014);
nand U13121 (N_13121,N_13036,N_13053);
and U13122 (N_13122,N_13099,N_13073);
and U13123 (N_13123,N_13078,N_13066);
or U13124 (N_13124,N_13035,N_13018);
or U13125 (N_13125,N_13091,N_13067);
nand U13126 (N_13126,N_13098,N_13089);
and U13127 (N_13127,N_13088,N_13023);
nand U13128 (N_13128,N_13074,N_12961);
nor U13129 (N_13129,N_13049,N_12976);
nand U13130 (N_13130,N_13046,N_13101);
and U13131 (N_13131,N_13076,N_13002);
xnor U13132 (N_13132,N_13079,N_12970);
nor U13133 (N_13133,N_13034,N_13058);
nand U13134 (N_13134,N_13059,N_13011);
nand U13135 (N_13135,N_13119,N_13062);
nor U13136 (N_13136,N_13107,N_13008);
xnor U13137 (N_13137,N_12988,N_13081);
xnor U13138 (N_13138,N_12977,N_13004);
nand U13139 (N_13139,N_13031,N_13103);
nor U13140 (N_13140,N_12968,N_13096);
nor U13141 (N_13141,N_13116,N_12998);
or U13142 (N_13142,N_13080,N_13020);
nor U13143 (N_13143,N_13001,N_12983);
nand U13144 (N_13144,N_12996,N_13012);
nor U13145 (N_13145,N_12963,N_12964);
nand U13146 (N_13146,N_12991,N_12995);
and U13147 (N_13147,N_12990,N_13111);
or U13148 (N_13148,N_13108,N_13041);
and U13149 (N_13149,N_13075,N_13006);
nor U13150 (N_13150,N_13069,N_12973);
and U13151 (N_13151,N_13113,N_13115);
or U13152 (N_13152,N_13092,N_13022);
xnor U13153 (N_13153,N_13044,N_13095);
nor U13154 (N_13154,N_13028,N_13112);
and U13155 (N_13155,N_12975,N_13070);
or U13156 (N_13156,N_13043,N_13077);
nand U13157 (N_13157,N_13106,N_13032);
or U13158 (N_13158,N_12978,N_13013);
xnor U13159 (N_13159,N_13054,N_13042);
xnor U13160 (N_13160,N_13068,N_13010);
and U13161 (N_13161,N_13033,N_12994);
or U13162 (N_13162,N_13085,N_13021);
nor U13163 (N_13163,N_13051,N_12987);
or U13164 (N_13164,N_13114,N_12974);
xnor U13165 (N_13165,N_13037,N_13064);
and U13166 (N_13166,N_13060,N_13086);
or U13167 (N_13167,N_12997,N_13015);
xnor U13168 (N_13168,N_12993,N_12966);
nand U13169 (N_13169,N_12989,N_13057);
nor U13170 (N_13170,N_13029,N_13100);
or U13171 (N_13171,N_12985,N_13087);
or U13172 (N_13172,N_12981,N_13072);
nand U13173 (N_13173,N_13102,N_13007);
or U13174 (N_13174,N_13052,N_12984);
xor U13175 (N_13175,N_13000,N_13055);
and U13176 (N_13176,N_13083,N_13097);
and U13177 (N_13177,N_12972,N_13093);
xor U13178 (N_13178,N_12979,N_13027);
nor U13179 (N_13179,N_12960,N_13048);
nand U13180 (N_13180,N_13065,N_13117);
nor U13181 (N_13181,N_13025,N_13090);
and U13182 (N_13182,N_13118,N_13084);
nand U13183 (N_13183,N_13039,N_13071);
xnor U13184 (N_13184,N_13061,N_13050);
or U13185 (N_13185,N_12969,N_13105);
nor U13186 (N_13186,N_13110,N_13104);
and U13187 (N_13187,N_12967,N_13094);
or U13188 (N_13188,N_13026,N_13030);
xor U13189 (N_13189,N_13016,N_12965);
or U13190 (N_13190,N_12971,N_13009);
or U13191 (N_13191,N_13017,N_12986);
nor U13192 (N_13192,N_12992,N_13024);
xor U13193 (N_13193,N_12980,N_13019);
or U13194 (N_13194,N_13082,N_13040);
xnor U13195 (N_13195,N_13038,N_13003);
xor U13196 (N_13196,N_12999,N_13047);
xor U13197 (N_13197,N_12982,N_13005);
nor U13198 (N_13198,N_13045,N_12962);
or U13199 (N_13199,N_13109,N_13063);
and U13200 (N_13200,N_13083,N_13067);
xor U13201 (N_13201,N_13009,N_13000);
xnor U13202 (N_13202,N_13021,N_13061);
and U13203 (N_13203,N_13091,N_13117);
nand U13204 (N_13204,N_13035,N_13098);
and U13205 (N_13205,N_12976,N_13080);
and U13206 (N_13206,N_12967,N_13114);
nand U13207 (N_13207,N_13075,N_12990);
xnor U13208 (N_13208,N_13107,N_12962);
and U13209 (N_13209,N_13093,N_13116);
or U13210 (N_13210,N_13071,N_12975);
and U13211 (N_13211,N_13068,N_12965);
nor U13212 (N_13212,N_13071,N_12965);
nand U13213 (N_13213,N_13017,N_12974);
nor U13214 (N_13214,N_13042,N_13036);
or U13215 (N_13215,N_13004,N_13045);
or U13216 (N_13216,N_12968,N_13086);
nand U13217 (N_13217,N_12965,N_12991);
nand U13218 (N_13218,N_12993,N_13061);
nor U13219 (N_13219,N_13111,N_13054);
nand U13220 (N_13220,N_13102,N_13042);
or U13221 (N_13221,N_13086,N_13052);
and U13222 (N_13222,N_13032,N_13033);
or U13223 (N_13223,N_13028,N_13023);
or U13224 (N_13224,N_13043,N_13074);
xor U13225 (N_13225,N_13108,N_13007);
and U13226 (N_13226,N_13035,N_13012);
nand U13227 (N_13227,N_13097,N_13003);
nor U13228 (N_13228,N_13057,N_13013);
or U13229 (N_13229,N_12962,N_12999);
xor U13230 (N_13230,N_13080,N_13100);
or U13231 (N_13231,N_13075,N_12987);
or U13232 (N_13232,N_12972,N_13049);
and U13233 (N_13233,N_12968,N_13076);
xor U13234 (N_13234,N_12966,N_13068);
nor U13235 (N_13235,N_13058,N_13062);
or U13236 (N_13236,N_13046,N_13084);
nand U13237 (N_13237,N_13061,N_13043);
or U13238 (N_13238,N_13117,N_13039);
nand U13239 (N_13239,N_13023,N_13055);
xnor U13240 (N_13240,N_13116,N_13060);
nor U13241 (N_13241,N_13022,N_13015);
and U13242 (N_13242,N_13027,N_13064);
nand U13243 (N_13243,N_13013,N_12975);
and U13244 (N_13244,N_12962,N_13109);
nand U13245 (N_13245,N_12980,N_13082);
nor U13246 (N_13246,N_12973,N_13000);
nor U13247 (N_13247,N_13010,N_12966);
nand U13248 (N_13248,N_13111,N_13040);
and U13249 (N_13249,N_13087,N_12986);
xnor U13250 (N_13250,N_13055,N_13040);
or U13251 (N_13251,N_13060,N_13075);
and U13252 (N_13252,N_13114,N_12983);
and U13253 (N_13253,N_12990,N_12986);
nor U13254 (N_13254,N_13117,N_12996);
nand U13255 (N_13255,N_13046,N_12978);
and U13256 (N_13256,N_12971,N_13017);
and U13257 (N_13257,N_12985,N_13002);
nand U13258 (N_13258,N_13103,N_13065);
or U13259 (N_13259,N_13046,N_13094);
nor U13260 (N_13260,N_13016,N_13117);
nor U13261 (N_13261,N_12981,N_13009);
nand U13262 (N_13262,N_13119,N_13076);
and U13263 (N_13263,N_12970,N_12991);
and U13264 (N_13264,N_13019,N_13112);
or U13265 (N_13265,N_12970,N_13076);
and U13266 (N_13266,N_13020,N_13066);
nand U13267 (N_13267,N_13041,N_13051);
and U13268 (N_13268,N_13080,N_13115);
and U13269 (N_13269,N_12973,N_12995);
and U13270 (N_13270,N_12977,N_13020);
and U13271 (N_13271,N_13074,N_13041);
xor U13272 (N_13272,N_13047,N_13006);
nor U13273 (N_13273,N_12973,N_13019);
xor U13274 (N_13274,N_12995,N_12998);
or U13275 (N_13275,N_13005,N_13098);
or U13276 (N_13276,N_12977,N_13078);
xor U13277 (N_13277,N_12981,N_13036);
nor U13278 (N_13278,N_12977,N_13051);
nand U13279 (N_13279,N_13058,N_13041);
and U13280 (N_13280,N_13176,N_13195);
nand U13281 (N_13281,N_13143,N_13130);
xnor U13282 (N_13282,N_13262,N_13148);
or U13283 (N_13283,N_13249,N_13182);
nor U13284 (N_13284,N_13158,N_13159);
nand U13285 (N_13285,N_13202,N_13234);
and U13286 (N_13286,N_13154,N_13172);
xor U13287 (N_13287,N_13198,N_13122);
or U13288 (N_13288,N_13131,N_13136);
nand U13289 (N_13289,N_13203,N_13173);
xnor U13290 (N_13290,N_13253,N_13192);
xor U13291 (N_13291,N_13137,N_13178);
nand U13292 (N_13292,N_13208,N_13126);
nand U13293 (N_13293,N_13144,N_13146);
xnor U13294 (N_13294,N_13248,N_13270);
xor U13295 (N_13295,N_13170,N_13211);
or U13296 (N_13296,N_13169,N_13240);
and U13297 (N_13297,N_13232,N_13269);
or U13298 (N_13298,N_13247,N_13220);
nor U13299 (N_13299,N_13121,N_13163);
xor U13300 (N_13300,N_13171,N_13256);
nor U13301 (N_13301,N_13227,N_13167);
xnor U13302 (N_13302,N_13205,N_13230);
nor U13303 (N_13303,N_13161,N_13251);
xnor U13304 (N_13304,N_13155,N_13194);
or U13305 (N_13305,N_13209,N_13207);
xor U13306 (N_13306,N_13162,N_13175);
nand U13307 (N_13307,N_13177,N_13224);
nor U13308 (N_13308,N_13246,N_13212);
or U13309 (N_13309,N_13165,N_13257);
xnor U13310 (N_13310,N_13245,N_13204);
nor U13311 (N_13311,N_13201,N_13250);
xnor U13312 (N_13312,N_13185,N_13156);
and U13313 (N_13313,N_13254,N_13123);
or U13314 (N_13314,N_13275,N_13186);
and U13315 (N_13315,N_13164,N_13229);
and U13316 (N_13316,N_13189,N_13141);
nor U13317 (N_13317,N_13222,N_13157);
nand U13318 (N_13318,N_13221,N_13268);
nor U13319 (N_13319,N_13225,N_13183);
nor U13320 (N_13320,N_13133,N_13277);
nor U13321 (N_13321,N_13150,N_13142);
nor U13322 (N_13322,N_13196,N_13197);
xnor U13323 (N_13323,N_13279,N_13266);
nor U13324 (N_13324,N_13235,N_13274);
or U13325 (N_13325,N_13124,N_13140);
or U13326 (N_13326,N_13184,N_13242);
nor U13327 (N_13327,N_13271,N_13139);
or U13328 (N_13328,N_13226,N_13135);
and U13329 (N_13329,N_13191,N_13236);
xnor U13330 (N_13330,N_13168,N_13187);
nor U13331 (N_13331,N_13193,N_13129);
and U13332 (N_13332,N_13120,N_13252);
or U13333 (N_13333,N_13128,N_13267);
nor U13334 (N_13334,N_13179,N_13160);
nand U13335 (N_13335,N_13174,N_13152);
and U13336 (N_13336,N_13218,N_13223);
xnor U13337 (N_13337,N_13149,N_13265);
or U13338 (N_13338,N_13166,N_13243);
nand U13339 (N_13339,N_13276,N_13216);
nor U13340 (N_13340,N_13199,N_13138);
nand U13341 (N_13341,N_13258,N_13239);
nor U13342 (N_13342,N_13238,N_13259);
xor U13343 (N_13343,N_13278,N_13214);
xnor U13344 (N_13344,N_13180,N_13153);
and U13345 (N_13345,N_13237,N_13206);
nand U13346 (N_13346,N_13233,N_13263);
nor U13347 (N_13347,N_13190,N_13147);
nor U13348 (N_13348,N_13228,N_13145);
nand U13349 (N_13349,N_13188,N_13261);
xor U13350 (N_13350,N_13272,N_13132);
nor U13351 (N_13351,N_13219,N_13213);
nor U13352 (N_13352,N_13200,N_13210);
and U13353 (N_13353,N_13134,N_13231);
xor U13354 (N_13354,N_13181,N_13127);
xnor U13355 (N_13355,N_13273,N_13151);
nor U13356 (N_13356,N_13255,N_13241);
and U13357 (N_13357,N_13125,N_13217);
nor U13358 (N_13358,N_13244,N_13215);
and U13359 (N_13359,N_13260,N_13264);
or U13360 (N_13360,N_13122,N_13179);
or U13361 (N_13361,N_13277,N_13270);
and U13362 (N_13362,N_13259,N_13146);
nor U13363 (N_13363,N_13168,N_13253);
and U13364 (N_13364,N_13141,N_13213);
or U13365 (N_13365,N_13270,N_13128);
xnor U13366 (N_13366,N_13274,N_13272);
nor U13367 (N_13367,N_13215,N_13165);
nand U13368 (N_13368,N_13174,N_13172);
or U13369 (N_13369,N_13215,N_13147);
xnor U13370 (N_13370,N_13129,N_13250);
or U13371 (N_13371,N_13203,N_13245);
xnor U13372 (N_13372,N_13264,N_13208);
or U13373 (N_13373,N_13260,N_13145);
or U13374 (N_13374,N_13236,N_13239);
nor U13375 (N_13375,N_13199,N_13160);
or U13376 (N_13376,N_13161,N_13268);
and U13377 (N_13377,N_13131,N_13189);
xnor U13378 (N_13378,N_13175,N_13186);
xor U13379 (N_13379,N_13219,N_13163);
and U13380 (N_13380,N_13175,N_13170);
nor U13381 (N_13381,N_13161,N_13137);
nor U13382 (N_13382,N_13270,N_13165);
nor U13383 (N_13383,N_13265,N_13193);
nand U13384 (N_13384,N_13151,N_13174);
nor U13385 (N_13385,N_13241,N_13212);
nand U13386 (N_13386,N_13259,N_13178);
nand U13387 (N_13387,N_13240,N_13228);
nor U13388 (N_13388,N_13226,N_13192);
and U13389 (N_13389,N_13159,N_13238);
xnor U13390 (N_13390,N_13127,N_13254);
or U13391 (N_13391,N_13249,N_13188);
and U13392 (N_13392,N_13121,N_13216);
and U13393 (N_13393,N_13228,N_13193);
nand U13394 (N_13394,N_13166,N_13220);
nand U13395 (N_13395,N_13252,N_13239);
and U13396 (N_13396,N_13120,N_13173);
nand U13397 (N_13397,N_13219,N_13212);
nand U13398 (N_13398,N_13147,N_13274);
nand U13399 (N_13399,N_13181,N_13141);
or U13400 (N_13400,N_13272,N_13204);
or U13401 (N_13401,N_13195,N_13273);
xor U13402 (N_13402,N_13272,N_13248);
or U13403 (N_13403,N_13274,N_13203);
xor U13404 (N_13404,N_13192,N_13221);
nand U13405 (N_13405,N_13258,N_13163);
and U13406 (N_13406,N_13163,N_13133);
or U13407 (N_13407,N_13135,N_13224);
nor U13408 (N_13408,N_13213,N_13191);
or U13409 (N_13409,N_13240,N_13170);
or U13410 (N_13410,N_13124,N_13194);
nand U13411 (N_13411,N_13243,N_13146);
nor U13412 (N_13412,N_13175,N_13199);
and U13413 (N_13413,N_13231,N_13165);
nor U13414 (N_13414,N_13133,N_13152);
or U13415 (N_13415,N_13124,N_13166);
or U13416 (N_13416,N_13273,N_13257);
xnor U13417 (N_13417,N_13161,N_13136);
nor U13418 (N_13418,N_13220,N_13152);
xnor U13419 (N_13419,N_13171,N_13145);
and U13420 (N_13420,N_13148,N_13242);
and U13421 (N_13421,N_13174,N_13179);
nor U13422 (N_13422,N_13175,N_13195);
nand U13423 (N_13423,N_13181,N_13172);
xnor U13424 (N_13424,N_13263,N_13158);
nor U13425 (N_13425,N_13137,N_13205);
or U13426 (N_13426,N_13250,N_13210);
or U13427 (N_13427,N_13159,N_13260);
xnor U13428 (N_13428,N_13252,N_13142);
xnor U13429 (N_13429,N_13218,N_13235);
nand U13430 (N_13430,N_13145,N_13269);
nand U13431 (N_13431,N_13180,N_13164);
or U13432 (N_13432,N_13125,N_13186);
nor U13433 (N_13433,N_13148,N_13140);
or U13434 (N_13434,N_13250,N_13258);
nor U13435 (N_13435,N_13264,N_13217);
nand U13436 (N_13436,N_13204,N_13207);
nand U13437 (N_13437,N_13162,N_13262);
and U13438 (N_13438,N_13220,N_13162);
nand U13439 (N_13439,N_13274,N_13156);
xor U13440 (N_13440,N_13397,N_13416);
and U13441 (N_13441,N_13323,N_13371);
nand U13442 (N_13442,N_13300,N_13421);
nor U13443 (N_13443,N_13410,N_13420);
xor U13444 (N_13444,N_13318,N_13301);
nand U13445 (N_13445,N_13435,N_13373);
or U13446 (N_13446,N_13297,N_13370);
nor U13447 (N_13447,N_13303,N_13401);
xnor U13448 (N_13448,N_13292,N_13426);
or U13449 (N_13449,N_13411,N_13293);
xor U13450 (N_13450,N_13415,N_13384);
nand U13451 (N_13451,N_13417,N_13307);
nand U13452 (N_13452,N_13389,N_13290);
xor U13453 (N_13453,N_13349,N_13310);
and U13454 (N_13454,N_13322,N_13386);
or U13455 (N_13455,N_13340,N_13359);
nand U13456 (N_13456,N_13330,N_13342);
or U13457 (N_13457,N_13332,N_13422);
nand U13458 (N_13458,N_13324,N_13352);
or U13459 (N_13459,N_13403,N_13368);
nand U13460 (N_13460,N_13394,N_13406);
or U13461 (N_13461,N_13383,N_13317);
nor U13462 (N_13462,N_13355,N_13432);
and U13463 (N_13463,N_13284,N_13306);
nand U13464 (N_13464,N_13280,N_13358);
nand U13465 (N_13465,N_13296,N_13378);
or U13466 (N_13466,N_13337,N_13412);
xnor U13467 (N_13467,N_13428,N_13391);
and U13468 (N_13468,N_13379,N_13302);
and U13469 (N_13469,N_13354,N_13424);
nand U13470 (N_13470,N_13305,N_13376);
nor U13471 (N_13471,N_13336,N_13309);
and U13472 (N_13472,N_13429,N_13436);
xor U13473 (N_13473,N_13427,N_13404);
nor U13474 (N_13474,N_13388,N_13304);
nand U13475 (N_13475,N_13419,N_13314);
nand U13476 (N_13476,N_13291,N_13347);
xnor U13477 (N_13477,N_13430,N_13283);
nand U13478 (N_13478,N_13335,N_13327);
nand U13479 (N_13479,N_13282,N_13295);
or U13480 (N_13480,N_13341,N_13367);
nor U13481 (N_13481,N_13413,N_13374);
nor U13482 (N_13482,N_13339,N_13438);
and U13483 (N_13483,N_13380,N_13294);
or U13484 (N_13484,N_13328,N_13329);
and U13485 (N_13485,N_13361,N_13363);
and U13486 (N_13486,N_13287,N_13423);
nand U13487 (N_13487,N_13392,N_13313);
and U13488 (N_13488,N_13326,N_13408);
nand U13489 (N_13489,N_13311,N_13405);
and U13490 (N_13490,N_13418,N_13299);
or U13491 (N_13491,N_13395,N_13316);
nand U13492 (N_13492,N_13369,N_13325);
and U13493 (N_13493,N_13320,N_13407);
nand U13494 (N_13494,N_13437,N_13312);
and U13495 (N_13495,N_13315,N_13393);
and U13496 (N_13496,N_13385,N_13346);
or U13497 (N_13497,N_13402,N_13356);
xor U13498 (N_13498,N_13319,N_13399);
or U13499 (N_13499,N_13344,N_13345);
or U13500 (N_13500,N_13382,N_13362);
and U13501 (N_13501,N_13364,N_13439);
nor U13502 (N_13502,N_13431,N_13353);
nand U13503 (N_13503,N_13433,N_13334);
or U13504 (N_13504,N_13414,N_13333);
or U13505 (N_13505,N_13400,N_13348);
xor U13506 (N_13506,N_13338,N_13298);
or U13507 (N_13507,N_13375,N_13366);
xnor U13508 (N_13508,N_13360,N_13377);
and U13509 (N_13509,N_13387,N_13286);
xnor U13510 (N_13510,N_13321,N_13288);
nand U13511 (N_13511,N_13351,N_13409);
nand U13512 (N_13512,N_13285,N_13365);
or U13513 (N_13513,N_13331,N_13372);
xnor U13514 (N_13514,N_13308,N_13289);
xnor U13515 (N_13515,N_13281,N_13425);
nand U13516 (N_13516,N_13396,N_13357);
nand U13517 (N_13517,N_13343,N_13390);
xor U13518 (N_13518,N_13350,N_13398);
xnor U13519 (N_13519,N_13381,N_13434);
and U13520 (N_13520,N_13281,N_13286);
nor U13521 (N_13521,N_13378,N_13404);
xnor U13522 (N_13522,N_13390,N_13401);
and U13523 (N_13523,N_13314,N_13369);
xor U13524 (N_13524,N_13297,N_13366);
nor U13525 (N_13525,N_13324,N_13439);
nand U13526 (N_13526,N_13329,N_13410);
and U13527 (N_13527,N_13355,N_13418);
xnor U13528 (N_13528,N_13373,N_13375);
or U13529 (N_13529,N_13393,N_13331);
nor U13530 (N_13530,N_13298,N_13366);
nand U13531 (N_13531,N_13294,N_13389);
nand U13532 (N_13532,N_13320,N_13410);
and U13533 (N_13533,N_13370,N_13317);
xnor U13534 (N_13534,N_13376,N_13400);
and U13535 (N_13535,N_13327,N_13316);
or U13536 (N_13536,N_13360,N_13361);
or U13537 (N_13537,N_13409,N_13426);
and U13538 (N_13538,N_13295,N_13330);
and U13539 (N_13539,N_13285,N_13314);
nand U13540 (N_13540,N_13317,N_13314);
and U13541 (N_13541,N_13342,N_13432);
nor U13542 (N_13542,N_13286,N_13405);
nor U13543 (N_13543,N_13320,N_13293);
xnor U13544 (N_13544,N_13352,N_13396);
or U13545 (N_13545,N_13300,N_13325);
nand U13546 (N_13546,N_13293,N_13285);
nand U13547 (N_13547,N_13367,N_13387);
or U13548 (N_13548,N_13397,N_13408);
xor U13549 (N_13549,N_13355,N_13280);
nor U13550 (N_13550,N_13325,N_13329);
xnor U13551 (N_13551,N_13424,N_13411);
nor U13552 (N_13552,N_13285,N_13325);
nor U13553 (N_13553,N_13291,N_13325);
xor U13554 (N_13554,N_13332,N_13386);
and U13555 (N_13555,N_13311,N_13411);
or U13556 (N_13556,N_13285,N_13404);
and U13557 (N_13557,N_13404,N_13419);
or U13558 (N_13558,N_13326,N_13311);
or U13559 (N_13559,N_13385,N_13325);
or U13560 (N_13560,N_13300,N_13331);
xnor U13561 (N_13561,N_13333,N_13374);
nand U13562 (N_13562,N_13280,N_13324);
and U13563 (N_13563,N_13433,N_13283);
nand U13564 (N_13564,N_13439,N_13421);
nand U13565 (N_13565,N_13307,N_13291);
nand U13566 (N_13566,N_13378,N_13420);
and U13567 (N_13567,N_13304,N_13395);
or U13568 (N_13568,N_13345,N_13310);
or U13569 (N_13569,N_13358,N_13343);
nor U13570 (N_13570,N_13348,N_13345);
nor U13571 (N_13571,N_13408,N_13329);
or U13572 (N_13572,N_13285,N_13439);
nand U13573 (N_13573,N_13439,N_13376);
nor U13574 (N_13574,N_13368,N_13335);
nand U13575 (N_13575,N_13363,N_13315);
xor U13576 (N_13576,N_13304,N_13334);
nand U13577 (N_13577,N_13364,N_13300);
and U13578 (N_13578,N_13357,N_13318);
nor U13579 (N_13579,N_13360,N_13302);
xor U13580 (N_13580,N_13296,N_13402);
or U13581 (N_13581,N_13413,N_13322);
nand U13582 (N_13582,N_13377,N_13338);
nor U13583 (N_13583,N_13379,N_13287);
and U13584 (N_13584,N_13432,N_13319);
and U13585 (N_13585,N_13315,N_13370);
or U13586 (N_13586,N_13333,N_13331);
nor U13587 (N_13587,N_13417,N_13364);
and U13588 (N_13588,N_13412,N_13352);
xnor U13589 (N_13589,N_13384,N_13407);
nor U13590 (N_13590,N_13291,N_13357);
or U13591 (N_13591,N_13280,N_13393);
or U13592 (N_13592,N_13435,N_13288);
nor U13593 (N_13593,N_13299,N_13347);
nand U13594 (N_13594,N_13423,N_13390);
xnor U13595 (N_13595,N_13433,N_13385);
or U13596 (N_13596,N_13317,N_13303);
nor U13597 (N_13597,N_13414,N_13385);
nand U13598 (N_13598,N_13413,N_13375);
xor U13599 (N_13599,N_13294,N_13297);
or U13600 (N_13600,N_13516,N_13542);
or U13601 (N_13601,N_13462,N_13586);
nand U13602 (N_13602,N_13587,N_13463);
nand U13603 (N_13603,N_13574,N_13511);
or U13604 (N_13604,N_13530,N_13464);
or U13605 (N_13605,N_13555,N_13580);
xor U13606 (N_13606,N_13577,N_13576);
and U13607 (N_13607,N_13581,N_13451);
and U13608 (N_13608,N_13459,N_13566);
xnor U13609 (N_13609,N_13519,N_13529);
xnor U13610 (N_13610,N_13489,N_13460);
xor U13611 (N_13611,N_13467,N_13441);
or U13612 (N_13612,N_13536,N_13598);
or U13613 (N_13613,N_13554,N_13453);
nand U13614 (N_13614,N_13589,N_13483);
and U13615 (N_13615,N_13477,N_13445);
nand U13616 (N_13616,N_13579,N_13492);
and U13617 (N_13617,N_13535,N_13571);
xor U13618 (N_13618,N_13550,N_13540);
and U13619 (N_13619,N_13545,N_13474);
or U13620 (N_13620,N_13565,N_13495);
or U13621 (N_13621,N_13564,N_13480);
nand U13622 (N_13622,N_13497,N_13570);
nand U13623 (N_13623,N_13446,N_13484);
or U13624 (N_13624,N_13491,N_13595);
nor U13625 (N_13625,N_13582,N_13557);
xor U13626 (N_13626,N_13493,N_13449);
and U13627 (N_13627,N_13520,N_13454);
and U13628 (N_13628,N_13599,N_13584);
nand U13629 (N_13629,N_13538,N_13585);
nor U13630 (N_13630,N_13503,N_13455);
and U13631 (N_13631,N_13515,N_13551);
or U13632 (N_13632,N_13468,N_13563);
xor U13633 (N_13633,N_13525,N_13509);
or U13634 (N_13634,N_13560,N_13440);
xnor U13635 (N_13635,N_13479,N_13593);
and U13636 (N_13636,N_13524,N_13457);
xnor U13637 (N_13637,N_13458,N_13573);
nand U13638 (N_13638,N_13522,N_13537);
and U13639 (N_13639,N_13465,N_13561);
xor U13640 (N_13640,N_13471,N_13517);
or U13641 (N_13641,N_13442,N_13568);
nand U13642 (N_13642,N_13447,N_13578);
and U13643 (N_13643,N_13508,N_13498);
nand U13644 (N_13644,N_13473,N_13443);
xor U13645 (N_13645,N_13583,N_13481);
nor U13646 (N_13646,N_13528,N_13518);
nor U13647 (N_13647,N_13590,N_13504);
and U13648 (N_13648,N_13521,N_13547);
or U13649 (N_13649,N_13549,N_13539);
and U13650 (N_13650,N_13534,N_13562);
xnor U13651 (N_13651,N_13532,N_13448);
xor U13652 (N_13652,N_13500,N_13487);
nor U13653 (N_13653,N_13548,N_13514);
nor U13654 (N_13654,N_13472,N_13502);
nor U13655 (N_13655,N_13569,N_13507);
xnor U13656 (N_13656,N_13501,N_13588);
nor U13657 (N_13657,N_13450,N_13526);
nor U13658 (N_13658,N_13469,N_13470);
or U13659 (N_13659,N_13496,N_13556);
xnor U13660 (N_13660,N_13461,N_13553);
nor U13661 (N_13661,N_13531,N_13478);
nand U13662 (N_13662,N_13490,N_13466);
xnor U13663 (N_13663,N_13567,N_13486);
or U13664 (N_13664,N_13559,N_13512);
or U13665 (N_13665,N_13527,N_13543);
nand U13666 (N_13666,N_13488,N_13541);
nand U13667 (N_13667,N_13558,N_13594);
xor U13668 (N_13668,N_13452,N_13482);
xor U13669 (N_13669,N_13552,N_13506);
or U13670 (N_13670,N_13513,N_13523);
nor U13671 (N_13671,N_13485,N_13456);
and U13672 (N_13672,N_13505,N_13475);
and U13673 (N_13673,N_13444,N_13575);
nand U13674 (N_13674,N_13596,N_13572);
xor U13675 (N_13675,N_13510,N_13494);
nor U13676 (N_13676,N_13592,N_13499);
nor U13677 (N_13677,N_13597,N_13533);
or U13678 (N_13678,N_13591,N_13476);
nor U13679 (N_13679,N_13544,N_13546);
nor U13680 (N_13680,N_13549,N_13458);
and U13681 (N_13681,N_13490,N_13562);
xor U13682 (N_13682,N_13519,N_13483);
xnor U13683 (N_13683,N_13563,N_13561);
and U13684 (N_13684,N_13525,N_13466);
or U13685 (N_13685,N_13596,N_13537);
nor U13686 (N_13686,N_13540,N_13558);
nor U13687 (N_13687,N_13464,N_13589);
nor U13688 (N_13688,N_13567,N_13508);
nor U13689 (N_13689,N_13461,N_13542);
nand U13690 (N_13690,N_13548,N_13562);
xor U13691 (N_13691,N_13501,N_13576);
nand U13692 (N_13692,N_13554,N_13468);
nor U13693 (N_13693,N_13498,N_13575);
or U13694 (N_13694,N_13497,N_13481);
or U13695 (N_13695,N_13449,N_13516);
nand U13696 (N_13696,N_13576,N_13550);
nand U13697 (N_13697,N_13484,N_13554);
nor U13698 (N_13698,N_13497,N_13508);
nor U13699 (N_13699,N_13450,N_13444);
xor U13700 (N_13700,N_13507,N_13536);
and U13701 (N_13701,N_13569,N_13448);
or U13702 (N_13702,N_13442,N_13562);
xnor U13703 (N_13703,N_13456,N_13516);
and U13704 (N_13704,N_13563,N_13524);
or U13705 (N_13705,N_13577,N_13489);
nor U13706 (N_13706,N_13476,N_13471);
and U13707 (N_13707,N_13486,N_13525);
and U13708 (N_13708,N_13545,N_13554);
nor U13709 (N_13709,N_13588,N_13528);
and U13710 (N_13710,N_13450,N_13459);
nor U13711 (N_13711,N_13441,N_13542);
xnor U13712 (N_13712,N_13444,N_13506);
or U13713 (N_13713,N_13456,N_13534);
xor U13714 (N_13714,N_13555,N_13592);
and U13715 (N_13715,N_13474,N_13533);
and U13716 (N_13716,N_13520,N_13495);
xnor U13717 (N_13717,N_13462,N_13560);
nand U13718 (N_13718,N_13581,N_13570);
or U13719 (N_13719,N_13567,N_13583);
or U13720 (N_13720,N_13572,N_13588);
nand U13721 (N_13721,N_13578,N_13460);
nor U13722 (N_13722,N_13500,N_13576);
nor U13723 (N_13723,N_13587,N_13561);
and U13724 (N_13724,N_13445,N_13492);
nor U13725 (N_13725,N_13477,N_13461);
and U13726 (N_13726,N_13450,N_13449);
or U13727 (N_13727,N_13498,N_13545);
nor U13728 (N_13728,N_13597,N_13482);
nand U13729 (N_13729,N_13581,N_13459);
xor U13730 (N_13730,N_13584,N_13464);
xor U13731 (N_13731,N_13509,N_13593);
nor U13732 (N_13732,N_13519,N_13464);
or U13733 (N_13733,N_13544,N_13597);
xor U13734 (N_13734,N_13456,N_13567);
or U13735 (N_13735,N_13598,N_13490);
nand U13736 (N_13736,N_13468,N_13517);
nor U13737 (N_13737,N_13492,N_13497);
nor U13738 (N_13738,N_13571,N_13466);
nor U13739 (N_13739,N_13548,N_13483);
and U13740 (N_13740,N_13528,N_13466);
and U13741 (N_13741,N_13543,N_13525);
nand U13742 (N_13742,N_13505,N_13479);
or U13743 (N_13743,N_13575,N_13591);
and U13744 (N_13744,N_13590,N_13543);
and U13745 (N_13745,N_13546,N_13512);
nand U13746 (N_13746,N_13475,N_13558);
or U13747 (N_13747,N_13576,N_13535);
xor U13748 (N_13748,N_13507,N_13494);
xor U13749 (N_13749,N_13498,N_13455);
nand U13750 (N_13750,N_13501,N_13449);
or U13751 (N_13751,N_13594,N_13452);
nor U13752 (N_13752,N_13540,N_13496);
xnor U13753 (N_13753,N_13592,N_13451);
nor U13754 (N_13754,N_13557,N_13499);
nor U13755 (N_13755,N_13549,N_13520);
nand U13756 (N_13756,N_13556,N_13444);
nor U13757 (N_13757,N_13514,N_13444);
nand U13758 (N_13758,N_13570,N_13517);
nand U13759 (N_13759,N_13519,N_13541);
nand U13760 (N_13760,N_13735,N_13749);
nand U13761 (N_13761,N_13618,N_13600);
or U13762 (N_13762,N_13742,N_13734);
xnor U13763 (N_13763,N_13638,N_13623);
nor U13764 (N_13764,N_13673,N_13661);
nor U13765 (N_13765,N_13696,N_13739);
xnor U13766 (N_13766,N_13677,N_13603);
and U13767 (N_13767,N_13645,N_13681);
xor U13768 (N_13768,N_13684,N_13699);
nand U13769 (N_13769,N_13701,N_13616);
nand U13770 (N_13770,N_13624,N_13604);
xor U13771 (N_13771,N_13729,N_13695);
nand U13772 (N_13772,N_13757,N_13721);
or U13773 (N_13773,N_13607,N_13708);
nand U13774 (N_13774,N_13746,N_13644);
xor U13775 (N_13775,N_13724,N_13690);
xnor U13776 (N_13776,N_13732,N_13610);
xnor U13777 (N_13777,N_13743,N_13647);
or U13778 (N_13778,N_13631,N_13714);
nor U13779 (N_13779,N_13754,N_13637);
and U13780 (N_13780,N_13656,N_13633);
nand U13781 (N_13781,N_13665,N_13628);
nand U13782 (N_13782,N_13731,N_13651);
xor U13783 (N_13783,N_13745,N_13671);
nor U13784 (N_13784,N_13630,N_13700);
and U13785 (N_13785,N_13640,N_13682);
nand U13786 (N_13786,N_13641,N_13626);
nor U13787 (N_13787,N_13726,N_13691);
and U13788 (N_13788,N_13635,N_13722);
or U13789 (N_13789,N_13759,N_13702);
nor U13790 (N_13790,N_13715,N_13639);
and U13791 (N_13791,N_13613,N_13723);
or U13792 (N_13792,N_13711,N_13755);
and U13793 (N_13793,N_13718,N_13636);
nand U13794 (N_13794,N_13752,N_13649);
nand U13795 (N_13795,N_13625,N_13683);
and U13796 (N_13796,N_13713,N_13679);
xor U13797 (N_13797,N_13685,N_13663);
xor U13798 (N_13798,N_13704,N_13697);
and U13799 (N_13799,N_13614,N_13741);
xnor U13800 (N_13800,N_13693,N_13632);
or U13801 (N_13801,N_13717,N_13712);
or U13802 (N_13802,N_13687,N_13688);
nand U13803 (N_13803,N_13669,N_13716);
or U13804 (N_13804,N_13605,N_13747);
nor U13805 (N_13805,N_13620,N_13666);
or U13806 (N_13806,N_13689,N_13672);
nor U13807 (N_13807,N_13660,N_13608);
xor U13808 (N_13808,N_13675,N_13642);
nor U13809 (N_13809,N_13692,N_13733);
or U13810 (N_13810,N_13740,N_13686);
or U13811 (N_13811,N_13706,N_13621);
or U13812 (N_13812,N_13748,N_13676);
or U13813 (N_13813,N_13667,N_13727);
xnor U13814 (N_13814,N_13674,N_13670);
or U13815 (N_13815,N_13646,N_13709);
nor U13816 (N_13816,N_13627,N_13606);
and U13817 (N_13817,N_13659,N_13662);
or U13818 (N_13818,N_13615,N_13705);
xnor U13819 (N_13819,N_13629,N_13728);
xnor U13820 (N_13820,N_13758,N_13744);
nor U13821 (N_13821,N_13736,N_13668);
and U13822 (N_13822,N_13703,N_13707);
or U13823 (N_13823,N_13619,N_13680);
nor U13824 (N_13824,N_13652,N_13725);
nand U13825 (N_13825,N_13678,N_13657);
xor U13826 (N_13826,N_13750,N_13738);
nor U13827 (N_13827,N_13650,N_13654);
nor U13828 (N_13828,N_13609,N_13710);
xnor U13829 (N_13829,N_13694,N_13719);
nand U13830 (N_13830,N_13648,N_13602);
xnor U13831 (N_13831,N_13751,N_13611);
nand U13832 (N_13832,N_13753,N_13730);
xnor U13833 (N_13833,N_13653,N_13655);
nand U13834 (N_13834,N_13698,N_13617);
and U13835 (N_13835,N_13622,N_13601);
or U13836 (N_13836,N_13643,N_13737);
xor U13837 (N_13837,N_13634,N_13756);
and U13838 (N_13838,N_13612,N_13720);
and U13839 (N_13839,N_13658,N_13664);
and U13840 (N_13840,N_13714,N_13756);
nand U13841 (N_13841,N_13655,N_13755);
xor U13842 (N_13842,N_13621,N_13601);
nor U13843 (N_13843,N_13748,N_13738);
or U13844 (N_13844,N_13724,N_13615);
or U13845 (N_13845,N_13604,N_13681);
xor U13846 (N_13846,N_13629,N_13676);
and U13847 (N_13847,N_13668,N_13621);
xnor U13848 (N_13848,N_13628,N_13608);
and U13849 (N_13849,N_13717,N_13649);
nor U13850 (N_13850,N_13718,N_13615);
nand U13851 (N_13851,N_13610,N_13677);
nand U13852 (N_13852,N_13644,N_13694);
nand U13853 (N_13853,N_13605,N_13625);
or U13854 (N_13854,N_13607,N_13752);
nand U13855 (N_13855,N_13707,N_13605);
nand U13856 (N_13856,N_13699,N_13726);
nor U13857 (N_13857,N_13698,N_13653);
xor U13858 (N_13858,N_13667,N_13708);
and U13859 (N_13859,N_13741,N_13754);
and U13860 (N_13860,N_13617,N_13703);
and U13861 (N_13861,N_13634,N_13612);
nor U13862 (N_13862,N_13757,N_13734);
nand U13863 (N_13863,N_13623,N_13631);
or U13864 (N_13864,N_13646,N_13614);
xnor U13865 (N_13865,N_13607,N_13749);
xnor U13866 (N_13866,N_13713,N_13641);
xor U13867 (N_13867,N_13607,N_13726);
xnor U13868 (N_13868,N_13717,N_13618);
and U13869 (N_13869,N_13702,N_13721);
and U13870 (N_13870,N_13749,N_13672);
nand U13871 (N_13871,N_13715,N_13731);
or U13872 (N_13872,N_13644,N_13603);
xor U13873 (N_13873,N_13737,N_13758);
or U13874 (N_13874,N_13729,N_13752);
nor U13875 (N_13875,N_13669,N_13742);
nor U13876 (N_13876,N_13644,N_13691);
and U13877 (N_13877,N_13754,N_13702);
nor U13878 (N_13878,N_13672,N_13710);
nor U13879 (N_13879,N_13680,N_13600);
and U13880 (N_13880,N_13660,N_13604);
nand U13881 (N_13881,N_13622,N_13605);
nand U13882 (N_13882,N_13613,N_13757);
and U13883 (N_13883,N_13692,N_13676);
xnor U13884 (N_13884,N_13643,N_13742);
or U13885 (N_13885,N_13657,N_13752);
and U13886 (N_13886,N_13662,N_13607);
nor U13887 (N_13887,N_13706,N_13615);
or U13888 (N_13888,N_13734,N_13744);
xor U13889 (N_13889,N_13749,N_13739);
nor U13890 (N_13890,N_13622,N_13682);
xnor U13891 (N_13891,N_13758,N_13704);
or U13892 (N_13892,N_13697,N_13713);
xnor U13893 (N_13893,N_13755,N_13660);
xor U13894 (N_13894,N_13668,N_13676);
nand U13895 (N_13895,N_13661,N_13708);
nand U13896 (N_13896,N_13749,N_13606);
and U13897 (N_13897,N_13642,N_13724);
nor U13898 (N_13898,N_13637,N_13746);
or U13899 (N_13899,N_13653,N_13666);
or U13900 (N_13900,N_13639,N_13718);
and U13901 (N_13901,N_13651,N_13712);
nand U13902 (N_13902,N_13675,N_13742);
nor U13903 (N_13903,N_13711,N_13625);
nand U13904 (N_13904,N_13621,N_13707);
and U13905 (N_13905,N_13660,N_13717);
and U13906 (N_13906,N_13751,N_13677);
nand U13907 (N_13907,N_13681,N_13633);
and U13908 (N_13908,N_13684,N_13628);
or U13909 (N_13909,N_13759,N_13728);
xor U13910 (N_13910,N_13757,N_13609);
xnor U13911 (N_13911,N_13678,N_13681);
xnor U13912 (N_13912,N_13677,N_13622);
and U13913 (N_13913,N_13615,N_13690);
nor U13914 (N_13914,N_13670,N_13635);
nor U13915 (N_13915,N_13704,N_13615);
nor U13916 (N_13916,N_13640,N_13707);
xor U13917 (N_13917,N_13741,N_13610);
nor U13918 (N_13918,N_13609,N_13737);
xnor U13919 (N_13919,N_13609,N_13601);
xor U13920 (N_13920,N_13859,N_13796);
and U13921 (N_13921,N_13809,N_13771);
or U13922 (N_13922,N_13886,N_13909);
xor U13923 (N_13923,N_13849,N_13778);
nand U13924 (N_13924,N_13895,N_13835);
and U13925 (N_13925,N_13917,N_13904);
or U13926 (N_13926,N_13913,N_13916);
xnor U13927 (N_13927,N_13897,N_13903);
nor U13928 (N_13928,N_13877,N_13802);
xor U13929 (N_13929,N_13779,N_13889);
xnor U13930 (N_13930,N_13881,N_13797);
nand U13931 (N_13931,N_13892,N_13838);
and U13932 (N_13932,N_13828,N_13861);
nand U13933 (N_13933,N_13775,N_13788);
or U13934 (N_13934,N_13882,N_13815);
nand U13935 (N_13935,N_13840,N_13898);
nand U13936 (N_13936,N_13846,N_13764);
nor U13937 (N_13937,N_13787,N_13801);
xnor U13938 (N_13938,N_13906,N_13768);
nand U13939 (N_13939,N_13890,N_13833);
nand U13940 (N_13940,N_13847,N_13832);
xnor U13941 (N_13941,N_13883,N_13762);
nand U13942 (N_13942,N_13869,N_13765);
xnor U13943 (N_13943,N_13781,N_13839);
xnor U13944 (N_13944,N_13866,N_13767);
and U13945 (N_13945,N_13805,N_13760);
xor U13946 (N_13946,N_13893,N_13800);
or U13947 (N_13947,N_13836,N_13769);
and U13948 (N_13948,N_13915,N_13848);
nor U13949 (N_13949,N_13865,N_13885);
nor U13950 (N_13950,N_13777,N_13891);
nand U13951 (N_13951,N_13783,N_13867);
or U13952 (N_13952,N_13845,N_13776);
xor U13953 (N_13953,N_13808,N_13824);
and U13954 (N_13954,N_13878,N_13790);
nor U13955 (N_13955,N_13841,N_13894);
and U13956 (N_13956,N_13795,N_13887);
and U13957 (N_13957,N_13870,N_13819);
and U13958 (N_13958,N_13884,N_13856);
and U13959 (N_13959,N_13818,N_13905);
nor U13960 (N_13960,N_13851,N_13902);
or U13961 (N_13961,N_13873,N_13914);
and U13962 (N_13962,N_13912,N_13774);
xnor U13963 (N_13963,N_13860,N_13812);
xor U13964 (N_13964,N_13785,N_13766);
and U13965 (N_13965,N_13871,N_13780);
nor U13966 (N_13966,N_13763,N_13784);
or U13967 (N_13967,N_13872,N_13830);
nand U13968 (N_13968,N_13789,N_13829);
nor U13969 (N_13969,N_13794,N_13852);
or U13970 (N_13970,N_13864,N_13798);
and U13971 (N_13971,N_13854,N_13806);
or U13972 (N_13972,N_13817,N_13857);
xor U13973 (N_13973,N_13814,N_13834);
nand U13974 (N_13974,N_13772,N_13799);
and U13975 (N_13975,N_13807,N_13825);
and U13976 (N_13976,N_13910,N_13761);
nand U13977 (N_13977,N_13907,N_13804);
or U13978 (N_13978,N_13858,N_13853);
nor U13979 (N_13979,N_13842,N_13813);
nor U13980 (N_13980,N_13843,N_13822);
nor U13981 (N_13981,N_13786,N_13811);
nor U13982 (N_13982,N_13911,N_13855);
nand U13983 (N_13983,N_13908,N_13803);
or U13984 (N_13984,N_13880,N_13826);
or U13985 (N_13985,N_13850,N_13919);
and U13986 (N_13986,N_13791,N_13863);
or U13987 (N_13987,N_13831,N_13844);
or U13988 (N_13988,N_13876,N_13901);
xor U13989 (N_13989,N_13837,N_13899);
nand U13990 (N_13990,N_13821,N_13810);
or U13991 (N_13991,N_13820,N_13868);
or U13992 (N_13992,N_13896,N_13792);
nor U13993 (N_13993,N_13862,N_13900);
or U13994 (N_13994,N_13879,N_13770);
and U13995 (N_13995,N_13918,N_13793);
nand U13996 (N_13996,N_13816,N_13782);
xor U13997 (N_13997,N_13773,N_13874);
nor U13998 (N_13998,N_13823,N_13827);
and U13999 (N_13999,N_13888,N_13875);
nand U14000 (N_14000,N_13829,N_13813);
nor U14001 (N_14001,N_13849,N_13776);
and U14002 (N_14002,N_13834,N_13795);
and U14003 (N_14003,N_13858,N_13786);
or U14004 (N_14004,N_13820,N_13796);
nor U14005 (N_14005,N_13801,N_13916);
or U14006 (N_14006,N_13809,N_13877);
nor U14007 (N_14007,N_13772,N_13873);
or U14008 (N_14008,N_13797,N_13843);
xnor U14009 (N_14009,N_13860,N_13761);
and U14010 (N_14010,N_13800,N_13871);
or U14011 (N_14011,N_13868,N_13888);
nor U14012 (N_14012,N_13809,N_13847);
nand U14013 (N_14013,N_13918,N_13863);
nor U14014 (N_14014,N_13770,N_13878);
nor U14015 (N_14015,N_13820,N_13909);
or U14016 (N_14016,N_13905,N_13912);
xnor U14017 (N_14017,N_13809,N_13780);
nand U14018 (N_14018,N_13770,N_13781);
nor U14019 (N_14019,N_13823,N_13773);
nor U14020 (N_14020,N_13843,N_13826);
nor U14021 (N_14021,N_13795,N_13874);
or U14022 (N_14022,N_13838,N_13909);
or U14023 (N_14023,N_13883,N_13853);
and U14024 (N_14024,N_13913,N_13883);
or U14025 (N_14025,N_13866,N_13834);
nand U14026 (N_14026,N_13844,N_13797);
and U14027 (N_14027,N_13886,N_13883);
nand U14028 (N_14028,N_13915,N_13824);
nor U14029 (N_14029,N_13877,N_13864);
nor U14030 (N_14030,N_13837,N_13810);
or U14031 (N_14031,N_13898,N_13813);
xnor U14032 (N_14032,N_13838,N_13825);
nor U14033 (N_14033,N_13819,N_13880);
nand U14034 (N_14034,N_13861,N_13775);
or U14035 (N_14035,N_13875,N_13866);
or U14036 (N_14036,N_13832,N_13915);
xor U14037 (N_14037,N_13906,N_13831);
xnor U14038 (N_14038,N_13835,N_13896);
or U14039 (N_14039,N_13812,N_13822);
and U14040 (N_14040,N_13802,N_13790);
or U14041 (N_14041,N_13808,N_13807);
or U14042 (N_14042,N_13835,N_13819);
nand U14043 (N_14043,N_13871,N_13900);
and U14044 (N_14044,N_13823,N_13822);
or U14045 (N_14045,N_13832,N_13815);
xor U14046 (N_14046,N_13773,N_13911);
and U14047 (N_14047,N_13874,N_13872);
nand U14048 (N_14048,N_13781,N_13871);
and U14049 (N_14049,N_13837,N_13828);
nand U14050 (N_14050,N_13913,N_13843);
or U14051 (N_14051,N_13764,N_13808);
nor U14052 (N_14052,N_13832,N_13770);
or U14053 (N_14053,N_13804,N_13918);
and U14054 (N_14054,N_13795,N_13814);
nor U14055 (N_14055,N_13872,N_13873);
nor U14056 (N_14056,N_13833,N_13823);
nand U14057 (N_14057,N_13792,N_13778);
nand U14058 (N_14058,N_13779,N_13821);
nand U14059 (N_14059,N_13787,N_13867);
xor U14060 (N_14060,N_13805,N_13827);
nor U14061 (N_14061,N_13874,N_13856);
xor U14062 (N_14062,N_13790,N_13761);
nand U14063 (N_14063,N_13787,N_13863);
xor U14064 (N_14064,N_13906,N_13870);
xnor U14065 (N_14065,N_13821,N_13898);
xor U14066 (N_14066,N_13795,N_13885);
nor U14067 (N_14067,N_13893,N_13888);
or U14068 (N_14068,N_13860,N_13914);
xor U14069 (N_14069,N_13841,N_13822);
or U14070 (N_14070,N_13859,N_13915);
xnor U14071 (N_14071,N_13905,N_13910);
xnor U14072 (N_14072,N_13881,N_13879);
nor U14073 (N_14073,N_13769,N_13805);
and U14074 (N_14074,N_13888,N_13820);
xnor U14075 (N_14075,N_13883,N_13859);
nand U14076 (N_14076,N_13898,N_13764);
and U14077 (N_14077,N_13798,N_13849);
nor U14078 (N_14078,N_13874,N_13842);
xor U14079 (N_14079,N_13806,N_13917);
xor U14080 (N_14080,N_14069,N_14037);
nand U14081 (N_14081,N_13999,N_14065);
nor U14082 (N_14082,N_14030,N_13963);
nand U14083 (N_14083,N_13983,N_14054);
nor U14084 (N_14084,N_13953,N_13939);
nor U14085 (N_14085,N_13989,N_14060);
xnor U14086 (N_14086,N_13940,N_14053);
or U14087 (N_14087,N_13938,N_13952);
xor U14088 (N_14088,N_13945,N_13948);
or U14089 (N_14089,N_14041,N_13970);
and U14090 (N_14090,N_13976,N_14006);
or U14091 (N_14091,N_13974,N_14018);
nand U14092 (N_14092,N_14062,N_14023);
nor U14093 (N_14093,N_14040,N_13922);
nand U14094 (N_14094,N_13987,N_14033);
or U14095 (N_14095,N_13931,N_14002);
nor U14096 (N_14096,N_13977,N_13942);
nor U14097 (N_14097,N_14070,N_13930);
nand U14098 (N_14098,N_14077,N_13975);
or U14099 (N_14099,N_13933,N_14051);
nor U14100 (N_14100,N_13965,N_13980);
and U14101 (N_14101,N_13962,N_14059);
xnor U14102 (N_14102,N_14003,N_13928);
nand U14103 (N_14103,N_14057,N_13950);
or U14104 (N_14104,N_13972,N_13926);
nand U14105 (N_14105,N_14019,N_14067);
and U14106 (N_14106,N_13927,N_14031);
nand U14107 (N_14107,N_13992,N_13979);
xnor U14108 (N_14108,N_14049,N_13969);
nor U14109 (N_14109,N_13967,N_14008);
and U14110 (N_14110,N_13964,N_13921);
and U14111 (N_14111,N_14029,N_13986);
xor U14112 (N_14112,N_13978,N_13929);
nand U14113 (N_14113,N_13958,N_14048);
or U14114 (N_14114,N_13995,N_14079);
and U14115 (N_14115,N_14052,N_13985);
and U14116 (N_14116,N_14038,N_13946);
xor U14117 (N_14117,N_14055,N_13971);
nand U14118 (N_14118,N_13924,N_14072);
xnor U14119 (N_14119,N_13981,N_13955);
or U14120 (N_14120,N_13949,N_13968);
and U14121 (N_14121,N_14000,N_14021);
nor U14122 (N_14122,N_13988,N_13943);
or U14123 (N_14123,N_14043,N_14005);
nor U14124 (N_14124,N_13997,N_14013);
or U14125 (N_14125,N_14016,N_13973);
and U14126 (N_14126,N_14056,N_13920);
and U14127 (N_14127,N_14007,N_14004);
or U14128 (N_14128,N_13996,N_14073);
nor U14129 (N_14129,N_13984,N_13935);
xor U14130 (N_14130,N_13961,N_14022);
nor U14131 (N_14131,N_13991,N_13959);
or U14132 (N_14132,N_14044,N_14064);
nand U14133 (N_14133,N_13994,N_14061);
nor U14134 (N_14134,N_14034,N_14035);
xor U14135 (N_14135,N_14050,N_13954);
nor U14136 (N_14136,N_14074,N_14015);
and U14137 (N_14137,N_14001,N_13966);
or U14138 (N_14138,N_13998,N_14027);
or U14139 (N_14139,N_14068,N_13957);
nor U14140 (N_14140,N_14076,N_14047);
nand U14141 (N_14141,N_14028,N_14032);
and U14142 (N_14142,N_14066,N_14011);
xor U14143 (N_14143,N_14063,N_14039);
and U14144 (N_14144,N_14058,N_14017);
nor U14145 (N_14145,N_13956,N_13951);
or U14146 (N_14146,N_14036,N_13944);
nand U14147 (N_14147,N_13932,N_13925);
nor U14148 (N_14148,N_14010,N_14046);
and U14149 (N_14149,N_14025,N_14071);
xnor U14150 (N_14150,N_14042,N_13941);
and U14151 (N_14151,N_13937,N_14012);
or U14152 (N_14152,N_14078,N_14014);
xor U14153 (N_14153,N_14045,N_13982);
nor U14154 (N_14154,N_13990,N_14009);
nand U14155 (N_14155,N_13960,N_14024);
or U14156 (N_14156,N_13934,N_13947);
and U14157 (N_14157,N_14075,N_13936);
or U14158 (N_14158,N_13923,N_13993);
xnor U14159 (N_14159,N_14026,N_14020);
nand U14160 (N_14160,N_13980,N_14041);
nor U14161 (N_14161,N_14077,N_14020);
or U14162 (N_14162,N_13965,N_13956);
nand U14163 (N_14163,N_13985,N_13933);
or U14164 (N_14164,N_14046,N_13923);
and U14165 (N_14165,N_13938,N_14006);
nand U14166 (N_14166,N_13924,N_13935);
nor U14167 (N_14167,N_14009,N_14046);
or U14168 (N_14168,N_14016,N_14025);
or U14169 (N_14169,N_14050,N_13944);
xnor U14170 (N_14170,N_13956,N_13989);
nor U14171 (N_14171,N_13944,N_14005);
or U14172 (N_14172,N_14050,N_13986);
and U14173 (N_14173,N_13943,N_14074);
xor U14174 (N_14174,N_13980,N_14055);
and U14175 (N_14175,N_14047,N_13941);
nand U14176 (N_14176,N_14037,N_13937);
nand U14177 (N_14177,N_14058,N_13968);
or U14178 (N_14178,N_13984,N_14017);
and U14179 (N_14179,N_13949,N_13976);
nand U14180 (N_14180,N_13940,N_14040);
or U14181 (N_14181,N_13941,N_14023);
or U14182 (N_14182,N_13928,N_14011);
nand U14183 (N_14183,N_13980,N_14053);
nor U14184 (N_14184,N_13921,N_13985);
nor U14185 (N_14185,N_13975,N_14003);
and U14186 (N_14186,N_14058,N_13936);
and U14187 (N_14187,N_14035,N_14007);
xnor U14188 (N_14188,N_13991,N_14058);
nor U14189 (N_14189,N_13935,N_14006);
nand U14190 (N_14190,N_14030,N_14000);
nand U14191 (N_14191,N_14021,N_13998);
nand U14192 (N_14192,N_13943,N_14039);
and U14193 (N_14193,N_14009,N_13934);
and U14194 (N_14194,N_14052,N_13931);
nor U14195 (N_14195,N_13944,N_13951);
xor U14196 (N_14196,N_14063,N_14060);
nor U14197 (N_14197,N_14003,N_13931);
nor U14198 (N_14198,N_13927,N_13934);
or U14199 (N_14199,N_13939,N_14000);
and U14200 (N_14200,N_14034,N_13942);
nand U14201 (N_14201,N_13922,N_13938);
xor U14202 (N_14202,N_14078,N_14073);
nor U14203 (N_14203,N_13921,N_14020);
and U14204 (N_14204,N_14064,N_13979);
and U14205 (N_14205,N_14023,N_13951);
and U14206 (N_14206,N_14033,N_13935);
or U14207 (N_14207,N_14058,N_13967);
or U14208 (N_14208,N_13921,N_13994);
nor U14209 (N_14209,N_14078,N_14001);
or U14210 (N_14210,N_14043,N_13968);
xnor U14211 (N_14211,N_14017,N_14043);
nor U14212 (N_14212,N_13972,N_14073);
nor U14213 (N_14213,N_14010,N_13960);
xor U14214 (N_14214,N_14065,N_14002);
nor U14215 (N_14215,N_14075,N_13968);
or U14216 (N_14216,N_13955,N_13934);
and U14217 (N_14217,N_13961,N_13996);
nand U14218 (N_14218,N_13999,N_14059);
or U14219 (N_14219,N_13951,N_14037);
xor U14220 (N_14220,N_13941,N_13944);
nor U14221 (N_14221,N_13953,N_14018);
or U14222 (N_14222,N_14026,N_13932);
nand U14223 (N_14223,N_14055,N_14029);
xor U14224 (N_14224,N_13949,N_13969);
or U14225 (N_14225,N_13989,N_13972);
nor U14226 (N_14226,N_14068,N_14038);
nor U14227 (N_14227,N_14063,N_13957);
xor U14228 (N_14228,N_14074,N_13978);
or U14229 (N_14229,N_13936,N_14048);
nand U14230 (N_14230,N_14053,N_13967);
nand U14231 (N_14231,N_13940,N_14028);
and U14232 (N_14232,N_13941,N_13934);
xor U14233 (N_14233,N_14026,N_13990);
or U14234 (N_14234,N_13956,N_14005);
nand U14235 (N_14235,N_13948,N_14051);
nand U14236 (N_14236,N_14007,N_14011);
or U14237 (N_14237,N_13953,N_13978);
and U14238 (N_14238,N_14039,N_13981);
and U14239 (N_14239,N_14046,N_13925);
xnor U14240 (N_14240,N_14198,N_14168);
xnor U14241 (N_14241,N_14227,N_14203);
nor U14242 (N_14242,N_14229,N_14143);
xnor U14243 (N_14243,N_14189,N_14104);
nand U14244 (N_14244,N_14127,N_14144);
nand U14245 (N_14245,N_14163,N_14138);
nand U14246 (N_14246,N_14132,N_14207);
or U14247 (N_14247,N_14134,N_14233);
and U14248 (N_14248,N_14215,N_14235);
xor U14249 (N_14249,N_14108,N_14112);
and U14250 (N_14250,N_14224,N_14161);
nor U14251 (N_14251,N_14188,N_14223);
xnor U14252 (N_14252,N_14171,N_14094);
nand U14253 (N_14253,N_14085,N_14210);
nor U14254 (N_14254,N_14157,N_14120);
nand U14255 (N_14255,N_14200,N_14169);
and U14256 (N_14256,N_14084,N_14220);
nor U14257 (N_14257,N_14178,N_14238);
or U14258 (N_14258,N_14147,N_14125);
and U14259 (N_14259,N_14121,N_14231);
xor U14260 (N_14260,N_14133,N_14192);
or U14261 (N_14261,N_14098,N_14096);
and U14262 (N_14262,N_14237,N_14119);
xnor U14263 (N_14263,N_14150,N_14184);
or U14264 (N_14264,N_14088,N_14142);
nand U14265 (N_14265,N_14141,N_14151);
xnor U14266 (N_14266,N_14175,N_14089);
xnor U14267 (N_14267,N_14149,N_14211);
or U14268 (N_14268,N_14232,N_14239);
nor U14269 (N_14269,N_14199,N_14204);
nand U14270 (N_14270,N_14162,N_14128);
or U14271 (N_14271,N_14201,N_14106);
or U14272 (N_14272,N_14086,N_14214);
xor U14273 (N_14273,N_14187,N_14131);
xnor U14274 (N_14274,N_14115,N_14217);
xor U14275 (N_14275,N_14156,N_14190);
xor U14276 (N_14276,N_14109,N_14110);
nor U14277 (N_14277,N_14111,N_14228);
nor U14278 (N_14278,N_14212,N_14221);
xnor U14279 (N_14279,N_14202,N_14166);
nor U14280 (N_14280,N_14116,N_14183);
or U14281 (N_14281,N_14124,N_14170);
nand U14282 (N_14282,N_14087,N_14126);
nand U14283 (N_14283,N_14090,N_14103);
nor U14284 (N_14284,N_14185,N_14130);
and U14285 (N_14285,N_14135,N_14219);
nor U14286 (N_14286,N_14099,N_14176);
and U14287 (N_14287,N_14146,N_14172);
nor U14288 (N_14288,N_14165,N_14180);
nand U14289 (N_14289,N_14083,N_14145);
nand U14290 (N_14290,N_14186,N_14136);
nand U14291 (N_14291,N_14177,N_14164);
or U14292 (N_14292,N_14118,N_14154);
and U14293 (N_14293,N_14191,N_14195);
nor U14294 (N_14294,N_14174,N_14082);
nand U14295 (N_14295,N_14206,N_14091);
xor U14296 (N_14296,N_14148,N_14114);
and U14297 (N_14297,N_14205,N_14105);
nor U14298 (N_14298,N_14117,N_14225);
nor U14299 (N_14299,N_14234,N_14100);
and U14300 (N_14300,N_14095,N_14222);
or U14301 (N_14301,N_14159,N_14194);
nor U14302 (N_14302,N_14140,N_14216);
nand U14303 (N_14303,N_14152,N_14129);
nor U14304 (N_14304,N_14139,N_14101);
or U14305 (N_14305,N_14193,N_14208);
nand U14306 (N_14306,N_14160,N_14113);
xnor U14307 (N_14307,N_14179,N_14167);
nor U14308 (N_14308,N_14081,N_14213);
and U14309 (N_14309,N_14230,N_14102);
or U14310 (N_14310,N_14123,N_14196);
or U14311 (N_14311,N_14155,N_14092);
xnor U14312 (N_14312,N_14182,N_14236);
or U14313 (N_14313,N_14173,N_14097);
or U14314 (N_14314,N_14153,N_14080);
xor U14315 (N_14315,N_14226,N_14158);
nor U14316 (N_14316,N_14137,N_14197);
or U14317 (N_14317,N_14093,N_14181);
nand U14318 (N_14318,N_14218,N_14122);
xor U14319 (N_14319,N_14209,N_14107);
nand U14320 (N_14320,N_14096,N_14128);
and U14321 (N_14321,N_14089,N_14087);
and U14322 (N_14322,N_14190,N_14140);
and U14323 (N_14323,N_14119,N_14098);
nand U14324 (N_14324,N_14234,N_14167);
nor U14325 (N_14325,N_14151,N_14127);
nor U14326 (N_14326,N_14138,N_14127);
nor U14327 (N_14327,N_14101,N_14160);
nor U14328 (N_14328,N_14173,N_14147);
and U14329 (N_14329,N_14144,N_14155);
or U14330 (N_14330,N_14208,N_14162);
xnor U14331 (N_14331,N_14161,N_14217);
xor U14332 (N_14332,N_14102,N_14136);
and U14333 (N_14333,N_14154,N_14185);
nor U14334 (N_14334,N_14201,N_14108);
nor U14335 (N_14335,N_14207,N_14203);
nor U14336 (N_14336,N_14234,N_14182);
xnor U14337 (N_14337,N_14165,N_14104);
nand U14338 (N_14338,N_14131,N_14104);
nand U14339 (N_14339,N_14231,N_14156);
nor U14340 (N_14340,N_14105,N_14183);
xnor U14341 (N_14341,N_14171,N_14198);
or U14342 (N_14342,N_14220,N_14162);
xor U14343 (N_14343,N_14138,N_14232);
xnor U14344 (N_14344,N_14204,N_14128);
and U14345 (N_14345,N_14151,N_14139);
or U14346 (N_14346,N_14125,N_14239);
nor U14347 (N_14347,N_14217,N_14193);
and U14348 (N_14348,N_14096,N_14169);
xnor U14349 (N_14349,N_14099,N_14175);
nand U14350 (N_14350,N_14183,N_14126);
or U14351 (N_14351,N_14155,N_14172);
xnor U14352 (N_14352,N_14144,N_14224);
or U14353 (N_14353,N_14100,N_14189);
nor U14354 (N_14354,N_14200,N_14090);
or U14355 (N_14355,N_14236,N_14238);
xor U14356 (N_14356,N_14195,N_14093);
and U14357 (N_14357,N_14237,N_14081);
nand U14358 (N_14358,N_14205,N_14090);
and U14359 (N_14359,N_14117,N_14183);
nand U14360 (N_14360,N_14110,N_14137);
or U14361 (N_14361,N_14123,N_14184);
nor U14362 (N_14362,N_14190,N_14139);
xnor U14363 (N_14363,N_14133,N_14083);
or U14364 (N_14364,N_14086,N_14131);
xor U14365 (N_14365,N_14198,N_14159);
nand U14366 (N_14366,N_14199,N_14130);
nor U14367 (N_14367,N_14147,N_14171);
nor U14368 (N_14368,N_14185,N_14158);
xor U14369 (N_14369,N_14094,N_14160);
or U14370 (N_14370,N_14219,N_14194);
or U14371 (N_14371,N_14122,N_14111);
nor U14372 (N_14372,N_14236,N_14189);
nand U14373 (N_14373,N_14208,N_14232);
or U14374 (N_14374,N_14135,N_14194);
and U14375 (N_14375,N_14217,N_14132);
nor U14376 (N_14376,N_14215,N_14176);
xnor U14377 (N_14377,N_14145,N_14147);
nand U14378 (N_14378,N_14234,N_14142);
xnor U14379 (N_14379,N_14096,N_14147);
and U14380 (N_14380,N_14110,N_14090);
or U14381 (N_14381,N_14107,N_14186);
nor U14382 (N_14382,N_14198,N_14136);
and U14383 (N_14383,N_14236,N_14084);
nor U14384 (N_14384,N_14199,N_14146);
nand U14385 (N_14385,N_14184,N_14154);
and U14386 (N_14386,N_14187,N_14162);
nor U14387 (N_14387,N_14194,N_14230);
or U14388 (N_14388,N_14139,N_14199);
nor U14389 (N_14389,N_14229,N_14129);
xor U14390 (N_14390,N_14128,N_14207);
nand U14391 (N_14391,N_14219,N_14191);
xnor U14392 (N_14392,N_14142,N_14193);
xor U14393 (N_14393,N_14197,N_14125);
nand U14394 (N_14394,N_14160,N_14193);
or U14395 (N_14395,N_14082,N_14084);
and U14396 (N_14396,N_14212,N_14136);
nor U14397 (N_14397,N_14204,N_14110);
or U14398 (N_14398,N_14187,N_14133);
nand U14399 (N_14399,N_14081,N_14088);
nand U14400 (N_14400,N_14246,N_14276);
nand U14401 (N_14401,N_14335,N_14343);
nor U14402 (N_14402,N_14325,N_14322);
nor U14403 (N_14403,N_14347,N_14350);
and U14404 (N_14404,N_14262,N_14281);
nor U14405 (N_14405,N_14249,N_14328);
nor U14406 (N_14406,N_14360,N_14336);
or U14407 (N_14407,N_14379,N_14386);
nor U14408 (N_14408,N_14363,N_14300);
nor U14409 (N_14409,N_14345,N_14331);
nand U14410 (N_14410,N_14398,N_14310);
xor U14411 (N_14411,N_14308,N_14355);
nand U14412 (N_14412,N_14356,N_14301);
and U14413 (N_14413,N_14318,N_14351);
nor U14414 (N_14414,N_14260,N_14326);
and U14415 (N_14415,N_14334,N_14275);
and U14416 (N_14416,N_14383,N_14270);
xor U14417 (N_14417,N_14307,N_14394);
nor U14418 (N_14418,N_14259,N_14257);
nand U14419 (N_14419,N_14380,N_14302);
xor U14420 (N_14420,N_14365,N_14397);
nand U14421 (N_14421,N_14309,N_14327);
or U14422 (N_14422,N_14287,N_14255);
nand U14423 (N_14423,N_14278,N_14254);
or U14424 (N_14424,N_14315,N_14264);
nor U14425 (N_14425,N_14251,N_14253);
or U14426 (N_14426,N_14361,N_14248);
and U14427 (N_14427,N_14242,N_14273);
and U14428 (N_14428,N_14298,N_14339);
nand U14429 (N_14429,N_14277,N_14258);
and U14430 (N_14430,N_14294,N_14368);
and U14431 (N_14431,N_14284,N_14387);
nand U14432 (N_14432,N_14241,N_14311);
and U14433 (N_14433,N_14381,N_14352);
or U14434 (N_14434,N_14297,N_14319);
nor U14435 (N_14435,N_14372,N_14268);
xnor U14436 (N_14436,N_14324,N_14385);
or U14437 (N_14437,N_14330,N_14369);
nand U14438 (N_14438,N_14342,N_14265);
or U14439 (N_14439,N_14269,N_14299);
or U14440 (N_14440,N_14382,N_14354);
or U14441 (N_14441,N_14395,N_14333);
nand U14442 (N_14442,N_14295,N_14286);
and U14443 (N_14443,N_14272,N_14340);
and U14444 (N_14444,N_14312,N_14353);
nor U14445 (N_14445,N_14375,N_14390);
and U14446 (N_14446,N_14250,N_14341);
nand U14447 (N_14447,N_14285,N_14282);
nor U14448 (N_14448,N_14263,N_14370);
and U14449 (N_14449,N_14261,N_14267);
or U14450 (N_14450,N_14289,N_14303);
xor U14451 (N_14451,N_14374,N_14377);
or U14452 (N_14452,N_14274,N_14316);
xnor U14453 (N_14453,N_14366,N_14367);
xnor U14454 (N_14454,N_14256,N_14384);
or U14455 (N_14455,N_14329,N_14349);
nand U14456 (N_14456,N_14346,N_14371);
and U14457 (N_14457,N_14288,N_14338);
nor U14458 (N_14458,N_14362,N_14323);
nand U14459 (N_14459,N_14357,N_14388);
nand U14460 (N_14460,N_14320,N_14240);
xnor U14461 (N_14461,N_14252,N_14376);
xor U14462 (N_14462,N_14305,N_14280);
and U14463 (N_14463,N_14244,N_14291);
or U14464 (N_14464,N_14391,N_14313);
nor U14465 (N_14465,N_14373,N_14271);
nand U14466 (N_14466,N_14243,N_14314);
and U14467 (N_14467,N_14358,N_14279);
or U14468 (N_14468,N_14266,N_14392);
nor U14469 (N_14469,N_14344,N_14292);
nor U14470 (N_14470,N_14378,N_14337);
xor U14471 (N_14471,N_14321,N_14290);
nor U14472 (N_14472,N_14399,N_14283);
nand U14473 (N_14473,N_14293,N_14317);
nor U14474 (N_14474,N_14332,N_14296);
and U14475 (N_14475,N_14396,N_14247);
or U14476 (N_14476,N_14245,N_14359);
nand U14477 (N_14477,N_14393,N_14348);
nor U14478 (N_14478,N_14306,N_14304);
and U14479 (N_14479,N_14364,N_14389);
nor U14480 (N_14480,N_14312,N_14263);
or U14481 (N_14481,N_14280,N_14263);
or U14482 (N_14482,N_14263,N_14372);
or U14483 (N_14483,N_14292,N_14297);
nor U14484 (N_14484,N_14376,N_14307);
or U14485 (N_14485,N_14278,N_14376);
and U14486 (N_14486,N_14249,N_14338);
nand U14487 (N_14487,N_14241,N_14341);
and U14488 (N_14488,N_14267,N_14366);
or U14489 (N_14489,N_14294,N_14319);
nor U14490 (N_14490,N_14313,N_14271);
or U14491 (N_14491,N_14283,N_14338);
nor U14492 (N_14492,N_14328,N_14336);
or U14493 (N_14493,N_14397,N_14359);
xnor U14494 (N_14494,N_14378,N_14338);
xnor U14495 (N_14495,N_14381,N_14262);
or U14496 (N_14496,N_14274,N_14362);
nand U14497 (N_14497,N_14346,N_14362);
or U14498 (N_14498,N_14283,N_14275);
xnor U14499 (N_14499,N_14347,N_14324);
nand U14500 (N_14500,N_14314,N_14398);
nand U14501 (N_14501,N_14357,N_14350);
nand U14502 (N_14502,N_14264,N_14277);
nand U14503 (N_14503,N_14260,N_14325);
xnor U14504 (N_14504,N_14292,N_14260);
xnor U14505 (N_14505,N_14313,N_14266);
nand U14506 (N_14506,N_14339,N_14280);
and U14507 (N_14507,N_14244,N_14243);
and U14508 (N_14508,N_14396,N_14255);
xnor U14509 (N_14509,N_14252,N_14299);
nor U14510 (N_14510,N_14322,N_14373);
or U14511 (N_14511,N_14291,N_14333);
or U14512 (N_14512,N_14314,N_14317);
or U14513 (N_14513,N_14281,N_14276);
xor U14514 (N_14514,N_14316,N_14286);
and U14515 (N_14515,N_14313,N_14338);
or U14516 (N_14516,N_14341,N_14252);
nand U14517 (N_14517,N_14297,N_14286);
nand U14518 (N_14518,N_14336,N_14388);
xor U14519 (N_14519,N_14304,N_14366);
or U14520 (N_14520,N_14309,N_14352);
nand U14521 (N_14521,N_14349,N_14398);
or U14522 (N_14522,N_14366,N_14387);
and U14523 (N_14523,N_14336,N_14297);
xor U14524 (N_14524,N_14247,N_14351);
or U14525 (N_14525,N_14361,N_14391);
or U14526 (N_14526,N_14372,N_14374);
nor U14527 (N_14527,N_14328,N_14295);
nand U14528 (N_14528,N_14295,N_14323);
or U14529 (N_14529,N_14306,N_14277);
xor U14530 (N_14530,N_14378,N_14288);
xnor U14531 (N_14531,N_14343,N_14391);
and U14532 (N_14532,N_14358,N_14302);
and U14533 (N_14533,N_14268,N_14297);
xnor U14534 (N_14534,N_14352,N_14334);
xor U14535 (N_14535,N_14358,N_14398);
nor U14536 (N_14536,N_14246,N_14286);
and U14537 (N_14537,N_14266,N_14335);
and U14538 (N_14538,N_14334,N_14369);
xor U14539 (N_14539,N_14343,N_14376);
xnor U14540 (N_14540,N_14362,N_14276);
or U14541 (N_14541,N_14324,N_14352);
nor U14542 (N_14542,N_14274,N_14302);
nor U14543 (N_14543,N_14319,N_14368);
and U14544 (N_14544,N_14310,N_14283);
and U14545 (N_14545,N_14301,N_14369);
nor U14546 (N_14546,N_14242,N_14343);
nand U14547 (N_14547,N_14290,N_14315);
and U14548 (N_14548,N_14389,N_14373);
and U14549 (N_14549,N_14248,N_14399);
xnor U14550 (N_14550,N_14307,N_14252);
xnor U14551 (N_14551,N_14350,N_14394);
and U14552 (N_14552,N_14346,N_14305);
nand U14553 (N_14553,N_14295,N_14320);
nor U14554 (N_14554,N_14309,N_14251);
xor U14555 (N_14555,N_14252,N_14284);
nand U14556 (N_14556,N_14393,N_14280);
and U14557 (N_14557,N_14381,N_14264);
and U14558 (N_14558,N_14340,N_14284);
xor U14559 (N_14559,N_14321,N_14319);
xnor U14560 (N_14560,N_14443,N_14424);
nor U14561 (N_14561,N_14402,N_14540);
nor U14562 (N_14562,N_14480,N_14481);
or U14563 (N_14563,N_14550,N_14521);
or U14564 (N_14564,N_14473,N_14477);
nand U14565 (N_14565,N_14499,N_14490);
and U14566 (N_14566,N_14418,N_14409);
nor U14567 (N_14567,N_14414,N_14432);
xnor U14568 (N_14568,N_14435,N_14539);
and U14569 (N_14569,N_14534,N_14479);
nor U14570 (N_14570,N_14447,N_14517);
nor U14571 (N_14571,N_14406,N_14448);
or U14572 (N_14572,N_14413,N_14417);
or U14573 (N_14573,N_14441,N_14536);
nand U14574 (N_14574,N_14497,N_14436);
nor U14575 (N_14575,N_14549,N_14530);
nand U14576 (N_14576,N_14466,N_14468);
nand U14577 (N_14577,N_14526,N_14469);
xor U14578 (N_14578,N_14545,N_14484);
xnor U14579 (N_14579,N_14453,N_14425);
nand U14580 (N_14580,N_14401,N_14513);
nand U14581 (N_14581,N_14488,N_14487);
nand U14582 (N_14582,N_14500,N_14518);
xnor U14583 (N_14583,N_14404,N_14444);
and U14584 (N_14584,N_14552,N_14515);
xnor U14585 (N_14585,N_14486,N_14535);
and U14586 (N_14586,N_14430,N_14554);
nor U14587 (N_14587,N_14507,N_14419);
nor U14588 (N_14588,N_14529,N_14555);
xnor U14589 (N_14589,N_14508,N_14492);
or U14590 (N_14590,N_14463,N_14504);
nor U14591 (N_14591,N_14506,N_14527);
nand U14592 (N_14592,N_14475,N_14433);
xor U14593 (N_14593,N_14405,N_14478);
nand U14594 (N_14594,N_14491,N_14464);
or U14595 (N_14595,N_14454,N_14408);
nor U14596 (N_14596,N_14450,N_14494);
nand U14597 (N_14597,N_14489,N_14411);
and U14598 (N_14598,N_14427,N_14421);
and U14599 (N_14599,N_14455,N_14531);
nand U14600 (N_14600,N_14471,N_14524);
nand U14601 (N_14601,N_14551,N_14462);
nor U14602 (N_14602,N_14416,N_14557);
xnor U14603 (N_14603,N_14451,N_14428);
nor U14604 (N_14604,N_14485,N_14474);
xnor U14605 (N_14605,N_14440,N_14556);
or U14606 (N_14606,N_14544,N_14403);
or U14607 (N_14607,N_14525,N_14519);
nand U14608 (N_14608,N_14446,N_14548);
nand U14609 (N_14609,N_14512,N_14482);
nand U14610 (N_14610,N_14547,N_14431);
nor U14611 (N_14611,N_14410,N_14472);
nor U14612 (N_14612,N_14538,N_14467);
xor U14613 (N_14613,N_14493,N_14498);
nand U14614 (N_14614,N_14407,N_14422);
nand U14615 (N_14615,N_14445,N_14465);
xor U14616 (N_14616,N_14452,N_14400);
xor U14617 (N_14617,N_14434,N_14426);
xnor U14618 (N_14618,N_14415,N_14546);
or U14619 (N_14619,N_14532,N_14520);
and U14620 (N_14620,N_14459,N_14509);
or U14621 (N_14621,N_14523,N_14458);
nand U14622 (N_14622,N_14495,N_14420);
nor U14623 (N_14623,N_14541,N_14514);
and U14624 (N_14624,N_14437,N_14423);
or U14625 (N_14625,N_14456,N_14522);
nand U14626 (N_14626,N_14528,N_14510);
nand U14627 (N_14627,N_14533,N_14470);
nand U14628 (N_14628,N_14439,N_14558);
and U14629 (N_14629,N_14442,N_14438);
and U14630 (N_14630,N_14543,N_14553);
or U14631 (N_14631,N_14505,N_14537);
or U14632 (N_14632,N_14516,N_14496);
nor U14633 (N_14633,N_14502,N_14476);
nand U14634 (N_14634,N_14542,N_14457);
and U14635 (N_14635,N_14511,N_14460);
nand U14636 (N_14636,N_14429,N_14461);
and U14637 (N_14637,N_14501,N_14449);
and U14638 (N_14638,N_14412,N_14483);
or U14639 (N_14639,N_14503,N_14559);
nor U14640 (N_14640,N_14506,N_14479);
or U14641 (N_14641,N_14491,N_14446);
and U14642 (N_14642,N_14546,N_14487);
and U14643 (N_14643,N_14434,N_14517);
nand U14644 (N_14644,N_14402,N_14554);
and U14645 (N_14645,N_14487,N_14513);
nor U14646 (N_14646,N_14406,N_14534);
nor U14647 (N_14647,N_14479,N_14408);
nor U14648 (N_14648,N_14535,N_14551);
nand U14649 (N_14649,N_14491,N_14410);
nor U14650 (N_14650,N_14532,N_14470);
and U14651 (N_14651,N_14518,N_14544);
or U14652 (N_14652,N_14495,N_14400);
nor U14653 (N_14653,N_14494,N_14417);
nand U14654 (N_14654,N_14469,N_14432);
nor U14655 (N_14655,N_14513,N_14478);
xor U14656 (N_14656,N_14416,N_14447);
and U14657 (N_14657,N_14435,N_14462);
and U14658 (N_14658,N_14474,N_14512);
nand U14659 (N_14659,N_14442,N_14514);
or U14660 (N_14660,N_14409,N_14543);
and U14661 (N_14661,N_14427,N_14528);
and U14662 (N_14662,N_14484,N_14468);
or U14663 (N_14663,N_14475,N_14516);
nor U14664 (N_14664,N_14472,N_14494);
or U14665 (N_14665,N_14414,N_14556);
nor U14666 (N_14666,N_14506,N_14460);
nand U14667 (N_14667,N_14425,N_14497);
nor U14668 (N_14668,N_14440,N_14545);
and U14669 (N_14669,N_14442,N_14414);
xnor U14670 (N_14670,N_14557,N_14472);
or U14671 (N_14671,N_14528,N_14403);
or U14672 (N_14672,N_14445,N_14492);
nand U14673 (N_14673,N_14485,N_14402);
nor U14674 (N_14674,N_14413,N_14477);
nor U14675 (N_14675,N_14462,N_14438);
nand U14676 (N_14676,N_14429,N_14543);
nor U14677 (N_14677,N_14495,N_14409);
and U14678 (N_14678,N_14499,N_14481);
nor U14679 (N_14679,N_14490,N_14418);
nand U14680 (N_14680,N_14528,N_14518);
or U14681 (N_14681,N_14413,N_14494);
nand U14682 (N_14682,N_14490,N_14402);
xnor U14683 (N_14683,N_14512,N_14430);
nand U14684 (N_14684,N_14532,N_14512);
or U14685 (N_14685,N_14423,N_14524);
xnor U14686 (N_14686,N_14514,N_14502);
xor U14687 (N_14687,N_14534,N_14429);
or U14688 (N_14688,N_14534,N_14530);
or U14689 (N_14689,N_14537,N_14482);
nor U14690 (N_14690,N_14549,N_14402);
or U14691 (N_14691,N_14473,N_14471);
or U14692 (N_14692,N_14414,N_14450);
or U14693 (N_14693,N_14522,N_14405);
xor U14694 (N_14694,N_14512,N_14483);
and U14695 (N_14695,N_14441,N_14466);
nand U14696 (N_14696,N_14485,N_14451);
and U14697 (N_14697,N_14436,N_14551);
nor U14698 (N_14698,N_14555,N_14524);
and U14699 (N_14699,N_14428,N_14443);
nand U14700 (N_14700,N_14526,N_14406);
xor U14701 (N_14701,N_14423,N_14473);
and U14702 (N_14702,N_14553,N_14541);
xnor U14703 (N_14703,N_14407,N_14502);
nor U14704 (N_14704,N_14455,N_14502);
or U14705 (N_14705,N_14523,N_14535);
and U14706 (N_14706,N_14449,N_14534);
nand U14707 (N_14707,N_14428,N_14515);
nand U14708 (N_14708,N_14534,N_14521);
xor U14709 (N_14709,N_14448,N_14404);
or U14710 (N_14710,N_14519,N_14459);
nand U14711 (N_14711,N_14479,N_14403);
xnor U14712 (N_14712,N_14408,N_14538);
and U14713 (N_14713,N_14519,N_14450);
xnor U14714 (N_14714,N_14481,N_14430);
xnor U14715 (N_14715,N_14464,N_14532);
xor U14716 (N_14716,N_14547,N_14413);
xor U14717 (N_14717,N_14492,N_14429);
and U14718 (N_14718,N_14512,N_14521);
and U14719 (N_14719,N_14411,N_14541);
and U14720 (N_14720,N_14630,N_14706);
or U14721 (N_14721,N_14597,N_14562);
or U14722 (N_14722,N_14578,N_14606);
or U14723 (N_14723,N_14664,N_14687);
or U14724 (N_14724,N_14698,N_14676);
or U14725 (N_14725,N_14662,N_14680);
xnor U14726 (N_14726,N_14640,N_14584);
nor U14727 (N_14727,N_14611,N_14712);
nor U14728 (N_14728,N_14691,N_14595);
nor U14729 (N_14729,N_14586,N_14697);
xnor U14730 (N_14730,N_14564,N_14689);
nor U14731 (N_14731,N_14651,N_14677);
nand U14732 (N_14732,N_14717,N_14669);
xnor U14733 (N_14733,N_14609,N_14667);
xor U14734 (N_14734,N_14695,N_14678);
xor U14735 (N_14735,N_14700,N_14693);
xnor U14736 (N_14736,N_14604,N_14598);
nand U14737 (N_14737,N_14670,N_14711);
or U14738 (N_14738,N_14590,N_14563);
nand U14739 (N_14739,N_14653,N_14599);
or U14740 (N_14740,N_14568,N_14573);
nand U14741 (N_14741,N_14569,N_14668);
or U14742 (N_14742,N_14709,N_14626);
nor U14743 (N_14743,N_14694,N_14656);
nor U14744 (N_14744,N_14631,N_14612);
or U14745 (N_14745,N_14625,N_14675);
and U14746 (N_14746,N_14605,N_14623);
nor U14747 (N_14747,N_14634,N_14657);
and U14748 (N_14748,N_14613,N_14594);
and U14749 (N_14749,N_14707,N_14663);
or U14750 (N_14750,N_14637,N_14682);
nand U14751 (N_14751,N_14692,N_14565);
or U14752 (N_14752,N_14659,N_14591);
or U14753 (N_14753,N_14660,N_14628);
nand U14754 (N_14754,N_14638,N_14618);
and U14755 (N_14755,N_14671,N_14672);
and U14756 (N_14756,N_14593,N_14635);
or U14757 (N_14757,N_14614,N_14639);
nor U14758 (N_14758,N_14703,N_14575);
and U14759 (N_14759,N_14610,N_14636);
nor U14760 (N_14760,N_14577,N_14571);
nor U14761 (N_14761,N_14632,N_14674);
nand U14762 (N_14762,N_14579,N_14716);
and U14763 (N_14763,N_14690,N_14615);
and U14764 (N_14764,N_14683,N_14650);
or U14765 (N_14765,N_14620,N_14576);
or U14766 (N_14766,N_14619,N_14686);
nand U14767 (N_14767,N_14688,N_14710);
xor U14768 (N_14768,N_14685,N_14696);
or U14769 (N_14769,N_14679,N_14681);
xnor U14770 (N_14770,N_14718,N_14572);
xor U14771 (N_14771,N_14629,N_14684);
xor U14772 (N_14772,N_14624,N_14574);
xnor U14773 (N_14773,N_14654,N_14607);
nand U14774 (N_14774,N_14647,N_14622);
or U14775 (N_14775,N_14673,N_14596);
xnor U14776 (N_14776,N_14701,N_14600);
nand U14777 (N_14777,N_14642,N_14713);
and U14778 (N_14778,N_14661,N_14648);
or U14779 (N_14779,N_14699,N_14658);
and U14780 (N_14780,N_14585,N_14602);
xnor U14781 (N_14781,N_14627,N_14592);
nor U14782 (N_14782,N_14649,N_14589);
or U14783 (N_14783,N_14580,N_14583);
or U14784 (N_14784,N_14616,N_14708);
nor U14785 (N_14785,N_14601,N_14561);
or U14786 (N_14786,N_14652,N_14646);
nor U14787 (N_14787,N_14621,N_14641);
or U14788 (N_14788,N_14567,N_14704);
nor U14789 (N_14789,N_14655,N_14582);
nand U14790 (N_14790,N_14560,N_14702);
and U14791 (N_14791,N_14719,N_14603);
and U14792 (N_14792,N_14643,N_14566);
nand U14793 (N_14793,N_14617,N_14581);
nand U14794 (N_14794,N_14588,N_14666);
xor U14795 (N_14795,N_14665,N_14645);
nand U14796 (N_14796,N_14633,N_14644);
and U14797 (N_14797,N_14715,N_14714);
xor U14798 (N_14798,N_14587,N_14705);
xor U14799 (N_14799,N_14570,N_14608);
and U14800 (N_14800,N_14672,N_14685);
nand U14801 (N_14801,N_14577,N_14569);
nor U14802 (N_14802,N_14638,N_14673);
nand U14803 (N_14803,N_14576,N_14662);
and U14804 (N_14804,N_14677,N_14615);
or U14805 (N_14805,N_14661,N_14592);
and U14806 (N_14806,N_14639,N_14586);
or U14807 (N_14807,N_14605,N_14574);
nor U14808 (N_14808,N_14674,N_14574);
nor U14809 (N_14809,N_14621,N_14685);
and U14810 (N_14810,N_14576,N_14710);
xor U14811 (N_14811,N_14608,N_14705);
or U14812 (N_14812,N_14591,N_14665);
and U14813 (N_14813,N_14692,N_14714);
xor U14814 (N_14814,N_14589,N_14632);
xor U14815 (N_14815,N_14650,N_14603);
or U14816 (N_14816,N_14667,N_14643);
nand U14817 (N_14817,N_14635,N_14703);
nor U14818 (N_14818,N_14713,N_14629);
nor U14819 (N_14819,N_14706,N_14642);
or U14820 (N_14820,N_14676,N_14678);
and U14821 (N_14821,N_14624,N_14637);
xor U14822 (N_14822,N_14669,N_14689);
xor U14823 (N_14823,N_14578,N_14691);
xor U14824 (N_14824,N_14670,N_14644);
xnor U14825 (N_14825,N_14610,N_14594);
or U14826 (N_14826,N_14576,N_14599);
nor U14827 (N_14827,N_14576,N_14650);
nand U14828 (N_14828,N_14681,N_14635);
and U14829 (N_14829,N_14568,N_14695);
or U14830 (N_14830,N_14670,N_14671);
and U14831 (N_14831,N_14589,N_14614);
xor U14832 (N_14832,N_14712,N_14718);
and U14833 (N_14833,N_14572,N_14645);
xor U14834 (N_14834,N_14691,N_14573);
nor U14835 (N_14835,N_14684,N_14689);
xnor U14836 (N_14836,N_14589,N_14620);
nand U14837 (N_14837,N_14627,N_14562);
or U14838 (N_14838,N_14590,N_14585);
nor U14839 (N_14839,N_14628,N_14642);
and U14840 (N_14840,N_14673,N_14699);
or U14841 (N_14841,N_14699,N_14562);
xor U14842 (N_14842,N_14629,N_14689);
and U14843 (N_14843,N_14590,N_14699);
nand U14844 (N_14844,N_14626,N_14576);
xnor U14845 (N_14845,N_14702,N_14579);
nor U14846 (N_14846,N_14650,N_14690);
nor U14847 (N_14847,N_14620,N_14639);
nand U14848 (N_14848,N_14647,N_14661);
and U14849 (N_14849,N_14592,N_14707);
xnor U14850 (N_14850,N_14628,N_14622);
xnor U14851 (N_14851,N_14600,N_14700);
or U14852 (N_14852,N_14693,N_14642);
xnor U14853 (N_14853,N_14568,N_14664);
nand U14854 (N_14854,N_14662,N_14632);
xor U14855 (N_14855,N_14685,N_14647);
xnor U14856 (N_14856,N_14701,N_14562);
or U14857 (N_14857,N_14598,N_14661);
and U14858 (N_14858,N_14710,N_14619);
nor U14859 (N_14859,N_14565,N_14677);
nor U14860 (N_14860,N_14642,N_14652);
xnor U14861 (N_14861,N_14681,N_14634);
and U14862 (N_14862,N_14654,N_14626);
nor U14863 (N_14863,N_14602,N_14576);
and U14864 (N_14864,N_14683,N_14663);
and U14865 (N_14865,N_14697,N_14621);
xnor U14866 (N_14866,N_14626,N_14624);
xor U14867 (N_14867,N_14689,N_14598);
xnor U14868 (N_14868,N_14641,N_14606);
nand U14869 (N_14869,N_14638,N_14690);
and U14870 (N_14870,N_14661,N_14690);
or U14871 (N_14871,N_14626,N_14653);
nand U14872 (N_14872,N_14611,N_14577);
nor U14873 (N_14873,N_14695,N_14676);
nand U14874 (N_14874,N_14704,N_14715);
and U14875 (N_14875,N_14686,N_14638);
nand U14876 (N_14876,N_14712,N_14668);
and U14877 (N_14877,N_14657,N_14716);
xnor U14878 (N_14878,N_14619,N_14579);
and U14879 (N_14879,N_14694,N_14571);
or U14880 (N_14880,N_14742,N_14748);
xnor U14881 (N_14881,N_14812,N_14763);
nor U14882 (N_14882,N_14819,N_14856);
xnor U14883 (N_14883,N_14828,N_14831);
nand U14884 (N_14884,N_14784,N_14874);
xor U14885 (N_14885,N_14849,N_14759);
and U14886 (N_14886,N_14878,N_14788);
xnor U14887 (N_14887,N_14833,N_14848);
and U14888 (N_14888,N_14838,N_14771);
nand U14889 (N_14889,N_14845,N_14794);
nor U14890 (N_14890,N_14854,N_14760);
and U14891 (N_14891,N_14769,N_14852);
nand U14892 (N_14892,N_14746,N_14775);
or U14893 (N_14893,N_14726,N_14758);
and U14894 (N_14894,N_14821,N_14737);
or U14895 (N_14895,N_14822,N_14862);
xor U14896 (N_14896,N_14750,N_14736);
nand U14897 (N_14897,N_14868,N_14827);
and U14898 (N_14898,N_14879,N_14780);
nor U14899 (N_14899,N_14738,N_14860);
xor U14900 (N_14900,N_14809,N_14813);
nand U14901 (N_14901,N_14840,N_14807);
nand U14902 (N_14902,N_14728,N_14811);
and U14903 (N_14903,N_14850,N_14839);
nand U14904 (N_14904,N_14744,N_14743);
and U14905 (N_14905,N_14815,N_14734);
or U14906 (N_14906,N_14783,N_14774);
nand U14907 (N_14907,N_14847,N_14871);
nand U14908 (N_14908,N_14859,N_14740);
nand U14909 (N_14909,N_14865,N_14835);
nand U14910 (N_14910,N_14723,N_14801);
nand U14911 (N_14911,N_14803,N_14837);
nand U14912 (N_14912,N_14732,N_14867);
and U14913 (N_14913,N_14730,N_14834);
and U14914 (N_14914,N_14781,N_14722);
and U14915 (N_14915,N_14751,N_14772);
and U14916 (N_14916,N_14802,N_14808);
or U14917 (N_14917,N_14830,N_14836);
nor U14918 (N_14918,N_14832,N_14757);
and U14919 (N_14919,N_14731,N_14786);
or U14920 (N_14920,N_14762,N_14741);
or U14921 (N_14921,N_14824,N_14825);
nand U14922 (N_14922,N_14857,N_14872);
or U14923 (N_14923,N_14804,N_14778);
nor U14924 (N_14924,N_14823,N_14761);
or U14925 (N_14925,N_14795,N_14739);
nand U14926 (N_14926,N_14843,N_14851);
nand U14927 (N_14927,N_14826,N_14805);
nor U14928 (N_14928,N_14765,N_14817);
nand U14929 (N_14929,N_14841,N_14870);
xnor U14930 (N_14930,N_14747,N_14729);
xnor U14931 (N_14931,N_14877,N_14764);
nand U14932 (N_14932,N_14855,N_14785);
or U14933 (N_14933,N_14767,N_14720);
and U14934 (N_14934,N_14721,N_14768);
nor U14935 (N_14935,N_14829,N_14770);
nor U14936 (N_14936,N_14727,N_14773);
and U14937 (N_14937,N_14755,N_14816);
nor U14938 (N_14938,N_14853,N_14864);
nor U14939 (N_14939,N_14806,N_14776);
and U14940 (N_14940,N_14793,N_14869);
nand U14941 (N_14941,N_14844,N_14745);
nor U14942 (N_14942,N_14818,N_14875);
or U14943 (N_14943,N_14766,N_14797);
nor U14944 (N_14944,N_14733,N_14790);
or U14945 (N_14945,N_14735,N_14777);
nand U14946 (N_14946,N_14752,N_14858);
xor U14947 (N_14947,N_14842,N_14754);
nand U14948 (N_14948,N_14796,N_14846);
or U14949 (N_14949,N_14753,N_14800);
or U14950 (N_14950,N_14789,N_14791);
or U14951 (N_14951,N_14787,N_14749);
xnor U14952 (N_14952,N_14873,N_14799);
nor U14953 (N_14953,N_14876,N_14779);
nor U14954 (N_14954,N_14861,N_14820);
nand U14955 (N_14955,N_14814,N_14782);
nor U14956 (N_14956,N_14724,N_14863);
and U14957 (N_14957,N_14798,N_14792);
xor U14958 (N_14958,N_14725,N_14810);
nand U14959 (N_14959,N_14756,N_14866);
or U14960 (N_14960,N_14852,N_14808);
and U14961 (N_14961,N_14845,N_14735);
and U14962 (N_14962,N_14799,N_14753);
and U14963 (N_14963,N_14730,N_14798);
or U14964 (N_14964,N_14757,N_14848);
xor U14965 (N_14965,N_14857,N_14817);
nand U14966 (N_14966,N_14735,N_14811);
or U14967 (N_14967,N_14832,N_14815);
or U14968 (N_14968,N_14767,N_14877);
or U14969 (N_14969,N_14874,N_14780);
nor U14970 (N_14970,N_14828,N_14827);
or U14971 (N_14971,N_14838,N_14855);
or U14972 (N_14972,N_14842,N_14757);
nand U14973 (N_14973,N_14810,N_14782);
or U14974 (N_14974,N_14726,N_14856);
xnor U14975 (N_14975,N_14800,N_14777);
nor U14976 (N_14976,N_14832,N_14744);
and U14977 (N_14977,N_14784,N_14849);
nor U14978 (N_14978,N_14786,N_14765);
nor U14979 (N_14979,N_14807,N_14738);
xnor U14980 (N_14980,N_14815,N_14755);
or U14981 (N_14981,N_14793,N_14850);
xor U14982 (N_14982,N_14867,N_14848);
xor U14983 (N_14983,N_14874,N_14863);
nand U14984 (N_14984,N_14760,N_14830);
xnor U14985 (N_14985,N_14753,N_14851);
xor U14986 (N_14986,N_14796,N_14818);
nor U14987 (N_14987,N_14749,N_14851);
or U14988 (N_14988,N_14876,N_14866);
xnor U14989 (N_14989,N_14781,N_14802);
nand U14990 (N_14990,N_14721,N_14864);
nand U14991 (N_14991,N_14874,N_14787);
and U14992 (N_14992,N_14729,N_14831);
or U14993 (N_14993,N_14837,N_14825);
nand U14994 (N_14994,N_14816,N_14820);
and U14995 (N_14995,N_14824,N_14753);
and U14996 (N_14996,N_14814,N_14823);
xor U14997 (N_14997,N_14778,N_14801);
or U14998 (N_14998,N_14774,N_14805);
nor U14999 (N_14999,N_14785,N_14727);
nor U15000 (N_15000,N_14807,N_14858);
or U15001 (N_15001,N_14748,N_14849);
and U15002 (N_15002,N_14749,N_14739);
xnor U15003 (N_15003,N_14732,N_14856);
and U15004 (N_15004,N_14816,N_14722);
or U15005 (N_15005,N_14878,N_14760);
and U15006 (N_15006,N_14834,N_14778);
or U15007 (N_15007,N_14796,N_14838);
and U15008 (N_15008,N_14838,N_14849);
and U15009 (N_15009,N_14849,N_14863);
nand U15010 (N_15010,N_14733,N_14844);
nand U15011 (N_15011,N_14847,N_14739);
and U15012 (N_15012,N_14833,N_14834);
and U15013 (N_15013,N_14832,N_14789);
nand U15014 (N_15014,N_14745,N_14820);
nand U15015 (N_15015,N_14841,N_14847);
xnor U15016 (N_15016,N_14738,N_14766);
xnor U15017 (N_15017,N_14846,N_14854);
xor U15018 (N_15018,N_14784,N_14846);
or U15019 (N_15019,N_14754,N_14775);
nand U15020 (N_15020,N_14785,N_14723);
nand U15021 (N_15021,N_14797,N_14763);
nand U15022 (N_15022,N_14769,N_14734);
and U15023 (N_15023,N_14821,N_14784);
xnor U15024 (N_15024,N_14762,N_14753);
or U15025 (N_15025,N_14787,N_14803);
nand U15026 (N_15026,N_14743,N_14860);
and U15027 (N_15027,N_14855,N_14815);
xnor U15028 (N_15028,N_14739,N_14724);
nand U15029 (N_15029,N_14773,N_14815);
or U15030 (N_15030,N_14725,N_14813);
nor U15031 (N_15031,N_14741,N_14834);
nand U15032 (N_15032,N_14851,N_14850);
or U15033 (N_15033,N_14816,N_14781);
nand U15034 (N_15034,N_14788,N_14805);
and U15035 (N_15035,N_14817,N_14789);
nand U15036 (N_15036,N_14868,N_14736);
xnor U15037 (N_15037,N_14774,N_14848);
nand U15038 (N_15038,N_14782,N_14752);
xnor U15039 (N_15039,N_14775,N_14734);
and U15040 (N_15040,N_15003,N_14895);
nand U15041 (N_15041,N_14919,N_14884);
and U15042 (N_15042,N_15036,N_14955);
nand U15043 (N_15043,N_14931,N_14907);
nand U15044 (N_15044,N_14950,N_15009);
or U15045 (N_15045,N_15002,N_14891);
nor U15046 (N_15046,N_14910,N_14989);
xor U15047 (N_15047,N_14984,N_14932);
and U15048 (N_15048,N_14975,N_14914);
nor U15049 (N_15049,N_15037,N_14949);
xnor U15050 (N_15050,N_15012,N_14917);
nand U15051 (N_15051,N_14925,N_14994);
and U15052 (N_15052,N_14942,N_14982);
or U15053 (N_15053,N_14896,N_14892);
nand U15054 (N_15054,N_14936,N_14908);
nor U15055 (N_15055,N_14981,N_14885);
xnor U15056 (N_15056,N_14933,N_14893);
nand U15057 (N_15057,N_14903,N_14920);
and U15058 (N_15058,N_14995,N_14913);
nor U15059 (N_15059,N_15026,N_14962);
or U15060 (N_15060,N_14963,N_14969);
xnor U15061 (N_15061,N_14901,N_15000);
xnor U15062 (N_15062,N_15004,N_14944);
nor U15063 (N_15063,N_14940,N_14945);
nor U15064 (N_15064,N_15032,N_15033);
and U15065 (N_15065,N_14946,N_14888);
or U15066 (N_15066,N_14992,N_14985);
and U15067 (N_15067,N_15005,N_14977);
nor U15068 (N_15068,N_14886,N_15023);
and U15069 (N_15069,N_14923,N_14934);
nor U15070 (N_15070,N_14998,N_14948);
and U15071 (N_15071,N_15013,N_15039);
nor U15072 (N_15072,N_14947,N_14905);
and U15073 (N_15073,N_14990,N_14909);
nand U15074 (N_15074,N_14973,N_15035);
nand U15075 (N_15075,N_14976,N_14971);
or U15076 (N_15076,N_14993,N_15028);
and U15077 (N_15077,N_14957,N_15029);
or U15078 (N_15078,N_14930,N_14960);
xnor U15079 (N_15079,N_14935,N_14883);
or U15080 (N_15080,N_14966,N_14997);
and U15081 (N_15081,N_14926,N_14978);
nor U15082 (N_15082,N_15019,N_14938);
xor U15083 (N_15083,N_14952,N_14974);
xor U15084 (N_15084,N_14999,N_15011);
nor U15085 (N_15085,N_15014,N_15031);
nor U15086 (N_15086,N_14937,N_14911);
nand U15087 (N_15087,N_14882,N_15022);
and U15088 (N_15088,N_14958,N_14970);
xnor U15089 (N_15089,N_15010,N_14956);
xor U15090 (N_15090,N_14929,N_14991);
xor U15091 (N_15091,N_15008,N_14983);
or U15092 (N_15092,N_14967,N_15020);
and U15093 (N_15093,N_14918,N_14972);
and U15094 (N_15094,N_14953,N_14939);
or U15095 (N_15095,N_14959,N_15016);
nor U15096 (N_15096,N_14902,N_15030);
xor U15097 (N_15097,N_14988,N_14887);
and U15098 (N_15098,N_14900,N_14927);
nor U15099 (N_15099,N_15017,N_14898);
or U15100 (N_15100,N_15018,N_14964);
xnor U15101 (N_15101,N_14899,N_15007);
and U15102 (N_15102,N_14965,N_14916);
or U15103 (N_15103,N_14915,N_15015);
and U15104 (N_15104,N_14889,N_14890);
xor U15105 (N_15105,N_14928,N_14922);
or U15106 (N_15106,N_14961,N_15001);
and U15107 (N_15107,N_15006,N_14979);
xor U15108 (N_15108,N_15038,N_14921);
and U15109 (N_15109,N_15025,N_14881);
nand U15110 (N_15110,N_14904,N_14894);
nand U15111 (N_15111,N_15034,N_15021);
and U15112 (N_15112,N_14897,N_14980);
or U15113 (N_15113,N_14906,N_15027);
nor U15114 (N_15114,N_14996,N_14924);
nand U15115 (N_15115,N_14968,N_14943);
and U15116 (N_15116,N_14987,N_14951);
and U15117 (N_15117,N_14880,N_14954);
and U15118 (N_15118,N_15024,N_14912);
or U15119 (N_15119,N_14986,N_14941);
and U15120 (N_15120,N_14929,N_14905);
xor U15121 (N_15121,N_15008,N_14997);
and U15122 (N_15122,N_14945,N_14906);
or U15123 (N_15123,N_14936,N_14897);
xnor U15124 (N_15124,N_14955,N_14997);
or U15125 (N_15125,N_14887,N_15020);
nand U15126 (N_15126,N_14962,N_14903);
xnor U15127 (N_15127,N_15009,N_14890);
nand U15128 (N_15128,N_14939,N_14982);
nor U15129 (N_15129,N_14943,N_14969);
and U15130 (N_15130,N_14969,N_15036);
nor U15131 (N_15131,N_14961,N_15000);
or U15132 (N_15132,N_14984,N_15022);
xor U15133 (N_15133,N_14918,N_14892);
nand U15134 (N_15134,N_14993,N_14905);
or U15135 (N_15135,N_14892,N_14960);
xor U15136 (N_15136,N_14953,N_14955);
xnor U15137 (N_15137,N_14932,N_15032);
and U15138 (N_15138,N_14910,N_15007);
nor U15139 (N_15139,N_14926,N_14967);
or U15140 (N_15140,N_14935,N_15018);
nor U15141 (N_15141,N_14917,N_15008);
xnor U15142 (N_15142,N_14902,N_14950);
xnor U15143 (N_15143,N_14894,N_14968);
and U15144 (N_15144,N_14904,N_15024);
nor U15145 (N_15145,N_14932,N_14897);
or U15146 (N_15146,N_14933,N_15025);
xnor U15147 (N_15147,N_14984,N_14902);
xnor U15148 (N_15148,N_15031,N_14943);
xnor U15149 (N_15149,N_14988,N_15000);
or U15150 (N_15150,N_14891,N_14887);
or U15151 (N_15151,N_14935,N_14976);
or U15152 (N_15152,N_15019,N_14880);
nand U15153 (N_15153,N_14948,N_15034);
or U15154 (N_15154,N_15037,N_15035);
nand U15155 (N_15155,N_15006,N_15016);
nand U15156 (N_15156,N_14905,N_15033);
nand U15157 (N_15157,N_14888,N_14927);
and U15158 (N_15158,N_14952,N_14906);
and U15159 (N_15159,N_14999,N_15006);
nor U15160 (N_15160,N_14994,N_15037);
xor U15161 (N_15161,N_14910,N_14892);
xor U15162 (N_15162,N_14918,N_15019);
or U15163 (N_15163,N_14915,N_15030);
nand U15164 (N_15164,N_14902,N_14898);
and U15165 (N_15165,N_14968,N_14932);
xnor U15166 (N_15166,N_14976,N_14947);
xor U15167 (N_15167,N_14987,N_14919);
xor U15168 (N_15168,N_14982,N_15019);
or U15169 (N_15169,N_14998,N_14984);
and U15170 (N_15170,N_15022,N_14890);
nor U15171 (N_15171,N_15012,N_14970);
or U15172 (N_15172,N_15016,N_14968);
xor U15173 (N_15173,N_15031,N_14930);
nor U15174 (N_15174,N_15012,N_15039);
nand U15175 (N_15175,N_14881,N_15032);
nor U15176 (N_15176,N_14910,N_14937);
and U15177 (N_15177,N_14987,N_14994);
nand U15178 (N_15178,N_14980,N_14947);
nor U15179 (N_15179,N_15021,N_14898);
and U15180 (N_15180,N_14898,N_14921);
nor U15181 (N_15181,N_15015,N_15008);
nand U15182 (N_15182,N_15006,N_14892);
nand U15183 (N_15183,N_14916,N_14883);
nor U15184 (N_15184,N_14919,N_15014);
and U15185 (N_15185,N_14977,N_15008);
nand U15186 (N_15186,N_15009,N_14920);
xor U15187 (N_15187,N_14880,N_15036);
xnor U15188 (N_15188,N_14942,N_14881);
and U15189 (N_15189,N_14881,N_14994);
nand U15190 (N_15190,N_14932,N_14991);
nor U15191 (N_15191,N_14988,N_15008);
xnor U15192 (N_15192,N_14938,N_15010);
xor U15193 (N_15193,N_14981,N_15036);
and U15194 (N_15194,N_14902,N_14976);
xnor U15195 (N_15195,N_14927,N_14971);
nor U15196 (N_15196,N_14905,N_14957);
and U15197 (N_15197,N_14969,N_15007);
or U15198 (N_15198,N_14904,N_14961);
xnor U15199 (N_15199,N_15032,N_14937);
xnor U15200 (N_15200,N_15077,N_15065);
xor U15201 (N_15201,N_15118,N_15047);
nand U15202 (N_15202,N_15151,N_15049);
nor U15203 (N_15203,N_15098,N_15148);
nand U15204 (N_15204,N_15193,N_15113);
xor U15205 (N_15205,N_15162,N_15119);
and U15206 (N_15206,N_15196,N_15129);
or U15207 (N_15207,N_15096,N_15104);
or U15208 (N_15208,N_15045,N_15150);
and U15209 (N_15209,N_15195,N_15176);
xor U15210 (N_15210,N_15068,N_15182);
xnor U15211 (N_15211,N_15199,N_15088);
xnor U15212 (N_15212,N_15177,N_15126);
and U15213 (N_15213,N_15120,N_15124);
nand U15214 (N_15214,N_15114,N_15108);
xor U15215 (N_15215,N_15076,N_15056);
or U15216 (N_15216,N_15084,N_15155);
and U15217 (N_15217,N_15180,N_15090);
xnor U15218 (N_15218,N_15188,N_15178);
and U15219 (N_15219,N_15189,N_15042);
nand U15220 (N_15220,N_15050,N_15044);
nand U15221 (N_15221,N_15170,N_15168);
or U15222 (N_15222,N_15112,N_15198);
and U15223 (N_15223,N_15183,N_15095);
or U15224 (N_15224,N_15145,N_15153);
nand U15225 (N_15225,N_15064,N_15190);
and U15226 (N_15226,N_15133,N_15160);
or U15227 (N_15227,N_15079,N_15191);
xor U15228 (N_15228,N_15125,N_15131);
and U15229 (N_15229,N_15138,N_15106);
and U15230 (N_15230,N_15128,N_15097);
xor U15231 (N_15231,N_15194,N_15173);
nand U15232 (N_15232,N_15179,N_15101);
or U15233 (N_15233,N_15144,N_15109);
and U15234 (N_15234,N_15091,N_15086);
nand U15235 (N_15235,N_15063,N_15083);
nor U15236 (N_15236,N_15142,N_15141);
nand U15237 (N_15237,N_15149,N_15067);
nand U15238 (N_15238,N_15048,N_15053);
nand U15239 (N_15239,N_15167,N_15174);
nand U15240 (N_15240,N_15099,N_15165);
nand U15241 (N_15241,N_15159,N_15043);
xor U15242 (N_15242,N_15181,N_15057);
nor U15243 (N_15243,N_15054,N_15105);
and U15244 (N_15244,N_15156,N_15111);
or U15245 (N_15245,N_15040,N_15081);
xor U15246 (N_15246,N_15134,N_15139);
or U15247 (N_15247,N_15061,N_15157);
nand U15248 (N_15248,N_15073,N_15116);
nor U15249 (N_15249,N_15169,N_15185);
and U15250 (N_15250,N_15192,N_15166);
or U15251 (N_15251,N_15059,N_15172);
and U15252 (N_15252,N_15152,N_15085);
xor U15253 (N_15253,N_15171,N_15135);
or U15254 (N_15254,N_15052,N_15132);
or U15255 (N_15255,N_15122,N_15158);
nor U15256 (N_15256,N_15130,N_15154);
or U15257 (N_15257,N_15074,N_15187);
or U15258 (N_15258,N_15046,N_15051);
nor U15259 (N_15259,N_15110,N_15075);
xnor U15260 (N_15260,N_15100,N_15066);
nand U15261 (N_15261,N_15058,N_15071);
or U15262 (N_15262,N_15163,N_15140);
nand U15263 (N_15263,N_15060,N_15184);
nand U15264 (N_15264,N_15186,N_15078);
or U15265 (N_15265,N_15080,N_15069);
or U15266 (N_15266,N_15055,N_15146);
xnor U15267 (N_15267,N_15175,N_15115);
nand U15268 (N_15268,N_15070,N_15121);
or U15269 (N_15269,N_15164,N_15089);
or U15270 (N_15270,N_15117,N_15197);
and U15271 (N_15271,N_15072,N_15161);
nor U15272 (N_15272,N_15137,N_15062);
nor U15273 (N_15273,N_15143,N_15123);
and U15274 (N_15274,N_15082,N_15093);
nor U15275 (N_15275,N_15102,N_15103);
nor U15276 (N_15276,N_15041,N_15087);
nor U15277 (N_15277,N_15094,N_15092);
or U15278 (N_15278,N_15127,N_15147);
or U15279 (N_15279,N_15107,N_15136);
and U15280 (N_15280,N_15127,N_15137);
and U15281 (N_15281,N_15104,N_15150);
xor U15282 (N_15282,N_15044,N_15088);
nor U15283 (N_15283,N_15125,N_15066);
nor U15284 (N_15284,N_15187,N_15145);
nor U15285 (N_15285,N_15050,N_15049);
nor U15286 (N_15286,N_15084,N_15069);
xnor U15287 (N_15287,N_15076,N_15149);
or U15288 (N_15288,N_15081,N_15101);
or U15289 (N_15289,N_15150,N_15117);
nand U15290 (N_15290,N_15075,N_15097);
or U15291 (N_15291,N_15128,N_15133);
nor U15292 (N_15292,N_15078,N_15113);
and U15293 (N_15293,N_15068,N_15066);
or U15294 (N_15294,N_15101,N_15120);
nor U15295 (N_15295,N_15072,N_15124);
nor U15296 (N_15296,N_15079,N_15046);
xor U15297 (N_15297,N_15152,N_15174);
or U15298 (N_15298,N_15115,N_15125);
or U15299 (N_15299,N_15121,N_15061);
and U15300 (N_15300,N_15114,N_15174);
or U15301 (N_15301,N_15151,N_15194);
nor U15302 (N_15302,N_15124,N_15134);
xor U15303 (N_15303,N_15129,N_15132);
nor U15304 (N_15304,N_15195,N_15159);
and U15305 (N_15305,N_15137,N_15102);
nand U15306 (N_15306,N_15194,N_15158);
nor U15307 (N_15307,N_15045,N_15176);
xnor U15308 (N_15308,N_15141,N_15199);
nor U15309 (N_15309,N_15044,N_15117);
nand U15310 (N_15310,N_15107,N_15152);
nand U15311 (N_15311,N_15120,N_15107);
nor U15312 (N_15312,N_15072,N_15097);
or U15313 (N_15313,N_15192,N_15051);
or U15314 (N_15314,N_15171,N_15078);
nand U15315 (N_15315,N_15132,N_15093);
nor U15316 (N_15316,N_15054,N_15142);
xor U15317 (N_15317,N_15190,N_15062);
or U15318 (N_15318,N_15087,N_15052);
nor U15319 (N_15319,N_15081,N_15155);
xnor U15320 (N_15320,N_15088,N_15189);
xor U15321 (N_15321,N_15115,N_15105);
or U15322 (N_15322,N_15181,N_15080);
xnor U15323 (N_15323,N_15110,N_15121);
or U15324 (N_15324,N_15161,N_15147);
xnor U15325 (N_15325,N_15156,N_15110);
and U15326 (N_15326,N_15183,N_15160);
nor U15327 (N_15327,N_15103,N_15090);
nor U15328 (N_15328,N_15102,N_15099);
nor U15329 (N_15329,N_15147,N_15143);
nand U15330 (N_15330,N_15085,N_15103);
xor U15331 (N_15331,N_15055,N_15073);
nand U15332 (N_15332,N_15113,N_15188);
nor U15333 (N_15333,N_15137,N_15096);
or U15334 (N_15334,N_15096,N_15129);
xnor U15335 (N_15335,N_15148,N_15179);
and U15336 (N_15336,N_15042,N_15085);
and U15337 (N_15337,N_15140,N_15043);
nand U15338 (N_15338,N_15093,N_15185);
and U15339 (N_15339,N_15106,N_15134);
nor U15340 (N_15340,N_15109,N_15164);
nor U15341 (N_15341,N_15136,N_15080);
nor U15342 (N_15342,N_15082,N_15063);
nor U15343 (N_15343,N_15159,N_15194);
xnor U15344 (N_15344,N_15101,N_15046);
xnor U15345 (N_15345,N_15087,N_15116);
nor U15346 (N_15346,N_15189,N_15193);
nor U15347 (N_15347,N_15134,N_15158);
xor U15348 (N_15348,N_15197,N_15113);
or U15349 (N_15349,N_15090,N_15084);
or U15350 (N_15350,N_15057,N_15101);
xor U15351 (N_15351,N_15044,N_15107);
or U15352 (N_15352,N_15100,N_15052);
nand U15353 (N_15353,N_15048,N_15154);
and U15354 (N_15354,N_15054,N_15068);
nand U15355 (N_15355,N_15069,N_15109);
xnor U15356 (N_15356,N_15061,N_15195);
xor U15357 (N_15357,N_15198,N_15157);
or U15358 (N_15358,N_15070,N_15164);
nand U15359 (N_15359,N_15186,N_15172);
and U15360 (N_15360,N_15330,N_15302);
or U15361 (N_15361,N_15288,N_15272);
nand U15362 (N_15362,N_15346,N_15203);
and U15363 (N_15363,N_15348,N_15314);
or U15364 (N_15364,N_15263,N_15331);
xnor U15365 (N_15365,N_15236,N_15262);
nand U15366 (N_15366,N_15283,N_15355);
and U15367 (N_15367,N_15258,N_15305);
xnor U15368 (N_15368,N_15353,N_15217);
nor U15369 (N_15369,N_15318,N_15220);
or U15370 (N_15370,N_15234,N_15256);
xor U15371 (N_15371,N_15252,N_15303);
nor U15372 (N_15372,N_15301,N_15257);
and U15373 (N_15373,N_15213,N_15218);
nor U15374 (N_15374,N_15357,N_15202);
nor U15375 (N_15375,N_15299,N_15259);
nand U15376 (N_15376,N_15343,N_15273);
nand U15377 (N_15377,N_15358,N_15344);
nand U15378 (N_15378,N_15322,N_15237);
or U15379 (N_15379,N_15227,N_15329);
and U15380 (N_15380,N_15292,N_15233);
nor U15381 (N_15381,N_15205,N_15327);
nand U15382 (N_15382,N_15351,N_15328);
xor U15383 (N_15383,N_15249,N_15210);
nor U15384 (N_15384,N_15287,N_15352);
xnor U15385 (N_15385,N_15266,N_15356);
nand U15386 (N_15386,N_15300,N_15267);
nand U15387 (N_15387,N_15320,N_15214);
and U15388 (N_15388,N_15223,N_15294);
xnor U15389 (N_15389,N_15245,N_15226);
xor U15390 (N_15390,N_15270,N_15333);
nor U15391 (N_15391,N_15219,N_15271);
or U15392 (N_15392,N_15354,N_15204);
xnor U15393 (N_15393,N_15228,N_15297);
nand U15394 (N_15394,N_15311,N_15250);
xnor U15395 (N_15395,N_15268,N_15286);
or U15396 (N_15396,N_15246,N_15265);
nor U15397 (N_15397,N_15221,N_15308);
xnor U15398 (N_15398,N_15274,N_15335);
nor U15399 (N_15399,N_15295,N_15285);
xor U15400 (N_15400,N_15209,N_15304);
or U15401 (N_15401,N_15281,N_15238);
nand U15402 (N_15402,N_15326,N_15342);
nand U15403 (N_15403,N_15216,N_15350);
nand U15404 (N_15404,N_15312,N_15254);
nor U15405 (N_15405,N_15278,N_15359);
xor U15406 (N_15406,N_15319,N_15201);
nor U15407 (N_15407,N_15279,N_15260);
or U15408 (N_15408,N_15289,N_15231);
xor U15409 (N_15409,N_15323,N_15232);
or U15410 (N_15410,N_15211,N_15224);
or U15411 (N_15411,N_15212,N_15282);
or U15412 (N_15412,N_15321,N_15244);
and U15413 (N_15413,N_15248,N_15307);
or U15414 (N_15414,N_15336,N_15261);
nand U15415 (N_15415,N_15277,N_15206);
and U15416 (N_15416,N_15316,N_15284);
and U15417 (N_15417,N_15317,N_15296);
nand U15418 (N_15418,N_15332,N_15290);
xnor U15419 (N_15419,N_15225,N_15208);
nor U15420 (N_15420,N_15324,N_15325);
nand U15421 (N_15421,N_15230,N_15309);
or U15422 (N_15422,N_15253,N_15347);
nand U15423 (N_15423,N_15229,N_15240);
or U15424 (N_15424,N_15241,N_15291);
nor U15425 (N_15425,N_15306,N_15349);
nor U15426 (N_15426,N_15276,N_15251);
xnor U15427 (N_15427,N_15269,N_15215);
xnor U15428 (N_15428,N_15200,N_15337);
or U15429 (N_15429,N_15345,N_15235);
xor U15430 (N_15430,N_15239,N_15280);
nand U15431 (N_15431,N_15334,N_15275);
nor U15432 (N_15432,N_15340,N_15264);
nor U15433 (N_15433,N_15338,N_15293);
nor U15434 (N_15434,N_15222,N_15341);
and U15435 (N_15435,N_15310,N_15207);
or U15436 (N_15436,N_15313,N_15255);
and U15437 (N_15437,N_15315,N_15339);
xor U15438 (N_15438,N_15247,N_15242);
and U15439 (N_15439,N_15298,N_15243);
nand U15440 (N_15440,N_15228,N_15335);
xor U15441 (N_15441,N_15243,N_15266);
and U15442 (N_15442,N_15205,N_15307);
nand U15443 (N_15443,N_15322,N_15325);
nand U15444 (N_15444,N_15203,N_15258);
nor U15445 (N_15445,N_15335,N_15230);
nand U15446 (N_15446,N_15273,N_15237);
nor U15447 (N_15447,N_15294,N_15262);
nor U15448 (N_15448,N_15336,N_15308);
nor U15449 (N_15449,N_15293,N_15278);
or U15450 (N_15450,N_15325,N_15296);
nand U15451 (N_15451,N_15208,N_15276);
or U15452 (N_15452,N_15266,N_15214);
xnor U15453 (N_15453,N_15348,N_15310);
nor U15454 (N_15454,N_15278,N_15309);
xnor U15455 (N_15455,N_15260,N_15248);
and U15456 (N_15456,N_15207,N_15215);
and U15457 (N_15457,N_15326,N_15270);
and U15458 (N_15458,N_15240,N_15280);
nand U15459 (N_15459,N_15316,N_15207);
xnor U15460 (N_15460,N_15279,N_15262);
nand U15461 (N_15461,N_15337,N_15248);
or U15462 (N_15462,N_15261,N_15285);
or U15463 (N_15463,N_15233,N_15275);
nor U15464 (N_15464,N_15359,N_15298);
or U15465 (N_15465,N_15213,N_15327);
nor U15466 (N_15466,N_15343,N_15325);
nor U15467 (N_15467,N_15305,N_15353);
and U15468 (N_15468,N_15325,N_15262);
or U15469 (N_15469,N_15250,N_15257);
or U15470 (N_15470,N_15245,N_15324);
nor U15471 (N_15471,N_15313,N_15207);
or U15472 (N_15472,N_15306,N_15303);
and U15473 (N_15473,N_15230,N_15339);
or U15474 (N_15474,N_15312,N_15310);
nor U15475 (N_15475,N_15230,N_15324);
nand U15476 (N_15476,N_15233,N_15333);
nand U15477 (N_15477,N_15242,N_15318);
nor U15478 (N_15478,N_15267,N_15284);
or U15479 (N_15479,N_15202,N_15280);
or U15480 (N_15480,N_15345,N_15323);
nand U15481 (N_15481,N_15227,N_15300);
nor U15482 (N_15482,N_15357,N_15289);
nand U15483 (N_15483,N_15292,N_15326);
xor U15484 (N_15484,N_15323,N_15245);
or U15485 (N_15485,N_15212,N_15306);
and U15486 (N_15486,N_15348,N_15315);
nor U15487 (N_15487,N_15252,N_15219);
and U15488 (N_15488,N_15264,N_15285);
nor U15489 (N_15489,N_15305,N_15324);
nor U15490 (N_15490,N_15293,N_15276);
and U15491 (N_15491,N_15247,N_15327);
or U15492 (N_15492,N_15331,N_15306);
nor U15493 (N_15493,N_15213,N_15261);
or U15494 (N_15494,N_15303,N_15313);
and U15495 (N_15495,N_15336,N_15208);
xor U15496 (N_15496,N_15204,N_15202);
or U15497 (N_15497,N_15224,N_15341);
or U15498 (N_15498,N_15201,N_15265);
nand U15499 (N_15499,N_15290,N_15334);
or U15500 (N_15500,N_15225,N_15269);
xnor U15501 (N_15501,N_15213,N_15232);
nand U15502 (N_15502,N_15273,N_15281);
nor U15503 (N_15503,N_15343,N_15268);
nor U15504 (N_15504,N_15311,N_15256);
nand U15505 (N_15505,N_15247,N_15305);
or U15506 (N_15506,N_15230,N_15310);
or U15507 (N_15507,N_15201,N_15357);
nand U15508 (N_15508,N_15345,N_15251);
or U15509 (N_15509,N_15239,N_15318);
nor U15510 (N_15510,N_15349,N_15325);
or U15511 (N_15511,N_15236,N_15238);
and U15512 (N_15512,N_15352,N_15356);
nand U15513 (N_15513,N_15310,N_15285);
xnor U15514 (N_15514,N_15266,N_15203);
or U15515 (N_15515,N_15287,N_15212);
and U15516 (N_15516,N_15204,N_15319);
and U15517 (N_15517,N_15338,N_15307);
nor U15518 (N_15518,N_15349,N_15340);
and U15519 (N_15519,N_15211,N_15336);
xnor U15520 (N_15520,N_15480,N_15508);
nor U15521 (N_15521,N_15421,N_15396);
nand U15522 (N_15522,N_15448,N_15416);
nor U15523 (N_15523,N_15436,N_15362);
and U15524 (N_15524,N_15499,N_15382);
and U15525 (N_15525,N_15517,N_15476);
nor U15526 (N_15526,N_15497,N_15397);
or U15527 (N_15527,N_15368,N_15507);
or U15528 (N_15528,N_15440,N_15371);
nor U15529 (N_15529,N_15365,N_15447);
xnor U15530 (N_15530,N_15445,N_15381);
nand U15531 (N_15531,N_15427,N_15449);
nand U15532 (N_15532,N_15474,N_15426);
xor U15533 (N_15533,N_15428,N_15363);
nand U15534 (N_15534,N_15384,N_15398);
nand U15535 (N_15535,N_15478,N_15514);
xnor U15536 (N_15536,N_15366,N_15410);
nor U15537 (N_15537,N_15404,N_15361);
and U15538 (N_15538,N_15439,N_15438);
and U15539 (N_15539,N_15360,N_15466);
or U15540 (N_15540,N_15490,N_15388);
nand U15541 (N_15541,N_15463,N_15495);
nor U15542 (N_15542,N_15377,N_15369);
xnor U15543 (N_15543,N_15393,N_15433);
xor U15544 (N_15544,N_15506,N_15511);
and U15545 (N_15545,N_15485,N_15467);
or U15546 (N_15546,N_15394,N_15457);
and U15547 (N_15547,N_15435,N_15451);
and U15548 (N_15548,N_15408,N_15479);
xor U15549 (N_15549,N_15505,N_15389);
and U15550 (N_15550,N_15450,N_15460);
nand U15551 (N_15551,N_15444,N_15489);
and U15552 (N_15552,N_15458,N_15378);
nand U15553 (N_15553,N_15415,N_15403);
nand U15554 (N_15554,N_15441,N_15446);
and U15555 (N_15555,N_15512,N_15380);
xnor U15556 (N_15556,N_15468,N_15493);
and U15557 (N_15557,N_15407,N_15477);
nand U15558 (N_15558,N_15471,N_15443);
nand U15559 (N_15559,N_15375,N_15412);
or U15560 (N_15560,N_15417,N_15425);
and U15561 (N_15561,N_15469,N_15420);
nor U15562 (N_15562,N_15364,N_15494);
nor U15563 (N_15563,N_15515,N_15395);
nand U15564 (N_15564,N_15510,N_15430);
nor U15565 (N_15565,N_15385,N_15484);
nand U15566 (N_15566,N_15486,N_15429);
nor U15567 (N_15567,N_15461,N_15372);
and U15568 (N_15568,N_15411,N_15424);
xor U15569 (N_15569,N_15481,N_15503);
nand U15570 (N_15570,N_15473,N_15423);
or U15571 (N_15571,N_15452,N_15422);
nor U15572 (N_15572,N_15376,N_15370);
nand U15573 (N_15573,N_15392,N_15431);
nor U15574 (N_15574,N_15492,N_15373);
and U15575 (N_15575,N_15519,N_15491);
nor U15576 (N_15576,N_15482,N_15367);
and U15577 (N_15577,N_15432,N_15472);
nor U15578 (N_15578,N_15516,N_15475);
nand U15579 (N_15579,N_15391,N_15509);
xor U15580 (N_15580,N_15453,N_15418);
nor U15581 (N_15581,N_15504,N_15379);
xor U15582 (N_15582,N_15399,N_15454);
nor U15583 (N_15583,N_15464,N_15434);
and U15584 (N_15584,N_15483,N_15500);
xnor U15585 (N_15585,N_15387,N_15513);
nand U15586 (N_15586,N_15413,N_15459);
and U15587 (N_15587,N_15487,N_15390);
and U15588 (N_15588,N_15386,N_15498);
nor U15589 (N_15589,N_15442,N_15462);
or U15590 (N_15590,N_15488,N_15383);
nand U15591 (N_15591,N_15502,N_15518);
nand U15592 (N_15592,N_15405,N_15465);
nand U15593 (N_15593,N_15419,N_15401);
or U15594 (N_15594,N_15409,N_15400);
nor U15595 (N_15595,N_15496,N_15501);
nor U15596 (N_15596,N_15456,N_15414);
or U15597 (N_15597,N_15402,N_15470);
or U15598 (N_15598,N_15374,N_15406);
nand U15599 (N_15599,N_15455,N_15437);
xor U15600 (N_15600,N_15423,N_15494);
nand U15601 (N_15601,N_15504,N_15441);
or U15602 (N_15602,N_15422,N_15491);
or U15603 (N_15603,N_15366,N_15501);
nor U15604 (N_15604,N_15426,N_15504);
nand U15605 (N_15605,N_15385,N_15436);
or U15606 (N_15606,N_15467,N_15415);
or U15607 (N_15607,N_15447,N_15478);
or U15608 (N_15608,N_15508,N_15512);
nor U15609 (N_15609,N_15519,N_15408);
nor U15610 (N_15610,N_15401,N_15374);
nor U15611 (N_15611,N_15365,N_15412);
and U15612 (N_15612,N_15488,N_15422);
and U15613 (N_15613,N_15367,N_15445);
nand U15614 (N_15614,N_15443,N_15394);
xor U15615 (N_15615,N_15499,N_15481);
nor U15616 (N_15616,N_15491,N_15498);
nor U15617 (N_15617,N_15477,N_15392);
and U15618 (N_15618,N_15476,N_15442);
xnor U15619 (N_15619,N_15424,N_15360);
nand U15620 (N_15620,N_15375,N_15376);
or U15621 (N_15621,N_15423,N_15382);
or U15622 (N_15622,N_15386,N_15424);
and U15623 (N_15623,N_15364,N_15443);
or U15624 (N_15624,N_15423,N_15496);
or U15625 (N_15625,N_15375,N_15425);
xnor U15626 (N_15626,N_15475,N_15491);
nor U15627 (N_15627,N_15426,N_15395);
xor U15628 (N_15628,N_15385,N_15398);
or U15629 (N_15629,N_15429,N_15405);
xnor U15630 (N_15630,N_15508,N_15478);
nand U15631 (N_15631,N_15402,N_15469);
and U15632 (N_15632,N_15516,N_15463);
nand U15633 (N_15633,N_15397,N_15404);
xor U15634 (N_15634,N_15509,N_15518);
xnor U15635 (N_15635,N_15416,N_15384);
and U15636 (N_15636,N_15494,N_15378);
xor U15637 (N_15637,N_15380,N_15372);
nor U15638 (N_15638,N_15408,N_15410);
nand U15639 (N_15639,N_15473,N_15458);
or U15640 (N_15640,N_15461,N_15441);
xor U15641 (N_15641,N_15433,N_15474);
or U15642 (N_15642,N_15419,N_15363);
nor U15643 (N_15643,N_15404,N_15380);
or U15644 (N_15644,N_15494,N_15501);
nand U15645 (N_15645,N_15419,N_15463);
nor U15646 (N_15646,N_15479,N_15429);
or U15647 (N_15647,N_15473,N_15440);
nand U15648 (N_15648,N_15484,N_15470);
and U15649 (N_15649,N_15450,N_15432);
or U15650 (N_15650,N_15518,N_15445);
nand U15651 (N_15651,N_15510,N_15450);
nor U15652 (N_15652,N_15380,N_15427);
and U15653 (N_15653,N_15519,N_15481);
nand U15654 (N_15654,N_15402,N_15446);
xor U15655 (N_15655,N_15373,N_15497);
or U15656 (N_15656,N_15450,N_15516);
and U15657 (N_15657,N_15473,N_15389);
or U15658 (N_15658,N_15393,N_15372);
and U15659 (N_15659,N_15492,N_15503);
nand U15660 (N_15660,N_15482,N_15443);
or U15661 (N_15661,N_15504,N_15416);
nand U15662 (N_15662,N_15396,N_15388);
and U15663 (N_15663,N_15496,N_15386);
or U15664 (N_15664,N_15511,N_15398);
or U15665 (N_15665,N_15398,N_15470);
and U15666 (N_15666,N_15370,N_15478);
xnor U15667 (N_15667,N_15385,N_15488);
xor U15668 (N_15668,N_15461,N_15443);
xnor U15669 (N_15669,N_15514,N_15398);
or U15670 (N_15670,N_15371,N_15417);
and U15671 (N_15671,N_15388,N_15444);
nor U15672 (N_15672,N_15519,N_15418);
nand U15673 (N_15673,N_15505,N_15403);
nand U15674 (N_15674,N_15451,N_15495);
and U15675 (N_15675,N_15379,N_15479);
and U15676 (N_15676,N_15383,N_15507);
nand U15677 (N_15677,N_15437,N_15505);
nor U15678 (N_15678,N_15384,N_15386);
and U15679 (N_15679,N_15446,N_15390);
nor U15680 (N_15680,N_15613,N_15523);
or U15681 (N_15681,N_15579,N_15664);
and U15682 (N_15682,N_15548,N_15627);
or U15683 (N_15683,N_15586,N_15526);
xnor U15684 (N_15684,N_15629,N_15666);
xnor U15685 (N_15685,N_15552,N_15520);
and U15686 (N_15686,N_15678,N_15658);
nand U15687 (N_15687,N_15542,N_15604);
nor U15688 (N_15688,N_15673,N_15618);
nand U15689 (N_15689,N_15644,N_15569);
xnor U15690 (N_15690,N_15553,N_15573);
xnor U15691 (N_15691,N_15625,N_15584);
or U15692 (N_15692,N_15608,N_15558);
nor U15693 (N_15693,N_15653,N_15530);
and U15694 (N_15694,N_15655,N_15540);
and U15695 (N_15695,N_15667,N_15631);
nor U15696 (N_15696,N_15633,N_15643);
nand U15697 (N_15697,N_15599,N_15626);
nand U15698 (N_15698,N_15525,N_15601);
nor U15699 (N_15699,N_15641,N_15669);
nor U15700 (N_15700,N_15605,N_15594);
or U15701 (N_15701,N_15535,N_15639);
and U15702 (N_15702,N_15581,N_15539);
nand U15703 (N_15703,N_15671,N_15538);
nand U15704 (N_15704,N_15621,N_15616);
nor U15705 (N_15705,N_15528,N_15521);
and U15706 (N_15706,N_15642,N_15591);
nand U15707 (N_15707,N_15566,N_15544);
or U15708 (N_15708,N_15546,N_15632);
xor U15709 (N_15709,N_15549,N_15563);
xnor U15710 (N_15710,N_15596,N_15559);
xor U15711 (N_15711,N_15531,N_15677);
or U15712 (N_15712,N_15628,N_15598);
or U15713 (N_15713,N_15668,N_15652);
nor U15714 (N_15714,N_15537,N_15676);
and U15715 (N_15715,N_15679,N_15646);
and U15716 (N_15716,N_15534,N_15555);
xor U15717 (N_15717,N_15576,N_15656);
or U15718 (N_15718,N_15600,N_15532);
or U15719 (N_15719,N_15572,N_15587);
nand U15720 (N_15720,N_15615,N_15657);
or U15721 (N_15721,N_15610,N_15557);
or U15722 (N_15722,N_15556,N_15645);
and U15723 (N_15723,N_15565,N_15662);
and U15724 (N_15724,N_15571,N_15654);
nand U15725 (N_15725,N_15589,N_15672);
nor U15726 (N_15726,N_15607,N_15578);
and U15727 (N_15727,N_15636,N_15562);
and U15728 (N_15728,N_15614,N_15536);
and U15729 (N_15729,N_15580,N_15670);
or U15730 (N_15730,N_15635,N_15606);
nand U15731 (N_15731,N_15647,N_15622);
and U15732 (N_15732,N_15612,N_15648);
nor U15733 (N_15733,N_15543,N_15663);
and U15734 (N_15734,N_15590,N_15550);
nor U15735 (N_15735,N_15529,N_15533);
or U15736 (N_15736,N_15659,N_15649);
xor U15737 (N_15737,N_15623,N_15547);
nor U15738 (N_15738,N_15597,N_15619);
and U15739 (N_15739,N_15582,N_15637);
and U15740 (N_15740,N_15551,N_15675);
or U15741 (N_15741,N_15617,N_15624);
and U15742 (N_15742,N_15592,N_15630);
nor U15743 (N_15743,N_15660,N_15609);
nand U15744 (N_15744,N_15564,N_15595);
nand U15745 (N_15745,N_15585,N_15634);
nand U15746 (N_15746,N_15575,N_15588);
or U15747 (N_15747,N_15603,N_15541);
or U15748 (N_15748,N_15651,N_15554);
and U15749 (N_15749,N_15640,N_15665);
xnor U15750 (N_15750,N_15620,N_15545);
nand U15751 (N_15751,N_15593,N_15638);
and U15752 (N_15752,N_15524,N_15583);
and U15753 (N_15753,N_15674,N_15574);
nand U15754 (N_15754,N_15650,N_15567);
and U15755 (N_15755,N_15602,N_15661);
nand U15756 (N_15756,N_15522,N_15527);
or U15757 (N_15757,N_15568,N_15577);
xor U15758 (N_15758,N_15570,N_15560);
nand U15759 (N_15759,N_15611,N_15561);
nand U15760 (N_15760,N_15552,N_15675);
nor U15761 (N_15761,N_15644,N_15572);
nor U15762 (N_15762,N_15566,N_15604);
nand U15763 (N_15763,N_15606,N_15627);
nand U15764 (N_15764,N_15633,N_15552);
nand U15765 (N_15765,N_15677,N_15569);
or U15766 (N_15766,N_15557,N_15550);
xnor U15767 (N_15767,N_15526,N_15661);
nor U15768 (N_15768,N_15601,N_15659);
nand U15769 (N_15769,N_15617,N_15620);
nor U15770 (N_15770,N_15643,N_15661);
nand U15771 (N_15771,N_15562,N_15590);
xnor U15772 (N_15772,N_15588,N_15598);
or U15773 (N_15773,N_15552,N_15539);
nor U15774 (N_15774,N_15556,N_15575);
xnor U15775 (N_15775,N_15601,N_15534);
and U15776 (N_15776,N_15532,N_15639);
nand U15777 (N_15777,N_15528,N_15549);
nand U15778 (N_15778,N_15670,N_15608);
and U15779 (N_15779,N_15565,N_15607);
xnor U15780 (N_15780,N_15609,N_15652);
or U15781 (N_15781,N_15624,N_15541);
or U15782 (N_15782,N_15542,N_15658);
xor U15783 (N_15783,N_15553,N_15653);
xor U15784 (N_15784,N_15608,N_15550);
nor U15785 (N_15785,N_15546,N_15542);
nor U15786 (N_15786,N_15553,N_15663);
nor U15787 (N_15787,N_15573,N_15543);
nor U15788 (N_15788,N_15581,N_15607);
and U15789 (N_15789,N_15580,N_15564);
or U15790 (N_15790,N_15565,N_15619);
nor U15791 (N_15791,N_15666,N_15620);
and U15792 (N_15792,N_15637,N_15555);
or U15793 (N_15793,N_15602,N_15558);
or U15794 (N_15794,N_15561,N_15575);
and U15795 (N_15795,N_15572,N_15609);
and U15796 (N_15796,N_15572,N_15522);
nor U15797 (N_15797,N_15645,N_15613);
xor U15798 (N_15798,N_15643,N_15677);
or U15799 (N_15799,N_15654,N_15634);
xor U15800 (N_15800,N_15549,N_15546);
and U15801 (N_15801,N_15663,N_15629);
nand U15802 (N_15802,N_15548,N_15552);
nand U15803 (N_15803,N_15666,N_15529);
and U15804 (N_15804,N_15634,N_15643);
nand U15805 (N_15805,N_15651,N_15674);
xor U15806 (N_15806,N_15580,N_15656);
nor U15807 (N_15807,N_15647,N_15542);
nor U15808 (N_15808,N_15573,N_15619);
nor U15809 (N_15809,N_15522,N_15622);
nand U15810 (N_15810,N_15660,N_15530);
xnor U15811 (N_15811,N_15667,N_15562);
or U15812 (N_15812,N_15608,N_15536);
xor U15813 (N_15813,N_15606,N_15672);
and U15814 (N_15814,N_15553,N_15527);
and U15815 (N_15815,N_15569,N_15596);
xnor U15816 (N_15816,N_15533,N_15610);
and U15817 (N_15817,N_15553,N_15520);
or U15818 (N_15818,N_15605,N_15643);
xnor U15819 (N_15819,N_15561,N_15554);
nor U15820 (N_15820,N_15602,N_15549);
nor U15821 (N_15821,N_15542,N_15569);
nor U15822 (N_15822,N_15652,N_15588);
nand U15823 (N_15823,N_15521,N_15663);
nor U15824 (N_15824,N_15644,N_15642);
and U15825 (N_15825,N_15575,N_15586);
nand U15826 (N_15826,N_15614,N_15628);
nand U15827 (N_15827,N_15543,N_15561);
nor U15828 (N_15828,N_15639,N_15660);
xnor U15829 (N_15829,N_15580,N_15583);
nor U15830 (N_15830,N_15578,N_15656);
nand U15831 (N_15831,N_15538,N_15582);
xor U15832 (N_15832,N_15652,N_15672);
nand U15833 (N_15833,N_15675,N_15522);
or U15834 (N_15834,N_15576,N_15520);
nor U15835 (N_15835,N_15619,N_15647);
nand U15836 (N_15836,N_15602,N_15557);
or U15837 (N_15837,N_15667,N_15655);
or U15838 (N_15838,N_15657,N_15573);
xor U15839 (N_15839,N_15659,N_15611);
nand U15840 (N_15840,N_15736,N_15821);
nand U15841 (N_15841,N_15711,N_15782);
xor U15842 (N_15842,N_15722,N_15702);
or U15843 (N_15843,N_15797,N_15683);
nand U15844 (N_15844,N_15786,N_15777);
and U15845 (N_15845,N_15775,N_15788);
xor U15846 (N_15846,N_15812,N_15822);
and U15847 (N_15847,N_15759,N_15705);
or U15848 (N_15848,N_15698,N_15749);
or U15849 (N_15849,N_15738,N_15793);
nand U15850 (N_15850,N_15817,N_15774);
and U15851 (N_15851,N_15828,N_15730);
nor U15852 (N_15852,N_15816,N_15834);
and U15853 (N_15853,N_15796,N_15684);
nand U15854 (N_15854,N_15723,N_15699);
xor U15855 (N_15855,N_15779,N_15805);
nor U15856 (N_15856,N_15742,N_15792);
xor U15857 (N_15857,N_15762,N_15745);
nand U15858 (N_15858,N_15688,N_15700);
or U15859 (N_15859,N_15696,N_15686);
xnor U15860 (N_15860,N_15740,N_15827);
or U15861 (N_15861,N_15758,N_15756);
nor U15862 (N_15862,N_15706,N_15685);
or U15863 (N_15863,N_15772,N_15743);
and U15864 (N_15864,N_15781,N_15720);
nor U15865 (N_15865,N_15728,N_15717);
or U15866 (N_15866,N_15754,N_15818);
and U15867 (N_15867,N_15704,N_15833);
or U15868 (N_15868,N_15773,N_15692);
and U15869 (N_15869,N_15731,N_15750);
and U15870 (N_15870,N_15697,N_15787);
and U15871 (N_15871,N_15824,N_15703);
xnor U15872 (N_15872,N_15733,N_15727);
nand U15873 (N_15873,N_15790,N_15721);
nor U15874 (N_15874,N_15752,N_15690);
nor U15875 (N_15875,N_15811,N_15836);
or U15876 (N_15876,N_15829,N_15729);
nor U15877 (N_15877,N_15799,N_15794);
xnor U15878 (N_15878,N_15746,N_15707);
or U15879 (N_15879,N_15785,N_15693);
and U15880 (N_15880,N_15732,N_15766);
nor U15881 (N_15881,N_15804,N_15708);
nor U15882 (N_15882,N_15783,N_15763);
nor U15883 (N_15883,N_15764,N_15769);
nor U15884 (N_15884,N_15709,N_15784);
nand U15885 (N_15885,N_15682,N_15832);
xnor U15886 (N_15886,N_15765,N_15780);
xnor U15887 (N_15887,N_15687,N_15802);
and U15888 (N_15888,N_15760,N_15809);
nand U15889 (N_15889,N_15798,N_15791);
nor U15890 (N_15890,N_15737,N_15681);
nor U15891 (N_15891,N_15748,N_15718);
nand U15892 (N_15892,N_15831,N_15753);
nand U15893 (N_15893,N_15757,N_15725);
nor U15894 (N_15894,N_15826,N_15778);
nand U15895 (N_15895,N_15815,N_15823);
or U15896 (N_15896,N_15771,N_15789);
xnor U15897 (N_15897,N_15767,N_15837);
xnor U15898 (N_15898,N_15795,N_15755);
nor U15899 (N_15899,N_15715,N_15776);
nand U15900 (N_15900,N_15710,N_15735);
nor U15901 (N_15901,N_15761,N_15830);
nor U15902 (N_15902,N_15807,N_15719);
nand U15903 (N_15903,N_15713,N_15825);
or U15904 (N_15904,N_15810,N_15751);
xor U15905 (N_15905,N_15747,N_15739);
nand U15906 (N_15906,N_15835,N_15691);
nor U15907 (N_15907,N_15689,N_15712);
xor U15908 (N_15908,N_15714,N_15695);
and U15909 (N_15909,N_15726,N_15770);
and U15910 (N_15910,N_15734,N_15680);
and U15911 (N_15911,N_15744,N_15701);
nor U15912 (N_15912,N_15694,N_15741);
nor U15913 (N_15913,N_15838,N_15724);
xor U15914 (N_15914,N_15839,N_15813);
xor U15915 (N_15915,N_15801,N_15814);
or U15916 (N_15916,N_15820,N_15800);
and U15917 (N_15917,N_15819,N_15806);
and U15918 (N_15918,N_15808,N_15716);
nor U15919 (N_15919,N_15803,N_15768);
nand U15920 (N_15920,N_15828,N_15823);
and U15921 (N_15921,N_15744,N_15834);
xnor U15922 (N_15922,N_15683,N_15733);
or U15923 (N_15923,N_15825,N_15698);
and U15924 (N_15924,N_15793,N_15726);
and U15925 (N_15925,N_15693,N_15720);
xor U15926 (N_15926,N_15820,N_15776);
xnor U15927 (N_15927,N_15780,N_15690);
nor U15928 (N_15928,N_15827,N_15707);
nand U15929 (N_15929,N_15787,N_15722);
xor U15930 (N_15930,N_15688,N_15730);
and U15931 (N_15931,N_15832,N_15800);
and U15932 (N_15932,N_15837,N_15772);
and U15933 (N_15933,N_15691,N_15722);
xnor U15934 (N_15934,N_15826,N_15791);
nand U15935 (N_15935,N_15717,N_15806);
nor U15936 (N_15936,N_15767,N_15727);
nand U15937 (N_15937,N_15681,N_15735);
nand U15938 (N_15938,N_15773,N_15785);
nand U15939 (N_15939,N_15816,N_15818);
xor U15940 (N_15940,N_15700,N_15749);
and U15941 (N_15941,N_15807,N_15729);
and U15942 (N_15942,N_15695,N_15760);
xor U15943 (N_15943,N_15814,N_15733);
xor U15944 (N_15944,N_15801,N_15818);
nand U15945 (N_15945,N_15763,N_15735);
nor U15946 (N_15946,N_15691,N_15795);
nor U15947 (N_15947,N_15740,N_15764);
nand U15948 (N_15948,N_15805,N_15793);
nand U15949 (N_15949,N_15702,N_15808);
nand U15950 (N_15950,N_15714,N_15806);
or U15951 (N_15951,N_15753,N_15807);
xnor U15952 (N_15952,N_15785,N_15834);
and U15953 (N_15953,N_15784,N_15761);
nor U15954 (N_15954,N_15811,N_15734);
and U15955 (N_15955,N_15764,N_15811);
nor U15956 (N_15956,N_15688,N_15788);
nor U15957 (N_15957,N_15789,N_15819);
or U15958 (N_15958,N_15821,N_15766);
xor U15959 (N_15959,N_15688,N_15714);
or U15960 (N_15960,N_15828,N_15819);
or U15961 (N_15961,N_15696,N_15829);
nor U15962 (N_15962,N_15799,N_15802);
or U15963 (N_15963,N_15680,N_15754);
nor U15964 (N_15964,N_15799,N_15786);
or U15965 (N_15965,N_15774,N_15719);
and U15966 (N_15966,N_15708,N_15768);
or U15967 (N_15967,N_15766,N_15782);
nand U15968 (N_15968,N_15764,N_15832);
and U15969 (N_15969,N_15721,N_15692);
or U15970 (N_15970,N_15762,N_15786);
and U15971 (N_15971,N_15759,N_15745);
and U15972 (N_15972,N_15719,N_15752);
nand U15973 (N_15973,N_15827,N_15739);
nand U15974 (N_15974,N_15789,N_15788);
nand U15975 (N_15975,N_15765,N_15738);
and U15976 (N_15976,N_15693,N_15798);
and U15977 (N_15977,N_15690,N_15702);
and U15978 (N_15978,N_15685,N_15741);
xor U15979 (N_15979,N_15729,N_15780);
xor U15980 (N_15980,N_15689,N_15754);
nor U15981 (N_15981,N_15733,N_15706);
and U15982 (N_15982,N_15764,N_15699);
and U15983 (N_15983,N_15805,N_15696);
or U15984 (N_15984,N_15698,N_15812);
nor U15985 (N_15985,N_15757,N_15785);
nand U15986 (N_15986,N_15786,N_15688);
or U15987 (N_15987,N_15697,N_15793);
and U15988 (N_15988,N_15834,N_15746);
and U15989 (N_15989,N_15723,N_15817);
xor U15990 (N_15990,N_15714,N_15792);
or U15991 (N_15991,N_15748,N_15762);
and U15992 (N_15992,N_15739,N_15706);
and U15993 (N_15993,N_15808,N_15811);
nor U15994 (N_15994,N_15752,N_15814);
nor U15995 (N_15995,N_15786,N_15726);
and U15996 (N_15996,N_15828,N_15805);
nor U15997 (N_15997,N_15778,N_15695);
nand U15998 (N_15998,N_15832,N_15831);
or U15999 (N_15999,N_15805,N_15683);
nor U16000 (N_16000,N_15995,N_15962);
or U16001 (N_16001,N_15944,N_15875);
xor U16002 (N_16002,N_15928,N_15888);
nor U16003 (N_16003,N_15881,N_15885);
nand U16004 (N_16004,N_15924,N_15952);
or U16005 (N_16005,N_15884,N_15909);
nand U16006 (N_16006,N_15900,N_15939);
nand U16007 (N_16007,N_15948,N_15898);
and U16008 (N_16008,N_15979,N_15935);
nor U16009 (N_16009,N_15883,N_15983);
and U16010 (N_16010,N_15937,N_15877);
and U16011 (N_16011,N_15990,N_15968);
nand U16012 (N_16012,N_15861,N_15874);
nand U16013 (N_16013,N_15840,N_15889);
or U16014 (N_16014,N_15986,N_15927);
and U16015 (N_16015,N_15961,N_15904);
nand U16016 (N_16016,N_15858,N_15870);
xor U16017 (N_16017,N_15926,N_15955);
nor U16018 (N_16018,N_15963,N_15940);
xnor U16019 (N_16019,N_15950,N_15908);
xnor U16020 (N_16020,N_15994,N_15906);
nor U16021 (N_16021,N_15988,N_15933);
and U16022 (N_16022,N_15993,N_15982);
or U16023 (N_16023,N_15984,N_15907);
or U16024 (N_16024,N_15911,N_15845);
and U16025 (N_16025,N_15864,N_15953);
or U16026 (N_16026,N_15880,N_15917);
or U16027 (N_16027,N_15863,N_15997);
nand U16028 (N_16028,N_15918,N_15970);
or U16029 (N_16029,N_15841,N_15854);
or U16030 (N_16030,N_15873,N_15886);
nand U16031 (N_16031,N_15949,N_15905);
or U16032 (N_16032,N_15887,N_15852);
and U16033 (N_16033,N_15947,N_15848);
or U16034 (N_16034,N_15857,N_15876);
or U16035 (N_16035,N_15922,N_15971);
xor U16036 (N_16036,N_15932,N_15882);
or U16037 (N_16037,N_15910,N_15871);
nand U16038 (N_16038,N_15936,N_15853);
and U16039 (N_16039,N_15945,N_15978);
nor U16040 (N_16040,N_15920,N_15919);
and U16041 (N_16041,N_15902,N_15903);
xnor U16042 (N_16042,N_15856,N_15980);
and U16043 (N_16043,N_15915,N_15862);
and U16044 (N_16044,N_15957,N_15956);
nor U16045 (N_16045,N_15991,N_15943);
xor U16046 (N_16046,N_15843,N_15916);
or U16047 (N_16047,N_15878,N_15895);
nand U16048 (N_16048,N_15896,N_15872);
xnor U16049 (N_16049,N_15967,N_15942);
nor U16050 (N_16050,N_15989,N_15977);
or U16051 (N_16051,N_15929,N_15844);
or U16052 (N_16052,N_15899,N_15930);
nand U16053 (N_16053,N_15869,N_15913);
xnor U16054 (N_16054,N_15923,N_15985);
nor U16055 (N_16055,N_15901,N_15891);
xnor U16056 (N_16056,N_15941,N_15859);
or U16057 (N_16057,N_15964,N_15849);
and U16058 (N_16058,N_15976,N_15879);
and U16059 (N_16059,N_15851,N_15966);
xnor U16060 (N_16060,N_15868,N_15890);
nor U16061 (N_16061,N_15972,N_15959);
nand U16062 (N_16062,N_15847,N_15998);
nand U16063 (N_16063,N_15846,N_15850);
or U16064 (N_16064,N_15975,N_15974);
nand U16065 (N_16065,N_15921,N_15934);
or U16066 (N_16066,N_15931,N_15892);
xnor U16067 (N_16067,N_15897,N_15894);
xor U16068 (N_16068,N_15965,N_15960);
or U16069 (N_16069,N_15999,N_15973);
and U16070 (N_16070,N_15996,N_15969);
nor U16071 (N_16071,N_15866,N_15914);
and U16072 (N_16072,N_15987,N_15865);
xor U16073 (N_16073,N_15867,N_15893);
nor U16074 (N_16074,N_15958,N_15946);
or U16075 (N_16075,N_15925,N_15981);
or U16076 (N_16076,N_15954,N_15912);
and U16077 (N_16077,N_15842,N_15860);
xnor U16078 (N_16078,N_15951,N_15938);
or U16079 (N_16079,N_15855,N_15992);
nor U16080 (N_16080,N_15884,N_15976);
and U16081 (N_16081,N_15905,N_15893);
and U16082 (N_16082,N_15922,N_15915);
xor U16083 (N_16083,N_15971,N_15921);
and U16084 (N_16084,N_15866,N_15870);
or U16085 (N_16085,N_15916,N_15869);
xor U16086 (N_16086,N_15913,N_15868);
nor U16087 (N_16087,N_15847,N_15918);
nand U16088 (N_16088,N_15842,N_15950);
nor U16089 (N_16089,N_15991,N_15992);
or U16090 (N_16090,N_15865,N_15988);
or U16091 (N_16091,N_15842,N_15943);
nor U16092 (N_16092,N_15932,N_15900);
or U16093 (N_16093,N_15963,N_15919);
xnor U16094 (N_16094,N_15937,N_15858);
xor U16095 (N_16095,N_15967,N_15971);
nor U16096 (N_16096,N_15885,N_15902);
or U16097 (N_16097,N_15951,N_15841);
nor U16098 (N_16098,N_15972,N_15856);
nand U16099 (N_16099,N_15863,N_15892);
xnor U16100 (N_16100,N_15871,N_15971);
xnor U16101 (N_16101,N_15949,N_15897);
xor U16102 (N_16102,N_15935,N_15932);
xnor U16103 (N_16103,N_15975,N_15970);
nand U16104 (N_16104,N_15969,N_15975);
nor U16105 (N_16105,N_15900,N_15993);
xnor U16106 (N_16106,N_15975,N_15871);
nand U16107 (N_16107,N_15925,N_15983);
xnor U16108 (N_16108,N_15856,N_15864);
nand U16109 (N_16109,N_15845,N_15982);
and U16110 (N_16110,N_15849,N_15991);
nor U16111 (N_16111,N_15949,N_15849);
xnor U16112 (N_16112,N_15897,N_15850);
nand U16113 (N_16113,N_15909,N_15922);
xnor U16114 (N_16114,N_15924,N_15966);
or U16115 (N_16115,N_15899,N_15853);
nor U16116 (N_16116,N_15994,N_15999);
nand U16117 (N_16117,N_15910,N_15920);
and U16118 (N_16118,N_15844,N_15918);
nand U16119 (N_16119,N_15997,N_15983);
nor U16120 (N_16120,N_15856,N_15892);
and U16121 (N_16121,N_15870,N_15955);
and U16122 (N_16122,N_15885,N_15876);
or U16123 (N_16123,N_15890,N_15969);
or U16124 (N_16124,N_15842,N_15926);
nor U16125 (N_16125,N_15969,N_15985);
nor U16126 (N_16126,N_15901,N_15917);
and U16127 (N_16127,N_15861,N_15923);
xor U16128 (N_16128,N_15974,N_15876);
nor U16129 (N_16129,N_15897,N_15916);
or U16130 (N_16130,N_15891,N_15873);
nor U16131 (N_16131,N_15988,N_15945);
and U16132 (N_16132,N_15926,N_15883);
xor U16133 (N_16133,N_15854,N_15869);
or U16134 (N_16134,N_15975,N_15917);
xor U16135 (N_16135,N_15852,N_15996);
or U16136 (N_16136,N_15878,N_15981);
nand U16137 (N_16137,N_15980,N_15840);
and U16138 (N_16138,N_15925,N_15896);
xor U16139 (N_16139,N_15991,N_15929);
or U16140 (N_16140,N_15943,N_15857);
and U16141 (N_16141,N_15879,N_15870);
xor U16142 (N_16142,N_15938,N_15943);
or U16143 (N_16143,N_15930,N_15978);
or U16144 (N_16144,N_15911,N_15905);
nand U16145 (N_16145,N_15995,N_15987);
and U16146 (N_16146,N_15952,N_15967);
nor U16147 (N_16147,N_15904,N_15856);
nor U16148 (N_16148,N_15888,N_15920);
xnor U16149 (N_16149,N_15958,N_15970);
and U16150 (N_16150,N_15938,N_15979);
nand U16151 (N_16151,N_15979,N_15842);
xor U16152 (N_16152,N_15844,N_15891);
and U16153 (N_16153,N_15980,N_15897);
nand U16154 (N_16154,N_15880,N_15949);
and U16155 (N_16155,N_15914,N_15952);
nand U16156 (N_16156,N_15973,N_15890);
and U16157 (N_16157,N_15937,N_15956);
nor U16158 (N_16158,N_15975,N_15840);
nand U16159 (N_16159,N_15929,N_15978);
nor U16160 (N_16160,N_16147,N_16002);
and U16161 (N_16161,N_16069,N_16048);
xor U16162 (N_16162,N_16138,N_16033);
and U16163 (N_16163,N_16018,N_16053);
nor U16164 (N_16164,N_16067,N_16117);
or U16165 (N_16165,N_16115,N_16060);
nand U16166 (N_16166,N_16128,N_16106);
and U16167 (N_16167,N_16111,N_16052);
nand U16168 (N_16168,N_16021,N_16009);
or U16169 (N_16169,N_16058,N_16133);
nor U16170 (N_16170,N_16046,N_16030);
nand U16171 (N_16171,N_16157,N_16113);
xor U16172 (N_16172,N_16050,N_16097);
and U16173 (N_16173,N_16015,N_16129);
and U16174 (N_16174,N_16061,N_16103);
and U16175 (N_16175,N_16063,N_16098);
or U16176 (N_16176,N_16076,N_16070);
and U16177 (N_16177,N_16012,N_16159);
nand U16178 (N_16178,N_16084,N_16094);
nor U16179 (N_16179,N_16123,N_16026);
nand U16180 (N_16180,N_16125,N_16145);
nor U16181 (N_16181,N_16007,N_16051);
and U16182 (N_16182,N_16055,N_16149);
or U16183 (N_16183,N_16119,N_16095);
or U16184 (N_16184,N_16116,N_16062);
xor U16185 (N_16185,N_16107,N_16132);
nand U16186 (N_16186,N_16082,N_16093);
xor U16187 (N_16187,N_16102,N_16074);
nand U16188 (N_16188,N_16150,N_16137);
nor U16189 (N_16189,N_16045,N_16153);
nor U16190 (N_16190,N_16025,N_16031);
and U16191 (N_16191,N_16014,N_16008);
or U16192 (N_16192,N_16131,N_16118);
nor U16193 (N_16193,N_16088,N_16042);
or U16194 (N_16194,N_16152,N_16081);
or U16195 (N_16195,N_16109,N_16114);
and U16196 (N_16196,N_16049,N_16037);
or U16197 (N_16197,N_16141,N_16020);
and U16198 (N_16198,N_16127,N_16100);
and U16199 (N_16199,N_16038,N_16073);
xnor U16200 (N_16200,N_16108,N_16112);
and U16201 (N_16201,N_16005,N_16003);
and U16202 (N_16202,N_16126,N_16075);
xnor U16203 (N_16203,N_16104,N_16087);
xnor U16204 (N_16204,N_16091,N_16121);
or U16205 (N_16205,N_16155,N_16077);
and U16206 (N_16206,N_16023,N_16032);
and U16207 (N_16207,N_16024,N_16022);
or U16208 (N_16208,N_16059,N_16154);
nor U16209 (N_16209,N_16146,N_16151);
nand U16210 (N_16210,N_16099,N_16143);
nor U16211 (N_16211,N_16122,N_16158);
nor U16212 (N_16212,N_16001,N_16054);
nor U16213 (N_16213,N_16096,N_16065);
xnor U16214 (N_16214,N_16034,N_16090);
xor U16215 (N_16215,N_16072,N_16019);
xnor U16216 (N_16216,N_16083,N_16057);
and U16217 (N_16217,N_16142,N_16120);
and U16218 (N_16218,N_16044,N_16004);
nand U16219 (N_16219,N_16105,N_16110);
nand U16220 (N_16220,N_16013,N_16156);
nor U16221 (N_16221,N_16039,N_16078);
xnor U16222 (N_16222,N_16043,N_16085);
nand U16223 (N_16223,N_16066,N_16080);
nor U16224 (N_16224,N_16089,N_16064);
xnor U16225 (N_16225,N_16136,N_16101);
nand U16226 (N_16226,N_16139,N_16010);
xnor U16227 (N_16227,N_16000,N_16006);
nor U16228 (N_16228,N_16040,N_16140);
and U16229 (N_16229,N_16079,N_16056);
or U16230 (N_16230,N_16086,N_16124);
and U16231 (N_16231,N_16035,N_16092);
and U16232 (N_16232,N_16071,N_16017);
and U16233 (N_16233,N_16144,N_16130);
and U16234 (N_16234,N_16134,N_16041);
and U16235 (N_16235,N_16028,N_16036);
xnor U16236 (N_16236,N_16027,N_16011);
or U16237 (N_16237,N_16029,N_16068);
xor U16238 (N_16238,N_16016,N_16135);
and U16239 (N_16239,N_16148,N_16047);
or U16240 (N_16240,N_16061,N_16028);
nand U16241 (N_16241,N_16033,N_16133);
nor U16242 (N_16242,N_16125,N_16026);
nand U16243 (N_16243,N_16026,N_16039);
or U16244 (N_16244,N_16097,N_16152);
nand U16245 (N_16245,N_16019,N_16155);
or U16246 (N_16246,N_16094,N_16000);
or U16247 (N_16247,N_16050,N_16039);
and U16248 (N_16248,N_16122,N_16097);
nor U16249 (N_16249,N_16014,N_16047);
nor U16250 (N_16250,N_16062,N_16040);
nand U16251 (N_16251,N_16073,N_16112);
or U16252 (N_16252,N_16105,N_16109);
xor U16253 (N_16253,N_16110,N_16157);
and U16254 (N_16254,N_16151,N_16075);
and U16255 (N_16255,N_16095,N_16000);
or U16256 (N_16256,N_16001,N_16056);
and U16257 (N_16257,N_16037,N_16012);
or U16258 (N_16258,N_16157,N_16011);
nand U16259 (N_16259,N_16126,N_16017);
and U16260 (N_16260,N_16085,N_16100);
nand U16261 (N_16261,N_16002,N_16127);
or U16262 (N_16262,N_16037,N_16089);
nor U16263 (N_16263,N_16131,N_16146);
nor U16264 (N_16264,N_16090,N_16025);
or U16265 (N_16265,N_16071,N_16038);
xor U16266 (N_16266,N_16076,N_16085);
xnor U16267 (N_16267,N_16122,N_16085);
nand U16268 (N_16268,N_16046,N_16098);
and U16269 (N_16269,N_16027,N_16024);
nor U16270 (N_16270,N_16124,N_16152);
xnor U16271 (N_16271,N_16075,N_16015);
xor U16272 (N_16272,N_16013,N_16159);
or U16273 (N_16273,N_16115,N_16007);
and U16274 (N_16274,N_16025,N_16083);
and U16275 (N_16275,N_16151,N_16152);
or U16276 (N_16276,N_16120,N_16001);
nor U16277 (N_16277,N_16135,N_16035);
and U16278 (N_16278,N_16157,N_16128);
nor U16279 (N_16279,N_16057,N_16151);
or U16280 (N_16280,N_16158,N_16006);
nand U16281 (N_16281,N_16098,N_16133);
xnor U16282 (N_16282,N_16064,N_16142);
and U16283 (N_16283,N_16048,N_16116);
nand U16284 (N_16284,N_16110,N_16070);
xor U16285 (N_16285,N_16117,N_16013);
and U16286 (N_16286,N_16057,N_16009);
xor U16287 (N_16287,N_16068,N_16027);
and U16288 (N_16288,N_16064,N_16023);
nand U16289 (N_16289,N_16115,N_16131);
nor U16290 (N_16290,N_16047,N_16038);
or U16291 (N_16291,N_16101,N_16048);
nand U16292 (N_16292,N_16096,N_16093);
nor U16293 (N_16293,N_16035,N_16141);
nand U16294 (N_16294,N_16142,N_16154);
and U16295 (N_16295,N_16100,N_16112);
nand U16296 (N_16296,N_16073,N_16081);
nor U16297 (N_16297,N_16096,N_16024);
and U16298 (N_16298,N_16133,N_16025);
nand U16299 (N_16299,N_16038,N_16143);
and U16300 (N_16300,N_16051,N_16127);
nor U16301 (N_16301,N_16138,N_16037);
xor U16302 (N_16302,N_16132,N_16084);
nor U16303 (N_16303,N_16076,N_16022);
or U16304 (N_16304,N_16072,N_16087);
nand U16305 (N_16305,N_16040,N_16135);
or U16306 (N_16306,N_16058,N_16080);
nand U16307 (N_16307,N_16116,N_16016);
and U16308 (N_16308,N_16112,N_16071);
nor U16309 (N_16309,N_16122,N_16031);
nor U16310 (N_16310,N_16095,N_16132);
nand U16311 (N_16311,N_16103,N_16006);
nand U16312 (N_16312,N_16139,N_16109);
nand U16313 (N_16313,N_16042,N_16131);
nand U16314 (N_16314,N_16005,N_16043);
xnor U16315 (N_16315,N_16041,N_16154);
xnor U16316 (N_16316,N_16128,N_16137);
or U16317 (N_16317,N_16092,N_16048);
or U16318 (N_16318,N_16036,N_16076);
nor U16319 (N_16319,N_16120,N_16056);
and U16320 (N_16320,N_16268,N_16163);
nand U16321 (N_16321,N_16277,N_16302);
nand U16322 (N_16322,N_16247,N_16171);
or U16323 (N_16323,N_16231,N_16172);
nor U16324 (N_16324,N_16295,N_16313);
nand U16325 (N_16325,N_16173,N_16276);
nor U16326 (N_16326,N_16300,N_16297);
xnor U16327 (N_16327,N_16209,N_16176);
and U16328 (N_16328,N_16265,N_16291);
nand U16329 (N_16329,N_16308,N_16304);
nand U16330 (N_16330,N_16298,N_16273);
and U16331 (N_16331,N_16292,N_16279);
nand U16332 (N_16332,N_16278,N_16233);
or U16333 (N_16333,N_16286,N_16315);
or U16334 (N_16334,N_16167,N_16262);
nand U16335 (N_16335,N_16183,N_16222);
nor U16336 (N_16336,N_16217,N_16160);
nand U16337 (N_16337,N_16256,N_16214);
nor U16338 (N_16338,N_16283,N_16178);
nand U16339 (N_16339,N_16177,N_16165);
and U16340 (N_16340,N_16230,N_16274);
nor U16341 (N_16341,N_16208,N_16210);
or U16342 (N_16342,N_16319,N_16311);
and U16343 (N_16343,N_16179,N_16185);
or U16344 (N_16344,N_16245,N_16285);
nand U16345 (N_16345,N_16267,N_16250);
nand U16346 (N_16346,N_16246,N_16249);
xor U16347 (N_16347,N_16296,N_16260);
or U16348 (N_16348,N_16161,N_16257);
or U16349 (N_16349,N_16166,N_16306);
or U16350 (N_16350,N_16175,N_16213);
and U16351 (N_16351,N_16248,N_16187);
nand U16352 (N_16352,N_16201,N_16221);
and U16353 (N_16353,N_16228,N_16318);
nand U16354 (N_16354,N_16216,N_16272);
and U16355 (N_16355,N_16182,N_16164);
nand U16356 (N_16356,N_16303,N_16237);
and U16357 (N_16357,N_16263,N_16219);
and U16358 (N_16358,N_16266,N_16241);
nand U16359 (N_16359,N_16189,N_16215);
nand U16360 (N_16360,N_16211,N_16314);
and U16361 (N_16361,N_16280,N_16199);
and U16362 (N_16362,N_16204,N_16261);
and U16363 (N_16363,N_16243,N_16238);
xnor U16364 (N_16364,N_16220,N_16229);
nor U16365 (N_16365,N_16271,N_16253);
nand U16366 (N_16366,N_16290,N_16312);
and U16367 (N_16367,N_16305,N_16316);
and U16368 (N_16368,N_16240,N_16224);
nor U16369 (N_16369,N_16317,N_16259);
or U16370 (N_16370,N_16293,N_16270);
xnor U16371 (N_16371,N_16301,N_16299);
nor U16372 (N_16372,N_16195,N_16168);
nand U16373 (N_16373,N_16307,N_16170);
nand U16374 (N_16374,N_16186,N_16288);
xor U16375 (N_16375,N_16232,N_16206);
and U16376 (N_16376,N_16212,N_16198);
and U16377 (N_16377,N_16207,N_16287);
nor U16378 (N_16378,N_16239,N_16200);
or U16379 (N_16379,N_16196,N_16281);
xor U16380 (N_16380,N_16310,N_16227);
nand U16381 (N_16381,N_16252,N_16236);
and U16382 (N_16382,N_16202,N_16194);
nor U16383 (N_16383,N_16169,N_16275);
nand U16384 (N_16384,N_16226,N_16190);
or U16385 (N_16385,N_16255,N_16203);
nand U16386 (N_16386,N_16258,N_16174);
nand U16387 (N_16387,N_16192,N_16180);
xnor U16388 (N_16388,N_16284,N_16188);
nor U16389 (N_16389,N_16162,N_16289);
nand U16390 (N_16390,N_16242,N_16294);
or U16391 (N_16391,N_16264,N_16282);
nor U16392 (N_16392,N_16225,N_16269);
nor U16393 (N_16393,N_16197,N_16251);
xor U16394 (N_16394,N_16191,N_16244);
or U16395 (N_16395,N_16205,N_16254);
and U16396 (N_16396,N_16181,N_16184);
nor U16397 (N_16397,N_16235,N_16218);
or U16398 (N_16398,N_16309,N_16234);
or U16399 (N_16399,N_16223,N_16193);
or U16400 (N_16400,N_16216,N_16185);
and U16401 (N_16401,N_16263,N_16210);
and U16402 (N_16402,N_16287,N_16218);
xor U16403 (N_16403,N_16308,N_16223);
nor U16404 (N_16404,N_16293,N_16165);
nand U16405 (N_16405,N_16269,N_16302);
and U16406 (N_16406,N_16296,N_16166);
nand U16407 (N_16407,N_16287,N_16236);
or U16408 (N_16408,N_16278,N_16236);
nor U16409 (N_16409,N_16286,N_16248);
nand U16410 (N_16410,N_16201,N_16183);
nor U16411 (N_16411,N_16169,N_16310);
nor U16412 (N_16412,N_16247,N_16168);
nand U16413 (N_16413,N_16209,N_16182);
or U16414 (N_16414,N_16192,N_16170);
or U16415 (N_16415,N_16300,N_16200);
nand U16416 (N_16416,N_16177,N_16237);
nand U16417 (N_16417,N_16200,N_16175);
xnor U16418 (N_16418,N_16292,N_16264);
nand U16419 (N_16419,N_16228,N_16301);
nand U16420 (N_16420,N_16241,N_16308);
or U16421 (N_16421,N_16245,N_16169);
nor U16422 (N_16422,N_16238,N_16244);
nand U16423 (N_16423,N_16228,N_16299);
nand U16424 (N_16424,N_16318,N_16302);
nor U16425 (N_16425,N_16287,N_16244);
and U16426 (N_16426,N_16304,N_16188);
nor U16427 (N_16427,N_16187,N_16297);
xor U16428 (N_16428,N_16176,N_16201);
nand U16429 (N_16429,N_16196,N_16234);
xor U16430 (N_16430,N_16193,N_16244);
xnor U16431 (N_16431,N_16254,N_16281);
or U16432 (N_16432,N_16302,N_16191);
nand U16433 (N_16433,N_16302,N_16237);
xnor U16434 (N_16434,N_16219,N_16258);
or U16435 (N_16435,N_16313,N_16165);
nand U16436 (N_16436,N_16196,N_16171);
or U16437 (N_16437,N_16273,N_16251);
nand U16438 (N_16438,N_16285,N_16215);
or U16439 (N_16439,N_16317,N_16194);
nor U16440 (N_16440,N_16205,N_16194);
nor U16441 (N_16441,N_16292,N_16244);
and U16442 (N_16442,N_16249,N_16221);
and U16443 (N_16443,N_16232,N_16241);
nor U16444 (N_16444,N_16268,N_16232);
or U16445 (N_16445,N_16205,N_16240);
nor U16446 (N_16446,N_16227,N_16234);
nor U16447 (N_16447,N_16197,N_16319);
nand U16448 (N_16448,N_16319,N_16290);
nor U16449 (N_16449,N_16289,N_16252);
nor U16450 (N_16450,N_16216,N_16240);
nor U16451 (N_16451,N_16302,N_16213);
or U16452 (N_16452,N_16223,N_16244);
nand U16453 (N_16453,N_16202,N_16179);
nand U16454 (N_16454,N_16198,N_16240);
xor U16455 (N_16455,N_16315,N_16230);
nor U16456 (N_16456,N_16235,N_16187);
xor U16457 (N_16457,N_16250,N_16187);
or U16458 (N_16458,N_16317,N_16191);
xnor U16459 (N_16459,N_16259,N_16172);
and U16460 (N_16460,N_16251,N_16188);
and U16461 (N_16461,N_16203,N_16282);
xnor U16462 (N_16462,N_16214,N_16202);
and U16463 (N_16463,N_16244,N_16263);
xor U16464 (N_16464,N_16246,N_16239);
and U16465 (N_16465,N_16303,N_16195);
nand U16466 (N_16466,N_16319,N_16249);
nand U16467 (N_16467,N_16183,N_16265);
and U16468 (N_16468,N_16206,N_16184);
or U16469 (N_16469,N_16317,N_16252);
or U16470 (N_16470,N_16198,N_16179);
or U16471 (N_16471,N_16273,N_16170);
nor U16472 (N_16472,N_16213,N_16178);
and U16473 (N_16473,N_16198,N_16237);
nor U16474 (N_16474,N_16306,N_16252);
or U16475 (N_16475,N_16183,N_16163);
nor U16476 (N_16476,N_16177,N_16304);
or U16477 (N_16477,N_16315,N_16272);
nand U16478 (N_16478,N_16183,N_16319);
nand U16479 (N_16479,N_16247,N_16170);
and U16480 (N_16480,N_16409,N_16350);
or U16481 (N_16481,N_16421,N_16441);
xnor U16482 (N_16482,N_16369,N_16433);
xor U16483 (N_16483,N_16334,N_16354);
xor U16484 (N_16484,N_16321,N_16331);
nor U16485 (N_16485,N_16457,N_16419);
nand U16486 (N_16486,N_16403,N_16473);
and U16487 (N_16487,N_16469,N_16393);
nand U16488 (N_16488,N_16351,N_16320);
nor U16489 (N_16489,N_16366,N_16358);
or U16490 (N_16490,N_16423,N_16324);
nand U16491 (N_16491,N_16442,N_16396);
nand U16492 (N_16492,N_16322,N_16456);
nor U16493 (N_16493,N_16459,N_16417);
xor U16494 (N_16494,N_16328,N_16323);
nand U16495 (N_16495,N_16385,N_16426);
or U16496 (N_16496,N_16411,N_16340);
nand U16497 (N_16497,N_16335,N_16438);
or U16498 (N_16498,N_16355,N_16451);
nand U16499 (N_16499,N_16439,N_16364);
and U16500 (N_16500,N_16341,N_16363);
xor U16501 (N_16501,N_16425,N_16461);
or U16502 (N_16502,N_16389,N_16388);
nor U16503 (N_16503,N_16443,N_16359);
nor U16504 (N_16504,N_16436,N_16477);
or U16505 (N_16505,N_16434,N_16376);
nand U16506 (N_16506,N_16375,N_16404);
nor U16507 (N_16507,N_16325,N_16468);
nor U16508 (N_16508,N_16410,N_16378);
xnor U16509 (N_16509,N_16336,N_16418);
nand U16510 (N_16510,N_16394,N_16420);
nand U16511 (N_16511,N_16383,N_16400);
xnor U16512 (N_16512,N_16380,N_16356);
or U16513 (N_16513,N_16395,N_16478);
and U16514 (N_16514,N_16445,N_16475);
nand U16515 (N_16515,N_16344,N_16472);
or U16516 (N_16516,N_16357,N_16384);
xnor U16517 (N_16517,N_16450,N_16402);
or U16518 (N_16518,N_16405,N_16416);
or U16519 (N_16519,N_16386,N_16353);
nor U16520 (N_16520,N_16329,N_16377);
xnor U16521 (N_16521,N_16365,N_16455);
nor U16522 (N_16522,N_16352,N_16337);
nand U16523 (N_16523,N_16346,N_16467);
nor U16524 (N_16524,N_16429,N_16348);
and U16525 (N_16525,N_16454,N_16427);
nand U16526 (N_16526,N_16448,N_16367);
xnor U16527 (N_16527,N_16339,N_16407);
nand U16528 (N_16528,N_16474,N_16447);
xor U16529 (N_16529,N_16338,N_16412);
xnor U16530 (N_16530,N_16440,N_16430);
nor U16531 (N_16531,N_16373,N_16479);
and U16532 (N_16532,N_16361,N_16462);
xnor U16533 (N_16533,N_16332,N_16437);
and U16534 (N_16534,N_16414,N_16428);
nor U16535 (N_16535,N_16342,N_16471);
xnor U16536 (N_16536,N_16374,N_16415);
xor U16537 (N_16537,N_16382,N_16449);
and U16538 (N_16538,N_16431,N_16371);
nand U16539 (N_16539,N_16333,N_16452);
xor U16540 (N_16540,N_16381,N_16330);
xor U16541 (N_16541,N_16387,N_16343);
xnor U16542 (N_16542,N_16326,N_16347);
nand U16543 (N_16543,N_16463,N_16397);
nand U16544 (N_16544,N_16372,N_16401);
nand U16545 (N_16545,N_16422,N_16406);
nand U16546 (N_16546,N_16460,N_16349);
nor U16547 (N_16547,N_16398,N_16413);
nand U16548 (N_16548,N_16432,N_16464);
or U16549 (N_16549,N_16390,N_16408);
or U16550 (N_16550,N_16360,N_16458);
or U16551 (N_16551,N_16446,N_16453);
nand U16552 (N_16552,N_16399,N_16379);
or U16553 (N_16553,N_16466,N_16444);
xor U16554 (N_16554,N_16435,N_16370);
and U16555 (N_16555,N_16424,N_16327);
or U16556 (N_16556,N_16391,N_16476);
nand U16557 (N_16557,N_16392,N_16362);
nand U16558 (N_16558,N_16345,N_16368);
nand U16559 (N_16559,N_16470,N_16465);
nand U16560 (N_16560,N_16472,N_16448);
nand U16561 (N_16561,N_16442,N_16388);
nor U16562 (N_16562,N_16476,N_16435);
and U16563 (N_16563,N_16338,N_16329);
nor U16564 (N_16564,N_16375,N_16449);
nor U16565 (N_16565,N_16321,N_16421);
xnor U16566 (N_16566,N_16337,N_16331);
or U16567 (N_16567,N_16464,N_16447);
or U16568 (N_16568,N_16432,N_16389);
and U16569 (N_16569,N_16391,N_16390);
xor U16570 (N_16570,N_16393,N_16366);
xnor U16571 (N_16571,N_16374,N_16400);
xnor U16572 (N_16572,N_16477,N_16435);
nand U16573 (N_16573,N_16444,N_16441);
nor U16574 (N_16574,N_16467,N_16441);
nand U16575 (N_16575,N_16469,N_16410);
nand U16576 (N_16576,N_16327,N_16454);
nand U16577 (N_16577,N_16320,N_16470);
and U16578 (N_16578,N_16434,N_16449);
or U16579 (N_16579,N_16456,N_16371);
nand U16580 (N_16580,N_16397,N_16376);
xor U16581 (N_16581,N_16396,N_16424);
nand U16582 (N_16582,N_16335,N_16368);
nor U16583 (N_16583,N_16427,N_16389);
nor U16584 (N_16584,N_16429,N_16323);
nand U16585 (N_16585,N_16398,N_16461);
nor U16586 (N_16586,N_16459,N_16354);
nor U16587 (N_16587,N_16422,N_16420);
nor U16588 (N_16588,N_16393,N_16424);
nor U16589 (N_16589,N_16478,N_16466);
xor U16590 (N_16590,N_16465,N_16440);
xnor U16591 (N_16591,N_16382,N_16394);
or U16592 (N_16592,N_16386,N_16457);
and U16593 (N_16593,N_16338,N_16444);
xnor U16594 (N_16594,N_16467,N_16442);
xnor U16595 (N_16595,N_16433,N_16411);
or U16596 (N_16596,N_16372,N_16371);
or U16597 (N_16597,N_16335,N_16406);
or U16598 (N_16598,N_16381,N_16459);
and U16599 (N_16599,N_16389,N_16397);
and U16600 (N_16600,N_16360,N_16425);
or U16601 (N_16601,N_16433,N_16322);
xnor U16602 (N_16602,N_16326,N_16337);
and U16603 (N_16603,N_16411,N_16358);
nor U16604 (N_16604,N_16354,N_16322);
and U16605 (N_16605,N_16351,N_16403);
nor U16606 (N_16606,N_16365,N_16475);
or U16607 (N_16607,N_16429,N_16430);
and U16608 (N_16608,N_16460,N_16382);
nor U16609 (N_16609,N_16361,N_16477);
nor U16610 (N_16610,N_16384,N_16393);
xor U16611 (N_16611,N_16432,N_16362);
xor U16612 (N_16612,N_16365,N_16354);
xnor U16613 (N_16613,N_16445,N_16388);
nand U16614 (N_16614,N_16406,N_16389);
and U16615 (N_16615,N_16334,N_16337);
or U16616 (N_16616,N_16428,N_16321);
nor U16617 (N_16617,N_16351,N_16333);
and U16618 (N_16618,N_16349,N_16457);
or U16619 (N_16619,N_16406,N_16332);
nor U16620 (N_16620,N_16353,N_16453);
xor U16621 (N_16621,N_16401,N_16329);
and U16622 (N_16622,N_16411,N_16452);
nor U16623 (N_16623,N_16421,N_16331);
and U16624 (N_16624,N_16374,N_16406);
nand U16625 (N_16625,N_16375,N_16410);
and U16626 (N_16626,N_16347,N_16450);
xor U16627 (N_16627,N_16478,N_16404);
nand U16628 (N_16628,N_16378,N_16347);
and U16629 (N_16629,N_16343,N_16420);
xor U16630 (N_16630,N_16380,N_16385);
or U16631 (N_16631,N_16440,N_16417);
nor U16632 (N_16632,N_16405,N_16426);
nand U16633 (N_16633,N_16423,N_16328);
or U16634 (N_16634,N_16320,N_16399);
nor U16635 (N_16635,N_16447,N_16386);
and U16636 (N_16636,N_16408,N_16333);
and U16637 (N_16637,N_16425,N_16323);
nand U16638 (N_16638,N_16407,N_16476);
nand U16639 (N_16639,N_16408,N_16410);
xor U16640 (N_16640,N_16510,N_16483);
nand U16641 (N_16641,N_16590,N_16517);
nand U16642 (N_16642,N_16627,N_16482);
nor U16643 (N_16643,N_16575,N_16624);
nand U16644 (N_16644,N_16528,N_16531);
nor U16645 (N_16645,N_16509,N_16552);
xnor U16646 (N_16646,N_16586,N_16619);
or U16647 (N_16647,N_16617,N_16579);
nand U16648 (N_16648,N_16566,N_16615);
nand U16649 (N_16649,N_16563,N_16634);
nor U16650 (N_16650,N_16535,N_16609);
nor U16651 (N_16651,N_16606,N_16582);
xnor U16652 (N_16652,N_16537,N_16522);
and U16653 (N_16653,N_16625,N_16505);
xnor U16654 (N_16654,N_16564,N_16519);
nor U16655 (N_16655,N_16636,N_16507);
and U16656 (N_16656,N_16592,N_16530);
xnor U16657 (N_16657,N_16596,N_16536);
and U16658 (N_16658,N_16570,N_16577);
nor U16659 (N_16659,N_16623,N_16554);
nand U16660 (N_16660,N_16626,N_16589);
xnor U16661 (N_16661,N_16631,N_16557);
xnor U16662 (N_16662,N_16493,N_16565);
nor U16663 (N_16663,N_16559,N_16605);
or U16664 (N_16664,N_16578,N_16608);
and U16665 (N_16665,N_16513,N_16548);
or U16666 (N_16666,N_16489,N_16639);
xnor U16667 (N_16667,N_16511,N_16602);
and U16668 (N_16668,N_16599,N_16540);
and U16669 (N_16669,N_16543,N_16572);
and U16670 (N_16670,N_16629,N_16583);
xor U16671 (N_16671,N_16499,N_16614);
xnor U16672 (N_16672,N_16516,N_16593);
nand U16673 (N_16673,N_16546,N_16492);
and U16674 (N_16674,N_16635,N_16491);
xor U16675 (N_16675,N_16598,N_16594);
xnor U16676 (N_16676,N_16562,N_16628);
and U16677 (N_16677,N_16485,N_16553);
nand U16678 (N_16678,N_16480,N_16607);
nand U16679 (N_16679,N_16534,N_16560);
xor U16680 (N_16680,N_16585,N_16527);
and U16681 (N_16681,N_16620,N_16568);
nor U16682 (N_16682,N_16576,N_16514);
or U16683 (N_16683,N_16630,N_16584);
nor U16684 (N_16684,N_16501,N_16547);
nor U16685 (N_16685,N_16542,N_16588);
and U16686 (N_16686,N_16616,N_16612);
nand U16687 (N_16687,N_16632,N_16498);
and U16688 (N_16688,N_16488,N_16529);
nand U16689 (N_16689,N_16539,N_16613);
nand U16690 (N_16690,N_16622,N_16504);
and U16691 (N_16691,N_16541,N_16621);
or U16692 (N_16692,N_16580,N_16497);
or U16693 (N_16693,N_16486,N_16512);
or U16694 (N_16694,N_16496,N_16525);
nor U16695 (N_16695,N_16494,N_16487);
nor U16696 (N_16696,N_16597,N_16544);
and U16697 (N_16697,N_16500,N_16603);
xnor U16698 (N_16698,N_16545,N_16521);
or U16699 (N_16699,N_16611,N_16569);
or U16700 (N_16700,N_16571,N_16600);
or U16701 (N_16701,N_16595,N_16508);
or U16702 (N_16702,N_16555,N_16574);
nor U16703 (N_16703,N_16573,N_16550);
and U16704 (N_16704,N_16633,N_16532);
nand U16705 (N_16705,N_16523,N_16549);
nor U16706 (N_16706,N_16518,N_16524);
or U16707 (N_16707,N_16618,N_16533);
or U16708 (N_16708,N_16502,N_16591);
nor U16709 (N_16709,N_16561,N_16503);
or U16710 (N_16710,N_16538,N_16637);
or U16711 (N_16711,N_16587,N_16558);
nor U16712 (N_16712,N_16610,N_16495);
or U16713 (N_16713,N_16506,N_16604);
or U16714 (N_16714,N_16551,N_16481);
and U16715 (N_16715,N_16515,N_16638);
nor U16716 (N_16716,N_16526,N_16556);
nor U16717 (N_16717,N_16484,N_16490);
xnor U16718 (N_16718,N_16567,N_16520);
or U16719 (N_16719,N_16601,N_16581);
nand U16720 (N_16720,N_16565,N_16498);
or U16721 (N_16721,N_16600,N_16633);
nor U16722 (N_16722,N_16616,N_16509);
nand U16723 (N_16723,N_16610,N_16580);
nor U16724 (N_16724,N_16519,N_16597);
and U16725 (N_16725,N_16631,N_16510);
xnor U16726 (N_16726,N_16499,N_16575);
nand U16727 (N_16727,N_16531,N_16511);
or U16728 (N_16728,N_16517,N_16617);
or U16729 (N_16729,N_16574,N_16492);
or U16730 (N_16730,N_16527,N_16561);
or U16731 (N_16731,N_16637,N_16572);
and U16732 (N_16732,N_16480,N_16507);
xnor U16733 (N_16733,N_16527,N_16486);
or U16734 (N_16734,N_16510,N_16505);
nor U16735 (N_16735,N_16523,N_16542);
or U16736 (N_16736,N_16538,N_16598);
and U16737 (N_16737,N_16487,N_16601);
xnor U16738 (N_16738,N_16594,N_16612);
and U16739 (N_16739,N_16552,N_16487);
or U16740 (N_16740,N_16518,N_16516);
or U16741 (N_16741,N_16517,N_16532);
and U16742 (N_16742,N_16522,N_16595);
nand U16743 (N_16743,N_16512,N_16545);
nor U16744 (N_16744,N_16565,N_16578);
or U16745 (N_16745,N_16516,N_16521);
nand U16746 (N_16746,N_16540,N_16558);
nand U16747 (N_16747,N_16506,N_16521);
and U16748 (N_16748,N_16499,N_16600);
nand U16749 (N_16749,N_16495,N_16522);
nor U16750 (N_16750,N_16511,N_16596);
or U16751 (N_16751,N_16505,N_16578);
and U16752 (N_16752,N_16599,N_16510);
nand U16753 (N_16753,N_16514,N_16540);
nor U16754 (N_16754,N_16572,N_16525);
or U16755 (N_16755,N_16557,N_16560);
and U16756 (N_16756,N_16588,N_16625);
or U16757 (N_16757,N_16579,N_16533);
nor U16758 (N_16758,N_16594,N_16631);
nor U16759 (N_16759,N_16561,N_16636);
nand U16760 (N_16760,N_16587,N_16522);
and U16761 (N_16761,N_16542,N_16569);
nand U16762 (N_16762,N_16504,N_16519);
nand U16763 (N_16763,N_16512,N_16521);
nor U16764 (N_16764,N_16569,N_16605);
and U16765 (N_16765,N_16490,N_16524);
nand U16766 (N_16766,N_16605,N_16519);
and U16767 (N_16767,N_16560,N_16554);
or U16768 (N_16768,N_16566,N_16525);
nor U16769 (N_16769,N_16520,N_16585);
or U16770 (N_16770,N_16601,N_16529);
nor U16771 (N_16771,N_16612,N_16548);
and U16772 (N_16772,N_16522,N_16585);
and U16773 (N_16773,N_16624,N_16617);
and U16774 (N_16774,N_16587,N_16638);
xor U16775 (N_16775,N_16533,N_16632);
nor U16776 (N_16776,N_16636,N_16554);
nor U16777 (N_16777,N_16486,N_16621);
and U16778 (N_16778,N_16570,N_16503);
xnor U16779 (N_16779,N_16494,N_16574);
and U16780 (N_16780,N_16538,N_16558);
and U16781 (N_16781,N_16506,N_16536);
nand U16782 (N_16782,N_16623,N_16563);
and U16783 (N_16783,N_16490,N_16491);
nor U16784 (N_16784,N_16610,N_16489);
nand U16785 (N_16785,N_16609,N_16501);
xor U16786 (N_16786,N_16536,N_16627);
and U16787 (N_16787,N_16626,N_16602);
nand U16788 (N_16788,N_16502,N_16539);
nor U16789 (N_16789,N_16490,N_16481);
and U16790 (N_16790,N_16483,N_16607);
nor U16791 (N_16791,N_16578,N_16585);
and U16792 (N_16792,N_16568,N_16610);
nor U16793 (N_16793,N_16548,N_16497);
or U16794 (N_16794,N_16502,N_16635);
xnor U16795 (N_16795,N_16493,N_16601);
nand U16796 (N_16796,N_16603,N_16588);
or U16797 (N_16797,N_16516,N_16509);
or U16798 (N_16798,N_16553,N_16548);
nor U16799 (N_16799,N_16519,N_16551);
xnor U16800 (N_16800,N_16697,N_16795);
xnor U16801 (N_16801,N_16673,N_16725);
and U16802 (N_16802,N_16664,N_16737);
and U16803 (N_16803,N_16742,N_16779);
nor U16804 (N_16804,N_16693,N_16690);
nand U16805 (N_16805,N_16659,N_16705);
or U16806 (N_16806,N_16712,N_16796);
or U16807 (N_16807,N_16759,N_16711);
or U16808 (N_16808,N_16760,N_16658);
nor U16809 (N_16809,N_16793,N_16723);
and U16810 (N_16810,N_16738,N_16700);
and U16811 (N_16811,N_16672,N_16676);
nor U16812 (N_16812,N_16698,N_16791);
xor U16813 (N_16813,N_16765,N_16713);
nor U16814 (N_16814,N_16655,N_16643);
nor U16815 (N_16815,N_16644,N_16758);
or U16816 (N_16816,N_16652,N_16767);
nor U16817 (N_16817,N_16718,N_16721);
and U16818 (N_16818,N_16744,N_16692);
and U16819 (N_16819,N_16716,N_16772);
xnor U16820 (N_16820,N_16774,N_16743);
and U16821 (N_16821,N_16787,N_16694);
or U16822 (N_16822,N_16683,N_16670);
xor U16823 (N_16823,N_16726,N_16657);
nor U16824 (N_16824,N_16691,N_16769);
nor U16825 (N_16825,N_16794,N_16717);
or U16826 (N_16826,N_16747,N_16654);
nor U16827 (N_16827,N_16651,N_16753);
or U16828 (N_16828,N_16750,N_16665);
nand U16829 (N_16829,N_16732,N_16646);
nand U16830 (N_16830,N_16666,N_16682);
nor U16831 (N_16831,N_16730,N_16797);
nor U16832 (N_16832,N_16704,N_16688);
nand U16833 (N_16833,N_16776,N_16780);
or U16834 (N_16834,N_16728,N_16669);
or U16835 (N_16835,N_16689,N_16660);
or U16836 (N_16836,N_16731,N_16739);
and U16837 (N_16837,N_16695,N_16663);
nand U16838 (N_16838,N_16798,N_16770);
or U16839 (N_16839,N_16746,N_16761);
nor U16840 (N_16840,N_16755,N_16680);
nor U16841 (N_16841,N_16778,N_16773);
xnor U16842 (N_16842,N_16771,N_16786);
xnor U16843 (N_16843,N_16714,N_16679);
nand U16844 (N_16844,N_16649,N_16645);
or U16845 (N_16845,N_16648,N_16668);
xor U16846 (N_16846,N_16764,N_16667);
xor U16847 (N_16847,N_16707,N_16642);
nand U16848 (N_16848,N_16671,N_16662);
or U16849 (N_16849,N_16782,N_16789);
nand U16850 (N_16850,N_16745,N_16729);
nor U16851 (N_16851,N_16741,N_16681);
xnor U16852 (N_16852,N_16661,N_16762);
xnor U16853 (N_16853,N_16696,N_16763);
or U16854 (N_16854,N_16653,N_16751);
xor U16855 (N_16855,N_16685,N_16715);
and U16856 (N_16856,N_16788,N_16701);
nor U16857 (N_16857,N_16790,N_16784);
xnor U16858 (N_16858,N_16684,N_16720);
and U16859 (N_16859,N_16677,N_16733);
and U16860 (N_16860,N_16709,N_16647);
or U16861 (N_16861,N_16699,N_16766);
or U16862 (N_16862,N_16768,N_16703);
and U16863 (N_16863,N_16687,N_16706);
nor U16864 (N_16864,N_16675,N_16640);
xnor U16865 (N_16865,N_16736,N_16777);
xor U16866 (N_16866,N_16749,N_16710);
and U16867 (N_16867,N_16781,N_16727);
or U16868 (N_16868,N_16775,N_16740);
nor U16869 (N_16869,N_16735,N_16678);
and U16870 (N_16870,N_16656,N_16754);
nor U16871 (N_16871,N_16799,N_16686);
nor U16872 (N_16872,N_16724,N_16719);
nor U16873 (N_16873,N_16702,N_16783);
xnor U16874 (N_16874,N_16785,N_16674);
and U16875 (N_16875,N_16757,N_16752);
or U16876 (N_16876,N_16650,N_16722);
nand U16877 (N_16877,N_16641,N_16756);
xnor U16878 (N_16878,N_16734,N_16708);
nor U16879 (N_16879,N_16748,N_16792);
nor U16880 (N_16880,N_16648,N_16746);
and U16881 (N_16881,N_16785,N_16742);
and U16882 (N_16882,N_16757,N_16642);
nor U16883 (N_16883,N_16721,N_16731);
nand U16884 (N_16884,N_16712,N_16787);
xor U16885 (N_16885,N_16797,N_16690);
nand U16886 (N_16886,N_16782,N_16768);
xnor U16887 (N_16887,N_16690,N_16763);
nor U16888 (N_16888,N_16712,N_16662);
nand U16889 (N_16889,N_16712,N_16791);
xor U16890 (N_16890,N_16766,N_16799);
nor U16891 (N_16891,N_16703,N_16788);
or U16892 (N_16892,N_16715,N_16750);
and U16893 (N_16893,N_16747,N_16684);
or U16894 (N_16894,N_16698,N_16737);
or U16895 (N_16895,N_16719,N_16739);
or U16896 (N_16896,N_16705,N_16715);
or U16897 (N_16897,N_16649,N_16719);
nor U16898 (N_16898,N_16731,N_16655);
nand U16899 (N_16899,N_16706,N_16698);
and U16900 (N_16900,N_16674,N_16683);
nor U16901 (N_16901,N_16716,N_16667);
nor U16902 (N_16902,N_16748,N_16753);
and U16903 (N_16903,N_16778,N_16766);
nand U16904 (N_16904,N_16758,N_16658);
nand U16905 (N_16905,N_16679,N_16761);
nand U16906 (N_16906,N_16721,N_16674);
nand U16907 (N_16907,N_16689,N_16671);
nor U16908 (N_16908,N_16756,N_16767);
xor U16909 (N_16909,N_16670,N_16781);
nand U16910 (N_16910,N_16703,N_16692);
xor U16911 (N_16911,N_16642,N_16769);
or U16912 (N_16912,N_16753,N_16772);
and U16913 (N_16913,N_16658,N_16737);
or U16914 (N_16914,N_16672,N_16655);
or U16915 (N_16915,N_16671,N_16685);
and U16916 (N_16916,N_16787,N_16641);
or U16917 (N_16917,N_16751,N_16788);
or U16918 (N_16918,N_16766,N_16656);
nand U16919 (N_16919,N_16781,N_16756);
xnor U16920 (N_16920,N_16796,N_16737);
and U16921 (N_16921,N_16742,N_16720);
xor U16922 (N_16922,N_16771,N_16649);
xnor U16923 (N_16923,N_16640,N_16695);
nand U16924 (N_16924,N_16702,N_16706);
nand U16925 (N_16925,N_16726,N_16647);
nand U16926 (N_16926,N_16643,N_16779);
and U16927 (N_16927,N_16661,N_16791);
nor U16928 (N_16928,N_16706,N_16797);
or U16929 (N_16929,N_16650,N_16771);
or U16930 (N_16930,N_16726,N_16768);
nor U16931 (N_16931,N_16790,N_16654);
nand U16932 (N_16932,N_16644,N_16709);
xnor U16933 (N_16933,N_16787,N_16719);
and U16934 (N_16934,N_16648,N_16720);
or U16935 (N_16935,N_16689,N_16737);
nor U16936 (N_16936,N_16727,N_16789);
nor U16937 (N_16937,N_16707,N_16732);
and U16938 (N_16938,N_16724,N_16734);
nand U16939 (N_16939,N_16767,N_16788);
nand U16940 (N_16940,N_16729,N_16688);
and U16941 (N_16941,N_16736,N_16707);
nand U16942 (N_16942,N_16791,N_16683);
and U16943 (N_16943,N_16667,N_16761);
nor U16944 (N_16944,N_16650,N_16647);
and U16945 (N_16945,N_16796,N_16720);
nor U16946 (N_16946,N_16750,N_16788);
or U16947 (N_16947,N_16696,N_16793);
nor U16948 (N_16948,N_16690,N_16689);
and U16949 (N_16949,N_16793,N_16645);
and U16950 (N_16950,N_16759,N_16792);
nand U16951 (N_16951,N_16648,N_16684);
nand U16952 (N_16952,N_16725,N_16691);
and U16953 (N_16953,N_16781,N_16797);
nand U16954 (N_16954,N_16757,N_16713);
or U16955 (N_16955,N_16641,N_16758);
nor U16956 (N_16956,N_16643,N_16664);
or U16957 (N_16957,N_16752,N_16666);
nor U16958 (N_16958,N_16785,N_16770);
xor U16959 (N_16959,N_16691,N_16714);
and U16960 (N_16960,N_16820,N_16930);
nor U16961 (N_16961,N_16816,N_16875);
xor U16962 (N_16962,N_16865,N_16948);
and U16963 (N_16963,N_16831,N_16897);
nand U16964 (N_16964,N_16886,N_16841);
xnor U16965 (N_16965,N_16837,N_16913);
and U16966 (N_16966,N_16942,N_16805);
nor U16967 (N_16967,N_16952,N_16864);
and U16968 (N_16968,N_16927,N_16843);
or U16969 (N_16969,N_16945,N_16850);
nor U16970 (N_16970,N_16924,N_16933);
or U16971 (N_16971,N_16825,N_16856);
nand U16972 (N_16972,N_16898,N_16908);
nor U16973 (N_16973,N_16903,N_16809);
nand U16974 (N_16974,N_16951,N_16862);
xor U16975 (N_16975,N_16955,N_16828);
and U16976 (N_16976,N_16815,N_16920);
and U16977 (N_16977,N_16880,N_16851);
nand U16978 (N_16978,N_16925,N_16946);
xnor U16979 (N_16979,N_16804,N_16943);
xnor U16980 (N_16980,N_16909,N_16817);
or U16981 (N_16981,N_16863,N_16802);
nand U16982 (N_16982,N_16896,N_16867);
and U16983 (N_16983,N_16823,N_16860);
and U16984 (N_16984,N_16822,N_16879);
xnor U16985 (N_16985,N_16826,N_16894);
or U16986 (N_16986,N_16824,N_16885);
and U16987 (N_16987,N_16949,N_16891);
nor U16988 (N_16988,N_16890,N_16857);
nor U16989 (N_16989,N_16959,N_16842);
and U16990 (N_16990,N_16905,N_16819);
and U16991 (N_16991,N_16931,N_16953);
and U16992 (N_16992,N_16835,N_16878);
nand U16993 (N_16993,N_16902,N_16844);
and U16994 (N_16994,N_16957,N_16868);
and U16995 (N_16995,N_16892,N_16893);
nand U16996 (N_16996,N_16855,N_16883);
and U16997 (N_16997,N_16910,N_16919);
or U16998 (N_16998,N_16830,N_16888);
nand U16999 (N_16999,N_16916,N_16838);
or U17000 (N_17000,N_16818,N_16836);
xor U17001 (N_17001,N_16956,N_16950);
xor U17002 (N_17002,N_16901,N_16846);
and U17003 (N_17003,N_16859,N_16872);
xor U17004 (N_17004,N_16833,N_16944);
and U17005 (N_17005,N_16803,N_16932);
or U17006 (N_17006,N_16811,N_16889);
xor U17007 (N_17007,N_16884,N_16926);
xnor U17008 (N_17008,N_16914,N_16839);
or U17009 (N_17009,N_16801,N_16870);
xnor U17010 (N_17010,N_16941,N_16881);
xnor U17011 (N_17011,N_16906,N_16807);
nand U17012 (N_17012,N_16882,N_16939);
or U17013 (N_17013,N_16813,N_16847);
nor U17014 (N_17014,N_16900,N_16907);
and U17015 (N_17015,N_16827,N_16904);
nor U17016 (N_17016,N_16940,N_16917);
nand U17017 (N_17017,N_16934,N_16874);
nor U17018 (N_17018,N_16869,N_16832);
and U17019 (N_17019,N_16873,N_16806);
xor U17020 (N_17020,N_16814,N_16936);
nand U17021 (N_17021,N_16852,N_16922);
xnor U17022 (N_17022,N_16866,N_16821);
and U17023 (N_17023,N_16928,N_16853);
and U17024 (N_17024,N_16921,N_16915);
and U17025 (N_17025,N_16911,N_16834);
xnor U17026 (N_17026,N_16845,N_16854);
nand U17027 (N_17027,N_16848,N_16858);
xnor U17028 (N_17028,N_16876,N_16887);
or U17029 (N_17029,N_16935,N_16808);
nor U17030 (N_17030,N_16895,N_16861);
and U17031 (N_17031,N_16912,N_16812);
nor U17032 (N_17032,N_16929,N_16918);
and U17033 (N_17033,N_16871,N_16947);
or U17034 (N_17034,N_16923,N_16877);
xor U17035 (N_17035,N_16810,N_16840);
and U17036 (N_17036,N_16937,N_16954);
xnor U17037 (N_17037,N_16829,N_16958);
or U17038 (N_17038,N_16938,N_16800);
and U17039 (N_17039,N_16899,N_16849);
nand U17040 (N_17040,N_16899,N_16916);
xnor U17041 (N_17041,N_16884,N_16805);
or U17042 (N_17042,N_16917,N_16958);
and U17043 (N_17043,N_16830,N_16918);
and U17044 (N_17044,N_16836,N_16891);
and U17045 (N_17045,N_16871,N_16938);
or U17046 (N_17046,N_16803,N_16878);
nand U17047 (N_17047,N_16902,N_16939);
and U17048 (N_17048,N_16843,N_16916);
and U17049 (N_17049,N_16919,N_16854);
nor U17050 (N_17050,N_16925,N_16821);
nor U17051 (N_17051,N_16877,N_16931);
and U17052 (N_17052,N_16863,N_16818);
or U17053 (N_17053,N_16805,N_16886);
or U17054 (N_17054,N_16827,N_16800);
or U17055 (N_17055,N_16802,N_16905);
xnor U17056 (N_17056,N_16824,N_16880);
xnor U17057 (N_17057,N_16868,N_16801);
xor U17058 (N_17058,N_16865,N_16833);
and U17059 (N_17059,N_16903,N_16825);
or U17060 (N_17060,N_16875,N_16802);
xnor U17061 (N_17061,N_16838,N_16847);
and U17062 (N_17062,N_16943,N_16919);
nand U17063 (N_17063,N_16921,N_16900);
and U17064 (N_17064,N_16856,N_16912);
or U17065 (N_17065,N_16896,N_16800);
nor U17066 (N_17066,N_16954,N_16949);
xnor U17067 (N_17067,N_16852,N_16806);
or U17068 (N_17068,N_16836,N_16831);
nand U17069 (N_17069,N_16843,N_16853);
nor U17070 (N_17070,N_16826,N_16898);
xnor U17071 (N_17071,N_16823,N_16928);
xnor U17072 (N_17072,N_16919,N_16801);
xor U17073 (N_17073,N_16923,N_16904);
nand U17074 (N_17074,N_16846,N_16853);
nand U17075 (N_17075,N_16911,N_16859);
nand U17076 (N_17076,N_16887,N_16842);
nor U17077 (N_17077,N_16807,N_16806);
xor U17078 (N_17078,N_16944,N_16959);
or U17079 (N_17079,N_16917,N_16918);
and U17080 (N_17080,N_16890,N_16823);
xor U17081 (N_17081,N_16938,N_16918);
nand U17082 (N_17082,N_16944,N_16824);
and U17083 (N_17083,N_16828,N_16854);
nand U17084 (N_17084,N_16877,N_16818);
nand U17085 (N_17085,N_16878,N_16925);
or U17086 (N_17086,N_16831,N_16800);
nand U17087 (N_17087,N_16806,N_16836);
xor U17088 (N_17088,N_16871,N_16831);
or U17089 (N_17089,N_16826,N_16873);
nand U17090 (N_17090,N_16812,N_16911);
xor U17091 (N_17091,N_16857,N_16826);
nand U17092 (N_17092,N_16886,N_16954);
xnor U17093 (N_17093,N_16952,N_16853);
xor U17094 (N_17094,N_16945,N_16886);
nor U17095 (N_17095,N_16932,N_16806);
or U17096 (N_17096,N_16857,N_16836);
or U17097 (N_17097,N_16880,N_16945);
xnor U17098 (N_17098,N_16953,N_16861);
and U17099 (N_17099,N_16953,N_16857);
or U17100 (N_17100,N_16851,N_16845);
and U17101 (N_17101,N_16884,N_16804);
and U17102 (N_17102,N_16892,N_16812);
nand U17103 (N_17103,N_16900,N_16814);
nand U17104 (N_17104,N_16811,N_16867);
or U17105 (N_17105,N_16874,N_16811);
or U17106 (N_17106,N_16854,N_16870);
nor U17107 (N_17107,N_16890,N_16932);
or U17108 (N_17108,N_16845,N_16903);
and U17109 (N_17109,N_16934,N_16958);
or U17110 (N_17110,N_16895,N_16853);
nand U17111 (N_17111,N_16803,N_16880);
and U17112 (N_17112,N_16903,N_16818);
or U17113 (N_17113,N_16880,N_16810);
nand U17114 (N_17114,N_16912,N_16815);
nor U17115 (N_17115,N_16861,N_16869);
xor U17116 (N_17116,N_16942,N_16815);
nand U17117 (N_17117,N_16820,N_16917);
nand U17118 (N_17118,N_16923,N_16888);
nand U17119 (N_17119,N_16806,N_16954);
or U17120 (N_17120,N_16993,N_17111);
xor U17121 (N_17121,N_16976,N_17061);
xor U17122 (N_17122,N_17010,N_16981);
and U17123 (N_17123,N_17050,N_16960);
or U17124 (N_17124,N_16967,N_17099);
xnor U17125 (N_17125,N_17100,N_17006);
xor U17126 (N_17126,N_17118,N_17011);
or U17127 (N_17127,N_16964,N_17027);
and U17128 (N_17128,N_16970,N_17065);
nor U17129 (N_17129,N_16991,N_17063);
xor U17130 (N_17130,N_16972,N_17003);
and U17131 (N_17131,N_17064,N_17102);
or U17132 (N_17132,N_16998,N_17021);
or U17133 (N_17133,N_17093,N_16982);
nor U17134 (N_17134,N_16969,N_17101);
xor U17135 (N_17135,N_17070,N_17001);
nor U17136 (N_17136,N_16999,N_17092);
or U17137 (N_17137,N_17016,N_16996);
nand U17138 (N_17138,N_17052,N_17029);
nor U17139 (N_17139,N_17051,N_16977);
nand U17140 (N_17140,N_17081,N_17038);
nor U17141 (N_17141,N_17025,N_17071);
nand U17142 (N_17142,N_17053,N_17107);
nand U17143 (N_17143,N_16975,N_17077);
xnor U17144 (N_17144,N_17043,N_17087);
nor U17145 (N_17145,N_17067,N_17008);
xnor U17146 (N_17146,N_17096,N_17110);
xnor U17147 (N_17147,N_17091,N_17002);
nand U17148 (N_17148,N_16988,N_16978);
or U17149 (N_17149,N_17073,N_16994);
nand U17150 (N_17150,N_17035,N_17045);
and U17151 (N_17151,N_17088,N_17116);
nor U17152 (N_17152,N_17036,N_16973);
nor U17153 (N_17153,N_16965,N_17031);
or U17154 (N_17154,N_16968,N_17047);
or U17155 (N_17155,N_17098,N_16997);
nand U17156 (N_17156,N_17095,N_16974);
nor U17157 (N_17157,N_16990,N_17058);
nor U17158 (N_17158,N_17033,N_17028);
and U17159 (N_17159,N_17117,N_17005);
nor U17160 (N_17160,N_16986,N_17072);
nand U17161 (N_17161,N_16961,N_17076);
nor U17162 (N_17162,N_17040,N_16984);
xnor U17163 (N_17163,N_17037,N_17032);
or U17164 (N_17164,N_17044,N_17039);
xor U17165 (N_17165,N_17049,N_17082);
xnor U17166 (N_17166,N_17115,N_17094);
or U17167 (N_17167,N_17004,N_17057);
nand U17168 (N_17168,N_16971,N_17119);
nand U17169 (N_17169,N_17020,N_17034);
or U17170 (N_17170,N_17060,N_17069);
nand U17171 (N_17171,N_16987,N_17078);
or U17172 (N_17172,N_17023,N_17113);
or U17173 (N_17173,N_17009,N_17018);
or U17174 (N_17174,N_17086,N_16962);
nor U17175 (N_17175,N_17024,N_17103);
xor U17176 (N_17176,N_17066,N_17022);
nand U17177 (N_17177,N_17083,N_16963);
or U17178 (N_17178,N_17068,N_17090);
nand U17179 (N_17179,N_17108,N_16995);
xor U17180 (N_17180,N_17104,N_17079);
and U17181 (N_17181,N_17012,N_17026);
nor U17182 (N_17182,N_17056,N_16992);
and U17183 (N_17183,N_17017,N_17084);
nor U17184 (N_17184,N_17041,N_17080);
nor U17185 (N_17185,N_16979,N_16985);
or U17186 (N_17186,N_17085,N_17042);
nand U17187 (N_17187,N_17097,N_17048);
nor U17188 (N_17188,N_17054,N_16983);
nor U17189 (N_17189,N_17014,N_17105);
xnor U17190 (N_17190,N_17109,N_17019);
and U17191 (N_17191,N_17062,N_17000);
or U17192 (N_17192,N_17106,N_16980);
xor U17193 (N_17193,N_17059,N_16989);
nor U17194 (N_17194,N_17015,N_17030);
xor U17195 (N_17195,N_17089,N_17114);
nor U17196 (N_17196,N_17075,N_17074);
or U17197 (N_17197,N_17007,N_16966);
and U17198 (N_17198,N_17112,N_17055);
xor U17199 (N_17199,N_17013,N_17046);
or U17200 (N_17200,N_17044,N_17035);
nor U17201 (N_17201,N_17055,N_17048);
nand U17202 (N_17202,N_16996,N_17105);
nor U17203 (N_17203,N_17001,N_17085);
and U17204 (N_17204,N_17062,N_17079);
xnor U17205 (N_17205,N_17107,N_17113);
nor U17206 (N_17206,N_17095,N_17000);
xor U17207 (N_17207,N_17096,N_16970);
and U17208 (N_17208,N_17086,N_17117);
and U17209 (N_17209,N_17119,N_17049);
nand U17210 (N_17210,N_17078,N_16964);
nor U17211 (N_17211,N_16999,N_17062);
nor U17212 (N_17212,N_17067,N_17070);
nand U17213 (N_17213,N_16967,N_17113);
and U17214 (N_17214,N_16992,N_17073);
and U17215 (N_17215,N_17021,N_17025);
or U17216 (N_17216,N_17081,N_17044);
and U17217 (N_17217,N_17000,N_16979);
nor U17218 (N_17218,N_17092,N_17033);
or U17219 (N_17219,N_17051,N_17115);
nor U17220 (N_17220,N_17069,N_17062);
xnor U17221 (N_17221,N_17097,N_16999);
or U17222 (N_17222,N_17091,N_17078);
nand U17223 (N_17223,N_16994,N_17041);
or U17224 (N_17224,N_17091,N_16964);
nor U17225 (N_17225,N_16990,N_17114);
and U17226 (N_17226,N_17062,N_16991);
nand U17227 (N_17227,N_17083,N_17009);
or U17228 (N_17228,N_17047,N_16966);
nor U17229 (N_17229,N_16998,N_17067);
xnor U17230 (N_17230,N_17056,N_17110);
nand U17231 (N_17231,N_17050,N_17093);
or U17232 (N_17232,N_17053,N_17007);
and U17233 (N_17233,N_17072,N_17059);
nor U17234 (N_17234,N_16988,N_16965);
or U17235 (N_17235,N_16992,N_17101);
xor U17236 (N_17236,N_17079,N_17084);
xor U17237 (N_17237,N_17018,N_17040);
and U17238 (N_17238,N_17051,N_17021);
xnor U17239 (N_17239,N_17036,N_17043);
nand U17240 (N_17240,N_17036,N_16996);
and U17241 (N_17241,N_17119,N_16974);
xnor U17242 (N_17242,N_17019,N_17026);
nor U17243 (N_17243,N_17018,N_16974);
or U17244 (N_17244,N_17045,N_17030);
and U17245 (N_17245,N_17046,N_17075);
nand U17246 (N_17246,N_16981,N_17080);
and U17247 (N_17247,N_17080,N_16992);
xor U17248 (N_17248,N_17102,N_17096);
or U17249 (N_17249,N_16996,N_17011);
nand U17250 (N_17250,N_16960,N_16996);
or U17251 (N_17251,N_17034,N_17102);
and U17252 (N_17252,N_17017,N_17050);
xnor U17253 (N_17253,N_17030,N_17081);
or U17254 (N_17254,N_17115,N_17113);
or U17255 (N_17255,N_17083,N_17049);
nand U17256 (N_17256,N_16995,N_17003);
and U17257 (N_17257,N_17010,N_17039);
xnor U17258 (N_17258,N_17057,N_16987);
xor U17259 (N_17259,N_17083,N_16970);
or U17260 (N_17260,N_16969,N_16995);
nand U17261 (N_17261,N_16998,N_16968);
nor U17262 (N_17262,N_17009,N_17002);
and U17263 (N_17263,N_17079,N_17037);
nor U17264 (N_17264,N_17101,N_17065);
and U17265 (N_17265,N_17056,N_16977);
and U17266 (N_17266,N_16980,N_17008);
and U17267 (N_17267,N_17087,N_16979);
xor U17268 (N_17268,N_17035,N_16993);
nor U17269 (N_17269,N_17029,N_17079);
or U17270 (N_17270,N_16978,N_17015);
nor U17271 (N_17271,N_17013,N_17062);
nor U17272 (N_17272,N_17013,N_17100);
nand U17273 (N_17273,N_17110,N_17022);
nor U17274 (N_17274,N_16978,N_16960);
or U17275 (N_17275,N_16987,N_16969);
xnor U17276 (N_17276,N_17058,N_17000);
nand U17277 (N_17277,N_17098,N_17058);
nor U17278 (N_17278,N_17057,N_17050);
or U17279 (N_17279,N_17002,N_17051);
nor U17280 (N_17280,N_17169,N_17160);
and U17281 (N_17281,N_17146,N_17157);
nor U17282 (N_17282,N_17184,N_17245);
xnor U17283 (N_17283,N_17234,N_17209);
nand U17284 (N_17284,N_17170,N_17208);
nand U17285 (N_17285,N_17173,N_17154);
nand U17286 (N_17286,N_17125,N_17165);
nand U17287 (N_17287,N_17152,N_17229);
xor U17288 (N_17288,N_17195,N_17134);
xnor U17289 (N_17289,N_17132,N_17238);
nand U17290 (N_17290,N_17270,N_17274);
or U17291 (N_17291,N_17262,N_17232);
nor U17292 (N_17292,N_17167,N_17181);
and U17293 (N_17293,N_17228,N_17139);
nor U17294 (N_17294,N_17264,N_17244);
or U17295 (N_17295,N_17137,N_17136);
or U17296 (N_17296,N_17135,N_17242);
xnor U17297 (N_17297,N_17226,N_17158);
nor U17298 (N_17298,N_17194,N_17256);
xor U17299 (N_17299,N_17269,N_17258);
or U17300 (N_17300,N_17176,N_17163);
nor U17301 (N_17301,N_17252,N_17259);
or U17302 (N_17302,N_17235,N_17183);
and U17303 (N_17303,N_17166,N_17123);
or U17304 (N_17304,N_17149,N_17240);
and U17305 (N_17305,N_17192,N_17178);
or U17306 (N_17306,N_17272,N_17273);
xnor U17307 (N_17307,N_17187,N_17250);
or U17308 (N_17308,N_17239,N_17161);
nor U17309 (N_17309,N_17214,N_17253);
and U17310 (N_17310,N_17279,N_17126);
nand U17311 (N_17311,N_17130,N_17122);
nand U17312 (N_17312,N_17260,N_17222);
nand U17313 (N_17313,N_17241,N_17121);
nor U17314 (N_17314,N_17221,N_17144);
nand U17315 (N_17315,N_17202,N_17205);
and U17316 (N_17316,N_17153,N_17265);
and U17317 (N_17317,N_17162,N_17268);
and U17318 (N_17318,N_17248,N_17147);
and U17319 (N_17319,N_17142,N_17217);
or U17320 (N_17320,N_17247,N_17257);
nor U17321 (N_17321,N_17156,N_17174);
nand U17322 (N_17322,N_17215,N_17190);
nor U17323 (N_17323,N_17180,N_17278);
xnor U17324 (N_17324,N_17197,N_17172);
nor U17325 (N_17325,N_17138,N_17150);
and U17326 (N_17326,N_17218,N_17206);
nand U17327 (N_17327,N_17225,N_17255);
nand U17328 (N_17328,N_17230,N_17277);
nor U17329 (N_17329,N_17151,N_17236);
or U17330 (N_17330,N_17124,N_17219);
nor U17331 (N_17331,N_17212,N_17220);
or U17332 (N_17332,N_17128,N_17243);
nand U17333 (N_17333,N_17155,N_17196);
nor U17334 (N_17334,N_17182,N_17177);
xnor U17335 (N_17335,N_17164,N_17276);
or U17336 (N_17336,N_17246,N_17127);
xnor U17337 (N_17337,N_17120,N_17275);
nand U17338 (N_17338,N_17193,N_17200);
or U17339 (N_17339,N_17168,N_17141);
xor U17340 (N_17340,N_17233,N_17261);
and U17341 (N_17341,N_17251,N_17224);
and U17342 (N_17342,N_17249,N_17203);
xor U17343 (N_17343,N_17171,N_17231);
and U17344 (N_17344,N_17263,N_17143);
or U17345 (N_17345,N_17159,N_17129);
or U17346 (N_17346,N_17213,N_17133);
xnor U17347 (N_17347,N_17216,N_17188);
and U17348 (N_17348,N_17131,N_17204);
xnor U17349 (N_17349,N_17140,N_17266);
nand U17350 (N_17350,N_17191,N_17179);
or U17351 (N_17351,N_17199,N_17185);
nor U17352 (N_17352,N_17237,N_17223);
nor U17353 (N_17353,N_17201,N_17254);
or U17354 (N_17354,N_17175,N_17189);
and U17355 (N_17355,N_17148,N_17211);
nand U17356 (N_17356,N_17186,N_17267);
or U17357 (N_17357,N_17198,N_17207);
or U17358 (N_17358,N_17271,N_17210);
or U17359 (N_17359,N_17227,N_17145);
nor U17360 (N_17360,N_17195,N_17133);
and U17361 (N_17361,N_17154,N_17202);
nor U17362 (N_17362,N_17270,N_17182);
nand U17363 (N_17363,N_17267,N_17142);
and U17364 (N_17364,N_17267,N_17126);
and U17365 (N_17365,N_17270,N_17228);
xor U17366 (N_17366,N_17196,N_17165);
nor U17367 (N_17367,N_17143,N_17274);
xor U17368 (N_17368,N_17173,N_17195);
nand U17369 (N_17369,N_17202,N_17251);
or U17370 (N_17370,N_17198,N_17195);
or U17371 (N_17371,N_17121,N_17184);
nor U17372 (N_17372,N_17127,N_17190);
or U17373 (N_17373,N_17237,N_17279);
xnor U17374 (N_17374,N_17268,N_17225);
nand U17375 (N_17375,N_17163,N_17223);
and U17376 (N_17376,N_17173,N_17244);
and U17377 (N_17377,N_17272,N_17143);
xor U17378 (N_17378,N_17201,N_17149);
and U17379 (N_17379,N_17161,N_17246);
xor U17380 (N_17380,N_17136,N_17255);
xor U17381 (N_17381,N_17195,N_17207);
and U17382 (N_17382,N_17171,N_17238);
nor U17383 (N_17383,N_17273,N_17148);
or U17384 (N_17384,N_17243,N_17234);
nand U17385 (N_17385,N_17204,N_17216);
nor U17386 (N_17386,N_17238,N_17239);
nand U17387 (N_17387,N_17163,N_17268);
nand U17388 (N_17388,N_17239,N_17273);
or U17389 (N_17389,N_17270,N_17165);
and U17390 (N_17390,N_17275,N_17207);
nor U17391 (N_17391,N_17249,N_17235);
nand U17392 (N_17392,N_17157,N_17121);
nor U17393 (N_17393,N_17162,N_17191);
or U17394 (N_17394,N_17139,N_17165);
or U17395 (N_17395,N_17183,N_17236);
and U17396 (N_17396,N_17210,N_17202);
nor U17397 (N_17397,N_17147,N_17277);
and U17398 (N_17398,N_17156,N_17265);
or U17399 (N_17399,N_17152,N_17132);
and U17400 (N_17400,N_17142,N_17277);
nand U17401 (N_17401,N_17149,N_17249);
or U17402 (N_17402,N_17155,N_17247);
xor U17403 (N_17403,N_17141,N_17250);
nor U17404 (N_17404,N_17253,N_17259);
and U17405 (N_17405,N_17136,N_17190);
nand U17406 (N_17406,N_17204,N_17260);
xor U17407 (N_17407,N_17190,N_17238);
xor U17408 (N_17408,N_17226,N_17128);
nand U17409 (N_17409,N_17266,N_17264);
nand U17410 (N_17410,N_17239,N_17200);
xor U17411 (N_17411,N_17244,N_17271);
xnor U17412 (N_17412,N_17158,N_17195);
nand U17413 (N_17413,N_17174,N_17148);
nand U17414 (N_17414,N_17163,N_17233);
nand U17415 (N_17415,N_17185,N_17165);
or U17416 (N_17416,N_17168,N_17185);
xnor U17417 (N_17417,N_17240,N_17177);
or U17418 (N_17418,N_17215,N_17133);
xor U17419 (N_17419,N_17134,N_17144);
nand U17420 (N_17420,N_17120,N_17255);
and U17421 (N_17421,N_17163,N_17231);
and U17422 (N_17422,N_17212,N_17150);
and U17423 (N_17423,N_17216,N_17138);
nand U17424 (N_17424,N_17131,N_17172);
nor U17425 (N_17425,N_17254,N_17181);
and U17426 (N_17426,N_17127,N_17165);
xor U17427 (N_17427,N_17127,N_17132);
nor U17428 (N_17428,N_17144,N_17223);
xnor U17429 (N_17429,N_17247,N_17217);
nand U17430 (N_17430,N_17127,N_17227);
and U17431 (N_17431,N_17224,N_17166);
xnor U17432 (N_17432,N_17149,N_17277);
or U17433 (N_17433,N_17123,N_17223);
nor U17434 (N_17434,N_17150,N_17167);
nor U17435 (N_17435,N_17149,N_17158);
or U17436 (N_17436,N_17150,N_17240);
nor U17437 (N_17437,N_17197,N_17248);
or U17438 (N_17438,N_17165,N_17273);
xnor U17439 (N_17439,N_17211,N_17255);
nor U17440 (N_17440,N_17390,N_17396);
nand U17441 (N_17441,N_17401,N_17336);
and U17442 (N_17442,N_17324,N_17316);
nor U17443 (N_17443,N_17338,N_17373);
xor U17444 (N_17444,N_17410,N_17293);
or U17445 (N_17445,N_17395,N_17351);
or U17446 (N_17446,N_17439,N_17381);
xor U17447 (N_17447,N_17391,N_17436);
nor U17448 (N_17448,N_17307,N_17429);
xor U17449 (N_17449,N_17302,N_17416);
xor U17450 (N_17450,N_17327,N_17413);
nor U17451 (N_17451,N_17286,N_17418);
xnor U17452 (N_17452,N_17386,N_17389);
or U17453 (N_17453,N_17420,N_17438);
or U17454 (N_17454,N_17354,N_17406);
or U17455 (N_17455,N_17350,N_17320);
nand U17456 (N_17456,N_17311,N_17367);
nand U17457 (N_17457,N_17362,N_17353);
nand U17458 (N_17458,N_17310,N_17281);
or U17459 (N_17459,N_17408,N_17411);
nand U17460 (N_17460,N_17403,N_17394);
nand U17461 (N_17461,N_17375,N_17347);
nor U17462 (N_17462,N_17342,N_17330);
and U17463 (N_17463,N_17318,N_17332);
nor U17464 (N_17464,N_17392,N_17405);
and U17465 (N_17465,N_17326,N_17321);
nand U17466 (N_17466,N_17363,N_17341);
xnor U17467 (N_17467,N_17368,N_17393);
nor U17468 (N_17468,N_17319,N_17382);
xnor U17469 (N_17469,N_17372,N_17397);
xor U17470 (N_17470,N_17300,N_17377);
and U17471 (N_17471,N_17304,N_17427);
nor U17472 (N_17472,N_17322,N_17346);
and U17473 (N_17473,N_17407,N_17366);
and U17474 (N_17474,N_17313,N_17371);
or U17475 (N_17475,N_17325,N_17361);
nand U17476 (N_17476,N_17296,N_17305);
nand U17477 (N_17477,N_17387,N_17365);
nand U17478 (N_17478,N_17308,N_17331);
nor U17479 (N_17479,N_17352,N_17328);
and U17480 (N_17480,N_17376,N_17432);
and U17481 (N_17481,N_17399,N_17380);
nand U17482 (N_17482,N_17434,N_17423);
or U17483 (N_17483,N_17359,N_17426);
or U17484 (N_17484,N_17345,N_17433);
xor U17485 (N_17485,N_17417,N_17385);
nand U17486 (N_17486,N_17398,N_17283);
nand U17487 (N_17487,N_17284,N_17412);
nand U17488 (N_17488,N_17297,N_17337);
xnor U17489 (N_17489,N_17355,N_17340);
nand U17490 (N_17490,N_17298,N_17388);
xor U17491 (N_17491,N_17369,N_17312);
or U17492 (N_17492,N_17435,N_17414);
or U17493 (N_17493,N_17409,N_17335);
and U17494 (N_17494,N_17437,N_17384);
nand U17495 (N_17495,N_17428,N_17292);
nor U17496 (N_17496,N_17317,N_17333);
nand U17497 (N_17497,N_17287,N_17379);
xnor U17498 (N_17498,N_17400,N_17364);
or U17499 (N_17499,N_17370,N_17289);
and U17500 (N_17500,N_17285,N_17344);
nand U17501 (N_17501,N_17309,N_17314);
xnor U17502 (N_17502,N_17356,N_17339);
or U17503 (N_17503,N_17357,N_17349);
nand U17504 (N_17504,N_17334,N_17280);
nand U17505 (N_17505,N_17301,N_17378);
or U17506 (N_17506,N_17383,N_17295);
nor U17507 (N_17507,N_17299,N_17323);
nand U17508 (N_17508,N_17282,N_17404);
nand U17509 (N_17509,N_17421,N_17430);
or U17510 (N_17510,N_17431,N_17348);
nand U17511 (N_17511,N_17415,N_17329);
and U17512 (N_17512,N_17288,N_17422);
nor U17513 (N_17513,N_17315,N_17294);
or U17514 (N_17514,N_17424,N_17374);
xor U17515 (N_17515,N_17291,N_17303);
xor U17516 (N_17516,N_17343,N_17402);
or U17517 (N_17517,N_17290,N_17360);
and U17518 (N_17518,N_17358,N_17425);
nand U17519 (N_17519,N_17306,N_17419);
or U17520 (N_17520,N_17322,N_17310);
and U17521 (N_17521,N_17384,N_17436);
nor U17522 (N_17522,N_17437,N_17389);
or U17523 (N_17523,N_17328,N_17325);
xnor U17524 (N_17524,N_17317,N_17360);
nand U17525 (N_17525,N_17313,N_17412);
nor U17526 (N_17526,N_17326,N_17431);
and U17527 (N_17527,N_17358,N_17426);
nand U17528 (N_17528,N_17300,N_17344);
or U17529 (N_17529,N_17295,N_17380);
nand U17530 (N_17530,N_17421,N_17387);
and U17531 (N_17531,N_17328,N_17437);
nand U17532 (N_17532,N_17325,N_17307);
nor U17533 (N_17533,N_17322,N_17439);
nand U17534 (N_17534,N_17366,N_17336);
or U17535 (N_17535,N_17291,N_17379);
nand U17536 (N_17536,N_17365,N_17297);
nand U17537 (N_17537,N_17383,N_17336);
xnor U17538 (N_17538,N_17387,N_17406);
nor U17539 (N_17539,N_17339,N_17308);
and U17540 (N_17540,N_17393,N_17435);
nand U17541 (N_17541,N_17376,N_17302);
or U17542 (N_17542,N_17294,N_17310);
nand U17543 (N_17543,N_17320,N_17364);
nand U17544 (N_17544,N_17432,N_17403);
nand U17545 (N_17545,N_17298,N_17412);
or U17546 (N_17546,N_17401,N_17416);
and U17547 (N_17547,N_17392,N_17400);
and U17548 (N_17548,N_17388,N_17412);
nand U17549 (N_17549,N_17314,N_17354);
nand U17550 (N_17550,N_17368,N_17347);
nor U17551 (N_17551,N_17333,N_17301);
nor U17552 (N_17552,N_17325,N_17434);
nor U17553 (N_17553,N_17417,N_17373);
nor U17554 (N_17554,N_17364,N_17402);
or U17555 (N_17555,N_17370,N_17409);
xor U17556 (N_17556,N_17411,N_17353);
and U17557 (N_17557,N_17290,N_17395);
and U17558 (N_17558,N_17355,N_17304);
or U17559 (N_17559,N_17353,N_17437);
nand U17560 (N_17560,N_17430,N_17426);
nor U17561 (N_17561,N_17296,N_17308);
nand U17562 (N_17562,N_17325,N_17401);
or U17563 (N_17563,N_17351,N_17363);
nand U17564 (N_17564,N_17362,N_17303);
nand U17565 (N_17565,N_17397,N_17409);
nor U17566 (N_17566,N_17312,N_17359);
xor U17567 (N_17567,N_17305,N_17291);
nand U17568 (N_17568,N_17337,N_17341);
and U17569 (N_17569,N_17308,N_17317);
or U17570 (N_17570,N_17300,N_17434);
and U17571 (N_17571,N_17433,N_17373);
or U17572 (N_17572,N_17438,N_17351);
and U17573 (N_17573,N_17408,N_17434);
nand U17574 (N_17574,N_17353,N_17427);
nand U17575 (N_17575,N_17410,N_17321);
nor U17576 (N_17576,N_17292,N_17338);
or U17577 (N_17577,N_17362,N_17342);
or U17578 (N_17578,N_17359,N_17433);
and U17579 (N_17579,N_17357,N_17352);
and U17580 (N_17580,N_17438,N_17300);
xor U17581 (N_17581,N_17403,N_17385);
or U17582 (N_17582,N_17338,N_17375);
and U17583 (N_17583,N_17367,N_17316);
xor U17584 (N_17584,N_17301,N_17385);
nor U17585 (N_17585,N_17381,N_17301);
and U17586 (N_17586,N_17323,N_17302);
and U17587 (N_17587,N_17350,N_17426);
nor U17588 (N_17588,N_17412,N_17392);
or U17589 (N_17589,N_17299,N_17378);
nand U17590 (N_17590,N_17292,N_17311);
nor U17591 (N_17591,N_17391,N_17421);
nand U17592 (N_17592,N_17338,N_17303);
nor U17593 (N_17593,N_17314,N_17419);
xnor U17594 (N_17594,N_17373,N_17283);
nand U17595 (N_17595,N_17354,N_17383);
nor U17596 (N_17596,N_17433,N_17305);
nand U17597 (N_17597,N_17362,N_17434);
and U17598 (N_17598,N_17280,N_17314);
and U17599 (N_17599,N_17367,N_17428);
nor U17600 (N_17600,N_17447,N_17572);
nand U17601 (N_17601,N_17518,N_17584);
or U17602 (N_17602,N_17473,N_17596);
nand U17603 (N_17603,N_17570,N_17482);
xor U17604 (N_17604,N_17485,N_17543);
and U17605 (N_17605,N_17597,N_17449);
nor U17606 (N_17606,N_17554,N_17452);
nand U17607 (N_17607,N_17571,N_17458);
nand U17608 (N_17608,N_17581,N_17493);
and U17609 (N_17609,N_17537,N_17462);
nand U17610 (N_17610,N_17488,N_17490);
nand U17611 (N_17611,N_17467,N_17511);
and U17612 (N_17612,N_17509,N_17475);
or U17613 (N_17613,N_17507,N_17534);
nor U17614 (N_17614,N_17594,N_17464);
xor U17615 (N_17615,N_17499,N_17539);
or U17616 (N_17616,N_17491,N_17561);
or U17617 (N_17617,N_17536,N_17598);
or U17618 (N_17618,N_17589,N_17495);
nand U17619 (N_17619,N_17540,N_17528);
nand U17620 (N_17620,N_17472,N_17592);
and U17621 (N_17621,N_17496,N_17522);
nand U17622 (N_17622,N_17586,N_17574);
xor U17623 (N_17623,N_17544,N_17483);
nor U17624 (N_17624,N_17446,N_17550);
and U17625 (N_17625,N_17497,N_17577);
nand U17626 (N_17626,N_17578,N_17564);
and U17627 (N_17627,N_17532,N_17448);
and U17628 (N_17628,N_17521,N_17551);
nor U17629 (N_17629,N_17484,N_17548);
xor U17630 (N_17630,N_17530,N_17531);
or U17631 (N_17631,N_17588,N_17508);
xnor U17632 (N_17632,N_17468,N_17479);
xor U17633 (N_17633,N_17580,N_17444);
xnor U17634 (N_17634,N_17525,N_17535);
xnor U17635 (N_17635,N_17465,N_17556);
nor U17636 (N_17636,N_17503,N_17579);
nor U17637 (N_17637,N_17529,N_17524);
and U17638 (N_17638,N_17494,N_17587);
nor U17639 (N_17639,N_17478,N_17593);
or U17640 (N_17640,N_17568,N_17516);
nand U17641 (N_17641,N_17480,N_17533);
and U17642 (N_17642,N_17560,N_17454);
nor U17643 (N_17643,N_17456,N_17471);
or U17644 (N_17644,N_17585,N_17517);
and U17645 (N_17645,N_17569,N_17498);
xnor U17646 (N_17646,N_17559,N_17591);
and U17647 (N_17647,N_17443,N_17575);
and U17648 (N_17648,N_17545,N_17466);
nor U17649 (N_17649,N_17546,N_17576);
nand U17650 (N_17650,N_17504,N_17451);
xnor U17651 (N_17651,N_17502,N_17514);
nand U17652 (N_17652,N_17526,N_17541);
xnor U17653 (N_17653,N_17573,N_17510);
and U17654 (N_17654,N_17557,N_17523);
or U17655 (N_17655,N_17527,N_17453);
and U17656 (N_17656,N_17565,N_17590);
and U17657 (N_17657,N_17455,N_17552);
nor U17658 (N_17658,N_17520,N_17599);
xnor U17659 (N_17659,N_17549,N_17460);
xor U17660 (N_17660,N_17547,N_17558);
nand U17661 (N_17661,N_17440,N_17489);
or U17662 (N_17662,N_17463,N_17486);
nand U17663 (N_17663,N_17505,N_17487);
or U17664 (N_17664,N_17519,N_17567);
or U17665 (N_17665,N_17470,N_17542);
xor U17666 (N_17666,N_17595,N_17492);
or U17667 (N_17667,N_17538,N_17515);
or U17668 (N_17668,N_17461,N_17512);
and U17669 (N_17669,N_17562,N_17506);
nand U17670 (N_17670,N_17563,N_17501);
or U17671 (N_17671,N_17553,N_17500);
nand U17672 (N_17672,N_17459,N_17469);
nand U17673 (N_17673,N_17477,N_17445);
nand U17674 (N_17674,N_17441,N_17476);
xor U17675 (N_17675,N_17481,N_17555);
nor U17676 (N_17676,N_17474,N_17450);
xnor U17677 (N_17677,N_17442,N_17582);
or U17678 (N_17678,N_17457,N_17513);
nand U17679 (N_17679,N_17566,N_17583);
nand U17680 (N_17680,N_17544,N_17484);
nor U17681 (N_17681,N_17476,N_17529);
nand U17682 (N_17682,N_17479,N_17482);
nor U17683 (N_17683,N_17493,N_17450);
nand U17684 (N_17684,N_17474,N_17452);
nand U17685 (N_17685,N_17499,N_17579);
nand U17686 (N_17686,N_17549,N_17570);
nor U17687 (N_17687,N_17580,N_17466);
and U17688 (N_17688,N_17596,N_17482);
nor U17689 (N_17689,N_17588,N_17502);
xnor U17690 (N_17690,N_17534,N_17524);
nand U17691 (N_17691,N_17508,N_17553);
or U17692 (N_17692,N_17574,N_17519);
nand U17693 (N_17693,N_17486,N_17511);
nand U17694 (N_17694,N_17590,N_17563);
xor U17695 (N_17695,N_17588,N_17451);
nand U17696 (N_17696,N_17584,N_17536);
or U17697 (N_17697,N_17475,N_17469);
or U17698 (N_17698,N_17466,N_17473);
and U17699 (N_17699,N_17456,N_17457);
xor U17700 (N_17700,N_17542,N_17585);
or U17701 (N_17701,N_17498,N_17554);
or U17702 (N_17702,N_17546,N_17520);
nor U17703 (N_17703,N_17453,N_17505);
nand U17704 (N_17704,N_17510,N_17451);
or U17705 (N_17705,N_17531,N_17573);
and U17706 (N_17706,N_17523,N_17575);
and U17707 (N_17707,N_17461,N_17462);
and U17708 (N_17708,N_17560,N_17500);
or U17709 (N_17709,N_17515,N_17469);
or U17710 (N_17710,N_17450,N_17445);
nor U17711 (N_17711,N_17465,N_17555);
and U17712 (N_17712,N_17452,N_17542);
nor U17713 (N_17713,N_17563,N_17537);
nand U17714 (N_17714,N_17477,N_17440);
nor U17715 (N_17715,N_17461,N_17593);
nor U17716 (N_17716,N_17470,N_17597);
or U17717 (N_17717,N_17478,N_17453);
nand U17718 (N_17718,N_17517,N_17456);
nor U17719 (N_17719,N_17584,N_17454);
nand U17720 (N_17720,N_17471,N_17579);
nor U17721 (N_17721,N_17491,N_17484);
nor U17722 (N_17722,N_17567,N_17497);
and U17723 (N_17723,N_17484,N_17474);
nand U17724 (N_17724,N_17597,N_17590);
nor U17725 (N_17725,N_17455,N_17479);
nor U17726 (N_17726,N_17556,N_17565);
or U17727 (N_17727,N_17577,N_17512);
xnor U17728 (N_17728,N_17480,N_17561);
xnor U17729 (N_17729,N_17596,N_17528);
nand U17730 (N_17730,N_17521,N_17440);
nor U17731 (N_17731,N_17479,N_17461);
nand U17732 (N_17732,N_17494,N_17497);
or U17733 (N_17733,N_17552,N_17534);
and U17734 (N_17734,N_17544,N_17497);
nor U17735 (N_17735,N_17477,N_17540);
nand U17736 (N_17736,N_17527,N_17536);
nand U17737 (N_17737,N_17549,N_17541);
xor U17738 (N_17738,N_17596,N_17493);
nand U17739 (N_17739,N_17568,N_17571);
and U17740 (N_17740,N_17443,N_17539);
and U17741 (N_17741,N_17480,N_17449);
or U17742 (N_17742,N_17484,N_17594);
nand U17743 (N_17743,N_17487,N_17492);
nor U17744 (N_17744,N_17440,N_17536);
xor U17745 (N_17745,N_17444,N_17557);
and U17746 (N_17746,N_17526,N_17459);
nor U17747 (N_17747,N_17471,N_17512);
or U17748 (N_17748,N_17540,N_17465);
nor U17749 (N_17749,N_17494,N_17558);
nor U17750 (N_17750,N_17498,N_17551);
nand U17751 (N_17751,N_17584,N_17592);
nor U17752 (N_17752,N_17441,N_17532);
xnor U17753 (N_17753,N_17513,N_17526);
and U17754 (N_17754,N_17578,N_17591);
and U17755 (N_17755,N_17441,N_17442);
xnor U17756 (N_17756,N_17470,N_17448);
and U17757 (N_17757,N_17474,N_17493);
nand U17758 (N_17758,N_17576,N_17572);
nand U17759 (N_17759,N_17597,N_17488);
or U17760 (N_17760,N_17669,N_17690);
and U17761 (N_17761,N_17677,N_17665);
and U17762 (N_17762,N_17718,N_17613);
or U17763 (N_17763,N_17643,N_17639);
and U17764 (N_17764,N_17619,N_17750);
nor U17765 (N_17765,N_17658,N_17603);
xnor U17766 (N_17766,N_17663,N_17615);
and U17767 (N_17767,N_17701,N_17736);
nand U17768 (N_17768,N_17621,N_17753);
nand U17769 (N_17769,N_17654,N_17749);
xor U17770 (N_17770,N_17723,N_17726);
and U17771 (N_17771,N_17634,N_17672);
nor U17772 (N_17772,N_17644,N_17678);
and U17773 (N_17773,N_17693,N_17631);
xor U17774 (N_17774,N_17670,N_17671);
or U17775 (N_17775,N_17687,N_17704);
and U17776 (N_17776,N_17675,N_17695);
or U17777 (N_17777,N_17661,N_17752);
nor U17778 (N_17778,N_17630,N_17698);
nand U17779 (N_17779,N_17689,N_17744);
xnor U17780 (N_17780,N_17612,N_17739);
and U17781 (N_17781,N_17728,N_17700);
and U17782 (N_17782,N_17746,N_17651);
nand U17783 (N_17783,N_17696,N_17721);
nor U17784 (N_17784,N_17722,N_17601);
nand U17785 (N_17785,N_17636,N_17679);
xor U17786 (N_17786,N_17712,N_17714);
xnor U17787 (N_17787,N_17743,N_17727);
nor U17788 (N_17788,N_17691,N_17650);
nand U17789 (N_17789,N_17606,N_17640);
or U17790 (N_17790,N_17666,N_17686);
or U17791 (N_17791,N_17681,N_17662);
xor U17792 (N_17792,N_17664,N_17713);
or U17793 (N_17793,N_17759,N_17637);
and U17794 (N_17794,N_17667,N_17625);
xor U17795 (N_17795,N_17688,N_17729);
nor U17796 (N_17796,N_17755,N_17649);
nand U17797 (N_17797,N_17605,N_17600);
xnor U17798 (N_17798,N_17706,N_17748);
nor U17799 (N_17799,N_17707,N_17633);
nand U17800 (N_17800,N_17638,N_17699);
nand U17801 (N_17801,N_17610,N_17705);
xor U17802 (N_17802,N_17674,N_17646);
nor U17803 (N_17803,N_17611,N_17604);
nand U17804 (N_17804,N_17641,N_17738);
or U17805 (N_17805,N_17608,N_17692);
or U17806 (N_17806,N_17632,N_17660);
xor U17807 (N_17807,N_17628,N_17754);
nor U17808 (N_17808,N_17708,N_17653);
nor U17809 (N_17809,N_17709,N_17684);
xor U17810 (N_17810,N_17673,N_17626);
xnor U17811 (N_17811,N_17609,N_17710);
and U17812 (N_17812,N_17756,N_17694);
or U17813 (N_17813,N_17607,N_17624);
xor U17814 (N_17814,N_17740,N_17733);
and U17815 (N_17815,N_17745,N_17620);
xnor U17816 (N_17816,N_17724,N_17623);
nor U17817 (N_17817,N_17703,N_17741);
or U17818 (N_17818,N_17676,N_17648);
xnor U17819 (N_17819,N_17751,N_17657);
and U17820 (N_17820,N_17719,N_17725);
and U17821 (N_17821,N_17737,N_17685);
and U17822 (N_17822,N_17735,N_17711);
nor U17823 (N_17823,N_17682,N_17702);
nor U17824 (N_17824,N_17731,N_17717);
and U17825 (N_17825,N_17616,N_17720);
and U17826 (N_17826,N_17652,N_17683);
and U17827 (N_17827,N_17716,N_17642);
or U17828 (N_17828,N_17730,N_17635);
nor U17829 (N_17829,N_17680,N_17617);
or U17830 (N_17830,N_17659,N_17655);
or U17831 (N_17831,N_17618,N_17656);
and U17832 (N_17832,N_17602,N_17742);
xnor U17833 (N_17833,N_17668,N_17647);
nand U17834 (N_17834,N_17645,N_17734);
nor U17835 (N_17835,N_17747,N_17622);
nand U17836 (N_17836,N_17627,N_17757);
nor U17837 (N_17837,N_17614,N_17697);
xor U17838 (N_17838,N_17732,N_17629);
xor U17839 (N_17839,N_17758,N_17715);
or U17840 (N_17840,N_17671,N_17636);
and U17841 (N_17841,N_17712,N_17702);
and U17842 (N_17842,N_17719,N_17608);
nand U17843 (N_17843,N_17656,N_17634);
or U17844 (N_17844,N_17665,N_17755);
nand U17845 (N_17845,N_17697,N_17624);
or U17846 (N_17846,N_17619,N_17661);
nand U17847 (N_17847,N_17617,N_17666);
or U17848 (N_17848,N_17656,N_17725);
nand U17849 (N_17849,N_17621,N_17755);
nand U17850 (N_17850,N_17611,N_17671);
nor U17851 (N_17851,N_17642,N_17647);
xnor U17852 (N_17852,N_17704,N_17654);
nand U17853 (N_17853,N_17697,N_17661);
nand U17854 (N_17854,N_17705,N_17642);
xnor U17855 (N_17855,N_17671,N_17624);
xor U17856 (N_17856,N_17692,N_17758);
xnor U17857 (N_17857,N_17643,N_17748);
or U17858 (N_17858,N_17737,N_17628);
or U17859 (N_17859,N_17697,N_17690);
nor U17860 (N_17860,N_17732,N_17658);
and U17861 (N_17861,N_17745,N_17757);
nor U17862 (N_17862,N_17692,N_17700);
xor U17863 (N_17863,N_17697,N_17743);
nor U17864 (N_17864,N_17607,N_17676);
and U17865 (N_17865,N_17702,N_17725);
nor U17866 (N_17866,N_17727,N_17630);
xnor U17867 (N_17867,N_17710,N_17656);
or U17868 (N_17868,N_17636,N_17756);
or U17869 (N_17869,N_17715,N_17619);
xor U17870 (N_17870,N_17711,N_17662);
and U17871 (N_17871,N_17688,N_17719);
xor U17872 (N_17872,N_17705,N_17648);
nand U17873 (N_17873,N_17687,N_17665);
xnor U17874 (N_17874,N_17717,N_17601);
xnor U17875 (N_17875,N_17608,N_17652);
and U17876 (N_17876,N_17650,N_17627);
or U17877 (N_17877,N_17704,N_17667);
nand U17878 (N_17878,N_17643,N_17753);
nand U17879 (N_17879,N_17718,N_17627);
or U17880 (N_17880,N_17696,N_17735);
nor U17881 (N_17881,N_17739,N_17747);
nor U17882 (N_17882,N_17638,N_17686);
or U17883 (N_17883,N_17657,N_17629);
nand U17884 (N_17884,N_17739,N_17605);
nor U17885 (N_17885,N_17691,N_17608);
nor U17886 (N_17886,N_17661,N_17737);
and U17887 (N_17887,N_17669,N_17685);
nand U17888 (N_17888,N_17684,N_17698);
and U17889 (N_17889,N_17619,N_17723);
xnor U17890 (N_17890,N_17636,N_17739);
or U17891 (N_17891,N_17642,N_17633);
and U17892 (N_17892,N_17738,N_17666);
nand U17893 (N_17893,N_17628,N_17615);
xnor U17894 (N_17894,N_17709,N_17633);
and U17895 (N_17895,N_17607,N_17642);
nand U17896 (N_17896,N_17659,N_17728);
xor U17897 (N_17897,N_17622,N_17689);
or U17898 (N_17898,N_17675,N_17604);
or U17899 (N_17899,N_17641,N_17617);
xnor U17900 (N_17900,N_17603,N_17679);
or U17901 (N_17901,N_17604,N_17615);
xor U17902 (N_17902,N_17717,N_17662);
or U17903 (N_17903,N_17679,N_17729);
nand U17904 (N_17904,N_17743,N_17652);
nor U17905 (N_17905,N_17736,N_17751);
nor U17906 (N_17906,N_17656,N_17627);
and U17907 (N_17907,N_17633,N_17732);
nand U17908 (N_17908,N_17667,N_17663);
xnor U17909 (N_17909,N_17729,N_17757);
xnor U17910 (N_17910,N_17634,N_17657);
nor U17911 (N_17911,N_17700,N_17686);
and U17912 (N_17912,N_17731,N_17617);
nor U17913 (N_17913,N_17625,N_17656);
nand U17914 (N_17914,N_17720,N_17730);
nor U17915 (N_17915,N_17705,N_17600);
xor U17916 (N_17916,N_17630,N_17728);
and U17917 (N_17917,N_17754,N_17713);
and U17918 (N_17918,N_17751,N_17705);
and U17919 (N_17919,N_17753,N_17697);
xor U17920 (N_17920,N_17764,N_17821);
and U17921 (N_17921,N_17866,N_17762);
nand U17922 (N_17922,N_17849,N_17886);
xnor U17923 (N_17923,N_17915,N_17855);
nand U17924 (N_17924,N_17803,N_17781);
or U17925 (N_17925,N_17818,N_17847);
and U17926 (N_17926,N_17868,N_17913);
nor U17927 (N_17927,N_17899,N_17771);
nor U17928 (N_17928,N_17840,N_17844);
and U17929 (N_17929,N_17894,N_17869);
xor U17930 (N_17930,N_17763,N_17862);
or U17931 (N_17931,N_17768,N_17906);
nand U17932 (N_17932,N_17895,N_17856);
and U17933 (N_17933,N_17772,N_17810);
or U17934 (N_17934,N_17777,N_17882);
nand U17935 (N_17935,N_17871,N_17808);
or U17936 (N_17936,N_17831,N_17864);
nor U17937 (N_17937,N_17826,N_17907);
and U17938 (N_17938,N_17800,N_17825);
xnor U17939 (N_17939,N_17767,N_17900);
xor U17940 (N_17940,N_17910,N_17873);
xor U17941 (N_17941,N_17850,N_17795);
and U17942 (N_17942,N_17893,N_17784);
and U17943 (N_17943,N_17901,N_17828);
nor U17944 (N_17944,N_17793,N_17766);
nor U17945 (N_17945,N_17919,N_17911);
xnor U17946 (N_17946,N_17878,N_17872);
or U17947 (N_17947,N_17852,N_17885);
xor U17948 (N_17948,N_17880,N_17916);
nor U17949 (N_17949,N_17807,N_17813);
or U17950 (N_17950,N_17820,N_17833);
xor U17951 (N_17951,N_17838,N_17897);
nand U17952 (N_17952,N_17814,N_17794);
nand U17953 (N_17953,N_17775,N_17822);
xor U17954 (N_17954,N_17827,N_17799);
nor U17955 (N_17955,N_17791,N_17829);
xnor U17956 (N_17956,N_17909,N_17785);
and U17957 (N_17957,N_17917,N_17816);
nor U17958 (N_17958,N_17760,N_17787);
xor U17959 (N_17959,N_17790,N_17857);
and U17960 (N_17960,N_17765,N_17903);
xnor U17961 (N_17961,N_17902,N_17843);
nand U17962 (N_17962,N_17780,N_17783);
xnor U17963 (N_17963,N_17892,N_17789);
nand U17964 (N_17964,N_17835,N_17858);
or U17965 (N_17965,N_17788,N_17842);
or U17966 (N_17966,N_17904,N_17802);
nor U17967 (N_17967,N_17770,N_17837);
nor U17968 (N_17968,N_17786,N_17854);
nand U17969 (N_17969,N_17841,N_17774);
nand U17970 (N_17970,N_17839,N_17881);
and U17971 (N_17971,N_17846,N_17798);
nand U17972 (N_17972,N_17811,N_17806);
or U17973 (N_17973,N_17853,N_17801);
or U17974 (N_17974,N_17809,N_17863);
and U17975 (N_17975,N_17823,N_17817);
or U17976 (N_17976,N_17890,N_17805);
xnor U17977 (N_17977,N_17874,N_17834);
xor U17978 (N_17978,N_17832,N_17815);
xor U17979 (N_17979,N_17888,N_17761);
xnor U17980 (N_17980,N_17865,N_17796);
or U17981 (N_17981,N_17884,N_17877);
xnor U17982 (N_17982,N_17879,N_17848);
xor U17983 (N_17983,N_17887,N_17797);
nand U17984 (N_17984,N_17883,N_17860);
and U17985 (N_17985,N_17792,N_17804);
nand U17986 (N_17986,N_17769,N_17836);
nor U17987 (N_17987,N_17889,N_17908);
or U17988 (N_17988,N_17896,N_17867);
nand U17989 (N_17989,N_17830,N_17861);
and U17990 (N_17990,N_17905,N_17891);
nor U17991 (N_17991,N_17776,N_17851);
or U17992 (N_17992,N_17859,N_17875);
nand U17993 (N_17993,N_17773,N_17914);
nand U17994 (N_17994,N_17819,N_17779);
or U17995 (N_17995,N_17912,N_17845);
or U17996 (N_17996,N_17824,N_17778);
or U17997 (N_17997,N_17918,N_17898);
xnor U17998 (N_17998,N_17870,N_17812);
or U17999 (N_17999,N_17782,N_17876);
nand U18000 (N_18000,N_17909,N_17840);
nand U18001 (N_18001,N_17904,N_17850);
or U18002 (N_18002,N_17884,N_17792);
nor U18003 (N_18003,N_17891,N_17799);
and U18004 (N_18004,N_17796,N_17768);
nand U18005 (N_18005,N_17828,N_17790);
and U18006 (N_18006,N_17791,N_17871);
nor U18007 (N_18007,N_17855,N_17890);
xnor U18008 (N_18008,N_17888,N_17780);
nor U18009 (N_18009,N_17904,N_17827);
nor U18010 (N_18010,N_17792,N_17904);
nor U18011 (N_18011,N_17906,N_17893);
nor U18012 (N_18012,N_17898,N_17820);
and U18013 (N_18013,N_17797,N_17799);
nor U18014 (N_18014,N_17862,N_17873);
xnor U18015 (N_18015,N_17897,N_17907);
and U18016 (N_18016,N_17844,N_17762);
or U18017 (N_18017,N_17882,N_17783);
or U18018 (N_18018,N_17890,N_17799);
nand U18019 (N_18019,N_17915,N_17892);
and U18020 (N_18020,N_17909,N_17873);
or U18021 (N_18021,N_17875,N_17905);
xnor U18022 (N_18022,N_17853,N_17844);
nor U18023 (N_18023,N_17765,N_17889);
nand U18024 (N_18024,N_17836,N_17900);
or U18025 (N_18025,N_17765,N_17857);
or U18026 (N_18026,N_17775,N_17774);
or U18027 (N_18027,N_17841,N_17799);
nand U18028 (N_18028,N_17878,N_17868);
xnor U18029 (N_18029,N_17908,N_17841);
nor U18030 (N_18030,N_17915,N_17913);
nand U18031 (N_18031,N_17837,N_17901);
xnor U18032 (N_18032,N_17838,N_17794);
nor U18033 (N_18033,N_17792,N_17887);
and U18034 (N_18034,N_17832,N_17818);
nand U18035 (N_18035,N_17822,N_17837);
nand U18036 (N_18036,N_17853,N_17815);
or U18037 (N_18037,N_17874,N_17907);
xnor U18038 (N_18038,N_17779,N_17815);
xor U18039 (N_18039,N_17762,N_17793);
or U18040 (N_18040,N_17805,N_17798);
nor U18041 (N_18041,N_17779,N_17902);
and U18042 (N_18042,N_17781,N_17860);
nand U18043 (N_18043,N_17900,N_17788);
nand U18044 (N_18044,N_17902,N_17770);
nor U18045 (N_18045,N_17763,N_17818);
and U18046 (N_18046,N_17760,N_17840);
nand U18047 (N_18047,N_17786,N_17860);
or U18048 (N_18048,N_17839,N_17763);
and U18049 (N_18049,N_17815,N_17879);
or U18050 (N_18050,N_17760,N_17798);
nor U18051 (N_18051,N_17870,N_17770);
and U18052 (N_18052,N_17862,N_17832);
and U18053 (N_18053,N_17859,N_17869);
and U18054 (N_18054,N_17874,N_17896);
nand U18055 (N_18055,N_17822,N_17798);
or U18056 (N_18056,N_17861,N_17856);
nor U18057 (N_18057,N_17799,N_17824);
nor U18058 (N_18058,N_17800,N_17829);
or U18059 (N_18059,N_17792,N_17800);
xor U18060 (N_18060,N_17774,N_17860);
nor U18061 (N_18061,N_17835,N_17902);
nor U18062 (N_18062,N_17842,N_17847);
nand U18063 (N_18063,N_17873,N_17827);
nor U18064 (N_18064,N_17786,N_17880);
or U18065 (N_18065,N_17792,N_17862);
xor U18066 (N_18066,N_17783,N_17824);
nand U18067 (N_18067,N_17805,N_17775);
and U18068 (N_18068,N_17782,N_17826);
or U18069 (N_18069,N_17809,N_17915);
nand U18070 (N_18070,N_17890,N_17763);
nor U18071 (N_18071,N_17826,N_17764);
xnor U18072 (N_18072,N_17825,N_17902);
xnor U18073 (N_18073,N_17857,N_17859);
xnor U18074 (N_18074,N_17825,N_17824);
and U18075 (N_18075,N_17912,N_17833);
and U18076 (N_18076,N_17774,N_17869);
nor U18077 (N_18077,N_17802,N_17899);
nor U18078 (N_18078,N_17828,N_17916);
nand U18079 (N_18079,N_17780,N_17851);
nor U18080 (N_18080,N_17969,N_18060);
and U18081 (N_18081,N_18001,N_17963);
xnor U18082 (N_18082,N_17943,N_18000);
nor U18083 (N_18083,N_17995,N_17993);
xor U18084 (N_18084,N_18030,N_17933);
or U18085 (N_18085,N_18061,N_18033);
nand U18086 (N_18086,N_17994,N_17981);
or U18087 (N_18087,N_17928,N_17959);
nand U18088 (N_18088,N_17951,N_17949);
nor U18089 (N_18089,N_18055,N_17942);
nor U18090 (N_18090,N_18020,N_18063);
xor U18091 (N_18091,N_18023,N_18065);
xor U18092 (N_18092,N_17996,N_17975);
or U18093 (N_18093,N_18044,N_17992);
or U18094 (N_18094,N_18064,N_18039);
or U18095 (N_18095,N_17970,N_18042);
and U18096 (N_18096,N_18037,N_17956);
and U18097 (N_18097,N_17997,N_17998);
nand U18098 (N_18098,N_18051,N_18017);
nand U18099 (N_18099,N_18045,N_18046);
nand U18100 (N_18100,N_17989,N_18029);
nand U18101 (N_18101,N_17920,N_17973);
or U18102 (N_18102,N_17924,N_17954);
or U18103 (N_18103,N_18015,N_17988);
or U18104 (N_18104,N_17983,N_17965);
and U18105 (N_18105,N_17932,N_18057);
xnor U18106 (N_18106,N_17971,N_17958);
and U18107 (N_18107,N_17950,N_18040);
nand U18108 (N_18108,N_17944,N_18066);
or U18109 (N_18109,N_18010,N_18048);
xor U18110 (N_18110,N_18011,N_18073);
or U18111 (N_18111,N_17936,N_17957);
nor U18112 (N_18112,N_17940,N_17964);
xor U18113 (N_18113,N_18006,N_17922);
xnor U18114 (N_18114,N_18019,N_18034);
xor U18115 (N_18115,N_18075,N_18069);
nor U18116 (N_18116,N_18018,N_18043);
xor U18117 (N_18117,N_18071,N_17953);
nor U18118 (N_18118,N_18013,N_17972);
or U18119 (N_18119,N_18002,N_18012);
nor U18120 (N_18120,N_18021,N_18028);
and U18121 (N_18121,N_17999,N_17927);
and U18122 (N_18122,N_18059,N_18009);
nor U18123 (N_18123,N_18036,N_17968);
or U18124 (N_18124,N_17986,N_18050);
or U18125 (N_18125,N_17925,N_17974);
and U18126 (N_18126,N_18031,N_18041);
and U18127 (N_18127,N_17923,N_17955);
nand U18128 (N_18128,N_17979,N_17952);
xor U18129 (N_18129,N_18022,N_17977);
xor U18130 (N_18130,N_17938,N_18027);
nor U18131 (N_18131,N_18068,N_18062);
nor U18132 (N_18132,N_18008,N_17991);
or U18133 (N_18133,N_17980,N_17931);
or U18134 (N_18134,N_18078,N_18058);
xor U18135 (N_18135,N_18072,N_17990);
nand U18136 (N_18136,N_18049,N_18035);
nand U18137 (N_18137,N_17930,N_18025);
xor U18138 (N_18138,N_17929,N_17939);
or U18139 (N_18139,N_18032,N_17962);
and U18140 (N_18140,N_17945,N_17967);
or U18141 (N_18141,N_18052,N_17984);
nor U18142 (N_18142,N_18014,N_17941);
xnor U18143 (N_18143,N_17947,N_18024);
or U18144 (N_18144,N_18067,N_17976);
nand U18145 (N_18145,N_17960,N_18074);
nor U18146 (N_18146,N_18076,N_17987);
and U18147 (N_18147,N_18038,N_17985);
and U18148 (N_18148,N_18016,N_17921);
nand U18149 (N_18149,N_18054,N_18007);
nand U18150 (N_18150,N_18005,N_17946);
nor U18151 (N_18151,N_17934,N_17937);
nor U18152 (N_18152,N_17961,N_18004);
and U18153 (N_18153,N_17926,N_17966);
nand U18154 (N_18154,N_18053,N_17982);
nor U18155 (N_18155,N_18077,N_18047);
and U18156 (N_18156,N_18026,N_17935);
nand U18157 (N_18157,N_18056,N_17978);
nand U18158 (N_18158,N_17948,N_18003);
and U18159 (N_18159,N_18079,N_18070);
xor U18160 (N_18160,N_17951,N_17952);
or U18161 (N_18161,N_17949,N_18028);
nor U18162 (N_18162,N_17985,N_17991);
or U18163 (N_18163,N_18065,N_17962);
or U18164 (N_18164,N_17930,N_17964);
and U18165 (N_18165,N_17983,N_17924);
nor U18166 (N_18166,N_18063,N_17979);
or U18167 (N_18167,N_17933,N_17980);
and U18168 (N_18168,N_17981,N_17985);
nor U18169 (N_18169,N_18032,N_17978);
and U18170 (N_18170,N_18066,N_18021);
or U18171 (N_18171,N_18008,N_17983);
or U18172 (N_18172,N_18076,N_18038);
or U18173 (N_18173,N_17928,N_17935);
and U18174 (N_18174,N_18040,N_18046);
and U18175 (N_18175,N_17926,N_18017);
or U18176 (N_18176,N_18012,N_18054);
nand U18177 (N_18177,N_17937,N_18056);
or U18178 (N_18178,N_18000,N_18012);
or U18179 (N_18179,N_17989,N_17933);
and U18180 (N_18180,N_18013,N_17937);
nand U18181 (N_18181,N_17924,N_18052);
xor U18182 (N_18182,N_17997,N_18055);
and U18183 (N_18183,N_18041,N_17939);
nor U18184 (N_18184,N_18041,N_17958);
nand U18185 (N_18185,N_18007,N_18023);
nor U18186 (N_18186,N_18022,N_18013);
nand U18187 (N_18187,N_17946,N_18048);
nand U18188 (N_18188,N_18071,N_18060);
and U18189 (N_18189,N_18079,N_17974);
xnor U18190 (N_18190,N_17982,N_17947);
nand U18191 (N_18191,N_17939,N_17955);
and U18192 (N_18192,N_17985,N_18056);
nor U18193 (N_18193,N_18015,N_18069);
nor U18194 (N_18194,N_18055,N_17928);
xor U18195 (N_18195,N_17932,N_18000);
or U18196 (N_18196,N_17991,N_17971);
nor U18197 (N_18197,N_18029,N_18046);
or U18198 (N_18198,N_17927,N_18010);
or U18199 (N_18199,N_17947,N_17944);
nand U18200 (N_18200,N_18000,N_17969);
and U18201 (N_18201,N_18067,N_17953);
nand U18202 (N_18202,N_18002,N_18019);
or U18203 (N_18203,N_18077,N_17953);
xnor U18204 (N_18204,N_18058,N_18074);
nand U18205 (N_18205,N_18038,N_17978);
nand U18206 (N_18206,N_18040,N_17956);
or U18207 (N_18207,N_18040,N_18060);
or U18208 (N_18208,N_17987,N_18022);
nand U18209 (N_18209,N_18050,N_17959);
nor U18210 (N_18210,N_18058,N_17970);
nor U18211 (N_18211,N_17982,N_18054);
and U18212 (N_18212,N_17938,N_17957);
or U18213 (N_18213,N_18006,N_18076);
and U18214 (N_18214,N_18048,N_18062);
xnor U18215 (N_18215,N_18054,N_18047);
nor U18216 (N_18216,N_17928,N_17974);
or U18217 (N_18217,N_17975,N_18045);
or U18218 (N_18218,N_18022,N_18065);
nor U18219 (N_18219,N_18021,N_18054);
and U18220 (N_18220,N_18008,N_17953);
nor U18221 (N_18221,N_18062,N_17995);
nor U18222 (N_18222,N_17939,N_17966);
and U18223 (N_18223,N_18062,N_17973);
and U18224 (N_18224,N_18019,N_18036);
xnor U18225 (N_18225,N_18016,N_18027);
nor U18226 (N_18226,N_17954,N_17990);
or U18227 (N_18227,N_17966,N_18049);
or U18228 (N_18228,N_18027,N_18068);
nand U18229 (N_18229,N_18005,N_17992);
nand U18230 (N_18230,N_18039,N_18047);
and U18231 (N_18231,N_18007,N_18009);
nand U18232 (N_18232,N_17988,N_17935);
and U18233 (N_18233,N_18032,N_17966);
and U18234 (N_18234,N_17962,N_17922);
or U18235 (N_18235,N_17939,N_17977);
and U18236 (N_18236,N_18059,N_17983);
nand U18237 (N_18237,N_17950,N_18028);
nand U18238 (N_18238,N_18034,N_17993);
xnor U18239 (N_18239,N_18054,N_18015);
nand U18240 (N_18240,N_18210,N_18105);
and U18241 (N_18241,N_18202,N_18190);
nand U18242 (N_18242,N_18086,N_18147);
or U18243 (N_18243,N_18082,N_18204);
xor U18244 (N_18244,N_18239,N_18191);
and U18245 (N_18245,N_18101,N_18115);
or U18246 (N_18246,N_18169,N_18158);
xnor U18247 (N_18247,N_18194,N_18126);
or U18248 (N_18248,N_18174,N_18176);
nor U18249 (N_18249,N_18220,N_18123);
and U18250 (N_18250,N_18128,N_18094);
and U18251 (N_18251,N_18118,N_18165);
nand U18252 (N_18252,N_18233,N_18138);
nor U18253 (N_18253,N_18163,N_18142);
and U18254 (N_18254,N_18208,N_18121);
or U18255 (N_18255,N_18183,N_18155);
nor U18256 (N_18256,N_18226,N_18170);
nor U18257 (N_18257,N_18135,N_18122);
nor U18258 (N_18258,N_18237,N_18196);
xnor U18259 (N_18259,N_18185,N_18132);
nand U18260 (N_18260,N_18108,N_18186);
nor U18261 (N_18261,N_18168,N_18110);
nor U18262 (N_18262,N_18205,N_18144);
and U18263 (N_18263,N_18230,N_18154);
or U18264 (N_18264,N_18234,N_18187);
nor U18265 (N_18265,N_18216,N_18227);
xnor U18266 (N_18266,N_18112,N_18189);
xnor U18267 (N_18267,N_18206,N_18146);
xnor U18268 (N_18268,N_18218,N_18229);
and U18269 (N_18269,N_18085,N_18087);
nor U18270 (N_18270,N_18192,N_18203);
nor U18271 (N_18271,N_18219,N_18116);
and U18272 (N_18272,N_18214,N_18106);
or U18273 (N_18273,N_18084,N_18137);
nand U18274 (N_18274,N_18093,N_18175);
and U18275 (N_18275,N_18199,N_18179);
or U18276 (N_18276,N_18207,N_18130);
xnor U18277 (N_18277,N_18188,N_18092);
and U18278 (N_18278,N_18197,N_18172);
xnor U18279 (N_18279,N_18222,N_18117);
nor U18280 (N_18280,N_18091,N_18151);
xor U18281 (N_18281,N_18134,N_18193);
xor U18282 (N_18282,N_18145,N_18127);
and U18283 (N_18283,N_18136,N_18152);
nor U18284 (N_18284,N_18097,N_18088);
or U18285 (N_18285,N_18111,N_18232);
and U18286 (N_18286,N_18164,N_18236);
or U18287 (N_18287,N_18177,N_18180);
nor U18288 (N_18288,N_18156,N_18181);
xor U18289 (N_18289,N_18223,N_18109);
nor U18290 (N_18290,N_18178,N_18139);
nand U18291 (N_18291,N_18213,N_18125);
or U18292 (N_18292,N_18159,N_18184);
and U18293 (N_18293,N_18090,N_18238);
nand U18294 (N_18294,N_18149,N_18166);
or U18295 (N_18295,N_18173,N_18160);
nand U18296 (N_18296,N_18198,N_18133);
nor U18297 (N_18297,N_18102,N_18215);
xnor U18298 (N_18298,N_18221,N_18200);
nand U18299 (N_18299,N_18129,N_18182);
xor U18300 (N_18300,N_18148,N_18161);
nand U18301 (N_18301,N_18114,N_18098);
and U18302 (N_18302,N_18089,N_18150);
or U18303 (N_18303,N_18201,N_18095);
xor U18304 (N_18304,N_18235,N_18195);
nand U18305 (N_18305,N_18113,N_18104);
xor U18306 (N_18306,N_18157,N_18224);
or U18307 (N_18307,N_18228,N_18100);
and U18308 (N_18308,N_18211,N_18083);
and U18309 (N_18309,N_18225,N_18096);
nand U18310 (N_18310,N_18153,N_18171);
and U18311 (N_18311,N_18143,N_18119);
or U18312 (N_18312,N_18162,N_18212);
nor U18313 (N_18313,N_18107,N_18120);
nand U18314 (N_18314,N_18131,N_18081);
and U18315 (N_18315,N_18167,N_18080);
xnor U18316 (N_18316,N_18217,N_18141);
xnor U18317 (N_18317,N_18231,N_18209);
and U18318 (N_18318,N_18099,N_18103);
or U18319 (N_18319,N_18140,N_18124);
nand U18320 (N_18320,N_18140,N_18192);
nand U18321 (N_18321,N_18238,N_18218);
and U18322 (N_18322,N_18236,N_18215);
nor U18323 (N_18323,N_18202,N_18118);
nand U18324 (N_18324,N_18182,N_18146);
and U18325 (N_18325,N_18205,N_18172);
and U18326 (N_18326,N_18204,N_18113);
or U18327 (N_18327,N_18232,N_18128);
and U18328 (N_18328,N_18183,N_18199);
xnor U18329 (N_18329,N_18082,N_18087);
nand U18330 (N_18330,N_18123,N_18141);
nor U18331 (N_18331,N_18144,N_18115);
or U18332 (N_18332,N_18201,N_18224);
nand U18333 (N_18333,N_18114,N_18200);
or U18334 (N_18334,N_18111,N_18219);
nand U18335 (N_18335,N_18223,N_18165);
xnor U18336 (N_18336,N_18119,N_18220);
nand U18337 (N_18337,N_18100,N_18171);
and U18338 (N_18338,N_18183,N_18140);
nor U18339 (N_18339,N_18229,N_18105);
nor U18340 (N_18340,N_18123,N_18207);
nand U18341 (N_18341,N_18112,N_18153);
or U18342 (N_18342,N_18237,N_18206);
nor U18343 (N_18343,N_18150,N_18098);
xor U18344 (N_18344,N_18195,N_18222);
xor U18345 (N_18345,N_18142,N_18194);
nor U18346 (N_18346,N_18144,N_18127);
nand U18347 (N_18347,N_18135,N_18229);
or U18348 (N_18348,N_18096,N_18208);
and U18349 (N_18349,N_18095,N_18120);
xor U18350 (N_18350,N_18164,N_18224);
nor U18351 (N_18351,N_18200,N_18102);
and U18352 (N_18352,N_18158,N_18192);
and U18353 (N_18353,N_18209,N_18182);
nand U18354 (N_18354,N_18203,N_18087);
and U18355 (N_18355,N_18186,N_18227);
nor U18356 (N_18356,N_18207,N_18214);
nor U18357 (N_18357,N_18116,N_18236);
or U18358 (N_18358,N_18137,N_18152);
xnor U18359 (N_18359,N_18207,N_18202);
nand U18360 (N_18360,N_18193,N_18190);
and U18361 (N_18361,N_18118,N_18088);
nor U18362 (N_18362,N_18107,N_18134);
nand U18363 (N_18363,N_18155,N_18176);
nor U18364 (N_18364,N_18146,N_18108);
xnor U18365 (N_18365,N_18093,N_18107);
and U18366 (N_18366,N_18083,N_18188);
xnor U18367 (N_18367,N_18121,N_18187);
nand U18368 (N_18368,N_18154,N_18083);
or U18369 (N_18369,N_18103,N_18088);
and U18370 (N_18370,N_18092,N_18212);
nor U18371 (N_18371,N_18098,N_18234);
or U18372 (N_18372,N_18206,N_18236);
nand U18373 (N_18373,N_18107,N_18124);
nand U18374 (N_18374,N_18174,N_18113);
xnor U18375 (N_18375,N_18144,N_18212);
and U18376 (N_18376,N_18148,N_18151);
xor U18377 (N_18377,N_18235,N_18209);
and U18378 (N_18378,N_18120,N_18235);
xor U18379 (N_18379,N_18172,N_18084);
xnor U18380 (N_18380,N_18094,N_18100);
and U18381 (N_18381,N_18139,N_18146);
or U18382 (N_18382,N_18202,N_18083);
nand U18383 (N_18383,N_18199,N_18093);
nand U18384 (N_18384,N_18125,N_18134);
nand U18385 (N_18385,N_18166,N_18196);
nand U18386 (N_18386,N_18169,N_18218);
nor U18387 (N_18387,N_18217,N_18102);
nor U18388 (N_18388,N_18209,N_18214);
or U18389 (N_18389,N_18081,N_18187);
and U18390 (N_18390,N_18096,N_18237);
xor U18391 (N_18391,N_18209,N_18151);
xnor U18392 (N_18392,N_18228,N_18159);
nor U18393 (N_18393,N_18154,N_18112);
nand U18394 (N_18394,N_18209,N_18179);
or U18395 (N_18395,N_18130,N_18180);
or U18396 (N_18396,N_18145,N_18107);
nor U18397 (N_18397,N_18192,N_18223);
nand U18398 (N_18398,N_18232,N_18191);
nor U18399 (N_18399,N_18083,N_18089);
xnor U18400 (N_18400,N_18344,N_18271);
and U18401 (N_18401,N_18387,N_18252);
xor U18402 (N_18402,N_18308,N_18347);
and U18403 (N_18403,N_18327,N_18397);
or U18404 (N_18404,N_18357,N_18285);
nand U18405 (N_18405,N_18368,N_18288);
xnor U18406 (N_18406,N_18328,N_18376);
xor U18407 (N_18407,N_18241,N_18330);
and U18408 (N_18408,N_18307,N_18309);
nand U18409 (N_18409,N_18331,N_18295);
nor U18410 (N_18410,N_18398,N_18369);
or U18411 (N_18411,N_18379,N_18386);
nor U18412 (N_18412,N_18258,N_18270);
or U18413 (N_18413,N_18353,N_18313);
nand U18414 (N_18414,N_18374,N_18378);
or U18415 (N_18415,N_18390,N_18290);
nor U18416 (N_18416,N_18277,N_18247);
nor U18417 (N_18417,N_18272,N_18286);
nor U18418 (N_18418,N_18346,N_18391);
nor U18419 (N_18419,N_18292,N_18249);
and U18420 (N_18420,N_18370,N_18281);
xnor U18421 (N_18421,N_18282,N_18259);
or U18422 (N_18422,N_18382,N_18362);
nand U18423 (N_18423,N_18248,N_18299);
and U18424 (N_18424,N_18336,N_18296);
xor U18425 (N_18425,N_18337,N_18338);
and U18426 (N_18426,N_18396,N_18377);
xnor U18427 (N_18427,N_18312,N_18301);
and U18428 (N_18428,N_18303,N_18365);
nand U18429 (N_18429,N_18385,N_18373);
and U18430 (N_18430,N_18273,N_18367);
and U18431 (N_18431,N_18254,N_18334);
nor U18432 (N_18432,N_18371,N_18350);
or U18433 (N_18433,N_18359,N_18316);
nor U18434 (N_18434,N_18266,N_18304);
nand U18435 (N_18435,N_18279,N_18340);
xnor U18436 (N_18436,N_18323,N_18389);
xor U18437 (N_18437,N_18394,N_18264);
nand U18438 (N_18438,N_18375,N_18250);
nor U18439 (N_18439,N_18318,N_18294);
and U18440 (N_18440,N_18324,N_18320);
or U18441 (N_18441,N_18322,N_18268);
or U18442 (N_18442,N_18246,N_18306);
and U18443 (N_18443,N_18341,N_18399);
and U18444 (N_18444,N_18384,N_18319);
or U18445 (N_18445,N_18300,N_18356);
or U18446 (N_18446,N_18381,N_18329);
or U18447 (N_18447,N_18317,N_18363);
nor U18448 (N_18448,N_18343,N_18358);
xnor U18449 (N_18449,N_18260,N_18345);
nor U18450 (N_18450,N_18297,N_18364);
nor U18451 (N_18451,N_18335,N_18244);
nor U18452 (N_18452,N_18388,N_18253);
xnor U18453 (N_18453,N_18245,N_18242);
or U18454 (N_18454,N_18269,N_18298);
nand U18455 (N_18455,N_18314,N_18351);
or U18456 (N_18456,N_18257,N_18278);
or U18457 (N_18457,N_18325,N_18284);
and U18458 (N_18458,N_18276,N_18261);
or U18459 (N_18459,N_18289,N_18321);
xor U18460 (N_18460,N_18267,N_18348);
and U18461 (N_18461,N_18280,N_18310);
nand U18462 (N_18462,N_18291,N_18305);
nor U18463 (N_18463,N_18366,N_18360);
nor U18464 (N_18464,N_18240,N_18354);
xor U18465 (N_18465,N_18275,N_18383);
xor U18466 (N_18466,N_18255,N_18380);
and U18467 (N_18467,N_18311,N_18352);
xor U18468 (N_18468,N_18251,N_18274);
nand U18469 (N_18469,N_18339,N_18342);
xnor U18470 (N_18470,N_18355,N_18265);
or U18471 (N_18471,N_18395,N_18262);
and U18472 (N_18472,N_18333,N_18326);
and U18473 (N_18473,N_18361,N_18392);
or U18474 (N_18474,N_18263,N_18332);
nor U18475 (N_18475,N_18372,N_18393);
or U18476 (N_18476,N_18349,N_18283);
nand U18477 (N_18477,N_18287,N_18293);
and U18478 (N_18478,N_18302,N_18315);
nor U18479 (N_18479,N_18256,N_18243);
nor U18480 (N_18480,N_18263,N_18393);
and U18481 (N_18481,N_18250,N_18354);
xnor U18482 (N_18482,N_18373,N_18258);
or U18483 (N_18483,N_18368,N_18370);
and U18484 (N_18484,N_18362,N_18395);
xnor U18485 (N_18485,N_18391,N_18245);
nor U18486 (N_18486,N_18392,N_18323);
nand U18487 (N_18487,N_18288,N_18256);
xor U18488 (N_18488,N_18240,N_18322);
nand U18489 (N_18489,N_18298,N_18372);
and U18490 (N_18490,N_18297,N_18316);
nand U18491 (N_18491,N_18343,N_18242);
or U18492 (N_18492,N_18382,N_18377);
nor U18493 (N_18493,N_18328,N_18360);
nor U18494 (N_18494,N_18344,N_18336);
xor U18495 (N_18495,N_18271,N_18260);
or U18496 (N_18496,N_18384,N_18241);
nor U18497 (N_18497,N_18345,N_18300);
or U18498 (N_18498,N_18339,N_18303);
and U18499 (N_18499,N_18261,N_18350);
nand U18500 (N_18500,N_18382,N_18384);
nor U18501 (N_18501,N_18352,N_18340);
xor U18502 (N_18502,N_18262,N_18349);
nand U18503 (N_18503,N_18340,N_18388);
xor U18504 (N_18504,N_18346,N_18279);
and U18505 (N_18505,N_18382,N_18355);
nor U18506 (N_18506,N_18308,N_18358);
nor U18507 (N_18507,N_18375,N_18281);
and U18508 (N_18508,N_18240,N_18276);
xnor U18509 (N_18509,N_18350,N_18270);
xnor U18510 (N_18510,N_18330,N_18323);
nand U18511 (N_18511,N_18265,N_18370);
nor U18512 (N_18512,N_18391,N_18373);
or U18513 (N_18513,N_18391,N_18353);
nor U18514 (N_18514,N_18284,N_18337);
nor U18515 (N_18515,N_18319,N_18298);
xnor U18516 (N_18516,N_18298,N_18275);
xor U18517 (N_18517,N_18285,N_18319);
or U18518 (N_18518,N_18358,N_18299);
nor U18519 (N_18519,N_18288,N_18242);
nor U18520 (N_18520,N_18396,N_18318);
nand U18521 (N_18521,N_18325,N_18264);
xnor U18522 (N_18522,N_18351,N_18328);
xnor U18523 (N_18523,N_18285,N_18326);
nor U18524 (N_18524,N_18351,N_18363);
and U18525 (N_18525,N_18265,N_18308);
or U18526 (N_18526,N_18302,N_18244);
and U18527 (N_18527,N_18284,N_18311);
nor U18528 (N_18528,N_18279,N_18398);
or U18529 (N_18529,N_18244,N_18254);
nor U18530 (N_18530,N_18289,N_18367);
or U18531 (N_18531,N_18338,N_18330);
xnor U18532 (N_18532,N_18294,N_18349);
and U18533 (N_18533,N_18344,N_18323);
xnor U18534 (N_18534,N_18360,N_18362);
nand U18535 (N_18535,N_18341,N_18396);
xnor U18536 (N_18536,N_18310,N_18357);
or U18537 (N_18537,N_18367,N_18319);
nand U18538 (N_18538,N_18269,N_18377);
or U18539 (N_18539,N_18371,N_18328);
or U18540 (N_18540,N_18249,N_18366);
or U18541 (N_18541,N_18391,N_18291);
nor U18542 (N_18542,N_18292,N_18333);
and U18543 (N_18543,N_18356,N_18289);
and U18544 (N_18544,N_18376,N_18356);
nor U18545 (N_18545,N_18383,N_18302);
nand U18546 (N_18546,N_18268,N_18346);
or U18547 (N_18547,N_18381,N_18278);
xnor U18548 (N_18548,N_18279,N_18331);
nor U18549 (N_18549,N_18342,N_18349);
nor U18550 (N_18550,N_18286,N_18271);
or U18551 (N_18551,N_18310,N_18335);
xnor U18552 (N_18552,N_18387,N_18382);
xor U18553 (N_18553,N_18330,N_18374);
nand U18554 (N_18554,N_18288,N_18304);
and U18555 (N_18555,N_18326,N_18354);
or U18556 (N_18556,N_18284,N_18389);
or U18557 (N_18557,N_18316,N_18350);
nand U18558 (N_18558,N_18297,N_18337);
or U18559 (N_18559,N_18316,N_18337);
and U18560 (N_18560,N_18556,N_18537);
or U18561 (N_18561,N_18425,N_18431);
and U18562 (N_18562,N_18522,N_18553);
nand U18563 (N_18563,N_18492,N_18508);
xnor U18564 (N_18564,N_18460,N_18496);
xor U18565 (N_18565,N_18495,N_18410);
nor U18566 (N_18566,N_18472,N_18447);
or U18567 (N_18567,N_18533,N_18416);
xor U18568 (N_18568,N_18477,N_18517);
xor U18569 (N_18569,N_18407,N_18555);
xnor U18570 (N_18570,N_18421,N_18414);
xnor U18571 (N_18571,N_18549,N_18459);
xor U18572 (N_18572,N_18434,N_18551);
nor U18573 (N_18573,N_18475,N_18493);
nand U18574 (N_18574,N_18455,N_18461);
or U18575 (N_18575,N_18510,N_18498);
nor U18576 (N_18576,N_18526,N_18516);
xnor U18577 (N_18577,N_18506,N_18546);
or U18578 (N_18578,N_18535,N_18505);
nor U18579 (N_18579,N_18439,N_18543);
or U18580 (N_18580,N_18449,N_18423);
nor U18581 (N_18581,N_18524,N_18512);
xor U18582 (N_18582,N_18419,N_18465);
nand U18583 (N_18583,N_18415,N_18521);
and U18584 (N_18584,N_18507,N_18541);
and U18585 (N_18585,N_18446,N_18518);
nand U18586 (N_18586,N_18557,N_18443);
and U18587 (N_18587,N_18411,N_18474);
xor U18588 (N_18588,N_18404,N_18490);
and U18589 (N_18589,N_18432,N_18440);
nor U18590 (N_18590,N_18538,N_18473);
and U18591 (N_18591,N_18545,N_18457);
nand U18592 (N_18592,N_18400,N_18471);
nand U18593 (N_18593,N_18532,N_18509);
nand U18594 (N_18594,N_18540,N_18456);
xnor U18595 (N_18595,N_18435,N_18428);
nand U18596 (N_18596,N_18427,N_18453);
nand U18597 (N_18597,N_18534,N_18547);
and U18598 (N_18598,N_18408,N_18468);
nand U18599 (N_18599,N_18429,N_18478);
xor U18600 (N_18600,N_18463,N_18502);
nor U18601 (N_18601,N_18406,N_18485);
xnor U18602 (N_18602,N_18528,N_18504);
and U18603 (N_18603,N_18514,N_18479);
nor U18604 (N_18604,N_18501,N_18458);
or U18605 (N_18605,N_18402,N_18529);
and U18606 (N_18606,N_18466,N_18527);
and U18607 (N_18607,N_18470,N_18437);
nand U18608 (N_18608,N_18558,N_18464);
nor U18609 (N_18609,N_18536,N_18511);
or U18610 (N_18610,N_18523,N_18482);
nor U18611 (N_18611,N_18480,N_18424);
xor U18612 (N_18612,N_18539,N_18497);
or U18613 (N_18613,N_18452,N_18483);
nand U18614 (N_18614,N_18552,N_18418);
nand U18615 (N_18615,N_18488,N_18550);
xnor U18616 (N_18616,N_18548,N_18503);
nor U18617 (N_18617,N_18422,N_18476);
nand U18618 (N_18618,N_18417,N_18520);
or U18619 (N_18619,N_18467,N_18481);
or U18620 (N_18620,N_18525,N_18542);
or U18621 (N_18621,N_18420,N_18499);
nor U18622 (N_18622,N_18430,N_18489);
or U18623 (N_18623,N_18484,N_18559);
nor U18624 (N_18624,N_18450,N_18515);
xor U18625 (N_18625,N_18442,N_18426);
or U18626 (N_18626,N_18448,N_18469);
xor U18627 (N_18627,N_18462,N_18409);
xnor U18628 (N_18628,N_18513,N_18530);
or U18629 (N_18629,N_18500,N_18487);
or U18630 (N_18630,N_18519,N_18441);
or U18631 (N_18631,N_18486,N_18444);
nand U18632 (N_18632,N_18412,N_18454);
or U18633 (N_18633,N_18433,N_18554);
nand U18634 (N_18634,N_18438,N_18445);
and U18635 (N_18635,N_18413,N_18544);
nor U18636 (N_18636,N_18403,N_18451);
nor U18637 (N_18637,N_18531,N_18436);
or U18638 (N_18638,N_18405,N_18401);
nand U18639 (N_18639,N_18491,N_18494);
xnor U18640 (N_18640,N_18433,N_18530);
nand U18641 (N_18641,N_18453,N_18407);
nand U18642 (N_18642,N_18483,N_18427);
or U18643 (N_18643,N_18432,N_18449);
nor U18644 (N_18644,N_18438,N_18402);
xnor U18645 (N_18645,N_18433,N_18471);
or U18646 (N_18646,N_18465,N_18489);
xnor U18647 (N_18647,N_18440,N_18476);
or U18648 (N_18648,N_18426,N_18538);
or U18649 (N_18649,N_18443,N_18428);
nand U18650 (N_18650,N_18451,N_18443);
nand U18651 (N_18651,N_18474,N_18477);
xnor U18652 (N_18652,N_18409,N_18516);
xnor U18653 (N_18653,N_18518,N_18508);
nand U18654 (N_18654,N_18499,N_18402);
or U18655 (N_18655,N_18493,N_18436);
or U18656 (N_18656,N_18490,N_18531);
or U18657 (N_18657,N_18554,N_18551);
nor U18658 (N_18658,N_18401,N_18558);
and U18659 (N_18659,N_18435,N_18432);
nor U18660 (N_18660,N_18470,N_18431);
or U18661 (N_18661,N_18418,N_18547);
nor U18662 (N_18662,N_18475,N_18420);
nand U18663 (N_18663,N_18538,N_18405);
or U18664 (N_18664,N_18520,N_18419);
nand U18665 (N_18665,N_18488,N_18520);
xor U18666 (N_18666,N_18402,N_18541);
xnor U18667 (N_18667,N_18529,N_18460);
and U18668 (N_18668,N_18493,N_18439);
nand U18669 (N_18669,N_18502,N_18552);
xnor U18670 (N_18670,N_18509,N_18478);
or U18671 (N_18671,N_18544,N_18400);
xnor U18672 (N_18672,N_18435,N_18514);
and U18673 (N_18673,N_18423,N_18404);
xnor U18674 (N_18674,N_18448,N_18537);
nand U18675 (N_18675,N_18446,N_18536);
and U18676 (N_18676,N_18447,N_18513);
nand U18677 (N_18677,N_18420,N_18403);
nor U18678 (N_18678,N_18404,N_18496);
nand U18679 (N_18679,N_18470,N_18461);
or U18680 (N_18680,N_18453,N_18511);
and U18681 (N_18681,N_18527,N_18407);
xor U18682 (N_18682,N_18473,N_18438);
nor U18683 (N_18683,N_18459,N_18518);
nand U18684 (N_18684,N_18417,N_18522);
or U18685 (N_18685,N_18503,N_18434);
nor U18686 (N_18686,N_18414,N_18466);
nor U18687 (N_18687,N_18524,N_18518);
nand U18688 (N_18688,N_18407,N_18519);
or U18689 (N_18689,N_18489,N_18408);
nand U18690 (N_18690,N_18419,N_18526);
nand U18691 (N_18691,N_18509,N_18558);
or U18692 (N_18692,N_18555,N_18494);
and U18693 (N_18693,N_18417,N_18554);
nor U18694 (N_18694,N_18500,N_18551);
xnor U18695 (N_18695,N_18417,N_18416);
xnor U18696 (N_18696,N_18453,N_18499);
nor U18697 (N_18697,N_18417,N_18439);
or U18698 (N_18698,N_18487,N_18457);
and U18699 (N_18699,N_18466,N_18408);
nor U18700 (N_18700,N_18402,N_18497);
nor U18701 (N_18701,N_18418,N_18510);
or U18702 (N_18702,N_18473,N_18502);
and U18703 (N_18703,N_18511,N_18407);
and U18704 (N_18704,N_18401,N_18533);
nand U18705 (N_18705,N_18530,N_18519);
or U18706 (N_18706,N_18462,N_18495);
or U18707 (N_18707,N_18553,N_18536);
nor U18708 (N_18708,N_18474,N_18447);
nand U18709 (N_18709,N_18432,N_18522);
nand U18710 (N_18710,N_18548,N_18478);
nor U18711 (N_18711,N_18539,N_18409);
and U18712 (N_18712,N_18536,N_18465);
nand U18713 (N_18713,N_18490,N_18406);
nand U18714 (N_18714,N_18435,N_18520);
nor U18715 (N_18715,N_18430,N_18558);
nand U18716 (N_18716,N_18404,N_18412);
nor U18717 (N_18717,N_18524,N_18422);
nor U18718 (N_18718,N_18495,N_18530);
nor U18719 (N_18719,N_18529,N_18528);
nand U18720 (N_18720,N_18718,N_18628);
xor U18721 (N_18721,N_18614,N_18619);
xnor U18722 (N_18722,N_18711,N_18677);
xor U18723 (N_18723,N_18570,N_18686);
nand U18724 (N_18724,N_18562,N_18661);
nor U18725 (N_18725,N_18585,N_18712);
xor U18726 (N_18726,N_18567,N_18581);
xor U18727 (N_18727,N_18580,N_18583);
nor U18728 (N_18728,N_18589,N_18704);
nor U18729 (N_18729,N_18707,N_18702);
and U18730 (N_18730,N_18641,N_18605);
and U18731 (N_18731,N_18615,N_18633);
xnor U18732 (N_18732,N_18664,N_18660);
and U18733 (N_18733,N_18698,N_18595);
xnor U18734 (N_18734,N_18634,N_18577);
and U18735 (N_18735,N_18690,N_18651);
xor U18736 (N_18736,N_18561,N_18649);
nor U18737 (N_18737,N_18671,N_18688);
nor U18738 (N_18738,N_18719,N_18640);
or U18739 (N_18739,N_18574,N_18624);
nor U18740 (N_18740,N_18708,N_18679);
or U18741 (N_18741,N_18575,N_18608);
and U18742 (N_18742,N_18610,N_18683);
and U18743 (N_18743,N_18716,N_18710);
nand U18744 (N_18744,N_18714,N_18611);
nor U18745 (N_18745,N_18684,N_18672);
and U18746 (N_18746,N_18604,N_18693);
nand U18747 (N_18747,N_18616,N_18715);
xnor U18748 (N_18748,N_18652,N_18717);
and U18749 (N_18749,N_18673,N_18668);
or U18750 (N_18750,N_18586,N_18601);
nand U18751 (N_18751,N_18682,N_18568);
nor U18752 (N_18752,N_18689,N_18676);
or U18753 (N_18753,N_18643,N_18658);
nor U18754 (N_18754,N_18592,N_18630);
or U18755 (N_18755,N_18594,N_18560);
xnor U18756 (N_18756,N_18579,N_18588);
or U18757 (N_18757,N_18666,N_18587);
and U18758 (N_18758,N_18621,N_18697);
or U18759 (N_18759,N_18590,N_18636);
and U18760 (N_18760,N_18631,N_18687);
and U18761 (N_18761,N_18655,N_18646);
nand U18762 (N_18762,N_18653,N_18565);
nand U18763 (N_18763,N_18665,N_18596);
or U18764 (N_18764,N_18670,N_18569);
nor U18765 (N_18765,N_18618,N_18617);
nand U18766 (N_18766,N_18642,N_18662);
nor U18767 (N_18767,N_18602,N_18680);
and U18768 (N_18768,N_18627,N_18576);
and U18769 (N_18769,N_18656,N_18591);
nand U18770 (N_18770,N_18609,N_18696);
nand U18771 (N_18771,N_18667,N_18582);
or U18772 (N_18772,N_18564,N_18681);
or U18773 (N_18773,N_18600,N_18678);
nand U18774 (N_18774,N_18659,N_18571);
nor U18775 (N_18775,N_18572,N_18705);
and U18776 (N_18776,N_18637,N_18700);
and U18777 (N_18777,N_18623,N_18675);
and U18778 (N_18778,N_18573,N_18692);
and U18779 (N_18779,N_18645,N_18629);
nor U18780 (N_18780,N_18593,N_18644);
nor U18781 (N_18781,N_18691,N_18695);
and U18782 (N_18782,N_18635,N_18647);
nor U18783 (N_18783,N_18663,N_18657);
or U18784 (N_18784,N_18599,N_18578);
and U18785 (N_18785,N_18694,N_18607);
or U18786 (N_18786,N_18685,N_18612);
nand U18787 (N_18787,N_18626,N_18654);
and U18788 (N_18788,N_18669,N_18648);
or U18789 (N_18789,N_18597,N_18706);
and U18790 (N_18790,N_18709,N_18603);
xnor U18791 (N_18791,N_18639,N_18613);
or U18792 (N_18792,N_18713,N_18699);
nand U18793 (N_18793,N_18598,N_18622);
and U18794 (N_18794,N_18632,N_18563);
and U18795 (N_18795,N_18703,N_18625);
and U18796 (N_18796,N_18701,N_18584);
xnor U18797 (N_18797,N_18674,N_18620);
nand U18798 (N_18798,N_18566,N_18650);
or U18799 (N_18799,N_18638,N_18606);
nand U18800 (N_18800,N_18626,N_18704);
nand U18801 (N_18801,N_18716,N_18625);
nor U18802 (N_18802,N_18663,N_18609);
and U18803 (N_18803,N_18621,N_18671);
and U18804 (N_18804,N_18679,N_18633);
nand U18805 (N_18805,N_18580,N_18700);
nand U18806 (N_18806,N_18570,N_18678);
nand U18807 (N_18807,N_18574,N_18700);
xnor U18808 (N_18808,N_18670,N_18707);
nand U18809 (N_18809,N_18589,N_18612);
xor U18810 (N_18810,N_18578,N_18634);
nand U18811 (N_18811,N_18616,N_18643);
xnor U18812 (N_18812,N_18623,N_18659);
nor U18813 (N_18813,N_18637,N_18646);
nor U18814 (N_18814,N_18589,N_18674);
nand U18815 (N_18815,N_18702,N_18704);
nor U18816 (N_18816,N_18686,N_18709);
nand U18817 (N_18817,N_18563,N_18674);
xor U18818 (N_18818,N_18563,N_18644);
and U18819 (N_18819,N_18700,N_18684);
nor U18820 (N_18820,N_18598,N_18597);
nor U18821 (N_18821,N_18587,N_18708);
xnor U18822 (N_18822,N_18674,N_18693);
nand U18823 (N_18823,N_18571,N_18658);
and U18824 (N_18824,N_18629,N_18639);
and U18825 (N_18825,N_18564,N_18619);
nand U18826 (N_18826,N_18652,N_18676);
and U18827 (N_18827,N_18695,N_18651);
xnor U18828 (N_18828,N_18683,N_18658);
nand U18829 (N_18829,N_18687,N_18692);
and U18830 (N_18830,N_18568,N_18655);
or U18831 (N_18831,N_18596,N_18648);
and U18832 (N_18832,N_18631,N_18692);
nor U18833 (N_18833,N_18576,N_18633);
nor U18834 (N_18834,N_18617,N_18690);
or U18835 (N_18835,N_18571,N_18650);
and U18836 (N_18836,N_18715,N_18661);
nor U18837 (N_18837,N_18687,N_18670);
nand U18838 (N_18838,N_18710,N_18568);
xor U18839 (N_18839,N_18706,N_18615);
nor U18840 (N_18840,N_18575,N_18631);
nand U18841 (N_18841,N_18663,N_18647);
nor U18842 (N_18842,N_18584,N_18654);
or U18843 (N_18843,N_18704,N_18593);
xnor U18844 (N_18844,N_18629,N_18614);
and U18845 (N_18845,N_18589,N_18682);
or U18846 (N_18846,N_18626,N_18633);
and U18847 (N_18847,N_18671,N_18628);
and U18848 (N_18848,N_18696,N_18680);
nor U18849 (N_18849,N_18639,N_18690);
nand U18850 (N_18850,N_18671,N_18680);
or U18851 (N_18851,N_18620,N_18614);
and U18852 (N_18852,N_18671,N_18636);
nand U18853 (N_18853,N_18661,N_18595);
nor U18854 (N_18854,N_18641,N_18600);
nor U18855 (N_18855,N_18574,N_18610);
or U18856 (N_18856,N_18590,N_18622);
nor U18857 (N_18857,N_18615,N_18686);
nor U18858 (N_18858,N_18604,N_18573);
nand U18859 (N_18859,N_18575,N_18663);
or U18860 (N_18860,N_18630,N_18625);
nor U18861 (N_18861,N_18660,N_18582);
nor U18862 (N_18862,N_18598,N_18632);
and U18863 (N_18863,N_18671,N_18617);
nor U18864 (N_18864,N_18591,N_18637);
or U18865 (N_18865,N_18618,N_18651);
or U18866 (N_18866,N_18582,N_18611);
or U18867 (N_18867,N_18658,N_18622);
nor U18868 (N_18868,N_18596,N_18641);
nand U18869 (N_18869,N_18656,N_18665);
xor U18870 (N_18870,N_18666,N_18677);
nor U18871 (N_18871,N_18610,N_18579);
or U18872 (N_18872,N_18650,N_18608);
xor U18873 (N_18873,N_18683,N_18607);
xor U18874 (N_18874,N_18706,N_18628);
nor U18875 (N_18875,N_18696,N_18692);
xor U18876 (N_18876,N_18691,N_18693);
nand U18877 (N_18877,N_18717,N_18618);
nor U18878 (N_18878,N_18642,N_18644);
nor U18879 (N_18879,N_18662,N_18633);
xnor U18880 (N_18880,N_18822,N_18769);
nor U18881 (N_18881,N_18837,N_18772);
nor U18882 (N_18882,N_18754,N_18730);
nand U18883 (N_18883,N_18818,N_18801);
nand U18884 (N_18884,N_18722,N_18815);
xor U18885 (N_18885,N_18835,N_18824);
xor U18886 (N_18886,N_18846,N_18843);
nand U18887 (N_18887,N_18839,N_18743);
nand U18888 (N_18888,N_18762,N_18753);
nor U18889 (N_18889,N_18850,N_18793);
nor U18890 (N_18890,N_18774,N_18776);
nand U18891 (N_18891,N_18795,N_18814);
and U18892 (N_18892,N_18777,N_18831);
or U18893 (N_18893,N_18851,N_18834);
or U18894 (N_18894,N_18724,N_18859);
or U18895 (N_18895,N_18782,N_18790);
nand U18896 (N_18896,N_18844,N_18853);
xor U18897 (N_18897,N_18808,N_18875);
and U18898 (N_18898,N_18852,N_18784);
and U18899 (N_18899,N_18735,N_18797);
xor U18900 (N_18900,N_18826,N_18825);
xor U18901 (N_18901,N_18840,N_18868);
xnor U18902 (N_18902,N_18761,N_18766);
and U18903 (N_18903,N_18849,N_18873);
or U18904 (N_18904,N_18729,N_18727);
nand U18905 (N_18905,N_18847,N_18745);
or U18906 (N_18906,N_18781,N_18785);
and U18907 (N_18907,N_18802,N_18759);
or U18908 (N_18908,N_18836,N_18721);
or U18909 (N_18909,N_18866,N_18828);
xnor U18910 (N_18910,N_18751,N_18794);
or U18911 (N_18911,N_18755,N_18812);
or U18912 (N_18912,N_18804,N_18783);
or U18913 (N_18913,N_18750,N_18775);
and U18914 (N_18914,N_18756,N_18857);
nand U18915 (N_18915,N_18813,N_18865);
nand U18916 (N_18916,N_18823,N_18732);
xor U18917 (N_18917,N_18788,N_18821);
nand U18918 (N_18918,N_18767,N_18771);
or U18919 (N_18919,N_18879,N_18746);
or U18920 (N_18920,N_18838,N_18747);
xor U18921 (N_18921,N_18741,N_18787);
or U18922 (N_18922,N_18737,N_18768);
or U18923 (N_18923,N_18734,N_18749);
or U18924 (N_18924,N_18806,N_18858);
nor U18925 (N_18925,N_18848,N_18792);
nand U18926 (N_18926,N_18817,N_18803);
nor U18927 (N_18927,N_18752,N_18763);
xor U18928 (N_18928,N_18760,N_18829);
nand U18929 (N_18929,N_18874,N_18878);
nor U18930 (N_18930,N_18786,N_18740);
nor U18931 (N_18931,N_18871,N_18739);
and U18932 (N_18932,N_18861,N_18830);
or U18933 (N_18933,N_18733,N_18799);
xor U18934 (N_18934,N_18800,N_18728);
or U18935 (N_18935,N_18807,N_18872);
or U18936 (N_18936,N_18791,N_18778);
nor U18937 (N_18937,N_18736,N_18876);
or U18938 (N_18938,N_18842,N_18796);
nor U18939 (N_18939,N_18725,N_18757);
xnor U18940 (N_18940,N_18869,N_18870);
xor U18941 (N_18941,N_18811,N_18773);
or U18942 (N_18942,N_18833,N_18805);
or U18943 (N_18943,N_18832,N_18862);
nand U18944 (N_18944,N_18723,N_18731);
or U18945 (N_18945,N_18867,N_18758);
nor U18946 (N_18946,N_18810,N_18780);
and U18947 (N_18947,N_18748,N_18779);
and U18948 (N_18948,N_18854,N_18820);
nor U18949 (N_18949,N_18738,N_18856);
xnor U18950 (N_18950,N_18855,N_18841);
and U18951 (N_18951,N_18864,N_18860);
or U18952 (N_18952,N_18764,N_18726);
xor U18953 (N_18953,N_18827,N_18770);
and U18954 (N_18954,N_18798,N_18819);
and U18955 (N_18955,N_18789,N_18877);
and U18956 (N_18956,N_18816,N_18845);
xnor U18957 (N_18957,N_18744,N_18765);
xor U18958 (N_18958,N_18809,N_18742);
and U18959 (N_18959,N_18863,N_18720);
nand U18960 (N_18960,N_18833,N_18821);
xor U18961 (N_18961,N_18842,N_18788);
or U18962 (N_18962,N_18757,N_18862);
nor U18963 (N_18963,N_18848,N_18861);
or U18964 (N_18964,N_18756,N_18783);
nor U18965 (N_18965,N_18720,N_18873);
and U18966 (N_18966,N_18865,N_18822);
and U18967 (N_18967,N_18754,N_18876);
nor U18968 (N_18968,N_18829,N_18849);
or U18969 (N_18969,N_18847,N_18856);
xnor U18970 (N_18970,N_18788,N_18781);
or U18971 (N_18971,N_18786,N_18844);
and U18972 (N_18972,N_18824,N_18878);
nor U18973 (N_18973,N_18861,N_18844);
or U18974 (N_18974,N_18851,N_18862);
or U18975 (N_18975,N_18730,N_18751);
nand U18976 (N_18976,N_18772,N_18728);
or U18977 (N_18977,N_18814,N_18855);
nor U18978 (N_18978,N_18879,N_18778);
and U18979 (N_18979,N_18757,N_18794);
or U18980 (N_18980,N_18737,N_18866);
nand U18981 (N_18981,N_18724,N_18771);
xor U18982 (N_18982,N_18748,N_18814);
xnor U18983 (N_18983,N_18728,N_18852);
xnor U18984 (N_18984,N_18825,N_18862);
xnor U18985 (N_18985,N_18746,N_18874);
nand U18986 (N_18986,N_18819,N_18797);
and U18987 (N_18987,N_18865,N_18733);
and U18988 (N_18988,N_18835,N_18721);
or U18989 (N_18989,N_18724,N_18845);
and U18990 (N_18990,N_18767,N_18822);
and U18991 (N_18991,N_18841,N_18774);
and U18992 (N_18992,N_18802,N_18768);
nor U18993 (N_18993,N_18752,N_18815);
xor U18994 (N_18994,N_18810,N_18792);
xnor U18995 (N_18995,N_18804,N_18812);
nand U18996 (N_18996,N_18826,N_18869);
xor U18997 (N_18997,N_18753,N_18739);
or U18998 (N_18998,N_18833,N_18773);
nand U18999 (N_18999,N_18748,N_18781);
nand U19000 (N_19000,N_18751,N_18783);
and U19001 (N_19001,N_18850,N_18747);
xor U19002 (N_19002,N_18778,N_18818);
and U19003 (N_19003,N_18878,N_18772);
nor U19004 (N_19004,N_18748,N_18791);
nor U19005 (N_19005,N_18767,N_18783);
xor U19006 (N_19006,N_18761,N_18852);
or U19007 (N_19007,N_18777,N_18771);
xnor U19008 (N_19008,N_18770,N_18855);
nand U19009 (N_19009,N_18828,N_18781);
or U19010 (N_19010,N_18828,N_18746);
xnor U19011 (N_19011,N_18762,N_18812);
nor U19012 (N_19012,N_18751,N_18737);
and U19013 (N_19013,N_18770,N_18737);
or U19014 (N_19014,N_18766,N_18726);
nor U19015 (N_19015,N_18816,N_18796);
xor U19016 (N_19016,N_18820,N_18817);
or U19017 (N_19017,N_18856,N_18860);
nand U19018 (N_19018,N_18860,N_18806);
nand U19019 (N_19019,N_18834,N_18846);
xor U19020 (N_19020,N_18770,N_18835);
and U19021 (N_19021,N_18795,N_18853);
nand U19022 (N_19022,N_18759,N_18862);
xor U19023 (N_19023,N_18817,N_18868);
and U19024 (N_19024,N_18724,N_18757);
nor U19025 (N_19025,N_18825,N_18747);
and U19026 (N_19026,N_18783,N_18849);
xor U19027 (N_19027,N_18733,N_18782);
xor U19028 (N_19028,N_18801,N_18823);
nor U19029 (N_19029,N_18817,N_18774);
nor U19030 (N_19030,N_18758,N_18877);
or U19031 (N_19031,N_18868,N_18786);
nand U19032 (N_19032,N_18749,N_18808);
nand U19033 (N_19033,N_18828,N_18845);
nor U19034 (N_19034,N_18852,N_18822);
xor U19035 (N_19035,N_18752,N_18759);
nand U19036 (N_19036,N_18878,N_18819);
and U19037 (N_19037,N_18829,N_18812);
or U19038 (N_19038,N_18787,N_18790);
xor U19039 (N_19039,N_18741,N_18771);
xor U19040 (N_19040,N_18890,N_18917);
or U19041 (N_19041,N_19015,N_18921);
xor U19042 (N_19042,N_18898,N_18900);
xnor U19043 (N_19043,N_18974,N_18887);
or U19044 (N_19044,N_18936,N_18983);
and U19045 (N_19045,N_18994,N_18992);
nor U19046 (N_19046,N_18981,N_18989);
and U19047 (N_19047,N_18958,N_18970);
xor U19048 (N_19048,N_18987,N_19014);
xor U19049 (N_19049,N_18937,N_18904);
and U19050 (N_19050,N_19019,N_18961);
or U19051 (N_19051,N_19005,N_18930);
nand U19052 (N_19052,N_18991,N_18903);
or U19053 (N_19053,N_19011,N_18929);
xnor U19054 (N_19054,N_18977,N_18988);
xor U19055 (N_19055,N_18942,N_19028);
nor U19056 (N_19056,N_18998,N_19029);
and U19057 (N_19057,N_18955,N_19038);
nand U19058 (N_19058,N_18911,N_18882);
nor U19059 (N_19059,N_19001,N_19004);
and U19060 (N_19060,N_18984,N_18923);
nor U19061 (N_19061,N_18949,N_19023);
or U19062 (N_19062,N_18894,N_19039);
and U19063 (N_19063,N_18956,N_18966);
and U19064 (N_19064,N_19013,N_18924);
nor U19065 (N_19065,N_18971,N_18914);
or U19066 (N_19066,N_18928,N_18922);
and U19067 (N_19067,N_19017,N_19016);
nand U19068 (N_19068,N_18881,N_19018);
xor U19069 (N_19069,N_18886,N_18931);
nor U19070 (N_19070,N_19007,N_18938);
and U19071 (N_19071,N_19032,N_18905);
nor U19072 (N_19072,N_19022,N_18941);
xor U19073 (N_19073,N_18950,N_19037);
or U19074 (N_19074,N_18979,N_18968);
nor U19075 (N_19075,N_18909,N_19035);
nand U19076 (N_19076,N_18932,N_18885);
or U19077 (N_19077,N_18940,N_18964);
nor U19078 (N_19078,N_18888,N_18954);
xor U19079 (N_19079,N_18915,N_18920);
or U19080 (N_19080,N_18916,N_18933);
or U19081 (N_19081,N_18960,N_18897);
nand U19082 (N_19082,N_18980,N_18906);
nor U19083 (N_19083,N_18884,N_18926);
or U19084 (N_19084,N_18990,N_18925);
xor U19085 (N_19085,N_18918,N_18953);
xor U19086 (N_19086,N_18996,N_19025);
xor U19087 (N_19087,N_18943,N_18899);
and U19088 (N_19088,N_18893,N_18913);
xnor U19089 (N_19089,N_18957,N_19020);
or U19090 (N_19090,N_18976,N_18993);
and U19091 (N_19091,N_19003,N_19034);
and U19092 (N_19092,N_18967,N_18962);
and U19093 (N_19093,N_18978,N_19009);
nor U19094 (N_19094,N_18997,N_18946);
xor U19095 (N_19095,N_19021,N_19024);
nand U19096 (N_19096,N_18889,N_18908);
or U19097 (N_19097,N_18901,N_19012);
and U19098 (N_19098,N_18969,N_18944);
nand U19099 (N_19099,N_18999,N_18895);
xor U19100 (N_19100,N_18985,N_19030);
or U19101 (N_19101,N_19006,N_18907);
xor U19102 (N_19102,N_18965,N_19010);
xor U19103 (N_19103,N_18963,N_18912);
xnor U19104 (N_19104,N_19000,N_18995);
nor U19105 (N_19105,N_18959,N_18927);
nor U19106 (N_19106,N_18951,N_18919);
xor U19107 (N_19107,N_18934,N_18892);
nand U19108 (N_19108,N_18973,N_18947);
or U19109 (N_19109,N_18891,N_18896);
or U19110 (N_19110,N_18883,N_18948);
nand U19111 (N_19111,N_19031,N_18939);
nor U19112 (N_19112,N_18880,N_18952);
nand U19113 (N_19113,N_19008,N_19033);
and U19114 (N_19114,N_18975,N_19036);
nand U19115 (N_19115,N_18972,N_18986);
or U19116 (N_19116,N_19026,N_18982);
xnor U19117 (N_19117,N_18902,N_18945);
nand U19118 (N_19118,N_19002,N_18910);
nand U19119 (N_19119,N_18935,N_19027);
and U19120 (N_19120,N_18990,N_19019);
nand U19121 (N_19121,N_18959,N_19029);
or U19122 (N_19122,N_18996,N_18950);
or U19123 (N_19123,N_18994,N_18971);
nor U19124 (N_19124,N_19035,N_18903);
and U19125 (N_19125,N_18975,N_18989);
nand U19126 (N_19126,N_19007,N_18996);
nor U19127 (N_19127,N_18900,N_18932);
xnor U19128 (N_19128,N_18971,N_18935);
nand U19129 (N_19129,N_18976,N_18943);
nor U19130 (N_19130,N_18995,N_18956);
or U19131 (N_19131,N_18884,N_18993);
nor U19132 (N_19132,N_18961,N_18968);
or U19133 (N_19133,N_18945,N_18960);
or U19134 (N_19134,N_18967,N_19002);
and U19135 (N_19135,N_18907,N_18880);
or U19136 (N_19136,N_18894,N_18950);
nand U19137 (N_19137,N_19035,N_18955);
nand U19138 (N_19138,N_18987,N_19028);
nor U19139 (N_19139,N_19035,N_18927);
nand U19140 (N_19140,N_18919,N_18880);
nand U19141 (N_19141,N_18907,N_18902);
or U19142 (N_19142,N_19017,N_18960);
xnor U19143 (N_19143,N_18971,N_18903);
or U19144 (N_19144,N_18927,N_18989);
or U19145 (N_19145,N_18947,N_18910);
and U19146 (N_19146,N_18958,N_19009);
xnor U19147 (N_19147,N_19028,N_18887);
nand U19148 (N_19148,N_18984,N_18893);
and U19149 (N_19149,N_18965,N_18893);
or U19150 (N_19150,N_19030,N_19006);
xnor U19151 (N_19151,N_18913,N_18934);
xor U19152 (N_19152,N_18895,N_18918);
and U19153 (N_19153,N_18895,N_19026);
or U19154 (N_19154,N_18992,N_18984);
or U19155 (N_19155,N_18960,N_18991);
xnor U19156 (N_19156,N_18965,N_18966);
xnor U19157 (N_19157,N_18994,N_18921);
xnor U19158 (N_19158,N_18914,N_18894);
nand U19159 (N_19159,N_19036,N_18924);
nand U19160 (N_19160,N_18896,N_18927);
xnor U19161 (N_19161,N_18924,N_18935);
and U19162 (N_19162,N_19004,N_18958);
and U19163 (N_19163,N_18912,N_19031);
or U19164 (N_19164,N_19000,N_18886);
xor U19165 (N_19165,N_18921,N_19006);
and U19166 (N_19166,N_19002,N_19018);
and U19167 (N_19167,N_18894,N_18964);
nand U19168 (N_19168,N_19027,N_18928);
xnor U19169 (N_19169,N_19032,N_18943);
nor U19170 (N_19170,N_19006,N_18905);
or U19171 (N_19171,N_19004,N_19024);
nand U19172 (N_19172,N_18950,N_18897);
or U19173 (N_19173,N_18951,N_19008);
nand U19174 (N_19174,N_19021,N_18925);
nand U19175 (N_19175,N_18914,N_18905);
nor U19176 (N_19176,N_18971,N_18988);
or U19177 (N_19177,N_18901,N_19001);
and U19178 (N_19178,N_18914,N_18955);
and U19179 (N_19179,N_19038,N_18949);
xnor U19180 (N_19180,N_18953,N_18905);
nor U19181 (N_19181,N_18974,N_18965);
xor U19182 (N_19182,N_18987,N_18999);
xnor U19183 (N_19183,N_18908,N_18918);
or U19184 (N_19184,N_18963,N_18966);
and U19185 (N_19185,N_19011,N_18882);
xor U19186 (N_19186,N_19031,N_18913);
nand U19187 (N_19187,N_18921,N_18908);
xnor U19188 (N_19188,N_18902,N_18895);
or U19189 (N_19189,N_18935,N_18989);
and U19190 (N_19190,N_18984,N_18927);
nand U19191 (N_19191,N_19032,N_18906);
nor U19192 (N_19192,N_19019,N_18978);
xnor U19193 (N_19193,N_19028,N_18965);
nor U19194 (N_19194,N_18966,N_19033);
and U19195 (N_19195,N_18991,N_18985);
nor U19196 (N_19196,N_18932,N_18921);
nor U19197 (N_19197,N_18906,N_18944);
or U19198 (N_19198,N_18894,N_18997);
and U19199 (N_19199,N_18957,N_18884);
nand U19200 (N_19200,N_19045,N_19160);
nand U19201 (N_19201,N_19170,N_19081);
nor U19202 (N_19202,N_19115,N_19069);
nand U19203 (N_19203,N_19190,N_19098);
or U19204 (N_19204,N_19168,N_19118);
nand U19205 (N_19205,N_19151,N_19086);
and U19206 (N_19206,N_19048,N_19172);
nand U19207 (N_19207,N_19145,N_19054);
nand U19208 (N_19208,N_19181,N_19062);
and U19209 (N_19209,N_19096,N_19191);
or U19210 (N_19210,N_19042,N_19084);
or U19211 (N_19211,N_19197,N_19165);
xnor U19212 (N_19212,N_19169,N_19199);
nand U19213 (N_19213,N_19156,N_19043);
and U19214 (N_19214,N_19051,N_19056);
or U19215 (N_19215,N_19067,N_19150);
xor U19216 (N_19216,N_19125,N_19159);
and U19217 (N_19217,N_19180,N_19095);
or U19218 (N_19218,N_19102,N_19093);
or U19219 (N_19219,N_19107,N_19133);
xnor U19220 (N_19220,N_19140,N_19104);
nand U19221 (N_19221,N_19182,N_19076);
and U19222 (N_19222,N_19153,N_19198);
xor U19223 (N_19223,N_19193,N_19132);
or U19224 (N_19224,N_19103,N_19113);
or U19225 (N_19225,N_19094,N_19055);
nor U19226 (N_19226,N_19164,N_19126);
and U19227 (N_19227,N_19099,N_19143);
or U19228 (N_19228,N_19087,N_19174);
nand U19229 (N_19229,N_19058,N_19152);
and U19230 (N_19230,N_19137,N_19173);
and U19231 (N_19231,N_19163,N_19158);
nor U19232 (N_19232,N_19171,N_19135);
xnor U19233 (N_19233,N_19085,N_19123);
nand U19234 (N_19234,N_19092,N_19109);
and U19235 (N_19235,N_19189,N_19046);
nor U19236 (N_19236,N_19120,N_19097);
xor U19237 (N_19237,N_19090,N_19077);
xnor U19238 (N_19238,N_19078,N_19074);
and U19239 (N_19239,N_19179,N_19186);
nand U19240 (N_19240,N_19116,N_19129);
xor U19241 (N_19241,N_19079,N_19065);
and U19242 (N_19242,N_19155,N_19060);
nand U19243 (N_19243,N_19148,N_19177);
and U19244 (N_19244,N_19161,N_19080);
xnor U19245 (N_19245,N_19138,N_19157);
nor U19246 (N_19246,N_19112,N_19053);
and U19247 (N_19247,N_19057,N_19128);
or U19248 (N_19248,N_19059,N_19185);
nor U19249 (N_19249,N_19187,N_19070);
and U19250 (N_19250,N_19121,N_19044);
xor U19251 (N_19251,N_19127,N_19088);
nor U19252 (N_19252,N_19183,N_19188);
nand U19253 (N_19253,N_19111,N_19131);
or U19254 (N_19254,N_19147,N_19040);
and U19255 (N_19255,N_19146,N_19068);
nand U19256 (N_19256,N_19089,N_19117);
or U19257 (N_19257,N_19082,N_19091);
xnor U19258 (N_19258,N_19162,N_19144);
or U19259 (N_19259,N_19052,N_19105);
and U19260 (N_19260,N_19141,N_19108);
nor U19261 (N_19261,N_19119,N_19195);
or U19262 (N_19262,N_19075,N_19130);
xnor U19263 (N_19263,N_19184,N_19178);
xor U19264 (N_19264,N_19100,N_19110);
nand U19265 (N_19265,N_19101,N_19106);
xnor U19266 (N_19266,N_19167,N_19154);
or U19267 (N_19267,N_19192,N_19136);
nor U19268 (N_19268,N_19071,N_19061);
nand U19269 (N_19269,N_19134,N_19196);
nor U19270 (N_19270,N_19142,N_19047);
xor U19271 (N_19271,N_19122,N_19194);
nor U19272 (N_19272,N_19176,N_19114);
or U19273 (N_19273,N_19064,N_19066);
nand U19274 (N_19274,N_19139,N_19049);
nor U19275 (N_19275,N_19050,N_19149);
and U19276 (N_19276,N_19073,N_19041);
or U19277 (N_19277,N_19072,N_19083);
nand U19278 (N_19278,N_19063,N_19175);
and U19279 (N_19279,N_19124,N_19166);
and U19280 (N_19280,N_19078,N_19082);
or U19281 (N_19281,N_19109,N_19182);
nand U19282 (N_19282,N_19072,N_19196);
nor U19283 (N_19283,N_19053,N_19097);
or U19284 (N_19284,N_19041,N_19064);
or U19285 (N_19285,N_19159,N_19066);
and U19286 (N_19286,N_19135,N_19113);
xnor U19287 (N_19287,N_19048,N_19072);
nand U19288 (N_19288,N_19120,N_19192);
nor U19289 (N_19289,N_19096,N_19060);
xor U19290 (N_19290,N_19067,N_19186);
nor U19291 (N_19291,N_19144,N_19108);
or U19292 (N_19292,N_19083,N_19070);
xor U19293 (N_19293,N_19127,N_19064);
nor U19294 (N_19294,N_19154,N_19061);
and U19295 (N_19295,N_19186,N_19121);
and U19296 (N_19296,N_19102,N_19191);
nand U19297 (N_19297,N_19138,N_19190);
nor U19298 (N_19298,N_19194,N_19134);
or U19299 (N_19299,N_19163,N_19137);
or U19300 (N_19300,N_19186,N_19087);
or U19301 (N_19301,N_19197,N_19055);
xnor U19302 (N_19302,N_19198,N_19184);
or U19303 (N_19303,N_19059,N_19116);
or U19304 (N_19304,N_19115,N_19134);
and U19305 (N_19305,N_19104,N_19128);
or U19306 (N_19306,N_19189,N_19044);
or U19307 (N_19307,N_19172,N_19083);
xor U19308 (N_19308,N_19077,N_19154);
nor U19309 (N_19309,N_19185,N_19101);
and U19310 (N_19310,N_19152,N_19102);
and U19311 (N_19311,N_19046,N_19183);
nand U19312 (N_19312,N_19056,N_19145);
nand U19313 (N_19313,N_19192,N_19102);
nor U19314 (N_19314,N_19126,N_19069);
xnor U19315 (N_19315,N_19152,N_19143);
and U19316 (N_19316,N_19188,N_19131);
and U19317 (N_19317,N_19077,N_19091);
xnor U19318 (N_19318,N_19175,N_19195);
or U19319 (N_19319,N_19151,N_19192);
nand U19320 (N_19320,N_19154,N_19081);
nor U19321 (N_19321,N_19116,N_19118);
nor U19322 (N_19322,N_19097,N_19046);
nand U19323 (N_19323,N_19053,N_19099);
xnor U19324 (N_19324,N_19086,N_19152);
xor U19325 (N_19325,N_19159,N_19195);
nor U19326 (N_19326,N_19152,N_19147);
nand U19327 (N_19327,N_19181,N_19096);
nor U19328 (N_19328,N_19165,N_19068);
nor U19329 (N_19329,N_19132,N_19080);
and U19330 (N_19330,N_19068,N_19162);
and U19331 (N_19331,N_19081,N_19049);
nand U19332 (N_19332,N_19057,N_19077);
nor U19333 (N_19333,N_19168,N_19185);
or U19334 (N_19334,N_19066,N_19092);
or U19335 (N_19335,N_19170,N_19171);
nor U19336 (N_19336,N_19169,N_19181);
nand U19337 (N_19337,N_19151,N_19113);
and U19338 (N_19338,N_19135,N_19087);
and U19339 (N_19339,N_19135,N_19121);
xnor U19340 (N_19340,N_19127,N_19190);
or U19341 (N_19341,N_19142,N_19191);
nor U19342 (N_19342,N_19144,N_19069);
and U19343 (N_19343,N_19127,N_19101);
xor U19344 (N_19344,N_19064,N_19117);
nand U19345 (N_19345,N_19073,N_19198);
xor U19346 (N_19346,N_19082,N_19164);
nand U19347 (N_19347,N_19161,N_19118);
xor U19348 (N_19348,N_19114,N_19174);
xnor U19349 (N_19349,N_19083,N_19064);
nand U19350 (N_19350,N_19090,N_19155);
xor U19351 (N_19351,N_19049,N_19197);
or U19352 (N_19352,N_19085,N_19115);
and U19353 (N_19353,N_19140,N_19147);
and U19354 (N_19354,N_19066,N_19190);
nor U19355 (N_19355,N_19166,N_19044);
xor U19356 (N_19356,N_19115,N_19130);
nand U19357 (N_19357,N_19073,N_19114);
xnor U19358 (N_19358,N_19124,N_19059);
and U19359 (N_19359,N_19141,N_19056);
or U19360 (N_19360,N_19306,N_19232);
or U19361 (N_19361,N_19256,N_19337);
and U19362 (N_19362,N_19210,N_19237);
nor U19363 (N_19363,N_19273,N_19223);
xnor U19364 (N_19364,N_19291,N_19341);
nor U19365 (N_19365,N_19285,N_19312);
and U19366 (N_19366,N_19319,N_19204);
nor U19367 (N_19367,N_19202,N_19243);
nor U19368 (N_19368,N_19288,N_19229);
xnor U19369 (N_19369,N_19203,N_19205);
nor U19370 (N_19370,N_19263,N_19310);
xnor U19371 (N_19371,N_19258,N_19259);
nor U19372 (N_19372,N_19290,N_19340);
nand U19373 (N_19373,N_19280,N_19287);
nor U19374 (N_19374,N_19222,N_19283);
nand U19375 (N_19375,N_19294,N_19220);
xnor U19376 (N_19376,N_19267,N_19209);
or U19377 (N_19377,N_19356,N_19239);
or U19378 (N_19378,N_19292,N_19269);
and U19379 (N_19379,N_19355,N_19246);
nor U19380 (N_19380,N_19307,N_19255);
nand U19381 (N_19381,N_19298,N_19231);
nor U19382 (N_19382,N_19211,N_19226);
or U19383 (N_19383,N_19215,N_19260);
and U19384 (N_19384,N_19349,N_19245);
nand U19385 (N_19385,N_19224,N_19329);
or U19386 (N_19386,N_19354,N_19304);
or U19387 (N_19387,N_19324,N_19225);
and U19388 (N_19388,N_19328,N_19279);
nor U19389 (N_19389,N_19317,N_19271);
or U19390 (N_19390,N_19212,N_19200);
xor U19391 (N_19391,N_19253,N_19270);
nand U19392 (N_19392,N_19353,N_19216);
or U19393 (N_19393,N_19327,N_19321);
nand U19394 (N_19394,N_19228,N_19330);
xor U19395 (N_19395,N_19272,N_19289);
nand U19396 (N_19396,N_19357,N_19325);
xnor U19397 (N_19397,N_19251,N_19303);
nand U19398 (N_19398,N_19282,N_19208);
nor U19399 (N_19399,N_19248,N_19331);
xnor U19400 (N_19400,N_19350,N_19238);
nor U19401 (N_19401,N_19301,N_19320);
nor U19402 (N_19402,N_19266,N_19352);
nor U19403 (N_19403,N_19316,N_19326);
nand U19404 (N_19404,N_19300,N_19305);
and U19405 (N_19405,N_19274,N_19242);
xor U19406 (N_19406,N_19250,N_19261);
or U19407 (N_19407,N_19213,N_19240);
and U19408 (N_19408,N_19234,N_19315);
nor U19409 (N_19409,N_19351,N_19227);
nand U19410 (N_19410,N_19342,N_19257);
xnor U19411 (N_19411,N_19302,N_19334);
xor U19412 (N_19412,N_19233,N_19268);
nor U19413 (N_19413,N_19346,N_19275);
nor U19414 (N_19414,N_19244,N_19265);
and U19415 (N_19415,N_19347,N_19235);
and U19416 (N_19416,N_19241,N_19201);
or U19417 (N_19417,N_19309,N_19335);
xor U19418 (N_19418,N_19308,N_19214);
nor U19419 (N_19419,N_19348,N_19219);
xnor U19420 (N_19420,N_19344,N_19249);
xnor U19421 (N_19421,N_19336,N_19339);
or U19422 (N_19422,N_19318,N_19230);
nor U19423 (N_19423,N_19359,N_19276);
xnor U19424 (N_19424,N_19333,N_19296);
nand U19425 (N_19425,N_19277,N_19252);
and U19426 (N_19426,N_19278,N_19358);
or U19427 (N_19427,N_19284,N_19313);
nor U19428 (N_19428,N_19247,N_19207);
nand U19429 (N_19429,N_19286,N_19323);
xnor U19430 (N_19430,N_19322,N_19338);
or U19431 (N_19431,N_19343,N_19254);
xor U19432 (N_19432,N_19221,N_19299);
and U19433 (N_19433,N_19314,N_19217);
xor U19434 (N_19434,N_19264,N_19281);
nand U19435 (N_19435,N_19295,N_19297);
and U19436 (N_19436,N_19218,N_19236);
nand U19437 (N_19437,N_19332,N_19345);
nand U19438 (N_19438,N_19262,N_19293);
or U19439 (N_19439,N_19311,N_19206);
xnor U19440 (N_19440,N_19348,N_19323);
and U19441 (N_19441,N_19356,N_19301);
xor U19442 (N_19442,N_19279,N_19254);
nor U19443 (N_19443,N_19208,N_19221);
xor U19444 (N_19444,N_19280,N_19293);
and U19445 (N_19445,N_19295,N_19310);
nand U19446 (N_19446,N_19228,N_19247);
nand U19447 (N_19447,N_19293,N_19359);
or U19448 (N_19448,N_19350,N_19266);
xor U19449 (N_19449,N_19201,N_19344);
xnor U19450 (N_19450,N_19233,N_19351);
xor U19451 (N_19451,N_19265,N_19268);
nand U19452 (N_19452,N_19317,N_19214);
xnor U19453 (N_19453,N_19322,N_19241);
nand U19454 (N_19454,N_19305,N_19236);
nand U19455 (N_19455,N_19207,N_19333);
nand U19456 (N_19456,N_19346,N_19228);
nand U19457 (N_19457,N_19206,N_19232);
xor U19458 (N_19458,N_19274,N_19275);
or U19459 (N_19459,N_19309,N_19259);
xor U19460 (N_19460,N_19324,N_19208);
nor U19461 (N_19461,N_19241,N_19211);
nand U19462 (N_19462,N_19326,N_19299);
and U19463 (N_19463,N_19273,N_19326);
and U19464 (N_19464,N_19263,N_19207);
nand U19465 (N_19465,N_19216,N_19257);
and U19466 (N_19466,N_19294,N_19270);
nand U19467 (N_19467,N_19322,N_19201);
and U19468 (N_19468,N_19328,N_19213);
nand U19469 (N_19469,N_19207,N_19348);
xnor U19470 (N_19470,N_19356,N_19229);
and U19471 (N_19471,N_19226,N_19286);
and U19472 (N_19472,N_19235,N_19348);
or U19473 (N_19473,N_19251,N_19280);
xnor U19474 (N_19474,N_19338,N_19340);
nor U19475 (N_19475,N_19206,N_19321);
or U19476 (N_19476,N_19312,N_19226);
nand U19477 (N_19477,N_19258,N_19231);
and U19478 (N_19478,N_19284,N_19291);
nor U19479 (N_19479,N_19305,N_19313);
and U19480 (N_19480,N_19299,N_19267);
xnor U19481 (N_19481,N_19335,N_19212);
nor U19482 (N_19482,N_19313,N_19258);
nor U19483 (N_19483,N_19253,N_19267);
nand U19484 (N_19484,N_19244,N_19269);
and U19485 (N_19485,N_19316,N_19292);
or U19486 (N_19486,N_19222,N_19227);
xnor U19487 (N_19487,N_19245,N_19313);
and U19488 (N_19488,N_19285,N_19304);
xnor U19489 (N_19489,N_19330,N_19224);
or U19490 (N_19490,N_19292,N_19301);
and U19491 (N_19491,N_19297,N_19280);
nand U19492 (N_19492,N_19216,N_19266);
nor U19493 (N_19493,N_19339,N_19312);
or U19494 (N_19494,N_19242,N_19217);
nand U19495 (N_19495,N_19231,N_19357);
and U19496 (N_19496,N_19237,N_19247);
xor U19497 (N_19497,N_19337,N_19277);
or U19498 (N_19498,N_19254,N_19313);
nand U19499 (N_19499,N_19284,N_19273);
nand U19500 (N_19500,N_19291,N_19312);
and U19501 (N_19501,N_19356,N_19216);
and U19502 (N_19502,N_19249,N_19298);
nor U19503 (N_19503,N_19289,N_19319);
or U19504 (N_19504,N_19216,N_19250);
and U19505 (N_19505,N_19350,N_19282);
or U19506 (N_19506,N_19292,N_19330);
and U19507 (N_19507,N_19320,N_19219);
xnor U19508 (N_19508,N_19354,N_19301);
and U19509 (N_19509,N_19236,N_19315);
xnor U19510 (N_19510,N_19204,N_19302);
xor U19511 (N_19511,N_19277,N_19255);
nor U19512 (N_19512,N_19229,N_19238);
and U19513 (N_19513,N_19237,N_19226);
xnor U19514 (N_19514,N_19327,N_19302);
nand U19515 (N_19515,N_19247,N_19240);
nand U19516 (N_19516,N_19262,N_19358);
nand U19517 (N_19517,N_19214,N_19213);
and U19518 (N_19518,N_19289,N_19239);
nand U19519 (N_19519,N_19312,N_19250);
and U19520 (N_19520,N_19418,N_19429);
xor U19521 (N_19521,N_19403,N_19407);
xnor U19522 (N_19522,N_19462,N_19496);
xor U19523 (N_19523,N_19380,N_19374);
nand U19524 (N_19524,N_19420,N_19430);
xnor U19525 (N_19525,N_19465,N_19397);
nor U19526 (N_19526,N_19364,N_19449);
nand U19527 (N_19527,N_19367,N_19393);
or U19528 (N_19528,N_19417,N_19401);
nand U19529 (N_19529,N_19428,N_19415);
and U19530 (N_19530,N_19375,N_19504);
nor U19531 (N_19531,N_19461,N_19498);
and U19532 (N_19532,N_19410,N_19435);
nor U19533 (N_19533,N_19368,N_19477);
and U19534 (N_19534,N_19492,N_19457);
and U19535 (N_19535,N_19505,N_19489);
nand U19536 (N_19536,N_19455,N_19445);
nor U19537 (N_19537,N_19454,N_19386);
or U19538 (N_19538,N_19361,N_19436);
or U19539 (N_19539,N_19499,N_19510);
nor U19540 (N_19540,N_19458,N_19399);
and U19541 (N_19541,N_19478,N_19405);
and U19542 (N_19542,N_19424,N_19441);
and U19543 (N_19543,N_19422,N_19379);
nor U19544 (N_19544,N_19451,N_19395);
or U19545 (N_19545,N_19475,N_19377);
and U19546 (N_19546,N_19448,N_19452);
nor U19547 (N_19547,N_19463,N_19385);
or U19548 (N_19548,N_19438,N_19400);
nand U19549 (N_19549,N_19450,N_19517);
or U19550 (N_19550,N_19466,N_19446);
and U19551 (N_19551,N_19431,N_19440);
and U19552 (N_19552,N_19432,N_19437);
or U19553 (N_19553,N_19490,N_19444);
or U19554 (N_19554,N_19508,N_19483);
or U19555 (N_19555,N_19502,N_19409);
nand U19556 (N_19556,N_19390,N_19456);
or U19557 (N_19557,N_19442,N_19371);
or U19558 (N_19558,N_19495,N_19468);
and U19559 (N_19559,N_19479,N_19392);
or U19560 (N_19560,N_19387,N_19481);
or U19561 (N_19561,N_19493,N_19394);
or U19562 (N_19562,N_19516,N_19427);
nor U19563 (N_19563,N_19416,N_19376);
nand U19564 (N_19564,N_19373,N_19500);
nor U19565 (N_19565,N_19443,N_19503);
nand U19566 (N_19566,N_19509,N_19414);
nor U19567 (N_19567,N_19411,N_19402);
nand U19568 (N_19568,N_19469,N_19511);
and U19569 (N_19569,N_19384,N_19363);
nand U19570 (N_19570,N_19515,N_19470);
or U19571 (N_19571,N_19472,N_19453);
nand U19572 (N_19572,N_19513,N_19425);
nor U19573 (N_19573,N_19366,N_19388);
and U19574 (N_19574,N_19412,N_19467);
xor U19575 (N_19575,N_19518,N_19473);
nor U19576 (N_19576,N_19426,N_19507);
or U19577 (N_19577,N_19460,N_19362);
and U19578 (N_19578,N_19396,N_19391);
nand U19579 (N_19579,N_19439,N_19497);
and U19580 (N_19580,N_19434,N_19484);
nand U19581 (N_19581,N_19519,N_19423);
nor U19582 (N_19582,N_19506,N_19408);
and U19583 (N_19583,N_19383,N_19413);
or U19584 (N_19584,N_19491,N_19421);
xnor U19585 (N_19585,N_19485,N_19389);
or U19586 (N_19586,N_19370,N_19433);
and U19587 (N_19587,N_19381,N_19365);
nor U19588 (N_19588,N_19372,N_19382);
nand U19589 (N_19589,N_19378,N_19464);
xnor U19590 (N_19590,N_19501,N_19447);
xor U19591 (N_19591,N_19419,N_19360);
or U19592 (N_19592,N_19476,N_19514);
nor U19593 (N_19593,N_19369,N_19480);
nand U19594 (N_19594,N_19406,N_19487);
or U19595 (N_19595,N_19486,N_19398);
nand U19596 (N_19596,N_19482,N_19488);
and U19597 (N_19597,N_19494,N_19474);
xnor U19598 (N_19598,N_19459,N_19471);
or U19599 (N_19599,N_19512,N_19404);
nand U19600 (N_19600,N_19413,N_19360);
and U19601 (N_19601,N_19425,N_19468);
nor U19602 (N_19602,N_19361,N_19404);
nor U19603 (N_19603,N_19459,N_19517);
nor U19604 (N_19604,N_19482,N_19469);
or U19605 (N_19605,N_19506,N_19439);
nor U19606 (N_19606,N_19427,N_19366);
xnor U19607 (N_19607,N_19499,N_19498);
or U19608 (N_19608,N_19444,N_19361);
nand U19609 (N_19609,N_19470,N_19476);
or U19610 (N_19610,N_19419,N_19413);
nand U19611 (N_19611,N_19370,N_19377);
and U19612 (N_19612,N_19396,N_19449);
nand U19613 (N_19613,N_19479,N_19483);
nand U19614 (N_19614,N_19511,N_19405);
nand U19615 (N_19615,N_19392,N_19453);
xnor U19616 (N_19616,N_19453,N_19405);
nor U19617 (N_19617,N_19513,N_19419);
and U19618 (N_19618,N_19440,N_19469);
or U19619 (N_19619,N_19448,N_19473);
nand U19620 (N_19620,N_19452,N_19425);
nand U19621 (N_19621,N_19499,N_19466);
nand U19622 (N_19622,N_19368,N_19519);
or U19623 (N_19623,N_19379,N_19413);
xnor U19624 (N_19624,N_19463,N_19449);
or U19625 (N_19625,N_19475,N_19411);
nand U19626 (N_19626,N_19409,N_19388);
or U19627 (N_19627,N_19376,N_19422);
or U19628 (N_19628,N_19434,N_19460);
xnor U19629 (N_19629,N_19519,N_19393);
or U19630 (N_19630,N_19503,N_19379);
or U19631 (N_19631,N_19382,N_19434);
nand U19632 (N_19632,N_19392,N_19475);
or U19633 (N_19633,N_19372,N_19390);
nand U19634 (N_19634,N_19368,N_19414);
nor U19635 (N_19635,N_19438,N_19393);
nand U19636 (N_19636,N_19396,N_19498);
or U19637 (N_19637,N_19403,N_19511);
and U19638 (N_19638,N_19511,N_19415);
or U19639 (N_19639,N_19451,N_19457);
or U19640 (N_19640,N_19440,N_19377);
nor U19641 (N_19641,N_19409,N_19481);
nor U19642 (N_19642,N_19466,N_19425);
and U19643 (N_19643,N_19368,N_19397);
nor U19644 (N_19644,N_19382,N_19414);
nor U19645 (N_19645,N_19436,N_19363);
nor U19646 (N_19646,N_19365,N_19367);
or U19647 (N_19647,N_19478,N_19372);
nand U19648 (N_19648,N_19410,N_19423);
and U19649 (N_19649,N_19436,N_19496);
xnor U19650 (N_19650,N_19375,N_19428);
or U19651 (N_19651,N_19384,N_19452);
and U19652 (N_19652,N_19417,N_19492);
nand U19653 (N_19653,N_19381,N_19427);
and U19654 (N_19654,N_19365,N_19366);
xor U19655 (N_19655,N_19384,N_19502);
nand U19656 (N_19656,N_19517,N_19504);
nand U19657 (N_19657,N_19409,N_19494);
or U19658 (N_19658,N_19456,N_19387);
nand U19659 (N_19659,N_19429,N_19376);
or U19660 (N_19660,N_19427,N_19417);
or U19661 (N_19661,N_19493,N_19449);
nand U19662 (N_19662,N_19512,N_19437);
nor U19663 (N_19663,N_19480,N_19410);
nor U19664 (N_19664,N_19508,N_19426);
nand U19665 (N_19665,N_19505,N_19372);
nand U19666 (N_19666,N_19501,N_19426);
nand U19667 (N_19667,N_19460,N_19443);
nor U19668 (N_19668,N_19428,N_19379);
nor U19669 (N_19669,N_19430,N_19394);
nor U19670 (N_19670,N_19455,N_19431);
nor U19671 (N_19671,N_19519,N_19508);
nor U19672 (N_19672,N_19423,N_19483);
and U19673 (N_19673,N_19421,N_19394);
or U19674 (N_19674,N_19495,N_19421);
or U19675 (N_19675,N_19451,N_19449);
xnor U19676 (N_19676,N_19513,N_19500);
nand U19677 (N_19677,N_19368,N_19373);
and U19678 (N_19678,N_19459,N_19475);
or U19679 (N_19679,N_19445,N_19425);
xor U19680 (N_19680,N_19643,N_19638);
nand U19681 (N_19681,N_19653,N_19637);
nor U19682 (N_19682,N_19609,N_19522);
xor U19683 (N_19683,N_19644,N_19646);
nor U19684 (N_19684,N_19624,N_19599);
nand U19685 (N_19685,N_19550,N_19548);
nand U19686 (N_19686,N_19594,N_19555);
nor U19687 (N_19687,N_19613,N_19543);
xor U19688 (N_19688,N_19662,N_19540);
and U19689 (N_19689,N_19604,N_19631);
or U19690 (N_19690,N_19554,N_19593);
nand U19691 (N_19691,N_19587,N_19607);
or U19692 (N_19692,N_19610,N_19538);
or U19693 (N_19693,N_19619,N_19634);
nor U19694 (N_19694,N_19532,N_19535);
or U19695 (N_19695,N_19645,N_19650);
or U19696 (N_19696,N_19660,N_19561);
and U19697 (N_19697,N_19564,N_19675);
xor U19698 (N_19698,N_19663,N_19545);
or U19699 (N_19699,N_19605,N_19580);
and U19700 (N_19700,N_19616,N_19531);
or U19701 (N_19701,N_19576,N_19617);
nand U19702 (N_19702,N_19556,N_19529);
nand U19703 (N_19703,N_19567,N_19539);
nor U19704 (N_19704,N_19520,N_19591);
nand U19705 (N_19705,N_19665,N_19592);
and U19706 (N_19706,N_19666,N_19589);
or U19707 (N_19707,N_19647,N_19537);
and U19708 (N_19708,N_19523,N_19670);
or U19709 (N_19709,N_19559,N_19602);
nor U19710 (N_19710,N_19575,N_19571);
and U19711 (N_19711,N_19530,N_19661);
nand U19712 (N_19712,N_19611,N_19669);
nor U19713 (N_19713,N_19590,N_19648);
xnor U19714 (N_19714,N_19626,N_19557);
xor U19715 (N_19715,N_19621,N_19572);
and U19716 (N_19716,N_19640,N_19549);
or U19717 (N_19717,N_19521,N_19582);
or U19718 (N_19718,N_19639,N_19632);
nor U19719 (N_19719,N_19652,N_19568);
nor U19720 (N_19720,N_19596,N_19544);
xnor U19721 (N_19721,N_19651,N_19566);
or U19722 (N_19722,N_19668,N_19612);
nor U19723 (N_19723,N_19657,N_19565);
nor U19724 (N_19724,N_19608,N_19581);
nor U19725 (N_19725,N_19678,N_19542);
xnor U19726 (N_19726,N_19658,N_19672);
xor U19727 (N_19727,N_19620,N_19546);
and U19728 (N_19728,N_19563,N_19577);
nand U19729 (N_19729,N_19569,N_19614);
or U19730 (N_19730,N_19671,N_19524);
nand U19731 (N_19731,N_19585,N_19527);
xor U19732 (N_19732,N_19667,N_19601);
nand U19733 (N_19733,N_19558,N_19534);
xor U19734 (N_19734,N_19525,N_19541);
or U19735 (N_19735,N_19654,N_19595);
and U19736 (N_19736,N_19655,N_19600);
and U19737 (N_19737,N_19635,N_19625);
xor U19738 (N_19738,N_19560,N_19664);
xor U19739 (N_19739,N_19578,N_19573);
xor U19740 (N_19740,N_19676,N_19629);
nor U19741 (N_19741,N_19536,N_19627);
xnor U19742 (N_19742,N_19674,N_19533);
and U19743 (N_19743,N_19641,N_19633);
nand U19744 (N_19744,N_19586,N_19618);
or U19745 (N_19745,N_19679,N_19598);
nor U19746 (N_19746,N_19628,N_19579);
and U19747 (N_19747,N_19574,N_19597);
and U19748 (N_19748,N_19553,N_19636);
xor U19749 (N_19749,N_19659,N_19526);
xnor U19750 (N_19750,N_19656,N_19588);
or U19751 (N_19751,N_19528,N_19603);
nand U19752 (N_19752,N_19552,N_19615);
xnor U19753 (N_19753,N_19562,N_19623);
and U19754 (N_19754,N_19630,N_19547);
xnor U19755 (N_19755,N_19622,N_19606);
nor U19756 (N_19756,N_19642,N_19677);
or U19757 (N_19757,N_19584,N_19551);
xnor U19758 (N_19758,N_19583,N_19649);
nor U19759 (N_19759,N_19570,N_19673);
nor U19760 (N_19760,N_19554,N_19563);
and U19761 (N_19761,N_19593,N_19649);
and U19762 (N_19762,N_19609,N_19600);
or U19763 (N_19763,N_19607,N_19603);
nor U19764 (N_19764,N_19569,N_19650);
xor U19765 (N_19765,N_19555,N_19599);
nand U19766 (N_19766,N_19570,N_19532);
xor U19767 (N_19767,N_19593,N_19602);
nor U19768 (N_19768,N_19626,N_19673);
nand U19769 (N_19769,N_19627,N_19651);
and U19770 (N_19770,N_19536,N_19663);
or U19771 (N_19771,N_19636,N_19574);
nand U19772 (N_19772,N_19653,N_19590);
or U19773 (N_19773,N_19634,N_19642);
xnor U19774 (N_19774,N_19551,N_19657);
or U19775 (N_19775,N_19612,N_19618);
xor U19776 (N_19776,N_19537,N_19624);
xor U19777 (N_19777,N_19548,N_19558);
nand U19778 (N_19778,N_19571,N_19629);
nor U19779 (N_19779,N_19653,N_19597);
and U19780 (N_19780,N_19569,N_19529);
and U19781 (N_19781,N_19613,N_19598);
and U19782 (N_19782,N_19655,N_19583);
and U19783 (N_19783,N_19643,N_19567);
nor U19784 (N_19784,N_19635,N_19568);
nand U19785 (N_19785,N_19641,N_19629);
nor U19786 (N_19786,N_19542,N_19602);
and U19787 (N_19787,N_19618,N_19678);
xnor U19788 (N_19788,N_19601,N_19522);
and U19789 (N_19789,N_19576,N_19670);
nand U19790 (N_19790,N_19538,N_19622);
xor U19791 (N_19791,N_19568,N_19554);
or U19792 (N_19792,N_19639,N_19571);
and U19793 (N_19793,N_19665,N_19565);
or U19794 (N_19794,N_19635,N_19575);
xor U19795 (N_19795,N_19596,N_19655);
xnor U19796 (N_19796,N_19568,N_19590);
nor U19797 (N_19797,N_19583,N_19530);
xor U19798 (N_19798,N_19594,N_19582);
xor U19799 (N_19799,N_19529,N_19607);
and U19800 (N_19800,N_19640,N_19596);
nor U19801 (N_19801,N_19647,N_19674);
or U19802 (N_19802,N_19574,N_19594);
and U19803 (N_19803,N_19622,N_19561);
or U19804 (N_19804,N_19637,N_19561);
or U19805 (N_19805,N_19582,N_19618);
or U19806 (N_19806,N_19607,N_19540);
nand U19807 (N_19807,N_19523,N_19644);
xnor U19808 (N_19808,N_19544,N_19547);
nand U19809 (N_19809,N_19679,N_19575);
and U19810 (N_19810,N_19645,N_19570);
and U19811 (N_19811,N_19648,N_19582);
nor U19812 (N_19812,N_19580,N_19658);
xor U19813 (N_19813,N_19626,N_19679);
nor U19814 (N_19814,N_19601,N_19622);
and U19815 (N_19815,N_19617,N_19545);
or U19816 (N_19816,N_19570,N_19629);
nor U19817 (N_19817,N_19597,N_19583);
nand U19818 (N_19818,N_19561,N_19672);
or U19819 (N_19819,N_19588,N_19646);
nor U19820 (N_19820,N_19664,N_19673);
nand U19821 (N_19821,N_19654,N_19524);
and U19822 (N_19822,N_19529,N_19565);
xnor U19823 (N_19823,N_19531,N_19611);
nor U19824 (N_19824,N_19523,N_19521);
or U19825 (N_19825,N_19597,N_19599);
xor U19826 (N_19826,N_19656,N_19646);
and U19827 (N_19827,N_19520,N_19593);
nand U19828 (N_19828,N_19627,N_19535);
nand U19829 (N_19829,N_19631,N_19675);
nand U19830 (N_19830,N_19528,N_19634);
nor U19831 (N_19831,N_19586,N_19551);
nand U19832 (N_19832,N_19545,N_19668);
xnor U19833 (N_19833,N_19650,N_19595);
xnor U19834 (N_19834,N_19538,N_19592);
or U19835 (N_19835,N_19536,N_19586);
and U19836 (N_19836,N_19674,N_19622);
and U19837 (N_19837,N_19665,N_19542);
xnor U19838 (N_19838,N_19564,N_19583);
or U19839 (N_19839,N_19535,N_19596);
xor U19840 (N_19840,N_19709,N_19770);
or U19841 (N_19841,N_19763,N_19800);
nor U19842 (N_19842,N_19805,N_19792);
nor U19843 (N_19843,N_19736,N_19782);
nand U19844 (N_19844,N_19825,N_19707);
nand U19845 (N_19845,N_19704,N_19807);
and U19846 (N_19846,N_19758,N_19822);
nor U19847 (N_19847,N_19780,N_19689);
nand U19848 (N_19848,N_19814,N_19701);
and U19849 (N_19849,N_19731,N_19683);
or U19850 (N_19850,N_19754,N_19796);
nand U19851 (N_19851,N_19708,N_19712);
or U19852 (N_19852,N_19795,N_19793);
xnor U19853 (N_19853,N_19804,N_19775);
and U19854 (N_19854,N_19742,N_19741);
nor U19855 (N_19855,N_19747,N_19786);
and U19856 (N_19856,N_19749,N_19695);
xor U19857 (N_19857,N_19785,N_19729);
xnor U19858 (N_19858,N_19759,N_19691);
or U19859 (N_19859,N_19687,N_19810);
nand U19860 (N_19860,N_19692,N_19788);
nor U19861 (N_19861,N_19718,N_19812);
nor U19862 (N_19862,N_19752,N_19688);
or U19863 (N_19863,N_19756,N_19799);
and U19864 (N_19864,N_19818,N_19737);
xnor U19865 (N_19865,N_19835,N_19738);
nand U19866 (N_19866,N_19686,N_19722);
nand U19867 (N_19867,N_19798,N_19783);
xor U19868 (N_19868,N_19779,N_19784);
and U19869 (N_19869,N_19716,N_19831);
or U19870 (N_19870,N_19816,N_19781);
nor U19871 (N_19871,N_19821,N_19791);
nand U19872 (N_19872,N_19713,N_19829);
nand U19873 (N_19873,N_19778,N_19750);
nor U19874 (N_19874,N_19836,N_19787);
or U19875 (N_19875,N_19817,N_19802);
or U19876 (N_19876,N_19745,N_19790);
and U19877 (N_19877,N_19813,N_19751);
and U19878 (N_19878,N_19703,N_19832);
xor U19879 (N_19879,N_19815,N_19766);
nor U19880 (N_19880,N_19755,N_19808);
and U19881 (N_19881,N_19711,N_19710);
and U19882 (N_19882,N_19803,N_19681);
xor U19883 (N_19883,N_19828,N_19682);
nand U19884 (N_19884,N_19777,N_19839);
nand U19885 (N_19885,N_19762,N_19702);
or U19886 (N_19886,N_19733,N_19757);
and U19887 (N_19887,N_19760,N_19705);
nand U19888 (N_19888,N_19830,N_19684);
or U19889 (N_19889,N_19753,N_19680);
nor U19890 (N_19890,N_19748,N_19726);
or U19891 (N_19891,N_19820,N_19771);
or U19892 (N_19892,N_19697,N_19723);
nand U19893 (N_19893,N_19797,N_19826);
and U19894 (N_19894,N_19724,N_19730);
or U19895 (N_19895,N_19833,N_19706);
or U19896 (N_19896,N_19761,N_19834);
xor U19897 (N_19897,N_19769,N_19740);
nand U19898 (N_19898,N_19714,N_19789);
nand U19899 (N_19899,N_19764,N_19728);
nor U19900 (N_19900,N_19767,N_19698);
nand U19901 (N_19901,N_19720,N_19719);
xor U19902 (N_19902,N_19732,N_19685);
nor U19903 (N_19903,N_19838,N_19693);
xor U19904 (N_19904,N_19774,N_19739);
and U19905 (N_19905,N_19721,N_19837);
xor U19906 (N_19906,N_19823,N_19811);
or U19907 (N_19907,N_19765,N_19735);
and U19908 (N_19908,N_19743,N_19694);
or U19909 (N_19909,N_19824,N_19696);
nand U19910 (N_19910,N_19734,N_19819);
and U19911 (N_19911,N_19776,N_19727);
nor U19912 (N_19912,N_19809,N_19717);
xnor U19913 (N_19913,N_19801,N_19827);
and U19914 (N_19914,N_19725,N_19768);
nand U19915 (N_19915,N_19715,N_19699);
xnor U19916 (N_19916,N_19746,N_19806);
or U19917 (N_19917,N_19773,N_19700);
and U19918 (N_19918,N_19772,N_19744);
nor U19919 (N_19919,N_19690,N_19794);
nand U19920 (N_19920,N_19790,N_19688);
or U19921 (N_19921,N_19688,N_19786);
xnor U19922 (N_19922,N_19730,N_19763);
xnor U19923 (N_19923,N_19775,N_19833);
and U19924 (N_19924,N_19781,N_19837);
nand U19925 (N_19925,N_19697,N_19749);
nor U19926 (N_19926,N_19824,N_19748);
and U19927 (N_19927,N_19742,N_19701);
and U19928 (N_19928,N_19681,N_19770);
nor U19929 (N_19929,N_19764,N_19754);
nor U19930 (N_19930,N_19702,N_19742);
and U19931 (N_19931,N_19780,N_19688);
or U19932 (N_19932,N_19780,N_19800);
and U19933 (N_19933,N_19728,N_19838);
and U19934 (N_19934,N_19709,N_19830);
nor U19935 (N_19935,N_19830,N_19739);
xnor U19936 (N_19936,N_19752,N_19807);
or U19937 (N_19937,N_19704,N_19716);
and U19938 (N_19938,N_19837,N_19766);
nand U19939 (N_19939,N_19782,N_19723);
nor U19940 (N_19940,N_19838,N_19699);
nor U19941 (N_19941,N_19819,N_19750);
and U19942 (N_19942,N_19730,N_19820);
or U19943 (N_19943,N_19744,N_19781);
and U19944 (N_19944,N_19788,N_19777);
nand U19945 (N_19945,N_19777,N_19832);
and U19946 (N_19946,N_19719,N_19816);
or U19947 (N_19947,N_19796,N_19779);
nand U19948 (N_19948,N_19736,N_19738);
nand U19949 (N_19949,N_19751,N_19682);
and U19950 (N_19950,N_19831,N_19765);
xnor U19951 (N_19951,N_19688,N_19825);
nor U19952 (N_19952,N_19797,N_19684);
or U19953 (N_19953,N_19803,N_19785);
xor U19954 (N_19954,N_19813,N_19703);
and U19955 (N_19955,N_19714,N_19722);
or U19956 (N_19956,N_19699,N_19759);
and U19957 (N_19957,N_19811,N_19821);
nand U19958 (N_19958,N_19812,N_19725);
or U19959 (N_19959,N_19747,N_19727);
nand U19960 (N_19960,N_19813,N_19767);
or U19961 (N_19961,N_19701,N_19687);
xnor U19962 (N_19962,N_19756,N_19753);
or U19963 (N_19963,N_19726,N_19765);
nand U19964 (N_19964,N_19814,N_19790);
and U19965 (N_19965,N_19806,N_19714);
xnor U19966 (N_19966,N_19710,N_19783);
nor U19967 (N_19967,N_19796,N_19727);
or U19968 (N_19968,N_19691,N_19686);
xor U19969 (N_19969,N_19777,N_19766);
nand U19970 (N_19970,N_19740,N_19800);
nand U19971 (N_19971,N_19729,N_19698);
xor U19972 (N_19972,N_19687,N_19782);
nor U19973 (N_19973,N_19836,N_19732);
xor U19974 (N_19974,N_19823,N_19754);
xnor U19975 (N_19975,N_19721,N_19828);
and U19976 (N_19976,N_19736,N_19804);
xor U19977 (N_19977,N_19755,N_19706);
xnor U19978 (N_19978,N_19756,N_19716);
nor U19979 (N_19979,N_19805,N_19793);
nand U19980 (N_19980,N_19829,N_19779);
nand U19981 (N_19981,N_19810,N_19773);
nor U19982 (N_19982,N_19759,N_19833);
and U19983 (N_19983,N_19789,N_19806);
xnor U19984 (N_19984,N_19798,N_19772);
and U19985 (N_19985,N_19707,N_19691);
xnor U19986 (N_19986,N_19772,N_19721);
xnor U19987 (N_19987,N_19768,N_19729);
nor U19988 (N_19988,N_19712,N_19789);
nor U19989 (N_19989,N_19838,N_19750);
nand U19990 (N_19990,N_19831,N_19712);
nor U19991 (N_19991,N_19784,N_19793);
nor U19992 (N_19992,N_19758,N_19773);
and U19993 (N_19993,N_19826,N_19693);
and U19994 (N_19994,N_19699,N_19773);
nand U19995 (N_19995,N_19823,N_19738);
nor U19996 (N_19996,N_19764,N_19717);
xor U19997 (N_19997,N_19739,N_19821);
nand U19998 (N_19998,N_19748,N_19730);
nor U19999 (N_19999,N_19814,N_19773);
xor UO_0 (O_0,N_19886,N_19843);
or UO_1 (O_1,N_19877,N_19879);
nand UO_2 (O_2,N_19899,N_19991);
nor UO_3 (O_3,N_19890,N_19895);
xor UO_4 (O_4,N_19876,N_19869);
or UO_5 (O_5,N_19903,N_19984);
nor UO_6 (O_6,N_19878,N_19936);
xor UO_7 (O_7,N_19957,N_19953);
nand UO_8 (O_8,N_19977,N_19857);
or UO_9 (O_9,N_19929,N_19996);
nand UO_10 (O_10,N_19943,N_19864);
nand UO_11 (O_11,N_19938,N_19845);
nor UO_12 (O_12,N_19997,N_19891);
nor UO_13 (O_13,N_19889,N_19853);
xnor UO_14 (O_14,N_19884,N_19873);
and UO_15 (O_15,N_19948,N_19999);
nand UO_16 (O_16,N_19990,N_19969);
and UO_17 (O_17,N_19900,N_19874);
nor UO_18 (O_18,N_19954,N_19970);
xnor UO_19 (O_19,N_19961,N_19920);
nor UO_20 (O_20,N_19897,N_19922);
or UO_21 (O_21,N_19987,N_19937);
xnor UO_22 (O_22,N_19978,N_19855);
nand UO_23 (O_23,N_19946,N_19940);
nand UO_24 (O_24,N_19983,N_19915);
nor UO_25 (O_25,N_19882,N_19910);
nand UO_26 (O_26,N_19958,N_19973);
nand UO_27 (O_27,N_19887,N_19945);
nor UO_28 (O_28,N_19902,N_19858);
nand UO_29 (O_29,N_19947,N_19971);
or UO_30 (O_30,N_19912,N_19932);
or UO_31 (O_31,N_19911,N_19914);
xor UO_32 (O_32,N_19979,N_19859);
xor UO_33 (O_33,N_19974,N_19840);
xor UO_34 (O_34,N_19944,N_19955);
nand UO_35 (O_35,N_19880,N_19986);
and UO_36 (O_36,N_19941,N_19898);
or UO_37 (O_37,N_19951,N_19863);
or UO_38 (O_38,N_19989,N_19933);
and UO_39 (O_39,N_19975,N_19885);
xnor UO_40 (O_40,N_19993,N_19988);
xor UO_41 (O_41,N_19956,N_19842);
or UO_42 (O_42,N_19994,N_19949);
xor UO_43 (O_43,N_19906,N_19847);
and UO_44 (O_44,N_19925,N_19856);
xnor UO_45 (O_45,N_19868,N_19872);
and UO_46 (O_46,N_19942,N_19992);
and UO_47 (O_47,N_19883,N_19901);
nand UO_48 (O_48,N_19867,N_19927);
nor UO_49 (O_49,N_19963,N_19921);
xor UO_50 (O_50,N_19981,N_19862);
nor UO_51 (O_51,N_19917,N_19908);
or UO_52 (O_52,N_19923,N_19950);
nor UO_53 (O_53,N_19904,N_19870);
xor UO_54 (O_54,N_19967,N_19854);
and UO_55 (O_55,N_19875,N_19968);
or UO_56 (O_56,N_19959,N_19844);
and UO_57 (O_57,N_19964,N_19960);
and UO_58 (O_58,N_19888,N_19935);
or UO_59 (O_59,N_19965,N_19928);
nand UO_60 (O_60,N_19860,N_19985);
or UO_61 (O_61,N_19892,N_19934);
or UO_62 (O_62,N_19861,N_19966);
nand UO_63 (O_63,N_19907,N_19918);
nor UO_64 (O_64,N_19998,N_19952);
xor UO_65 (O_65,N_19893,N_19852);
xor UO_66 (O_66,N_19850,N_19841);
and UO_67 (O_67,N_19846,N_19930);
xor UO_68 (O_68,N_19926,N_19913);
and UO_69 (O_69,N_19916,N_19894);
xor UO_70 (O_70,N_19976,N_19995);
and UO_71 (O_71,N_19972,N_19848);
nor UO_72 (O_72,N_19982,N_19939);
nand UO_73 (O_73,N_19851,N_19896);
or UO_74 (O_74,N_19924,N_19866);
and UO_75 (O_75,N_19905,N_19962);
and UO_76 (O_76,N_19849,N_19871);
or UO_77 (O_77,N_19909,N_19865);
and UO_78 (O_78,N_19980,N_19919);
xor UO_79 (O_79,N_19931,N_19881);
and UO_80 (O_80,N_19969,N_19861);
nor UO_81 (O_81,N_19943,N_19856);
nor UO_82 (O_82,N_19843,N_19903);
nand UO_83 (O_83,N_19929,N_19855);
or UO_84 (O_84,N_19947,N_19932);
or UO_85 (O_85,N_19880,N_19876);
nor UO_86 (O_86,N_19866,N_19958);
and UO_87 (O_87,N_19939,N_19998);
xnor UO_88 (O_88,N_19948,N_19856);
or UO_89 (O_89,N_19942,N_19874);
nor UO_90 (O_90,N_19956,N_19851);
nor UO_91 (O_91,N_19908,N_19900);
and UO_92 (O_92,N_19897,N_19998);
xor UO_93 (O_93,N_19891,N_19895);
xnor UO_94 (O_94,N_19891,N_19847);
and UO_95 (O_95,N_19876,N_19925);
nor UO_96 (O_96,N_19892,N_19983);
and UO_97 (O_97,N_19976,N_19991);
or UO_98 (O_98,N_19855,N_19882);
xor UO_99 (O_99,N_19990,N_19912);
nor UO_100 (O_100,N_19916,N_19842);
nand UO_101 (O_101,N_19867,N_19879);
or UO_102 (O_102,N_19891,N_19843);
or UO_103 (O_103,N_19971,N_19924);
and UO_104 (O_104,N_19933,N_19898);
nand UO_105 (O_105,N_19919,N_19894);
and UO_106 (O_106,N_19936,N_19911);
nand UO_107 (O_107,N_19967,N_19894);
or UO_108 (O_108,N_19849,N_19900);
and UO_109 (O_109,N_19949,N_19929);
xor UO_110 (O_110,N_19910,N_19923);
or UO_111 (O_111,N_19936,N_19958);
nor UO_112 (O_112,N_19922,N_19935);
nand UO_113 (O_113,N_19969,N_19892);
or UO_114 (O_114,N_19999,N_19895);
and UO_115 (O_115,N_19985,N_19960);
or UO_116 (O_116,N_19909,N_19912);
nor UO_117 (O_117,N_19887,N_19885);
or UO_118 (O_118,N_19965,N_19952);
or UO_119 (O_119,N_19942,N_19905);
nor UO_120 (O_120,N_19912,N_19936);
xor UO_121 (O_121,N_19852,N_19926);
xnor UO_122 (O_122,N_19920,N_19971);
xnor UO_123 (O_123,N_19909,N_19977);
nand UO_124 (O_124,N_19970,N_19884);
nand UO_125 (O_125,N_19977,N_19879);
xnor UO_126 (O_126,N_19944,N_19935);
or UO_127 (O_127,N_19901,N_19856);
and UO_128 (O_128,N_19850,N_19997);
or UO_129 (O_129,N_19943,N_19851);
nand UO_130 (O_130,N_19947,N_19840);
or UO_131 (O_131,N_19949,N_19882);
nand UO_132 (O_132,N_19855,N_19918);
and UO_133 (O_133,N_19933,N_19967);
nor UO_134 (O_134,N_19901,N_19911);
nor UO_135 (O_135,N_19990,N_19920);
nand UO_136 (O_136,N_19870,N_19897);
or UO_137 (O_137,N_19869,N_19947);
nor UO_138 (O_138,N_19895,N_19954);
xor UO_139 (O_139,N_19867,N_19942);
or UO_140 (O_140,N_19872,N_19898);
or UO_141 (O_141,N_19974,N_19898);
and UO_142 (O_142,N_19989,N_19927);
or UO_143 (O_143,N_19990,N_19864);
or UO_144 (O_144,N_19875,N_19856);
xnor UO_145 (O_145,N_19906,N_19886);
nor UO_146 (O_146,N_19886,N_19961);
and UO_147 (O_147,N_19966,N_19905);
xor UO_148 (O_148,N_19871,N_19842);
or UO_149 (O_149,N_19902,N_19853);
xor UO_150 (O_150,N_19888,N_19882);
nand UO_151 (O_151,N_19865,N_19846);
and UO_152 (O_152,N_19978,N_19915);
nand UO_153 (O_153,N_19943,N_19886);
nor UO_154 (O_154,N_19995,N_19929);
or UO_155 (O_155,N_19840,N_19883);
or UO_156 (O_156,N_19968,N_19930);
or UO_157 (O_157,N_19872,N_19935);
nor UO_158 (O_158,N_19936,N_19855);
nor UO_159 (O_159,N_19895,N_19845);
nor UO_160 (O_160,N_19890,N_19873);
nor UO_161 (O_161,N_19841,N_19963);
and UO_162 (O_162,N_19896,N_19903);
and UO_163 (O_163,N_19851,N_19938);
or UO_164 (O_164,N_19883,N_19855);
xor UO_165 (O_165,N_19884,N_19947);
and UO_166 (O_166,N_19963,N_19913);
or UO_167 (O_167,N_19977,N_19970);
nor UO_168 (O_168,N_19987,N_19890);
nor UO_169 (O_169,N_19882,N_19912);
nor UO_170 (O_170,N_19852,N_19952);
nand UO_171 (O_171,N_19949,N_19857);
or UO_172 (O_172,N_19870,N_19889);
nand UO_173 (O_173,N_19841,N_19864);
nor UO_174 (O_174,N_19937,N_19968);
xor UO_175 (O_175,N_19856,N_19858);
nor UO_176 (O_176,N_19998,N_19862);
nor UO_177 (O_177,N_19943,N_19991);
and UO_178 (O_178,N_19960,N_19949);
or UO_179 (O_179,N_19975,N_19974);
nand UO_180 (O_180,N_19931,N_19869);
xor UO_181 (O_181,N_19996,N_19964);
nand UO_182 (O_182,N_19963,N_19869);
xnor UO_183 (O_183,N_19883,N_19847);
or UO_184 (O_184,N_19866,N_19907);
xor UO_185 (O_185,N_19892,N_19926);
xnor UO_186 (O_186,N_19978,N_19951);
nand UO_187 (O_187,N_19969,N_19989);
xor UO_188 (O_188,N_19962,N_19843);
xor UO_189 (O_189,N_19984,N_19906);
and UO_190 (O_190,N_19995,N_19869);
and UO_191 (O_191,N_19938,N_19843);
nor UO_192 (O_192,N_19852,N_19862);
xnor UO_193 (O_193,N_19843,N_19974);
nor UO_194 (O_194,N_19968,N_19941);
or UO_195 (O_195,N_19848,N_19857);
nand UO_196 (O_196,N_19890,N_19989);
or UO_197 (O_197,N_19989,N_19844);
nor UO_198 (O_198,N_19989,N_19889);
and UO_199 (O_199,N_19961,N_19916);
xnor UO_200 (O_200,N_19911,N_19912);
nor UO_201 (O_201,N_19869,N_19872);
and UO_202 (O_202,N_19949,N_19861);
and UO_203 (O_203,N_19841,N_19918);
xor UO_204 (O_204,N_19860,N_19991);
nand UO_205 (O_205,N_19933,N_19841);
nand UO_206 (O_206,N_19931,N_19954);
and UO_207 (O_207,N_19971,N_19894);
xor UO_208 (O_208,N_19954,N_19912);
and UO_209 (O_209,N_19935,N_19893);
or UO_210 (O_210,N_19893,N_19983);
nand UO_211 (O_211,N_19924,N_19948);
nor UO_212 (O_212,N_19961,N_19963);
xor UO_213 (O_213,N_19870,N_19946);
and UO_214 (O_214,N_19887,N_19857);
nor UO_215 (O_215,N_19990,N_19985);
nor UO_216 (O_216,N_19986,N_19927);
nand UO_217 (O_217,N_19881,N_19983);
or UO_218 (O_218,N_19856,N_19900);
nand UO_219 (O_219,N_19987,N_19902);
xnor UO_220 (O_220,N_19888,N_19956);
and UO_221 (O_221,N_19894,N_19974);
xor UO_222 (O_222,N_19870,N_19913);
nand UO_223 (O_223,N_19937,N_19913);
or UO_224 (O_224,N_19967,N_19889);
nand UO_225 (O_225,N_19872,N_19847);
nor UO_226 (O_226,N_19986,N_19911);
nor UO_227 (O_227,N_19996,N_19983);
nor UO_228 (O_228,N_19919,N_19952);
xnor UO_229 (O_229,N_19924,N_19933);
xnor UO_230 (O_230,N_19994,N_19948);
nand UO_231 (O_231,N_19971,N_19917);
or UO_232 (O_232,N_19973,N_19931);
and UO_233 (O_233,N_19923,N_19904);
nor UO_234 (O_234,N_19923,N_19986);
nor UO_235 (O_235,N_19858,N_19950);
xor UO_236 (O_236,N_19963,N_19851);
or UO_237 (O_237,N_19978,N_19895);
and UO_238 (O_238,N_19864,N_19972);
and UO_239 (O_239,N_19900,N_19929);
or UO_240 (O_240,N_19966,N_19928);
xor UO_241 (O_241,N_19864,N_19949);
xor UO_242 (O_242,N_19930,N_19972);
or UO_243 (O_243,N_19861,N_19891);
or UO_244 (O_244,N_19882,N_19989);
nand UO_245 (O_245,N_19916,N_19904);
nor UO_246 (O_246,N_19986,N_19906);
or UO_247 (O_247,N_19963,N_19857);
xnor UO_248 (O_248,N_19902,N_19894);
xnor UO_249 (O_249,N_19854,N_19886);
nand UO_250 (O_250,N_19947,N_19885);
or UO_251 (O_251,N_19991,N_19869);
nand UO_252 (O_252,N_19979,N_19942);
nor UO_253 (O_253,N_19846,N_19847);
nor UO_254 (O_254,N_19933,N_19997);
or UO_255 (O_255,N_19910,N_19855);
and UO_256 (O_256,N_19857,N_19953);
nor UO_257 (O_257,N_19921,N_19923);
and UO_258 (O_258,N_19913,N_19910);
nand UO_259 (O_259,N_19969,N_19992);
and UO_260 (O_260,N_19888,N_19951);
and UO_261 (O_261,N_19889,N_19892);
nand UO_262 (O_262,N_19930,N_19997);
nor UO_263 (O_263,N_19992,N_19915);
or UO_264 (O_264,N_19923,N_19851);
nand UO_265 (O_265,N_19840,N_19916);
and UO_266 (O_266,N_19843,N_19893);
or UO_267 (O_267,N_19940,N_19887);
nor UO_268 (O_268,N_19840,N_19959);
nand UO_269 (O_269,N_19905,N_19912);
or UO_270 (O_270,N_19875,N_19909);
or UO_271 (O_271,N_19866,N_19869);
or UO_272 (O_272,N_19968,N_19848);
xor UO_273 (O_273,N_19943,N_19968);
nor UO_274 (O_274,N_19842,N_19937);
nand UO_275 (O_275,N_19942,N_19978);
and UO_276 (O_276,N_19948,N_19889);
or UO_277 (O_277,N_19920,N_19881);
or UO_278 (O_278,N_19847,N_19977);
and UO_279 (O_279,N_19907,N_19900);
and UO_280 (O_280,N_19940,N_19947);
nand UO_281 (O_281,N_19848,N_19903);
nand UO_282 (O_282,N_19885,N_19984);
or UO_283 (O_283,N_19881,N_19972);
and UO_284 (O_284,N_19847,N_19998);
nor UO_285 (O_285,N_19878,N_19978);
nor UO_286 (O_286,N_19988,N_19977);
xor UO_287 (O_287,N_19934,N_19929);
and UO_288 (O_288,N_19974,N_19916);
nor UO_289 (O_289,N_19958,N_19944);
nand UO_290 (O_290,N_19903,N_19908);
xor UO_291 (O_291,N_19919,N_19973);
or UO_292 (O_292,N_19933,N_19958);
and UO_293 (O_293,N_19889,N_19925);
or UO_294 (O_294,N_19910,N_19875);
and UO_295 (O_295,N_19914,N_19843);
nor UO_296 (O_296,N_19998,N_19948);
and UO_297 (O_297,N_19887,N_19951);
nand UO_298 (O_298,N_19947,N_19962);
and UO_299 (O_299,N_19957,N_19879);
or UO_300 (O_300,N_19906,N_19989);
nand UO_301 (O_301,N_19942,N_19915);
and UO_302 (O_302,N_19867,N_19953);
nand UO_303 (O_303,N_19907,N_19977);
or UO_304 (O_304,N_19919,N_19884);
xnor UO_305 (O_305,N_19973,N_19942);
and UO_306 (O_306,N_19891,N_19850);
nand UO_307 (O_307,N_19849,N_19935);
nor UO_308 (O_308,N_19949,N_19917);
and UO_309 (O_309,N_19844,N_19866);
or UO_310 (O_310,N_19971,N_19975);
xnor UO_311 (O_311,N_19864,N_19925);
or UO_312 (O_312,N_19842,N_19858);
xor UO_313 (O_313,N_19965,N_19962);
and UO_314 (O_314,N_19928,N_19980);
xnor UO_315 (O_315,N_19961,N_19929);
or UO_316 (O_316,N_19929,N_19953);
or UO_317 (O_317,N_19888,N_19877);
nand UO_318 (O_318,N_19883,N_19958);
nor UO_319 (O_319,N_19980,N_19962);
xnor UO_320 (O_320,N_19960,N_19931);
nand UO_321 (O_321,N_19956,N_19844);
nand UO_322 (O_322,N_19896,N_19866);
nand UO_323 (O_323,N_19956,N_19954);
and UO_324 (O_324,N_19980,N_19979);
xor UO_325 (O_325,N_19985,N_19949);
nand UO_326 (O_326,N_19939,N_19974);
or UO_327 (O_327,N_19946,N_19964);
nor UO_328 (O_328,N_19871,N_19861);
nand UO_329 (O_329,N_19996,N_19854);
xor UO_330 (O_330,N_19840,N_19917);
xor UO_331 (O_331,N_19957,N_19844);
nand UO_332 (O_332,N_19966,N_19866);
nand UO_333 (O_333,N_19857,N_19884);
and UO_334 (O_334,N_19987,N_19914);
nand UO_335 (O_335,N_19965,N_19877);
nor UO_336 (O_336,N_19852,N_19913);
xnor UO_337 (O_337,N_19925,N_19986);
nand UO_338 (O_338,N_19944,N_19940);
nor UO_339 (O_339,N_19952,N_19989);
or UO_340 (O_340,N_19972,N_19979);
nand UO_341 (O_341,N_19925,N_19884);
xnor UO_342 (O_342,N_19873,N_19858);
nor UO_343 (O_343,N_19966,N_19869);
or UO_344 (O_344,N_19889,N_19982);
xor UO_345 (O_345,N_19864,N_19980);
xor UO_346 (O_346,N_19972,N_19977);
xor UO_347 (O_347,N_19932,N_19915);
and UO_348 (O_348,N_19930,N_19874);
nand UO_349 (O_349,N_19910,N_19983);
and UO_350 (O_350,N_19980,N_19902);
and UO_351 (O_351,N_19999,N_19997);
and UO_352 (O_352,N_19872,N_19865);
nand UO_353 (O_353,N_19877,N_19878);
or UO_354 (O_354,N_19847,N_19954);
xnor UO_355 (O_355,N_19966,N_19958);
nand UO_356 (O_356,N_19930,N_19840);
nand UO_357 (O_357,N_19889,N_19840);
nand UO_358 (O_358,N_19875,N_19945);
or UO_359 (O_359,N_19955,N_19991);
nor UO_360 (O_360,N_19973,N_19966);
and UO_361 (O_361,N_19905,N_19915);
and UO_362 (O_362,N_19899,N_19950);
nor UO_363 (O_363,N_19918,N_19944);
or UO_364 (O_364,N_19931,N_19917);
nor UO_365 (O_365,N_19962,N_19873);
nor UO_366 (O_366,N_19879,N_19847);
and UO_367 (O_367,N_19929,N_19984);
or UO_368 (O_368,N_19993,N_19978);
xnor UO_369 (O_369,N_19949,N_19940);
and UO_370 (O_370,N_19958,N_19849);
or UO_371 (O_371,N_19897,N_19844);
or UO_372 (O_372,N_19874,N_19940);
and UO_373 (O_373,N_19931,N_19873);
and UO_374 (O_374,N_19865,N_19954);
and UO_375 (O_375,N_19984,N_19982);
nand UO_376 (O_376,N_19848,N_19959);
nor UO_377 (O_377,N_19930,N_19947);
and UO_378 (O_378,N_19851,N_19889);
nor UO_379 (O_379,N_19870,N_19879);
or UO_380 (O_380,N_19942,N_19916);
or UO_381 (O_381,N_19966,N_19923);
nand UO_382 (O_382,N_19947,N_19861);
xnor UO_383 (O_383,N_19989,N_19968);
nand UO_384 (O_384,N_19977,N_19952);
nand UO_385 (O_385,N_19996,N_19959);
xnor UO_386 (O_386,N_19953,N_19919);
nor UO_387 (O_387,N_19877,N_19849);
or UO_388 (O_388,N_19861,N_19919);
nor UO_389 (O_389,N_19945,N_19964);
and UO_390 (O_390,N_19985,N_19962);
or UO_391 (O_391,N_19948,N_19917);
nor UO_392 (O_392,N_19906,N_19915);
nor UO_393 (O_393,N_19922,N_19908);
xor UO_394 (O_394,N_19878,N_19934);
and UO_395 (O_395,N_19847,N_19947);
nand UO_396 (O_396,N_19934,N_19952);
or UO_397 (O_397,N_19985,N_19996);
nor UO_398 (O_398,N_19903,N_19997);
nand UO_399 (O_399,N_19850,N_19968);
nor UO_400 (O_400,N_19918,N_19946);
xnor UO_401 (O_401,N_19938,N_19909);
nor UO_402 (O_402,N_19863,N_19963);
and UO_403 (O_403,N_19978,N_19930);
or UO_404 (O_404,N_19843,N_19915);
xor UO_405 (O_405,N_19997,N_19902);
or UO_406 (O_406,N_19973,N_19935);
or UO_407 (O_407,N_19978,N_19963);
and UO_408 (O_408,N_19890,N_19996);
nand UO_409 (O_409,N_19899,N_19984);
nor UO_410 (O_410,N_19920,N_19969);
and UO_411 (O_411,N_19936,N_19913);
nand UO_412 (O_412,N_19878,N_19890);
and UO_413 (O_413,N_19906,N_19845);
nor UO_414 (O_414,N_19898,N_19891);
xnor UO_415 (O_415,N_19924,N_19904);
nor UO_416 (O_416,N_19863,N_19922);
or UO_417 (O_417,N_19957,N_19887);
nor UO_418 (O_418,N_19881,N_19862);
nand UO_419 (O_419,N_19914,N_19869);
xor UO_420 (O_420,N_19852,N_19920);
nor UO_421 (O_421,N_19934,N_19982);
nor UO_422 (O_422,N_19899,N_19983);
and UO_423 (O_423,N_19848,N_19934);
or UO_424 (O_424,N_19897,N_19886);
nor UO_425 (O_425,N_19967,N_19998);
and UO_426 (O_426,N_19873,N_19889);
and UO_427 (O_427,N_19960,N_19894);
xnor UO_428 (O_428,N_19882,N_19963);
and UO_429 (O_429,N_19847,N_19909);
nand UO_430 (O_430,N_19865,N_19907);
xnor UO_431 (O_431,N_19874,N_19865);
nor UO_432 (O_432,N_19885,N_19897);
nand UO_433 (O_433,N_19927,N_19877);
or UO_434 (O_434,N_19870,N_19925);
xnor UO_435 (O_435,N_19943,N_19981);
xor UO_436 (O_436,N_19883,N_19982);
nand UO_437 (O_437,N_19901,N_19895);
and UO_438 (O_438,N_19878,N_19969);
xor UO_439 (O_439,N_19869,N_19867);
and UO_440 (O_440,N_19864,N_19929);
nand UO_441 (O_441,N_19980,N_19991);
nand UO_442 (O_442,N_19975,N_19933);
or UO_443 (O_443,N_19880,N_19927);
nor UO_444 (O_444,N_19987,N_19977);
and UO_445 (O_445,N_19903,N_19972);
xor UO_446 (O_446,N_19940,N_19920);
or UO_447 (O_447,N_19874,N_19992);
and UO_448 (O_448,N_19991,N_19959);
and UO_449 (O_449,N_19922,N_19973);
nand UO_450 (O_450,N_19892,N_19868);
nand UO_451 (O_451,N_19912,N_19993);
nand UO_452 (O_452,N_19924,N_19912);
and UO_453 (O_453,N_19969,N_19914);
xnor UO_454 (O_454,N_19841,N_19961);
or UO_455 (O_455,N_19928,N_19859);
nand UO_456 (O_456,N_19951,N_19860);
and UO_457 (O_457,N_19848,N_19962);
nand UO_458 (O_458,N_19942,N_19946);
or UO_459 (O_459,N_19975,N_19988);
xor UO_460 (O_460,N_19874,N_19912);
and UO_461 (O_461,N_19978,N_19923);
nand UO_462 (O_462,N_19873,N_19940);
nor UO_463 (O_463,N_19844,N_19898);
and UO_464 (O_464,N_19884,N_19979);
xnor UO_465 (O_465,N_19928,N_19909);
nand UO_466 (O_466,N_19986,N_19957);
nor UO_467 (O_467,N_19981,N_19976);
and UO_468 (O_468,N_19876,N_19997);
xnor UO_469 (O_469,N_19967,N_19980);
and UO_470 (O_470,N_19982,N_19962);
nand UO_471 (O_471,N_19920,N_19911);
xnor UO_472 (O_472,N_19980,N_19916);
nand UO_473 (O_473,N_19919,N_19967);
nor UO_474 (O_474,N_19929,N_19911);
or UO_475 (O_475,N_19870,N_19841);
and UO_476 (O_476,N_19908,N_19984);
and UO_477 (O_477,N_19969,N_19868);
and UO_478 (O_478,N_19875,N_19892);
or UO_479 (O_479,N_19975,N_19904);
xnor UO_480 (O_480,N_19936,N_19962);
nor UO_481 (O_481,N_19903,N_19964);
xnor UO_482 (O_482,N_19945,N_19969);
and UO_483 (O_483,N_19947,N_19843);
nand UO_484 (O_484,N_19911,N_19899);
xor UO_485 (O_485,N_19991,N_19944);
and UO_486 (O_486,N_19848,N_19878);
and UO_487 (O_487,N_19870,N_19859);
xnor UO_488 (O_488,N_19995,N_19930);
nor UO_489 (O_489,N_19844,N_19988);
nor UO_490 (O_490,N_19872,N_19854);
nand UO_491 (O_491,N_19862,N_19931);
nand UO_492 (O_492,N_19872,N_19946);
xor UO_493 (O_493,N_19933,N_19876);
or UO_494 (O_494,N_19889,N_19929);
and UO_495 (O_495,N_19922,N_19972);
nor UO_496 (O_496,N_19927,N_19954);
or UO_497 (O_497,N_19852,N_19957);
xnor UO_498 (O_498,N_19841,N_19855);
and UO_499 (O_499,N_19911,N_19921);
or UO_500 (O_500,N_19904,N_19976);
or UO_501 (O_501,N_19882,N_19960);
nor UO_502 (O_502,N_19938,N_19940);
nand UO_503 (O_503,N_19893,N_19858);
nand UO_504 (O_504,N_19947,N_19975);
nand UO_505 (O_505,N_19909,N_19885);
nand UO_506 (O_506,N_19877,N_19891);
and UO_507 (O_507,N_19949,N_19916);
nor UO_508 (O_508,N_19982,N_19879);
and UO_509 (O_509,N_19876,N_19883);
or UO_510 (O_510,N_19957,N_19871);
nand UO_511 (O_511,N_19867,N_19915);
nor UO_512 (O_512,N_19841,N_19985);
nand UO_513 (O_513,N_19855,N_19990);
and UO_514 (O_514,N_19907,N_19858);
xnor UO_515 (O_515,N_19979,N_19994);
or UO_516 (O_516,N_19941,N_19986);
nand UO_517 (O_517,N_19933,N_19995);
xor UO_518 (O_518,N_19960,N_19976);
or UO_519 (O_519,N_19863,N_19904);
or UO_520 (O_520,N_19875,N_19905);
nand UO_521 (O_521,N_19864,N_19934);
nand UO_522 (O_522,N_19971,N_19961);
nand UO_523 (O_523,N_19934,N_19911);
and UO_524 (O_524,N_19983,N_19857);
and UO_525 (O_525,N_19962,N_19934);
xor UO_526 (O_526,N_19967,N_19861);
nand UO_527 (O_527,N_19926,N_19963);
nor UO_528 (O_528,N_19842,N_19882);
nand UO_529 (O_529,N_19848,N_19977);
nand UO_530 (O_530,N_19949,N_19850);
xor UO_531 (O_531,N_19923,N_19871);
or UO_532 (O_532,N_19854,N_19914);
xnor UO_533 (O_533,N_19953,N_19951);
xor UO_534 (O_534,N_19996,N_19972);
nand UO_535 (O_535,N_19960,N_19922);
xnor UO_536 (O_536,N_19966,N_19871);
or UO_537 (O_537,N_19955,N_19978);
and UO_538 (O_538,N_19984,N_19950);
nand UO_539 (O_539,N_19951,N_19942);
nor UO_540 (O_540,N_19971,N_19878);
nand UO_541 (O_541,N_19964,N_19921);
nor UO_542 (O_542,N_19953,N_19996);
and UO_543 (O_543,N_19896,N_19930);
xnor UO_544 (O_544,N_19843,N_19907);
nand UO_545 (O_545,N_19963,N_19964);
nand UO_546 (O_546,N_19964,N_19900);
or UO_547 (O_547,N_19851,N_19913);
nand UO_548 (O_548,N_19988,N_19866);
nand UO_549 (O_549,N_19847,N_19916);
and UO_550 (O_550,N_19860,N_19889);
xnor UO_551 (O_551,N_19870,N_19852);
and UO_552 (O_552,N_19976,N_19913);
or UO_553 (O_553,N_19941,N_19906);
nor UO_554 (O_554,N_19924,N_19846);
and UO_555 (O_555,N_19873,N_19979);
or UO_556 (O_556,N_19887,N_19950);
nand UO_557 (O_557,N_19952,N_19904);
nor UO_558 (O_558,N_19996,N_19884);
nand UO_559 (O_559,N_19841,N_19847);
or UO_560 (O_560,N_19972,N_19897);
or UO_561 (O_561,N_19954,N_19911);
nand UO_562 (O_562,N_19915,N_19861);
xnor UO_563 (O_563,N_19922,N_19848);
xnor UO_564 (O_564,N_19887,N_19872);
and UO_565 (O_565,N_19918,N_19864);
xor UO_566 (O_566,N_19871,N_19987);
xnor UO_567 (O_567,N_19931,N_19900);
nand UO_568 (O_568,N_19878,N_19913);
xnor UO_569 (O_569,N_19934,N_19891);
xnor UO_570 (O_570,N_19927,N_19922);
nand UO_571 (O_571,N_19990,N_19956);
nand UO_572 (O_572,N_19867,N_19970);
xnor UO_573 (O_573,N_19912,N_19943);
or UO_574 (O_574,N_19993,N_19855);
nand UO_575 (O_575,N_19858,N_19845);
and UO_576 (O_576,N_19846,N_19895);
or UO_577 (O_577,N_19987,N_19886);
or UO_578 (O_578,N_19883,N_19994);
nand UO_579 (O_579,N_19916,N_19896);
xor UO_580 (O_580,N_19848,N_19898);
or UO_581 (O_581,N_19864,N_19946);
xnor UO_582 (O_582,N_19857,N_19859);
nand UO_583 (O_583,N_19888,N_19962);
xnor UO_584 (O_584,N_19903,N_19941);
nand UO_585 (O_585,N_19919,N_19881);
nor UO_586 (O_586,N_19996,N_19863);
xnor UO_587 (O_587,N_19842,N_19952);
nand UO_588 (O_588,N_19865,N_19994);
or UO_589 (O_589,N_19975,N_19870);
or UO_590 (O_590,N_19915,N_19878);
xor UO_591 (O_591,N_19894,N_19850);
and UO_592 (O_592,N_19846,N_19929);
xnor UO_593 (O_593,N_19847,N_19960);
or UO_594 (O_594,N_19881,N_19971);
xor UO_595 (O_595,N_19957,N_19974);
nand UO_596 (O_596,N_19883,N_19894);
nand UO_597 (O_597,N_19970,N_19924);
nor UO_598 (O_598,N_19962,N_19916);
xnor UO_599 (O_599,N_19924,N_19930);
nor UO_600 (O_600,N_19896,N_19961);
xor UO_601 (O_601,N_19851,N_19928);
nand UO_602 (O_602,N_19861,N_19850);
xor UO_603 (O_603,N_19884,N_19893);
or UO_604 (O_604,N_19994,N_19868);
and UO_605 (O_605,N_19960,N_19978);
or UO_606 (O_606,N_19988,N_19949);
and UO_607 (O_607,N_19956,N_19845);
nand UO_608 (O_608,N_19866,N_19894);
or UO_609 (O_609,N_19881,N_19879);
and UO_610 (O_610,N_19846,N_19913);
or UO_611 (O_611,N_19893,N_19997);
xnor UO_612 (O_612,N_19958,N_19975);
or UO_613 (O_613,N_19889,N_19862);
nor UO_614 (O_614,N_19913,N_19893);
or UO_615 (O_615,N_19872,N_19893);
nor UO_616 (O_616,N_19954,N_19948);
or UO_617 (O_617,N_19891,N_19932);
nor UO_618 (O_618,N_19867,N_19893);
or UO_619 (O_619,N_19905,N_19997);
and UO_620 (O_620,N_19923,N_19897);
nor UO_621 (O_621,N_19962,N_19887);
nor UO_622 (O_622,N_19883,N_19932);
and UO_623 (O_623,N_19843,N_19862);
and UO_624 (O_624,N_19985,N_19941);
and UO_625 (O_625,N_19858,N_19897);
nand UO_626 (O_626,N_19916,N_19965);
nand UO_627 (O_627,N_19938,N_19924);
or UO_628 (O_628,N_19957,N_19893);
nand UO_629 (O_629,N_19870,N_19861);
nand UO_630 (O_630,N_19962,N_19924);
nor UO_631 (O_631,N_19985,N_19933);
or UO_632 (O_632,N_19888,N_19970);
and UO_633 (O_633,N_19988,N_19981);
xnor UO_634 (O_634,N_19887,N_19944);
and UO_635 (O_635,N_19980,N_19926);
nor UO_636 (O_636,N_19860,N_19904);
nor UO_637 (O_637,N_19905,N_19979);
and UO_638 (O_638,N_19870,N_19919);
xnor UO_639 (O_639,N_19967,N_19957);
nor UO_640 (O_640,N_19904,N_19990);
or UO_641 (O_641,N_19946,N_19913);
xor UO_642 (O_642,N_19987,N_19879);
or UO_643 (O_643,N_19900,N_19974);
and UO_644 (O_644,N_19945,N_19861);
or UO_645 (O_645,N_19993,N_19907);
nand UO_646 (O_646,N_19880,N_19978);
or UO_647 (O_647,N_19842,N_19953);
nor UO_648 (O_648,N_19964,N_19915);
and UO_649 (O_649,N_19915,N_19883);
nor UO_650 (O_650,N_19883,N_19897);
nor UO_651 (O_651,N_19938,N_19969);
xnor UO_652 (O_652,N_19889,N_19978);
xnor UO_653 (O_653,N_19881,N_19940);
xor UO_654 (O_654,N_19968,N_19920);
or UO_655 (O_655,N_19993,N_19931);
xor UO_656 (O_656,N_19864,N_19968);
nor UO_657 (O_657,N_19894,N_19951);
nand UO_658 (O_658,N_19844,N_19854);
nand UO_659 (O_659,N_19989,N_19998);
and UO_660 (O_660,N_19910,N_19994);
and UO_661 (O_661,N_19916,N_19970);
nor UO_662 (O_662,N_19864,N_19981);
and UO_663 (O_663,N_19846,N_19880);
nor UO_664 (O_664,N_19905,N_19983);
xnor UO_665 (O_665,N_19898,N_19983);
nor UO_666 (O_666,N_19890,N_19991);
or UO_667 (O_667,N_19925,N_19893);
nor UO_668 (O_668,N_19932,N_19993);
or UO_669 (O_669,N_19951,N_19950);
or UO_670 (O_670,N_19924,N_19898);
and UO_671 (O_671,N_19881,N_19961);
and UO_672 (O_672,N_19902,N_19895);
xor UO_673 (O_673,N_19892,N_19942);
or UO_674 (O_674,N_19946,N_19903);
nand UO_675 (O_675,N_19947,N_19983);
nor UO_676 (O_676,N_19933,N_19983);
or UO_677 (O_677,N_19844,N_19961);
xnor UO_678 (O_678,N_19944,N_19860);
or UO_679 (O_679,N_19866,N_19968);
xnor UO_680 (O_680,N_19944,N_19989);
nor UO_681 (O_681,N_19995,N_19911);
nand UO_682 (O_682,N_19930,N_19920);
xnor UO_683 (O_683,N_19951,N_19968);
and UO_684 (O_684,N_19901,N_19941);
nor UO_685 (O_685,N_19895,N_19865);
or UO_686 (O_686,N_19954,N_19900);
or UO_687 (O_687,N_19905,N_19914);
and UO_688 (O_688,N_19883,N_19949);
or UO_689 (O_689,N_19987,N_19852);
or UO_690 (O_690,N_19929,N_19895);
or UO_691 (O_691,N_19908,N_19886);
or UO_692 (O_692,N_19853,N_19897);
nor UO_693 (O_693,N_19871,N_19857);
and UO_694 (O_694,N_19895,N_19961);
or UO_695 (O_695,N_19945,N_19852);
nand UO_696 (O_696,N_19934,N_19969);
and UO_697 (O_697,N_19841,N_19909);
and UO_698 (O_698,N_19849,N_19959);
or UO_699 (O_699,N_19886,N_19956);
and UO_700 (O_700,N_19851,N_19947);
nand UO_701 (O_701,N_19975,N_19999);
nor UO_702 (O_702,N_19848,N_19967);
or UO_703 (O_703,N_19987,N_19950);
nor UO_704 (O_704,N_19997,N_19929);
and UO_705 (O_705,N_19973,N_19911);
xor UO_706 (O_706,N_19980,N_19857);
xor UO_707 (O_707,N_19878,N_19959);
nor UO_708 (O_708,N_19846,N_19926);
and UO_709 (O_709,N_19876,N_19904);
and UO_710 (O_710,N_19982,N_19840);
xor UO_711 (O_711,N_19895,N_19912);
nand UO_712 (O_712,N_19926,N_19864);
nand UO_713 (O_713,N_19840,N_19981);
and UO_714 (O_714,N_19995,N_19938);
and UO_715 (O_715,N_19842,N_19935);
nand UO_716 (O_716,N_19862,N_19992);
or UO_717 (O_717,N_19924,N_19936);
xnor UO_718 (O_718,N_19891,N_19918);
nand UO_719 (O_719,N_19963,N_19942);
nand UO_720 (O_720,N_19902,N_19871);
nor UO_721 (O_721,N_19986,N_19976);
nor UO_722 (O_722,N_19904,N_19910);
nand UO_723 (O_723,N_19991,N_19848);
nor UO_724 (O_724,N_19856,N_19860);
nor UO_725 (O_725,N_19874,N_19985);
and UO_726 (O_726,N_19928,N_19951);
or UO_727 (O_727,N_19910,N_19898);
nor UO_728 (O_728,N_19850,N_19875);
xor UO_729 (O_729,N_19894,N_19905);
or UO_730 (O_730,N_19842,N_19927);
xor UO_731 (O_731,N_19946,N_19989);
xor UO_732 (O_732,N_19986,N_19854);
xor UO_733 (O_733,N_19943,N_19858);
or UO_734 (O_734,N_19960,N_19947);
nand UO_735 (O_735,N_19852,N_19909);
or UO_736 (O_736,N_19909,N_19922);
xnor UO_737 (O_737,N_19847,N_19897);
nor UO_738 (O_738,N_19853,N_19859);
or UO_739 (O_739,N_19850,N_19960);
or UO_740 (O_740,N_19902,N_19951);
or UO_741 (O_741,N_19987,N_19958);
or UO_742 (O_742,N_19859,N_19883);
xor UO_743 (O_743,N_19926,N_19885);
nand UO_744 (O_744,N_19972,N_19958);
and UO_745 (O_745,N_19937,N_19906);
and UO_746 (O_746,N_19870,N_19862);
or UO_747 (O_747,N_19880,N_19975);
and UO_748 (O_748,N_19982,N_19857);
or UO_749 (O_749,N_19949,N_19952);
or UO_750 (O_750,N_19879,N_19846);
nand UO_751 (O_751,N_19972,N_19844);
or UO_752 (O_752,N_19968,N_19991);
nor UO_753 (O_753,N_19903,N_19895);
and UO_754 (O_754,N_19995,N_19952);
and UO_755 (O_755,N_19990,N_19949);
nor UO_756 (O_756,N_19871,N_19893);
or UO_757 (O_757,N_19906,N_19870);
or UO_758 (O_758,N_19910,N_19905);
and UO_759 (O_759,N_19935,N_19976);
or UO_760 (O_760,N_19944,N_19923);
or UO_761 (O_761,N_19906,N_19878);
xnor UO_762 (O_762,N_19981,N_19868);
and UO_763 (O_763,N_19917,N_19993);
nor UO_764 (O_764,N_19926,N_19843);
nor UO_765 (O_765,N_19973,N_19888);
and UO_766 (O_766,N_19846,N_19852);
or UO_767 (O_767,N_19887,N_19896);
nand UO_768 (O_768,N_19977,N_19849);
or UO_769 (O_769,N_19981,N_19934);
nor UO_770 (O_770,N_19991,N_19875);
nand UO_771 (O_771,N_19973,N_19975);
nand UO_772 (O_772,N_19872,N_19937);
xor UO_773 (O_773,N_19974,N_19992);
nor UO_774 (O_774,N_19880,N_19843);
or UO_775 (O_775,N_19885,N_19868);
and UO_776 (O_776,N_19982,N_19916);
and UO_777 (O_777,N_19919,N_19859);
or UO_778 (O_778,N_19979,N_19896);
xor UO_779 (O_779,N_19971,N_19845);
or UO_780 (O_780,N_19979,N_19902);
or UO_781 (O_781,N_19918,N_19852);
xnor UO_782 (O_782,N_19917,N_19944);
or UO_783 (O_783,N_19931,N_19987);
nand UO_784 (O_784,N_19916,N_19957);
or UO_785 (O_785,N_19903,N_19883);
xor UO_786 (O_786,N_19863,N_19927);
nand UO_787 (O_787,N_19894,N_19920);
nand UO_788 (O_788,N_19964,N_19999);
nand UO_789 (O_789,N_19920,N_19847);
nand UO_790 (O_790,N_19921,N_19966);
or UO_791 (O_791,N_19871,N_19894);
nor UO_792 (O_792,N_19862,N_19846);
nand UO_793 (O_793,N_19847,N_19989);
or UO_794 (O_794,N_19960,N_19996);
nor UO_795 (O_795,N_19949,N_19965);
or UO_796 (O_796,N_19857,N_19976);
nand UO_797 (O_797,N_19922,N_19989);
xnor UO_798 (O_798,N_19871,N_19927);
nand UO_799 (O_799,N_19951,N_19994);
xor UO_800 (O_800,N_19922,N_19995);
or UO_801 (O_801,N_19843,N_19964);
and UO_802 (O_802,N_19939,N_19994);
xnor UO_803 (O_803,N_19858,N_19862);
nand UO_804 (O_804,N_19991,N_19940);
and UO_805 (O_805,N_19867,N_19946);
or UO_806 (O_806,N_19898,N_19962);
and UO_807 (O_807,N_19970,N_19913);
and UO_808 (O_808,N_19841,N_19894);
and UO_809 (O_809,N_19956,N_19881);
xor UO_810 (O_810,N_19880,N_19903);
or UO_811 (O_811,N_19966,N_19979);
or UO_812 (O_812,N_19885,N_19895);
nand UO_813 (O_813,N_19986,N_19999);
and UO_814 (O_814,N_19979,N_19943);
xor UO_815 (O_815,N_19875,N_19926);
nand UO_816 (O_816,N_19890,N_19949);
and UO_817 (O_817,N_19990,N_19928);
nor UO_818 (O_818,N_19886,N_19965);
xor UO_819 (O_819,N_19855,N_19980);
nand UO_820 (O_820,N_19880,N_19937);
xor UO_821 (O_821,N_19862,N_19965);
xor UO_822 (O_822,N_19966,N_19951);
nand UO_823 (O_823,N_19843,N_19887);
xor UO_824 (O_824,N_19917,N_19954);
and UO_825 (O_825,N_19979,N_19951);
nand UO_826 (O_826,N_19988,N_19952);
xnor UO_827 (O_827,N_19932,N_19985);
nand UO_828 (O_828,N_19981,N_19841);
xor UO_829 (O_829,N_19843,N_19939);
nor UO_830 (O_830,N_19990,N_19963);
and UO_831 (O_831,N_19978,N_19974);
or UO_832 (O_832,N_19900,N_19864);
nor UO_833 (O_833,N_19951,N_19907);
and UO_834 (O_834,N_19934,N_19931);
nand UO_835 (O_835,N_19908,N_19977);
nor UO_836 (O_836,N_19989,N_19963);
nand UO_837 (O_837,N_19860,N_19912);
or UO_838 (O_838,N_19925,N_19989);
and UO_839 (O_839,N_19900,N_19938);
and UO_840 (O_840,N_19896,N_19915);
or UO_841 (O_841,N_19983,N_19943);
xor UO_842 (O_842,N_19921,N_19844);
nor UO_843 (O_843,N_19861,N_19889);
xnor UO_844 (O_844,N_19894,N_19910);
or UO_845 (O_845,N_19976,N_19871);
nor UO_846 (O_846,N_19998,N_19866);
nor UO_847 (O_847,N_19860,N_19992);
xnor UO_848 (O_848,N_19930,N_19935);
or UO_849 (O_849,N_19882,N_19887);
and UO_850 (O_850,N_19962,N_19882);
and UO_851 (O_851,N_19892,N_19872);
nor UO_852 (O_852,N_19850,N_19921);
nor UO_853 (O_853,N_19879,N_19903);
and UO_854 (O_854,N_19888,N_19986);
nor UO_855 (O_855,N_19847,N_19984);
or UO_856 (O_856,N_19998,N_19888);
and UO_857 (O_857,N_19969,N_19983);
xnor UO_858 (O_858,N_19846,N_19936);
nor UO_859 (O_859,N_19988,N_19996);
and UO_860 (O_860,N_19942,N_19895);
or UO_861 (O_861,N_19955,N_19970);
nor UO_862 (O_862,N_19925,N_19933);
or UO_863 (O_863,N_19969,N_19940);
or UO_864 (O_864,N_19949,N_19959);
or UO_865 (O_865,N_19849,N_19983);
or UO_866 (O_866,N_19940,N_19954);
nor UO_867 (O_867,N_19957,N_19996);
or UO_868 (O_868,N_19988,N_19929);
nand UO_869 (O_869,N_19977,N_19949);
xor UO_870 (O_870,N_19869,N_19983);
or UO_871 (O_871,N_19970,N_19926);
xnor UO_872 (O_872,N_19939,N_19860);
nor UO_873 (O_873,N_19913,N_19952);
nand UO_874 (O_874,N_19867,N_19967);
and UO_875 (O_875,N_19898,N_19902);
or UO_876 (O_876,N_19920,N_19910);
nand UO_877 (O_877,N_19921,N_19934);
and UO_878 (O_878,N_19928,N_19931);
nor UO_879 (O_879,N_19968,N_19999);
or UO_880 (O_880,N_19972,N_19892);
or UO_881 (O_881,N_19872,N_19942);
and UO_882 (O_882,N_19923,N_19965);
xnor UO_883 (O_883,N_19869,N_19885);
and UO_884 (O_884,N_19908,N_19972);
nand UO_885 (O_885,N_19853,N_19910);
nand UO_886 (O_886,N_19975,N_19907);
xor UO_887 (O_887,N_19975,N_19985);
or UO_888 (O_888,N_19851,N_19955);
nor UO_889 (O_889,N_19998,N_19875);
nor UO_890 (O_890,N_19953,N_19869);
nand UO_891 (O_891,N_19882,N_19900);
nor UO_892 (O_892,N_19984,N_19959);
and UO_893 (O_893,N_19910,N_19996);
nand UO_894 (O_894,N_19961,N_19902);
and UO_895 (O_895,N_19918,N_19872);
nor UO_896 (O_896,N_19843,N_19978);
and UO_897 (O_897,N_19987,N_19984);
and UO_898 (O_898,N_19955,N_19936);
or UO_899 (O_899,N_19993,N_19965);
xor UO_900 (O_900,N_19994,N_19944);
xor UO_901 (O_901,N_19975,N_19860);
or UO_902 (O_902,N_19910,N_19930);
nor UO_903 (O_903,N_19882,N_19883);
nor UO_904 (O_904,N_19884,N_19897);
and UO_905 (O_905,N_19853,N_19898);
xor UO_906 (O_906,N_19952,N_19869);
or UO_907 (O_907,N_19979,N_19948);
or UO_908 (O_908,N_19843,N_19924);
and UO_909 (O_909,N_19912,N_19857);
nor UO_910 (O_910,N_19988,N_19896);
nor UO_911 (O_911,N_19872,N_19936);
xor UO_912 (O_912,N_19881,N_19967);
nor UO_913 (O_913,N_19949,N_19926);
nor UO_914 (O_914,N_19962,N_19885);
and UO_915 (O_915,N_19846,N_19843);
or UO_916 (O_916,N_19894,N_19986);
nand UO_917 (O_917,N_19938,N_19847);
nor UO_918 (O_918,N_19890,N_19992);
or UO_919 (O_919,N_19959,N_19912);
or UO_920 (O_920,N_19942,N_19940);
and UO_921 (O_921,N_19995,N_19910);
or UO_922 (O_922,N_19880,N_19990);
nor UO_923 (O_923,N_19881,N_19992);
or UO_924 (O_924,N_19907,N_19885);
or UO_925 (O_925,N_19913,N_19915);
and UO_926 (O_926,N_19932,N_19850);
and UO_927 (O_927,N_19851,N_19869);
xor UO_928 (O_928,N_19897,N_19912);
nand UO_929 (O_929,N_19885,N_19912);
and UO_930 (O_930,N_19869,N_19970);
xnor UO_931 (O_931,N_19949,N_19874);
xor UO_932 (O_932,N_19998,N_19956);
or UO_933 (O_933,N_19994,N_19930);
xnor UO_934 (O_934,N_19949,N_19921);
xor UO_935 (O_935,N_19889,N_19908);
and UO_936 (O_936,N_19956,N_19979);
nand UO_937 (O_937,N_19874,N_19978);
xnor UO_938 (O_938,N_19944,N_19879);
nand UO_939 (O_939,N_19990,N_19889);
nor UO_940 (O_940,N_19851,N_19935);
xor UO_941 (O_941,N_19989,N_19914);
nor UO_942 (O_942,N_19973,N_19845);
nor UO_943 (O_943,N_19981,N_19962);
xnor UO_944 (O_944,N_19949,N_19932);
nand UO_945 (O_945,N_19922,N_19994);
nand UO_946 (O_946,N_19944,N_19962);
nand UO_947 (O_947,N_19870,N_19916);
nand UO_948 (O_948,N_19922,N_19993);
nor UO_949 (O_949,N_19988,N_19862);
nor UO_950 (O_950,N_19868,N_19989);
nor UO_951 (O_951,N_19860,N_19926);
or UO_952 (O_952,N_19986,N_19849);
nor UO_953 (O_953,N_19861,N_19995);
nor UO_954 (O_954,N_19880,N_19943);
and UO_955 (O_955,N_19843,N_19905);
xor UO_956 (O_956,N_19966,N_19887);
nand UO_957 (O_957,N_19840,N_19897);
or UO_958 (O_958,N_19946,N_19874);
xnor UO_959 (O_959,N_19958,N_19954);
xor UO_960 (O_960,N_19939,N_19903);
nand UO_961 (O_961,N_19914,N_19862);
xor UO_962 (O_962,N_19997,N_19941);
nand UO_963 (O_963,N_19860,N_19882);
and UO_964 (O_964,N_19957,N_19938);
nand UO_965 (O_965,N_19882,N_19964);
or UO_966 (O_966,N_19858,N_19894);
nand UO_967 (O_967,N_19850,N_19889);
or UO_968 (O_968,N_19964,N_19922);
or UO_969 (O_969,N_19952,N_19879);
xor UO_970 (O_970,N_19908,N_19933);
xnor UO_971 (O_971,N_19916,N_19861);
xor UO_972 (O_972,N_19885,N_19842);
nand UO_973 (O_973,N_19903,N_19956);
xor UO_974 (O_974,N_19969,N_19895);
and UO_975 (O_975,N_19958,N_19863);
xnor UO_976 (O_976,N_19965,N_19879);
and UO_977 (O_977,N_19906,N_19953);
nand UO_978 (O_978,N_19981,N_19963);
nand UO_979 (O_979,N_19945,N_19954);
and UO_980 (O_980,N_19967,N_19875);
xnor UO_981 (O_981,N_19904,N_19902);
xor UO_982 (O_982,N_19840,N_19979);
nor UO_983 (O_983,N_19916,N_19867);
or UO_984 (O_984,N_19865,N_19868);
nor UO_985 (O_985,N_19942,N_19868);
and UO_986 (O_986,N_19989,N_19918);
or UO_987 (O_987,N_19948,N_19962);
nand UO_988 (O_988,N_19853,N_19949);
xnor UO_989 (O_989,N_19967,N_19853);
nor UO_990 (O_990,N_19890,N_19868);
nor UO_991 (O_991,N_19867,N_19963);
and UO_992 (O_992,N_19921,N_19930);
nand UO_993 (O_993,N_19921,N_19914);
nand UO_994 (O_994,N_19853,N_19960);
or UO_995 (O_995,N_19948,N_19865);
or UO_996 (O_996,N_19909,N_19952);
xnor UO_997 (O_997,N_19936,N_19880);
xnor UO_998 (O_998,N_19904,N_19891);
and UO_999 (O_999,N_19954,N_19919);
nand UO_1000 (O_1000,N_19953,N_19888);
nor UO_1001 (O_1001,N_19901,N_19980);
and UO_1002 (O_1002,N_19841,N_19914);
xor UO_1003 (O_1003,N_19942,N_19902);
and UO_1004 (O_1004,N_19914,N_19840);
and UO_1005 (O_1005,N_19901,N_19861);
nand UO_1006 (O_1006,N_19906,N_19952);
and UO_1007 (O_1007,N_19865,N_19940);
xor UO_1008 (O_1008,N_19858,N_19927);
nor UO_1009 (O_1009,N_19880,N_19994);
and UO_1010 (O_1010,N_19999,N_19956);
nor UO_1011 (O_1011,N_19968,N_19998);
or UO_1012 (O_1012,N_19893,N_19882);
or UO_1013 (O_1013,N_19898,N_19867);
xor UO_1014 (O_1014,N_19849,N_19908);
and UO_1015 (O_1015,N_19939,N_19985);
and UO_1016 (O_1016,N_19856,N_19964);
nand UO_1017 (O_1017,N_19988,N_19969);
nand UO_1018 (O_1018,N_19899,N_19893);
xnor UO_1019 (O_1019,N_19943,N_19956);
nand UO_1020 (O_1020,N_19932,N_19984);
and UO_1021 (O_1021,N_19862,N_19929);
nand UO_1022 (O_1022,N_19864,N_19909);
or UO_1023 (O_1023,N_19881,N_19954);
and UO_1024 (O_1024,N_19993,N_19897);
and UO_1025 (O_1025,N_19944,N_19861);
xor UO_1026 (O_1026,N_19923,N_19881);
and UO_1027 (O_1027,N_19866,N_19895);
or UO_1028 (O_1028,N_19846,N_19973);
and UO_1029 (O_1029,N_19912,N_19963);
nand UO_1030 (O_1030,N_19995,N_19919);
nor UO_1031 (O_1031,N_19970,N_19992);
or UO_1032 (O_1032,N_19843,N_19870);
nor UO_1033 (O_1033,N_19849,N_19858);
nor UO_1034 (O_1034,N_19953,N_19997);
or UO_1035 (O_1035,N_19960,N_19932);
xnor UO_1036 (O_1036,N_19854,N_19916);
nor UO_1037 (O_1037,N_19979,N_19936);
xnor UO_1038 (O_1038,N_19984,N_19975);
nand UO_1039 (O_1039,N_19929,N_19885);
nor UO_1040 (O_1040,N_19861,N_19911);
nor UO_1041 (O_1041,N_19927,N_19992);
or UO_1042 (O_1042,N_19910,N_19907);
nand UO_1043 (O_1043,N_19846,N_19855);
nand UO_1044 (O_1044,N_19979,N_19842);
nor UO_1045 (O_1045,N_19906,N_19877);
and UO_1046 (O_1046,N_19994,N_19984);
or UO_1047 (O_1047,N_19884,N_19937);
and UO_1048 (O_1048,N_19875,N_19904);
nand UO_1049 (O_1049,N_19949,N_19987);
xor UO_1050 (O_1050,N_19888,N_19989);
or UO_1051 (O_1051,N_19892,N_19949);
xor UO_1052 (O_1052,N_19942,N_19887);
xor UO_1053 (O_1053,N_19874,N_19973);
and UO_1054 (O_1054,N_19992,N_19876);
nand UO_1055 (O_1055,N_19950,N_19948);
xnor UO_1056 (O_1056,N_19989,N_19991);
nand UO_1057 (O_1057,N_19916,N_19881);
and UO_1058 (O_1058,N_19960,N_19974);
or UO_1059 (O_1059,N_19998,N_19906);
nand UO_1060 (O_1060,N_19978,N_19906);
nor UO_1061 (O_1061,N_19865,N_19957);
nor UO_1062 (O_1062,N_19877,N_19952);
nor UO_1063 (O_1063,N_19902,N_19883);
xnor UO_1064 (O_1064,N_19909,N_19878);
nand UO_1065 (O_1065,N_19957,N_19856);
and UO_1066 (O_1066,N_19846,N_19955);
nand UO_1067 (O_1067,N_19891,N_19868);
and UO_1068 (O_1068,N_19924,N_19864);
nand UO_1069 (O_1069,N_19981,N_19957);
nor UO_1070 (O_1070,N_19947,N_19954);
nor UO_1071 (O_1071,N_19847,N_19945);
nand UO_1072 (O_1072,N_19971,N_19891);
or UO_1073 (O_1073,N_19889,N_19902);
xnor UO_1074 (O_1074,N_19981,N_19961);
and UO_1075 (O_1075,N_19991,N_19970);
or UO_1076 (O_1076,N_19921,N_19882);
nand UO_1077 (O_1077,N_19860,N_19974);
nand UO_1078 (O_1078,N_19889,N_19933);
nand UO_1079 (O_1079,N_19874,N_19960);
nand UO_1080 (O_1080,N_19911,N_19883);
and UO_1081 (O_1081,N_19866,N_19977);
xor UO_1082 (O_1082,N_19844,N_19856);
or UO_1083 (O_1083,N_19881,N_19965);
or UO_1084 (O_1084,N_19853,N_19888);
nor UO_1085 (O_1085,N_19955,N_19998);
or UO_1086 (O_1086,N_19910,N_19864);
nand UO_1087 (O_1087,N_19956,N_19874);
and UO_1088 (O_1088,N_19882,N_19916);
xor UO_1089 (O_1089,N_19865,N_19851);
xnor UO_1090 (O_1090,N_19841,N_19858);
or UO_1091 (O_1091,N_19981,N_19902);
nor UO_1092 (O_1092,N_19996,N_19846);
nand UO_1093 (O_1093,N_19929,N_19943);
xor UO_1094 (O_1094,N_19914,N_19844);
nand UO_1095 (O_1095,N_19949,N_19964);
nor UO_1096 (O_1096,N_19961,N_19884);
xor UO_1097 (O_1097,N_19949,N_19966);
xor UO_1098 (O_1098,N_19925,N_19975);
nand UO_1099 (O_1099,N_19943,N_19904);
and UO_1100 (O_1100,N_19867,N_19948);
and UO_1101 (O_1101,N_19971,N_19914);
and UO_1102 (O_1102,N_19929,N_19978);
and UO_1103 (O_1103,N_19884,N_19932);
xor UO_1104 (O_1104,N_19909,N_19846);
nand UO_1105 (O_1105,N_19882,N_19985);
xnor UO_1106 (O_1106,N_19848,N_19954);
xor UO_1107 (O_1107,N_19933,N_19987);
nand UO_1108 (O_1108,N_19903,N_19911);
or UO_1109 (O_1109,N_19961,N_19939);
or UO_1110 (O_1110,N_19921,N_19857);
or UO_1111 (O_1111,N_19992,N_19967);
and UO_1112 (O_1112,N_19880,N_19841);
nor UO_1113 (O_1113,N_19991,N_19933);
nand UO_1114 (O_1114,N_19987,N_19979);
and UO_1115 (O_1115,N_19902,N_19873);
and UO_1116 (O_1116,N_19883,N_19945);
xnor UO_1117 (O_1117,N_19930,N_19973);
nor UO_1118 (O_1118,N_19936,N_19995);
or UO_1119 (O_1119,N_19971,N_19895);
or UO_1120 (O_1120,N_19965,N_19922);
or UO_1121 (O_1121,N_19986,N_19964);
nor UO_1122 (O_1122,N_19928,N_19964);
nor UO_1123 (O_1123,N_19940,N_19998);
and UO_1124 (O_1124,N_19997,N_19868);
or UO_1125 (O_1125,N_19854,N_19840);
nor UO_1126 (O_1126,N_19925,N_19999);
and UO_1127 (O_1127,N_19904,N_19883);
nand UO_1128 (O_1128,N_19875,N_19950);
or UO_1129 (O_1129,N_19842,N_19975);
nand UO_1130 (O_1130,N_19994,N_19911);
or UO_1131 (O_1131,N_19896,N_19955);
or UO_1132 (O_1132,N_19979,N_19973);
xnor UO_1133 (O_1133,N_19853,N_19871);
and UO_1134 (O_1134,N_19970,N_19896);
nand UO_1135 (O_1135,N_19872,N_19992);
nor UO_1136 (O_1136,N_19909,N_19920);
xnor UO_1137 (O_1137,N_19993,N_19895);
xnor UO_1138 (O_1138,N_19882,N_19946);
nor UO_1139 (O_1139,N_19969,N_19949);
and UO_1140 (O_1140,N_19880,N_19958);
xnor UO_1141 (O_1141,N_19911,N_19985);
nor UO_1142 (O_1142,N_19967,N_19903);
nor UO_1143 (O_1143,N_19844,N_19951);
or UO_1144 (O_1144,N_19906,N_19924);
nor UO_1145 (O_1145,N_19953,N_19976);
nand UO_1146 (O_1146,N_19938,N_19852);
nor UO_1147 (O_1147,N_19898,N_19952);
xor UO_1148 (O_1148,N_19853,N_19864);
or UO_1149 (O_1149,N_19850,N_19924);
nand UO_1150 (O_1150,N_19901,N_19950);
and UO_1151 (O_1151,N_19861,N_19877);
xnor UO_1152 (O_1152,N_19893,N_19932);
and UO_1153 (O_1153,N_19952,N_19917);
xnor UO_1154 (O_1154,N_19865,N_19964);
and UO_1155 (O_1155,N_19910,N_19888);
xnor UO_1156 (O_1156,N_19979,N_19997);
and UO_1157 (O_1157,N_19920,N_19967);
nand UO_1158 (O_1158,N_19939,N_19897);
or UO_1159 (O_1159,N_19922,N_19934);
or UO_1160 (O_1160,N_19873,N_19883);
and UO_1161 (O_1161,N_19941,N_19945);
or UO_1162 (O_1162,N_19945,N_19873);
and UO_1163 (O_1163,N_19918,N_19883);
nand UO_1164 (O_1164,N_19863,N_19923);
nor UO_1165 (O_1165,N_19938,N_19911);
xnor UO_1166 (O_1166,N_19990,N_19846);
and UO_1167 (O_1167,N_19959,N_19972);
or UO_1168 (O_1168,N_19935,N_19938);
or UO_1169 (O_1169,N_19966,N_19924);
and UO_1170 (O_1170,N_19846,N_19918);
xor UO_1171 (O_1171,N_19844,N_19999);
nor UO_1172 (O_1172,N_19988,N_19934);
and UO_1173 (O_1173,N_19996,N_19853);
and UO_1174 (O_1174,N_19980,N_19947);
and UO_1175 (O_1175,N_19845,N_19857);
nand UO_1176 (O_1176,N_19879,N_19986);
and UO_1177 (O_1177,N_19928,N_19917);
nor UO_1178 (O_1178,N_19990,N_19975);
and UO_1179 (O_1179,N_19955,N_19889);
and UO_1180 (O_1180,N_19957,N_19855);
nor UO_1181 (O_1181,N_19868,N_19878);
nand UO_1182 (O_1182,N_19842,N_19905);
and UO_1183 (O_1183,N_19913,N_19898);
nand UO_1184 (O_1184,N_19900,N_19960);
nand UO_1185 (O_1185,N_19974,N_19930);
nor UO_1186 (O_1186,N_19920,N_19956);
and UO_1187 (O_1187,N_19913,N_19875);
or UO_1188 (O_1188,N_19909,N_19941);
nor UO_1189 (O_1189,N_19960,N_19920);
and UO_1190 (O_1190,N_19897,N_19916);
and UO_1191 (O_1191,N_19969,N_19841);
nand UO_1192 (O_1192,N_19985,N_19920);
and UO_1193 (O_1193,N_19853,N_19978);
nor UO_1194 (O_1194,N_19854,N_19931);
nand UO_1195 (O_1195,N_19984,N_19969);
nor UO_1196 (O_1196,N_19894,N_19985);
xor UO_1197 (O_1197,N_19881,N_19935);
and UO_1198 (O_1198,N_19986,N_19873);
nor UO_1199 (O_1199,N_19934,N_19980);
nand UO_1200 (O_1200,N_19857,N_19904);
nand UO_1201 (O_1201,N_19977,N_19911);
and UO_1202 (O_1202,N_19841,N_19920);
and UO_1203 (O_1203,N_19998,N_19859);
nor UO_1204 (O_1204,N_19975,N_19872);
or UO_1205 (O_1205,N_19901,N_19859);
and UO_1206 (O_1206,N_19927,N_19841);
or UO_1207 (O_1207,N_19889,N_19996);
nand UO_1208 (O_1208,N_19868,N_19931);
and UO_1209 (O_1209,N_19978,N_19859);
and UO_1210 (O_1210,N_19967,N_19948);
xnor UO_1211 (O_1211,N_19988,N_19920);
nand UO_1212 (O_1212,N_19898,N_19987);
nor UO_1213 (O_1213,N_19928,N_19868);
or UO_1214 (O_1214,N_19860,N_19901);
nand UO_1215 (O_1215,N_19901,N_19967);
nand UO_1216 (O_1216,N_19981,N_19938);
xor UO_1217 (O_1217,N_19845,N_19890);
or UO_1218 (O_1218,N_19875,N_19918);
xor UO_1219 (O_1219,N_19904,N_19849);
and UO_1220 (O_1220,N_19922,N_19957);
and UO_1221 (O_1221,N_19948,N_19982);
nand UO_1222 (O_1222,N_19917,N_19874);
and UO_1223 (O_1223,N_19948,N_19859);
nor UO_1224 (O_1224,N_19873,N_19977);
nor UO_1225 (O_1225,N_19986,N_19882);
and UO_1226 (O_1226,N_19932,N_19988);
or UO_1227 (O_1227,N_19995,N_19893);
and UO_1228 (O_1228,N_19914,N_19928);
xor UO_1229 (O_1229,N_19979,N_19939);
nand UO_1230 (O_1230,N_19996,N_19870);
nand UO_1231 (O_1231,N_19967,N_19935);
nor UO_1232 (O_1232,N_19985,N_19855);
or UO_1233 (O_1233,N_19869,N_19994);
xnor UO_1234 (O_1234,N_19963,N_19944);
xor UO_1235 (O_1235,N_19908,N_19882);
xnor UO_1236 (O_1236,N_19920,N_19958);
nor UO_1237 (O_1237,N_19869,N_19998);
and UO_1238 (O_1238,N_19933,N_19954);
or UO_1239 (O_1239,N_19888,N_19994);
nand UO_1240 (O_1240,N_19971,N_19969);
and UO_1241 (O_1241,N_19885,N_19981);
nor UO_1242 (O_1242,N_19944,N_19872);
or UO_1243 (O_1243,N_19913,N_19944);
or UO_1244 (O_1244,N_19919,N_19933);
or UO_1245 (O_1245,N_19886,N_19923);
xnor UO_1246 (O_1246,N_19877,N_19853);
nand UO_1247 (O_1247,N_19881,N_19974);
xnor UO_1248 (O_1248,N_19920,N_19888);
and UO_1249 (O_1249,N_19853,N_19903);
xnor UO_1250 (O_1250,N_19976,N_19886);
or UO_1251 (O_1251,N_19973,N_19887);
xnor UO_1252 (O_1252,N_19925,N_19914);
or UO_1253 (O_1253,N_19985,N_19916);
nand UO_1254 (O_1254,N_19881,N_19945);
xnor UO_1255 (O_1255,N_19850,N_19988);
nor UO_1256 (O_1256,N_19934,N_19889);
xor UO_1257 (O_1257,N_19857,N_19967);
nand UO_1258 (O_1258,N_19842,N_19930);
or UO_1259 (O_1259,N_19855,N_19872);
or UO_1260 (O_1260,N_19865,N_19944);
nor UO_1261 (O_1261,N_19937,N_19954);
or UO_1262 (O_1262,N_19924,N_19950);
or UO_1263 (O_1263,N_19963,N_19995);
and UO_1264 (O_1264,N_19842,N_19908);
nand UO_1265 (O_1265,N_19969,N_19869);
or UO_1266 (O_1266,N_19860,N_19999);
nand UO_1267 (O_1267,N_19872,N_19845);
or UO_1268 (O_1268,N_19980,N_19886);
xnor UO_1269 (O_1269,N_19895,N_19881);
nor UO_1270 (O_1270,N_19892,N_19987);
nor UO_1271 (O_1271,N_19975,N_19942);
xnor UO_1272 (O_1272,N_19865,N_19969);
xor UO_1273 (O_1273,N_19860,N_19986);
and UO_1274 (O_1274,N_19997,N_19844);
nand UO_1275 (O_1275,N_19872,N_19933);
nor UO_1276 (O_1276,N_19852,N_19901);
and UO_1277 (O_1277,N_19950,N_19960);
or UO_1278 (O_1278,N_19891,N_19906);
xor UO_1279 (O_1279,N_19972,N_19898);
nor UO_1280 (O_1280,N_19938,N_19961);
nand UO_1281 (O_1281,N_19841,N_19874);
nand UO_1282 (O_1282,N_19971,N_19929);
nor UO_1283 (O_1283,N_19869,N_19980);
xor UO_1284 (O_1284,N_19859,N_19943);
nor UO_1285 (O_1285,N_19932,N_19969);
and UO_1286 (O_1286,N_19998,N_19901);
or UO_1287 (O_1287,N_19922,N_19985);
xnor UO_1288 (O_1288,N_19913,N_19919);
xnor UO_1289 (O_1289,N_19959,N_19986);
and UO_1290 (O_1290,N_19944,N_19945);
xor UO_1291 (O_1291,N_19846,N_19841);
or UO_1292 (O_1292,N_19884,N_19895);
nand UO_1293 (O_1293,N_19982,N_19988);
xnor UO_1294 (O_1294,N_19911,N_19989);
xor UO_1295 (O_1295,N_19895,N_19958);
nand UO_1296 (O_1296,N_19855,N_19885);
xor UO_1297 (O_1297,N_19842,N_19918);
or UO_1298 (O_1298,N_19928,N_19944);
or UO_1299 (O_1299,N_19854,N_19940);
xor UO_1300 (O_1300,N_19997,N_19912);
or UO_1301 (O_1301,N_19970,N_19968);
or UO_1302 (O_1302,N_19858,N_19995);
and UO_1303 (O_1303,N_19969,N_19998);
xnor UO_1304 (O_1304,N_19843,N_19970);
xnor UO_1305 (O_1305,N_19891,N_19905);
nand UO_1306 (O_1306,N_19891,N_19992);
or UO_1307 (O_1307,N_19975,N_19951);
and UO_1308 (O_1308,N_19982,N_19935);
or UO_1309 (O_1309,N_19906,N_19930);
nand UO_1310 (O_1310,N_19917,N_19976);
or UO_1311 (O_1311,N_19934,N_19885);
or UO_1312 (O_1312,N_19941,N_19878);
and UO_1313 (O_1313,N_19914,N_19952);
nand UO_1314 (O_1314,N_19977,N_19967);
xor UO_1315 (O_1315,N_19936,N_19943);
nor UO_1316 (O_1316,N_19856,N_19977);
xor UO_1317 (O_1317,N_19878,N_19843);
and UO_1318 (O_1318,N_19990,N_19917);
xnor UO_1319 (O_1319,N_19910,N_19901);
and UO_1320 (O_1320,N_19966,N_19873);
nand UO_1321 (O_1321,N_19925,N_19840);
xor UO_1322 (O_1322,N_19849,N_19970);
or UO_1323 (O_1323,N_19905,N_19968);
xor UO_1324 (O_1324,N_19986,N_19842);
nor UO_1325 (O_1325,N_19870,N_19932);
or UO_1326 (O_1326,N_19907,N_19871);
xnor UO_1327 (O_1327,N_19921,N_19932);
and UO_1328 (O_1328,N_19885,N_19945);
xor UO_1329 (O_1329,N_19996,N_19981);
nand UO_1330 (O_1330,N_19995,N_19873);
nand UO_1331 (O_1331,N_19936,N_19897);
and UO_1332 (O_1332,N_19872,N_19977);
or UO_1333 (O_1333,N_19963,N_19960);
xor UO_1334 (O_1334,N_19905,N_19943);
and UO_1335 (O_1335,N_19914,N_19986);
nor UO_1336 (O_1336,N_19997,N_19966);
and UO_1337 (O_1337,N_19940,N_19907);
xnor UO_1338 (O_1338,N_19958,N_19963);
and UO_1339 (O_1339,N_19884,N_19890);
and UO_1340 (O_1340,N_19991,N_19905);
nand UO_1341 (O_1341,N_19940,N_19971);
nand UO_1342 (O_1342,N_19911,N_19972);
xnor UO_1343 (O_1343,N_19952,N_19958);
nand UO_1344 (O_1344,N_19842,N_19911);
nand UO_1345 (O_1345,N_19840,N_19845);
xnor UO_1346 (O_1346,N_19887,N_19884);
nand UO_1347 (O_1347,N_19858,N_19987);
and UO_1348 (O_1348,N_19855,N_19930);
nand UO_1349 (O_1349,N_19890,N_19866);
nand UO_1350 (O_1350,N_19925,N_19948);
nor UO_1351 (O_1351,N_19893,N_19918);
xor UO_1352 (O_1352,N_19966,N_19927);
nand UO_1353 (O_1353,N_19898,N_19840);
or UO_1354 (O_1354,N_19894,N_19957);
or UO_1355 (O_1355,N_19947,N_19989);
xor UO_1356 (O_1356,N_19874,N_19919);
or UO_1357 (O_1357,N_19851,N_19953);
nor UO_1358 (O_1358,N_19940,N_19856);
xnor UO_1359 (O_1359,N_19933,N_19861);
or UO_1360 (O_1360,N_19975,N_19970);
xnor UO_1361 (O_1361,N_19895,N_19975);
or UO_1362 (O_1362,N_19949,N_19904);
or UO_1363 (O_1363,N_19995,N_19914);
xnor UO_1364 (O_1364,N_19915,N_19873);
or UO_1365 (O_1365,N_19973,N_19994);
or UO_1366 (O_1366,N_19883,N_19956);
and UO_1367 (O_1367,N_19857,N_19924);
and UO_1368 (O_1368,N_19883,N_19963);
nand UO_1369 (O_1369,N_19866,N_19843);
nor UO_1370 (O_1370,N_19847,N_19928);
nor UO_1371 (O_1371,N_19959,N_19945);
or UO_1372 (O_1372,N_19997,N_19923);
nand UO_1373 (O_1373,N_19939,N_19908);
xor UO_1374 (O_1374,N_19923,N_19893);
xor UO_1375 (O_1375,N_19991,N_19988);
nor UO_1376 (O_1376,N_19881,N_19997);
and UO_1377 (O_1377,N_19917,N_19940);
or UO_1378 (O_1378,N_19923,N_19856);
nand UO_1379 (O_1379,N_19934,N_19999);
xor UO_1380 (O_1380,N_19927,N_19962);
or UO_1381 (O_1381,N_19875,N_19977);
nand UO_1382 (O_1382,N_19864,N_19984);
or UO_1383 (O_1383,N_19936,N_19843);
or UO_1384 (O_1384,N_19940,N_19884);
nand UO_1385 (O_1385,N_19854,N_19936);
nor UO_1386 (O_1386,N_19873,N_19875);
xnor UO_1387 (O_1387,N_19913,N_19873);
and UO_1388 (O_1388,N_19965,N_19858);
xor UO_1389 (O_1389,N_19948,N_19871);
nor UO_1390 (O_1390,N_19964,N_19897);
nand UO_1391 (O_1391,N_19960,N_19907);
or UO_1392 (O_1392,N_19860,N_19876);
nand UO_1393 (O_1393,N_19929,N_19991);
nand UO_1394 (O_1394,N_19975,N_19993);
xor UO_1395 (O_1395,N_19911,N_19859);
nand UO_1396 (O_1396,N_19938,N_19895);
or UO_1397 (O_1397,N_19981,N_19873);
nor UO_1398 (O_1398,N_19845,N_19874);
xnor UO_1399 (O_1399,N_19918,N_19851);
nand UO_1400 (O_1400,N_19915,N_19909);
nand UO_1401 (O_1401,N_19900,N_19968);
and UO_1402 (O_1402,N_19918,N_19890);
or UO_1403 (O_1403,N_19962,N_19847);
or UO_1404 (O_1404,N_19986,N_19954);
xor UO_1405 (O_1405,N_19931,N_19974);
nor UO_1406 (O_1406,N_19937,N_19997);
nor UO_1407 (O_1407,N_19933,N_19965);
nor UO_1408 (O_1408,N_19882,N_19841);
and UO_1409 (O_1409,N_19968,N_19859);
and UO_1410 (O_1410,N_19842,N_19963);
or UO_1411 (O_1411,N_19845,N_19979);
or UO_1412 (O_1412,N_19892,N_19985);
xor UO_1413 (O_1413,N_19908,N_19868);
and UO_1414 (O_1414,N_19857,N_19910);
nor UO_1415 (O_1415,N_19905,N_19872);
or UO_1416 (O_1416,N_19953,N_19966);
nand UO_1417 (O_1417,N_19852,N_19890);
nor UO_1418 (O_1418,N_19987,N_19848);
xnor UO_1419 (O_1419,N_19933,N_19911);
or UO_1420 (O_1420,N_19949,N_19847);
and UO_1421 (O_1421,N_19943,N_19963);
xor UO_1422 (O_1422,N_19887,N_19864);
nor UO_1423 (O_1423,N_19869,N_19988);
xor UO_1424 (O_1424,N_19997,N_19952);
and UO_1425 (O_1425,N_19876,N_19994);
or UO_1426 (O_1426,N_19896,N_19843);
nor UO_1427 (O_1427,N_19895,N_19983);
and UO_1428 (O_1428,N_19948,N_19965);
nor UO_1429 (O_1429,N_19960,N_19876);
or UO_1430 (O_1430,N_19959,N_19856);
or UO_1431 (O_1431,N_19849,N_19864);
and UO_1432 (O_1432,N_19860,N_19977);
or UO_1433 (O_1433,N_19906,N_19951);
xor UO_1434 (O_1434,N_19999,N_19913);
nor UO_1435 (O_1435,N_19934,N_19854);
and UO_1436 (O_1436,N_19964,N_19982);
or UO_1437 (O_1437,N_19851,N_19877);
nand UO_1438 (O_1438,N_19901,N_19944);
or UO_1439 (O_1439,N_19904,N_19963);
xnor UO_1440 (O_1440,N_19851,N_19854);
and UO_1441 (O_1441,N_19878,N_19851);
and UO_1442 (O_1442,N_19976,N_19969);
nor UO_1443 (O_1443,N_19867,N_19955);
nand UO_1444 (O_1444,N_19912,N_19979);
xnor UO_1445 (O_1445,N_19949,N_19946);
nand UO_1446 (O_1446,N_19902,N_19899);
or UO_1447 (O_1447,N_19915,N_19931);
nor UO_1448 (O_1448,N_19852,N_19841);
nor UO_1449 (O_1449,N_19841,N_19932);
nand UO_1450 (O_1450,N_19903,N_19986);
nand UO_1451 (O_1451,N_19986,N_19919);
or UO_1452 (O_1452,N_19925,N_19941);
xnor UO_1453 (O_1453,N_19879,N_19920);
nand UO_1454 (O_1454,N_19935,N_19995);
or UO_1455 (O_1455,N_19976,N_19987);
or UO_1456 (O_1456,N_19922,N_19869);
and UO_1457 (O_1457,N_19928,N_19950);
and UO_1458 (O_1458,N_19996,N_19899);
and UO_1459 (O_1459,N_19848,N_19980);
nand UO_1460 (O_1460,N_19909,N_19905);
xnor UO_1461 (O_1461,N_19971,N_19945);
xnor UO_1462 (O_1462,N_19869,N_19987);
nand UO_1463 (O_1463,N_19916,N_19887);
and UO_1464 (O_1464,N_19958,N_19847);
xnor UO_1465 (O_1465,N_19953,N_19992);
nand UO_1466 (O_1466,N_19858,N_19945);
nor UO_1467 (O_1467,N_19979,N_19957);
or UO_1468 (O_1468,N_19930,N_19942);
nand UO_1469 (O_1469,N_19986,N_19863);
nor UO_1470 (O_1470,N_19984,N_19858);
or UO_1471 (O_1471,N_19967,N_19997);
nor UO_1472 (O_1472,N_19909,N_19876);
or UO_1473 (O_1473,N_19866,N_19947);
nand UO_1474 (O_1474,N_19925,N_19944);
and UO_1475 (O_1475,N_19978,N_19987);
and UO_1476 (O_1476,N_19870,N_19991);
xnor UO_1477 (O_1477,N_19987,N_19938);
nand UO_1478 (O_1478,N_19935,N_19948);
xor UO_1479 (O_1479,N_19918,N_19983);
nand UO_1480 (O_1480,N_19847,N_19843);
nand UO_1481 (O_1481,N_19965,N_19844);
nand UO_1482 (O_1482,N_19909,N_19981);
and UO_1483 (O_1483,N_19842,N_19891);
nor UO_1484 (O_1484,N_19881,N_19857);
xnor UO_1485 (O_1485,N_19955,N_19918);
nor UO_1486 (O_1486,N_19974,N_19873);
nor UO_1487 (O_1487,N_19915,N_19868);
or UO_1488 (O_1488,N_19841,N_19944);
and UO_1489 (O_1489,N_19993,N_19851);
xor UO_1490 (O_1490,N_19944,N_19988);
nand UO_1491 (O_1491,N_19880,N_19918);
nand UO_1492 (O_1492,N_19978,N_19946);
nand UO_1493 (O_1493,N_19998,N_19974);
nor UO_1494 (O_1494,N_19976,N_19842);
or UO_1495 (O_1495,N_19960,N_19877);
or UO_1496 (O_1496,N_19856,N_19883);
and UO_1497 (O_1497,N_19871,N_19935);
nor UO_1498 (O_1498,N_19854,N_19980);
and UO_1499 (O_1499,N_19994,N_19947);
nand UO_1500 (O_1500,N_19878,N_19961);
nand UO_1501 (O_1501,N_19893,N_19955);
nor UO_1502 (O_1502,N_19884,N_19883);
nand UO_1503 (O_1503,N_19981,N_19966);
xor UO_1504 (O_1504,N_19997,N_19947);
or UO_1505 (O_1505,N_19904,N_19953);
and UO_1506 (O_1506,N_19950,N_19840);
or UO_1507 (O_1507,N_19917,N_19866);
and UO_1508 (O_1508,N_19859,N_19991);
nand UO_1509 (O_1509,N_19974,N_19875);
nand UO_1510 (O_1510,N_19879,N_19988);
nor UO_1511 (O_1511,N_19989,N_19923);
nand UO_1512 (O_1512,N_19872,N_19962);
xor UO_1513 (O_1513,N_19900,N_19940);
or UO_1514 (O_1514,N_19856,N_19843);
nor UO_1515 (O_1515,N_19851,N_19882);
and UO_1516 (O_1516,N_19910,N_19940);
and UO_1517 (O_1517,N_19891,N_19953);
or UO_1518 (O_1518,N_19974,N_19953);
and UO_1519 (O_1519,N_19999,N_19905);
or UO_1520 (O_1520,N_19861,N_19925);
xnor UO_1521 (O_1521,N_19970,N_19959);
xor UO_1522 (O_1522,N_19868,N_19972);
nand UO_1523 (O_1523,N_19938,N_19975);
or UO_1524 (O_1524,N_19915,N_19967);
nand UO_1525 (O_1525,N_19990,N_19857);
and UO_1526 (O_1526,N_19988,N_19840);
xnor UO_1527 (O_1527,N_19935,N_19870);
and UO_1528 (O_1528,N_19926,N_19953);
and UO_1529 (O_1529,N_19923,N_19955);
nor UO_1530 (O_1530,N_19923,N_19870);
and UO_1531 (O_1531,N_19931,N_19855);
xnor UO_1532 (O_1532,N_19949,N_19975);
nor UO_1533 (O_1533,N_19922,N_19905);
nor UO_1534 (O_1534,N_19892,N_19913);
or UO_1535 (O_1535,N_19969,N_19937);
nand UO_1536 (O_1536,N_19923,N_19975);
nand UO_1537 (O_1537,N_19855,N_19960);
nor UO_1538 (O_1538,N_19892,N_19857);
nand UO_1539 (O_1539,N_19968,N_19886);
xor UO_1540 (O_1540,N_19861,N_19929);
nand UO_1541 (O_1541,N_19929,N_19982);
or UO_1542 (O_1542,N_19960,N_19873);
nand UO_1543 (O_1543,N_19998,N_19966);
or UO_1544 (O_1544,N_19874,N_19886);
nand UO_1545 (O_1545,N_19892,N_19885);
xor UO_1546 (O_1546,N_19964,N_19908);
and UO_1547 (O_1547,N_19990,N_19898);
and UO_1548 (O_1548,N_19955,N_19879);
or UO_1549 (O_1549,N_19863,N_19846);
or UO_1550 (O_1550,N_19891,N_19969);
and UO_1551 (O_1551,N_19924,N_19859);
nand UO_1552 (O_1552,N_19898,N_19939);
xor UO_1553 (O_1553,N_19882,N_19856);
nand UO_1554 (O_1554,N_19841,N_19879);
nand UO_1555 (O_1555,N_19875,N_19990);
xnor UO_1556 (O_1556,N_19947,N_19972);
xor UO_1557 (O_1557,N_19867,N_19960);
nand UO_1558 (O_1558,N_19994,N_19942);
nor UO_1559 (O_1559,N_19964,N_19875);
nor UO_1560 (O_1560,N_19921,N_19982);
or UO_1561 (O_1561,N_19898,N_19955);
and UO_1562 (O_1562,N_19913,N_19917);
or UO_1563 (O_1563,N_19870,N_19965);
xnor UO_1564 (O_1564,N_19869,N_19926);
nor UO_1565 (O_1565,N_19896,N_19956);
xnor UO_1566 (O_1566,N_19991,N_19964);
and UO_1567 (O_1567,N_19885,N_19886);
nor UO_1568 (O_1568,N_19958,N_19879);
or UO_1569 (O_1569,N_19900,N_19987);
and UO_1570 (O_1570,N_19986,N_19861);
and UO_1571 (O_1571,N_19933,N_19934);
or UO_1572 (O_1572,N_19841,N_19916);
or UO_1573 (O_1573,N_19950,N_19941);
xor UO_1574 (O_1574,N_19861,N_19959);
nor UO_1575 (O_1575,N_19970,N_19976);
or UO_1576 (O_1576,N_19909,N_19935);
or UO_1577 (O_1577,N_19898,N_19940);
or UO_1578 (O_1578,N_19896,N_19873);
nand UO_1579 (O_1579,N_19964,N_19978);
or UO_1580 (O_1580,N_19948,N_19875);
xor UO_1581 (O_1581,N_19958,N_19960);
nor UO_1582 (O_1582,N_19870,N_19911);
nor UO_1583 (O_1583,N_19889,N_19981);
nor UO_1584 (O_1584,N_19887,N_19956);
and UO_1585 (O_1585,N_19951,N_19884);
nand UO_1586 (O_1586,N_19861,N_19928);
nand UO_1587 (O_1587,N_19872,N_19873);
or UO_1588 (O_1588,N_19983,N_19916);
nor UO_1589 (O_1589,N_19940,N_19999);
nor UO_1590 (O_1590,N_19901,N_19858);
or UO_1591 (O_1591,N_19884,N_19984);
and UO_1592 (O_1592,N_19935,N_19869);
and UO_1593 (O_1593,N_19932,N_19928);
nor UO_1594 (O_1594,N_19873,N_19842);
or UO_1595 (O_1595,N_19931,N_19970);
xor UO_1596 (O_1596,N_19990,N_19873);
nor UO_1597 (O_1597,N_19942,N_19966);
xnor UO_1598 (O_1598,N_19991,N_19941);
nor UO_1599 (O_1599,N_19956,N_19892);
and UO_1600 (O_1600,N_19939,N_19874);
or UO_1601 (O_1601,N_19926,N_19971);
xor UO_1602 (O_1602,N_19895,N_19987);
or UO_1603 (O_1603,N_19935,N_19924);
nand UO_1604 (O_1604,N_19921,N_19894);
or UO_1605 (O_1605,N_19858,N_19930);
or UO_1606 (O_1606,N_19898,N_19988);
nand UO_1607 (O_1607,N_19955,N_19888);
nor UO_1608 (O_1608,N_19857,N_19890);
nor UO_1609 (O_1609,N_19925,N_19961);
nand UO_1610 (O_1610,N_19888,N_19852);
or UO_1611 (O_1611,N_19871,N_19947);
xnor UO_1612 (O_1612,N_19961,N_19932);
or UO_1613 (O_1613,N_19976,N_19861);
or UO_1614 (O_1614,N_19858,N_19868);
xnor UO_1615 (O_1615,N_19958,N_19916);
xnor UO_1616 (O_1616,N_19955,N_19958);
nor UO_1617 (O_1617,N_19902,N_19875);
or UO_1618 (O_1618,N_19867,N_19933);
xnor UO_1619 (O_1619,N_19871,N_19845);
nand UO_1620 (O_1620,N_19867,N_19907);
nand UO_1621 (O_1621,N_19903,N_19950);
and UO_1622 (O_1622,N_19931,N_19936);
nand UO_1623 (O_1623,N_19981,N_19859);
or UO_1624 (O_1624,N_19868,N_19867);
and UO_1625 (O_1625,N_19915,N_19874);
nand UO_1626 (O_1626,N_19989,N_19883);
nor UO_1627 (O_1627,N_19918,N_19877);
nand UO_1628 (O_1628,N_19893,N_19877);
nand UO_1629 (O_1629,N_19946,N_19878);
and UO_1630 (O_1630,N_19870,N_19885);
nand UO_1631 (O_1631,N_19930,N_19898);
or UO_1632 (O_1632,N_19890,N_19846);
and UO_1633 (O_1633,N_19876,N_19867);
nor UO_1634 (O_1634,N_19887,N_19967);
and UO_1635 (O_1635,N_19877,N_19904);
nand UO_1636 (O_1636,N_19842,N_19898);
nand UO_1637 (O_1637,N_19885,N_19852);
nand UO_1638 (O_1638,N_19940,N_19843);
nand UO_1639 (O_1639,N_19968,N_19844);
xnor UO_1640 (O_1640,N_19991,N_19998);
nand UO_1641 (O_1641,N_19867,N_19913);
nand UO_1642 (O_1642,N_19958,N_19842);
and UO_1643 (O_1643,N_19853,N_19935);
nor UO_1644 (O_1644,N_19976,N_19954);
xor UO_1645 (O_1645,N_19942,N_19962);
nor UO_1646 (O_1646,N_19950,N_19868);
xor UO_1647 (O_1647,N_19853,N_19943);
and UO_1648 (O_1648,N_19989,N_19907);
nor UO_1649 (O_1649,N_19873,N_19978);
xnor UO_1650 (O_1650,N_19863,N_19918);
and UO_1651 (O_1651,N_19859,N_19890);
or UO_1652 (O_1652,N_19932,N_19967);
and UO_1653 (O_1653,N_19890,N_19896);
or UO_1654 (O_1654,N_19869,N_19944);
nor UO_1655 (O_1655,N_19978,N_19912);
and UO_1656 (O_1656,N_19908,N_19896);
and UO_1657 (O_1657,N_19912,N_19958);
and UO_1658 (O_1658,N_19919,N_19850);
xnor UO_1659 (O_1659,N_19946,N_19943);
and UO_1660 (O_1660,N_19967,N_19923);
nor UO_1661 (O_1661,N_19920,N_19925);
nand UO_1662 (O_1662,N_19966,N_19867);
or UO_1663 (O_1663,N_19950,N_19853);
or UO_1664 (O_1664,N_19979,N_19946);
or UO_1665 (O_1665,N_19932,N_19887);
and UO_1666 (O_1666,N_19867,N_19840);
or UO_1667 (O_1667,N_19999,N_19849);
nor UO_1668 (O_1668,N_19993,N_19919);
xnor UO_1669 (O_1669,N_19871,N_19918);
or UO_1670 (O_1670,N_19985,N_19998);
or UO_1671 (O_1671,N_19903,N_19998);
or UO_1672 (O_1672,N_19844,N_19859);
or UO_1673 (O_1673,N_19981,N_19991);
or UO_1674 (O_1674,N_19938,N_19918);
nand UO_1675 (O_1675,N_19883,N_19979);
nor UO_1676 (O_1676,N_19941,N_19916);
xor UO_1677 (O_1677,N_19983,N_19886);
nand UO_1678 (O_1678,N_19960,N_19999);
and UO_1679 (O_1679,N_19857,N_19919);
xnor UO_1680 (O_1680,N_19979,N_19996);
or UO_1681 (O_1681,N_19882,N_19889);
nand UO_1682 (O_1682,N_19960,N_19899);
nand UO_1683 (O_1683,N_19983,N_19954);
nand UO_1684 (O_1684,N_19893,N_19927);
nor UO_1685 (O_1685,N_19915,N_19985);
nor UO_1686 (O_1686,N_19904,N_19980);
nand UO_1687 (O_1687,N_19987,N_19939);
nor UO_1688 (O_1688,N_19927,N_19890);
and UO_1689 (O_1689,N_19936,N_19982);
nor UO_1690 (O_1690,N_19952,N_19932);
nor UO_1691 (O_1691,N_19969,N_19886);
or UO_1692 (O_1692,N_19959,N_19918);
xor UO_1693 (O_1693,N_19964,N_19888);
nand UO_1694 (O_1694,N_19876,N_19978);
and UO_1695 (O_1695,N_19854,N_19871);
nor UO_1696 (O_1696,N_19888,N_19851);
xnor UO_1697 (O_1697,N_19975,N_19922);
and UO_1698 (O_1698,N_19907,N_19969);
nand UO_1699 (O_1699,N_19863,N_19856);
nor UO_1700 (O_1700,N_19985,N_19857);
nand UO_1701 (O_1701,N_19890,N_19941);
nor UO_1702 (O_1702,N_19999,N_19928);
nor UO_1703 (O_1703,N_19887,N_19873);
and UO_1704 (O_1704,N_19846,N_19954);
nor UO_1705 (O_1705,N_19883,N_19969);
xor UO_1706 (O_1706,N_19885,N_19919);
xnor UO_1707 (O_1707,N_19936,N_19956);
xnor UO_1708 (O_1708,N_19947,N_19904);
nor UO_1709 (O_1709,N_19947,N_19854);
nor UO_1710 (O_1710,N_19943,N_19922);
nand UO_1711 (O_1711,N_19875,N_19866);
or UO_1712 (O_1712,N_19947,N_19988);
xnor UO_1713 (O_1713,N_19916,N_19994);
nand UO_1714 (O_1714,N_19872,N_19923);
and UO_1715 (O_1715,N_19951,N_19952);
xnor UO_1716 (O_1716,N_19975,N_19878);
xor UO_1717 (O_1717,N_19994,N_19971);
or UO_1718 (O_1718,N_19848,N_19886);
nor UO_1719 (O_1719,N_19905,N_19866);
or UO_1720 (O_1720,N_19876,N_19990);
or UO_1721 (O_1721,N_19893,N_19958);
and UO_1722 (O_1722,N_19890,N_19911);
nand UO_1723 (O_1723,N_19996,N_19980);
xor UO_1724 (O_1724,N_19943,N_19917);
and UO_1725 (O_1725,N_19847,N_19840);
and UO_1726 (O_1726,N_19967,N_19900);
nor UO_1727 (O_1727,N_19857,N_19975);
nor UO_1728 (O_1728,N_19949,N_19876);
and UO_1729 (O_1729,N_19870,N_19850);
nor UO_1730 (O_1730,N_19985,N_19900);
or UO_1731 (O_1731,N_19968,N_19862);
and UO_1732 (O_1732,N_19862,N_19966);
nand UO_1733 (O_1733,N_19982,N_19985);
xnor UO_1734 (O_1734,N_19846,N_19898);
and UO_1735 (O_1735,N_19954,N_19939);
xor UO_1736 (O_1736,N_19868,N_19853);
xnor UO_1737 (O_1737,N_19915,N_19846);
or UO_1738 (O_1738,N_19992,N_19950);
or UO_1739 (O_1739,N_19960,N_19912);
xnor UO_1740 (O_1740,N_19856,N_19849);
and UO_1741 (O_1741,N_19995,N_19971);
nand UO_1742 (O_1742,N_19965,N_19849);
and UO_1743 (O_1743,N_19857,N_19918);
nor UO_1744 (O_1744,N_19930,N_19841);
and UO_1745 (O_1745,N_19857,N_19858);
xor UO_1746 (O_1746,N_19915,N_19857);
and UO_1747 (O_1747,N_19968,N_19917);
and UO_1748 (O_1748,N_19939,N_19917);
and UO_1749 (O_1749,N_19867,N_19968);
nand UO_1750 (O_1750,N_19883,N_19891);
or UO_1751 (O_1751,N_19957,N_19976);
and UO_1752 (O_1752,N_19915,N_19893);
and UO_1753 (O_1753,N_19989,N_19859);
or UO_1754 (O_1754,N_19913,N_19882);
nand UO_1755 (O_1755,N_19972,N_19855);
xnor UO_1756 (O_1756,N_19948,N_19947);
nand UO_1757 (O_1757,N_19962,N_19899);
nor UO_1758 (O_1758,N_19897,N_19864);
xor UO_1759 (O_1759,N_19968,N_19956);
xor UO_1760 (O_1760,N_19942,N_19961);
xor UO_1761 (O_1761,N_19956,N_19952);
nand UO_1762 (O_1762,N_19971,N_19931);
xnor UO_1763 (O_1763,N_19926,N_19866);
and UO_1764 (O_1764,N_19946,N_19916);
xnor UO_1765 (O_1765,N_19931,N_19937);
and UO_1766 (O_1766,N_19990,N_19900);
nand UO_1767 (O_1767,N_19918,N_19905);
and UO_1768 (O_1768,N_19875,N_19931);
xnor UO_1769 (O_1769,N_19843,N_19867);
nor UO_1770 (O_1770,N_19869,N_19943);
nor UO_1771 (O_1771,N_19921,N_19953);
nand UO_1772 (O_1772,N_19973,N_19891);
and UO_1773 (O_1773,N_19872,N_19925);
and UO_1774 (O_1774,N_19854,N_19853);
xor UO_1775 (O_1775,N_19858,N_19850);
xnor UO_1776 (O_1776,N_19906,N_19888);
and UO_1777 (O_1777,N_19905,N_19870);
or UO_1778 (O_1778,N_19985,N_19971);
nor UO_1779 (O_1779,N_19933,N_19936);
and UO_1780 (O_1780,N_19988,N_19874);
nor UO_1781 (O_1781,N_19856,N_19894);
and UO_1782 (O_1782,N_19994,N_19902);
nor UO_1783 (O_1783,N_19976,N_19879);
xnor UO_1784 (O_1784,N_19895,N_19982);
nor UO_1785 (O_1785,N_19863,N_19898);
nand UO_1786 (O_1786,N_19979,N_19889);
and UO_1787 (O_1787,N_19961,N_19903);
nand UO_1788 (O_1788,N_19933,N_19996);
and UO_1789 (O_1789,N_19849,N_19998);
nor UO_1790 (O_1790,N_19946,N_19902);
nor UO_1791 (O_1791,N_19910,N_19973);
nand UO_1792 (O_1792,N_19908,N_19992);
nand UO_1793 (O_1793,N_19935,N_19987);
and UO_1794 (O_1794,N_19975,N_19899);
and UO_1795 (O_1795,N_19917,N_19849);
nor UO_1796 (O_1796,N_19967,N_19921);
nor UO_1797 (O_1797,N_19872,N_19959);
xnor UO_1798 (O_1798,N_19947,N_19973);
xnor UO_1799 (O_1799,N_19926,N_19951);
nand UO_1800 (O_1800,N_19954,N_19946);
and UO_1801 (O_1801,N_19914,N_19910);
nor UO_1802 (O_1802,N_19849,N_19961);
nor UO_1803 (O_1803,N_19991,N_19985);
and UO_1804 (O_1804,N_19957,N_19861);
xor UO_1805 (O_1805,N_19954,N_19943);
xor UO_1806 (O_1806,N_19924,N_19965);
xor UO_1807 (O_1807,N_19993,N_19983);
nor UO_1808 (O_1808,N_19846,N_19959);
nand UO_1809 (O_1809,N_19987,N_19901);
nand UO_1810 (O_1810,N_19964,N_19840);
nand UO_1811 (O_1811,N_19893,N_19919);
and UO_1812 (O_1812,N_19955,N_19996);
nand UO_1813 (O_1813,N_19843,N_19969);
or UO_1814 (O_1814,N_19906,N_19867);
nand UO_1815 (O_1815,N_19937,N_19902);
and UO_1816 (O_1816,N_19889,N_19897);
or UO_1817 (O_1817,N_19973,N_19923);
nor UO_1818 (O_1818,N_19898,N_19869);
nand UO_1819 (O_1819,N_19962,N_19969);
or UO_1820 (O_1820,N_19936,N_19883);
nand UO_1821 (O_1821,N_19932,N_19869);
nand UO_1822 (O_1822,N_19914,N_19994);
xnor UO_1823 (O_1823,N_19951,N_19847);
nor UO_1824 (O_1824,N_19848,N_19999);
and UO_1825 (O_1825,N_19863,N_19929);
or UO_1826 (O_1826,N_19888,N_19847);
xnor UO_1827 (O_1827,N_19951,N_19843);
nand UO_1828 (O_1828,N_19983,N_19841);
nand UO_1829 (O_1829,N_19850,N_19884);
and UO_1830 (O_1830,N_19918,N_19843);
and UO_1831 (O_1831,N_19866,N_19952);
or UO_1832 (O_1832,N_19923,N_19899);
nand UO_1833 (O_1833,N_19936,N_19847);
and UO_1834 (O_1834,N_19888,N_19846);
and UO_1835 (O_1835,N_19890,N_19935);
xor UO_1836 (O_1836,N_19856,N_19918);
nand UO_1837 (O_1837,N_19933,N_19990);
nor UO_1838 (O_1838,N_19934,N_19938);
nand UO_1839 (O_1839,N_19905,N_19924);
or UO_1840 (O_1840,N_19964,N_19848);
and UO_1841 (O_1841,N_19933,N_19930);
or UO_1842 (O_1842,N_19856,N_19967);
and UO_1843 (O_1843,N_19949,N_19862);
nor UO_1844 (O_1844,N_19899,N_19971);
xor UO_1845 (O_1845,N_19847,N_19983);
nor UO_1846 (O_1846,N_19959,N_19911);
and UO_1847 (O_1847,N_19931,N_19846);
nor UO_1848 (O_1848,N_19945,N_19877);
and UO_1849 (O_1849,N_19881,N_19853);
nor UO_1850 (O_1850,N_19866,N_19960);
nor UO_1851 (O_1851,N_19939,N_19946);
and UO_1852 (O_1852,N_19993,N_19930);
or UO_1853 (O_1853,N_19862,N_19991);
or UO_1854 (O_1854,N_19890,N_19999);
nor UO_1855 (O_1855,N_19972,N_19993);
nor UO_1856 (O_1856,N_19869,N_19962);
nand UO_1857 (O_1857,N_19993,N_19951);
or UO_1858 (O_1858,N_19987,N_19850);
xnor UO_1859 (O_1859,N_19966,N_19920);
and UO_1860 (O_1860,N_19856,N_19909);
nor UO_1861 (O_1861,N_19911,N_19982);
and UO_1862 (O_1862,N_19890,N_19905);
nand UO_1863 (O_1863,N_19895,N_19966);
nand UO_1864 (O_1864,N_19940,N_19930);
nor UO_1865 (O_1865,N_19933,N_19921);
and UO_1866 (O_1866,N_19942,N_19842);
or UO_1867 (O_1867,N_19963,N_19881);
nand UO_1868 (O_1868,N_19970,N_19974);
nor UO_1869 (O_1869,N_19939,N_19911);
and UO_1870 (O_1870,N_19913,N_19877);
and UO_1871 (O_1871,N_19983,N_19999);
xnor UO_1872 (O_1872,N_19883,N_19865);
xor UO_1873 (O_1873,N_19951,N_19891);
xor UO_1874 (O_1874,N_19975,N_19998);
nand UO_1875 (O_1875,N_19975,N_19987);
nand UO_1876 (O_1876,N_19947,N_19959);
nand UO_1877 (O_1877,N_19843,N_19990);
or UO_1878 (O_1878,N_19871,N_19932);
xnor UO_1879 (O_1879,N_19904,N_19951);
xnor UO_1880 (O_1880,N_19949,N_19993);
nand UO_1881 (O_1881,N_19920,N_19916);
nor UO_1882 (O_1882,N_19983,N_19935);
xnor UO_1883 (O_1883,N_19899,N_19935);
and UO_1884 (O_1884,N_19982,N_19885);
and UO_1885 (O_1885,N_19927,N_19980);
and UO_1886 (O_1886,N_19870,N_19976);
nor UO_1887 (O_1887,N_19863,N_19860);
or UO_1888 (O_1888,N_19906,N_19981);
xor UO_1889 (O_1889,N_19914,N_19919);
and UO_1890 (O_1890,N_19893,N_19854);
nand UO_1891 (O_1891,N_19859,N_19926);
nor UO_1892 (O_1892,N_19979,N_19916);
and UO_1893 (O_1893,N_19880,N_19929);
nor UO_1894 (O_1894,N_19891,N_19909);
nor UO_1895 (O_1895,N_19904,N_19942);
nand UO_1896 (O_1896,N_19944,N_19842);
and UO_1897 (O_1897,N_19989,N_19974);
and UO_1898 (O_1898,N_19972,N_19984);
nor UO_1899 (O_1899,N_19969,N_19987);
and UO_1900 (O_1900,N_19871,N_19997);
xor UO_1901 (O_1901,N_19917,N_19903);
nor UO_1902 (O_1902,N_19892,N_19855);
and UO_1903 (O_1903,N_19922,N_19981);
and UO_1904 (O_1904,N_19928,N_19856);
or UO_1905 (O_1905,N_19953,N_19913);
and UO_1906 (O_1906,N_19907,N_19990);
or UO_1907 (O_1907,N_19840,N_19862);
or UO_1908 (O_1908,N_19844,N_19925);
nor UO_1909 (O_1909,N_19965,N_19920);
or UO_1910 (O_1910,N_19950,N_19870);
or UO_1911 (O_1911,N_19946,N_19924);
xor UO_1912 (O_1912,N_19921,N_19958);
xnor UO_1913 (O_1913,N_19877,N_19863);
xor UO_1914 (O_1914,N_19940,N_19972);
nand UO_1915 (O_1915,N_19860,N_19920);
or UO_1916 (O_1916,N_19976,N_19980);
xnor UO_1917 (O_1917,N_19909,N_19997);
xnor UO_1918 (O_1918,N_19970,N_19886);
nor UO_1919 (O_1919,N_19995,N_19982);
and UO_1920 (O_1920,N_19895,N_19964);
nor UO_1921 (O_1921,N_19896,N_19867);
and UO_1922 (O_1922,N_19921,N_19861);
and UO_1923 (O_1923,N_19879,N_19915);
nand UO_1924 (O_1924,N_19914,N_19872);
and UO_1925 (O_1925,N_19950,N_19993);
nor UO_1926 (O_1926,N_19873,N_19964);
nor UO_1927 (O_1927,N_19981,N_19856);
and UO_1928 (O_1928,N_19843,N_19897);
nor UO_1929 (O_1929,N_19912,N_19972);
nor UO_1930 (O_1930,N_19973,N_19969);
and UO_1931 (O_1931,N_19949,N_19912);
xnor UO_1932 (O_1932,N_19989,N_19857);
xor UO_1933 (O_1933,N_19922,N_19916);
xnor UO_1934 (O_1934,N_19905,N_19861);
nand UO_1935 (O_1935,N_19995,N_19949);
or UO_1936 (O_1936,N_19950,N_19847);
or UO_1937 (O_1937,N_19901,N_19891);
nor UO_1938 (O_1938,N_19887,N_19929);
nor UO_1939 (O_1939,N_19894,N_19948);
or UO_1940 (O_1940,N_19881,N_19960);
and UO_1941 (O_1941,N_19873,N_19939);
nor UO_1942 (O_1942,N_19961,N_19959);
nor UO_1943 (O_1943,N_19957,N_19956);
or UO_1944 (O_1944,N_19873,N_19970);
xnor UO_1945 (O_1945,N_19928,N_19973);
or UO_1946 (O_1946,N_19957,N_19920);
and UO_1947 (O_1947,N_19971,N_19873);
nand UO_1948 (O_1948,N_19915,N_19934);
and UO_1949 (O_1949,N_19916,N_19924);
nand UO_1950 (O_1950,N_19849,N_19967);
nor UO_1951 (O_1951,N_19945,N_19896);
nand UO_1952 (O_1952,N_19940,N_19981);
or UO_1953 (O_1953,N_19927,N_19912);
nand UO_1954 (O_1954,N_19925,N_19865);
nor UO_1955 (O_1955,N_19989,N_19941);
nor UO_1956 (O_1956,N_19932,N_19929);
xor UO_1957 (O_1957,N_19928,N_19969);
and UO_1958 (O_1958,N_19937,N_19853);
nand UO_1959 (O_1959,N_19979,N_19890);
xor UO_1960 (O_1960,N_19844,N_19880);
or UO_1961 (O_1961,N_19998,N_19979);
and UO_1962 (O_1962,N_19981,N_19950);
xor UO_1963 (O_1963,N_19973,N_19968);
or UO_1964 (O_1964,N_19878,N_19887);
nor UO_1965 (O_1965,N_19994,N_19887);
xor UO_1966 (O_1966,N_19905,N_19913);
or UO_1967 (O_1967,N_19850,N_19935);
nor UO_1968 (O_1968,N_19926,N_19957);
and UO_1969 (O_1969,N_19847,N_19953);
xnor UO_1970 (O_1970,N_19946,N_19862);
xor UO_1971 (O_1971,N_19943,N_19896);
and UO_1972 (O_1972,N_19911,N_19865);
nand UO_1973 (O_1973,N_19844,N_19945);
and UO_1974 (O_1974,N_19900,N_19995);
xor UO_1975 (O_1975,N_19955,N_19979);
and UO_1976 (O_1976,N_19869,N_19992);
or UO_1977 (O_1977,N_19933,N_19848);
or UO_1978 (O_1978,N_19853,N_19873);
nand UO_1979 (O_1979,N_19847,N_19964);
nand UO_1980 (O_1980,N_19876,N_19866);
xnor UO_1981 (O_1981,N_19934,N_19945);
nand UO_1982 (O_1982,N_19989,N_19999);
xnor UO_1983 (O_1983,N_19947,N_19925);
xnor UO_1984 (O_1984,N_19946,N_19968);
nor UO_1985 (O_1985,N_19893,N_19978);
nor UO_1986 (O_1986,N_19969,N_19948);
and UO_1987 (O_1987,N_19877,N_19948);
nand UO_1988 (O_1988,N_19886,N_19865);
or UO_1989 (O_1989,N_19855,N_19927);
xnor UO_1990 (O_1990,N_19988,N_19871);
nor UO_1991 (O_1991,N_19932,N_19900);
nor UO_1992 (O_1992,N_19984,N_19955);
nor UO_1993 (O_1993,N_19855,N_19926);
xor UO_1994 (O_1994,N_19923,N_19982);
and UO_1995 (O_1995,N_19970,N_19986);
nand UO_1996 (O_1996,N_19849,N_19924);
or UO_1997 (O_1997,N_19888,N_19862);
or UO_1998 (O_1998,N_19927,N_19996);
xnor UO_1999 (O_1999,N_19937,N_19927);
nor UO_2000 (O_2000,N_19897,N_19951);
xnor UO_2001 (O_2001,N_19986,N_19853);
xor UO_2002 (O_2002,N_19917,N_19927);
nand UO_2003 (O_2003,N_19993,N_19883);
and UO_2004 (O_2004,N_19858,N_19972);
xnor UO_2005 (O_2005,N_19977,N_19973);
and UO_2006 (O_2006,N_19931,N_19872);
nand UO_2007 (O_2007,N_19884,N_19966);
and UO_2008 (O_2008,N_19893,N_19846);
xnor UO_2009 (O_2009,N_19970,N_19973);
nand UO_2010 (O_2010,N_19880,N_19840);
and UO_2011 (O_2011,N_19849,N_19973);
nand UO_2012 (O_2012,N_19908,N_19902);
or UO_2013 (O_2013,N_19883,N_19937);
or UO_2014 (O_2014,N_19897,N_19928);
nor UO_2015 (O_2015,N_19856,N_19954);
nand UO_2016 (O_2016,N_19960,N_19903);
xnor UO_2017 (O_2017,N_19965,N_19921);
nand UO_2018 (O_2018,N_19990,N_19891);
nor UO_2019 (O_2019,N_19915,N_19865);
and UO_2020 (O_2020,N_19988,N_19883);
and UO_2021 (O_2021,N_19902,N_19926);
nand UO_2022 (O_2022,N_19843,N_19981);
and UO_2023 (O_2023,N_19904,N_19928);
nor UO_2024 (O_2024,N_19902,N_19993);
or UO_2025 (O_2025,N_19994,N_19983);
nand UO_2026 (O_2026,N_19884,N_19941);
xor UO_2027 (O_2027,N_19911,N_19925);
nand UO_2028 (O_2028,N_19881,N_19938);
or UO_2029 (O_2029,N_19975,N_19844);
and UO_2030 (O_2030,N_19976,N_19930);
nand UO_2031 (O_2031,N_19855,N_19934);
nand UO_2032 (O_2032,N_19895,N_19935);
nor UO_2033 (O_2033,N_19990,N_19971);
or UO_2034 (O_2034,N_19877,N_19856);
and UO_2035 (O_2035,N_19931,N_19848);
xor UO_2036 (O_2036,N_19909,N_19969);
nand UO_2037 (O_2037,N_19980,N_19894);
nor UO_2038 (O_2038,N_19898,N_19954);
and UO_2039 (O_2039,N_19986,N_19908);
xnor UO_2040 (O_2040,N_19894,N_19906);
or UO_2041 (O_2041,N_19870,N_19851);
or UO_2042 (O_2042,N_19872,N_19840);
and UO_2043 (O_2043,N_19845,N_19918);
and UO_2044 (O_2044,N_19884,N_19871);
xor UO_2045 (O_2045,N_19842,N_19855);
nand UO_2046 (O_2046,N_19956,N_19980);
xnor UO_2047 (O_2047,N_19965,N_19986);
nor UO_2048 (O_2048,N_19852,N_19981);
and UO_2049 (O_2049,N_19872,N_19881);
and UO_2050 (O_2050,N_19940,N_19896);
nand UO_2051 (O_2051,N_19990,N_19849);
or UO_2052 (O_2052,N_19971,N_19860);
and UO_2053 (O_2053,N_19920,N_19885);
and UO_2054 (O_2054,N_19940,N_19879);
and UO_2055 (O_2055,N_19898,N_19980);
nor UO_2056 (O_2056,N_19893,N_19968);
nor UO_2057 (O_2057,N_19989,N_19871);
and UO_2058 (O_2058,N_19960,N_19856);
xor UO_2059 (O_2059,N_19882,N_19901);
or UO_2060 (O_2060,N_19898,N_19991);
nand UO_2061 (O_2061,N_19922,N_19867);
xnor UO_2062 (O_2062,N_19878,N_19893);
nand UO_2063 (O_2063,N_19924,N_19881);
xnor UO_2064 (O_2064,N_19959,N_19863);
xnor UO_2065 (O_2065,N_19940,N_19852);
or UO_2066 (O_2066,N_19888,N_19985);
or UO_2067 (O_2067,N_19975,N_19950);
nand UO_2068 (O_2068,N_19911,N_19896);
nor UO_2069 (O_2069,N_19889,N_19903);
nand UO_2070 (O_2070,N_19885,N_19935);
and UO_2071 (O_2071,N_19868,N_19996);
nand UO_2072 (O_2072,N_19919,N_19867);
nor UO_2073 (O_2073,N_19857,N_19973);
nand UO_2074 (O_2074,N_19999,N_19972);
or UO_2075 (O_2075,N_19958,N_19997);
and UO_2076 (O_2076,N_19845,N_19943);
xor UO_2077 (O_2077,N_19920,N_19866);
and UO_2078 (O_2078,N_19937,N_19950);
nand UO_2079 (O_2079,N_19868,N_19914);
or UO_2080 (O_2080,N_19983,N_19840);
nor UO_2081 (O_2081,N_19946,N_19927);
or UO_2082 (O_2082,N_19873,N_19969);
or UO_2083 (O_2083,N_19870,N_19963);
xnor UO_2084 (O_2084,N_19956,N_19934);
xnor UO_2085 (O_2085,N_19999,N_19871);
nand UO_2086 (O_2086,N_19961,N_19965);
and UO_2087 (O_2087,N_19865,N_19867);
xnor UO_2088 (O_2088,N_19929,N_19854);
or UO_2089 (O_2089,N_19864,N_19953);
nand UO_2090 (O_2090,N_19934,N_19861);
nand UO_2091 (O_2091,N_19872,N_19858);
xnor UO_2092 (O_2092,N_19967,N_19981);
and UO_2093 (O_2093,N_19914,N_19990);
xor UO_2094 (O_2094,N_19935,N_19963);
nor UO_2095 (O_2095,N_19845,N_19878);
or UO_2096 (O_2096,N_19906,N_19968);
nor UO_2097 (O_2097,N_19907,N_19957);
or UO_2098 (O_2098,N_19843,N_19868);
nand UO_2099 (O_2099,N_19950,N_19962);
or UO_2100 (O_2100,N_19952,N_19925);
nand UO_2101 (O_2101,N_19885,N_19883);
or UO_2102 (O_2102,N_19905,N_19993);
or UO_2103 (O_2103,N_19930,N_19984);
xnor UO_2104 (O_2104,N_19981,N_19895);
nand UO_2105 (O_2105,N_19906,N_19920);
nor UO_2106 (O_2106,N_19846,N_19860);
nand UO_2107 (O_2107,N_19950,N_19913);
nor UO_2108 (O_2108,N_19926,N_19962);
and UO_2109 (O_2109,N_19986,N_19876);
and UO_2110 (O_2110,N_19842,N_19982);
and UO_2111 (O_2111,N_19904,N_19888);
or UO_2112 (O_2112,N_19918,N_19889);
and UO_2113 (O_2113,N_19868,N_19900);
or UO_2114 (O_2114,N_19895,N_19861);
xnor UO_2115 (O_2115,N_19864,N_19994);
or UO_2116 (O_2116,N_19849,N_19868);
nand UO_2117 (O_2117,N_19853,N_19932);
or UO_2118 (O_2118,N_19974,N_19949);
xnor UO_2119 (O_2119,N_19879,N_19925);
nor UO_2120 (O_2120,N_19919,N_19909);
or UO_2121 (O_2121,N_19879,N_19919);
and UO_2122 (O_2122,N_19932,N_19846);
and UO_2123 (O_2123,N_19950,N_19860);
nand UO_2124 (O_2124,N_19876,N_19996);
or UO_2125 (O_2125,N_19970,N_19989);
nand UO_2126 (O_2126,N_19870,N_19927);
or UO_2127 (O_2127,N_19992,N_19922);
nor UO_2128 (O_2128,N_19845,N_19954);
xor UO_2129 (O_2129,N_19860,N_19932);
nand UO_2130 (O_2130,N_19842,N_19884);
nand UO_2131 (O_2131,N_19883,N_19924);
xnor UO_2132 (O_2132,N_19967,N_19896);
xor UO_2133 (O_2133,N_19910,N_19892);
or UO_2134 (O_2134,N_19972,N_19951);
or UO_2135 (O_2135,N_19949,N_19860);
nand UO_2136 (O_2136,N_19996,N_19873);
nor UO_2137 (O_2137,N_19997,N_19993);
or UO_2138 (O_2138,N_19862,N_19896);
nand UO_2139 (O_2139,N_19871,N_19972);
nand UO_2140 (O_2140,N_19853,N_19860);
and UO_2141 (O_2141,N_19931,N_19980);
xnor UO_2142 (O_2142,N_19928,N_19949);
or UO_2143 (O_2143,N_19846,N_19892);
and UO_2144 (O_2144,N_19950,N_19859);
and UO_2145 (O_2145,N_19868,N_19949);
nor UO_2146 (O_2146,N_19894,N_19975);
and UO_2147 (O_2147,N_19886,N_19919);
and UO_2148 (O_2148,N_19931,N_19926);
nor UO_2149 (O_2149,N_19919,N_19856);
and UO_2150 (O_2150,N_19854,N_19977);
nand UO_2151 (O_2151,N_19988,N_19966);
and UO_2152 (O_2152,N_19970,N_19932);
nor UO_2153 (O_2153,N_19951,N_19899);
and UO_2154 (O_2154,N_19952,N_19986);
or UO_2155 (O_2155,N_19968,N_19846);
or UO_2156 (O_2156,N_19857,N_19885);
nand UO_2157 (O_2157,N_19938,N_19947);
xnor UO_2158 (O_2158,N_19988,N_19868);
xnor UO_2159 (O_2159,N_19983,N_19962);
nand UO_2160 (O_2160,N_19948,N_19907);
or UO_2161 (O_2161,N_19983,N_19884);
nor UO_2162 (O_2162,N_19972,N_19888);
or UO_2163 (O_2163,N_19942,N_19956);
or UO_2164 (O_2164,N_19975,N_19944);
xnor UO_2165 (O_2165,N_19989,N_19876);
nand UO_2166 (O_2166,N_19911,N_19907);
nor UO_2167 (O_2167,N_19972,N_19975);
nor UO_2168 (O_2168,N_19993,N_19854);
and UO_2169 (O_2169,N_19958,N_19979);
xor UO_2170 (O_2170,N_19917,N_19893);
xor UO_2171 (O_2171,N_19925,N_19901);
nand UO_2172 (O_2172,N_19915,N_19938);
nor UO_2173 (O_2173,N_19924,N_19951);
and UO_2174 (O_2174,N_19846,N_19848);
or UO_2175 (O_2175,N_19982,N_19932);
and UO_2176 (O_2176,N_19961,N_19853);
nand UO_2177 (O_2177,N_19961,N_19870);
nand UO_2178 (O_2178,N_19868,N_19873);
nor UO_2179 (O_2179,N_19842,N_19932);
xor UO_2180 (O_2180,N_19873,N_19982);
and UO_2181 (O_2181,N_19899,N_19867);
nand UO_2182 (O_2182,N_19919,N_19897);
xnor UO_2183 (O_2183,N_19926,N_19901);
and UO_2184 (O_2184,N_19974,N_19968);
and UO_2185 (O_2185,N_19992,N_19932);
or UO_2186 (O_2186,N_19981,N_19911);
and UO_2187 (O_2187,N_19981,N_19993);
nor UO_2188 (O_2188,N_19856,N_19896);
or UO_2189 (O_2189,N_19981,N_19930);
or UO_2190 (O_2190,N_19881,N_19851);
nand UO_2191 (O_2191,N_19988,N_19878);
or UO_2192 (O_2192,N_19972,N_19878);
or UO_2193 (O_2193,N_19971,N_19842);
or UO_2194 (O_2194,N_19991,N_19958);
nor UO_2195 (O_2195,N_19986,N_19847);
nand UO_2196 (O_2196,N_19951,N_19990);
xnor UO_2197 (O_2197,N_19948,N_19858);
or UO_2198 (O_2198,N_19884,N_19841);
and UO_2199 (O_2199,N_19854,N_19882);
nor UO_2200 (O_2200,N_19896,N_19976);
nand UO_2201 (O_2201,N_19985,N_19974);
nand UO_2202 (O_2202,N_19869,N_19882);
nand UO_2203 (O_2203,N_19999,N_19971);
or UO_2204 (O_2204,N_19967,N_19864);
and UO_2205 (O_2205,N_19864,N_19846);
nand UO_2206 (O_2206,N_19998,N_19923);
and UO_2207 (O_2207,N_19969,N_19963);
nand UO_2208 (O_2208,N_19897,N_19873);
nor UO_2209 (O_2209,N_19861,N_19918);
or UO_2210 (O_2210,N_19993,N_19842);
and UO_2211 (O_2211,N_19967,N_19908);
nand UO_2212 (O_2212,N_19897,N_19954);
nor UO_2213 (O_2213,N_19953,N_19961);
nor UO_2214 (O_2214,N_19969,N_19991);
and UO_2215 (O_2215,N_19887,N_19995);
xnor UO_2216 (O_2216,N_19991,N_19948);
nor UO_2217 (O_2217,N_19879,N_19948);
or UO_2218 (O_2218,N_19932,N_19878);
or UO_2219 (O_2219,N_19916,N_19855);
or UO_2220 (O_2220,N_19933,N_19855);
or UO_2221 (O_2221,N_19980,N_19880);
nor UO_2222 (O_2222,N_19872,N_19986);
and UO_2223 (O_2223,N_19909,N_19985);
xor UO_2224 (O_2224,N_19846,N_19986);
nand UO_2225 (O_2225,N_19963,N_19936);
nand UO_2226 (O_2226,N_19927,N_19991);
nand UO_2227 (O_2227,N_19963,N_19874);
or UO_2228 (O_2228,N_19969,N_19980);
xnor UO_2229 (O_2229,N_19957,N_19925);
and UO_2230 (O_2230,N_19945,N_19905);
xor UO_2231 (O_2231,N_19932,N_19852);
and UO_2232 (O_2232,N_19909,N_19911);
or UO_2233 (O_2233,N_19854,N_19870);
nand UO_2234 (O_2234,N_19900,N_19958);
nor UO_2235 (O_2235,N_19881,N_19889);
nand UO_2236 (O_2236,N_19948,N_19975);
xnor UO_2237 (O_2237,N_19864,N_19963);
and UO_2238 (O_2238,N_19932,N_19971);
and UO_2239 (O_2239,N_19842,N_19868);
xor UO_2240 (O_2240,N_19921,N_19946);
nor UO_2241 (O_2241,N_19899,N_19845);
nand UO_2242 (O_2242,N_19934,N_19985);
or UO_2243 (O_2243,N_19891,N_19914);
and UO_2244 (O_2244,N_19976,N_19851);
or UO_2245 (O_2245,N_19934,N_19989);
or UO_2246 (O_2246,N_19987,N_19919);
nor UO_2247 (O_2247,N_19998,N_19957);
xor UO_2248 (O_2248,N_19934,N_19968);
nor UO_2249 (O_2249,N_19917,N_19856);
xnor UO_2250 (O_2250,N_19992,N_19966);
nor UO_2251 (O_2251,N_19956,N_19965);
nor UO_2252 (O_2252,N_19924,N_19952);
xnor UO_2253 (O_2253,N_19961,N_19926);
xor UO_2254 (O_2254,N_19968,N_19964);
nor UO_2255 (O_2255,N_19868,N_19951);
nor UO_2256 (O_2256,N_19854,N_19958);
or UO_2257 (O_2257,N_19878,N_19870);
nand UO_2258 (O_2258,N_19887,N_19924);
xnor UO_2259 (O_2259,N_19863,N_19867);
nor UO_2260 (O_2260,N_19945,N_19882);
or UO_2261 (O_2261,N_19905,N_19865);
nand UO_2262 (O_2262,N_19898,N_19897);
or UO_2263 (O_2263,N_19925,N_19958);
nand UO_2264 (O_2264,N_19939,N_19905);
and UO_2265 (O_2265,N_19888,N_19927);
nand UO_2266 (O_2266,N_19902,N_19892);
nor UO_2267 (O_2267,N_19965,N_19846);
xor UO_2268 (O_2268,N_19867,N_19897);
nand UO_2269 (O_2269,N_19996,N_19901);
nand UO_2270 (O_2270,N_19915,N_19982);
nor UO_2271 (O_2271,N_19894,N_19887);
and UO_2272 (O_2272,N_19921,N_19867);
and UO_2273 (O_2273,N_19963,N_19847);
nand UO_2274 (O_2274,N_19929,N_19935);
xnor UO_2275 (O_2275,N_19931,N_19903);
nand UO_2276 (O_2276,N_19886,N_19934);
and UO_2277 (O_2277,N_19944,N_19856);
or UO_2278 (O_2278,N_19885,N_19969);
or UO_2279 (O_2279,N_19887,N_19895);
or UO_2280 (O_2280,N_19888,N_19930);
nand UO_2281 (O_2281,N_19904,N_19842);
or UO_2282 (O_2282,N_19940,N_19966);
xor UO_2283 (O_2283,N_19936,N_19895);
or UO_2284 (O_2284,N_19898,N_19901);
nand UO_2285 (O_2285,N_19899,N_19943);
or UO_2286 (O_2286,N_19846,N_19896);
nand UO_2287 (O_2287,N_19916,N_19997);
or UO_2288 (O_2288,N_19856,N_19915);
nand UO_2289 (O_2289,N_19977,N_19851);
nand UO_2290 (O_2290,N_19874,N_19961);
nor UO_2291 (O_2291,N_19921,N_19904);
xor UO_2292 (O_2292,N_19997,N_19859);
nor UO_2293 (O_2293,N_19869,N_19959);
nand UO_2294 (O_2294,N_19889,N_19998);
and UO_2295 (O_2295,N_19969,N_19970);
or UO_2296 (O_2296,N_19912,N_19891);
and UO_2297 (O_2297,N_19973,N_19907);
xor UO_2298 (O_2298,N_19909,N_19964);
and UO_2299 (O_2299,N_19910,N_19891);
nand UO_2300 (O_2300,N_19954,N_19916);
or UO_2301 (O_2301,N_19991,N_19872);
or UO_2302 (O_2302,N_19860,N_19930);
nand UO_2303 (O_2303,N_19844,N_19843);
and UO_2304 (O_2304,N_19869,N_19967);
and UO_2305 (O_2305,N_19992,N_19960);
xnor UO_2306 (O_2306,N_19877,N_19970);
or UO_2307 (O_2307,N_19964,N_19866);
xnor UO_2308 (O_2308,N_19874,N_19957);
nor UO_2309 (O_2309,N_19992,N_19929);
xnor UO_2310 (O_2310,N_19908,N_19936);
or UO_2311 (O_2311,N_19900,N_19906);
nand UO_2312 (O_2312,N_19994,N_19904);
nand UO_2313 (O_2313,N_19954,N_19861);
xnor UO_2314 (O_2314,N_19924,N_19969);
nor UO_2315 (O_2315,N_19930,N_19878);
and UO_2316 (O_2316,N_19846,N_19905);
xor UO_2317 (O_2317,N_19849,N_19921);
or UO_2318 (O_2318,N_19904,N_19907);
or UO_2319 (O_2319,N_19864,N_19905);
xor UO_2320 (O_2320,N_19874,N_19972);
nor UO_2321 (O_2321,N_19878,N_19997);
and UO_2322 (O_2322,N_19866,N_19931);
or UO_2323 (O_2323,N_19848,N_19891);
and UO_2324 (O_2324,N_19954,N_19899);
nor UO_2325 (O_2325,N_19977,N_19887);
and UO_2326 (O_2326,N_19984,N_19840);
and UO_2327 (O_2327,N_19878,N_19908);
and UO_2328 (O_2328,N_19846,N_19993);
nor UO_2329 (O_2329,N_19870,N_19853);
and UO_2330 (O_2330,N_19853,N_19965);
nand UO_2331 (O_2331,N_19918,N_19984);
nor UO_2332 (O_2332,N_19988,N_19863);
and UO_2333 (O_2333,N_19894,N_19840);
or UO_2334 (O_2334,N_19885,N_19977);
xnor UO_2335 (O_2335,N_19861,N_19875);
nand UO_2336 (O_2336,N_19907,N_19929);
and UO_2337 (O_2337,N_19941,N_19864);
nand UO_2338 (O_2338,N_19985,N_19955);
and UO_2339 (O_2339,N_19853,N_19976);
and UO_2340 (O_2340,N_19921,N_19879);
nor UO_2341 (O_2341,N_19995,N_19894);
nand UO_2342 (O_2342,N_19995,N_19941);
nor UO_2343 (O_2343,N_19973,N_19963);
nor UO_2344 (O_2344,N_19880,N_19860);
or UO_2345 (O_2345,N_19975,N_19840);
or UO_2346 (O_2346,N_19967,N_19956);
and UO_2347 (O_2347,N_19959,N_19982);
nor UO_2348 (O_2348,N_19982,N_19846);
xor UO_2349 (O_2349,N_19933,N_19901);
and UO_2350 (O_2350,N_19896,N_19865);
nand UO_2351 (O_2351,N_19891,N_19851);
and UO_2352 (O_2352,N_19902,N_19986);
or UO_2353 (O_2353,N_19878,N_19903);
and UO_2354 (O_2354,N_19928,N_19959);
nand UO_2355 (O_2355,N_19842,N_19889);
and UO_2356 (O_2356,N_19952,N_19964);
nor UO_2357 (O_2357,N_19931,N_19962);
or UO_2358 (O_2358,N_19867,N_19849);
xor UO_2359 (O_2359,N_19869,N_19960);
xor UO_2360 (O_2360,N_19997,N_19841);
nand UO_2361 (O_2361,N_19964,N_19916);
and UO_2362 (O_2362,N_19972,N_19941);
and UO_2363 (O_2363,N_19914,N_19970);
xor UO_2364 (O_2364,N_19843,N_19922);
or UO_2365 (O_2365,N_19925,N_19845);
xnor UO_2366 (O_2366,N_19926,N_19965);
nand UO_2367 (O_2367,N_19873,N_19984);
nand UO_2368 (O_2368,N_19884,N_19865);
nor UO_2369 (O_2369,N_19981,N_19939);
nor UO_2370 (O_2370,N_19895,N_19879);
and UO_2371 (O_2371,N_19984,N_19842);
nor UO_2372 (O_2372,N_19923,N_19891);
and UO_2373 (O_2373,N_19880,N_19919);
and UO_2374 (O_2374,N_19943,N_19911);
nor UO_2375 (O_2375,N_19942,N_19908);
nand UO_2376 (O_2376,N_19921,N_19944);
nand UO_2377 (O_2377,N_19978,N_19842);
or UO_2378 (O_2378,N_19854,N_19963);
nor UO_2379 (O_2379,N_19910,N_19906);
xor UO_2380 (O_2380,N_19871,N_19994);
and UO_2381 (O_2381,N_19995,N_19843);
or UO_2382 (O_2382,N_19953,N_19949);
nor UO_2383 (O_2383,N_19894,N_19949);
nor UO_2384 (O_2384,N_19842,N_19941);
nand UO_2385 (O_2385,N_19964,N_19973);
nor UO_2386 (O_2386,N_19909,N_19944);
xor UO_2387 (O_2387,N_19957,N_19881);
xor UO_2388 (O_2388,N_19944,N_19866);
nor UO_2389 (O_2389,N_19930,N_19877);
and UO_2390 (O_2390,N_19950,N_19967);
and UO_2391 (O_2391,N_19931,N_19911);
nand UO_2392 (O_2392,N_19856,N_19846);
nand UO_2393 (O_2393,N_19950,N_19958);
or UO_2394 (O_2394,N_19994,N_19981);
nor UO_2395 (O_2395,N_19875,N_19867);
or UO_2396 (O_2396,N_19946,N_19941);
xnor UO_2397 (O_2397,N_19985,N_19844);
nor UO_2398 (O_2398,N_19970,N_19859);
or UO_2399 (O_2399,N_19965,N_19942);
xnor UO_2400 (O_2400,N_19868,N_19992);
xnor UO_2401 (O_2401,N_19926,N_19856);
or UO_2402 (O_2402,N_19953,N_19902);
and UO_2403 (O_2403,N_19962,N_19906);
xnor UO_2404 (O_2404,N_19863,N_19841);
and UO_2405 (O_2405,N_19999,N_19994);
xor UO_2406 (O_2406,N_19900,N_19883);
nor UO_2407 (O_2407,N_19905,N_19908);
xnor UO_2408 (O_2408,N_19956,N_19926);
or UO_2409 (O_2409,N_19951,N_19961);
xor UO_2410 (O_2410,N_19904,N_19890);
xor UO_2411 (O_2411,N_19869,N_19942);
nor UO_2412 (O_2412,N_19874,N_19982);
or UO_2413 (O_2413,N_19889,N_19911);
nor UO_2414 (O_2414,N_19999,N_19976);
or UO_2415 (O_2415,N_19854,N_19920);
nor UO_2416 (O_2416,N_19842,N_19928);
xor UO_2417 (O_2417,N_19871,N_19931);
or UO_2418 (O_2418,N_19998,N_19918);
and UO_2419 (O_2419,N_19906,N_19876);
and UO_2420 (O_2420,N_19984,N_19878);
or UO_2421 (O_2421,N_19858,N_19942);
nor UO_2422 (O_2422,N_19983,N_19903);
nor UO_2423 (O_2423,N_19965,N_19900);
nor UO_2424 (O_2424,N_19919,N_19994);
nand UO_2425 (O_2425,N_19991,N_19971);
xor UO_2426 (O_2426,N_19983,N_19913);
xor UO_2427 (O_2427,N_19884,N_19920);
nand UO_2428 (O_2428,N_19937,N_19864);
nor UO_2429 (O_2429,N_19994,N_19952);
nand UO_2430 (O_2430,N_19943,N_19937);
nand UO_2431 (O_2431,N_19856,N_19978);
and UO_2432 (O_2432,N_19853,N_19948);
xor UO_2433 (O_2433,N_19882,N_19840);
nor UO_2434 (O_2434,N_19992,N_19866);
or UO_2435 (O_2435,N_19872,N_19955);
or UO_2436 (O_2436,N_19849,N_19944);
nand UO_2437 (O_2437,N_19956,N_19975);
xnor UO_2438 (O_2438,N_19918,N_19849);
xnor UO_2439 (O_2439,N_19904,N_19911);
and UO_2440 (O_2440,N_19859,N_19903);
nor UO_2441 (O_2441,N_19855,N_19915);
xnor UO_2442 (O_2442,N_19882,N_19974);
nand UO_2443 (O_2443,N_19953,N_19898);
or UO_2444 (O_2444,N_19994,N_19924);
xor UO_2445 (O_2445,N_19953,N_19912);
xnor UO_2446 (O_2446,N_19886,N_19864);
or UO_2447 (O_2447,N_19865,N_19858);
or UO_2448 (O_2448,N_19949,N_19843);
nand UO_2449 (O_2449,N_19845,N_19902);
or UO_2450 (O_2450,N_19866,N_19942);
xnor UO_2451 (O_2451,N_19994,N_19931);
or UO_2452 (O_2452,N_19930,N_19864);
nor UO_2453 (O_2453,N_19967,N_19931);
and UO_2454 (O_2454,N_19958,N_19897);
and UO_2455 (O_2455,N_19968,N_19874);
nor UO_2456 (O_2456,N_19937,N_19865);
xnor UO_2457 (O_2457,N_19876,N_19882);
or UO_2458 (O_2458,N_19923,N_19911);
xor UO_2459 (O_2459,N_19851,N_19992);
and UO_2460 (O_2460,N_19955,N_19908);
xor UO_2461 (O_2461,N_19984,N_19945);
nand UO_2462 (O_2462,N_19841,N_19876);
nor UO_2463 (O_2463,N_19923,N_19877);
and UO_2464 (O_2464,N_19999,N_19907);
xor UO_2465 (O_2465,N_19958,N_19902);
and UO_2466 (O_2466,N_19985,N_19979);
and UO_2467 (O_2467,N_19939,N_19919);
nand UO_2468 (O_2468,N_19990,N_19927);
or UO_2469 (O_2469,N_19881,N_19899);
nor UO_2470 (O_2470,N_19956,N_19878);
nand UO_2471 (O_2471,N_19862,N_19854);
or UO_2472 (O_2472,N_19915,N_19960);
xnor UO_2473 (O_2473,N_19869,N_19936);
and UO_2474 (O_2474,N_19977,N_19947);
nand UO_2475 (O_2475,N_19958,N_19906);
xor UO_2476 (O_2476,N_19974,N_19938);
xor UO_2477 (O_2477,N_19986,N_19870);
nand UO_2478 (O_2478,N_19916,N_19944);
nand UO_2479 (O_2479,N_19843,N_19857);
nand UO_2480 (O_2480,N_19942,N_19847);
nand UO_2481 (O_2481,N_19918,N_19935);
nor UO_2482 (O_2482,N_19988,N_19927);
nand UO_2483 (O_2483,N_19952,N_19908);
or UO_2484 (O_2484,N_19890,N_19876);
and UO_2485 (O_2485,N_19875,N_19925);
nand UO_2486 (O_2486,N_19852,N_19867);
xnor UO_2487 (O_2487,N_19977,N_19922);
or UO_2488 (O_2488,N_19922,N_19958);
nand UO_2489 (O_2489,N_19892,N_19975);
nand UO_2490 (O_2490,N_19924,N_19923);
and UO_2491 (O_2491,N_19841,N_19908);
or UO_2492 (O_2492,N_19995,N_19939);
nor UO_2493 (O_2493,N_19914,N_19867);
or UO_2494 (O_2494,N_19848,N_19845);
and UO_2495 (O_2495,N_19965,N_19842);
nand UO_2496 (O_2496,N_19981,N_19884);
xnor UO_2497 (O_2497,N_19961,N_19954);
xor UO_2498 (O_2498,N_19897,N_19874);
xnor UO_2499 (O_2499,N_19856,N_19945);
endmodule