module basic_2500_25000_3000_20_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_755,In_2201);
xor U1 (N_1,In_1071,In_1011);
xor U2 (N_2,In_1974,In_2380);
xor U3 (N_3,In_187,In_1704);
nor U4 (N_4,In_986,In_2325);
and U5 (N_5,In_573,In_1492);
or U6 (N_6,In_183,In_1920);
xor U7 (N_7,In_1989,In_112);
nand U8 (N_8,In_884,In_1389);
or U9 (N_9,In_2357,In_1568);
nor U10 (N_10,In_366,In_338);
xnor U11 (N_11,In_1225,In_2081);
xnor U12 (N_12,In_1404,In_423);
nand U13 (N_13,In_2249,In_199);
nand U14 (N_14,In_135,In_1136);
xnor U15 (N_15,In_632,In_1713);
xnor U16 (N_16,In_2389,In_2328);
nand U17 (N_17,In_1447,In_1841);
nor U18 (N_18,In_335,In_2332);
and U19 (N_19,In_358,In_1517);
and U20 (N_20,In_470,In_2075);
and U21 (N_21,In_491,In_16);
xor U22 (N_22,In_1628,In_1432);
and U23 (N_23,In_1045,In_203);
nor U24 (N_24,In_98,In_1294);
nand U25 (N_25,In_1824,In_1097);
nor U26 (N_26,In_1852,In_1388);
nand U27 (N_27,In_1394,In_1348);
nand U28 (N_28,In_2442,In_1602);
nor U29 (N_29,In_1134,In_1816);
and U30 (N_30,In_118,In_416);
xnor U31 (N_31,In_1689,In_2352);
and U32 (N_32,In_608,In_718);
nor U33 (N_33,In_1622,In_723);
xnor U34 (N_34,In_62,In_2436);
xnor U35 (N_35,In_1399,In_2018);
or U36 (N_36,In_933,In_61);
nor U37 (N_37,In_1060,In_2388);
xor U38 (N_38,In_294,In_209);
and U39 (N_39,In_2405,In_2205);
nand U40 (N_40,In_984,In_2029);
nand U41 (N_41,In_1983,In_1112);
or U42 (N_42,In_1257,In_1355);
nand U43 (N_43,In_2354,In_328);
xnor U44 (N_44,In_1769,In_2307);
and U45 (N_45,In_2045,In_2023);
nand U46 (N_46,In_2272,In_545);
nor U47 (N_47,In_259,In_529);
or U48 (N_48,In_891,In_288);
nor U49 (N_49,In_78,In_805);
or U50 (N_50,In_461,In_300);
and U51 (N_51,In_1712,In_1169);
or U52 (N_52,In_1352,In_652);
and U53 (N_53,In_524,In_269);
or U54 (N_54,In_2225,In_1125);
xnor U55 (N_55,In_57,In_1898);
nand U56 (N_56,In_541,In_1793);
xor U57 (N_57,In_830,In_694);
or U58 (N_58,In_872,In_1349);
nand U59 (N_59,In_1849,In_1900);
xnor U60 (N_60,In_2052,In_1213);
and U61 (N_61,In_111,In_854);
and U62 (N_62,In_1444,In_838);
nand U63 (N_63,In_1838,In_794);
xnor U64 (N_64,In_782,In_296);
xor U65 (N_65,In_665,In_397);
and U66 (N_66,In_858,In_1066);
or U67 (N_67,In_2217,In_1981);
xnor U68 (N_68,In_2320,In_720);
nand U69 (N_69,In_2243,In_954);
or U70 (N_70,In_1437,In_932);
nand U71 (N_71,In_2266,In_2251);
xor U72 (N_72,In_2410,In_1552);
nand U73 (N_73,In_1637,In_522);
nor U74 (N_74,In_121,In_584);
xnor U75 (N_75,In_173,In_152);
or U76 (N_76,In_433,In_389);
nand U77 (N_77,In_407,In_1907);
xnor U78 (N_78,In_2024,In_156);
xor U79 (N_79,In_721,In_907);
xnor U80 (N_80,In_1,In_1839);
and U81 (N_81,In_1113,In_474);
nor U82 (N_82,In_1052,In_2093);
nand U83 (N_83,In_2284,In_2079);
or U84 (N_84,In_1048,In_88);
nor U85 (N_85,In_2413,In_19);
or U86 (N_86,In_866,In_251);
xor U87 (N_87,In_1947,In_1980);
xor U88 (N_88,In_1668,In_310);
and U89 (N_89,In_1328,In_52);
nand U90 (N_90,In_1187,In_644);
or U91 (N_91,In_1290,In_1534);
nand U92 (N_92,In_1670,In_509);
xor U93 (N_93,In_946,In_1175);
nor U94 (N_94,In_427,In_55);
nand U95 (N_95,In_309,In_2438);
xnor U96 (N_96,In_717,In_2126);
and U97 (N_97,In_2398,In_768);
nor U98 (N_98,In_1227,In_117);
xor U99 (N_99,In_446,In_1876);
and U100 (N_100,In_816,In_798);
or U101 (N_101,In_765,In_2250);
nor U102 (N_102,In_2309,In_1716);
nand U103 (N_103,In_961,In_581);
or U104 (N_104,In_1992,In_1724);
xor U105 (N_105,In_886,In_589);
nand U106 (N_106,In_297,In_2115);
and U107 (N_107,In_2055,In_323);
and U108 (N_108,In_1463,In_32);
and U109 (N_109,In_2037,In_33);
xnor U110 (N_110,In_2064,In_2431);
and U111 (N_111,In_1997,In_1240);
nand U112 (N_112,In_85,In_651);
and U113 (N_113,In_204,In_2375);
xnor U114 (N_114,In_20,In_1829);
and U115 (N_115,In_669,In_1660);
and U116 (N_116,In_1267,In_1197);
nor U117 (N_117,In_2254,In_0);
xnor U118 (N_118,In_662,In_2218);
nor U119 (N_119,In_2020,In_2222);
xor U120 (N_120,In_585,In_218);
nand U121 (N_121,In_526,In_21);
nor U122 (N_122,In_2103,In_2187);
nand U123 (N_123,In_2348,In_2206);
nor U124 (N_124,In_2471,In_686);
and U125 (N_125,In_1596,In_1206);
or U126 (N_126,In_1319,In_1555);
or U127 (N_127,In_1528,In_1218);
or U128 (N_128,In_2042,In_1832);
xnor U129 (N_129,In_527,In_1866);
nand U130 (N_130,In_1597,In_1697);
or U131 (N_131,In_1135,In_992);
or U132 (N_132,In_708,In_1371);
nor U133 (N_133,In_1666,In_658);
nor U134 (N_134,In_2152,In_2276);
nor U135 (N_135,In_1033,In_1254);
or U136 (N_136,In_2083,In_1952);
xnor U137 (N_137,In_284,In_844);
nor U138 (N_138,In_908,In_690);
xnor U139 (N_139,In_136,In_466);
or U140 (N_140,In_1152,In_1093);
nor U141 (N_141,In_46,In_1853);
and U142 (N_142,In_1021,In_1835);
nor U143 (N_143,In_177,In_1721);
xnor U144 (N_144,In_889,In_2495);
nor U145 (N_145,In_2032,In_2453);
nor U146 (N_146,In_1305,In_1657);
xor U147 (N_147,In_1344,In_1639);
and U148 (N_148,In_2232,In_2401);
or U149 (N_149,In_2128,In_508);
nand U150 (N_150,In_155,In_1655);
nand U151 (N_151,In_1128,In_372);
xor U152 (N_152,In_2148,In_1896);
xnor U153 (N_153,In_1456,In_2268);
or U154 (N_154,In_459,In_894);
and U155 (N_155,In_2017,In_732);
nand U156 (N_156,In_878,In_941);
or U157 (N_157,In_1058,In_770);
and U158 (N_158,In_2224,In_197);
or U159 (N_159,In_50,In_2228);
nand U160 (N_160,In_1837,In_518);
or U161 (N_161,In_1902,In_370);
nand U162 (N_162,In_36,In_2382);
nand U163 (N_163,In_948,In_406);
and U164 (N_164,In_1229,In_2434);
nor U165 (N_165,In_863,In_641);
and U166 (N_166,In_2487,In_1424);
nand U167 (N_167,In_1467,In_1300);
nand U168 (N_168,In_1585,In_914);
nand U169 (N_169,In_639,In_1910);
and U170 (N_170,In_917,In_1111);
xor U171 (N_171,In_1559,In_1260);
nor U172 (N_172,In_1893,In_591);
nor U173 (N_173,In_724,In_702);
nand U174 (N_174,In_1787,In_523);
xnor U175 (N_175,In_1268,In_1583);
xnor U176 (N_176,In_521,In_54);
nand U177 (N_177,In_481,In_1809);
xnor U178 (N_178,In_2488,In_243);
and U179 (N_179,In_647,In_1198);
nand U180 (N_180,In_83,In_35);
nand U181 (N_181,In_745,In_711);
xnor U182 (N_182,In_555,In_63);
and U183 (N_183,In_701,In_1730);
xnor U184 (N_184,In_2233,In_2193);
xor U185 (N_185,In_1669,In_1353);
and U186 (N_186,In_1828,In_1358);
or U187 (N_187,In_1193,In_376);
and U188 (N_188,In_2447,In_1524);
nor U189 (N_189,In_354,In_2392);
nand U190 (N_190,In_1369,In_1548);
and U191 (N_191,In_1711,In_1422);
or U192 (N_192,In_493,In_1798);
nand U193 (N_193,In_2263,In_68);
nor U194 (N_194,In_1745,In_1376);
xor U195 (N_195,In_1298,In_1626);
xor U196 (N_196,In_1959,In_2166);
nor U197 (N_197,In_772,In_1101);
and U198 (N_198,In_2097,In_139);
nor U199 (N_199,In_657,In_1970);
and U200 (N_200,In_2489,In_713);
nand U201 (N_201,In_1004,In_2144);
nor U202 (N_202,In_549,In_1029);
nand U203 (N_203,In_1256,In_1943);
nand U204 (N_204,In_983,In_803);
xor U205 (N_205,In_1529,In_217);
nand U206 (N_206,In_1120,In_249);
nor U207 (N_207,In_725,In_248);
xnor U208 (N_208,In_2101,In_1149);
nand U209 (N_209,In_1690,In_1768);
or U210 (N_210,In_1307,In_1374);
or U211 (N_211,In_1095,In_2199);
nor U212 (N_212,In_993,In_229);
or U213 (N_213,In_2383,In_237);
xor U214 (N_214,In_2008,In_2295);
nand U215 (N_215,In_1204,In_1917);
nor U216 (N_216,In_2429,In_1402);
xnor U217 (N_217,In_1860,In_1221);
nand U218 (N_218,In_390,In_2421);
or U219 (N_219,In_1428,In_421);
xnor U220 (N_220,In_1379,In_937);
nor U221 (N_221,In_1522,In_51);
or U222 (N_222,In_377,In_222);
nand U223 (N_223,In_1926,In_314);
nand U224 (N_224,In_113,In_1776);
xnor U225 (N_225,In_4,In_2226);
and U226 (N_226,In_1693,In_326);
or U227 (N_227,In_385,In_2370);
nand U228 (N_228,In_1919,In_103);
nor U229 (N_229,In_257,In_2304);
nand U230 (N_230,In_2446,In_159);
and U231 (N_231,In_2270,In_90);
nor U232 (N_232,In_1698,In_2149);
nand U233 (N_233,In_679,In_2204);
nor U234 (N_234,In_42,In_538);
nand U235 (N_235,In_185,In_210);
and U236 (N_236,In_1117,In_1887);
nor U237 (N_237,In_2203,In_1990);
nor U238 (N_238,In_629,In_1347);
nor U239 (N_239,In_469,In_434);
and U240 (N_240,In_1251,In_2430);
nand U241 (N_241,In_2078,In_342);
nor U242 (N_242,In_81,In_892);
xnor U243 (N_243,In_1754,In_1479);
or U244 (N_244,In_1214,In_213);
and U245 (N_245,In_419,In_733);
nor U246 (N_246,In_1948,In_1792);
xnor U247 (N_247,In_640,In_1975);
and U248 (N_248,In_654,In_2001);
nand U249 (N_249,In_1874,In_264);
or U250 (N_250,In_211,In_1069);
xor U251 (N_251,In_120,In_2086);
nor U252 (N_252,In_2486,In_2132);
nor U253 (N_253,In_1400,In_1162);
xor U254 (N_254,In_938,In_618);
and U255 (N_255,In_2458,In_1387);
nand U256 (N_256,In_1936,In_2113);
nor U257 (N_257,In_164,In_308);
xnor U258 (N_258,In_1427,In_186);
or U259 (N_259,In_175,In_749);
or U260 (N_260,In_767,In_2036);
nand U261 (N_261,In_56,In_2192);
or U262 (N_262,In_356,In_2242);
nand U263 (N_263,In_2331,In_1501);
and U264 (N_264,In_1734,In_623);
and U265 (N_265,In_494,In_1827);
xnor U266 (N_266,In_1966,In_1130);
or U267 (N_267,In_600,In_1889);
and U268 (N_268,In_303,In_2402);
or U269 (N_269,In_1053,In_1965);
or U270 (N_270,In_40,In_448);
nor U271 (N_271,In_696,In_347);
or U272 (N_272,In_1336,In_754);
nand U273 (N_273,In_1085,In_769);
nand U274 (N_274,In_1018,In_375);
or U275 (N_275,In_329,In_2316);
xor U276 (N_276,In_599,In_2355);
and U277 (N_277,In_388,In_311);
and U278 (N_278,In_773,In_1744);
xor U279 (N_279,In_1497,In_2175);
and U280 (N_280,In_1265,In_1370);
or U281 (N_281,In_1846,In_2259);
nand U282 (N_282,In_633,In_1449);
xnor U283 (N_283,In_1418,In_1679);
nor U284 (N_284,In_265,In_2028);
and U285 (N_285,In_2283,In_1067);
nand U286 (N_286,In_622,In_1315);
and U287 (N_287,In_1001,In_2255);
nor U288 (N_288,In_2109,In_1147);
or U289 (N_289,In_2424,In_1211);
and U290 (N_290,In_806,In_671);
xor U291 (N_291,In_25,In_625);
nand U292 (N_292,In_715,In_1040);
and U293 (N_293,In_1865,In_2484);
nor U294 (N_294,In_1132,In_1024);
or U295 (N_295,In_661,In_254);
and U296 (N_296,In_2027,In_2450);
xnor U297 (N_297,In_1145,In_2121);
and U298 (N_298,In_2176,In_1831);
or U299 (N_299,In_402,In_1331);
or U300 (N_300,In_305,In_1115);
xnor U301 (N_301,In_1180,In_980);
and U302 (N_302,In_2245,In_1244);
nand U303 (N_303,In_1142,In_401);
and U304 (N_304,In_1223,In_1318);
nor U305 (N_305,In_1034,In_2296);
and U306 (N_306,In_1703,In_190);
nor U307 (N_307,In_2303,In_543);
and U308 (N_308,In_1278,In_1963);
or U309 (N_309,In_74,In_1423);
nand U310 (N_310,In_450,In_1238);
nor U311 (N_311,In_2427,In_2168);
nor U312 (N_312,In_2312,In_510);
nor U313 (N_313,In_2444,In_148);
or U314 (N_314,In_1789,In_1141);
and U315 (N_315,In_1114,In_59);
nor U316 (N_316,In_2007,In_1167);
nor U317 (N_317,In_2321,In_565);
and U318 (N_318,In_1311,In_2124);
and U319 (N_319,In_2170,In_1766);
xnor U320 (N_320,In_444,In_322);
or U321 (N_321,In_276,In_1633);
nand U322 (N_322,In_399,In_1280);
xor U323 (N_323,In_238,In_998);
nand U324 (N_324,In_2441,In_18);
or U325 (N_325,In_2318,In_1873);
xor U326 (N_326,In_1378,In_1202);
nor U327 (N_327,In_2319,In_1143);
nand U328 (N_328,In_2033,In_2433);
nor U329 (N_329,In_1102,In_1446);
nor U330 (N_330,In_77,In_557);
and U331 (N_331,In_691,In_438);
nand U332 (N_332,In_1028,In_2369);
and U333 (N_333,In_1195,In_1421);
or U334 (N_334,In_71,In_1511);
and U335 (N_335,In_987,In_743);
xnor U336 (N_336,In_1411,In_783);
xor U337 (N_337,In_2492,In_1475);
xnor U338 (N_338,In_1623,In_487);
xor U339 (N_339,In_28,In_53);
nand U340 (N_340,In_2305,In_2147);
or U341 (N_341,In_286,In_2237);
or U342 (N_342,In_64,In_344);
and U343 (N_343,In_1050,In_2183);
xnor U344 (N_344,In_605,In_31);
and U345 (N_345,In_813,In_1490);
nand U346 (N_346,In_412,In_915);
nor U347 (N_347,In_2143,In_531);
or U348 (N_348,In_1881,In_1473);
and U349 (N_349,In_533,In_682);
nor U350 (N_350,In_1042,In_1857);
or U351 (N_351,In_1561,In_823);
xnor U352 (N_352,In_1801,In_2374);
nand U353 (N_353,In_1715,In_1850);
nand U354 (N_354,In_2072,In_1087);
nor U355 (N_355,In_1954,In_2065);
xnor U356 (N_356,In_2476,In_1855);
or U357 (N_357,In_200,In_1314);
or U358 (N_358,In_1957,In_2000);
nor U359 (N_359,In_839,In_734);
or U360 (N_360,In_539,In_2269);
nor U361 (N_361,In_567,In_2498);
or U362 (N_362,In_1151,In_1357);
nor U363 (N_363,In_989,In_1398);
xor U364 (N_364,In_664,In_266);
nand U365 (N_365,In_1738,In_680);
nor U366 (N_366,In_1656,In_1939);
or U367 (N_367,In_579,In_1580);
xnor U368 (N_368,In_1185,In_964);
xnor U369 (N_369,In_2396,In_1468);
and U370 (N_370,In_105,In_1620);
xor U371 (N_371,In_1638,In_2173);
or U372 (N_372,In_2479,In_437);
and U373 (N_373,In_1591,In_666);
nand U374 (N_374,In_1338,In_764);
xnor U375 (N_375,In_2063,In_799);
nor U376 (N_376,In_351,In_1410);
nor U377 (N_377,In_1658,In_221);
nand U378 (N_378,In_1796,In_2098);
or U379 (N_379,In_1210,In_748);
and U380 (N_380,In_263,In_2418);
and U381 (N_381,In_2356,In_1505);
or U382 (N_382,In_472,In_2404);
xnor U383 (N_383,In_1217,In_2046);
xnor U384 (N_384,In_1822,In_157);
xnor U385 (N_385,In_1726,In_1036);
nand U386 (N_386,In_1600,In_1764);
and U387 (N_387,In_1535,In_1283);
or U388 (N_388,In_876,In_890);
or U389 (N_389,In_2297,In_610);
and U390 (N_390,In_2131,In_228);
nor U391 (N_391,In_1263,In_422);
nand U392 (N_392,In_2493,In_84);
or U393 (N_393,In_179,In_1106);
xor U394 (N_394,In_140,In_706);
nor U395 (N_395,In_410,In_1804);
nand U396 (N_396,In_325,In_1171);
or U397 (N_397,In_693,In_1779);
and U398 (N_398,In_1373,In_86);
nor U399 (N_399,In_1784,In_1527);
or U400 (N_400,In_2049,In_975);
nor U401 (N_401,In_239,In_498);
nor U402 (N_402,In_909,In_1105);
nor U403 (N_403,In_994,In_536);
nand U404 (N_404,In_1870,In_1599);
and U405 (N_405,In_1150,In_598);
nor U406 (N_406,In_2394,In_489);
nand U407 (N_407,In_988,In_879);
or U408 (N_408,In_1761,In_642);
xnor U409 (N_409,In_1339,In_1138);
nand U410 (N_410,In_405,In_781);
and U411 (N_411,In_1714,In_1380);
nor U412 (N_412,In_1709,In_275);
or U413 (N_413,In_2080,In_277);
nor U414 (N_414,In_2011,In_1790);
xor U415 (N_415,In_1567,In_821);
nand U416 (N_416,In_1047,In_1691);
xnor U417 (N_417,In_2308,In_233);
nor U418 (N_418,In_1196,In_575);
nand U419 (N_419,In_1993,In_1124);
or U420 (N_420,In_345,In_2373);
xnor U421 (N_421,In_2084,In_898);
nor U422 (N_422,In_638,In_1645);
and U423 (N_423,In_1820,In_1474);
or U424 (N_424,In_674,In_426);
or U425 (N_425,In_1718,In_1208);
nand U426 (N_426,In_1160,In_1063);
nand U427 (N_427,In_171,In_513);
xnor U428 (N_428,In_471,In_2422);
nor U429 (N_429,In_1081,In_1946);
nand U430 (N_430,In_802,In_1316);
nand U431 (N_431,In_2179,In_1692);
xor U432 (N_432,In_1562,In_1652);
and U433 (N_433,In_252,In_1867);
nor U434 (N_434,In_2219,In_2136);
and U435 (N_435,In_343,In_2169);
or U436 (N_436,In_1587,In_2091);
and U437 (N_437,In_1799,In_271);
nand U438 (N_438,In_1253,In_2230);
xnor U439 (N_439,In_227,In_1560);
and U440 (N_440,In_283,In_587);
nor U441 (N_441,In_1878,In_181);
nor U442 (N_442,In_2477,In_1273);
nand U443 (N_443,In_712,In_2013);
nor U444 (N_444,In_528,In_386);
nand U445 (N_445,In_1191,In_1930);
or U446 (N_446,In_2088,In_1519);
and U447 (N_447,In_958,In_899);
or U448 (N_448,In_1888,In_2194);
or U449 (N_449,In_1488,In_867);
or U450 (N_450,In_2129,In_2288);
nand U451 (N_451,In_2376,In_1771);
or U452 (N_452,In_492,In_468);
nand U453 (N_453,In_235,In_241);
nor U454 (N_454,In_594,In_1671);
nand U455 (N_455,In_726,In_2196);
nand U456 (N_456,In_1005,In_48);
nand U457 (N_457,In_663,In_999);
xor U458 (N_458,In_604,In_2390);
and U459 (N_459,In_668,In_1297);
nand U460 (N_460,In_815,In_89);
xnor U461 (N_461,In_1295,In_1436);
and U462 (N_462,In_2393,In_1220);
nand U463 (N_463,In_1003,In_1875);
xnor U464 (N_464,In_593,In_1755);
or U465 (N_465,In_947,In_1434);
or U466 (N_466,In_168,In_2154);
xor U467 (N_467,In_260,In_93);
xnor U468 (N_468,In_1588,In_381);
nor U469 (N_469,In_66,In_2289);
nor U470 (N_470,In_2151,In_1306);
nand U471 (N_471,In_2239,In_1250);
nand U472 (N_472,In_147,In_929);
and U473 (N_473,In_1359,In_1817);
nor U474 (N_474,In_127,In_562);
and U475 (N_475,In_2483,In_1915);
or U476 (N_476,In_396,In_506);
or U477 (N_477,In_2053,In_1186);
and U478 (N_478,In_2293,In_1430);
xor U479 (N_479,In_2435,In_104);
xnor U480 (N_480,In_1055,In_2473);
or U481 (N_481,In_1694,In_110);
xnor U482 (N_482,In_670,In_626);
nor U483 (N_483,In_612,In_842);
and U484 (N_484,In_1409,In_1531);
nand U485 (N_485,In_570,In_1025);
or U486 (N_486,In_1812,In_1759);
and U487 (N_487,In_801,In_182);
or U488 (N_488,In_1116,In_2158);
xor U489 (N_489,In_307,In_900);
and U490 (N_490,In_2366,In_158);
xnor U491 (N_491,In_1624,In_1163);
xor U492 (N_492,In_960,In_819);
xnor U493 (N_493,In_590,In_1261);
or U494 (N_494,In_2469,In_223);
nor U495 (N_495,In_2207,In_1343);
or U496 (N_496,In_2457,In_2253);
xnor U497 (N_497,In_548,In_2365);
nor U498 (N_498,In_476,In_1921);
or U499 (N_499,In_480,In_2344);
nor U500 (N_500,In_201,In_1617);
nor U501 (N_501,In_775,In_41);
and U502 (N_502,In_371,In_8);
nor U503 (N_503,In_888,In_2215);
and U504 (N_504,In_2360,In_1413);
or U505 (N_505,In_2050,In_1987);
xor U506 (N_506,In_1131,In_2258);
nor U507 (N_507,In_1941,In_1321);
and U508 (N_508,In_2333,In_2073);
or U509 (N_509,In_2326,In_1973);
xor U510 (N_510,In_1462,In_1908);
nor U511 (N_511,In_1485,In_2439);
and U512 (N_512,In_2160,In_403);
xnor U513 (N_513,In_1431,In_47);
nor U514 (N_514,In_1012,In_970);
xnor U515 (N_515,In_1178,In_2350);
nor U516 (N_516,In_1678,In_1582);
nand U517 (N_517,In_785,In_2227);
nor U518 (N_518,In_1397,In_571);
and U519 (N_519,In_580,In_1612);
nand U520 (N_520,In_1442,In_1070);
and U521 (N_521,In_1818,In_1493);
xor U522 (N_522,In_1303,In_1451);
xor U523 (N_523,In_1584,In_1453);
xnor U524 (N_524,In_272,In_128);
and U525 (N_525,In_162,In_26);
nor U526 (N_526,In_1086,In_2462);
or U527 (N_527,In_788,In_2116);
and U528 (N_528,In_699,In_2286);
nor U529 (N_529,In_192,In_484);
xnor U530 (N_530,In_1457,In_1884);
nor U531 (N_531,In_337,In_2403);
nor U532 (N_532,In_2087,In_1203);
and U533 (N_533,In_299,In_1687);
nand U534 (N_534,In_1046,In_614);
and U535 (N_535,In_1496,In_291);
nor U536 (N_536,In_362,In_1933);
xnor U537 (N_537,In_1351,In_787);
or U538 (N_538,In_287,In_116);
xor U539 (N_539,In_2290,In_659);
or U540 (N_540,In_1982,In_912);
or U541 (N_541,In_2451,In_943);
xor U542 (N_542,In_1014,In_73);
nor U543 (N_543,In_1526,In_2047);
nand U544 (N_544,In_174,In_2464);
nand U545 (N_545,In_1372,In_1550);
or U546 (N_546,In_124,In_851);
nand U547 (N_547,In_451,In_2130);
and U548 (N_548,In_80,In_2138);
nand U549 (N_549,In_1075,In_1439);
nor U550 (N_550,In_1891,In_2432);
or U551 (N_551,In_312,In_2010);
and U552 (N_552,In_1076,In_1931);
nor U553 (N_553,In_2343,In_1641);
nand U554 (N_554,In_2054,In_1886);
nor U555 (N_555,In_137,In_1673);
xor U556 (N_556,In_490,In_2163);
xnor U557 (N_557,In_793,In_1932);
xor U558 (N_558,In_2127,In_2278);
and U559 (N_559,In_153,In_1458);
xor U560 (N_560,In_383,In_1464);
and U561 (N_561,In_2122,In_315);
nor U562 (N_562,In_1649,In_106);
nand U563 (N_563,In_1189,In_1883);
xor U564 (N_564,In_1084,In_1068);
and U565 (N_565,In_756,In_643);
xor U566 (N_566,In_2244,In_332);
xnor U567 (N_567,In_2395,In_1484);
nor U568 (N_568,In_411,In_577);
xnor U569 (N_569,In_1940,In_298);
xor U570 (N_570,In_617,In_2353);
and U571 (N_571,In_373,In_1767);
nand U572 (N_572,In_1181,In_2359);
nor U573 (N_573,In_1895,In_911);
nand U574 (N_574,In_1292,In_968);
nor U575 (N_575,In_2338,In_2322);
or U576 (N_576,In_951,In_2185);
and U577 (N_577,In_1914,In_2311);
and U578 (N_578,In_2211,In_790);
nor U579 (N_579,In_231,In_91);
nor U580 (N_580,In_206,In_714);
xor U581 (N_581,In_1330,In_2314);
nor U582 (N_582,In_624,In_1538);
or U583 (N_583,In_2118,In_43);
nand U584 (N_584,In_1735,In_1869);
and U585 (N_585,In_1944,In_516);
xor U586 (N_586,In_1739,In_1200);
nor U587 (N_587,In_560,In_280);
xnor U588 (N_588,In_2460,In_1770);
or U589 (N_589,In_2082,In_1700);
xnor U590 (N_590,In_393,In_1502);
nor U591 (N_591,In_752,In_1736);
nand U592 (N_592,In_2100,In_1340);
xnor U593 (N_593,In_1455,In_576);
xnor U594 (N_594,In_2188,In_1412);
or U595 (N_595,In_1038,In_301);
or U596 (N_596,In_1619,In_1890);
or U597 (N_597,In_1471,In_895);
or U598 (N_598,In_515,In_1749);
and U599 (N_599,In_1565,In_58);
xor U600 (N_600,In_2449,In_453);
xnor U601 (N_601,In_603,In_100);
and U602 (N_602,In_2461,In_1478);
nor U603 (N_603,In_475,In_544);
or U604 (N_604,In_1074,In_1104);
nor U605 (N_605,In_1871,In_2174);
nor U606 (N_606,In_1750,In_1044);
and U607 (N_607,In_2235,In_365);
and U608 (N_608,In_488,In_928);
and U609 (N_609,In_758,In_537);
xnor U610 (N_610,In_1506,In_995);
and U611 (N_611,In_1507,In_963);
xnor U612 (N_612,In_452,In_1634);
or U613 (N_613,In_1616,In_1604);
or U614 (N_614,In_1435,In_1788);
nand U615 (N_615,In_131,In_552);
nor U616 (N_616,In_67,In_2267);
or U617 (N_617,In_1958,In_1172);
or U618 (N_618,In_969,In_455);
or U619 (N_619,In_361,In_556);
and U620 (N_620,In_141,In_1897);
or U621 (N_621,In_1406,In_519);
nor U622 (N_622,In_1190,In_1284);
nand U623 (N_623,In_1333,In_1262);
nand U624 (N_624,In_2133,In_1918);
nand U625 (N_625,In_1482,In_1969);
and U626 (N_626,In_1320,In_574);
nor U627 (N_627,In_2198,In_1847);
and U628 (N_628,In_2111,In_1441);
or U629 (N_629,In_688,In_1882);
xnor U630 (N_630,In_1635,In_2134);
nor U631 (N_631,In_1368,In_729);
or U632 (N_632,In_1127,In_457);
nor U633 (N_633,In_49,In_1964);
nor U634 (N_634,In_449,In_2420);
and U635 (N_635,In_1680,In_800);
nor U636 (N_636,In_1037,In_810);
nor U637 (N_637,In_971,In_1469);
xnor U638 (N_638,In_771,In_428);
nand U639 (N_639,In_796,In_1123);
or U640 (N_640,In_2378,In_391);
nand U641 (N_641,In_1662,In_1640);
nor U642 (N_642,In_2351,In_1245);
and U643 (N_643,In_1995,In_1729);
xnor U644 (N_644,In_1650,In_936);
nand U645 (N_645,In_1934,In_1797);
or U646 (N_646,In_635,In_1756);
or U647 (N_647,In_1426,In_2110);
and U648 (N_648,In_102,In_2367);
nand U649 (N_649,In_2060,In_1312);
nand U650 (N_650,In_1059,In_333);
xnor U651 (N_651,In_2034,In_837);
or U652 (N_652,In_1016,In_2472);
xnor U653 (N_653,In_384,In_2485);
nand U654 (N_654,In_132,In_1459);
and U655 (N_655,In_1530,In_2387);
xnor U656 (N_656,In_1549,In_1168);
nand U657 (N_657,In_219,In_2299);
xnor U658 (N_658,In_678,In_525);
xor U659 (N_659,In_1248,In_1537);
nand U660 (N_660,In_1753,In_824);
nand U661 (N_661,In_507,In_226);
nand U662 (N_662,In_2212,In_447);
nand U663 (N_663,In_1062,In_505);
and U664 (N_664,In_1651,In_462);
or U665 (N_665,In_1065,In_1073);
or U666 (N_666,In_982,In_864);
nand U667 (N_667,In_2335,In_1035);
and U668 (N_668,In_939,In_1508);
nor U669 (N_669,In_1546,In_1277);
nand U670 (N_670,In_212,In_92);
nand U671 (N_671,In_1688,In_2056);
nor U672 (N_672,In_2120,In_1777);
and U673 (N_673,In_2026,In_367);
nor U674 (N_674,In_619,In_1361);
and U675 (N_675,In_27,In_2066);
or U676 (N_676,In_2273,In_101);
or U677 (N_677,In_1592,In_79);
xnor U678 (N_678,In_2292,In_1851);
xnor U679 (N_679,In_1350,In_1148);
xnor U680 (N_680,In_1392,In_2349);
nand U681 (N_681,In_1782,In_1569);
xnor U682 (N_682,In_1119,In_1705);
nor U683 (N_683,In_119,In_1270);
and U684 (N_684,In_607,In_1416);
or U685 (N_685,In_1695,In_1999);
and U686 (N_686,In_675,In_2141);
nand U687 (N_687,In_172,In_2209);
nor U688 (N_688,In_318,In_304);
xnor U689 (N_689,In_990,In_1701);
nor U690 (N_690,In_1598,In_1108);
and U691 (N_691,In_859,In_195);
or U692 (N_692,In_840,In_107);
or U693 (N_693,In_1017,In_1605);
and U694 (N_694,In_1747,In_414);
or U695 (N_695,In_1916,In_123);
and U696 (N_696,In_2415,In_334);
xnor U697 (N_697,In_2181,In_784);
and U698 (N_698,In_676,In_13);
nor U699 (N_699,In_482,In_738);
and U700 (N_700,In_1672,In_2140);
and U701 (N_701,In_1481,In_700);
and U702 (N_702,In_1722,In_2409);
nand U703 (N_703,In_1525,In_1154);
and U704 (N_704,In_2164,In_2499);
nor U705 (N_705,In_2330,In_572);
and U706 (N_706,In_1702,In_835);
xor U707 (N_707,In_1201,In_1429);
xnor U708 (N_708,In_247,In_425);
xnor U709 (N_709,In_1872,In_766);
and U710 (N_710,In_1707,In_1346);
nor U711 (N_711,In_2108,In_1231);
and U712 (N_712,In_1614,In_1541);
xnor U713 (N_713,In_2162,In_1795);
nand U714 (N_714,In_1407,In_170);
xor U715 (N_715,In_2474,In_2391);
xnor U716 (N_716,In_234,In_1664);
or U717 (N_717,In_2408,In_1654);
nand U718 (N_718,In_1781,In_1360);
xnor U719 (N_719,In_1912,In_114);
or U720 (N_720,In_704,In_2346);
and U721 (N_721,In_1762,In_282);
or U722 (N_722,In_2171,In_2167);
or U723 (N_723,In_2195,In_1232);
nand U724 (N_724,In_1991,In_534);
nor U725 (N_725,In_2038,In_2363);
and U726 (N_726,In_550,In_2155);
or U727 (N_727,In_274,In_2039);
and U728 (N_728,In_2494,In_2099);
xnor U729 (N_729,In_1674,In_1057);
xor U730 (N_730,In_1285,In_1129);
and U731 (N_731,In_2280,In_1733);
or U732 (N_732,In_578,In_1621);
nor U733 (N_733,In_1433,In_1096);
and U734 (N_734,In_1727,In_1630);
xnor U735 (N_735,In_620,In_1553);
nand U736 (N_736,In_1518,In_1625);
and U737 (N_737,In_2294,In_1786);
xor U738 (N_738,In_739,In_1979);
and U739 (N_739,In_763,In_808);
or U740 (N_740,In_760,In_149);
xnor U741 (N_741,In_1039,In_762);
xnor U742 (N_742,In_1676,In_1390);
nor U743 (N_743,In_959,In_976);
and U744 (N_744,In_250,In_1222);
and U745 (N_745,In_497,In_1483);
or U746 (N_746,In_2459,In_2190);
and U747 (N_747,In_786,In_1741);
xor U748 (N_748,In_2327,In_129);
xnor U749 (N_749,In_940,In_1532);
nand U750 (N_750,In_1825,In_279);
nor U751 (N_751,In_1234,In_1159);
nor U752 (N_752,In_2426,In_1520);
or U753 (N_753,In_2282,In_267);
xor U754 (N_754,In_1309,In_1905);
nor U755 (N_755,In_1611,In_2021);
and U756 (N_756,In_1901,In_2301);
nor U757 (N_757,In_1544,In_1334);
and U758 (N_758,In_293,In_532);
xnor U759 (N_759,In_934,In_1155);
and U760 (N_760,In_1661,In_2480);
xnor U761 (N_761,In_956,In_278);
or U762 (N_762,In_684,In_1425);
or U763 (N_763,In_1504,In_1450);
and U764 (N_764,In_1968,In_216);
nand U765 (N_765,In_978,In_981);
nand U766 (N_766,In_849,In_1571);
xnor U767 (N_767,In_456,In_1845);
nor U768 (N_768,In_1815,In_1632);
and U769 (N_769,In_1420,In_1324);
and U770 (N_770,In_1576,In_653);
nand U771 (N_771,In_1020,In_1249);
nor U772 (N_772,In_1090,In_1859);
nand U773 (N_773,In_359,In_2336);
and U774 (N_774,In_695,In_208);
and U775 (N_775,In_2260,In_825);
xnor U776 (N_776,In_747,In_1445);
and U777 (N_777,In_1819,In_804);
xor U778 (N_778,In_827,In_707);
or U779 (N_779,In_1683,In_1089);
nor U780 (N_780,In_1382,In_962);
xnor U781 (N_781,In_2428,In_2482);
nand U782 (N_782,In_1601,In_1653);
nand U783 (N_783,In_566,In_1275);
or U784 (N_784,In_2182,In_553);
xor U785 (N_785,In_1731,In_499);
nor U786 (N_786,In_258,In_1513);
or U787 (N_787,In_319,In_1386);
xor U788 (N_788,In_34,In_979);
or U789 (N_789,In_776,In_2247);
or U790 (N_790,In_1603,In_2371);
nor U791 (N_791,In_458,In_2313);
nand U792 (N_792,In_316,In_709);
nand U793 (N_793,In_70,In_611);
xnor U794 (N_794,In_820,In_1746);
nor U795 (N_795,In_833,In_256);
nor U796 (N_796,In_1663,In_897);
xnor U797 (N_797,In_630,In_1494);
or U798 (N_798,In_146,In_1813);
nor U799 (N_799,In_2372,In_2012);
xnor U800 (N_800,In_1176,In_178);
xor U801 (N_801,In_1732,In_1009);
nand U802 (N_802,In_1332,In_432);
xnor U803 (N_803,In_413,In_1951);
nor U804 (N_804,In_744,In_1276);
nand U805 (N_805,In_205,In_39);
xnor U806 (N_806,In_360,In_1551);
nand U807 (N_807,In_2041,In_1092);
or U808 (N_808,In_757,In_923);
nor U809 (N_809,In_22,In_2256);
xnor U810 (N_810,In_1927,In_868);
nand U811 (N_811,In_2341,In_564);
nand U812 (N_812,In_1830,In_850);
nand U813 (N_813,In_672,In_2107);
xor U814 (N_814,In_2277,In_2153);
or U815 (N_815,In_1913,In_2090);
nand U816 (N_816,In_2015,In_1929);
nor U817 (N_817,In_420,In_2323);
nand U818 (N_818,In_1861,In_832);
nand U819 (N_819,In_336,In_1925);
nor U820 (N_820,In_1255,In_1184);
or U821 (N_821,In_1607,In_1911);
or U822 (N_822,In_445,In_225);
and U823 (N_823,In_512,In_1780);
xnor U824 (N_824,In_1252,In_1742);
nand U825 (N_825,In_1188,In_2094);
xnor U826 (N_826,In_865,In_2214);
xnor U827 (N_827,In_1978,In_1994);
or U828 (N_828,In_2399,In_2342);
nand U829 (N_829,In_780,In_69);
nand U830 (N_830,In_75,In_869);
xnor U831 (N_831,In_417,In_2347);
xnor U832 (N_832,In_920,In_1675);
nand U833 (N_833,In_2262,In_1041);
nand U834 (N_834,In_918,In_597);
xor U835 (N_835,In_1174,In_1536);
and U836 (N_836,In_1510,In_950);
and U837 (N_837,In_627,In_1183);
or U838 (N_838,In_1440,In_340);
xor U839 (N_839,In_1061,In_517);
and U840 (N_840,In_2092,In_1236);
xor U841 (N_841,In_1810,In_144);
or U842 (N_842,In_2416,In_1594);
or U843 (N_843,In_742,In_883);
nor U844 (N_844,In_327,In_1269);
nor U845 (N_845,In_392,In_1665);
and U846 (N_846,In_887,In_2058);
or U847 (N_847,In_2358,In_977);
xor U848 (N_848,In_2261,In_189);
and U849 (N_849,In_1823,In_355);
or U850 (N_850,In_1079,In_698);
xor U851 (N_851,In_143,In_1667);
and U852 (N_852,In_409,In_1219);
nand U853 (N_853,In_592,In_1182);
or U854 (N_854,In_23,In_1272);
and U855 (N_855,In_7,In_660);
nor U856 (N_856,In_15,In_10);
nor U857 (N_857,In_2178,In_38);
or U858 (N_858,In_646,In_65);
or U859 (N_859,In_2340,In_1216);
or U860 (N_860,In_778,In_2490);
nand U861 (N_861,In_1807,In_290);
or U862 (N_862,In_1586,In_1514);
xor U863 (N_863,In_1337,In_387);
or U864 (N_864,In_224,In_2334);
and U865 (N_865,In_1329,In_1862);
or U866 (N_866,In_165,In_2002);
xnor U867 (N_867,In_924,In_944);
xnor U868 (N_868,In_791,In_167);
or U869 (N_869,In_2125,In_331);
or U870 (N_870,In_2407,In_350);
xnor U871 (N_871,In_862,In_1362);
nand U872 (N_872,In_2425,In_1228);
and U873 (N_873,In_1773,In_814);
or U874 (N_874,In_436,In_2089);
nor U875 (N_875,In_1393,In_1906);
xor U876 (N_876,In_479,In_1923);
or U877 (N_877,In_2061,In_2040);
nor U878 (N_878,In_828,In_1521);
nor U879 (N_879,In_1325,In_1408);
nand U880 (N_880,In_1166,In_1470);
or U881 (N_881,In_1899,In_2470);
nand U882 (N_882,In_154,In_1791);
and U883 (N_883,In_1811,In_1976);
nor U884 (N_884,In_2216,In_161);
or U885 (N_885,In_727,In_2240);
or U886 (N_886,In_692,In_273);
or U887 (N_887,In_966,In_1962);
nand U888 (N_888,In_2411,In_1006);
nand U889 (N_889,In_925,In_797);
nand U890 (N_890,In_2440,In_751);
and U891 (N_891,In_363,In_483);
nand U892 (N_892,In_463,In_353);
and U893 (N_893,In_1725,In_1207);
or U894 (N_894,In_1967,In_2208);
or U895 (N_895,In_138,In_2197);
nand U896 (N_896,In_2044,In_1313);
nor U897 (N_897,In_1258,In_2069);
or U898 (N_898,In_1935,In_1192);
or U899 (N_899,In_430,In_2213);
nand U900 (N_900,In_2281,In_1153);
or U901 (N_901,In_1367,In_856);
nor U902 (N_902,In_1879,In_2385);
nand U903 (N_903,In_822,In_2031);
nor U904 (N_904,In_99,In_1401);
xnor U905 (N_905,In_1088,In_922);
nand U906 (N_906,In_2300,In_1438);
nand U907 (N_907,In_2202,In_1843);
nand U908 (N_908,In_2123,In_1083);
nand U909 (N_909,In_2386,In_2274);
or U910 (N_910,In_2105,In_740);
nand U911 (N_911,In_1022,In_1778);
and U912 (N_912,In_1495,In_953);
or U913 (N_913,In_1224,In_957);
and U914 (N_914,In_1243,In_1938);
or U915 (N_915,In_1636,In_1448);
nor U916 (N_916,In_722,In_230);
xor U917 (N_917,In_262,In_1026);
nor U918 (N_918,In_930,In_902);
nand U919 (N_919,In_1023,In_1466);
and U920 (N_920,In_596,In_5);
nor U921 (N_921,In_2009,In_648);
nor U922 (N_922,In_1685,In_1287);
xor U923 (N_923,In_1271,In_1774);
xnor U924 (N_924,In_1503,In_719);
nand U925 (N_925,In_1743,In_1008);
or U926 (N_926,In_418,In_1758);
nor U927 (N_927,In_2412,In_1877);
xnor U928 (N_928,In_1230,In_94);
and U929 (N_929,In_792,In_746);
nand U930 (N_930,In_339,In_1575);
and U931 (N_931,In_919,In_1205);
and U932 (N_932,In_2074,In_514);
xnor U933 (N_933,In_1121,In_606);
xor U934 (N_934,In_586,In_2455);
nor U935 (N_935,In_1013,In_852);
nor U936 (N_936,In_831,In_1646);
or U937 (N_937,In_1677,In_2317);
or U938 (N_938,In_1728,In_1547);
and U939 (N_939,In_1856,In_2156);
and U940 (N_940,In_220,In_795);
or U941 (N_941,In_1489,In_500);
or U942 (N_942,In_1629,In_1414);
xor U943 (N_943,In_1419,In_87);
nand U944 (N_944,In_761,In_1054);
nand U945 (N_945,In_511,In_730);
nor U946 (N_946,In_2071,In_1170);
or U947 (N_947,In_1581,In_1706);
and U948 (N_948,In_609,In_874);
nor U949 (N_949,In_160,In_1281);
nor U950 (N_950,In_2059,In_2229);
and U951 (N_951,In_2159,In_1880);
and U952 (N_952,In_1165,In_1094);
xnor U953 (N_953,In_236,In_677);
xor U954 (N_954,In_439,In_1757);
nor U955 (N_955,In_1627,In_949);
or U956 (N_956,In_1772,In_910);
and U957 (N_957,In_2339,In_559);
or U958 (N_958,In_1291,In_82);
xnor U959 (N_959,In_1103,In_1563);
and U960 (N_960,In_378,In_2139);
nand U961 (N_961,In_1391,In_408);
nand U962 (N_962,In_1589,In_1363);
nor U963 (N_963,In_2210,In_2478);
or U964 (N_964,In_1953,In_134);
nor U965 (N_965,In_1098,In_1577);
nor U966 (N_966,In_130,In_207);
and U967 (N_967,In_1684,In_2231);
or U968 (N_968,In_1615,In_1986);
nand U969 (N_969,In_2491,In_1985);
and U970 (N_970,In_2465,In_1118);
and U971 (N_971,In_542,In_394);
and U972 (N_972,In_1618,In_2003);
nor U973 (N_973,In_1107,In_973);
nor U974 (N_974,In_2241,In_30);
and U975 (N_975,In_502,In_1396);
nor U976 (N_976,In_1609,In_1554);
nor U977 (N_977,In_945,In_1606);
and U978 (N_978,In_1720,In_1960);
and U979 (N_979,In_1158,In_2265);
xnor U980 (N_980,In_2114,In_1015);
or U981 (N_981,In_1395,In_1928);
xor U982 (N_982,In_2102,In_441);
nor U983 (N_983,In_817,In_737);
xnor U984 (N_984,In_2279,In_836);
nand U985 (N_985,In_1235,In_1030);
and U986 (N_986,In_1239,In_1844);
nor U987 (N_987,In_2481,In_2467);
nor U988 (N_988,In_558,In_540);
xnor U989 (N_989,In_1775,In_1027);
nor U990 (N_990,In_1327,In_95);
or U991 (N_991,In_2022,In_636);
or U992 (N_992,In_2246,In_194);
nand U993 (N_993,In_1477,In_673);
or U994 (N_994,In_847,In_687);
nor U995 (N_995,In_631,In_926);
or U996 (N_996,In_44,In_1644);
nand U997 (N_997,In_2285,In_1737);
nor U998 (N_998,In_2302,In_880);
xnor U999 (N_999,In_927,In_2364);
xnor U1000 (N_1000,In_1945,In_348);
nand U1001 (N_1001,In_97,In_2298);
and U1002 (N_1002,In_1454,In_270);
or U1003 (N_1003,In_467,In_1177);
nor U1004 (N_1004,In_1543,In_1961);
or U1005 (N_1005,In_2291,In_108);
nand U1006 (N_1006,In_357,In_1282);
nand U1007 (N_1007,In_935,In_1500);
nand U1008 (N_1008,In_1956,In_198);
and U1009 (N_1009,In_145,In_240);
and U1010 (N_1010,In_655,In_2146);
nor U1011 (N_1011,In_1863,In_1834);
or U1012 (N_1012,In_1405,In_561);
or U1013 (N_1013,In_1836,In_826);
nand U1014 (N_1014,In_901,In_2180);
and U1015 (N_1015,In_563,In_991);
xor U1016 (N_1016,In_1110,In_431);
nor U1017 (N_1017,In_681,In_1937);
or U1018 (N_1018,In_731,In_2112);
or U1019 (N_1019,In_1019,In_853);
nor U1020 (N_1020,In_292,In_1540);
and U1021 (N_1021,In_1072,In_2119);
nor U1022 (N_1022,In_1137,In_2345);
nand U1023 (N_1023,In_1064,In_2221);
nand U1024 (N_1024,In_486,In_1144);
xnor U1025 (N_1025,In_244,In_628);
xnor U1026 (N_1026,In_621,In_404);
xor U1027 (N_1027,In_2104,In_1293);
and U1028 (N_1028,In_2315,In_2184);
nand U1029 (N_1029,In_1971,In_634);
and U1030 (N_1030,In_955,In_306);
or U1031 (N_1031,In_196,In_2257);
nor U1032 (N_1032,In_2014,In_1578);
and U1033 (N_1033,In_582,In_1487);
and U1034 (N_1034,In_330,In_1648);
xnor U1035 (N_1035,In_1752,In_317);
nand U1036 (N_1036,In_1686,In_504);
and U1037 (N_1037,In_779,In_896);
nor U1038 (N_1038,In_637,In_1010);
nand U1039 (N_1039,In_1302,In_2377);
or U1040 (N_1040,In_126,In_454);
xnor U1041 (N_1041,In_320,In_2271);
nand U1042 (N_1042,In_313,In_443);
and U1043 (N_1043,In_1122,In_1031);
nand U1044 (N_1044,In_2035,In_546);
xnor U1045 (N_1045,In_2452,In_997);
or U1046 (N_1046,In_812,In_1403);
nand U1047 (N_1047,In_741,In_2106);
and U1048 (N_1048,In_1765,In_232);
or U1049 (N_1049,In_17,In_1794);
or U1050 (N_1050,In_24,In_1613);
nor U1051 (N_1051,In_2095,In_789);
and U1052 (N_1052,In_1365,In_184);
or U1053 (N_1053,In_133,In_2142);
and U1054 (N_1054,In_1854,In_115);
nor U1055 (N_1055,In_2337,In_1215);
and U1056 (N_1056,In_913,In_380);
nand U1057 (N_1057,In_11,In_2172);
xor U1058 (N_1058,In_1805,In_1308);
and U1059 (N_1059,In_1708,In_1579);
xor U1060 (N_1060,In_1539,In_2397);
xnor U1061 (N_1061,In_45,In_667);
xor U1062 (N_1062,In_503,In_2048);
nor U1063 (N_1063,In_1043,In_2191);
xor U1064 (N_1064,In_861,In_142);
xnor U1065 (N_1065,In_1800,In_2067);
and U1066 (N_1066,In_369,In_2068);
nor U1067 (N_1067,In_645,In_1259);
or U1068 (N_1068,In_613,In_2454);
nor U1069 (N_1069,In_685,In_759);
xor U1070 (N_1070,In_656,In_429);
or U1071 (N_1071,In_845,In_2248);
xor U1072 (N_1072,In_1894,In_1556);
or U1073 (N_1073,In_893,In_2137);
xnor U1074 (N_1074,In_985,In_1091);
and U1075 (N_1075,In_2443,In_716);
or U1076 (N_1076,In_1864,In_1984);
and U1077 (N_1077,In_1140,In_485);
nor U1078 (N_1078,In_285,In_710);
or U1079 (N_1079,In_478,In_1476);
and U1080 (N_1080,In_1833,In_1342);
xnor U1081 (N_1081,In_176,In_1593);
and U1082 (N_1082,In_1164,In_1274);
nand U1083 (N_1083,In_1977,In_2417);
nand U1084 (N_1084,In_1002,In_530);
xnor U1085 (N_1085,In_2310,In_885);
nand U1086 (N_1086,In_2057,In_588);
or U1087 (N_1087,In_1631,In_903);
xnor U1088 (N_1088,In_1922,In_904);
xnor U1089 (N_1089,In_1608,In_1748);
nand U1090 (N_1090,In_916,In_1173);
or U1091 (N_1091,In_1322,In_460);
and U1092 (N_1092,In_2368,In_1377);
nor U1093 (N_1093,In_547,In_1533);
xnor U1094 (N_1094,In_2475,In_501);
and U1095 (N_1095,In_2361,In_1032);
xnor U1096 (N_1096,In_349,In_1082);
or U1097 (N_1097,In_60,In_1763);
nor U1098 (N_1098,In_29,In_1806);
xor U1099 (N_1099,In_1996,In_1950);
nor U1100 (N_1100,In_1696,In_352);
or U1101 (N_1101,In_76,In_841);
nand U1102 (N_1102,In_2200,In_440);
and U1103 (N_1103,In_2150,In_12);
xor U1104 (N_1104,In_1099,In_1000);
nand U1105 (N_1105,In_1512,In_2189);
and U1106 (N_1106,In_1826,In_1892);
xor U1107 (N_1107,In_1375,In_1242);
nor U1108 (N_1108,In_1317,In_169);
or U1109 (N_1109,In_2252,In_1381);
and U1110 (N_1110,In_807,In_1049);
nor U1111 (N_1111,In_601,In_1717);
xor U1112 (N_1112,In_1385,In_870);
or U1113 (N_1113,In_368,In_289);
nor U1114 (N_1114,In_424,In_268);
xor U1115 (N_1115,In_1610,In_974);
and U1116 (N_1116,In_2468,In_2379);
nand U1117 (N_1117,In_774,In_1509);
and U1118 (N_1118,In_1078,In_568);
and U1119 (N_1119,In_931,In_921);
and U1120 (N_1120,In_697,In_1233);
xor U1121 (N_1121,In_1723,In_1279);
or U1122 (N_1122,In_1740,In_2463);
and U1123 (N_1123,In_1642,In_2381);
or U1124 (N_1124,In_843,In_2287);
nand U1125 (N_1125,In_1924,In_1146);
and U1126 (N_1126,In_2384,In_1345);
and U1127 (N_1127,In_2019,In_1840);
nand U1128 (N_1128,In_1491,In_202);
xnor U1129 (N_1129,In_1803,In_2157);
nand U1130 (N_1130,In_2400,In_1139);
and U1131 (N_1131,In_2161,In_1056);
or U1132 (N_1132,In_1516,In_996);
xor U1133 (N_1133,In_6,In_2437);
nand U1134 (N_1134,In_595,In_2006);
or U1135 (N_1135,In_321,In_2445);
or U1136 (N_1136,In_1949,In_109);
xnor U1137 (N_1137,In_464,In_295);
xor U1138 (N_1138,In_400,In_1288);
nor U1139 (N_1139,In_1808,In_364);
xor U1140 (N_1140,In_952,In_1356);
or U1141 (N_1141,In_1465,In_1719);
xor U1142 (N_1142,In_2406,In_1858);
nor U1143 (N_1143,In_1051,In_2025);
nand U1144 (N_1144,In_215,In_1710);
xor U1145 (N_1145,In_14,In_703);
nor U1146 (N_1146,In_2275,In_1266);
xnor U1147 (N_1147,In_2165,In_873);
or U1148 (N_1148,In_1472,In_1304);
nor U1149 (N_1149,In_2,In_1998);
and U1150 (N_1150,In_1903,In_188);
or U1151 (N_1151,In_809,In_1647);
or U1152 (N_1152,In_1574,In_1972);
or U1153 (N_1153,In_860,In_1264);
xor U1154 (N_1154,In_1241,In_1751);
or U1155 (N_1155,In_166,In_2329);
xor U1156 (N_1156,In_1498,In_37);
xor U1157 (N_1157,In_972,In_1296);
xor U1158 (N_1158,In_1461,In_1194);
or U1159 (N_1159,In_2234,In_2220);
nand U1160 (N_1160,In_2043,In_2077);
xor U1161 (N_1161,In_2096,In_191);
or U1162 (N_1162,In_1942,In_255);
xor U1163 (N_1163,In_1109,In_2004);
nor U1164 (N_1164,In_1237,In_2236);
nor U1165 (N_1165,In_245,In_242);
nor U1166 (N_1166,In_1007,In_2117);
and U1167 (N_1167,In_2135,In_736);
nand U1168 (N_1168,In_1659,In_846);
nor U1169 (N_1169,In_1558,In_473);
nand U1170 (N_1170,In_193,In_2085);
nor U1171 (N_1171,In_2238,In_1885);
nand U1172 (N_1172,In_735,In_777);
or U1173 (N_1173,In_2306,In_96);
nand U1174 (N_1174,In_905,In_1415);
nand U1175 (N_1175,In_1486,In_1246);
nor U1176 (N_1176,In_818,In_1126);
and U1177 (N_1177,In_1904,In_967);
nor U1178 (N_1178,In_1209,In_1955);
or U1179 (N_1179,In_2466,In_650);
and U1180 (N_1180,In_9,In_881);
xor U1181 (N_1181,In_1564,In_382);
and U1182 (N_1182,In_1323,In_616);
nor U1183 (N_1183,In_875,In_1452);
nor U1184 (N_1184,In_1643,In_398);
nand U1185 (N_1185,In_72,In_1545);
xnor U1186 (N_1186,In_1179,In_495);
nand U1187 (N_1187,In_2186,In_1760);
or U1188 (N_1188,In_705,In_753);
xor U1189 (N_1189,In_1682,In_2051);
nor U1190 (N_1190,In_214,In_1212);
nand U1191 (N_1191,In_1161,In_1681);
nor U1192 (N_1192,In_442,In_1566);
xnor U1193 (N_1193,In_379,In_683);
xnor U1194 (N_1194,In_1595,In_2016);
xor U1195 (N_1195,In_496,In_834);
nor U1196 (N_1196,In_346,In_1299);
xor U1197 (N_1197,In_477,In_569);
nor U1198 (N_1198,In_324,In_1301);
nor U1199 (N_1199,In_1156,In_1842);
and U1200 (N_1200,In_871,In_1226);
or U1201 (N_1201,In_2076,In_855);
xor U1202 (N_1202,In_1783,In_1364);
or U1203 (N_1203,In_1417,In_1814);
xnor U1204 (N_1204,In_1354,In_374);
nand U1205 (N_1205,In_1499,In_857);
and U1206 (N_1206,In_1326,In_150);
nor U1207 (N_1207,In_829,In_877);
or U1208 (N_1208,In_180,In_750);
or U1209 (N_1209,In_281,In_1557);
and U1210 (N_1210,In_1821,In_1100);
nand U1211 (N_1211,In_2177,In_435);
and U1212 (N_1212,In_1384,In_1443);
and U1213 (N_1213,In_163,In_395);
nand U1214 (N_1214,In_1802,In_341);
or U1215 (N_1215,In_1542,In_2448);
or U1216 (N_1216,In_848,In_615);
and U1217 (N_1217,In_1570,In_253);
or U1218 (N_1218,In_535,In_246);
nor U1219 (N_1219,In_520,In_122);
or U1220 (N_1220,In_1573,In_2456);
xnor U1221 (N_1221,In_2005,In_1366);
and U1222 (N_1222,In_465,In_583);
and U1223 (N_1223,In_906,In_649);
xor U1224 (N_1224,In_1199,In_1383);
nor U1225 (N_1225,In_1909,In_2062);
nor U1226 (N_1226,In_125,In_1785);
xnor U1227 (N_1227,In_1286,In_3);
xnor U1228 (N_1228,In_302,In_2496);
and U1229 (N_1229,In_2324,In_551);
or U1230 (N_1230,In_689,In_1289);
xor U1231 (N_1231,In_554,In_1515);
nor U1232 (N_1232,In_1868,In_2030);
xnor U1233 (N_1233,In_1848,In_1247);
xnor U1234 (N_1234,In_2423,In_2419);
nor U1235 (N_1235,In_602,In_942);
and U1236 (N_1236,In_1341,In_1133);
and U1237 (N_1237,In_1077,In_882);
nand U1238 (N_1238,In_2070,In_965);
nand U1239 (N_1239,In_2223,In_151);
and U1240 (N_1240,In_1080,In_1699);
and U1241 (N_1241,In_1310,In_1590);
or U1242 (N_1242,In_2362,In_1157);
and U1243 (N_1243,In_1480,In_2145);
nand U1244 (N_1244,In_811,In_1523);
nor U1245 (N_1245,In_2414,In_2497);
nor U1246 (N_1246,In_1988,In_1460);
or U1247 (N_1247,In_1335,In_415);
nor U1248 (N_1248,In_1572,In_728);
or U1249 (N_1249,In_261,In_2264);
xnor U1250 (N_1250,N_615,N_1051);
or U1251 (N_1251,N_152,N_1081);
xnor U1252 (N_1252,N_196,N_449);
xnor U1253 (N_1253,N_1094,N_656);
nor U1254 (N_1254,N_210,N_93);
or U1255 (N_1255,N_648,N_249);
xor U1256 (N_1256,N_3,N_310);
xnor U1257 (N_1257,N_979,N_876);
nand U1258 (N_1258,N_805,N_198);
and U1259 (N_1259,N_398,N_544);
and U1260 (N_1260,N_42,N_146);
nand U1261 (N_1261,N_899,N_211);
or U1262 (N_1262,N_1182,N_965);
nand U1263 (N_1263,N_936,N_238);
nand U1264 (N_1264,N_387,N_241);
xor U1265 (N_1265,N_694,N_406);
nand U1266 (N_1266,N_10,N_135);
xor U1267 (N_1267,N_1199,N_415);
and U1268 (N_1268,N_930,N_914);
nand U1269 (N_1269,N_560,N_219);
or U1270 (N_1270,N_453,N_11);
xnor U1271 (N_1271,N_1083,N_1211);
nor U1272 (N_1272,N_263,N_651);
and U1273 (N_1273,N_131,N_520);
nand U1274 (N_1274,N_828,N_252);
nand U1275 (N_1275,N_773,N_117);
nand U1276 (N_1276,N_357,N_500);
nand U1277 (N_1277,N_348,N_1136);
nand U1278 (N_1278,N_1217,N_511);
xnor U1279 (N_1279,N_386,N_827);
nand U1280 (N_1280,N_32,N_138);
or U1281 (N_1281,N_153,N_507);
or U1282 (N_1282,N_854,N_1236);
nor U1283 (N_1283,N_162,N_354);
nor U1284 (N_1284,N_517,N_802);
and U1285 (N_1285,N_31,N_207);
or U1286 (N_1286,N_629,N_314);
xnor U1287 (N_1287,N_1041,N_705);
nand U1288 (N_1288,N_142,N_562);
nand U1289 (N_1289,N_1181,N_312);
or U1290 (N_1290,N_680,N_701);
nand U1291 (N_1291,N_785,N_1075);
nor U1292 (N_1292,N_139,N_659);
nand U1293 (N_1293,N_264,N_23);
and U1294 (N_1294,N_784,N_493);
nor U1295 (N_1295,N_897,N_525);
or U1296 (N_1296,N_477,N_97);
nor U1297 (N_1297,N_401,N_217);
nor U1298 (N_1298,N_1148,N_396);
nor U1299 (N_1299,N_450,N_541);
xor U1300 (N_1300,N_298,N_184);
nor U1301 (N_1301,N_916,N_1110);
and U1302 (N_1302,N_460,N_596);
nor U1303 (N_1303,N_879,N_474);
and U1304 (N_1304,N_815,N_1068);
or U1305 (N_1305,N_924,N_569);
or U1306 (N_1306,N_727,N_860);
nor U1307 (N_1307,N_350,N_951);
xor U1308 (N_1308,N_968,N_833);
xor U1309 (N_1309,N_48,N_794);
and U1310 (N_1310,N_228,N_1089);
xnor U1311 (N_1311,N_208,N_303);
nand U1312 (N_1312,N_1166,N_757);
and U1313 (N_1313,N_110,N_448);
xor U1314 (N_1314,N_990,N_1101);
or U1315 (N_1315,N_837,N_867);
and U1316 (N_1316,N_1018,N_851);
xor U1317 (N_1317,N_684,N_874);
and U1318 (N_1318,N_466,N_457);
nand U1319 (N_1319,N_818,N_334);
and U1320 (N_1320,N_1214,N_1011);
xor U1321 (N_1321,N_408,N_811);
nand U1322 (N_1322,N_942,N_692);
xor U1323 (N_1323,N_1047,N_1109);
nand U1324 (N_1324,N_443,N_693);
and U1325 (N_1325,N_1032,N_842);
nand U1326 (N_1326,N_284,N_1026);
nor U1327 (N_1327,N_452,N_940);
and U1328 (N_1328,N_463,N_1160);
nand U1329 (N_1329,N_649,N_149);
and U1330 (N_1330,N_344,N_1243);
nor U1331 (N_1331,N_133,N_67);
xor U1332 (N_1332,N_319,N_988);
nor U1333 (N_1333,N_148,N_294);
nand U1334 (N_1334,N_46,N_293);
nand U1335 (N_1335,N_253,N_166);
nand U1336 (N_1336,N_1052,N_880);
nand U1337 (N_1337,N_279,N_88);
or U1338 (N_1338,N_1138,N_515);
nor U1339 (N_1339,N_644,N_395);
xor U1340 (N_1340,N_235,N_365);
and U1341 (N_1341,N_480,N_1059);
nor U1342 (N_1342,N_559,N_617);
nor U1343 (N_1343,N_145,N_1050);
or U1344 (N_1344,N_1194,N_60);
xnor U1345 (N_1345,N_341,N_781);
and U1346 (N_1346,N_991,N_958);
nand U1347 (N_1347,N_1092,N_377);
nand U1348 (N_1348,N_804,N_425);
or U1349 (N_1349,N_972,N_335);
nor U1350 (N_1350,N_606,N_588);
xnor U1351 (N_1351,N_761,N_960);
and U1352 (N_1352,N_535,N_826);
xor U1353 (N_1353,N_150,N_782);
and U1354 (N_1354,N_445,N_963);
nor U1355 (N_1355,N_1223,N_6);
and U1356 (N_1356,N_885,N_668);
or U1357 (N_1357,N_130,N_1179);
or U1358 (N_1358,N_58,N_1014);
xnor U1359 (N_1359,N_671,N_502);
and U1360 (N_1360,N_462,N_28);
nand U1361 (N_1361,N_895,N_269);
xnor U1362 (N_1362,N_197,N_1150);
or U1363 (N_1363,N_550,N_571);
or U1364 (N_1364,N_667,N_376);
nand U1365 (N_1365,N_1029,N_928);
nand U1366 (N_1366,N_783,N_866);
or U1367 (N_1367,N_670,N_522);
xor U1368 (N_1368,N_1020,N_278);
and U1369 (N_1369,N_734,N_383);
xnor U1370 (N_1370,N_1095,N_388);
xnor U1371 (N_1371,N_1086,N_937);
or U1372 (N_1372,N_599,N_412);
or U1373 (N_1373,N_640,N_52);
xnor U1374 (N_1374,N_607,N_165);
xor U1375 (N_1375,N_608,N_161);
or U1376 (N_1376,N_498,N_178);
or U1377 (N_1377,N_961,N_1006);
nor U1378 (N_1378,N_1189,N_27);
nor U1379 (N_1379,N_1105,N_89);
nand U1380 (N_1380,N_364,N_1054);
nor U1381 (N_1381,N_191,N_652);
and U1382 (N_1382,N_430,N_1188);
nor U1383 (N_1383,N_246,N_459);
nor U1384 (N_1384,N_1120,N_531);
nor U1385 (N_1385,N_841,N_291);
nor U1386 (N_1386,N_724,N_1207);
or U1387 (N_1387,N_915,N_711);
and U1388 (N_1388,N_179,N_642);
and U1389 (N_1389,N_710,N_25);
nand U1390 (N_1390,N_1132,N_870);
and U1391 (N_1391,N_1146,N_814);
nor U1392 (N_1392,N_790,N_662);
or U1393 (N_1393,N_594,N_66);
nor U1394 (N_1394,N_664,N_1053);
nand U1395 (N_1395,N_168,N_352);
or U1396 (N_1396,N_1162,N_907);
xnor U1397 (N_1397,N_926,N_49);
or U1398 (N_1398,N_688,N_856);
and U1399 (N_1399,N_1111,N_809);
nor U1400 (N_1400,N_70,N_124);
xor U1401 (N_1401,N_1073,N_325);
xor U1402 (N_1402,N_318,N_496);
nand U1403 (N_1403,N_863,N_485);
xor U1404 (N_1404,N_24,N_484);
nor U1405 (N_1405,N_112,N_911);
xor U1406 (N_1406,N_182,N_1072);
and U1407 (N_1407,N_438,N_775);
xor U1408 (N_1408,N_1177,N_759);
xnor U1409 (N_1409,N_691,N_817);
nor U1410 (N_1410,N_796,N_1157);
xor U1411 (N_1411,N_609,N_1159);
and U1412 (N_1412,N_1098,N_546);
nand U1413 (N_1413,N_167,N_487);
nor U1414 (N_1414,N_43,N_1099);
and U1415 (N_1415,N_967,N_185);
or U1416 (N_1416,N_242,N_1155);
and U1417 (N_1417,N_812,N_543);
nor U1418 (N_1418,N_1209,N_1044);
xnor U1419 (N_1419,N_245,N_625);
nor U1420 (N_1420,N_317,N_465);
and U1421 (N_1421,N_679,N_225);
nand U1422 (N_1422,N_360,N_268);
and U1423 (N_1423,N_105,N_1002);
or U1424 (N_1424,N_702,N_1043);
nand U1425 (N_1425,N_250,N_1131);
nor U1426 (N_1426,N_221,N_925);
nand U1427 (N_1427,N_1233,N_714);
nand U1428 (N_1428,N_12,N_800);
and U1429 (N_1429,N_1001,N_1249);
nor U1430 (N_1430,N_94,N_14);
nor U1431 (N_1431,N_21,N_1009);
or U1432 (N_1432,N_33,N_905);
or U1433 (N_1433,N_247,N_313);
xnor U1434 (N_1434,N_855,N_125);
nor U1435 (N_1435,N_266,N_973);
or U1436 (N_1436,N_674,N_488);
and U1437 (N_1437,N_290,N_808);
or U1438 (N_1438,N_382,N_1016);
xnor U1439 (N_1439,N_332,N_427);
xnor U1440 (N_1440,N_1137,N_1142);
nand U1441 (N_1441,N_134,N_434);
and U1442 (N_1442,N_945,N_938);
xor U1443 (N_1443,N_78,N_444);
xor U1444 (N_1444,N_787,N_1208);
or U1445 (N_1445,N_338,N_1124);
xor U1446 (N_1446,N_810,N_1226);
and U1447 (N_1447,N_1064,N_984);
xor U1448 (N_1448,N_156,N_1088);
and U1449 (N_1449,N_657,N_76);
nor U1450 (N_1450,N_255,N_1170);
and U1451 (N_1451,N_995,N_813);
nand U1452 (N_1452,N_409,N_731);
and U1453 (N_1453,N_44,N_939);
nand U1454 (N_1454,N_129,N_1201);
or U1455 (N_1455,N_619,N_1063);
xor U1456 (N_1456,N_1205,N_499);
and U1457 (N_1457,N_1108,N_1235);
xor U1458 (N_1458,N_763,N_590);
nand U1459 (N_1459,N_326,N_1126);
nor U1460 (N_1460,N_1097,N_1225);
nand U1461 (N_1461,N_852,N_470);
nor U1462 (N_1462,N_283,N_144);
nand U1463 (N_1463,N_585,N_307);
xor U1464 (N_1464,N_276,N_512);
and U1465 (N_1465,N_47,N_1143);
nand U1466 (N_1466,N_65,N_935);
or U1467 (N_1467,N_2,N_1245);
nand U1468 (N_1468,N_548,N_737);
and U1469 (N_1469,N_270,N_524);
xnor U1470 (N_1470,N_1145,N_359);
xor U1471 (N_1471,N_473,N_1021);
or U1472 (N_1472,N_844,N_822);
nand U1473 (N_1473,N_795,N_71);
nand U1474 (N_1474,N_884,N_232);
nor U1475 (N_1475,N_1173,N_739);
or U1476 (N_1476,N_791,N_865);
nor U1477 (N_1477,N_713,N_1247);
xor U1478 (N_1478,N_1107,N_295);
or U1479 (N_1479,N_568,N_201);
nor U1480 (N_1480,N_140,N_725);
nor U1481 (N_1481,N_476,N_413);
or U1482 (N_1482,N_587,N_141);
or U1483 (N_1483,N_127,N_1234);
xor U1484 (N_1484,N_1195,N_765);
nand U1485 (N_1485,N_706,N_574);
nor U1486 (N_1486,N_723,N_119);
nand U1487 (N_1487,N_621,N_747);
nor U1488 (N_1488,N_402,N_170);
and U1489 (N_1489,N_921,N_34);
xor U1490 (N_1490,N_1154,N_405);
and U1491 (N_1491,N_416,N_454);
or U1492 (N_1492,N_1202,N_561);
xnor U1493 (N_1493,N_8,N_1172);
nor U1494 (N_1494,N_742,N_746);
xor U1495 (N_1495,N_760,N_581);
or U1496 (N_1496,N_859,N_1118);
or U1497 (N_1497,N_411,N_526);
xor U1498 (N_1498,N_1163,N_778);
nor U1499 (N_1499,N_55,N_857);
and U1500 (N_1500,N_749,N_41);
nand U1501 (N_1501,N_464,N_90);
xor U1502 (N_1502,N_205,N_1125);
or U1503 (N_1503,N_687,N_273);
xnor U1504 (N_1504,N_118,N_981);
and U1505 (N_1505,N_1175,N_107);
and U1506 (N_1506,N_189,N_927);
xor U1507 (N_1507,N_831,N_1074);
nand U1508 (N_1508,N_1027,N_40);
or U1509 (N_1509,N_558,N_910);
and U1510 (N_1510,N_573,N_1190);
and U1511 (N_1511,N_918,N_923);
nor U1512 (N_1512,N_489,N_1062);
and U1513 (N_1513,N_1048,N_1116);
and U1514 (N_1514,N_1010,N_986);
and U1515 (N_1515,N_203,N_697);
xnor U1516 (N_1516,N_733,N_100);
xor U1517 (N_1517,N_1219,N_1066);
xnor U1518 (N_1518,N_1114,N_175);
or U1519 (N_1519,N_686,N_390);
and U1520 (N_1520,N_384,N_431);
and U1521 (N_1521,N_906,N_698);
or U1522 (N_1522,N_639,N_901);
nand U1523 (N_1523,N_1206,N_285);
or U1524 (N_1524,N_977,N_77);
xnor U1525 (N_1525,N_735,N_439);
nor U1526 (N_1526,N_115,N_626);
or U1527 (N_1527,N_15,N_661);
nand U1528 (N_1528,N_1004,N_624);
nor U1529 (N_1529,N_952,N_1130);
or U1530 (N_1530,N_738,N_536);
or U1531 (N_1531,N_169,N_1129);
or U1532 (N_1532,N_638,N_770);
or U1533 (N_1533,N_299,N_497);
and U1534 (N_1534,N_302,N_685);
xor U1535 (N_1535,N_1035,N_799);
and U1536 (N_1536,N_964,N_1079);
or U1537 (N_1537,N_446,N_265);
nand U1538 (N_1538,N_780,N_595);
nand U1539 (N_1539,N_435,N_953);
nor U1540 (N_1540,N_69,N_188);
and U1541 (N_1541,N_171,N_776);
or U1542 (N_1542,N_922,N_966);
xor U1543 (N_1543,N_99,N_231);
nand U1544 (N_1544,N_1158,N_351);
or U1545 (N_1545,N_712,N_426);
xnor U1546 (N_1546,N_371,N_275);
and U1547 (N_1547,N_1085,N_985);
or U1548 (N_1548,N_367,N_1218);
xor U1549 (N_1549,N_904,N_92);
nand U1550 (N_1550,N_627,N_1210);
nand U1551 (N_1551,N_478,N_632);
xor U1552 (N_1552,N_1000,N_492);
nor U1553 (N_1553,N_164,N_955);
nand U1554 (N_1554,N_989,N_883);
and U1555 (N_1555,N_614,N_704);
and U1556 (N_1556,N_892,N_603);
nand U1557 (N_1557,N_190,N_946);
xor U1558 (N_1558,N_869,N_1119);
and U1559 (N_1559,N_375,N_437);
or U1560 (N_1560,N_518,N_1007);
nor U1561 (N_1561,N_159,N_533);
xnor U1562 (N_1562,N_240,N_666);
nor U1563 (N_1563,N_954,N_941);
nand U1564 (N_1564,N_1065,N_1008);
or U1565 (N_1565,N_873,N_1036);
and U1566 (N_1566,N_726,N_64);
and U1567 (N_1567,N_421,N_35);
nand U1568 (N_1568,N_1216,N_385);
nor U1569 (N_1569,N_336,N_447);
xor U1570 (N_1570,N_323,N_586);
and U1571 (N_1571,N_494,N_1045);
nand U1572 (N_1572,N_887,N_244);
nand U1573 (N_1573,N_552,N_137);
nand U1574 (N_1574,N_1039,N_163);
or U1575 (N_1575,N_766,N_1121);
nor U1576 (N_1576,N_1149,N_173);
and U1577 (N_1577,N_728,N_881);
or U1578 (N_1578,N_340,N_432);
xor U1579 (N_1579,N_251,N_913);
and U1580 (N_1580,N_700,N_155);
xnor U1581 (N_1581,N_222,N_829);
xor U1582 (N_1582,N_774,N_262);
and U1583 (N_1583,N_505,N_673);
nor U1584 (N_1584,N_0,N_575);
nand U1585 (N_1585,N_393,N_969);
or U1586 (N_1586,N_1187,N_529);
or U1587 (N_1587,N_902,N_637);
and U1588 (N_1588,N_1228,N_391);
xor U1589 (N_1589,N_944,N_1239);
xor U1590 (N_1590,N_779,N_1022);
xnor U1591 (N_1591,N_30,N_214);
or U1592 (N_1592,N_768,N_1003);
and U1593 (N_1593,N_120,N_19);
xnor U1594 (N_1594,N_1090,N_862);
or U1595 (N_1595,N_801,N_123);
and U1596 (N_1596,N_845,N_858);
nand U1597 (N_1597,N_327,N_379);
or U1598 (N_1598,N_17,N_86);
nand U1599 (N_1599,N_1174,N_890);
or U1600 (N_1600,N_423,N_750);
and U1601 (N_1601,N_1220,N_347);
xnor U1602 (N_1602,N_1030,N_1222);
or U1603 (N_1603,N_490,N_1013);
xnor U1604 (N_1604,N_1023,N_839);
and U1605 (N_1605,N_236,N_957);
nor U1606 (N_1606,N_51,N_151);
or U1607 (N_1607,N_337,N_920);
and U1608 (N_1608,N_286,N_226);
xor U1609 (N_1609,N_1198,N_878);
or U1610 (N_1610,N_719,N_730);
or U1611 (N_1611,N_20,N_424);
or U1612 (N_1612,N_1057,N_282);
nor U1613 (N_1613,N_1242,N_786);
nor U1614 (N_1614,N_767,N_81);
xor U1615 (N_1615,N_622,N_553);
nand U1616 (N_1616,N_257,N_847);
xor U1617 (N_1617,N_628,N_557);
nor U1618 (N_1618,N_308,N_180);
and U1619 (N_1619,N_1106,N_206);
xor U1620 (N_1620,N_1005,N_1134);
xnor U1621 (N_1621,N_1196,N_260);
nor U1622 (N_1622,N_160,N_756);
or U1623 (N_1623,N_917,N_523);
nor U1624 (N_1624,N_1197,N_655);
nand U1625 (N_1625,N_1031,N_633);
and U1626 (N_1626,N_732,N_63);
or U1627 (N_1627,N_440,N_147);
or U1628 (N_1628,N_258,N_374);
or U1629 (N_1629,N_194,N_1112);
xor U1630 (N_1630,N_932,N_1213);
xnor U1631 (N_1631,N_328,N_281);
and U1632 (N_1632,N_287,N_378);
nand U1633 (N_1633,N_975,N_72);
and U1634 (N_1634,N_708,N_1093);
and U1635 (N_1635,N_919,N_309);
nand U1636 (N_1636,N_1147,N_992);
nand U1637 (N_1637,N_136,N_1178);
xor U1638 (N_1638,N_634,N_122);
or U1639 (N_1639,N_1084,N_458);
nand U1640 (N_1640,N_539,N_271);
or U1641 (N_1641,N_399,N_613);
nand U1642 (N_1642,N_853,N_53);
and U1643 (N_1643,N_1080,N_433);
xor U1644 (N_1644,N_414,N_534);
and U1645 (N_1645,N_999,N_602);
nor U1646 (N_1646,N_563,N_506);
or U1647 (N_1647,N_1128,N_1091);
xnor U1648 (N_1648,N_1224,N_521);
nor U1649 (N_1649,N_7,N_948);
nor U1650 (N_1650,N_891,N_380);
and U1651 (N_1651,N_1153,N_983);
nand U1652 (N_1652,N_154,N_772);
nor U1653 (N_1653,N_663,N_912);
and U1654 (N_1654,N_600,N_358);
xnor U1655 (N_1655,N_947,N_95);
or U1656 (N_1656,N_669,N_530);
xor U1657 (N_1657,N_641,N_158);
nand U1658 (N_1658,N_567,N_516);
xnor U1659 (N_1659,N_545,N_343);
xor U1660 (N_1660,N_1071,N_132);
nor U1661 (N_1661,N_754,N_9);
nand U1662 (N_1662,N_508,N_549);
and U1663 (N_1663,N_1038,N_987);
or U1664 (N_1664,N_1028,N_1215);
nand U1665 (N_1665,N_1135,N_306);
xor U1666 (N_1666,N_1015,N_1244);
xnor U1667 (N_1667,N_239,N_356);
and U1668 (N_1668,N_540,N_200);
xnor U1669 (N_1669,N_324,N_475);
nand U1670 (N_1670,N_519,N_861);
nor U1671 (N_1671,N_1141,N_1203);
nor U1672 (N_1672,N_1204,N_1200);
and U1673 (N_1673,N_363,N_1248);
nand U1674 (N_1674,N_997,N_223);
nor U1675 (N_1675,N_931,N_1165);
and U1676 (N_1676,N_1104,N_849);
nor U1677 (N_1677,N_537,N_1169);
nand U1678 (N_1678,N_903,N_696);
nand U1679 (N_1679,N_106,N_816);
nor U1680 (N_1680,N_886,N_998);
or U1681 (N_1681,N_630,N_22);
or U1682 (N_1682,N_1161,N_1082);
nor U1683 (N_1683,N_1033,N_769);
nand U1684 (N_1684,N_116,N_830);
nand U1685 (N_1685,N_848,N_703);
xor U1686 (N_1686,N_486,N_102);
nor U1687 (N_1687,N_267,N_909);
nor U1688 (N_1688,N_1140,N_37);
nand U1689 (N_1689,N_894,N_1046);
xor U1690 (N_1690,N_1070,N_610);
xor U1691 (N_1691,N_1024,N_472);
or U1692 (N_1692,N_956,N_403);
nand U1693 (N_1693,N_45,N_584);
nor U1694 (N_1694,N_5,N_1164);
or U1695 (N_1695,N_612,N_740);
or U1696 (N_1696,N_16,N_39);
nand U1697 (N_1697,N_1238,N_777);
xor U1698 (N_1698,N_234,N_771);
or U1699 (N_1699,N_751,N_29);
or U1700 (N_1700,N_26,N_261);
xor U1701 (N_1701,N_803,N_311);
and U1702 (N_1702,N_576,N_1017);
nor U1703 (N_1703,N_1212,N_108);
or U1704 (N_1704,N_82,N_616);
and U1705 (N_1705,N_565,N_461);
nor U1706 (N_1706,N_1019,N_823);
xnor U1707 (N_1707,N_428,N_566);
and U1708 (N_1708,N_825,N_743);
xnor U1709 (N_1709,N_113,N_665);
nand U1710 (N_1710,N_838,N_397);
xnor U1711 (N_1711,N_736,N_748);
and U1712 (N_1712,N_591,N_755);
and U1713 (N_1713,N_220,N_442);
nand U1714 (N_1714,N_62,N_1040);
nor U1715 (N_1715,N_1113,N_193);
or U1716 (N_1716,N_321,N_346);
nor U1717 (N_1717,N_513,N_1069);
xor U1718 (N_1718,N_369,N_54);
nor U1719 (N_1719,N_943,N_1037);
or U1720 (N_1720,N_690,N_900);
or U1721 (N_1721,N_353,N_538);
or U1722 (N_1722,N_843,N_877);
nand U1723 (N_1723,N_882,N_419);
nand U1724 (N_1724,N_469,N_1144);
xor U1725 (N_1725,N_1025,N_788);
and U1726 (N_1726,N_57,N_889);
nand U1727 (N_1727,N_192,N_1087);
and U1728 (N_1728,N_1067,N_741);
xor U1729 (N_1729,N_73,N_84);
xor U1730 (N_1730,N_436,N_650);
or U1731 (N_1731,N_676,N_896);
xor U1732 (N_1732,N_1185,N_495);
or U1733 (N_1733,N_547,N_1061);
or U1734 (N_1734,N_707,N_798);
or U1735 (N_1735,N_38,N_1227);
nand U1736 (N_1736,N_229,N_933);
xor U1737 (N_1737,N_509,N_721);
or U1738 (N_1738,N_316,N_582);
nor U1739 (N_1739,N_392,N_745);
or U1740 (N_1740,N_128,N_87);
nor U1741 (N_1741,N_227,N_504);
xor U1742 (N_1742,N_1049,N_345);
nor U1743 (N_1743,N_83,N_592);
or U1744 (N_1744,N_248,N_611);
and U1745 (N_1745,N_555,N_368);
xnor U1746 (N_1746,N_176,N_59);
nor U1747 (N_1747,N_209,N_660);
nor U1748 (N_1748,N_583,N_501);
nand U1749 (N_1749,N_259,N_233);
nor U1750 (N_1750,N_570,N_304);
nor U1751 (N_1751,N_1012,N_836);
and U1752 (N_1752,N_681,N_564);
nand U1753 (N_1753,N_218,N_1139);
nor U1754 (N_1754,N_361,N_96);
or U1755 (N_1755,N_277,N_764);
xor U1756 (N_1756,N_1058,N_483);
or U1757 (N_1757,N_121,N_1167);
nor U1758 (N_1758,N_1122,N_601);
or U1759 (N_1759,N_18,N_126);
xor U1760 (N_1760,N_1151,N_556);
nor U1761 (N_1761,N_618,N_254);
xnor U1762 (N_1762,N_1034,N_579);
or U1763 (N_1763,N_1103,N_199);
or U1764 (N_1764,N_215,N_978);
and U1765 (N_1765,N_482,N_204);
nor U1766 (N_1766,N_1077,N_1176);
and U1767 (N_1767,N_330,N_195);
or U1768 (N_1768,N_417,N_467);
or U1769 (N_1769,N_551,N_1240);
nand U1770 (N_1770,N_850,N_762);
nor U1771 (N_1771,N_355,N_631);
nor U1772 (N_1772,N_1231,N_976);
nand U1773 (N_1773,N_373,N_908);
nor U1774 (N_1774,N_91,N_56);
nand U1775 (N_1775,N_349,N_1232);
nor U1776 (N_1776,N_456,N_85);
nor U1777 (N_1777,N_605,N_50);
nand U1778 (N_1778,N_394,N_1152);
xor U1779 (N_1779,N_274,N_74);
nor U1780 (N_1780,N_893,N_689);
nand U1781 (N_1781,N_542,N_98);
nand U1782 (N_1782,N_297,N_471);
and U1783 (N_1783,N_4,N_68);
or U1784 (N_1784,N_806,N_934);
and U1785 (N_1785,N_527,N_61);
nor U1786 (N_1786,N_658,N_481);
nand U1787 (N_1787,N_758,N_678);
nor U1788 (N_1788,N_709,N_333);
or U1789 (N_1789,N_871,N_807);
or U1790 (N_1790,N_418,N_720);
nor U1791 (N_1791,N_635,N_1180);
and U1792 (N_1792,N_109,N_329);
or U1793 (N_1793,N_1100,N_339);
and U1794 (N_1794,N_744,N_1237);
and U1795 (N_1795,N_1184,N_410);
nand U1796 (N_1796,N_111,N_832);
nand U1797 (N_1797,N_797,N_717);
or U1798 (N_1798,N_752,N_1115);
nor U1799 (N_1799,N_272,N_181);
xor U1800 (N_1800,N_420,N_503);
and U1801 (N_1801,N_1156,N_80);
and U1802 (N_1802,N_422,N_982);
and U1803 (N_1803,N_331,N_479);
or U1804 (N_1804,N_820,N_1078);
or U1805 (N_1805,N_1102,N_620);
or U1806 (N_1806,N_1230,N_230);
or U1807 (N_1807,N_1096,N_362);
or U1808 (N_1808,N_75,N_1171);
and U1809 (N_1809,N_971,N_578);
and U1810 (N_1810,N_36,N_996);
nor U1811 (N_1811,N_451,N_407);
nand U1812 (N_1812,N_875,N_224);
and U1813 (N_1813,N_532,N_672);
nand U1814 (N_1814,N_959,N_1123);
and U1815 (N_1815,N_1241,N_296);
xnor U1816 (N_1816,N_1042,N_645);
or U1817 (N_1817,N_683,N_288);
nor U1818 (N_1818,N_305,N_301);
and U1819 (N_1819,N_589,N_1186);
nor U1820 (N_1820,N_1191,N_1055);
or U1821 (N_1821,N_834,N_1117);
nor U1822 (N_1822,N_186,N_572);
nand U1823 (N_1823,N_699,N_593);
and U1824 (N_1824,N_1192,N_695);
and U1825 (N_1825,N_980,N_1076);
nor U1826 (N_1826,N_682,N_974);
xnor U1827 (N_1827,N_577,N_256);
nor U1828 (N_1828,N_792,N_623);
or U1829 (N_1829,N_718,N_636);
and U1830 (N_1830,N_289,N_962);
nand U1831 (N_1831,N_597,N_381);
nand U1832 (N_1832,N_342,N_835);
nand U1833 (N_1833,N_929,N_993);
nand U1834 (N_1834,N_819,N_1193);
nand U1835 (N_1835,N_646,N_187);
and U1836 (N_1836,N_202,N_970);
nor U1837 (N_1837,N_872,N_177);
and U1838 (N_1838,N_114,N_216);
and U1839 (N_1839,N_675,N_753);
nor U1840 (N_1840,N_994,N_300);
nand U1841 (N_1841,N_404,N_320);
nor U1842 (N_1842,N_1127,N_213);
nor U1843 (N_1843,N_280,N_514);
nor U1844 (N_1844,N_898,N_716);
nand U1845 (N_1845,N_653,N_950);
xor U1846 (N_1846,N_174,N_101);
and U1847 (N_1847,N_729,N_1229);
nand U1848 (N_1848,N_1060,N_715);
nor U1849 (N_1849,N_143,N_389);
and U1850 (N_1850,N_789,N_104);
nor U1851 (N_1851,N_554,N_1056);
nor U1852 (N_1852,N_212,N_888);
xnor U1853 (N_1853,N_468,N_372);
xnor U1854 (N_1854,N_793,N_846);
xor U1855 (N_1855,N_1,N_315);
xnor U1856 (N_1856,N_400,N_292);
xnor U1857 (N_1857,N_510,N_654);
or U1858 (N_1858,N_604,N_647);
nand U1859 (N_1859,N_13,N_322);
nor U1860 (N_1860,N_528,N_1133);
and U1861 (N_1861,N_441,N_643);
nor U1862 (N_1862,N_157,N_580);
nor U1863 (N_1863,N_1246,N_79);
and U1864 (N_1864,N_183,N_429);
nand U1865 (N_1865,N_824,N_172);
nand U1866 (N_1866,N_1168,N_1221);
and U1867 (N_1867,N_598,N_491);
nand U1868 (N_1868,N_237,N_949);
nand U1869 (N_1869,N_103,N_868);
or U1870 (N_1870,N_864,N_455);
nor U1871 (N_1871,N_370,N_677);
xnor U1872 (N_1872,N_840,N_366);
or U1873 (N_1873,N_821,N_722);
nand U1874 (N_1874,N_1183,N_243);
xnor U1875 (N_1875,N_294,N_504);
nand U1876 (N_1876,N_1207,N_146);
or U1877 (N_1877,N_660,N_1139);
xor U1878 (N_1878,N_688,N_428);
nor U1879 (N_1879,N_705,N_1118);
nand U1880 (N_1880,N_281,N_166);
xnor U1881 (N_1881,N_215,N_184);
xnor U1882 (N_1882,N_910,N_1163);
or U1883 (N_1883,N_235,N_229);
xnor U1884 (N_1884,N_37,N_514);
or U1885 (N_1885,N_764,N_1248);
and U1886 (N_1886,N_5,N_685);
nor U1887 (N_1887,N_1146,N_1166);
or U1888 (N_1888,N_442,N_786);
nor U1889 (N_1889,N_123,N_962);
nand U1890 (N_1890,N_744,N_1232);
nand U1891 (N_1891,N_1185,N_14);
nor U1892 (N_1892,N_1112,N_933);
nor U1893 (N_1893,N_288,N_539);
nor U1894 (N_1894,N_270,N_1069);
or U1895 (N_1895,N_978,N_102);
nand U1896 (N_1896,N_944,N_866);
xor U1897 (N_1897,N_991,N_279);
nor U1898 (N_1898,N_1088,N_444);
or U1899 (N_1899,N_896,N_241);
or U1900 (N_1900,N_388,N_463);
xnor U1901 (N_1901,N_379,N_189);
nor U1902 (N_1902,N_515,N_342);
or U1903 (N_1903,N_659,N_255);
nand U1904 (N_1904,N_536,N_450);
or U1905 (N_1905,N_988,N_499);
xnor U1906 (N_1906,N_103,N_383);
nor U1907 (N_1907,N_212,N_191);
xnor U1908 (N_1908,N_645,N_531);
or U1909 (N_1909,N_813,N_349);
xnor U1910 (N_1910,N_1245,N_1096);
or U1911 (N_1911,N_653,N_176);
and U1912 (N_1912,N_398,N_455);
or U1913 (N_1913,N_913,N_118);
nor U1914 (N_1914,N_728,N_1173);
or U1915 (N_1915,N_334,N_5);
nor U1916 (N_1916,N_498,N_969);
or U1917 (N_1917,N_30,N_894);
or U1918 (N_1918,N_839,N_953);
and U1919 (N_1919,N_489,N_640);
xnor U1920 (N_1920,N_527,N_1169);
nand U1921 (N_1921,N_538,N_3);
nor U1922 (N_1922,N_921,N_1238);
or U1923 (N_1923,N_156,N_482);
or U1924 (N_1924,N_1096,N_135);
xnor U1925 (N_1925,N_800,N_1142);
nand U1926 (N_1926,N_333,N_913);
and U1927 (N_1927,N_901,N_437);
nor U1928 (N_1928,N_813,N_987);
nand U1929 (N_1929,N_384,N_535);
xnor U1930 (N_1930,N_489,N_387);
xnor U1931 (N_1931,N_450,N_438);
xor U1932 (N_1932,N_1186,N_668);
xor U1933 (N_1933,N_961,N_371);
nor U1934 (N_1934,N_1029,N_778);
and U1935 (N_1935,N_447,N_139);
or U1936 (N_1936,N_153,N_236);
nor U1937 (N_1937,N_1121,N_108);
nor U1938 (N_1938,N_759,N_139);
xnor U1939 (N_1939,N_705,N_1200);
xor U1940 (N_1940,N_1150,N_971);
nand U1941 (N_1941,N_36,N_230);
or U1942 (N_1942,N_500,N_1206);
xnor U1943 (N_1943,N_168,N_856);
or U1944 (N_1944,N_592,N_664);
and U1945 (N_1945,N_88,N_11);
nand U1946 (N_1946,N_391,N_40);
and U1947 (N_1947,N_784,N_501);
nand U1948 (N_1948,N_660,N_103);
nor U1949 (N_1949,N_1170,N_507);
nor U1950 (N_1950,N_669,N_1006);
and U1951 (N_1951,N_933,N_948);
xnor U1952 (N_1952,N_704,N_130);
xnor U1953 (N_1953,N_139,N_549);
and U1954 (N_1954,N_191,N_873);
or U1955 (N_1955,N_1035,N_234);
nor U1956 (N_1956,N_482,N_135);
or U1957 (N_1957,N_482,N_25);
and U1958 (N_1958,N_556,N_307);
or U1959 (N_1959,N_34,N_905);
nand U1960 (N_1960,N_1199,N_820);
nor U1961 (N_1961,N_354,N_997);
nand U1962 (N_1962,N_903,N_998);
nor U1963 (N_1963,N_132,N_722);
xnor U1964 (N_1964,N_1249,N_393);
xnor U1965 (N_1965,N_814,N_470);
nand U1966 (N_1966,N_704,N_1140);
xnor U1967 (N_1967,N_433,N_950);
or U1968 (N_1968,N_111,N_838);
nand U1969 (N_1969,N_711,N_1044);
or U1970 (N_1970,N_793,N_955);
or U1971 (N_1971,N_514,N_1032);
and U1972 (N_1972,N_652,N_267);
xnor U1973 (N_1973,N_576,N_120);
nand U1974 (N_1974,N_433,N_924);
and U1975 (N_1975,N_1093,N_803);
and U1976 (N_1976,N_937,N_75);
xor U1977 (N_1977,N_529,N_756);
nand U1978 (N_1978,N_593,N_17);
xor U1979 (N_1979,N_818,N_365);
and U1980 (N_1980,N_236,N_1110);
or U1981 (N_1981,N_713,N_939);
or U1982 (N_1982,N_800,N_299);
nor U1983 (N_1983,N_691,N_1037);
or U1984 (N_1984,N_565,N_871);
nor U1985 (N_1985,N_727,N_16);
nand U1986 (N_1986,N_1188,N_984);
nor U1987 (N_1987,N_951,N_784);
nand U1988 (N_1988,N_108,N_512);
or U1989 (N_1989,N_634,N_120);
and U1990 (N_1990,N_1049,N_572);
and U1991 (N_1991,N_720,N_262);
xor U1992 (N_1992,N_864,N_577);
or U1993 (N_1993,N_613,N_364);
or U1994 (N_1994,N_790,N_719);
and U1995 (N_1995,N_20,N_289);
nand U1996 (N_1996,N_347,N_114);
nor U1997 (N_1997,N_560,N_505);
nor U1998 (N_1998,N_776,N_473);
or U1999 (N_1999,N_553,N_900);
or U2000 (N_2000,N_736,N_1187);
nor U2001 (N_2001,N_35,N_235);
or U2002 (N_2002,N_1170,N_1086);
and U2003 (N_2003,N_850,N_1225);
and U2004 (N_2004,N_758,N_780);
xor U2005 (N_2005,N_973,N_1104);
and U2006 (N_2006,N_1025,N_957);
nor U2007 (N_2007,N_111,N_726);
and U2008 (N_2008,N_217,N_1143);
or U2009 (N_2009,N_1183,N_494);
or U2010 (N_2010,N_636,N_1189);
nand U2011 (N_2011,N_195,N_1153);
nand U2012 (N_2012,N_194,N_1220);
nand U2013 (N_2013,N_630,N_651);
nor U2014 (N_2014,N_1,N_176);
xor U2015 (N_2015,N_226,N_1079);
nand U2016 (N_2016,N_499,N_1093);
or U2017 (N_2017,N_75,N_1116);
nor U2018 (N_2018,N_174,N_561);
and U2019 (N_2019,N_495,N_1067);
and U2020 (N_2020,N_304,N_896);
nand U2021 (N_2021,N_222,N_647);
or U2022 (N_2022,N_204,N_941);
nor U2023 (N_2023,N_232,N_1085);
xnor U2024 (N_2024,N_1134,N_1221);
and U2025 (N_2025,N_662,N_986);
or U2026 (N_2026,N_469,N_218);
or U2027 (N_2027,N_619,N_83);
xnor U2028 (N_2028,N_110,N_810);
nand U2029 (N_2029,N_1181,N_698);
nand U2030 (N_2030,N_637,N_359);
nor U2031 (N_2031,N_339,N_813);
nand U2032 (N_2032,N_364,N_131);
nand U2033 (N_2033,N_288,N_23);
xnor U2034 (N_2034,N_384,N_339);
xnor U2035 (N_2035,N_341,N_262);
and U2036 (N_2036,N_396,N_875);
or U2037 (N_2037,N_96,N_355);
nand U2038 (N_2038,N_363,N_1214);
nand U2039 (N_2039,N_967,N_123);
or U2040 (N_2040,N_232,N_691);
or U2041 (N_2041,N_1054,N_1091);
nand U2042 (N_2042,N_159,N_770);
xnor U2043 (N_2043,N_983,N_706);
nand U2044 (N_2044,N_1146,N_541);
xor U2045 (N_2045,N_320,N_803);
or U2046 (N_2046,N_829,N_1215);
or U2047 (N_2047,N_730,N_46);
nor U2048 (N_2048,N_390,N_961);
and U2049 (N_2049,N_273,N_548);
xor U2050 (N_2050,N_911,N_964);
nand U2051 (N_2051,N_1242,N_784);
or U2052 (N_2052,N_890,N_793);
or U2053 (N_2053,N_964,N_907);
and U2054 (N_2054,N_1236,N_797);
nand U2055 (N_2055,N_333,N_134);
or U2056 (N_2056,N_797,N_1054);
nor U2057 (N_2057,N_624,N_108);
and U2058 (N_2058,N_1161,N_707);
or U2059 (N_2059,N_615,N_1053);
nand U2060 (N_2060,N_935,N_646);
and U2061 (N_2061,N_1028,N_1056);
or U2062 (N_2062,N_843,N_983);
and U2063 (N_2063,N_573,N_1037);
nor U2064 (N_2064,N_236,N_727);
xor U2065 (N_2065,N_705,N_1224);
xnor U2066 (N_2066,N_1005,N_150);
xnor U2067 (N_2067,N_220,N_757);
nand U2068 (N_2068,N_412,N_44);
xnor U2069 (N_2069,N_658,N_547);
and U2070 (N_2070,N_973,N_1184);
xnor U2071 (N_2071,N_983,N_85);
nand U2072 (N_2072,N_229,N_986);
nor U2073 (N_2073,N_354,N_816);
nand U2074 (N_2074,N_984,N_709);
nand U2075 (N_2075,N_197,N_1085);
nor U2076 (N_2076,N_899,N_986);
nor U2077 (N_2077,N_1024,N_1043);
and U2078 (N_2078,N_1110,N_468);
and U2079 (N_2079,N_410,N_63);
or U2080 (N_2080,N_418,N_643);
or U2081 (N_2081,N_81,N_117);
nor U2082 (N_2082,N_1197,N_785);
and U2083 (N_2083,N_646,N_227);
or U2084 (N_2084,N_416,N_924);
nor U2085 (N_2085,N_392,N_1087);
nand U2086 (N_2086,N_27,N_894);
nor U2087 (N_2087,N_856,N_1075);
xor U2088 (N_2088,N_733,N_899);
and U2089 (N_2089,N_223,N_77);
or U2090 (N_2090,N_156,N_1087);
xnor U2091 (N_2091,N_268,N_1171);
xnor U2092 (N_2092,N_227,N_205);
nor U2093 (N_2093,N_575,N_1053);
xnor U2094 (N_2094,N_137,N_218);
nor U2095 (N_2095,N_1051,N_366);
nand U2096 (N_2096,N_273,N_703);
nand U2097 (N_2097,N_1221,N_130);
xor U2098 (N_2098,N_775,N_416);
or U2099 (N_2099,N_863,N_1249);
nor U2100 (N_2100,N_615,N_920);
and U2101 (N_2101,N_893,N_172);
and U2102 (N_2102,N_127,N_480);
and U2103 (N_2103,N_1159,N_840);
and U2104 (N_2104,N_716,N_458);
nand U2105 (N_2105,N_987,N_613);
xor U2106 (N_2106,N_184,N_1025);
nand U2107 (N_2107,N_288,N_513);
nand U2108 (N_2108,N_1024,N_495);
nand U2109 (N_2109,N_443,N_377);
xnor U2110 (N_2110,N_1063,N_494);
nor U2111 (N_2111,N_924,N_465);
xnor U2112 (N_2112,N_1035,N_64);
xnor U2113 (N_2113,N_496,N_559);
or U2114 (N_2114,N_642,N_1164);
nor U2115 (N_2115,N_381,N_736);
or U2116 (N_2116,N_474,N_535);
nor U2117 (N_2117,N_1186,N_1013);
or U2118 (N_2118,N_455,N_348);
xor U2119 (N_2119,N_1192,N_655);
and U2120 (N_2120,N_757,N_44);
nand U2121 (N_2121,N_1094,N_562);
xor U2122 (N_2122,N_1215,N_352);
or U2123 (N_2123,N_225,N_964);
and U2124 (N_2124,N_989,N_381);
xor U2125 (N_2125,N_13,N_303);
xnor U2126 (N_2126,N_795,N_98);
or U2127 (N_2127,N_727,N_155);
xnor U2128 (N_2128,N_477,N_569);
xor U2129 (N_2129,N_1047,N_575);
and U2130 (N_2130,N_753,N_1026);
or U2131 (N_2131,N_290,N_347);
and U2132 (N_2132,N_159,N_673);
xor U2133 (N_2133,N_202,N_957);
nand U2134 (N_2134,N_1000,N_926);
nor U2135 (N_2135,N_120,N_567);
nand U2136 (N_2136,N_264,N_145);
and U2137 (N_2137,N_273,N_77);
nor U2138 (N_2138,N_1229,N_577);
nor U2139 (N_2139,N_680,N_481);
nor U2140 (N_2140,N_337,N_19);
or U2141 (N_2141,N_1194,N_1045);
or U2142 (N_2142,N_718,N_1123);
xnor U2143 (N_2143,N_312,N_729);
xor U2144 (N_2144,N_71,N_459);
xnor U2145 (N_2145,N_347,N_147);
or U2146 (N_2146,N_401,N_738);
nand U2147 (N_2147,N_487,N_978);
nand U2148 (N_2148,N_446,N_582);
nand U2149 (N_2149,N_910,N_832);
nor U2150 (N_2150,N_135,N_251);
or U2151 (N_2151,N_380,N_227);
and U2152 (N_2152,N_991,N_1177);
and U2153 (N_2153,N_100,N_251);
or U2154 (N_2154,N_352,N_319);
or U2155 (N_2155,N_266,N_175);
nor U2156 (N_2156,N_505,N_1011);
xnor U2157 (N_2157,N_693,N_1204);
and U2158 (N_2158,N_332,N_730);
nand U2159 (N_2159,N_624,N_792);
and U2160 (N_2160,N_692,N_150);
and U2161 (N_2161,N_430,N_682);
nand U2162 (N_2162,N_697,N_186);
and U2163 (N_2163,N_542,N_353);
nand U2164 (N_2164,N_994,N_891);
nand U2165 (N_2165,N_724,N_1053);
nand U2166 (N_2166,N_813,N_362);
and U2167 (N_2167,N_1095,N_807);
nor U2168 (N_2168,N_389,N_757);
or U2169 (N_2169,N_188,N_932);
nand U2170 (N_2170,N_706,N_177);
or U2171 (N_2171,N_456,N_134);
or U2172 (N_2172,N_806,N_1134);
or U2173 (N_2173,N_1111,N_902);
nand U2174 (N_2174,N_278,N_757);
xnor U2175 (N_2175,N_896,N_552);
and U2176 (N_2176,N_842,N_776);
or U2177 (N_2177,N_720,N_800);
nand U2178 (N_2178,N_1029,N_103);
nand U2179 (N_2179,N_363,N_813);
xor U2180 (N_2180,N_157,N_587);
and U2181 (N_2181,N_820,N_617);
xnor U2182 (N_2182,N_1014,N_50);
nor U2183 (N_2183,N_612,N_813);
nor U2184 (N_2184,N_992,N_515);
and U2185 (N_2185,N_485,N_379);
nand U2186 (N_2186,N_322,N_253);
or U2187 (N_2187,N_197,N_676);
nand U2188 (N_2188,N_1069,N_248);
or U2189 (N_2189,N_1000,N_594);
xnor U2190 (N_2190,N_676,N_109);
or U2191 (N_2191,N_377,N_1226);
nand U2192 (N_2192,N_638,N_1121);
nor U2193 (N_2193,N_476,N_1048);
xnor U2194 (N_2194,N_486,N_906);
nand U2195 (N_2195,N_215,N_1167);
or U2196 (N_2196,N_709,N_1093);
and U2197 (N_2197,N_891,N_499);
or U2198 (N_2198,N_741,N_344);
and U2199 (N_2199,N_1089,N_207);
or U2200 (N_2200,N_659,N_346);
and U2201 (N_2201,N_156,N_243);
and U2202 (N_2202,N_450,N_780);
nand U2203 (N_2203,N_732,N_204);
xnor U2204 (N_2204,N_921,N_336);
xnor U2205 (N_2205,N_825,N_1045);
nor U2206 (N_2206,N_1140,N_1155);
and U2207 (N_2207,N_597,N_1199);
nor U2208 (N_2208,N_600,N_5);
xnor U2209 (N_2209,N_328,N_1248);
xor U2210 (N_2210,N_795,N_1140);
xor U2211 (N_2211,N_387,N_978);
nand U2212 (N_2212,N_466,N_1196);
nor U2213 (N_2213,N_6,N_436);
or U2214 (N_2214,N_549,N_859);
nor U2215 (N_2215,N_482,N_1034);
nand U2216 (N_2216,N_783,N_1064);
xnor U2217 (N_2217,N_62,N_407);
nand U2218 (N_2218,N_1112,N_1110);
xnor U2219 (N_2219,N_874,N_1184);
nor U2220 (N_2220,N_798,N_614);
or U2221 (N_2221,N_891,N_793);
nor U2222 (N_2222,N_1209,N_1098);
nand U2223 (N_2223,N_300,N_787);
or U2224 (N_2224,N_65,N_239);
nor U2225 (N_2225,N_647,N_6);
nor U2226 (N_2226,N_151,N_737);
and U2227 (N_2227,N_627,N_829);
xnor U2228 (N_2228,N_1149,N_1109);
xnor U2229 (N_2229,N_408,N_409);
and U2230 (N_2230,N_737,N_422);
xnor U2231 (N_2231,N_728,N_461);
nor U2232 (N_2232,N_249,N_340);
or U2233 (N_2233,N_770,N_469);
xnor U2234 (N_2234,N_884,N_399);
nor U2235 (N_2235,N_1235,N_145);
xnor U2236 (N_2236,N_207,N_1069);
and U2237 (N_2237,N_1053,N_897);
xor U2238 (N_2238,N_894,N_502);
nand U2239 (N_2239,N_665,N_215);
or U2240 (N_2240,N_651,N_831);
xor U2241 (N_2241,N_175,N_1036);
and U2242 (N_2242,N_89,N_92);
nand U2243 (N_2243,N_1191,N_436);
and U2244 (N_2244,N_95,N_704);
nand U2245 (N_2245,N_503,N_1018);
nor U2246 (N_2246,N_723,N_390);
nand U2247 (N_2247,N_763,N_1087);
or U2248 (N_2248,N_391,N_931);
and U2249 (N_2249,N_299,N_784);
or U2250 (N_2250,N_775,N_439);
or U2251 (N_2251,N_644,N_772);
nor U2252 (N_2252,N_889,N_1031);
or U2253 (N_2253,N_71,N_367);
xnor U2254 (N_2254,N_808,N_1181);
nand U2255 (N_2255,N_1060,N_1194);
or U2256 (N_2256,N_337,N_84);
nand U2257 (N_2257,N_446,N_1177);
or U2258 (N_2258,N_628,N_1147);
nor U2259 (N_2259,N_989,N_324);
and U2260 (N_2260,N_988,N_993);
and U2261 (N_2261,N_201,N_594);
and U2262 (N_2262,N_141,N_500);
nand U2263 (N_2263,N_344,N_1048);
and U2264 (N_2264,N_1096,N_1032);
xnor U2265 (N_2265,N_958,N_807);
xnor U2266 (N_2266,N_888,N_341);
xnor U2267 (N_2267,N_911,N_674);
and U2268 (N_2268,N_372,N_519);
nand U2269 (N_2269,N_469,N_53);
nor U2270 (N_2270,N_930,N_364);
nor U2271 (N_2271,N_377,N_81);
or U2272 (N_2272,N_306,N_505);
and U2273 (N_2273,N_1181,N_277);
nor U2274 (N_2274,N_1027,N_1026);
and U2275 (N_2275,N_655,N_149);
xnor U2276 (N_2276,N_820,N_816);
and U2277 (N_2277,N_1117,N_543);
or U2278 (N_2278,N_233,N_1058);
and U2279 (N_2279,N_264,N_529);
or U2280 (N_2280,N_540,N_865);
nand U2281 (N_2281,N_1,N_683);
nand U2282 (N_2282,N_82,N_938);
nand U2283 (N_2283,N_442,N_1169);
xor U2284 (N_2284,N_992,N_555);
nor U2285 (N_2285,N_520,N_977);
and U2286 (N_2286,N_202,N_686);
nand U2287 (N_2287,N_149,N_1220);
or U2288 (N_2288,N_588,N_704);
and U2289 (N_2289,N_602,N_75);
and U2290 (N_2290,N_501,N_75);
and U2291 (N_2291,N_491,N_478);
and U2292 (N_2292,N_613,N_287);
and U2293 (N_2293,N_202,N_631);
and U2294 (N_2294,N_672,N_1030);
and U2295 (N_2295,N_150,N_1055);
and U2296 (N_2296,N_702,N_911);
xor U2297 (N_2297,N_830,N_659);
or U2298 (N_2298,N_296,N_876);
nand U2299 (N_2299,N_800,N_1048);
nand U2300 (N_2300,N_1180,N_562);
nand U2301 (N_2301,N_1116,N_353);
or U2302 (N_2302,N_623,N_430);
xnor U2303 (N_2303,N_656,N_789);
nor U2304 (N_2304,N_933,N_224);
nand U2305 (N_2305,N_215,N_202);
or U2306 (N_2306,N_1186,N_394);
or U2307 (N_2307,N_281,N_301);
nor U2308 (N_2308,N_163,N_1186);
nand U2309 (N_2309,N_1173,N_140);
or U2310 (N_2310,N_455,N_788);
or U2311 (N_2311,N_432,N_728);
nand U2312 (N_2312,N_652,N_130);
nor U2313 (N_2313,N_407,N_1071);
or U2314 (N_2314,N_1190,N_227);
nor U2315 (N_2315,N_1202,N_575);
nor U2316 (N_2316,N_305,N_694);
nor U2317 (N_2317,N_1108,N_559);
nor U2318 (N_2318,N_324,N_877);
nand U2319 (N_2319,N_200,N_1246);
and U2320 (N_2320,N_696,N_191);
nand U2321 (N_2321,N_52,N_105);
nor U2322 (N_2322,N_1132,N_20);
or U2323 (N_2323,N_492,N_614);
or U2324 (N_2324,N_921,N_493);
or U2325 (N_2325,N_775,N_874);
and U2326 (N_2326,N_428,N_651);
or U2327 (N_2327,N_523,N_650);
nand U2328 (N_2328,N_670,N_861);
xor U2329 (N_2329,N_311,N_166);
xnor U2330 (N_2330,N_652,N_1099);
nor U2331 (N_2331,N_612,N_464);
nand U2332 (N_2332,N_541,N_1164);
or U2333 (N_2333,N_588,N_47);
or U2334 (N_2334,N_1130,N_869);
xnor U2335 (N_2335,N_744,N_20);
nor U2336 (N_2336,N_692,N_535);
nand U2337 (N_2337,N_523,N_178);
xnor U2338 (N_2338,N_542,N_906);
nor U2339 (N_2339,N_1200,N_1073);
or U2340 (N_2340,N_595,N_96);
or U2341 (N_2341,N_15,N_116);
and U2342 (N_2342,N_389,N_70);
and U2343 (N_2343,N_668,N_153);
nor U2344 (N_2344,N_949,N_1079);
and U2345 (N_2345,N_1008,N_440);
or U2346 (N_2346,N_102,N_214);
nand U2347 (N_2347,N_149,N_746);
nand U2348 (N_2348,N_1209,N_759);
xnor U2349 (N_2349,N_441,N_298);
xnor U2350 (N_2350,N_964,N_6);
and U2351 (N_2351,N_16,N_224);
xnor U2352 (N_2352,N_1155,N_1204);
or U2353 (N_2353,N_51,N_85);
nor U2354 (N_2354,N_35,N_979);
or U2355 (N_2355,N_1205,N_103);
nand U2356 (N_2356,N_1115,N_727);
xnor U2357 (N_2357,N_690,N_613);
or U2358 (N_2358,N_498,N_261);
xnor U2359 (N_2359,N_243,N_167);
nor U2360 (N_2360,N_319,N_1189);
nand U2361 (N_2361,N_683,N_1035);
nand U2362 (N_2362,N_727,N_742);
xnor U2363 (N_2363,N_399,N_162);
or U2364 (N_2364,N_310,N_713);
or U2365 (N_2365,N_1224,N_1019);
xnor U2366 (N_2366,N_992,N_652);
and U2367 (N_2367,N_958,N_1177);
or U2368 (N_2368,N_925,N_961);
or U2369 (N_2369,N_493,N_937);
xor U2370 (N_2370,N_644,N_948);
xnor U2371 (N_2371,N_1058,N_585);
nand U2372 (N_2372,N_658,N_1220);
xnor U2373 (N_2373,N_270,N_129);
and U2374 (N_2374,N_667,N_527);
nand U2375 (N_2375,N_503,N_1021);
and U2376 (N_2376,N_947,N_1244);
xnor U2377 (N_2377,N_474,N_991);
xor U2378 (N_2378,N_927,N_1245);
and U2379 (N_2379,N_516,N_542);
and U2380 (N_2380,N_1006,N_1030);
and U2381 (N_2381,N_485,N_781);
and U2382 (N_2382,N_771,N_16);
nor U2383 (N_2383,N_314,N_926);
nand U2384 (N_2384,N_1056,N_623);
and U2385 (N_2385,N_136,N_1148);
nand U2386 (N_2386,N_197,N_720);
xor U2387 (N_2387,N_417,N_0);
nor U2388 (N_2388,N_1223,N_69);
xnor U2389 (N_2389,N_127,N_606);
or U2390 (N_2390,N_776,N_534);
or U2391 (N_2391,N_476,N_646);
nand U2392 (N_2392,N_215,N_1107);
nor U2393 (N_2393,N_1188,N_1047);
or U2394 (N_2394,N_959,N_1050);
and U2395 (N_2395,N_334,N_615);
and U2396 (N_2396,N_792,N_476);
nor U2397 (N_2397,N_643,N_469);
and U2398 (N_2398,N_892,N_819);
or U2399 (N_2399,N_341,N_610);
nor U2400 (N_2400,N_694,N_871);
xnor U2401 (N_2401,N_1129,N_1016);
nor U2402 (N_2402,N_983,N_443);
nor U2403 (N_2403,N_894,N_407);
nor U2404 (N_2404,N_107,N_440);
xnor U2405 (N_2405,N_322,N_693);
and U2406 (N_2406,N_700,N_286);
xnor U2407 (N_2407,N_676,N_702);
and U2408 (N_2408,N_173,N_677);
or U2409 (N_2409,N_55,N_1019);
and U2410 (N_2410,N_1043,N_141);
or U2411 (N_2411,N_1108,N_199);
or U2412 (N_2412,N_165,N_462);
nand U2413 (N_2413,N_40,N_569);
xnor U2414 (N_2414,N_1226,N_1004);
nor U2415 (N_2415,N_823,N_832);
xnor U2416 (N_2416,N_1023,N_188);
nand U2417 (N_2417,N_731,N_539);
and U2418 (N_2418,N_274,N_629);
nor U2419 (N_2419,N_458,N_183);
and U2420 (N_2420,N_718,N_652);
nor U2421 (N_2421,N_874,N_357);
and U2422 (N_2422,N_970,N_352);
and U2423 (N_2423,N_195,N_40);
nand U2424 (N_2424,N_1156,N_824);
xor U2425 (N_2425,N_504,N_804);
nor U2426 (N_2426,N_583,N_639);
xor U2427 (N_2427,N_384,N_494);
nand U2428 (N_2428,N_555,N_780);
and U2429 (N_2429,N_264,N_234);
nand U2430 (N_2430,N_830,N_965);
or U2431 (N_2431,N_597,N_387);
and U2432 (N_2432,N_873,N_202);
or U2433 (N_2433,N_657,N_199);
xnor U2434 (N_2434,N_592,N_897);
or U2435 (N_2435,N_331,N_599);
nor U2436 (N_2436,N_956,N_832);
and U2437 (N_2437,N_257,N_376);
or U2438 (N_2438,N_840,N_974);
xnor U2439 (N_2439,N_512,N_686);
or U2440 (N_2440,N_1164,N_638);
nand U2441 (N_2441,N_321,N_40);
nor U2442 (N_2442,N_245,N_824);
or U2443 (N_2443,N_357,N_1064);
or U2444 (N_2444,N_410,N_353);
and U2445 (N_2445,N_243,N_509);
xnor U2446 (N_2446,N_1172,N_22);
nor U2447 (N_2447,N_331,N_273);
nand U2448 (N_2448,N_653,N_347);
and U2449 (N_2449,N_683,N_907);
nand U2450 (N_2450,N_800,N_597);
nor U2451 (N_2451,N_907,N_895);
nor U2452 (N_2452,N_975,N_1100);
xnor U2453 (N_2453,N_696,N_1240);
or U2454 (N_2454,N_291,N_132);
or U2455 (N_2455,N_847,N_621);
xor U2456 (N_2456,N_1138,N_647);
or U2457 (N_2457,N_71,N_1183);
nand U2458 (N_2458,N_216,N_597);
xnor U2459 (N_2459,N_1247,N_198);
or U2460 (N_2460,N_731,N_790);
and U2461 (N_2461,N_707,N_855);
nand U2462 (N_2462,N_363,N_408);
nor U2463 (N_2463,N_753,N_1000);
and U2464 (N_2464,N_210,N_196);
nand U2465 (N_2465,N_872,N_888);
nor U2466 (N_2466,N_513,N_989);
nand U2467 (N_2467,N_840,N_115);
nand U2468 (N_2468,N_225,N_604);
nor U2469 (N_2469,N_722,N_50);
xnor U2470 (N_2470,N_862,N_160);
nor U2471 (N_2471,N_242,N_311);
and U2472 (N_2472,N_816,N_1232);
nand U2473 (N_2473,N_49,N_501);
or U2474 (N_2474,N_864,N_1247);
and U2475 (N_2475,N_413,N_649);
and U2476 (N_2476,N_245,N_571);
nor U2477 (N_2477,N_724,N_539);
nand U2478 (N_2478,N_968,N_398);
or U2479 (N_2479,N_357,N_753);
and U2480 (N_2480,N_497,N_547);
nand U2481 (N_2481,N_523,N_155);
and U2482 (N_2482,N_467,N_861);
or U2483 (N_2483,N_243,N_216);
and U2484 (N_2484,N_32,N_439);
nand U2485 (N_2485,N_853,N_586);
nand U2486 (N_2486,N_210,N_605);
and U2487 (N_2487,N_157,N_683);
nor U2488 (N_2488,N_35,N_324);
or U2489 (N_2489,N_181,N_640);
and U2490 (N_2490,N_551,N_1131);
and U2491 (N_2491,N_860,N_1205);
and U2492 (N_2492,N_379,N_787);
and U2493 (N_2493,N_150,N_849);
xor U2494 (N_2494,N_872,N_324);
nor U2495 (N_2495,N_435,N_690);
xor U2496 (N_2496,N_18,N_583);
nand U2497 (N_2497,N_16,N_1156);
nand U2498 (N_2498,N_1248,N_1008);
or U2499 (N_2499,N_1175,N_1209);
xnor U2500 (N_2500,N_1701,N_1584);
and U2501 (N_2501,N_2009,N_2342);
nor U2502 (N_2502,N_2313,N_2394);
xor U2503 (N_2503,N_2455,N_2215);
nor U2504 (N_2504,N_1453,N_2475);
xnor U2505 (N_2505,N_1960,N_2037);
nand U2506 (N_2506,N_1900,N_1927);
and U2507 (N_2507,N_1355,N_1688);
and U2508 (N_2508,N_2376,N_2349);
xnor U2509 (N_2509,N_1503,N_2270);
nand U2510 (N_2510,N_2237,N_1567);
and U2511 (N_2511,N_2072,N_1597);
and U2512 (N_2512,N_2295,N_1410);
nand U2513 (N_2513,N_1865,N_1862);
xnor U2514 (N_2514,N_2188,N_2207);
nor U2515 (N_2515,N_2061,N_1808);
or U2516 (N_2516,N_2102,N_1450);
nand U2517 (N_2517,N_1792,N_2269);
nand U2518 (N_2518,N_2384,N_1649);
nor U2519 (N_2519,N_1756,N_2016);
nor U2520 (N_2520,N_1580,N_2370);
nand U2521 (N_2521,N_2348,N_2010);
xor U2522 (N_2522,N_1318,N_1325);
and U2523 (N_2523,N_1434,N_1754);
nor U2524 (N_2524,N_1314,N_1544);
or U2525 (N_2525,N_1476,N_1295);
and U2526 (N_2526,N_1441,N_1819);
nand U2527 (N_2527,N_1652,N_1802);
nand U2528 (N_2528,N_1704,N_1677);
nor U2529 (N_2529,N_2329,N_2162);
or U2530 (N_2530,N_1381,N_1499);
or U2531 (N_2531,N_2323,N_2347);
or U2532 (N_2532,N_1391,N_2052);
nor U2533 (N_2533,N_1257,N_1897);
nand U2534 (N_2534,N_2488,N_2400);
and U2535 (N_2535,N_1501,N_2148);
and U2536 (N_2536,N_1903,N_2195);
or U2537 (N_2537,N_1455,N_1870);
or U2538 (N_2538,N_1273,N_1623);
and U2539 (N_2539,N_2135,N_1626);
nor U2540 (N_2540,N_2401,N_2180);
nor U2541 (N_2541,N_1342,N_2186);
xnor U2542 (N_2542,N_2065,N_1463);
xor U2543 (N_2543,N_2049,N_2314);
xor U2544 (N_2544,N_2276,N_1738);
nor U2545 (N_2545,N_1469,N_1599);
and U2546 (N_2546,N_1291,N_2469);
and U2547 (N_2547,N_1685,N_1470);
or U2548 (N_2548,N_1497,N_1407);
and U2549 (N_2549,N_1696,N_1912);
xor U2550 (N_2550,N_2247,N_1561);
and U2551 (N_2551,N_1727,N_1767);
nand U2552 (N_2552,N_2260,N_1687);
xor U2553 (N_2553,N_2422,N_1262);
xor U2554 (N_2554,N_2234,N_2092);
and U2555 (N_2555,N_2147,N_2075);
nor U2556 (N_2556,N_2317,N_1421);
or U2557 (N_2557,N_1397,N_1762);
or U2558 (N_2558,N_1486,N_1904);
nor U2559 (N_2559,N_1574,N_1471);
and U2560 (N_2560,N_1929,N_1986);
or U2561 (N_2561,N_1483,N_1582);
nand U2562 (N_2562,N_2334,N_2132);
nand U2563 (N_2563,N_1964,N_2179);
nor U2564 (N_2564,N_1684,N_1285);
or U2565 (N_2565,N_1809,N_2425);
nor U2566 (N_2566,N_2171,N_1746);
nand U2567 (N_2567,N_1898,N_1866);
xor U2568 (N_2568,N_1399,N_2372);
nand U2569 (N_2569,N_1308,N_1581);
or U2570 (N_2570,N_1653,N_2141);
and U2571 (N_2571,N_1348,N_1961);
nand U2572 (N_2572,N_1735,N_1474);
and U2573 (N_2573,N_2249,N_1818);
nand U2574 (N_2574,N_2453,N_1915);
xnor U2575 (N_2575,N_1911,N_2096);
nor U2576 (N_2576,N_2273,N_1997);
and U2577 (N_2577,N_1692,N_2434);
nor U2578 (N_2578,N_1343,N_2373);
xor U2579 (N_2579,N_1557,N_1758);
nor U2580 (N_2580,N_2145,N_1628);
and U2581 (N_2581,N_1608,N_2446);
and U2582 (N_2582,N_2198,N_2278);
nand U2583 (N_2583,N_1783,N_1265);
and U2584 (N_2584,N_1383,N_1660);
xnor U2585 (N_2585,N_1366,N_1617);
or U2586 (N_2586,N_1297,N_1467);
xnor U2587 (N_2587,N_2417,N_1596);
and U2588 (N_2588,N_1806,N_1392);
and U2589 (N_2589,N_2374,N_1959);
and U2590 (N_2590,N_1638,N_2082);
nor U2591 (N_2591,N_2390,N_2003);
and U2592 (N_2592,N_1991,N_1344);
xnor U2593 (N_2593,N_1675,N_1769);
or U2594 (N_2594,N_2029,N_2134);
nor U2595 (N_2595,N_2078,N_1686);
nor U2596 (N_2596,N_1500,N_1951);
xor U2597 (N_2597,N_1872,N_2181);
and U2598 (N_2598,N_2210,N_1620);
nand U2599 (N_2599,N_1569,N_1251);
and U2600 (N_2600,N_2345,N_2059);
nor U2601 (N_2601,N_2423,N_1989);
xnor U2602 (N_2602,N_1563,N_2055);
and U2603 (N_2603,N_2025,N_1274);
or U2604 (N_2604,N_2456,N_1869);
nor U2605 (N_2605,N_1311,N_2333);
nor U2606 (N_2606,N_1349,N_1428);
nand U2607 (N_2607,N_2355,N_1836);
and U2608 (N_2608,N_1863,N_1408);
nand U2609 (N_2609,N_1981,N_2150);
nor U2610 (N_2610,N_1554,N_2245);
or U2611 (N_2611,N_2362,N_1970);
xnor U2612 (N_2612,N_2438,N_1681);
and U2613 (N_2613,N_1666,N_2033);
nor U2614 (N_2614,N_1782,N_1713);
nor U2615 (N_2615,N_2442,N_1846);
xor U2616 (N_2616,N_1683,N_1590);
and U2617 (N_2617,N_2375,N_2080);
nand U2618 (N_2618,N_1533,N_2208);
and U2619 (N_2619,N_1549,N_1320);
xnor U2620 (N_2620,N_1542,N_2077);
nand U2621 (N_2621,N_1445,N_2214);
or U2622 (N_2622,N_1941,N_2060);
or U2623 (N_2623,N_2243,N_1920);
or U2624 (N_2624,N_2309,N_2470);
or U2625 (N_2625,N_1859,N_2084);
xnor U2626 (N_2626,N_1322,N_1966);
nand U2627 (N_2627,N_1256,N_1531);
nor U2628 (N_2628,N_2499,N_1665);
xnor U2629 (N_2629,N_2023,N_1613);
xnor U2630 (N_2630,N_1824,N_1437);
and U2631 (N_2631,N_2290,N_2152);
and U2632 (N_2632,N_2086,N_2129);
or U2633 (N_2633,N_1269,N_1301);
nand U2634 (N_2634,N_1556,N_1460);
xnor U2635 (N_2635,N_1546,N_1456);
xor U2636 (N_2636,N_1919,N_1275);
nor U2637 (N_2637,N_1481,N_1370);
nand U2638 (N_2638,N_1384,N_2272);
nand U2639 (N_2639,N_1327,N_1926);
nand U2640 (N_2640,N_1700,N_1910);
nor U2641 (N_2641,N_2350,N_1404);
nor U2642 (N_2642,N_2196,N_1536);
nor U2643 (N_2643,N_1454,N_1588);
and U2644 (N_2644,N_1740,N_2358);
xor U2645 (N_2645,N_2182,N_2250);
or U2646 (N_2646,N_1770,N_2439);
nand U2647 (N_2647,N_1300,N_2451);
nor U2648 (N_2648,N_1832,N_1726);
nand U2649 (N_2649,N_2039,N_2218);
xnor U2650 (N_2650,N_1253,N_2274);
or U2651 (N_2651,N_1933,N_2353);
or U2652 (N_2652,N_2450,N_1893);
or U2653 (N_2653,N_2087,N_2476);
nand U2654 (N_2654,N_2429,N_2232);
nand U2655 (N_2655,N_1373,N_1350);
and U2656 (N_2656,N_1992,N_2261);
nand U2657 (N_2657,N_1988,N_1861);
xnor U2658 (N_2658,N_1447,N_1337);
nor U2659 (N_2659,N_1579,N_1644);
and U2660 (N_2660,N_1952,N_2103);
nor U2661 (N_2661,N_2254,N_1401);
and U2662 (N_2662,N_2011,N_2346);
nor U2663 (N_2663,N_1415,N_1993);
or U2664 (N_2664,N_1379,N_1939);
and U2665 (N_2665,N_1716,N_2448);
nor U2666 (N_2666,N_1489,N_1829);
and U2667 (N_2667,N_1303,N_2480);
nor U2668 (N_2668,N_1418,N_1833);
nor U2669 (N_2669,N_2263,N_2027);
and U2670 (N_2670,N_1795,N_2296);
nor U2671 (N_2671,N_1361,N_2287);
and U2672 (N_2672,N_1414,N_2233);
or U2673 (N_2673,N_2322,N_2357);
nand U2674 (N_2674,N_1494,N_1572);
or U2675 (N_2675,N_1508,N_2127);
and U2676 (N_2676,N_1413,N_2465);
and U2677 (N_2677,N_2415,N_2185);
or U2678 (N_2678,N_1743,N_2304);
and U2679 (N_2679,N_1945,N_1778);
nor U2680 (N_2680,N_2026,N_1834);
and U2681 (N_2681,N_1287,N_2340);
nor U2682 (N_2682,N_2221,N_1280);
or U2683 (N_2683,N_1510,N_1896);
or U2684 (N_2684,N_1635,N_1412);
nor U2685 (N_2685,N_2155,N_2191);
nor U2686 (N_2686,N_2256,N_2089);
and U2687 (N_2687,N_2280,N_1310);
nand U2688 (N_2688,N_2497,N_1409);
nand U2689 (N_2689,N_2163,N_1516);
nor U2690 (N_2690,N_1736,N_2165);
nor U2691 (N_2691,N_1715,N_1458);
xnor U2692 (N_2692,N_1942,N_2231);
and U2693 (N_2693,N_2397,N_2380);
nor U2694 (N_2694,N_1258,N_1312);
nor U2695 (N_2695,N_1761,N_1600);
or U2696 (N_2696,N_1321,N_2461);
xor U2697 (N_2697,N_1977,N_1934);
or U2698 (N_2698,N_1403,N_2140);
nor U2699 (N_2699,N_2217,N_1267);
nand U2700 (N_2700,N_1566,N_2020);
nand U2701 (N_2701,N_1520,N_1847);
nand U2702 (N_2702,N_1438,N_1794);
nor U2703 (N_2703,N_2169,N_2408);
and U2704 (N_2704,N_1659,N_2064);
and U2705 (N_2705,N_1773,N_1757);
nor U2706 (N_2706,N_2143,N_1969);
or U2707 (N_2707,N_2090,N_1521);
xor U2708 (N_2708,N_2406,N_1805);
xor U2709 (N_2709,N_1302,N_1967);
or U2710 (N_2710,N_1750,N_1540);
or U2711 (N_2711,N_2000,N_2354);
nand U2712 (N_2712,N_2298,N_1957);
and U2713 (N_2713,N_1739,N_1797);
nand U2714 (N_2714,N_2382,N_1576);
nor U2715 (N_2715,N_1680,N_2288);
xor U2716 (N_2716,N_2359,N_2149);
xnor U2717 (N_2717,N_1282,N_1822);
or U2718 (N_2718,N_1424,N_2428);
nor U2719 (N_2719,N_1877,N_1845);
or U2720 (N_2720,N_2111,N_2454);
nand U2721 (N_2721,N_1667,N_1645);
nor U2722 (N_2722,N_1543,N_2071);
or U2723 (N_2723,N_1266,N_1914);
nor U2724 (N_2724,N_2032,N_1947);
or U2725 (N_2725,N_2105,N_1316);
nand U2726 (N_2726,N_1524,N_1884);
nor U2727 (N_2727,N_2205,N_2458);
nor U2728 (N_2728,N_2431,N_1980);
and U2729 (N_2729,N_1615,N_2467);
nor U2730 (N_2730,N_2115,N_2413);
and U2731 (N_2731,N_1416,N_1760);
or U2732 (N_2732,N_1385,N_2161);
or U2733 (N_2733,N_1525,N_1948);
nand U2734 (N_2734,N_1710,N_1785);
nand U2735 (N_2735,N_1643,N_2410);
and U2736 (N_2736,N_1843,N_1772);
xor U2737 (N_2737,N_1374,N_2293);
xnor U2738 (N_2738,N_2216,N_1363);
xnor U2739 (N_2739,N_2447,N_1857);
nand U2740 (N_2740,N_1537,N_2030);
or U2741 (N_2741,N_2483,N_1364);
nand U2742 (N_2742,N_1706,N_1395);
xor U2743 (N_2743,N_1780,N_2318);
xnor U2744 (N_2744,N_2241,N_1842);
and U2745 (N_2745,N_2219,N_1490);
or U2746 (N_2746,N_2178,N_1526);
nand U2747 (N_2747,N_2076,N_1250);
nor U2748 (N_2748,N_1488,N_2002);
and U2749 (N_2749,N_1585,N_1281);
xnor U2750 (N_2750,N_2445,N_1478);
or U2751 (N_2751,N_1766,N_2238);
xnor U2752 (N_2752,N_1317,N_1850);
or U2753 (N_2753,N_1816,N_1786);
nor U2754 (N_2754,N_1506,N_1365);
nand U2755 (N_2755,N_1858,N_1646);
or U2756 (N_2756,N_2267,N_2282);
nand U2757 (N_2757,N_2262,N_2053);
or U2758 (N_2758,N_2042,N_1286);
or U2759 (N_2759,N_1283,N_1296);
nand U2760 (N_2760,N_1922,N_2137);
nand U2761 (N_2761,N_2266,N_1514);
and U2762 (N_2762,N_1662,N_1278);
nand U2763 (N_2763,N_1380,N_2139);
nand U2764 (N_2764,N_1360,N_2404);
nand U2765 (N_2765,N_1732,N_1661);
and U2766 (N_2766,N_2062,N_2441);
xor U2767 (N_2767,N_1930,N_1351);
or U2768 (N_2768,N_2389,N_2063);
nand U2769 (N_2769,N_2268,N_1553);
nand U2770 (N_2770,N_1633,N_1570);
or U2771 (N_2771,N_1482,N_1871);
nand U2772 (N_2772,N_1329,N_1636);
nand U2773 (N_2773,N_2478,N_1372);
xnor U2774 (N_2774,N_1509,N_1528);
xnor U2775 (N_2775,N_1552,N_1603);
nand U2776 (N_2776,N_1362,N_2324);
or U2777 (N_2777,N_2393,N_1548);
xor U2778 (N_2778,N_1431,N_1901);
nor U2779 (N_2779,N_1341,N_1465);
nor U2780 (N_2780,N_2183,N_2363);
xnor U2781 (N_2781,N_1963,N_2204);
nand U2782 (N_2782,N_1887,N_1810);
xnor U2783 (N_2783,N_2133,N_1932);
and U2784 (N_2784,N_1284,N_1304);
or U2785 (N_2785,N_1880,N_2074);
or U2786 (N_2786,N_2112,N_1731);
and U2787 (N_2787,N_2440,N_2106);
or U2788 (N_2788,N_2321,N_1535);
nand U2789 (N_2789,N_1909,N_1504);
nor U2790 (N_2790,N_1356,N_2083);
and U2791 (N_2791,N_2407,N_2457);
and U2792 (N_2792,N_2437,N_1711);
and U2793 (N_2793,N_1511,N_1522);
or U2794 (N_2794,N_2176,N_2302);
and U2795 (N_2795,N_1464,N_1689);
and U2796 (N_2796,N_1650,N_1496);
nand U2797 (N_2797,N_1475,N_1604);
or U2798 (N_2798,N_2405,N_2303);
nor U2799 (N_2799,N_2203,N_2160);
nor U2800 (N_2800,N_2279,N_1378);
nand U2801 (N_2801,N_2398,N_1899);
nand U2802 (N_2802,N_2367,N_2166);
xnor U2803 (N_2803,N_2197,N_2436);
xor U2804 (N_2804,N_1624,N_2396);
nand U2805 (N_2805,N_1678,N_2482);
or U2806 (N_2806,N_1825,N_2312);
nand U2807 (N_2807,N_1622,N_2144);
or U2808 (N_2808,N_2158,N_1357);
or U2809 (N_2809,N_1427,N_1639);
nand U2810 (N_2810,N_2184,N_1443);
or U2811 (N_2811,N_2311,N_2008);
nor U2812 (N_2812,N_2122,N_1406);
nand U2813 (N_2813,N_1294,N_1734);
or U2814 (N_2814,N_2294,N_1821);
nor U2815 (N_2815,N_1916,N_1405);
and U2816 (N_2816,N_2067,N_2388);
or U2817 (N_2817,N_1493,N_1505);
or U2818 (N_2818,N_2047,N_2048);
xor U2819 (N_2819,N_1601,N_2043);
xor U2820 (N_2820,N_2200,N_2173);
nand U2821 (N_2821,N_2138,N_2369);
xor U2822 (N_2822,N_2007,N_2494);
or U2823 (N_2823,N_1545,N_1400);
nand U2824 (N_2824,N_2190,N_1690);
and U2825 (N_2825,N_2131,N_1745);
or U2826 (N_2826,N_2069,N_2386);
nand U2827 (N_2827,N_2125,N_1562);
nand U2828 (N_2828,N_1324,N_2473);
nand U2829 (N_2829,N_2113,N_1479);
or U2830 (N_2830,N_1512,N_2325);
nand U2831 (N_2831,N_1423,N_1461);
nand U2832 (N_2832,N_1358,N_1254);
nand U2833 (N_2833,N_2236,N_2330);
or U2834 (N_2834,N_2174,N_2194);
or U2835 (N_2835,N_1800,N_2360);
nor U2836 (N_2836,N_2319,N_1532);
and U2837 (N_2837,N_1936,N_1837);
or U2838 (N_2838,N_1823,N_2253);
or U2839 (N_2839,N_1729,N_2057);
nand U2840 (N_2840,N_1527,N_1885);
nand U2841 (N_2841,N_2104,N_2391);
xor U2842 (N_2842,N_2109,N_1515);
xor U2843 (N_2843,N_1741,N_1326);
nor U2844 (N_2844,N_1831,N_1679);
xor U2845 (N_2845,N_1550,N_2046);
nand U2846 (N_2846,N_1717,N_1937);
nor U2847 (N_2847,N_1938,N_1425);
and U2848 (N_2848,N_1630,N_1737);
and U2849 (N_2849,N_2284,N_1663);
and U2850 (N_2850,N_2202,N_2193);
xnor U2851 (N_2851,N_2220,N_1398);
nand U2852 (N_2852,N_1820,N_1656);
nand U2853 (N_2853,N_2044,N_2275);
or U2854 (N_2854,N_1640,N_2433);
nor U2855 (N_2855,N_1905,N_2452);
nand U2856 (N_2856,N_1347,N_1519);
nor U2857 (N_2857,N_2310,N_1671);
and U2858 (N_2858,N_1634,N_1733);
nand U2859 (N_2859,N_1676,N_2005);
and U2860 (N_2860,N_1855,N_2299);
or U2861 (N_2861,N_1707,N_2306);
nand U2862 (N_2862,N_1340,N_1587);
or U2863 (N_2863,N_2130,N_1518);
and U2864 (N_2864,N_1974,N_1720);
nand U2865 (N_2865,N_1730,N_2056);
and U2866 (N_2866,N_1309,N_1804);
nor U2867 (N_2867,N_2093,N_2305);
or U2868 (N_2868,N_1728,N_1568);
nand U2869 (N_2869,N_2251,N_1387);
and U2870 (N_2870,N_1573,N_2107);
xor U2871 (N_2871,N_2301,N_1807);
or U2872 (N_2872,N_1339,N_1641);
nor U2873 (N_2873,N_2320,N_1994);
or U2874 (N_2874,N_2153,N_1288);
nor U2875 (N_2875,N_1946,N_2259);
nand U2876 (N_2876,N_1313,N_1695);
nand U2877 (N_2877,N_1925,N_1459);
nand U2878 (N_2878,N_1259,N_1614);
or U2879 (N_2879,N_2051,N_2013);
or U2880 (N_2880,N_1978,N_2019);
or U2881 (N_2881,N_1606,N_2432);
nor U2882 (N_2882,N_2209,N_1674);
nand U2883 (N_2883,N_2399,N_1979);
and U2884 (N_2884,N_2403,N_1375);
nor U2885 (N_2885,N_1529,N_1699);
or U2886 (N_2886,N_2164,N_1955);
and U2887 (N_2887,N_2477,N_1975);
nor U2888 (N_2888,N_1530,N_1513);
xor U2889 (N_2889,N_2490,N_2351);
nand U2890 (N_2890,N_1890,N_1703);
xor U2891 (N_2891,N_2421,N_1902);
nor U2892 (N_2892,N_1457,N_2230);
nand U2893 (N_2893,N_1473,N_2240);
or U2894 (N_2894,N_1801,N_1605);
nand U2895 (N_2895,N_1996,N_2392);
nand U2896 (N_2896,N_2227,N_1466);
or U2897 (N_2897,N_2239,N_2341);
and U2898 (N_2898,N_2085,N_2366);
nor U2899 (N_2899,N_1787,N_1878);
or U2900 (N_2900,N_2206,N_1323);
xor U2901 (N_2901,N_2229,N_2485);
nor U2902 (N_2902,N_2021,N_1971);
or U2903 (N_2903,N_2094,N_1875);
nor U2904 (N_2904,N_1538,N_1272);
xor U2905 (N_2905,N_1393,N_1389);
nand U2906 (N_2906,N_2189,N_1263);
xnor U2907 (N_2907,N_2308,N_1376);
or U2908 (N_2908,N_2379,N_2123);
nand U2909 (N_2909,N_1709,N_1779);
nand U2910 (N_2910,N_2471,N_2024);
nand U2911 (N_2911,N_2170,N_1571);
xor U2912 (N_2912,N_1973,N_1771);
nand U2913 (N_2913,N_1983,N_2242);
or U2914 (N_2914,N_2419,N_2081);
or U2915 (N_2915,N_2427,N_1592);
or U2916 (N_2916,N_2248,N_2058);
xor U2917 (N_2917,N_1371,N_1669);
and U2918 (N_2918,N_2283,N_1551);
nand U2919 (N_2919,N_2383,N_1958);
nor U2920 (N_2920,N_1648,N_1565);
and U2921 (N_2921,N_1411,N_1923);
or U2922 (N_2922,N_2496,N_1906);
nor U2923 (N_2923,N_2336,N_1331);
xor U2924 (N_2924,N_1886,N_2255);
or U2925 (N_2925,N_1765,N_2142);
nor U2926 (N_2926,N_1867,N_1293);
or U2927 (N_2927,N_1485,N_1828);
xnor U2928 (N_2928,N_1985,N_1744);
xor U2929 (N_2929,N_2099,N_1682);
or U2930 (N_2930,N_1338,N_1480);
or U2931 (N_2931,N_1873,N_2120);
and U2932 (N_2932,N_1359,N_2402);
nor U2933 (N_2933,N_2121,N_1725);
and U2934 (N_2934,N_2371,N_2070);
and U2935 (N_2935,N_2339,N_1712);
nor U2936 (N_2936,N_1439,N_1555);
nand U2937 (N_2937,N_1432,N_1864);
nor U2938 (N_2938,N_1752,N_2378);
or U2939 (N_2939,N_1618,N_2377);
nor U2940 (N_2940,N_1435,N_1776);
or U2941 (N_2941,N_2332,N_2352);
nor U2942 (N_2942,N_2154,N_2264);
and U2943 (N_2943,N_2012,N_1367);
nor U2944 (N_2944,N_1523,N_1307);
and U2945 (N_2945,N_1722,N_2034);
nand U2946 (N_2946,N_2484,N_1813);
and U2947 (N_2947,N_2035,N_1451);
nand U2948 (N_2948,N_1446,N_1539);
nand U2949 (N_2949,N_2443,N_1305);
xnor U2950 (N_2950,N_2292,N_2326);
or U2951 (N_2951,N_1292,N_1382);
or U2952 (N_2952,N_1702,N_2411);
nor U2953 (N_2953,N_2156,N_2213);
xor U2954 (N_2954,N_1817,N_2412);
nand U2955 (N_2955,N_1444,N_2387);
nand U2956 (N_2956,N_2265,N_1962);
or U2957 (N_2957,N_1984,N_1724);
or U2958 (N_2958,N_1844,N_1330);
xor U2959 (N_2959,N_2118,N_2381);
and U2960 (N_2960,N_1260,N_1607);
nand U2961 (N_2961,N_1999,N_2199);
nand U2962 (N_2962,N_2416,N_1276);
and U2963 (N_2963,N_1995,N_1426);
and U2964 (N_2964,N_1698,N_1839);
or U2965 (N_2965,N_2449,N_2495);
or U2966 (N_2966,N_2110,N_2014);
or U2967 (N_2967,N_1277,N_1616);
xnor U2968 (N_2968,N_1642,N_2136);
and U2969 (N_2969,N_1507,N_2050);
nor U2970 (N_2970,N_1972,N_2328);
or U2971 (N_2971,N_1924,N_2430);
and U2972 (N_2972,N_1908,N_1793);
xnor U2973 (N_2973,N_2228,N_1315);
xor U2974 (N_2974,N_1838,N_1788);
or U2975 (N_2975,N_2338,N_1811);
and U2976 (N_2976,N_1586,N_1881);
nor U2977 (N_2977,N_1612,N_1851);
and U2978 (N_2978,N_2316,N_2068);
nand U2979 (N_2979,N_1940,N_1252);
xnor U2980 (N_2980,N_1815,N_1390);
and U2981 (N_2981,N_2491,N_2041);
nand U2982 (N_2982,N_2006,N_2117);
or U2983 (N_2983,N_2493,N_2444);
xnor U2984 (N_2984,N_1714,N_1593);
and U2985 (N_2985,N_2172,N_2435);
xor U2986 (N_2986,N_2418,N_1889);
xnor U2987 (N_2987,N_2225,N_1637);
nor U2988 (N_2988,N_1270,N_1595);
nor U2989 (N_2989,N_1377,N_2101);
nor U2990 (N_2990,N_2114,N_1882);
xnor U2991 (N_2991,N_1547,N_2466);
xnor U2992 (N_2992,N_1577,N_2054);
or U2993 (N_2993,N_1353,N_1827);
or U2994 (N_2994,N_1559,N_1928);
nand U2995 (N_2995,N_1935,N_2119);
or U2996 (N_2996,N_1796,N_1723);
or U2997 (N_2997,N_1417,N_2492);
and U2998 (N_2998,N_2414,N_1517);
or U2999 (N_2999,N_1468,N_1791);
nor U3000 (N_3000,N_1849,N_2331);
or U3001 (N_3001,N_1279,N_1271);
nor U3002 (N_3002,N_1747,N_1560);
nand U3003 (N_3003,N_2192,N_1261);
or U3004 (N_3004,N_2168,N_2022);
or U3005 (N_3005,N_1907,N_2116);
nor U3006 (N_3006,N_1462,N_1721);
or U3007 (N_3007,N_1610,N_1668);
nor U3008 (N_3008,N_1602,N_2286);
and U3009 (N_3009,N_2045,N_1830);
or U3010 (N_3010,N_1589,N_1386);
and U3011 (N_3011,N_1697,N_2157);
nand U3012 (N_3012,N_1621,N_2066);
or U3013 (N_3013,N_2424,N_1632);
xnor U3014 (N_3014,N_1789,N_2258);
or U3015 (N_3015,N_1672,N_2244);
and U3016 (N_3016,N_1954,N_2252);
or U3017 (N_3017,N_2126,N_2146);
nor U3018 (N_3018,N_2223,N_1670);
or U3019 (N_3019,N_2462,N_1965);
nor U3020 (N_3020,N_1658,N_1657);
and U3021 (N_3021,N_1883,N_1753);
or U3022 (N_3022,N_2420,N_1627);
nand U3023 (N_3023,N_2015,N_1647);
or U3024 (N_3024,N_1673,N_2004);
and U3025 (N_3025,N_1918,N_1448);
and U3026 (N_3026,N_2212,N_1429);
and U3027 (N_3027,N_1629,N_1611);
nor U3028 (N_3028,N_2175,N_1289);
nand U3029 (N_3029,N_1860,N_2343);
xor U3030 (N_3030,N_2327,N_1333);
nor U3031 (N_3031,N_2361,N_2285);
nor U3032 (N_3032,N_1748,N_2291);
nand U3033 (N_3033,N_1755,N_1298);
nor U3034 (N_3034,N_1691,N_2038);
nand U3035 (N_3035,N_1319,N_1953);
xnor U3036 (N_3036,N_2097,N_2211);
nor U3037 (N_3037,N_1345,N_1598);
xor U3038 (N_3038,N_1891,N_1472);
and U3039 (N_3039,N_2036,N_1264);
and U3040 (N_3040,N_2368,N_1826);
and U3041 (N_3041,N_2395,N_2486);
xor U3042 (N_3042,N_2001,N_1781);
or U3043 (N_3043,N_1768,N_1255);
nor U3044 (N_3044,N_1803,N_1575);
or U3045 (N_3045,N_1369,N_2464);
xor U3046 (N_3046,N_1895,N_1354);
nor U3047 (N_3047,N_2017,N_1694);
xor U3048 (N_3048,N_1835,N_2246);
nor U3049 (N_3049,N_1921,N_1759);
nor U3050 (N_3050,N_1874,N_2337);
and U3051 (N_3051,N_1968,N_2100);
nor U3052 (N_3052,N_2088,N_2124);
or U3053 (N_3053,N_1763,N_1742);
and U3054 (N_3054,N_1868,N_1396);
xnor U3055 (N_3055,N_1534,N_1719);
or U3056 (N_3056,N_1440,N_2356);
nand U3057 (N_3057,N_1564,N_1495);
nand U3058 (N_3058,N_1332,N_1352);
nand U3059 (N_3059,N_1751,N_1982);
and U3060 (N_3060,N_1487,N_1879);
xor U3061 (N_3061,N_2277,N_1420);
nand U3062 (N_3062,N_1931,N_1894);
and U3063 (N_3063,N_1917,N_2222);
xor U3064 (N_3064,N_1693,N_1306);
and U3065 (N_3065,N_2300,N_2297);
or U3066 (N_3066,N_2167,N_1541);
and U3067 (N_3067,N_1814,N_1335);
xor U3068 (N_3068,N_1578,N_1774);
and U3069 (N_3069,N_1852,N_2257);
nor U3070 (N_3070,N_1799,N_1402);
nand U3071 (N_3071,N_2335,N_2201);
and U3072 (N_3072,N_2073,N_1394);
nand U3073 (N_3073,N_2489,N_2474);
nor U3074 (N_3074,N_1749,N_1976);
nor U3075 (N_3075,N_1840,N_1631);
and U3076 (N_3076,N_1583,N_2344);
and U3077 (N_3077,N_1913,N_1430);
nor U3078 (N_3078,N_1422,N_2098);
and U3079 (N_3079,N_2226,N_2289);
nor U3080 (N_3080,N_1328,N_2091);
nand U3081 (N_3081,N_1419,N_2365);
xnor U3082 (N_3082,N_1949,N_1764);
xnor U3083 (N_3083,N_2028,N_2498);
or U3084 (N_3084,N_1452,N_1848);
and U3085 (N_3085,N_1334,N_2409);
and U3086 (N_3086,N_1449,N_2271);
nand U3087 (N_3087,N_2224,N_1654);
nor U3088 (N_3088,N_1388,N_1609);
and U3089 (N_3089,N_2095,N_2481);
nor U3090 (N_3090,N_2385,N_1705);
xnor U3091 (N_3091,N_1558,N_2235);
xor U3092 (N_3092,N_1498,N_2487);
nor U3093 (N_3093,N_1346,N_2463);
and U3094 (N_3094,N_1892,N_2307);
nor U3095 (N_3095,N_1299,N_1484);
nor U3096 (N_3096,N_1790,N_1943);
nand U3097 (N_3097,N_2151,N_2479);
nand U3098 (N_3098,N_1876,N_2460);
or U3099 (N_3099,N_1888,N_1812);
nand U3100 (N_3100,N_1950,N_2159);
xor U3101 (N_3101,N_1775,N_1841);
or U3102 (N_3102,N_2364,N_1956);
nand U3103 (N_3103,N_2426,N_1502);
and U3104 (N_3104,N_1619,N_1718);
xor U3105 (N_3105,N_2281,N_1655);
and U3106 (N_3106,N_2040,N_1853);
xnor U3107 (N_3107,N_1492,N_1664);
xor U3108 (N_3108,N_2187,N_1784);
nand U3109 (N_3109,N_1290,N_1708);
nor U3110 (N_3110,N_1651,N_2108);
nand U3111 (N_3111,N_1854,N_1268);
or U3112 (N_3112,N_1368,N_1436);
xnor U3113 (N_3113,N_1856,N_2472);
and U3114 (N_3114,N_1594,N_1987);
nand U3115 (N_3115,N_1433,N_2031);
and U3116 (N_3116,N_1798,N_1477);
nand U3117 (N_3117,N_2128,N_1336);
nand U3118 (N_3118,N_1591,N_1990);
and U3119 (N_3119,N_2315,N_1944);
nand U3120 (N_3120,N_2177,N_1442);
nand U3121 (N_3121,N_1777,N_1625);
or U3122 (N_3122,N_1491,N_2079);
and U3123 (N_3123,N_2459,N_2018);
nand U3124 (N_3124,N_2468,N_1998);
and U3125 (N_3125,N_2243,N_2150);
or U3126 (N_3126,N_1760,N_1411);
or U3127 (N_3127,N_2172,N_2180);
xor U3128 (N_3128,N_1845,N_2308);
nor U3129 (N_3129,N_1632,N_1538);
nor U3130 (N_3130,N_1631,N_1615);
nand U3131 (N_3131,N_1593,N_1483);
nand U3132 (N_3132,N_2343,N_1415);
or U3133 (N_3133,N_1479,N_1944);
or U3134 (N_3134,N_1863,N_1330);
xnor U3135 (N_3135,N_1259,N_1421);
or U3136 (N_3136,N_1274,N_2438);
or U3137 (N_3137,N_1978,N_1782);
or U3138 (N_3138,N_1315,N_1485);
nand U3139 (N_3139,N_2344,N_1457);
and U3140 (N_3140,N_2334,N_1743);
xor U3141 (N_3141,N_1589,N_1706);
nand U3142 (N_3142,N_1261,N_1804);
or U3143 (N_3143,N_2052,N_2068);
and U3144 (N_3144,N_1535,N_1478);
or U3145 (N_3145,N_2325,N_1418);
nor U3146 (N_3146,N_1899,N_1582);
or U3147 (N_3147,N_2457,N_1867);
and U3148 (N_3148,N_2034,N_1485);
xor U3149 (N_3149,N_2259,N_1926);
and U3150 (N_3150,N_2482,N_2447);
xor U3151 (N_3151,N_1644,N_1622);
xnor U3152 (N_3152,N_1430,N_2280);
xor U3153 (N_3153,N_1910,N_1831);
and U3154 (N_3154,N_1892,N_1872);
nor U3155 (N_3155,N_2384,N_2292);
nand U3156 (N_3156,N_1270,N_2441);
and U3157 (N_3157,N_1891,N_2251);
nor U3158 (N_3158,N_2026,N_1622);
and U3159 (N_3159,N_1906,N_1568);
xnor U3160 (N_3160,N_2494,N_2186);
nor U3161 (N_3161,N_1945,N_1841);
nor U3162 (N_3162,N_2379,N_1346);
xor U3163 (N_3163,N_1953,N_1740);
nor U3164 (N_3164,N_1476,N_1291);
xnor U3165 (N_3165,N_2441,N_1567);
nor U3166 (N_3166,N_1802,N_1291);
nor U3167 (N_3167,N_1420,N_2435);
and U3168 (N_3168,N_2465,N_2159);
xnor U3169 (N_3169,N_1898,N_1491);
and U3170 (N_3170,N_1481,N_1702);
xnor U3171 (N_3171,N_1447,N_2491);
nor U3172 (N_3172,N_1631,N_1454);
nor U3173 (N_3173,N_1431,N_1690);
nor U3174 (N_3174,N_1384,N_1903);
xor U3175 (N_3175,N_1857,N_1684);
xnor U3176 (N_3176,N_1609,N_1432);
xor U3177 (N_3177,N_1659,N_1852);
and U3178 (N_3178,N_2170,N_2470);
and U3179 (N_3179,N_2405,N_1995);
or U3180 (N_3180,N_1608,N_1673);
nand U3181 (N_3181,N_2030,N_1288);
or U3182 (N_3182,N_2014,N_2300);
or U3183 (N_3183,N_2164,N_1537);
xor U3184 (N_3184,N_1570,N_1705);
or U3185 (N_3185,N_2273,N_2195);
nor U3186 (N_3186,N_1770,N_1748);
nand U3187 (N_3187,N_1926,N_2396);
or U3188 (N_3188,N_2484,N_1605);
xnor U3189 (N_3189,N_2468,N_2170);
and U3190 (N_3190,N_1932,N_1879);
and U3191 (N_3191,N_2401,N_1956);
xnor U3192 (N_3192,N_1755,N_2074);
or U3193 (N_3193,N_1956,N_1473);
nand U3194 (N_3194,N_1682,N_2037);
and U3195 (N_3195,N_1281,N_2073);
or U3196 (N_3196,N_2325,N_1514);
nor U3197 (N_3197,N_1654,N_1413);
xor U3198 (N_3198,N_1342,N_1814);
nand U3199 (N_3199,N_2341,N_2336);
nand U3200 (N_3200,N_2292,N_1685);
xor U3201 (N_3201,N_2483,N_1934);
or U3202 (N_3202,N_1341,N_1563);
nand U3203 (N_3203,N_1494,N_2330);
or U3204 (N_3204,N_2170,N_1906);
nor U3205 (N_3205,N_1761,N_2370);
xnor U3206 (N_3206,N_2108,N_1774);
and U3207 (N_3207,N_2260,N_1299);
or U3208 (N_3208,N_2028,N_1414);
or U3209 (N_3209,N_1809,N_1440);
and U3210 (N_3210,N_2435,N_2252);
and U3211 (N_3211,N_1381,N_2386);
xnor U3212 (N_3212,N_1326,N_1913);
nor U3213 (N_3213,N_2050,N_1548);
or U3214 (N_3214,N_1437,N_2079);
and U3215 (N_3215,N_2461,N_1862);
or U3216 (N_3216,N_2269,N_2311);
xor U3217 (N_3217,N_2341,N_2150);
nand U3218 (N_3218,N_2003,N_1541);
or U3219 (N_3219,N_1879,N_2432);
or U3220 (N_3220,N_1991,N_1371);
and U3221 (N_3221,N_2161,N_1880);
xnor U3222 (N_3222,N_2313,N_2044);
nand U3223 (N_3223,N_1922,N_1957);
nor U3224 (N_3224,N_2326,N_1922);
nor U3225 (N_3225,N_1480,N_2180);
nor U3226 (N_3226,N_1421,N_1343);
and U3227 (N_3227,N_1866,N_1622);
nor U3228 (N_3228,N_2286,N_1520);
or U3229 (N_3229,N_1331,N_1678);
or U3230 (N_3230,N_2470,N_1507);
and U3231 (N_3231,N_1760,N_2187);
and U3232 (N_3232,N_1538,N_1324);
and U3233 (N_3233,N_2475,N_1304);
nor U3234 (N_3234,N_1338,N_1862);
xor U3235 (N_3235,N_1717,N_2155);
nor U3236 (N_3236,N_1963,N_1823);
xor U3237 (N_3237,N_2053,N_2005);
xnor U3238 (N_3238,N_2386,N_2201);
or U3239 (N_3239,N_2091,N_1980);
and U3240 (N_3240,N_1649,N_1939);
and U3241 (N_3241,N_2459,N_1497);
xnor U3242 (N_3242,N_1474,N_1486);
and U3243 (N_3243,N_1690,N_2329);
xor U3244 (N_3244,N_1311,N_1755);
and U3245 (N_3245,N_1553,N_2065);
nand U3246 (N_3246,N_2266,N_2388);
xor U3247 (N_3247,N_1779,N_2365);
xor U3248 (N_3248,N_1543,N_1830);
and U3249 (N_3249,N_2127,N_2142);
xnor U3250 (N_3250,N_2014,N_2363);
and U3251 (N_3251,N_1451,N_2112);
nand U3252 (N_3252,N_1806,N_1771);
nor U3253 (N_3253,N_2398,N_1604);
or U3254 (N_3254,N_2350,N_2237);
nand U3255 (N_3255,N_2457,N_1300);
xnor U3256 (N_3256,N_2133,N_2170);
nand U3257 (N_3257,N_1380,N_2232);
or U3258 (N_3258,N_1712,N_2431);
or U3259 (N_3259,N_1528,N_2402);
or U3260 (N_3260,N_1451,N_2065);
xnor U3261 (N_3261,N_1897,N_1860);
and U3262 (N_3262,N_1527,N_1967);
and U3263 (N_3263,N_1995,N_2388);
xor U3264 (N_3264,N_2204,N_1824);
or U3265 (N_3265,N_2085,N_2296);
or U3266 (N_3266,N_1519,N_1309);
nor U3267 (N_3267,N_1444,N_1520);
xor U3268 (N_3268,N_2020,N_1713);
or U3269 (N_3269,N_2216,N_1644);
nor U3270 (N_3270,N_1604,N_1953);
or U3271 (N_3271,N_2241,N_1435);
nand U3272 (N_3272,N_1568,N_2249);
xnor U3273 (N_3273,N_1680,N_2401);
nor U3274 (N_3274,N_1462,N_2246);
or U3275 (N_3275,N_1400,N_1503);
nor U3276 (N_3276,N_2108,N_1414);
xor U3277 (N_3277,N_2277,N_2042);
nand U3278 (N_3278,N_2131,N_2343);
nor U3279 (N_3279,N_2012,N_2395);
nor U3280 (N_3280,N_2188,N_2027);
nor U3281 (N_3281,N_1350,N_2497);
nand U3282 (N_3282,N_1852,N_2220);
and U3283 (N_3283,N_2360,N_2391);
xnor U3284 (N_3284,N_2176,N_1341);
nand U3285 (N_3285,N_1762,N_2362);
or U3286 (N_3286,N_2207,N_1975);
or U3287 (N_3287,N_1989,N_1507);
and U3288 (N_3288,N_2215,N_2210);
xnor U3289 (N_3289,N_1723,N_1425);
and U3290 (N_3290,N_2051,N_1276);
nor U3291 (N_3291,N_1656,N_2194);
and U3292 (N_3292,N_1974,N_1762);
nand U3293 (N_3293,N_1770,N_1805);
xor U3294 (N_3294,N_1538,N_1860);
nor U3295 (N_3295,N_2087,N_2416);
xor U3296 (N_3296,N_1343,N_1308);
xor U3297 (N_3297,N_2223,N_2414);
nand U3298 (N_3298,N_1610,N_2414);
nor U3299 (N_3299,N_2452,N_1912);
nand U3300 (N_3300,N_1418,N_1876);
xor U3301 (N_3301,N_1664,N_1950);
or U3302 (N_3302,N_1966,N_2290);
nand U3303 (N_3303,N_1605,N_1444);
or U3304 (N_3304,N_1366,N_1843);
nor U3305 (N_3305,N_2399,N_2471);
or U3306 (N_3306,N_1951,N_1611);
and U3307 (N_3307,N_1991,N_2142);
xor U3308 (N_3308,N_1256,N_2222);
nand U3309 (N_3309,N_2120,N_1649);
xor U3310 (N_3310,N_2086,N_1719);
xnor U3311 (N_3311,N_1749,N_1293);
and U3312 (N_3312,N_1437,N_1478);
nand U3313 (N_3313,N_1677,N_2320);
nor U3314 (N_3314,N_1793,N_2078);
and U3315 (N_3315,N_2373,N_2308);
or U3316 (N_3316,N_1332,N_1575);
nand U3317 (N_3317,N_2498,N_1330);
nand U3318 (N_3318,N_1634,N_1482);
and U3319 (N_3319,N_2361,N_2468);
xnor U3320 (N_3320,N_1345,N_1263);
nor U3321 (N_3321,N_2252,N_2201);
nand U3322 (N_3322,N_1501,N_2188);
xor U3323 (N_3323,N_1950,N_1256);
nand U3324 (N_3324,N_1595,N_2252);
or U3325 (N_3325,N_1701,N_1358);
and U3326 (N_3326,N_1542,N_1280);
xor U3327 (N_3327,N_1588,N_1916);
or U3328 (N_3328,N_1384,N_2339);
nand U3329 (N_3329,N_1463,N_1623);
or U3330 (N_3330,N_1350,N_1437);
nand U3331 (N_3331,N_1642,N_2272);
nor U3332 (N_3332,N_2296,N_1677);
and U3333 (N_3333,N_2499,N_2225);
nor U3334 (N_3334,N_1463,N_1738);
and U3335 (N_3335,N_1365,N_1448);
nand U3336 (N_3336,N_1422,N_1729);
or U3337 (N_3337,N_2052,N_1433);
xor U3338 (N_3338,N_1825,N_2014);
xor U3339 (N_3339,N_2150,N_2065);
nor U3340 (N_3340,N_1962,N_2118);
nor U3341 (N_3341,N_1274,N_2123);
and U3342 (N_3342,N_2060,N_1518);
nand U3343 (N_3343,N_2358,N_2157);
nor U3344 (N_3344,N_2016,N_2421);
or U3345 (N_3345,N_1592,N_2381);
or U3346 (N_3346,N_1727,N_2474);
and U3347 (N_3347,N_2189,N_2167);
or U3348 (N_3348,N_1477,N_1810);
nor U3349 (N_3349,N_1901,N_1762);
or U3350 (N_3350,N_2260,N_2377);
and U3351 (N_3351,N_1761,N_1308);
nor U3352 (N_3352,N_1790,N_1807);
or U3353 (N_3353,N_1992,N_1524);
xnor U3354 (N_3354,N_1341,N_2147);
xnor U3355 (N_3355,N_2083,N_1990);
xor U3356 (N_3356,N_2263,N_1937);
nor U3357 (N_3357,N_2415,N_2192);
nor U3358 (N_3358,N_1564,N_1280);
nand U3359 (N_3359,N_2379,N_2218);
nor U3360 (N_3360,N_1449,N_1733);
xor U3361 (N_3361,N_1967,N_1266);
nand U3362 (N_3362,N_1654,N_2062);
xor U3363 (N_3363,N_2332,N_2164);
and U3364 (N_3364,N_2252,N_2421);
or U3365 (N_3365,N_2311,N_1969);
or U3366 (N_3366,N_1292,N_1842);
or U3367 (N_3367,N_2040,N_1258);
nand U3368 (N_3368,N_1684,N_2199);
or U3369 (N_3369,N_2271,N_2402);
nand U3370 (N_3370,N_1375,N_1428);
xnor U3371 (N_3371,N_2203,N_1827);
and U3372 (N_3372,N_2178,N_2078);
and U3373 (N_3373,N_1746,N_2036);
xnor U3374 (N_3374,N_2401,N_2286);
xor U3375 (N_3375,N_1928,N_1372);
nand U3376 (N_3376,N_2285,N_2331);
xnor U3377 (N_3377,N_1562,N_1635);
or U3378 (N_3378,N_1356,N_2171);
and U3379 (N_3379,N_1829,N_2248);
nor U3380 (N_3380,N_2141,N_1840);
xnor U3381 (N_3381,N_2154,N_2203);
nand U3382 (N_3382,N_1756,N_1893);
nand U3383 (N_3383,N_1424,N_2350);
and U3384 (N_3384,N_2019,N_1262);
or U3385 (N_3385,N_1315,N_1512);
nor U3386 (N_3386,N_2471,N_2081);
xnor U3387 (N_3387,N_1700,N_2171);
nand U3388 (N_3388,N_1839,N_1640);
xnor U3389 (N_3389,N_2159,N_1809);
nor U3390 (N_3390,N_2476,N_1293);
or U3391 (N_3391,N_1710,N_1438);
or U3392 (N_3392,N_2424,N_1426);
xnor U3393 (N_3393,N_2081,N_1729);
or U3394 (N_3394,N_2205,N_2232);
or U3395 (N_3395,N_2426,N_2253);
nand U3396 (N_3396,N_1409,N_2227);
or U3397 (N_3397,N_2414,N_2370);
nor U3398 (N_3398,N_2265,N_1481);
nor U3399 (N_3399,N_1444,N_1828);
and U3400 (N_3400,N_1306,N_1720);
or U3401 (N_3401,N_2222,N_1556);
xnor U3402 (N_3402,N_1302,N_1598);
and U3403 (N_3403,N_1446,N_2021);
nand U3404 (N_3404,N_1380,N_1396);
nor U3405 (N_3405,N_2035,N_2209);
nor U3406 (N_3406,N_2411,N_1906);
and U3407 (N_3407,N_2080,N_1874);
nand U3408 (N_3408,N_2238,N_1724);
or U3409 (N_3409,N_1503,N_2395);
nand U3410 (N_3410,N_2434,N_1486);
nor U3411 (N_3411,N_1752,N_1345);
or U3412 (N_3412,N_1509,N_1384);
nand U3413 (N_3413,N_1639,N_2304);
nand U3414 (N_3414,N_1867,N_2241);
and U3415 (N_3415,N_1269,N_1401);
or U3416 (N_3416,N_2233,N_2259);
and U3417 (N_3417,N_1798,N_2147);
or U3418 (N_3418,N_2096,N_2309);
or U3419 (N_3419,N_2166,N_2263);
or U3420 (N_3420,N_2347,N_2314);
and U3421 (N_3421,N_2438,N_1362);
and U3422 (N_3422,N_2303,N_2277);
xor U3423 (N_3423,N_2408,N_1461);
and U3424 (N_3424,N_1437,N_2196);
nor U3425 (N_3425,N_2355,N_1336);
nand U3426 (N_3426,N_2327,N_1431);
or U3427 (N_3427,N_2327,N_2198);
nand U3428 (N_3428,N_1919,N_2488);
nor U3429 (N_3429,N_2193,N_1683);
nor U3430 (N_3430,N_1860,N_2224);
or U3431 (N_3431,N_2250,N_2369);
nor U3432 (N_3432,N_2009,N_2055);
nand U3433 (N_3433,N_1687,N_2344);
or U3434 (N_3434,N_1300,N_1926);
and U3435 (N_3435,N_2150,N_2491);
or U3436 (N_3436,N_1273,N_2049);
nand U3437 (N_3437,N_2300,N_1496);
or U3438 (N_3438,N_2039,N_2189);
nor U3439 (N_3439,N_1927,N_1442);
nand U3440 (N_3440,N_1749,N_1861);
or U3441 (N_3441,N_2303,N_2447);
and U3442 (N_3442,N_1530,N_1394);
nor U3443 (N_3443,N_1826,N_1276);
xnor U3444 (N_3444,N_2058,N_1532);
or U3445 (N_3445,N_2204,N_1725);
nand U3446 (N_3446,N_1835,N_1877);
xnor U3447 (N_3447,N_2235,N_2271);
xor U3448 (N_3448,N_1416,N_1369);
xnor U3449 (N_3449,N_2098,N_1884);
or U3450 (N_3450,N_1386,N_2444);
and U3451 (N_3451,N_1533,N_1348);
or U3452 (N_3452,N_1546,N_2229);
or U3453 (N_3453,N_1896,N_1605);
nand U3454 (N_3454,N_1660,N_2261);
nand U3455 (N_3455,N_1280,N_1460);
or U3456 (N_3456,N_2054,N_2357);
nand U3457 (N_3457,N_2009,N_1796);
and U3458 (N_3458,N_1791,N_2374);
or U3459 (N_3459,N_1914,N_1544);
nand U3460 (N_3460,N_1843,N_1553);
nand U3461 (N_3461,N_2459,N_1839);
xor U3462 (N_3462,N_1425,N_1729);
and U3463 (N_3463,N_1459,N_1377);
nand U3464 (N_3464,N_2259,N_2058);
or U3465 (N_3465,N_1908,N_1690);
nand U3466 (N_3466,N_2311,N_2376);
and U3467 (N_3467,N_1935,N_2258);
and U3468 (N_3468,N_2086,N_1896);
or U3469 (N_3469,N_1556,N_2119);
nand U3470 (N_3470,N_1668,N_1577);
and U3471 (N_3471,N_2295,N_2369);
nand U3472 (N_3472,N_1568,N_1708);
or U3473 (N_3473,N_1350,N_1811);
and U3474 (N_3474,N_1771,N_1795);
xnor U3475 (N_3475,N_1977,N_1684);
nand U3476 (N_3476,N_1999,N_1899);
xnor U3477 (N_3477,N_2422,N_1592);
or U3478 (N_3478,N_2158,N_1692);
nor U3479 (N_3479,N_2490,N_1421);
nor U3480 (N_3480,N_2107,N_1374);
nor U3481 (N_3481,N_2473,N_2379);
nor U3482 (N_3482,N_1553,N_2082);
nand U3483 (N_3483,N_2464,N_1284);
or U3484 (N_3484,N_2497,N_1396);
nor U3485 (N_3485,N_1419,N_1646);
nand U3486 (N_3486,N_2114,N_1841);
and U3487 (N_3487,N_2186,N_1919);
and U3488 (N_3488,N_2249,N_1526);
nand U3489 (N_3489,N_1317,N_1525);
nand U3490 (N_3490,N_1395,N_1293);
nor U3491 (N_3491,N_1905,N_1952);
and U3492 (N_3492,N_1846,N_1739);
or U3493 (N_3493,N_2063,N_1875);
or U3494 (N_3494,N_1725,N_1905);
xnor U3495 (N_3495,N_2046,N_1797);
or U3496 (N_3496,N_1469,N_1870);
nand U3497 (N_3497,N_1557,N_1778);
nand U3498 (N_3498,N_1336,N_1900);
xnor U3499 (N_3499,N_2269,N_1529);
nand U3500 (N_3500,N_2228,N_1654);
nand U3501 (N_3501,N_2020,N_1360);
or U3502 (N_3502,N_1585,N_2388);
or U3503 (N_3503,N_2143,N_1255);
nor U3504 (N_3504,N_1535,N_1752);
nor U3505 (N_3505,N_1874,N_2482);
xor U3506 (N_3506,N_1550,N_1899);
or U3507 (N_3507,N_1809,N_2337);
xnor U3508 (N_3508,N_1778,N_2169);
and U3509 (N_3509,N_1572,N_2111);
or U3510 (N_3510,N_1941,N_2353);
nand U3511 (N_3511,N_2460,N_2279);
or U3512 (N_3512,N_2199,N_1766);
and U3513 (N_3513,N_1937,N_2340);
and U3514 (N_3514,N_1675,N_1433);
nor U3515 (N_3515,N_1774,N_2093);
nand U3516 (N_3516,N_1433,N_2372);
and U3517 (N_3517,N_1571,N_1778);
or U3518 (N_3518,N_1701,N_1250);
xnor U3519 (N_3519,N_1483,N_1904);
and U3520 (N_3520,N_1950,N_1593);
nor U3521 (N_3521,N_1680,N_2320);
or U3522 (N_3522,N_2298,N_2196);
xor U3523 (N_3523,N_1511,N_2332);
and U3524 (N_3524,N_1956,N_2155);
nor U3525 (N_3525,N_1443,N_1311);
and U3526 (N_3526,N_1453,N_1535);
and U3527 (N_3527,N_1690,N_2472);
xnor U3528 (N_3528,N_1724,N_2295);
and U3529 (N_3529,N_2439,N_1574);
xor U3530 (N_3530,N_1723,N_2287);
xnor U3531 (N_3531,N_2351,N_2051);
nand U3532 (N_3532,N_1509,N_2384);
xor U3533 (N_3533,N_1975,N_2377);
nand U3534 (N_3534,N_2472,N_1492);
and U3535 (N_3535,N_1928,N_2222);
and U3536 (N_3536,N_1593,N_1671);
or U3537 (N_3537,N_1539,N_2433);
and U3538 (N_3538,N_2358,N_2162);
and U3539 (N_3539,N_2066,N_1701);
and U3540 (N_3540,N_1472,N_1938);
nand U3541 (N_3541,N_1281,N_1802);
and U3542 (N_3542,N_1605,N_1478);
nor U3543 (N_3543,N_2302,N_1765);
xnor U3544 (N_3544,N_2018,N_2154);
and U3545 (N_3545,N_1350,N_1478);
and U3546 (N_3546,N_2022,N_2089);
nor U3547 (N_3547,N_1455,N_1964);
and U3548 (N_3548,N_1326,N_2226);
and U3549 (N_3549,N_2378,N_2360);
nand U3550 (N_3550,N_1416,N_2252);
and U3551 (N_3551,N_1735,N_2226);
or U3552 (N_3552,N_2035,N_1690);
nor U3553 (N_3553,N_2310,N_1804);
xnor U3554 (N_3554,N_1907,N_2480);
xor U3555 (N_3555,N_1472,N_1914);
nor U3556 (N_3556,N_1285,N_1588);
xor U3557 (N_3557,N_1871,N_1472);
xor U3558 (N_3558,N_1650,N_1352);
or U3559 (N_3559,N_1517,N_1635);
or U3560 (N_3560,N_1279,N_2363);
xnor U3561 (N_3561,N_1717,N_1966);
xnor U3562 (N_3562,N_1294,N_2142);
or U3563 (N_3563,N_2304,N_2317);
nand U3564 (N_3564,N_2347,N_1969);
and U3565 (N_3565,N_2387,N_2021);
nor U3566 (N_3566,N_2160,N_1342);
and U3567 (N_3567,N_1912,N_1669);
nor U3568 (N_3568,N_2087,N_1709);
nor U3569 (N_3569,N_1259,N_2131);
xor U3570 (N_3570,N_1335,N_2467);
and U3571 (N_3571,N_2045,N_1564);
and U3572 (N_3572,N_1719,N_2494);
xor U3573 (N_3573,N_1572,N_2391);
or U3574 (N_3574,N_2449,N_2097);
and U3575 (N_3575,N_1290,N_1598);
nor U3576 (N_3576,N_1971,N_1598);
nand U3577 (N_3577,N_1927,N_2363);
nand U3578 (N_3578,N_1884,N_2427);
nand U3579 (N_3579,N_1835,N_1706);
xor U3580 (N_3580,N_2318,N_2498);
nor U3581 (N_3581,N_2328,N_1767);
and U3582 (N_3582,N_2179,N_1510);
nor U3583 (N_3583,N_1661,N_1908);
and U3584 (N_3584,N_2275,N_2067);
nand U3585 (N_3585,N_2399,N_2131);
nand U3586 (N_3586,N_1665,N_2145);
nor U3587 (N_3587,N_1861,N_1545);
nor U3588 (N_3588,N_1640,N_1814);
nand U3589 (N_3589,N_2246,N_2189);
nand U3590 (N_3590,N_1896,N_2130);
and U3591 (N_3591,N_1490,N_1618);
nand U3592 (N_3592,N_1912,N_1397);
nor U3593 (N_3593,N_1526,N_1788);
nand U3594 (N_3594,N_1775,N_1634);
or U3595 (N_3595,N_2182,N_1286);
xor U3596 (N_3596,N_2362,N_1443);
and U3597 (N_3597,N_2135,N_1680);
and U3598 (N_3598,N_2048,N_1725);
and U3599 (N_3599,N_1809,N_1267);
and U3600 (N_3600,N_1776,N_2353);
nand U3601 (N_3601,N_2138,N_2242);
and U3602 (N_3602,N_1495,N_2019);
and U3603 (N_3603,N_2249,N_2312);
nand U3604 (N_3604,N_1944,N_1693);
xor U3605 (N_3605,N_2088,N_1762);
and U3606 (N_3606,N_2373,N_2309);
nand U3607 (N_3607,N_2148,N_1688);
and U3608 (N_3608,N_1322,N_2035);
nand U3609 (N_3609,N_1692,N_1354);
nand U3610 (N_3610,N_1309,N_1984);
and U3611 (N_3611,N_1897,N_1569);
nand U3612 (N_3612,N_2291,N_1900);
or U3613 (N_3613,N_2268,N_1759);
nand U3614 (N_3614,N_2410,N_1350);
or U3615 (N_3615,N_1896,N_1902);
nand U3616 (N_3616,N_1529,N_2425);
nand U3617 (N_3617,N_2010,N_2113);
and U3618 (N_3618,N_1631,N_2086);
or U3619 (N_3619,N_1535,N_2314);
nand U3620 (N_3620,N_1835,N_1952);
and U3621 (N_3621,N_1697,N_2487);
and U3622 (N_3622,N_1816,N_1984);
or U3623 (N_3623,N_1314,N_2254);
and U3624 (N_3624,N_2232,N_1776);
xnor U3625 (N_3625,N_1650,N_2398);
xor U3626 (N_3626,N_1934,N_1920);
nor U3627 (N_3627,N_1411,N_1426);
or U3628 (N_3628,N_1584,N_2021);
and U3629 (N_3629,N_2446,N_1787);
nor U3630 (N_3630,N_2314,N_2209);
nand U3631 (N_3631,N_2482,N_1738);
and U3632 (N_3632,N_1427,N_1470);
or U3633 (N_3633,N_2137,N_2195);
and U3634 (N_3634,N_1335,N_1473);
nand U3635 (N_3635,N_2119,N_2443);
or U3636 (N_3636,N_1929,N_1645);
nor U3637 (N_3637,N_2336,N_2497);
nor U3638 (N_3638,N_2129,N_2440);
nand U3639 (N_3639,N_1469,N_1585);
and U3640 (N_3640,N_2368,N_1908);
xor U3641 (N_3641,N_1599,N_2191);
xor U3642 (N_3642,N_1740,N_2403);
nand U3643 (N_3643,N_1904,N_1877);
nor U3644 (N_3644,N_1857,N_2024);
and U3645 (N_3645,N_1673,N_1851);
nand U3646 (N_3646,N_2104,N_2291);
and U3647 (N_3647,N_1643,N_2110);
or U3648 (N_3648,N_1927,N_1491);
and U3649 (N_3649,N_1675,N_2075);
nand U3650 (N_3650,N_1683,N_1953);
and U3651 (N_3651,N_1600,N_1440);
and U3652 (N_3652,N_1899,N_1690);
xnor U3653 (N_3653,N_1512,N_2089);
or U3654 (N_3654,N_2247,N_1985);
nor U3655 (N_3655,N_1912,N_2300);
xor U3656 (N_3656,N_1343,N_1960);
and U3657 (N_3657,N_1648,N_1653);
and U3658 (N_3658,N_1722,N_2049);
and U3659 (N_3659,N_2232,N_1400);
nor U3660 (N_3660,N_2026,N_1590);
or U3661 (N_3661,N_1900,N_2044);
and U3662 (N_3662,N_1937,N_2123);
and U3663 (N_3663,N_1473,N_1844);
and U3664 (N_3664,N_2038,N_2474);
xor U3665 (N_3665,N_1298,N_2384);
or U3666 (N_3666,N_2044,N_2478);
nand U3667 (N_3667,N_2254,N_1666);
xor U3668 (N_3668,N_1704,N_2125);
xor U3669 (N_3669,N_2118,N_1825);
nor U3670 (N_3670,N_1697,N_2387);
nand U3671 (N_3671,N_2185,N_1402);
nor U3672 (N_3672,N_1670,N_2328);
nand U3673 (N_3673,N_1631,N_1475);
nand U3674 (N_3674,N_1490,N_2283);
nand U3675 (N_3675,N_1731,N_2020);
nand U3676 (N_3676,N_2492,N_1688);
nor U3677 (N_3677,N_1463,N_1934);
nor U3678 (N_3678,N_1981,N_1855);
nand U3679 (N_3679,N_1428,N_2115);
and U3680 (N_3680,N_1261,N_2263);
nor U3681 (N_3681,N_2155,N_1467);
and U3682 (N_3682,N_1867,N_1454);
nor U3683 (N_3683,N_2237,N_1319);
or U3684 (N_3684,N_1813,N_2104);
nand U3685 (N_3685,N_1438,N_1951);
nand U3686 (N_3686,N_1827,N_1454);
or U3687 (N_3687,N_1783,N_1287);
or U3688 (N_3688,N_2099,N_1291);
xor U3689 (N_3689,N_2334,N_2192);
nor U3690 (N_3690,N_2401,N_1272);
nand U3691 (N_3691,N_2168,N_1863);
nor U3692 (N_3692,N_1515,N_2288);
and U3693 (N_3693,N_1767,N_1356);
xnor U3694 (N_3694,N_1333,N_1558);
or U3695 (N_3695,N_1573,N_1896);
or U3696 (N_3696,N_1412,N_2465);
and U3697 (N_3697,N_1706,N_1849);
xnor U3698 (N_3698,N_1361,N_1443);
xor U3699 (N_3699,N_1780,N_1450);
nor U3700 (N_3700,N_2054,N_1503);
or U3701 (N_3701,N_1357,N_2172);
nand U3702 (N_3702,N_1876,N_2291);
and U3703 (N_3703,N_2369,N_1955);
or U3704 (N_3704,N_2484,N_2389);
nor U3705 (N_3705,N_2335,N_2312);
and U3706 (N_3706,N_2034,N_1529);
nor U3707 (N_3707,N_1700,N_1278);
xor U3708 (N_3708,N_1455,N_1790);
nand U3709 (N_3709,N_1600,N_1976);
or U3710 (N_3710,N_1634,N_1919);
nand U3711 (N_3711,N_1855,N_2204);
nor U3712 (N_3712,N_1591,N_2012);
nor U3713 (N_3713,N_1474,N_1844);
nor U3714 (N_3714,N_1478,N_2275);
xnor U3715 (N_3715,N_1471,N_1525);
nor U3716 (N_3716,N_2092,N_1325);
or U3717 (N_3717,N_1984,N_1646);
xor U3718 (N_3718,N_2036,N_1578);
or U3719 (N_3719,N_1268,N_1858);
and U3720 (N_3720,N_1528,N_1511);
xnor U3721 (N_3721,N_1528,N_2210);
nand U3722 (N_3722,N_1311,N_1858);
xor U3723 (N_3723,N_2289,N_1634);
xnor U3724 (N_3724,N_2451,N_1335);
and U3725 (N_3725,N_1952,N_1440);
or U3726 (N_3726,N_1448,N_1295);
nor U3727 (N_3727,N_1647,N_2231);
xnor U3728 (N_3728,N_1960,N_2482);
nand U3729 (N_3729,N_1875,N_2455);
nand U3730 (N_3730,N_1662,N_2378);
nor U3731 (N_3731,N_1765,N_1342);
nor U3732 (N_3732,N_2304,N_1994);
nor U3733 (N_3733,N_1885,N_1662);
nor U3734 (N_3734,N_2238,N_1417);
or U3735 (N_3735,N_1895,N_1821);
and U3736 (N_3736,N_1687,N_2251);
or U3737 (N_3737,N_1824,N_1311);
nor U3738 (N_3738,N_2004,N_2316);
nor U3739 (N_3739,N_2207,N_1431);
xor U3740 (N_3740,N_1963,N_1488);
or U3741 (N_3741,N_2011,N_1555);
xor U3742 (N_3742,N_1951,N_2378);
nand U3743 (N_3743,N_1259,N_1429);
and U3744 (N_3744,N_1463,N_2420);
nand U3745 (N_3745,N_1517,N_1876);
nor U3746 (N_3746,N_1441,N_1486);
nand U3747 (N_3747,N_1582,N_1324);
and U3748 (N_3748,N_2023,N_1337);
nand U3749 (N_3749,N_2071,N_1470);
and U3750 (N_3750,N_2834,N_3347);
nand U3751 (N_3751,N_2617,N_3467);
or U3752 (N_3752,N_3358,N_3541);
xnor U3753 (N_3753,N_3498,N_3184);
xnor U3754 (N_3754,N_2668,N_2640);
nor U3755 (N_3755,N_3535,N_2928);
or U3756 (N_3756,N_2889,N_3082);
or U3757 (N_3757,N_3202,N_2576);
nand U3758 (N_3758,N_2633,N_2541);
and U3759 (N_3759,N_3552,N_3011);
xnor U3760 (N_3760,N_2872,N_2596);
or U3761 (N_3761,N_2887,N_2568);
and U3762 (N_3762,N_2980,N_2999);
nor U3763 (N_3763,N_3105,N_3651);
and U3764 (N_3764,N_2781,N_3282);
nor U3765 (N_3765,N_2672,N_3592);
and U3766 (N_3766,N_3086,N_3598);
nor U3767 (N_3767,N_3696,N_2918);
xnor U3768 (N_3768,N_3345,N_2560);
and U3769 (N_3769,N_2935,N_2610);
xor U3770 (N_3770,N_3269,N_2657);
nor U3771 (N_3771,N_2730,N_3477);
nor U3772 (N_3772,N_3146,N_3420);
nand U3773 (N_3773,N_2690,N_2595);
xor U3774 (N_3774,N_3609,N_2622);
nand U3775 (N_3775,N_3448,N_3447);
and U3776 (N_3776,N_3281,N_2826);
xor U3777 (N_3777,N_2804,N_2509);
and U3778 (N_3778,N_3719,N_2927);
nand U3779 (N_3779,N_3386,N_3581);
xor U3780 (N_3780,N_3302,N_3616);
and U3781 (N_3781,N_3741,N_3547);
or U3782 (N_3782,N_2749,N_3702);
and U3783 (N_3783,N_3349,N_3731);
and U3784 (N_3784,N_3267,N_2549);
nand U3785 (N_3785,N_3587,N_2620);
xor U3786 (N_3786,N_3605,N_2913);
or U3787 (N_3787,N_3486,N_3107);
xor U3788 (N_3788,N_2722,N_3318);
or U3789 (N_3789,N_2829,N_3357);
and U3790 (N_3790,N_3394,N_2925);
or U3791 (N_3791,N_3663,N_2791);
and U3792 (N_3792,N_2923,N_3571);
nand U3793 (N_3793,N_3660,N_3279);
nor U3794 (N_3794,N_3259,N_2848);
nor U3795 (N_3795,N_3230,N_3191);
or U3796 (N_3796,N_3740,N_3113);
and U3797 (N_3797,N_3375,N_3294);
and U3798 (N_3798,N_2900,N_3734);
xnor U3799 (N_3799,N_3028,N_3655);
nand U3800 (N_3800,N_3128,N_2685);
nor U3801 (N_3801,N_3261,N_3181);
nor U3802 (N_3802,N_3542,N_2841);
xor U3803 (N_3803,N_2914,N_2763);
nor U3804 (N_3804,N_2892,N_3101);
nand U3805 (N_3805,N_3201,N_3334);
nand U3806 (N_3806,N_2642,N_2952);
nand U3807 (N_3807,N_3732,N_3661);
nand U3808 (N_3808,N_2702,N_2592);
xnor U3809 (N_3809,N_2717,N_3133);
or U3810 (N_3810,N_2545,N_3317);
nor U3811 (N_3811,N_3724,N_3194);
or U3812 (N_3812,N_2566,N_3511);
or U3813 (N_3813,N_2714,N_3109);
nand U3814 (N_3814,N_2971,N_3159);
and U3815 (N_3815,N_2612,N_3610);
xor U3816 (N_3816,N_3460,N_3435);
xor U3817 (N_3817,N_3440,N_3182);
and U3818 (N_3818,N_3411,N_3033);
and U3819 (N_3819,N_3502,N_3630);
xnor U3820 (N_3820,N_3568,N_3672);
xor U3821 (N_3821,N_3627,N_2764);
and U3822 (N_3822,N_2823,N_2861);
or U3823 (N_3823,N_2983,N_3429);
nor U3824 (N_3824,N_3102,N_3353);
xnor U3825 (N_3825,N_3369,N_2931);
nor U3826 (N_3826,N_2856,N_3108);
nand U3827 (N_3827,N_3141,N_2740);
or U3828 (N_3828,N_3470,N_3255);
nor U3829 (N_3829,N_3703,N_2785);
and U3830 (N_3830,N_3152,N_2725);
nand U3831 (N_3831,N_2524,N_3584);
nor U3832 (N_3832,N_3254,N_3580);
nor U3833 (N_3833,N_3077,N_3260);
nor U3834 (N_3834,N_3166,N_3193);
nand U3835 (N_3835,N_3052,N_3468);
nand U3836 (N_3836,N_3250,N_3171);
or U3837 (N_3837,N_2845,N_2628);
nor U3838 (N_3838,N_2796,N_3023);
nand U3839 (N_3839,N_3197,N_3292);
or U3840 (N_3840,N_2648,N_3258);
nor U3841 (N_3841,N_3327,N_3218);
nor U3842 (N_3842,N_2575,N_2602);
nand U3843 (N_3843,N_3667,N_3398);
nand U3844 (N_3844,N_3325,N_3482);
nor U3845 (N_3845,N_2599,N_2924);
nor U3846 (N_3846,N_2881,N_2799);
or U3847 (N_3847,N_2586,N_2540);
nand U3848 (N_3848,N_3692,N_2650);
nand U3849 (N_3849,N_3528,N_2916);
xor U3850 (N_3850,N_2662,N_3209);
or U3851 (N_3851,N_3291,N_2994);
xnor U3852 (N_3852,N_3084,N_2526);
or U3853 (N_3853,N_3410,N_2720);
nand U3854 (N_3854,N_3065,N_2865);
nor U3855 (N_3855,N_2898,N_3022);
and U3856 (N_3856,N_2932,N_2572);
nor U3857 (N_3857,N_2786,N_2949);
xnor U3858 (N_3858,N_2552,N_2607);
or U3859 (N_3859,N_3559,N_3539);
nor U3860 (N_3860,N_2767,N_2992);
nand U3861 (N_3861,N_2854,N_2869);
and U3862 (N_3862,N_3381,N_2623);
and U3863 (N_3863,N_3681,N_3224);
nor U3864 (N_3864,N_2681,N_3290);
nor U3865 (N_3865,N_3241,N_3098);
or U3866 (N_3866,N_3729,N_3149);
or U3867 (N_3867,N_2705,N_3355);
nand U3868 (N_3868,N_3376,N_2891);
nor U3869 (N_3869,N_2557,N_3574);
nand U3870 (N_3870,N_2762,N_3705);
or U3871 (N_3871,N_2849,N_3577);
and U3872 (N_3872,N_3481,N_3677);
xor U3873 (N_3873,N_2563,N_3602);
or U3874 (N_3874,N_2525,N_3485);
or U3875 (N_3875,N_3196,N_2649);
nand U3876 (N_3876,N_3745,N_2538);
nor U3877 (N_3877,N_3186,N_3163);
nand U3878 (N_3878,N_2520,N_2930);
nor U3879 (N_3879,N_3306,N_3716);
nand U3880 (N_3880,N_3284,N_3335);
xor U3881 (N_3881,N_3097,N_2911);
and U3882 (N_3882,N_2522,N_3537);
xor U3883 (N_3883,N_2811,N_2656);
and U3884 (N_3884,N_3738,N_2917);
or U3885 (N_3885,N_2839,N_2864);
and U3886 (N_3886,N_3253,N_3348);
and U3887 (N_3887,N_3044,N_2573);
nor U3888 (N_3888,N_2726,N_3229);
and U3889 (N_3889,N_3054,N_3071);
or U3890 (N_3890,N_2544,N_2882);
nor U3891 (N_3891,N_3648,N_3646);
or U3892 (N_3892,N_3220,N_3005);
nand U3893 (N_3893,N_2696,N_3187);
or U3894 (N_3894,N_2735,N_3174);
xor U3895 (N_3895,N_3721,N_2684);
xor U3896 (N_3896,N_3314,N_3695);
nor U3897 (N_3897,N_3222,N_2609);
nand U3898 (N_3898,N_3168,N_3619);
and U3899 (N_3899,N_2974,N_3232);
xnor U3900 (N_3900,N_3089,N_2679);
and U3901 (N_3901,N_2943,N_2666);
or U3902 (N_3902,N_2895,N_3735);
xnor U3903 (N_3903,N_2970,N_3434);
nand U3904 (N_3904,N_2938,N_2588);
or U3905 (N_3905,N_2634,N_3623);
xnor U3906 (N_3906,N_2511,N_3137);
or U3907 (N_3907,N_2514,N_3138);
or U3908 (N_3908,N_2615,N_2537);
or U3909 (N_3909,N_3690,N_3576);
nor U3910 (N_3910,N_3096,N_3343);
nand U3911 (N_3911,N_2993,N_2682);
xor U3912 (N_3912,N_3673,N_3469);
and U3913 (N_3913,N_3236,N_2667);
or U3914 (N_3914,N_2597,N_3013);
xnor U3915 (N_3915,N_2953,N_3503);
or U3916 (N_3916,N_3228,N_3707);
nand U3917 (N_3917,N_2742,N_3175);
nand U3918 (N_3918,N_3134,N_3046);
nand U3919 (N_3919,N_2630,N_3736);
and U3920 (N_3920,N_2738,N_2756);
and U3921 (N_3921,N_3265,N_2523);
or U3922 (N_3922,N_3382,N_2700);
or U3923 (N_3923,N_3536,N_3390);
and U3924 (N_3924,N_2531,N_2871);
and U3925 (N_3925,N_3508,N_3656);
nor U3926 (N_3926,N_3612,N_3472);
or U3927 (N_3927,N_3608,N_3093);
nand U3928 (N_3928,N_2501,N_3387);
nand U3929 (N_3929,N_3216,N_3453);
and U3930 (N_3930,N_2951,N_2670);
xor U3931 (N_3931,N_2577,N_3513);
nor U3932 (N_3932,N_3252,N_2614);
or U3933 (N_3933,N_3017,N_3079);
nand U3934 (N_3934,N_3743,N_3037);
and U3935 (N_3935,N_3304,N_3589);
or U3936 (N_3936,N_2527,N_3564);
nor U3937 (N_3937,N_2761,N_3501);
and U3938 (N_3938,N_3212,N_2939);
nand U3939 (N_3939,N_2975,N_2831);
nand U3940 (N_3940,N_2774,N_2874);
and U3941 (N_3941,N_3670,N_3122);
and U3942 (N_3942,N_3072,N_3286);
or U3943 (N_3943,N_2777,N_3392);
xnor U3944 (N_3944,N_2616,N_2787);
nor U3945 (N_3945,N_3366,N_3523);
nor U3946 (N_3946,N_3653,N_2603);
xnor U3947 (N_3947,N_3517,N_2645);
and U3948 (N_3948,N_2734,N_3056);
and U3949 (N_3949,N_3263,N_2644);
nand U3950 (N_3950,N_3711,N_3395);
nor U3951 (N_3951,N_3590,N_2859);
xor U3952 (N_3952,N_3164,N_3615);
or U3953 (N_3953,N_3678,N_3288);
or U3954 (N_3954,N_2765,N_3035);
and U3955 (N_3955,N_3725,N_3313);
or U3956 (N_3956,N_3078,N_2948);
nand U3957 (N_3957,N_2536,N_3640);
or U3958 (N_3958,N_3051,N_2606);
and U3959 (N_3959,N_3717,N_2584);
or U3960 (N_3960,N_3632,N_3569);
nand U3961 (N_3961,N_3546,N_3362);
or U3962 (N_3962,N_2652,N_2678);
xor U3963 (N_3963,N_3525,N_3591);
nand U3964 (N_3964,N_3300,N_3243);
xor U3965 (N_3965,N_2539,N_2710);
xor U3966 (N_3966,N_2926,N_3720);
xnor U3967 (N_3967,N_3674,N_3328);
nor U3968 (N_3968,N_2736,N_3688);
nor U3969 (N_3969,N_2899,N_2556);
xnor U3970 (N_3970,N_3628,N_3007);
nand U3971 (N_3971,N_3019,N_3682);
or U3972 (N_3972,N_3123,N_3377);
and U3973 (N_3973,N_3700,N_3457);
nor U3974 (N_3974,N_3373,N_2625);
nand U3975 (N_3975,N_3520,N_3699);
nand U3976 (N_3976,N_2530,N_2870);
xnor U3977 (N_3977,N_3199,N_3280);
nor U3978 (N_3978,N_3200,N_2671);
and U3979 (N_3979,N_3103,N_2808);
nor U3980 (N_3980,N_2741,N_2775);
xor U3981 (N_3981,N_3087,N_2886);
xnor U3982 (N_3982,N_3004,N_3074);
xnor U3983 (N_3983,N_3183,N_3247);
and U3984 (N_3984,N_3715,N_3190);
nor U3985 (N_3985,N_2719,N_2550);
nand U3986 (N_3986,N_2825,N_2716);
nor U3987 (N_3987,N_3488,N_2608);
nor U3988 (N_3988,N_2833,N_2877);
xor U3989 (N_3989,N_2535,N_3350);
xor U3990 (N_3990,N_3686,N_3045);
xor U3991 (N_3991,N_3614,N_2835);
nor U3992 (N_3992,N_3425,N_3685);
nor U3993 (N_3993,N_2661,N_3642);
xnor U3994 (N_3994,N_3154,N_3710);
and U3995 (N_3995,N_2941,N_3746);
and U3996 (N_3996,N_3438,N_3049);
or U3997 (N_3997,N_3337,N_3647);
xor U3998 (N_3998,N_2843,N_3728);
nand U3999 (N_3999,N_3421,N_3179);
xor U4000 (N_4000,N_3723,N_3428);
xor U4001 (N_4001,N_2855,N_3322);
nand U4002 (N_4002,N_3323,N_3048);
or U4003 (N_4003,N_2950,N_2554);
nand U4004 (N_4004,N_3006,N_3295);
or U4005 (N_4005,N_3548,N_2807);
xnor U4006 (N_4006,N_2795,N_3203);
nor U4007 (N_4007,N_3050,N_3713);
xnor U4008 (N_4008,N_3586,N_3748);
and U4009 (N_4009,N_3008,N_2824);
and U4010 (N_4010,N_3389,N_2567);
xnor U4011 (N_4011,N_2922,N_3561);
xnor U4012 (N_4012,N_3749,N_3563);
nor U4013 (N_4013,N_3659,N_2707);
nor U4014 (N_4014,N_2915,N_2758);
or U4015 (N_4015,N_3492,N_2688);
or U4016 (N_4016,N_3550,N_3534);
xor U4017 (N_4017,N_2902,N_2770);
and U4018 (N_4018,N_2582,N_3264);
nand U4019 (N_4019,N_3208,N_3336);
or U4020 (N_4020,N_2844,N_3393);
and U4021 (N_4021,N_3319,N_3570);
nand U4022 (N_4022,N_2506,N_3061);
xor U4023 (N_4023,N_3445,N_2691);
nor U4024 (N_4024,N_3240,N_3400);
nand U4025 (N_4025,N_3573,N_2704);
or U4026 (N_4026,N_3622,N_3085);
and U4027 (N_4027,N_3474,N_3706);
nand U4028 (N_4028,N_2885,N_2507);
nand U4029 (N_4029,N_3491,N_2986);
nand U4030 (N_4030,N_2987,N_3634);
xnor U4031 (N_4031,N_2890,N_3148);
nor U4032 (N_4032,N_3683,N_3114);
or U4033 (N_4033,N_3227,N_3518);
or U4034 (N_4034,N_3471,N_2646);
xnor U4035 (N_4035,N_2853,N_2815);
nand U4036 (N_4036,N_3450,N_2789);
nor U4037 (N_4037,N_3494,N_2958);
xnor U4038 (N_4038,N_2565,N_2594);
nor U4039 (N_4039,N_3597,N_2718);
and U4040 (N_4040,N_3297,N_3578);
and U4041 (N_4041,N_2967,N_2706);
nand U4042 (N_4042,N_3709,N_3698);
nor U4043 (N_4043,N_2699,N_3268);
nand U4044 (N_4044,N_2559,N_3324);
nand U4045 (N_4045,N_3385,N_2500);
nand U4046 (N_4046,N_2793,N_3185);
nand U4047 (N_4047,N_3666,N_2940);
nor U4048 (N_4048,N_3636,N_2929);
nand U4049 (N_4049,N_2850,N_2604);
xor U4050 (N_4050,N_2981,N_2832);
nand U4051 (N_4051,N_3371,N_2581);
xor U4052 (N_4052,N_2698,N_3225);
and U4053 (N_4053,N_3426,N_3556);
xnor U4054 (N_4054,N_2748,N_3144);
xor U4055 (N_4055,N_3675,N_2757);
nand U4056 (N_4056,N_3139,N_3372);
or U4057 (N_4057,N_2518,N_3320);
and U4058 (N_4058,N_3730,N_3742);
xnor U4059 (N_4059,N_3431,N_3712);
nor U4060 (N_4060,N_3365,N_3157);
nor U4061 (N_4061,N_3031,N_2600);
xnor U4062 (N_4062,N_2627,N_2827);
or U4063 (N_4063,N_3067,N_2820);
xnor U4064 (N_4064,N_2579,N_3092);
nand U4065 (N_4065,N_3021,N_3572);
xor U4066 (N_4066,N_3315,N_3120);
nor U4067 (N_4067,N_2728,N_2766);
xnor U4068 (N_4068,N_3543,N_3565);
xor U4069 (N_4069,N_2972,N_2904);
xnor U4070 (N_4070,N_3354,N_3257);
and U4071 (N_4071,N_3599,N_2780);
or U4072 (N_4072,N_3364,N_3594);
or U4073 (N_4073,N_3361,N_3088);
nor U4074 (N_4074,N_3697,N_3497);
nor U4075 (N_4075,N_3495,N_2731);
xnor U4076 (N_4076,N_2959,N_3140);
and U4077 (N_4077,N_2921,N_3643);
and U4078 (N_4078,N_3427,N_3237);
or U4079 (N_4079,N_3654,N_2801);
or U4080 (N_4080,N_3125,N_2571);
nor U4081 (N_4081,N_2897,N_3244);
nor U4082 (N_4082,N_3432,N_2574);
and U4083 (N_4083,N_3650,N_2578);
xor U4084 (N_4084,N_3689,N_3370);
xnor U4085 (N_4085,N_2708,N_3451);
or U4086 (N_4086,N_3531,N_2673);
xnor U4087 (N_4087,N_2729,N_3030);
or U4088 (N_4088,N_3652,N_3476);
xor U4089 (N_4089,N_2973,N_3409);
nor U4090 (N_4090,N_2937,N_3423);
nand U4091 (N_4091,N_2703,N_3378);
xnor U4092 (N_4092,N_3223,N_3413);
nor U4093 (N_4093,N_3339,N_2768);
or U4094 (N_4094,N_2590,N_2580);
nand U4095 (N_4095,N_2979,N_3507);
or U4096 (N_4096,N_3239,N_2797);
nand U4097 (N_4097,N_3662,N_3490);
or U4098 (N_4098,N_3676,N_3496);
or U4099 (N_4099,N_3475,N_2908);
xor U4100 (N_4100,N_3283,N_3060);
xnor U4101 (N_4101,N_3277,N_3116);
xnor U4102 (N_4102,N_3701,N_2739);
nand U4103 (N_4103,N_2866,N_3509);
and U4104 (N_4104,N_3064,N_2945);
nand U4105 (N_4105,N_3235,N_2653);
nand U4106 (N_4106,N_3246,N_3463);
or U4107 (N_4107,N_2753,N_2641);
or U4108 (N_4108,N_3043,N_3360);
nor U4109 (N_4109,N_3566,N_3326);
xnor U4110 (N_4110,N_3036,N_3329);
or U4111 (N_4111,N_3532,N_3091);
or U4112 (N_4112,N_3342,N_3330);
nand U4113 (N_4113,N_3204,N_3233);
nor U4114 (N_4114,N_3579,N_3521);
xor U4115 (N_4115,N_3456,N_3003);
and U4116 (N_4116,N_2743,N_3397);
nand U4117 (N_4117,N_3424,N_3069);
and U4118 (N_4118,N_3161,N_3620);
or U4119 (N_4119,N_3744,N_3309);
or U4120 (N_4120,N_3458,N_2966);
xnor U4121 (N_4121,N_3039,N_2880);
nor U4122 (N_4122,N_3301,N_3726);
nor U4123 (N_4123,N_3693,N_2585);
nor U4124 (N_4124,N_3684,N_2956);
nor U4125 (N_4125,N_3242,N_3489);
or U4126 (N_4126,N_3226,N_2689);
and U4127 (N_4127,N_2860,N_2813);
nor U4128 (N_4128,N_2806,N_2711);
or U4129 (N_4129,N_2677,N_3526);
or U4130 (N_4130,N_3407,N_2905);
nand U4131 (N_4131,N_2773,N_3680);
nand U4132 (N_4132,N_3073,N_3178);
nor U4133 (N_4133,N_2990,N_2805);
nand U4134 (N_4134,N_2555,N_3063);
and U4135 (N_4135,N_3635,N_3665);
or U4136 (N_4136,N_3195,N_3638);
nand U4137 (N_4137,N_3156,N_3132);
nor U4138 (N_4138,N_3346,N_2894);
and U4139 (N_4139,N_3639,N_3285);
nor U4140 (N_4140,N_3047,N_2638);
nand U4141 (N_4141,N_3271,N_3436);
xor U4142 (N_4142,N_3131,N_3145);
or U4143 (N_4143,N_3505,N_2989);
nor U4144 (N_4144,N_3025,N_3419);
xnor U4145 (N_4145,N_2790,N_2942);
and U4146 (N_4146,N_3188,N_3691);
nor U4147 (N_4147,N_2611,N_3206);
xor U4148 (N_4148,N_3549,N_2794);
nor U4149 (N_4149,N_3504,N_2639);
or U4150 (N_4150,N_3529,N_3379);
nor U4151 (N_4151,N_3273,N_3538);
xor U4152 (N_4152,N_3351,N_2997);
nand U4153 (N_4153,N_3142,N_3384);
nor U4154 (N_4154,N_2760,N_2746);
nor U4155 (N_4155,N_3015,N_3624);
or U4156 (N_4156,N_3664,N_3582);
xor U4157 (N_4157,N_2977,N_3461);
nand U4158 (N_4158,N_2985,N_3617);
nor U4159 (N_4159,N_3210,N_2818);
or U4160 (N_4160,N_3135,N_3487);
and U4161 (N_4161,N_2548,N_3452);
nand U4162 (N_4162,N_3514,N_3739);
xnor U4163 (N_4163,N_3100,N_2876);
nand U4164 (N_4164,N_2919,N_3041);
nor U4165 (N_4165,N_2846,N_2553);
nor U4166 (N_4166,N_3213,N_2784);
xor U4167 (N_4167,N_3299,N_2814);
nor U4168 (N_4168,N_3066,N_3585);
and U4169 (N_4169,N_3180,N_2995);
or U4170 (N_4170,N_3147,N_3310);
and U4171 (N_4171,N_3173,N_3708);
and U4172 (N_4172,N_2654,N_2512);
nor U4173 (N_4173,N_3014,N_3668);
or U4174 (N_4174,N_2683,N_3245);
nor U4175 (N_4175,N_3406,N_2732);
xor U4176 (N_4176,N_3455,N_3551);
and U4177 (N_4177,N_3422,N_3669);
or U4178 (N_4178,N_2631,N_3626);
or U4179 (N_4179,N_2991,N_3303);
xor U4180 (N_4180,N_2605,N_2664);
nand U4181 (N_4181,N_2830,N_2516);
nor U4182 (N_4182,N_2663,N_2884);
and U4183 (N_4183,N_3401,N_2800);
nand U4184 (N_4184,N_2968,N_3115);
nor U4185 (N_4185,N_3058,N_3408);
xor U4186 (N_4186,N_3657,N_3296);
nand U4187 (N_4187,N_3256,N_2858);
and U4188 (N_4188,N_2637,N_3557);
or U4189 (N_4189,N_3625,N_3266);
nor U4190 (N_4190,N_2647,N_3544);
or U4191 (N_4191,N_3075,N_3444);
xnor U4192 (N_4192,N_3024,N_2798);
nand U4193 (N_4193,N_3433,N_3198);
nand U4194 (N_4194,N_2984,N_2840);
or U4195 (N_4195,N_2660,N_2542);
and U4196 (N_4196,N_2669,N_3106);
nor U4197 (N_4197,N_2505,N_2635);
nor U4198 (N_4198,N_2519,N_3649);
and U4199 (N_4199,N_3053,N_3443);
nor U4200 (N_4200,N_3276,N_3172);
xor U4201 (N_4201,N_2873,N_3344);
nor U4202 (N_4202,N_2562,N_2532);
and U4203 (N_4203,N_2933,N_3333);
xor U4204 (N_4204,N_2624,N_2836);
nand U4205 (N_4205,N_2998,N_3519);
nor U4206 (N_4206,N_2788,N_2619);
nand U4207 (N_4207,N_3633,N_3417);
and U4208 (N_4208,N_3070,N_3465);
nor U4209 (N_4209,N_3151,N_3032);
or U4210 (N_4210,N_2693,N_2883);
xor U4211 (N_4211,N_2629,N_3307);
and U4212 (N_4212,N_3391,N_3117);
nor U4213 (N_4213,N_3205,N_2515);
or U4214 (N_4214,N_3462,N_3441);
or U4215 (N_4215,N_2910,N_3510);
nand U4216 (N_4216,N_2715,N_2965);
nor U4217 (N_4217,N_3165,N_3221);
xor U4218 (N_4218,N_3160,N_3083);
xnor U4219 (N_4219,N_3118,N_2513);
nand U4220 (N_4220,N_3026,N_3418);
nand U4221 (N_4221,N_3499,N_2621);
and U4222 (N_4222,N_3484,N_3112);
xnor U4223 (N_4223,N_2517,N_3176);
nor U4224 (N_4224,N_3631,N_2751);
nand U4225 (N_4225,N_2962,N_3483);
xor U4226 (N_4226,N_3234,N_3402);
xnor U4227 (N_4227,N_2680,N_2838);
or U4228 (N_4228,N_2863,N_3057);
or U4229 (N_4229,N_3020,N_3545);
nor U4230 (N_4230,N_2857,N_2591);
nor U4231 (N_4231,N_2901,N_3356);
nand U4232 (N_4232,N_2821,N_2954);
or U4233 (N_4233,N_3403,N_3090);
xor U4234 (N_4234,N_3001,N_2564);
nand U4235 (N_4235,N_3012,N_3217);
xor U4236 (N_4236,N_2782,N_2744);
nor U4237 (N_4237,N_3104,N_2534);
or U4238 (N_4238,N_2802,N_3516);
xnor U4239 (N_4239,N_2508,N_2551);
nand U4240 (N_4240,N_3321,N_3583);
nor U4241 (N_4241,N_2934,N_3153);
xnor U4242 (N_4242,N_3311,N_3042);
xor U4243 (N_4243,N_2783,N_2817);
nand U4244 (N_4244,N_2547,N_2976);
xnor U4245 (N_4245,N_2721,N_2893);
xor U4246 (N_4246,N_3601,N_3553);
xor U4247 (N_4247,N_3368,N_2961);
nand U4248 (N_4248,N_2906,N_2842);
nor U4249 (N_4249,N_2947,N_3524);
nor U4250 (N_4250,N_2503,N_3383);
nand U4251 (N_4251,N_3238,N_3251);
or U4252 (N_4252,N_2963,N_3119);
or U4253 (N_4253,N_3416,N_2960);
nor U4254 (N_4254,N_3270,N_3136);
nand U4255 (N_4255,N_3658,N_3679);
nand U4256 (N_4256,N_2822,N_3002);
and U4257 (N_4257,N_3437,N_3733);
or U4258 (N_4258,N_3298,N_2724);
or U4259 (N_4259,N_3718,N_3081);
nand U4260 (N_4260,N_3169,N_2676);
or U4261 (N_4261,N_3466,N_3530);
nor U4262 (N_4262,N_2819,N_3687);
or U4263 (N_4263,N_3010,N_3500);
xnor U4264 (N_4264,N_2558,N_3641);
or U4265 (N_4265,N_3027,N_3515);
and U4266 (N_4266,N_2695,N_2709);
and U4267 (N_4267,N_3595,N_2867);
xor U4268 (N_4268,N_3287,N_2803);
and U4269 (N_4269,N_3527,N_2543);
xor U4270 (N_4270,N_3312,N_2828);
xnor U4271 (N_4271,N_2888,N_3192);
nand U4272 (N_4272,N_2851,N_3305);
nand U4273 (N_4273,N_3080,N_3396);
and U4274 (N_4274,N_2810,N_2847);
nand U4275 (N_4275,N_3480,N_2589);
nand U4276 (N_4276,N_2792,N_3127);
or U4277 (N_4277,N_3099,N_2988);
or U4278 (N_4278,N_3367,N_3111);
or U4279 (N_4279,N_3430,N_3737);
and U4280 (N_4280,N_3446,N_2754);
or U4281 (N_4281,N_2529,N_2982);
xnor U4282 (N_4282,N_2598,N_2755);
or U4283 (N_4283,N_3016,N_3621);
nor U4284 (N_4284,N_3562,N_3506);
or U4285 (N_4285,N_3645,N_2694);
nor U4286 (N_4286,N_2776,N_3167);
nor U4287 (N_4287,N_3604,N_2816);
nor U4288 (N_4288,N_3143,N_3308);
nand U4289 (N_4289,N_2618,N_2752);
nor U4290 (N_4290,N_3009,N_2659);
xnor U4291 (N_4291,N_3449,N_3512);
or U4292 (N_4292,N_2996,N_3554);
nand U4293 (N_4293,N_3533,N_2674);
or U4294 (N_4294,N_2903,N_2665);
nor U4295 (N_4295,N_2533,N_2907);
nor U4296 (N_4296,N_3603,N_3560);
and U4297 (N_4297,N_2759,N_2779);
or U4298 (N_4298,N_2686,N_3121);
nand U4299 (N_4299,N_2587,N_2936);
nor U4300 (N_4300,N_3600,N_3374);
nand U4301 (N_4301,N_3331,N_3076);
or U4302 (N_4302,N_3293,N_2583);
nor U4303 (N_4303,N_2636,N_3558);
or U4304 (N_4304,N_3207,N_3040);
and U4305 (N_4305,N_3278,N_2713);
xnor U4306 (N_4306,N_2651,N_3341);
xnor U4307 (N_4307,N_2502,N_3110);
xnor U4308 (N_4308,N_2712,N_2778);
nand U4309 (N_4309,N_3442,N_3211);
or U4310 (N_4310,N_3479,N_3214);
nor U4311 (N_4311,N_3155,N_3363);
nand U4312 (N_4312,N_3464,N_3352);
and U4313 (N_4313,N_2809,N_3274);
xor U4314 (N_4314,N_3380,N_3588);
or U4315 (N_4315,N_2912,N_3493);
nand U4316 (N_4316,N_2601,N_3000);
or U4317 (N_4317,N_2701,N_3055);
xnor U4318 (N_4318,N_3555,N_2546);
xor U4319 (N_4319,N_3727,N_3162);
nand U4320 (N_4320,N_3575,N_2687);
or U4321 (N_4321,N_3231,N_3029);
nor U4322 (N_4322,N_3522,N_2772);
xor U4323 (N_4323,N_3414,N_3637);
xnor U4324 (N_4324,N_3272,N_3611);
and U4325 (N_4325,N_3405,N_2593);
and U4326 (N_4326,N_3189,N_3059);
nand U4327 (N_4327,N_3415,N_2862);
nor U4328 (N_4328,N_3454,N_3170);
or U4329 (N_4329,N_2750,N_3332);
xnor U4330 (N_4330,N_3540,N_2528);
xor U4331 (N_4331,N_3613,N_3034);
xnor U4332 (N_4332,N_3094,N_3473);
xor U4333 (N_4333,N_2510,N_2632);
or U4334 (N_4334,N_3338,N_3150);
nor U4335 (N_4335,N_3018,N_3478);
nor U4336 (N_4336,N_3038,N_3722);
nand U4337 (N_4337,N_3388,N_3262);
and U4338 (N_4338,N_3124,N_2946);
and U4339 (N_4339,N_2521,N_3275);
xor U4340 (N_4340,N_2626,N_2561);
xor U4341 (N_4341,N_2868,N_3412);
xnor U4342 (N_4342,N_3747,N_3606);
nor U4343 (N_4343,N_3130,N_2978);
nand U4344 (N_4344,N_3593,N_3671);
or U4345 (N_4345,N_3126,N_3215);
nor U4346 (N_4346,N_3068,N_2969);
or U4347 (N_4347,N_3694,N_3404);
and U4348 (N_4348,N_2957,N_3249);
or U4349 (N_4349,N_2769,N_2944);
nand U4350 (N_4350,N_2655,N_2879);
or U4351 (N_4351,N_3459,N_2697);
and U4352 (N_4352,N_3095,N_3439);
or U4353 (N_4353,N_2875,N_3618);
or U4354 (N_4354,N_3219,N_3316);
nor U4355 (N_4355,N_2812,N_2643);
nor U4356 (N_4356,N_3714,N_3399);
nand U4357 (N_4357,N_3607,N_2733);
or U4358 (N_4358,N_2852,N_2955);
xor U4359 (N_4359,N_3289,N_2675);
nor U4360 (N_4360,N_3359,N_3129);
nor U4361 (N_4361,N_3567,N_2837);
nand U4362 (N_4362,N_3158,N_3704);
nand U4363 (N_4363,N_2569,N_2723);
xor U4364 (N_4364,N_2692,N_3248);
nor U4365 (N_4365,N_2964,N_3644);
or U4366 (N_4366,N_2658,N_2747);
nor U4367 (N_4367,N_2737,N_2727);
xor U4368 (N_4368,N_2504,N_3177);
or U4369 (N_4369,N_2771,N_2613);
xor U4370 (N_4370,N_3596,N_2896);
and U4371 (N_4371,N_2909,N_2878);
xnor U4372 (N_4372,N_3629,N_2745);
nor U4373 (N_4373,N_2570,N_3062);
and U4374 (N_4374,N_2920,N_3340);
xnor U4375 (N_4375,N_2915,N_2640);
nor U4376 (N_4376,N_2605,N_3364);
nand U4377 (N_4377,N_2688,N_3660);
or U4378 (N_4378,N_3104,N_3245);
or U4379 (N_4379,N_3570,N_2719);
xor U4380 (N_4380,N_3330,N_3684);
or U4381 (N_4381,N_2837,N_2646);
xnor U4382 (N_4382,N_2817,N_2971);
and U4383 (N_4383,N_2546,N_3403);
nor U4384 (N_4384,N_3441,N_3717);
xor U4385 (N_4385,N_3252,N_2855);
nor U4386 (N_4386,N_2637,N_3322);
nor U4387 (N_4387,N_3571,N_2645);
or U4388 (N_4388,N_3363,N_3582);
or U4389 (N_4389,N_3307,N_3038);
or U4390 (N_4390,N_3449,N_3546);
and U4391 (N_4391,N_3511,N_3402);
and U4392 (N_4392,N_2757,N_3707);
and U4393 (N_4393,N_2968,N_3155);
and U4394 (N_4394,N_3231,N_2538);
nor U4395 (N_4395,N_2893,N_3280);
nor U4396 (N_4396,N_3584,N_2814);
and U4397 (N_4397,N_3357,N_3493);
xor U4398 (N_4398,N_3302,N_3045);
nor U4399 (N_4399,N_3020,N_3199);
xnor U4400 (N_4400,N_2924,N_3365);
xor U4401 (N_4401,N_2863,N_2564);
nand U4402 (N_4402,N_2579,N_3005);
xor U4403 (N_4403,N_3277,N_3728);
or U4404 (N_4404,N_3460,N_3160);
or U4405 (N_4405,N_3339,N_2810);
and U4406 (N_4406,N_3590,N_2705);
xnor U4407 (N_4407,N_2865,N_3380);
nand U4408 (N_4408,N_3568,N_3630);
or U4409 (N_4409,N_3273,N_3396);
xor U4410 (N_4410,N_2571,N_3715);
nor U4411 (N_4411,N_3505,N_3616);
or U4412 (N_4412,N_2925,N_3152);
or U4413 (N_4413,N_2809,N_3673);
and U4414 (N_4414,N_3708,N_2962);
nand U4415 (N_4415,N_2888,N_3398);
nor U4416 (N_4416,N_3495,N_3668);
nand U4417 (N_4417,N_2909,N_2573);
or U4418 (N_4418,N_2538,N_3316);
or U4419 (N_4419,N_3409,N_3200);
nor U4420 (N_4420,N_2847,N_3728);
xnor U4421 (N_4421,N_3547,N_2929);
nor U4422 (N_4422,N_2694,N_3145);
nand U4423 (N_4423,N_2934,N_3547);
nand U4424 (N_4424,N_3682,N_3187);
nor U4425 (N_4425,N_2727,N_2689);
nand U4426 (N_4426,N_2938,N_2656);
or U4427 (N_4427,N_2746,N_3735);
nor U4428 (N_4428,N_3012,N_2769);
nor U4429 (N_4429,N_2682,N_2967);
nor U4430 (N_4430,N_2635,N_3436);
and U4431 (N_4431,N_2740,N_3458);
or U4432 (N_4432,N_2720,N_2653);
nor U4433 (N_4433,N_2549,N_2945);
or U4434 (N_4434,N_3577,N_3739);
or U4435 (N_4435,N_3069,N_3565);
and U4436 (N_4436,N_2617,N_2726);
xor U4437 (N_4437,N_3550,N_3571);
or U4438 (N_4438,N_2561,N_3504);
xnor U4439 (N_4439,N_3452,N_2925);
and U4440 (N_4440,N_2598,N_2838);
nor U4441 (N_4441,N_2856,N_2987);
and U4442 (N_4442,N_2944,N_2733);
nand U4443 (N_4443,N_2635,N_2793);
xor U4444 (N_4444,N_3479,N_3660);
xnor U4445 (N_4445,N_3353,N_2693);
nand U4446 (N_4446,N_2915,N_3708);
xnor U4447 (N_4447,N_3531,N_2541);
nand U4448 (N_4448,N_3560,N_3441);
nor U4449 (N_4449,N_3739,N_3479);
xnor U4450 (N_4450,N_2810,N_3276);
and U4451 (N_4451,N_2872,N_3676);
nor U4452 (N_4452,N_3059,N_2548);
nor U4453 (N_4453,N_3631,N_2940);
nor U4454 (N_4454,N_2931,N_3116);
and U4455 (N_4455,N_2874,N_2575);
nor U4456 (N_4456,N_2620,N_3525);
and U4457 (N_4457,N_3225,N_3273);
nand U4458 (N_4458,N_2564,N_2596);
or U4459 (N_4459,N_2688,N_3106);
nand U4460 (N_4460,N_2873,N_3645);
xnor U4461 (N_4461,N_3120,N_3493);
xnor U4462 (N_4462,N_3395,N_3238);
xor U4463 (N_4463,N_3172,N_3092);
and U4464 (N_4464,N_3491,N_3067);
and U4465 (N_4465,N_3094,N_2721);
or U4466 (N_4466,N_3135,N_3716);
and U4467 (N_4467,N_3046,N_2784);
nor U4468 (N_4468,N_2748,N_2919);
and U4469 (N_4469,N_2719,N_2929);
and U4470 (N_4470,N_3238,N_3159);
nor U4471 (N_4471,N_2599,N_2793);
xor U4472 (N_4472,N_3544,N_2869);
xor U4473 (N_4473,N_3575,N_2751);
nor U4474 (N_4474,N_2562,N_3034);
and U4475 (N_4475,N_2692,N_3455);
nor U4476 (N_4476,N_2614,N_3625);
nor U4477 (N_4477,N_3689,N_3416);
xnor U4478 (N_4478,N_3524,N_2546);
xnor U4479 (N_4479,N_3212,N_3591);
nand U4480 (N_4480,N_2622,N_3386);
xor U4481 (N_4481,N_2932,N_3415);
or U4482 (N_4482,N_3679,N_3744);
xor U4483 (N_4483,N_3396,N_3333);
xnor U4484 (N_4484,N_3265,N_3283);
and U4485 (N_4485,N_2650,N_3591);
nand U4486 (N_4486,N_3302,N_2783);
nor U4487 (N_4487,N_2789,N_3156);
nand U4488 (N_4488,N_3134,N_2779);
and U4489 (N_4489,N_2506,N_3689);
nor U4490 (N_4490,N_3531,N_3699);
or U4491 (N_4491,N_3047,N_3553);
and U4492 (N_4492,N_3472,N_3622);
nand U4493 (N_4493,N_2580,N_2832);
or U4494 (N_4494,N_3094,N_3033);
xnor U4495 (N_4495,N_2817,N_2906);
or U4496 (N_4496,N_2545,N_2701);
xnor U4497 (N_4497,N_2904,N_3674);
nor U4498 (N_4498,N_3399,N_2753);
and U4499 (N_4499,N_3301,N_2881);
xor U4500 (N_4500,N_3474,N_2940);
or U4501 (N_4501,N_3056,N_3422);
nor U4502 (N_4502,N_3596,N_2972);
and U4503 (N_4503,N_3327,N_2851);
nor U4504 (N_4504,N_2962,N_2868);
xnor U4505 (N_4505,N_3036,N_3516);
nor U4506 (N_4506,N_2720,N_3651);
xnor U4507 (N_4507,N_2580,N_2973);
or U4508 (N_4508,N_3587,N_3073);
or U4509 (N_4509,N_3127,N_2524);
and U4510 (N_4510,N_2910,N_2806);
and U4511 (N_4511,N_2579,N_3537);
xor U4512 (N_4512,N_3445,N_3334);
nor U4513 (N_4513,N_3239,N_2530);
or U4514 (N_4514,N_2832,N_2520);
xnor U4515 (N_4515,N_3187,N_2771);
or U4516 (N_4516,N_2907,N_2633);
xnor U4517 (N_4517,N_2638,N_2811);
or U4518 (N_4518,N_2607,N_2927);
nor U4519 (N_4519,N_3335,N_3415);
or U4520 (N_4520,N_2946,N_3082);
or U4521 (N_4521,N_3143,N_2761);
or U4522 (N_4522,N_3577,N_3235);
nor U4523 (N_4523,N_3159,N_3032);
nand U4524 (N_4524,N_3244,N_3283);
or U4525 (N_4525,N_2976,N_3467);
xor U4526 (N_4526,N_3723,N_2552);
xnor U4527 (N_4527,N_3732,N_3169);
nand U4528 (N_4528,N_2794,N_3220);
or U4529 (N_4529,N_3335,N_2939);
nor U4530 (N_4530,N_3268,N_3494);
nor U4531 (N_4531,N_2980,N_3061);
or U4532 (N_4532,N_2695,N_2750);
xor U4533 (N_4533,N_3497,N_3514);
and U4534 (N_4534,N_3317,N_3568);
nor U4535 (N_4535,N_2889,N_2702);
or U4536 (N_4536,N_2952,N_3154);
or U4537 (N_4537,N_2739,N_3431);
and U4538 (N_4538,N_2569,N_2558);
and U4539 (N_4539,N_3688,N_2724);
nor U4540 (N_4540,N_2652,N_2619);
nor U4541 (N_4541,N_3145,N_2733);
and U4542 (N_4542,N_2771,N_3583);
xor U4543 (N_4543,N_3402,N_3564);
nand U4544 (N_4544,N_2673,N_3164);
xnor U4545 (N_4545,N_3704,N_3680);
nand U4546 (N_4546,N_3685,N_3694);
nor U4547 (N_4547,N_2845,N_2584);
nor U4548 (N_4548,N_2983,N_2744);
nand U4549 (N_4549,N_3343,N_3562);
nor U4550 (N_4550,N_3413,N_3524);
xor U4551 (N_4551,N_2644,N_3038);
and U4552 (N_4552,N_2873,N_3532);
xor U4553 (N_4553,N_3567,N_3684);
or U4554 (N_4554,N_2835,N_3463);
nand U4555 (N_4555,N_3096,N_3011);
nor U4556 (N_4556,N_2956,N_2538);
or U4557 (N_4557,N_3243,N_2653);
nand U4558 (N_4558,N_3157,N_3537);
or U4559 (N_4559,N_3240,N_3271);
and U4560 (N_4560,N_3572,N_3371);
nor U4561 (N_4561,N_3613,N_3686);
or U4562 (N_4562,N_2692,N_2573);
xor U4563 (N_4563,N_2579,N_2576);
xor U4564 (N_4564,N_3611,N_2707);
nor U4565 (N_4565,N_3612,N_3271);
xnor U4566 (N_4566,N_3567,N_3145);
nand U4567 (N_4567,N_3581,N_3637);
xor U4568 (N_4568,N_3628,N_3728);
xor U4569 (N_4569,N_3380,N_2570);
nor U4570 (N_4570,N_2550,N_2873);
nand U4571 (N_4571,N_3413,N_3280);
xor U4572 (N_4572,N_2560,N_2945);
nand U4573 (N_4573,N_3255,N_2508);
nor U4574 (N_4574,N_3677,N_3672);
or U4575 (N_4575,N_2797,N_3063);
and U4576 (N_4576,N_3678,N_3748);
nor U4577 (N_4577,N_3469,N_3737);
and U4578 (N_4578,N_3571,N_2516);
nor U4579 (N_4579,N_2769,N_3270);
xor U4580 (N_4580,N_3311,N_3546);
or U4581 (N_4581,N_2544,N_2538);
nor U4582 (N_4582,N_3246,N_2816);
nand U4583 (N_4583,N_3498,N_3501);
nand U4584 (N_4584,N_2612,N_2574);
xnor U4585 (N_4585,N_3067,N_2933);
nand U4586 (N_4586,N_2640,N_3069);
nor U4587 (N_4587,N_2513,N_3123);
or U4588 (N_4588,N_3251,N_2692);
nand U4589 (N_4589,N_3748,N_3700);
xnor U4590 (N_4590,N_2986,N_3369);
and U4591 (N_4591,N_3031,N_3148);
nor U4592 (N_4592,N_3090,N_3264);
nor U4593 (N_4593,N_3626,N_3679);
xnor U4594 (N_4594,N_3463,N_2964);
nor U4595 (N_4595,N_3538,N_3126);
and U4596 (N_4596,N_3665,N_2803);
nand U4597 (N_4597,N_2515,N_3119);
or U4598 (N_4598,N_3602,N_3016);
and U4599 (N_4599,N_2930,N_3740);
nor U4600 (N_4600,N_2778,N_3673);
or U4601 (N_4601,N_2897,N_3344);
xnor U4602 (N_4602,N_3587,N_2684);
nand U4603 (N_4603,N_2653,N_2713);
nand U4604 (N_4604,N_3149,N_3089);
nor U4605 (N_4605,N_3023,N_2983);
or U4606 (N_4606,N_3220,N_2835);
or U4607 (N_4607,N_3523,N_3650);
xor U4608 (N_4608,N_2891,N_2808);
nor U4609 (N_4609,N_3456,N_3482);
or U4610 (N_4610,N_2686,N_3327);
nand U4611 (N_4611,N_3172,N_3258);
nand U4612 (N_4612,N_3570,N_3029);
xnor U4613 (N_4613,N_2833,N_2862);
and U4614 (N_4614,N_2933,N_3229);
nand U4615 (N_4615,N_3374,N_3183);
nand U4616 (N_4616,N_2986,N_2753);
and U4617 (N_4617,N_2665,N_3745);
xor U4618 (N_4618,N_2525,N_2909);
nor U4619 (N_4619,N_2852,N_2578);
xnor U4620 (N_4620,N_3708,N_2992);
xnor U4621 (N_4621,N_2841,N_3685);
and U4622 (N_4622,N_3576,N_3464);
nand U4623 (N_4623,N_3340,N_2847);
nor U4624 (N_4624,N_3113,N_3497);
xor U4625 (N_4625,N_3332,N_3479);
xor U4626 (N_4626,N_3039,N_3487);
xor U4627 (N_4627,N_3704,N_3007);
nand U4628 (N_4628,N_3089,N_2572);
or U4629 (N_4629,N_3431,N_2516);
xnor U4630 (N_4630,N_3120,N_3516);
nand U4631 (N_4631,N_2660,N_2864);
xor U4632 (N_4632,N_3019,N_2539);
or U4633 (N_4633,N_2508,N_3265);
and U4634 (N_4634,N_3128,N_2637);
or U4635 (N_4635,N_3428,N_3469);
and U4636 (N_4636,N_2853,N_2949);
xnor U4637 (N_4637,N_2789,N_3633);
and U4638 (N_4638,N_3484,N_3614);
and U4639 (N_4639,N_2600,N_3427);
and U4640 (N_4640,N_3540,N_3463);
nand U4641 (N_4641,N_3648,N_2806);
and U4642 (N_4642,N_3446,N_3746);
nand U4643 (N_4643,N_2887,N_3272);
xor U4644 (N_4644,N_3201,N_3180);
xnor U4645 (N_4645,N_3164,N_2611);
nand U4646 (N_4646,N_3698,N_3351);
xor U4647 (N_4647,N_3572,N_3139);
xnor U4648 (N_4648,N_2874,N_3130);
xnor U4649 (N_4649,N_2630,N_3479);
xnor U4650 (N_4650,N_3115,N_2909);
xor U4651 (N_4651,N_3522,N_2710);
nor U4652 (N_4652,N_2843,N_3749);
xnor U4653 (N_4653,N_2672,N_3124);
nand U4654 (N_4654,N_3021,N_3673);
nor U4655 (N_4655,N_2563,N_2731);
and U4656 (N_4656,N_3285,N_3279);
and U4657 (N_4657,N_3715,N_2849);
xnor U4658 (N_4658,N_3188,N_2520);
nand U4659 (N_4659,N_2895,N_2569);
and U4660 (N_4660,N_2915,N_3255);
or U4661 (N_4661,N_2586,N_3716);
nand U4662 (N_4662,N_3166,N_2989);
xor U4663 (N_4663,N_2926,N_3154);
nor U4664 (N_4664,N_2669,N_3570);
nor U4665 (N_4665,N_2582,N_3150);
xor U4666 (N_4666,N_3257,N_3737);
xor U4667 (N_4667,N_3441,N_3120);
nor U4668 (N_4668,N_2776,N_3724);
nand U4669 (N_4669,N_2585,N_3406);
nand U4670 (N_4670,N_3609,N_3211);
xnor U4671 (N_4671,N_2639,N_2653);
or U4672 (N_4672,N_2977,N_2966);
xor U4673 (N_4673,N_2591,N_2704);
and U4674 (N_4674,N_3331,N_3381);
or U4675 (N_4675,N_2791,N_3382);
and U4676 (N_4676,N_2996,N_3400);
and U4677 (N_4677,N_3439,N_2876);
xor U4678 (N_4678,N_3673,N_3258);
or U4679 (N_4679,N_2912,N_2997);
nor U4680 (N_4680,N_3641,N_3540);
xnor U4681 (N_4681,N_2585,N_3606);
nand U4682 (N_4682,N_3654,N_3204);
nor U4683 (N_4683,N_3597,N_3638);
nand U4684 (N_4684,N_3386,N_2641);
nor U4685 (N_4685,N_2665,N_2810);
nand U4686 (N_4686,N_3251,N_3184);
and U4687 (N_4687,N_2729,N_3676);
nand U4688 (N_4688,N_2723,N_2843);
nor U4689 (N_4689,N_2930,N_2567);
nand U4690 (N_4690,N_2554,N_3074);
nand U4691 (N_4691,N_3298,N_3292);
nor U4692 (N_4692,N_2781,N_3311);
or U4693 (N_4693,N_3022,N_2796);
or U4694 (N_4694,N_2638,N_2822);
xnor U4695 (N_4695,N_2687,N_2530);
nand U4696 (N_4696,N_3063,N_3611);
xor U4697 (N_4697,N_2834,N_3145);
nor U4698 (N_4698,N_3145,N_2862);
or U4699 (N_4699,N_2756,N_2553);
nor U4700 (N_4700,N_3231,N_3045);
xnor U4701 (N_4701,N_3528,N_3359);
nor U4702 (N_4702,N_2583,N_3168);
xnor U4703 (N_4703,N_3647,N_2914);
or U4704 (N_4704,N_2900,N_3049);
or U4705 (N_4705,N_2594,N_3666);
nor U4706 (N_4706,N_2736,N_2501);
nor U4707 (N_4707,N_2926,N_2876);
xnor U4708 (N_4708,N_3602,N_3287);
and U4709 (N_4709,N_3679,N_3556);
xor U4710 (N_4710,N_3579,N_2750);
nand U4711 (N_4711,N_3073,N_2971);
or U4712 (N_4712,N_2639,N_3558);
nor U4713 (N_4713,N_2845,N_3155);
nor U4714 (N_4714,N_3281,N_3467);
or U4715 (N_4715,N_3410,N_2508);
and U4716 (N_4716,N_2820,N_3240);
and U4717 (N_4717,N_2838,N_3368);
and U4718 (N_4718,N_2708,N_2583);
nand U4719 (N_4719,N_2625,N_2892);
nor U4720 (N_4720,N_3056,N_2623);
or U4721 (N_4721,N_3492,N_3410);
or U4722 (N_4722,N_2685,N_3695);
xor U4723 (N_4723,N_2553,N_3704);
xor U4724 (N_4724,N_3452,N_3278);
nand U4725 (N_4725,N_3180,N_3064);
and U4726 (N_4726,N_2710,N_2756);
xor U4727 (N_4727,N_3291,N_3535);
and U4728 (N_4728,N_2693,N_2919);
and U4729 (N_4729,N_3444,N_3614);
and U4730 (N_4730,N_2536,N_3222);
nor U4731 (N_4731,N_2857,N_3631);
xor U4732 (N_4732,N_3106,N_3281);
or U4733 (N_4733,N_3413,N_2955);
nor U4734 (N_4734,N_2939,N_2868);
or U4735 (N_4735,N_3001,N_3143);
nor U4736 (N_4736,N_3354,N_3722);
xnor U4737 (N_4737,N_2540,N_3030);
and U4738 (N_4738,N_3460,N_3228);
or U4739 (N_4739,N_3697,N_3227);
xor U4740 (N_4740,N_3191,N_3692);
nand U4741 (N_4741,N_2599,N_3043);
xnor U4742 (N_4742,N_3000,N_3542);
xor U4743 (N_4743,N_2554,N_3076);
xnor U4744 (N_4744,N_2672,N_3062);
xor U4745 (N_4745,N_3066,N_2811);
and U4746 (N_4746,N_3030,N_3472);
or U4747 (N_4747,N_3020,N_3664);
nor U4748 (N_4748,N_3472,N_2926);
and U4749 (N_4749,N_3234,N_2903);
or U4750 (N_4750,N_3462,N_3577);
xnor U4751 (N_4751,N_2543,N_2566);
nand U4752 (N_4752,N_2922,N_3256);
and U4753 (N_4753,N_3500,N_2856);
xor U4754 (N_4754,N_3747,N_3694);
or U4755 (N_4755,N_3066,N_2587);
and U4756 (N_4756,N_3692,N_3166);
or U4757 (N_4757,N_2614,N_3179);
and U4758 (N_4758,N_3613,N_3449);
or U4759 (N_4759,N_3055,N_3606);
or U4760 (N_4760,N_3473,N_2797);
nor U4761 (N_4761,N_3527,N_3194);
nor U4762 (N_4762,N_3746,N_3137);
xor U4763 (N_4763,N_3237,N_3299);
and U4764 (N_4764,N_2509,N_2888);
and U4765 (N_4765,N_3278,N_2926);
nor U4766 (N_4766,N_3507,N_3548);
nand U4767 (N_4767,N_3491,N_3202);
xnor U4768 (N_4768,N_2713,N_2919);
nand U4769 (N_4769,N_3449,N_2883);
xnor U4770 (N_4770,N_3380,N_3128);
xnor U4771 (N_4771,N_2768,N_3722);
xnor U4772 (N_4772,N_3190,N_2850);
and U4773 (N_4773,N_3507,N_2585);
or U4774 (N_4774,N_3280,N_3021);
and U4775 (N_4775,N_3408,N_3168);
xnor U4776 (N_4776,N_2578,N_2593);
or U4777 (N_4777,N_2956,N_2873);
and U4778 (N_4778,N_3118,N_2819);
or U4779 (N_4779,N_2594,N_3541);
or U4780 (N_4780,N_2977,N_3019);
and U4781 (N_4781,N_2664,N_3282);
and U4782 (N_4782,N_2568,N_2684);
xor U4783 (N_4783,N_2873,N_2895);
or U4784 (N_4784,N_3273,N_2509);
and U4785 (N_4785,N_2933,N_3594);
xnor U4786 (N_4786,N_2984,N_2971);
or U4787 (N_4787,N_2798,N_3348);
xnor U4788 (N_4788,N_2577,N_3287);
and U4789 (N_4789,N_3181,N_3056);
and U4790 (N_4790,N_3567,N_2690);
nand U4791 (N_4791,N_3081,N_3116);
nor U4792 (N_4792,N_3465,N_3350);
xnor U4793 (N_4793,N_3744,N_2993);
nand U4794 (N_4794,N_3222,N_3598);
or U4795 (N_4795,N_2677,N_3212);
xnor U4796 (N_4796,N_3361,N_3032);
or U4797 (N_4797,N_3162,N_3469);
xnor U4798 (N_4798,N_3748,N_2730);
and U4799 (N_4799,N_3398,N_2660);
or U4800 (N_4800,N_3464,N_2748);
nor U4801 (N_4801,N_2826,N_3135);
nor U4802 (N_4802,N_3473,N_2963);
and U4803 (N_4803,N_3191,N_3509);
nor U4804 (N_4804,N_2810,N_3569);
nand U4805 (N_4805,N_2721,N_3421);
and U4806 (N_4806,N_2800,N_3441);
nor U4807 (N_4807,N_3345,N_3445);
xnor U4808 (N_4808,N_3680,N_2891);
and U4809 (N_4809,N_2667,N_3458);
xnor U4810 (N_4810,N_2760,N_3261);
and U4811 (N_4811,N_3133,N_3229);
nand U4812 (N_4812,N_3430,N_2719);
xor U4813 (N_4813,N_3295,N_3275);
xor U4814 (N_4814,N_2551,N_3063);
and U4815 (N_4815,N_3554,N_2835);
nor U4816 (N_4816,N_3012,N_2683);
nor U4817 (N_4817,N_2823,N_3514);
xor U4818 (N_4818,N_3543,N_2812);
or U4819 (N_4819,N_3482,N_2678);
xnor U4820 (N_4820,N_2886,N_3436);
nor U4821 (N_4821,N_2989,N_3279);
nand U4822 (N_4822,N_2891,N_2719);
and U4823 (N_4823,N_2964,N_3012);
nor U4824 (N_4824,N_2949,N_3055);
nand U4825 (N_4825,N_2929,N_3194);
nor U4826 (N_4826,N_3270,N_3182);
or U4827 (N_4827,N_3433,N_2702);
xor U4828 (N_4828,N_3095,N_3443);
or U4829 (N_4829,N_3555,N_2780);
nand U4830 (N_4830,N_3039,N_2911);
or U4831 (N_4831,N_3738,N_3486);
and U4832 (N_4832,N_3256,N_2918);
nor U4833 (N_4833,N_2937,N_3467);
nor U4834 (N_4834,N_3426,N_3458);
xor U4835 (N_4835,N_3387,N_3188);
or U4836 (N_4836,N_3276,N_2633);
nor U4837 (N_4837,N_3227,N_2698);
xor U4838 (N_4838,N_2940,N_3726);
or U4839 (N_4839,N_2969,N_2653);
nor U4840 (N_4840,N_3496,N_3710);
xor U4841 (N_4841,N_2696,N_3515);
nand U4842 (N_4842,N_3225,N_2852);
nor U4843 (N_4843,N_2791,N_3712);
nand U4844 (N_4844,N_2523,N_3732);
nor U4845 (N_4845,N_3366,N_2885);
or U4846 (N_4846,N_3493,N_2995);
nor U4847 (N_4847,N_3348,N_3180);
nand U4848 (N_4848,N_2725,N_3255);
and U4849 (N_4849,N_3321,N_3482);
nand U4850 (N_4850,N_3357,N_2802);
xnor U4851 (N_4851,N_3080,N_3014);
or U4852 (N_4852,N_2628,N_3357);
xor U4853 (N_4853,N_3342,N_3129);
nor U4854 (N_4854,N_2798,N_2709);
and U4855 (N_4855,N_2768,N_2537);
or U4856 (N_4856,N_3248,N_2696);
and U4857 (N_4857,N_2840,N_3382);
nand U4858 (N_4858,N_3509,N_2943);
nand U4859 (N_4859,N_2880,N_3097);
and U4860 (N_4860,N_2961,N_3426);
nand U4861 (N_4861,N_2624,N_3046);
nor U4862 (N_4862,N_2500,N_3277);
nand U4863 (N_4863,N_3208,N_3399);
nand U4864 (N_4864,N_3552,N_3454);
and U4865 (N_4865,N_3401,N_3662);
and U4866 (N_4866,N_3340,N_2877);
xnor U4867 (N_4867,N_3306,N_2707);
and U4868 (N_4868,N_2974,N_3122);
or U4869 (N_4869,N_3468,N_2998);
nand U4870 (N_4870,N_2975,N_2690);
or U4871 (N_4871,N_3336,N_3581);
and U4872 (N_4872,N_3451,N_2629);
nand U4873 (N_4873,N_2519,N_3435);
nand U4874 (N_4874,N_2934,N_2865);
or U4875 (N_4875,N_2993,N_2981);
nand U4876 (N_4876,N_3279,N_2623);
nand U4877 (N_4877,N_3672,N_3247);
nor U4878 (N_4878,N_2881,N_2792);
nor U4879 (N_4879,N_3542,N_2717);
nand U4880 (N_4880,N_3227,N_2946);
or U4881 (N_4881,N_3008,N_3056);
xnor U4882 (N_4882,N_2948,N_2936);
xnor U4883 (N_4883,N_3658,N_3680);
nor U4884 (N_4884,N_2921,N_3081);
nand U4885 (N_4885,N_2884,N_3654);
nand U4886 (N_4886,N_2961,N_2654);
and U4887 (N_4887,N_2514,N_3518);
nor U4888 (N_4888,N_3265,N_2711);
xor U4889 (N_4889,N_3117,N_2744);
and U4890 (N_4890,N_3136,N_2660);
xor U4891 (N_4891,N_3443,N_3243);
or U4892 (N_4892,N_2605,N_2965);
and U4893 (N_4893,N_3518,N_3294);
and U4894 (N_4894,N_3637,N_2610);
or U4895 (N_4895,N_3172,N_3641);
nand U4896 (N_4896,N_3312,N_2815);
xor U4897 (N_4897,N_2554,N_3002);
or U4898 (N_4898,N_2892,N_3291);
and U4899 (N_4899,N_3244,N_3147);
and U4900 (N_4900,N_3562,N_2840);
xnor U4901 (N_4901,N_3212,N_3380);
and U4902 (N_4902,N_3446,N_3036);
nor U4903 (N_4903,N_3259,N_3693);
and U4904 (N_4904,N_3320,N_2805);
nand U4905 (N_4905,N_2535,N_2880);
xor U4906 (N_4906,N_3464,N_3131);
and U4907 (N_4907,N_3495,N_2543);
and U4908 (N_4908,N_3639,N_3071);
nand U4909 (N_4909,N_3556,N_3042);
nor U4910 (N_4910,N_2928,N_3619);
nor U4911 (N_4911,N_2647,N_3328);
nor U4912 (N_4912,N_2868,N_2637);
or U4913 (N_4913,N_2681,N_3658);
xnor U4914 (N_4914,N_2754,N_2559);
xnor U4915 (N_4915,N_3395,N_2707);
nor U4916 (N_4916,N_3090,N_3279);
and U4917 (N_4917,N_3705,N_3249);
xor U4918 (N_4918,N_3061,N_3322);
nand U4919 (N_4919,N_2953,N_2962);
nand U4920 (N_4920,N_2720,N_2526);
xor U4921 (N_4921,N_3548,N_2862);
nand U4922 (N_4922,N_2744,N_2913);
nor U4923 (N_4923,N_3627,N_3228);
nand U4924 (N_4924,N_3575,N_2964);
nor U4925 (N_4925,N_3599,N_3462);
nor U4926 (N_4926,N_3267,N_3517);
or U4927 (N_4927,N_3243,N_3622);
xor U4928 (N_4928,N_3617,N_2938);
or U4929 (N_4929,N_2903,N_2990);
xnor U4930 (N_4930,N_3595,N_3666);
nand U4931 (N_4931,N_2944,N_3507);
nor U4932 (N_4932,N_3021,N_3016);
or U4933 (N_4933,N_3444,N_3706);
or U4934 (N_4934,N_2956,N_3351);
and U4935 (N_4935,N_3272,N_2508);
or U4936 (N_4936,N_2913,N_2942);
and U4937 (N_4937,N_3167,N_3417);
nor U4938 (N_4938,N_3216,N_3575);
and U4939 (N_4939,N_2984,N_3224);
or U4940 (N_4940,N_3666,N_2723);
or U4941 (N_4941,N_3013,N_3218);
and U4942 (N_4942,N_3627,N_3258);
nor U4943 (N_4943,N_3226,N_2578);
nand U4944 (N_4944,N_3489,N_2878);
xnor U4945 (N_4945,N_2765,N_3486);
or U4946 (N_4946,N_2839,N_2854);
or U4947 (N_4947,N_3018,N_3446);
nor U4948 (N_4948,N_2964,N_2625);
nor U4949 (N_4949,N_3629,N_2978);
xnor U4950 (N_4950,N_3438,N_2919);
nand U4951 (N_4951,N_2604,N_2819);
xnor U4952 (N_4952,N_2704,N_3314);
or U4953 (N_4953,N_2646,N_2542);
nand U4954 (N_4954,N_3643,N_3437);
nand U4955 (N_4955,N_3229,N_3264);
and U4956 (N_4956,N_2932,N_3321);
nor U4957 (N_4957,N_3641,N_3703);
nand U4958 (N_4958,N_3445,N_3087);
nor U4959 (N_4959,N_3535,N_3725);
xor U4960 (N_4960,N_2570,N_3551);
nor U4961 (N_4961,N_2847,N_2502);
or U4962 (N_4962,N_2663,N_3143);
or U4963 (N_4963,N_3331,N_3046);
xor U4964 (N_4964,N_3293,N_2837);
nand U4965 (N_4965,N_3500,N_3538);
and U4966 (N_4966,N_3692,N_3064);
and U4967 (N_4967,N_2568,N_3161);
or U4968 (N_4968,N_3495,N_2871);
nor U4969 (N_4969,N_3339,N_3169);
xnor U4970 (N_4970,N_2829,N_3597);
or U4971 (N_4971,N_2803,N_2519);
or U4972 (N_4972,N_3021,N_3050);
xnor U4973 (N_4973,N_3567,N_2878);
nor U4974 (N_4974,N_3290,N_3198);
nand U4975 (N_4975,N_3553,N_3224);
and U4976 (N_4976,N_3470,N_3012);
or U4977 (N_4977,N_2659,N_3311);
and U4978 (N_4978,N_2687,N_2940);
xor U4979 (N_4979,N_3511,N_3593);
nand U4980 (N_4980,N_3297,N_3154);
nor U4981 (N_4981,N_2634,N_3645);
nand U4982 (N_4982,N_3328,N_3057);
or U4983 (N_4983,N_3526,N_3621);
xnor U4984 (N_4984,N_3412,N_3433);
xor U4985 (N_4985,N_3745,N_3348);
nor U4986 (N_4986,N_2841,N_3002);
nor U4987 (N_4987,N_3234,N_3365);
and U4988 (N_4988,N_3427,N_2698);
nor U4989 (N_4989,N_2510,N_3675);
and U4990 (N_4990,N_2648,N_2692);
nand U4991 (N_4991,N_3420,N_3227);
nand U4992 (N_4992,N_3502,N_3108);
xor U4993 (N_4993,N_3236,N_3693);
xor U4994 (N_4994,N_3006,N_3705);
nand U4995 (N_4995,N_3555,N_3425);
or U4996 (N_4996,N_2517,N_3018);
nor U4997 (N_4997,N_3587,N_2795);
xnor U4998 (N_4998,N_2513,N_3216);
or U4999 (N_4999,N_3054,N_2527);
or U5000 (N_5000,N_4139,N_4157);
nor U5001 (N_5001,N_4553,N_4035);
nor U5002 (N_5002,N_4839,N_4833);
nor U5003 (N_5003,N_4115,N_4718);
xor U5004 (N_5004,N_4779,N_4905);
and U5005 (N_5005,N_4025,N_4235);
and U5006 (N_5006,N_4254,N_4770);
or U5007 (N_5007,N_4564,N_4902);
and U5008 (N_5008,N_3971,N_4217);
xor U5009 (N_5009,N_4927,N_4335);
nand U5010 (N_5010,N_4530,N_4596);
nor U5011 (N_5011,N_4194,N_4636);
xnor U5012 (N_5012,N_3907,N_4768);
nor U5013 (N_5013,N_4411,N_4037);
nor U5014 (N_5014,N_4331,N_4527);
nor U5015 (N_5015,N_4844,N_4130);
or U5016 (N_5016,N_4283,N_3908);
xor U5017 (N_5017,N_4608,N_4952);
and U5018 (N_5018,N_3989,N_4987);
and U5019 (N_5019,N_4716,N_4074);
and U5020 (N_5020,N_4118,N_4357);
nand U5021 (N_5021,N_3833,N_4903);
xor U5022 (N_5022,N_4236,N_3934);
or U5023 (N_5023,N_3816,N_4670);
xor U5024 (N_5024,N_4843,N_4188);
or U5025 (N_5025,N_4699,N_4231);
nand U5026 (N_5026,N_4134,N_4268);
nor U5027 (N_5027,N_3813,N_4717);
nand U5028 (N_5028,N_4323,N_4767);
nor U5029 (N_5029,N_3964,N_4394);
nand U5030 (N_5030,N_4375,N_4016);
nor U5031 (N_5031,N_4280,N_3766);
or U5032 (N_5032,N_4090,N_4885);
nand U5033 (N_5033,N_4145,N_4834);
nor U5034 (N_5034,N_3928,N_3829);
nor U5035 (N_5035,N_3924,N_4351);
nand U5036 (N_5036,N_4733,N_4295);
xnor U5037 (N_5037,N_4956,N_4909);
and U5038 (N_5038,N_3945,N_4935);
nor U5039 (N_5039,N_4931,N_4749);
nand U5040 (N_5040,N_4001,N_4206);
or U5041 (N_5041,N_4598,N_4058);
nor U5042 (N_5042,N_3815,N_4079);
and U5043 (N_5043,N_3985,N_4817);
nand U5044 (N_5044,N_4831,N_4920);
xor U5045 (N_5045,N_4528,N_3846);
or U5046 (N_5046,N_3970,N_4019);
and U5047 (N_5047,N_4874,N_4406);
xor U5048 (N_5048,N_3903,N_4476);
and U5049 (N_5049,N_4451,N_4635);
and U5050 (N_5050,N_4329,N_4904);
or U5051 (N_5051,N_4128,N_4786);
and U5052 (N_5052,N_4223,N_4612);
nand U5053 (N_5053,N_4899,N_4923);
xnor U5054 (N_5054,N_4341,N_4032);
nand U5055 (N_5055,N_4298,N_3942);
nand U5056 (N_5056,N_4447,N_3892);
xor U5057 (N_5057,N_3859,N_4325);
or U5058 (N_5058,N_3993,N_4809);
nor U5059 (N_5059,N_4604,N_4473);
or U5060 (N_5060,N_4121,N_4264);
xor U5061 (N_5061,N_4477,N_4429);
and U5062 (N_5062,N_4321,N_4694);
nor U5063 (N_5063,N_4054,N_4419);
nand U5064 (N_5064,N_3952,N_4934);
or U5065 (N_5065,N_4728,N_4173);
xor U5066 (N_5066,N_4137,N_3818);
nor U5067 (N_5067,N_4774,N_4017);
nor U5068 (N_5068,N_4590,N_4291);
xnor U5069 (N_5069,N_3967,N_4972);
and U5070 (N_5070,N_4083,N_4624);
or U5071 (N_5071,N_4010,N_4637);
xnor U5072 (N_5072,N_4092,N_4089);
nand U5073 (N_5073,N_4234,N_4305);
nor U5074 (N_5074,N_4229,N_4174);
xor U5075 (N_5075,N_4866,N_3905);
and U5076 (N_5076,N_3780,N_4542);
xnor U5077 (N_5077,N_4474,N_4479);
and U5078 (N_5078,N_3773,N_3946);
xor U5079 (N_5079,N_3764,N_4973);
or U5080 (N_5080,N_4286,N_4353);
nor U5081 (N_5081,N_4125,N_4883);
nand U5082 (N_5082,N_3869,N_4135);
or U5083 (N_5083,N_4066,N_3873);
nor U5084 (N_5084,N_4342,N_3792);
nor U5085 (N_5085,N_4413,N_4896);
or U5086 (N_5086,N_4237,N_4819);
xnor U5087 (N_5087,N_4519,N_4020);
or U5088 (N_5088,N_4114,N_4712);
xnor U5089 (N_5089,N_4098,N_3936);
and U5090 (N_5090,N_4856,N_3986);
or U5091 (N_5091,N_4187,N_4769);
xor U5092 (N_5092,N_4766,N_4213);
and U5093 (N_5093,N_4751,N_4205);
or U5094 (N_5094,N_4415,N_4502);
or U5095 (N_5095,N_4651,N_4064);
or U5096 (N_5096,N_4991,N_4913);
nor U5097 (N_5097,N_4799,N_4685);
and U5098 (N_5098,N_4348,N_3949);
nand U5099 (N_5099,N_4386,N_4803);
nand U5100 (N_5100,N_4053,N_4155);
nor U5101 (N_5101,N_4172,N_4049);
and U5102 (N_5102,N_3870,N_4080);
or U5103 (N_5103,N_4452,N_4330);
nor U5104 (N_5104,N_3817,N_4928);
nand U5105 (N_5105,N_4692,N_3864);
nor U5106 (N_5106,N_4729,N_4674);
xor U5107 (N_5107,N_3927,N_4271);
nand U5108 (N_5108,N_4561,N_3957);
xnor U5109 (N_5109,N_4820,N_4185);
and U5110 (N_5110,N_4050,N_3983);
nor U5111 (N_5111,N_4701,N_4791);
or U5112 (N_5112,N_4028,N_4269);
nor U5113 (N_5113,N_3785,N_4732);
xor U5114 (N_5114,N_3787,N_4849);
or U5115 (N_5115,N_4320,N_3923);
xnor U5116 (N_5116,N_3809,N_4738);
nand U5117 (N_5117,N_4591,N_4499);
nor U5118 (N_5118,N_3755,N_4850);
nor U5119 (N_5119,N_3863,N_4152);
and U5120 (N_5120,N_4589,N_3968);
xor U5121 (N_5121,N_4789,N_4613);
xnor U5122 (N_5122,N_4181,N_4731);
xor U5123 (N_5123,N_4878,N_4763);
and U5124 (N_5124,N_4140,N_3757);
xnor U5125 (N_5125,N_4365,N_4262);
nand U5126 (N_5126,N_4493,N_4508);
xnor U5127 (N_5127,N_4463,N_4420);
nor U5128 (N_5128,N_4042,N_4541);
nand U5129 (N_5129,N_4397,N_4946);
or U5130 (N_5130,N_4912,N_4698);
or U5131 (N_5131,N_4399,N_3839);
nor U5132 (N_5132,N_4143,N_4714);
xor U5133 (N_5133,N_4450,N_4123);
and U5134 (N_5134,N_4607,N_4443);
nor U5135 (N_5135,N_3978,N_3888);
nor U5136 (N_5136,N_3834,N_4785);
and U5137 (N_5137,N_4200,N_4540);
nand U5138 (N_5138,N_4290,N_4507);
xor U5139 (N_5139,N_4706,N_3838);
and U5140 (N_5140,N_4018,N_3950);
xnor U5141 (N_5141,N_4802,N_4629);
or U5142 (N_5142,N_4610,N_4232);
or U5143 (N_5143,N_4576,N_4981);
xor U5144 (N_5144,N_4556,N_4898);
nand U5145 (N_5145,N_4322,N_4689);
and U5146 (N_5146,N_4457,N_3944);
xnor U5147 (N_5147,N_4518,N_4369);
nor U5148 (N_5148,N_4796,N_4183);
xor U5149 (N_5149,N_4841,N_3808);
or U5150 (N_5150,N_4675,N_4317);
nor U5151 (N_5151,N_4076,N_4256);
xnor U5152 (N_5152,N_3917,N_4772);
nand U5153 (N_5153,N_4566,N_3904);
nand U5154 (N_5154,N_4681,N_4277);
or U5155 (N_5155,N_4857,N_4086);
xnor U5156 (N_5156,N_4600,N_4823);
and U5157 (N_5157,N_4593,N_4897);
nand U5158 (N_5158,N_4884,N_3868);
or U5159 (N_5159,N_4512,N_4273);
and U5160 (N_5160,N_4662,N_4537);
nand U5161 (N_5161,N_4436,N_4797);
and U5162 (N_5162,N_3973,N_4975);
nand U5163 (N_5163,N_3932,N_4836);
and U5164 (N_5164,N_4208,N_4124);
or U5165 (N_5165,N_4555,N_4551);
nand U5166 (N_5166,N_4788,N_4778);
nor U5167 (N_5167,N_3754,N_4279);
nand U5168 (N_5168,N_4690,N_4048);
or U5169 (N_5169,N_4241,N_4951);
or U5170 (N_5170,N_4852,N_4379);
nand U5171 (N_5171,N_4739,N_3775);
xor U5172 (N_5172,N_4129,N_4459);
nor U5173 (N_5173,N_4059,N_4549);
nor U5174 (N_5174,N_3961,N_3980);
or U5175 (N_5175,N_4112,N_3913);
xnor U5176 (N_5176,N_4558,N_4201);
and U5177 (N_5177,N_3806,N_3953);
and U5178 (N_5178,N_4361,N_4759);
nor U5179 (N_5179,N_4614,N_4167);
nor U5180 (N_5180,N_3895,N_3777);
nor U5181 (N_5181,N_4940,N_4942);
and U5182 (N_5182,N_4830,N_4484);
xnor U5183 (N_5183,N_4248,N_4171);
or U5184 (N_5184,N_4434,N_4146);
xor U5185 (N_5185,N_4683,N_4122);
nor U5186 (N_5186,N_4383,N_4068);
xor U5187 (N_5187,N_4777,N_4472);
nor U5188 (N_5188,N_4319,N_4220);
and U5189 (N_5189,N_4426,N_3914);
xnor U5190 (N_5190,N_4469,N_4166);
xnor U5191 (N_5191,N_4390,N_4891);
xor U5192 (N_5192,N_4937,N_4713);
or U5193 (N_5193,N_4498,N_4314);
nor U5194 (N_5194,N_3879,N_4643);
or U5195 (N_5195,N_3848,N_3836);
and U5196 (N_5196,N_3795,N_4676);
nor U5197 (N_5197,N_4204,N_4022);
nand U5198 (N_5198,N_3992,N_4798);
nor U5199 (N_5199,N_4743,N_4030);
xnor U5200 (N_5200,N_3772,N_4582);
and U5201 (N_5201,N_3872,N_3759);
nand U5202 (N_5202,N_4156,N_3982);
or U5203 (N_5203,N_4615,N_4040);
nor U5204 (N_5204,N_4193,N_4218);
and U5205 (N_5205,N_4545,N_4299);
nand U5206 (N_5206,N_4827,N_4816);
and U5207 (N_5207,N_4832,N_4210);
or U5208 (N_5208,N_4585,N_4116);
nand U5209 (N_5209,N_4529,N_4918);
nand U5210 (N_5210,N_4992,N_4966);
xor U5211 (N_5211,N_4103,N_4313);
xnor U5212 (N_5212,N_4380,N_4368);
nor U5213 (N_5213,N_4707,N_4359);
and U5214 (N_5214,N_4258,N_4765);
or U5215 (N_5215,N_3793,N_3969);
or U5216 (N_5216,N_3857,N_3844);
xnor U5217 (N_5217,N_3786,N_4881);
or U5218 (N_5218,N_4251,N_3984);
nor U5219 (N_5219,N_4072,N_4691);
and U5220 (N_5220,N_4861,N_3791);
nand U5221 (N_5221,N_4672,N_4845);
and U5222 (N_5222,N_4136,N_4730);
xor U5223 (N_5223,N_4259,N_4976);
nand U5224 (N_5224,N_3954,N_4239);
or U5225 (N_5225,N_4316,N_4737);
xnor U5226 (N_5226,N_4653,N_3991);
xor U5227 (N_5227,N_4747,N_4742);
and U5228 (N_5228,N_4289,N_3830);
or U5229 (N_5229,N_4671,N_4606);
xnor U5230 (N_5230,N_4658,N_4538);
nand U5231 (N_5231,N_4075,N_4828);
or U5232 (N_5232,N_3893,N_4750);
or U5233 (N_5233,N_4969,N_4071);
nand U5234 (N_5234,N_3899,N_4013);
and U5235 (N_5235,N_4366,N_4374);
xnor U5236 (N_5236,N_3918,N_4175);
or U5237 (N_5237,N_4052,N_4811);
nand U5238 (N_5238,N_4177,N_4449);
nand U5239 (N_5239,N_4400,N_3958);
nor U5240 (N_5240,N_4311,N_4597);
and U5241 (N_5241,N_3751,N_3959);
or U5242 (N_5242,N_3956,N_4872);
nand U5243 (N_5243,N_3854,N_4933);
nor U5244 (N_5244,N_4352,N_4997);
nand U5245 (N_5245,N_4853,N_4044);
nor U5246 (N_5246,N_4611,N_4882);
xnor U5247 (N_5247,N_4900,N_4428);
nor U5248 (N_5248,N_4097,N_4081);
nor U5249 (N_5249,N_4702,N_3894);
xnor U5250 (N_5250,N_4875,N_3827);
nand U5251 (N_5251,N_3776,N_4734);
nor U5252 (N_5252,N_4483,N_3768);
and U5253 (N_5253,N_4043,N_4078);
nand U5254 (N_5254,N_4389,N_4332);
nor U5255 (N_5255,N_4027,N_4412);
and U5256 (N_5256,N_4002,N_4441);
and U5257 (N_5257,N_4801,N_4526);
nor U5258 (N_5258,N_3832,N_4535);
and U5259 (N_5259,N_3831,N_4021);
or U5260 (N_5260,N_3856,N_4800);
nand U5261 (N_5261,N_4253,N_4646);
xor U5262 (N_5262,N_3963,N_3911);
nor U5263 (N_5263,N_4039,N_4107);
nand U5264 (N_5264,N_4740,N_3814);
nor U5265 (N_5265,N_3765,N_4632);
nor U5266 (N_5266,N_4270,N_4127);
and U5267 (N_5267,N_4186,N_3998);
or U5268 (N_5268,N_4993,N_4189);
nand U5269 (N_5269,N_4260,N_4854);
xor U5270 (N_5270,N_4961,N_4063);
or U5271 (N_5271,N_3988,N_4805);
xor U5272 (N_5272,N_4669,N_4794);
and U5273 (N_5273,N_4810,N_3783);
nand U5274 (N_5274,N_4625,N_4423);
nor U5275 (N_5275,N_3925,N_4744);
and U5276 (N_5276,N_4522,N_4915);
xor U5277 (N_5277,N_4466,N_4509);
and U5278 (N_5278,N_3851,N_4087);
and U5279 (N_5279,N_3979,N_4641);
nand U5280 (N_5280,N_4438,N_3821);
and U5281 (N_5281,N_3767,N_4243);
or U5282 (N_5282,N_4906,N_4384);
or U5283 (N_5283,N_4131,N_4191);
and U5284 (N_5284,N_3760,N_4648);
or U5285 (N_5285,N_4574,N_4267);
nand U5286 (N_5286,N_4524,N_4471);
nor U5287 (N_5287,N_4084,N_4639);
nor U5288 (N_5288,N_4096,N_4288);
or U5289 (N_5289,N_4695,N_3850);
or U5290 (N_5290,N_4859,N_3941);
nand U5291 (N_5291,N_3805,N_4947);
or U5292 (N_5292,N_4132,N_4936);
and U5293 (N_5293,N_3915,N_3812);
nor U5294 (N_5294,N_4650,N_4403);
xnor U5295 (N_5295,N_4982,N_3782);
and U5296 (N_5296,N_4445,N_4988);
or U5297 (N_5297,N_4886,N_3883);
and U5298 (N_5298,N_4062,N_4228);
and U5299 (N_5299,N_4148,N_4184);
and U5300 (N_5300,N_4111,N_4974);
and U5301 (N_5301,N_3779,N_3855);
and U5302 (N_5302,N_4968,N_4977);
nor U5303 (N_5303,N_4462,N_4978);
or U5304 (N_5304,N_4346,N_4003);
nor U5305 (N_5305,N_4948,N_4563);
xnor U5306 (N_5306,N_3976,N_4657);
nand U5307 (N_5307,N_3865,N_4162);
nor U5308 (N_5308,N_4515,N_3898);
nor U5309 (N_5309,N_4696,N_4679);
nand U5310 (N_5310,N_4113,N_3940);
xnor U5311 (N_5311,N_4494,N_4647);
nand U5312 (N_5312,N_3930,N_4603);
xnor U5313 (N_5313,N_3916,N_4531);
xor U5314 (N_5314,N_3889,N_4281);
nand U5315 (N_5315,N_3900,N_4318);
and U5316 (N_5316,N_4703,N_4395);
nand U5317 (N_5317,N_3943,N_4340);
or U5318 (N_5318,N_4754,N_4285);
nand U5319 (N_5319,N_4626,N_4385);
nand U5320 (N_5320,N_4682,N_4726);
xnor U5321 (N_5321,N_3921,N_4761);
nand U5322 (N_5322,N_3987,N_4783);
nor U5323 (N_5323,N_4544,N_4024);
nor U5324 (N_5324,N_3802,N_4454);
xnor U5325 (N_5325,N_4921,N_4619);
nor U5326 (N_5326,N_4012,N_4294);
nand U5327 (N_5327,N_3866,N_3790);
or U5328 (N_5328,N_4709,N_4552);
or U5329 (N_5329,N_4150,N_4245);
nand U5330 (N_5330,N_4496,N_4922);
nor U5331 (N_5331,N_4572,N_4301);
or U5332 (N_5332,N_4873,N_4202);
nand U5333 (N_5333,N_4547,N_4067);
xnor U5334 (N_5334,N_4869,N_4414);
or U5335 (N_5335,N_4645,N_3796);
and U5336 (N_5336,N_4879,N_4980);
nand U5337 (N_5337,N_3871,N_4757);
nand U5338 (N_5338,N_4034,N_3887);
nand U5339 (N_5339,N_3794,N_3860);
nor U5340 (N_5340,N_3753,N_4578);
or U5341 (N_5341,N_3828,N_3845);
nand U5342 (N_5342,N_4337,N_4154);
xor U5343 (N_5343,N_4338,N_4465);
xor U5344 (N_5344,N_4656,N_3804);
or U5345 (N_5345,N_3789,N_3882);
xnor U5346 (N_5346,N_4310,N_3841);
and U5347 (N_5347,N_4138,N_4168);
and U5348 (N_5348,N_4848,N_4093);
or U5349 (N_5349,N_4704,N_4176);
or U5350 (N_5350,N_4345,N_4865);
nand U5351 (N_5351,N_4995,N_4160);
or U5352 (N_5352,N_4424,N_4986);
or U5353 (N_5353,N_4492,N_4257);
and U5354 (N_5354,N_4554,N_4312);
nand U5355 (N_5355,N_3819,N_4388);
or U5356 (N_5356,N_4930,N_4655);
and U5357 (N_5357,N_4667,N_4370);
or U5358 (N_5358,N_4282,N_4482);
and U5359 (N_5359,N_4488,N_4938);
and U5360 (N_5360,N_4687,N_4300);
nand U5361 (N_5361,N_4278,N_4047);
and U5362 (N_5362,N_4272,N_4199);
and U5363 (N_5363,N_4328,N_4350);
nor U5364 (N_5364,N_4023,N_4815);
nor U5365 (N_5365,N_4391,N_4943);
nor U5366 (N_5366,N_4621,N_4161);
and U5367 (N_5367,N_4967,N_4808);
nor U5368 (N_5368,N_4315,N_4534);
xnor U5369 (N_5369,N_4514,N_4179);
and U5370 (N_5370,N_4456,N_4439);
and U5371 (N_5371,N_3877,N_3807);
xnor U5372 (N_5372,N_4005,N_4159);
xor U5373 (N_5373,N_3843,N_4577);
nor U5374 (N_5374,N_4249,N_4654);
nand U5375 (N_5375,N_4077,N_4082);
or U5376 (N_5376,N_3762,N_4617);
or U5377 (N_5377,N_4782,N_4421);
nor U5378 (N_5378,N_4941,N_4233);
and U5379 (N_5379,N_3750,N_4334);
and U5380 (N_5380,N_3852,N_3974);
nand U5381 (N_5381,N_4065,N_3912);
xnor U5382 (N_5382,N_3853,N_4813);
and U5383 (N_5383,N_4000,N_4944);
nor U5384 (N_5384,N_4602,N_4356);
and U5385 (N_5385,N_4649,N_4627);
nand U5386 (N_5386,N_4026,N_4180);
or U5387 (N_5387,N_3822,N_4999);
nand U5388 (N_5388,N_4432,N_4601);
or U5389 (N_5389,N_4567,N_4503);
nand U5390 (N_5390,N_3896,N_4746);
nor U5391 (N_5391,N_4634,N_4101);
and U5392 (N_5392,N_3799,N_4762);
nor U5393 (N_5393,N_4680,N_4787);
xor U5394 (N_5394,N_3797,N_4387);
xor U5395 (N_5395,N_4971,N_4640);
xor U5396 (N_5396,N_3960,N_4868);
and U5397 (N_5397,N_4196,N_4818);
xnor U5398 (N_5398,N_4036,N_4207);
nand U5399 (N_5399,N_4442,N_4246);
nor U5400 (N_5400,N_4446,N_4994);
or U5401 (N_5401,N_4398,N_4141);
or U5402 (N_5402,N_4957,N_4425);
or U5403 (N_5403,N_4736,N_4829);
nand U5404 (N_5404,N_4893,N_4876);
or U5405 (N_5405,N_4989,N_4573);
or U5406 (N_5406,N_4410,N_3897);
or U5407 (N_5407,N_3966,N_4665);
xnor U5408 (N_5408,N_4758,N_4106);
and U5409 (N_5409,N_4008,N_4668);
xnor U5410 (N_5410,N_3774,N_4894);
or U5411 (N_5411,N_4812,N_4142);
nor U5412 (N_5412,N_4911,N_3922);
or U5413 (N_5413,N_3981,N_4720);
xnor U5414 (N_5414,N_4569,N_3965);
and U5415 (N_5415,N_3996,N_4919);
and U5416 (N_5416,N_4756,N_3935);
and U5417 (N_5417,N_4609,N_4073);
and U5418 (N_5418,N_4336,N_4453);
or U5419 (N_5419,N_4170,N_4725);
and U5420 (N_5420,N_3826,N_4265);
xor U5421 (N_5421,N_4292,N_4532);
nor U5422 (N_5422,N_4851,N_3752);
xor U5423 (N_5423,N_4673,N_4409);
nand U5424 (N_5424,N_3990,N_4748);
and U5425 (N_5425,N_3919,N_3840);
nor U5426 (N_5426,N_4784,N_4838);
nor U5427 (N_5427,N_4924,N_4562);
nor U5428 (N_5428,N_4623,N_4373);
xnor U5429 (N_5429,N_3798,N_4307);
nor U5430 (N_5430,N_4437,N_3837);
nand U5431 (N_5431,N_3769,N_4684);
or U5432 (N_5432,N_4580,N_4495);
nand U5433 (N_5433,N_4009,N_4983);
xor U5434 (N_5434,N_4060,N_4806);
or U5435 (N_5435,N_3929,N_4252);
nand U5436 (N_5436,N_4287,N_4950);
nand U5437 (N_5437,N_4929,N_4195);
nor U5438 (N_5438,N_4500,N_4458);
xor U5439 (N_5439,N_4901,N_4304);
nor U5440 (N_5440,N_4644,N_4945);
and U5441 (N_5441,N_4723,N_4004);
nand U5442 (N_5442,N_4460,N_3995);
nand U5443 (N_5443,N_3875,N_4085);
nor U5444 (N_5444,N_4362,N_3962);
xor U5445 (N_5445,N_4990,N_4333);
or U5446 (N_5446,N_4088,N_3781);
or U5447 (N_5447,N_4431,N_4792);
xnor U5448 (N_5448,N_4100,N_3886);
nor U5449 (N_5449,N_4405,N_4543);
xnor U5450 (N_5450,N_4825,N_4605);
or U5451 (N_5451,N_4953,N_4440);
and U5452 (N_5452,N_4877,N_4917);
xor U5453 (N_5453,N_4954,N_4014);
nand U5454 (N_5454,N_4343,N_4722);
or U5455 (N_5455,N_3876,N_4306);
and U5456 (N_5456,N_4594,N_3867);
xnor U5457 (N_5457,N_4029,N_3803);
nor U5458 (N_5458,N_3948,N_4302);
and U5459 (N_5459,N_3947,N_4192);
nand U5460 (N_5460,N_4491,N_4710);
and U5461 (N_5461,N_4964,N_4427);
nor U5462 (N_5462,N_4327,N_4771);
or U5463 (N_5463,N_4045,N_4163);
nand U5464 (N_5464,N_3820,N_4513);
xnor U5465 (N_5465,N_4571,N_4536);
nor U5466 (N_5466,N_4996,N_4117);
xnor U5467 (N_5467,N_3881,N_4664);
and U5468 (N_5468,N_3909,N_3824);
and U5469 (N_5469,N_4517,N_4764);
xor U5470 (N_5470,N_4046,N_4178);
and U5471 (N_5471,N_4686,N_3771);
xor U5472 (N_5472,N_4659,N_4926);
nor U5473 (N_5473,N_4102,N_4408);
nor U5474 (N_5474,N_4363,N_3977);
nand U5475 (N_5475,N_4211,N_4261);
and U5476 (N_5476,N_3931,N_4266);
xnor U5477 (N_5477,N_4925,N_3885);
xnor U5478 (N_5478,N_3939,N_4401);
xnor U5479 (N_5479,N_4914,N_3938);
or U5480 (N_5480,N_4416,N_4888);
and U5481 (N_5481,N_4480,N_4055);
or U5482 (N_5482,N_4381,N_4678);
nand U5483 (N_5483,N_4033,N_4119);
nor U5484 (N_5484,N_4583,N_4633);
and U5485 (N_5485,N_4599,N_4895);
and U5486 (N_5486,N_3847,N_4349);
xor U5487 (N_5487,N_4247,N_4781);
nand U5488 (N_5488,N_4505,N_3862);
nor U5489 (N_5489,N_4377,N_4727);
xor U5490 (N_5490,N_4430,N_4435);
nor U5491 (N_5491,N_4753,N_4516);
xnor U5492 (N_5492,N_4255,N_4705);
nand U5493 (N_5493,N_4916,N_4308);
and U5494 (N_5494,N_3951,N_4151);
and U5495 (N_5495,N_4070,N_4225);
or U5496 (N_5496,N_4560,N_3849);
and U5497 (N_5497,N_4095,N_4104);
xnor U5498 (N_5498,N_4949,N_4011);
xor U5499 (N_5499,N_3972,N_4015);
xor U5500 (N_5500,N_4226,N_4826);
nor U5501 (N_5501,N_4109,N_3884);
nand U5502 (N_5502,N_4481,N_4504);
nand U5503 (N_5503,N_4099,N_4979);
or U5504 (N_5504,N_4219,N_4837);
nor U5505 (N_5505,N_4570,N_4700);
nand U5506 (N_5506,N_3778,N_4889);
xnor U5507 (N_5507,N_4557,N_4711);
nor U5508 (N_5508,N_4719,N_3901);
and U5509 (N_5509,N_4932,N_4371);
nor U5510 (N_5510,N_3801,N_4110);
and U5511 (N_5511,N_4618,N_4203);
nor U5512 (N_5512,N_4263,N_4497);
xor U5513 (N_5513,N_4584,N_4959);
or U5514 (N_5514,N_4182,N_3810);
nand U5515 (N_5515,N_4840,N_4984);
or U5516 (N_5516,N_4297,N_4422);
and U5517 (N_5517,N_4858,N_4870);
and U5518 (N_5518,N_3994,N_3920);
nand U5519 (N_5519,N_4326,N_4120);
nand U5520 (N_5520,N_4907,N_4688);
and U5521 (N_5521,N_3784,N_4715);
or U5522 (N_5522,N_4533,N_4795);
or U5523 (N_5523,N_3861,N_4244);
nor U5524 (N_5524,N_3758,N_4478);
nand U5525 (N_5525,N_4444,N_4007);
or U5526 (N_5526,N_4216,N_4847);
or U5527 (N_5527,N_4775,N_4470);
nand U5528 (N_5528,N_4224,N_4487);
xnor U5529 (N_5529,N_4586,N_4910);
nor U5530 (N_5530,N_3756,N_4565);
xor U5531 (N_5531,N_4871,N_4324);
nor U5532 (N_5532,N_4250,N_4721);
and U5533 (N_5533,N_3880,N_4814);
and U5534 (N_5534,N_4393,N_4344);
nand U5535 (N_5535,N_4867,N_3763);
nor U5536 (N_5536,N_4568,N_4455);
nor U5537 (N_5537,N_4461,N_3878);
nor U5538 (N_5538,N_4660,N_4741);
or U5539 (N_5539,N_4041,N_4892);
nor U5540 (N_5540,N_4275,N_3823);
and U5541 (N_5541,N_4616,N_4031);
xor U5542 (N_5542,N_4539,N_4677);
or U5543 (N_5543,N_4367,N_4880);
or U5544 (N_5544,N_4396,N_4939);
xnor U5545 (N_5545,N_4051,N_4965);
nand U5546 (N_5546,N_4970,N_4793);
and U5547 (N_5547,N_4392,N_4887);
or U5548 (N_5548,N_4227,N_4355);
xor U5549 (N_5549,N_4588,N_4622);
or U5550 (N_5550,N_4222,N_3835);
or U5551 (N_5551,N_4376,N_3890);
nor U5552 (N_5552,N_4276,N_4056);
xnor U5553 (N_5553,N_3800,N_4382);
nor U5554 (N_5554,N_4506,N_4165);
nor U5555 (N_5555,N_4790,N_3858);
or U5556 (N_5556,N_4642,N_4581);
or U5557 (N_5557,N_4133,N_4548);
and U5558 (N_5558,N_4960,N_4293);
or U5559 (N_5559,N_4467,N_4807);
xor U5560 (N_5560,N_4697,N_4418);
nand U5561 (N_5561,N_4842,N_4475);
and U5562 (N_5562,N_4169,N_4628);
and U5563 (N_5563,N_4863,N_4105);
or U5564 (N_5564,N_4525,N_4755);
xnor U5565 (N_5565,N_4347,N_4198);
xor U5566 (N_5566,N_4860,N_4240);
or U5567 (N_5567,N_4214,N_4862);
nor U5568 (N_5568,N_4372,N_4587);
and U5569 (N_5569,N_4069,N_3770);
and U5570 (N_5570,N_4490,N_4575);
nor U5571 (N_5571,N_4520,N_3926);
or U5572 (N_5572,N_4864,N_4631);
nor U5573 (N_5573,N_4404,N_4358);
and U5574 (N_5574,N_4510,N_3902);
nand U5575 (N_5575,N_4804,N_3955);
or U5576 (N_5576,N_4284,N_4559);
nand U5577 (N_5577,N_4061,N_4745);
nor U5578 (N_5578,N_4407,N_4364);
or U5579 (N_5579,N_4652,N_4057);
or U5580 (N_5580,N_3891,N_3788);
or U5581 (N_5581,N_4855,N_4780);
nand U5582 (N_5582,N_3975,N_4164);
and U5583 (N_5583,N_4230,N_4448);
and U5584 (N_5584,N_4666,N_4752);
nor U5585 (N_5585,N_4821,N_4661);
and U5586 (N_5586,N_4890,N_4038);
xnor U5587 (N_5587,N_4592,N_4760);
and U5588 (N_5588,N_4091,N_3999);
xnor U5589 (N_5589,N_3825,N_4360);
or U5590 (N_5590,N_4663,N_4094);
or U5591 (N_5591,N_4776,N_4190);
xnor U5592 (N_5592,N_4501,N_4724);
nor U5593 (N_5593,N_4595,N_4242);
nand U5594 (N_5594,N_4309,N_4417);
nor U5595 (N_5595,N_4153,N_4523);
nand U5596 (N_5596,N_4486,N_4464);
xnor U5597 (N_5597,N_3997,N_4521);
and U5598 (N_5598,N_4638,N_4908);
nand U5599 (N_5599,N_4489,N_4354);
nor U5600 (N_5600,N_3842,N_4221);
or U5601 (N_5601,N_3761,N_4735);
nor U5602 (N_5602,N_4824,N_4998);
nand U5603 (N_5603,N_4579,N_4693);
nand U5604 (N_5604,N_4215,N_4846);
nor U5605 (N_5605,N_4303,N_4274);
nor U5606 (N_5606,N_4238,N_4822);
nor U5607 (N_5607,N_4402,N_4773);
or U5608 (N_5608,N_3937,N_4468);
and U5609 (N_5609,N_4835,N_4378);
or U5610 (N_5610,N_3874,N_3811);
nor U5611 (N_5611,N_4296,N_4546);
xnor U5612 (N_5612,N_4485,N_4962);
nor U5613 (N_5613,N_4108,N_4147);
xnor U5614 (N_5614,N_4126,N_4708);
xnor U5615 (N_5615,N_4212,N_4955);
or U5616 (N_5616,N_4630,N_4144);
nand U5617 (N_5617,N_4985,N_4511);
nor U5618 (N_5618,N_4149,N_4620);
and U5619 (N_5619,N_4963,N_4006);
or U5620 (N_5620,N_3910,N_4433);
nor U5621 (N_5621,N_4209,N_4197);
and U5622 (N_5622,N_4958,N_4339);
or U5623 (N_5623,N_3933,N_4158);
and U5624 (N_5624,N_3906,N_4550);
or U5625 (N_5625,N_3805,N_4270);
or U5626 (N_5626,N_4427,N_4718);
xor U5627 (N_5627,N_4433,N_4557);
nor U5628 (N_5628,N_4312,N_4547);
or U5629 (N_5629,N_4558,N_4163);
xnor U5630 (N_5630,N_4526,N_4315);
xnor U5631 (N_5631,N_4419,N_4629);
xnor U5632 (N_5632,N_4868,N_4050);
and U5633 (N_5633,N_4556,N_4652);
or U5634 (N_5634,N_4148,N_4303);
or U5635 (N_5635,N_3900,N_4776);
nand U5636 (N_5636,N_4620,N_3976);
nand U5637 (N_5637,N_4131,N_4147);
or U5638 (N_5638,N_4664,N_4152);
nor U5639 (N_5639,N_4558,N_4031);
nor U5640 (N_5640,N_4204,N_4384);
nand U5641 (N_5641,N_4897,N_4984);
nand U5642 (N_5642,N_4186,N_4165);
and U5643 (N_5643,N_4945,N_4355);
xor U5644 (N_5644,N_3890,N_4117);
nor U5645 (N_5645,N_4708,N_4882);
nand U5646 (N_5646,N_4695,N_4514);
nand U5647 (N_5647,N_4011,N_3999);
and U5648 (N_5648,N_4725,N_4582);
nor U5649 (N_5649,N_4822,N_4291);
nand U5650 (N_5650,N_4156,N_3862);
and U5651 (N_5651,N_3980,N_4004);
or U5652 (N_5652,N_4999,N_3977);
or U5653 (N_5653,N_4478,N_4578);
xnor U5654 (N_5654,N_4233,N_4129);
nand U5655 (N_5655,N_4063,N_4967);
xor U5656 (N_5656,N_4639,N_4614);
nand U5657 (N_5657,N_4238,N_4562);
nor U5658 (N_5658,N_3881,N_4230);
nand U5659 (N_5659,N_3977,N_4466);
nand U5660 (N_5660,N_4532,N_4670);
nor U5661 (N_5661,N_4781,N_4772);
nor U5662 (N_5662,N_4892,N_3904);
nor U5663 (N_5663,N_4385,N_3899);
xor U5664 (N_5664,N_4962,N_4689);
or U5665 (N_5665,N_4064,N_4166);
nor U5666 (N_5666,N_4434,N_4619);
xor U5667 (N_5667,N_3753,N_3750);
and U5668 (N_5668,N_4628,N_4215);
xnor U5669 (N_5669,N_3845,N_3968);
nand U5670 (N_5670,N_4102,N_4271);
nor U5671 (N_5671,N_4702,N_4798);
or U5672 (N_5672,N_4475,N_4379);
or U5673 (N_5673,N_4887,N_3935);
or U5674 (N_5674,N_3994,N_4493);
or U5675 (N_5675,N_4325,N_3771);
nand U5676 (N_5676,N_3837,N_4597);
nor U5677 (N_5677,N_4724,N_4272);
xor U5678 (N_5678,N_4480,N_4992);
nor U5679 (N_5679,N_4524,N_4377);
and U5680 (N_5680,N_4543,N_3851);
nand U5681 (N_5681,N_4309,N_4354);
nand U5682 (N_5682,N_4997,N_3758);
xor U5683 (N_5683,N_4235,N_4428);
or U5684 (N_5684,N_4481,N_4031);
xnor U5685 (N_5685,N_4595,N_3860);
nor U5686 (N_5686,N_4151,N_4624);
and U5687 (N_5687,N_4253,N_4265);
or U5688 (N_5688,N_4402,N_4944);
and U5689 (N_5689,N_3914,N_4106);
and U5690 (N_5690,N_4562,N_4436);
xor U5691 (N_5691,N_4475,N_4862);
xnor U5692 (N_5692,N_4727,N_4900);
and U5693 (N_5693,N_4313,N_4998);
nor U5694 (N_5694,N_4330,N_4438);
and U5695 (N_5695,N_4907,N_4555);
nor U5696 (N_5696,N_4647,N_4072);
nor U5697 (N_5697,N_4826,N_4914);
nor U5698 (N_5698,N_4847,N_4838);
xnor U5699 (N_5699,N_4156,N_4254);
or U5700 (N_5700,N_4274,N_4830);
nand U5701 (N_5701,N_4047,N_4408);
nor U5702 (N_5702,N_4862,N_4507);
and U5703 (N_5703,N_4073,N_4262);
nor U5704 (N_5704,N_4870,N_4668);
or U5705 (N_5705,N_4146,N_3900);
nor U5706 (N_5706,N_3843,N_4088);
or U5707 (N_5707,N_3837,N_4947);
nand U5708 (N_5708,N_4544,N_4579);
or U5709 (N_5709,N_4455,N_3822);
and U5710 (N_5710,N_4075,N_4604);
nor U5711 (N_5711,N_3918,N_4146);
nor U5712 (N_5712,N_3977,N_4331);
nand U5713 (N_5713,N_3895,N_4050);
xor U5714 (N_5714,N_3940,N_4867);
nor U5715 (N_5715,N_4897,N_4589);
or U5716 (N_5716,N_3815,N_3895);
xnor U5717 (N_5717,N_4718,N_4327);
nor U5718 (N_5718,N_4142,N_3805);
or U5719 (N_5719,N_3877,N_4596);
and U5720 (N_5720,N_4945,N_3905);
nand U5721 (N_5721,N_4234,N_4654);
nor U5722 (N_5722,N_3843,N_4579);
or U5723 (N_5723,N_4906,N_4810);
xor U5724 (N_5724,N_4567,N_4591);
nor U5725 (N_5725,N_4826,N_4207);
nand U5726 (N_5726,N_4392,N_3823);
nand U5727 (N_5727,N_4408,N_4793);
nand U5728 (N_5728,N_4957,N_4718);
xnor U5729 (N_5729,N_4541,N_4913);
and U5730 (N_5730,N_3762,N_4496);
xnor U5731 (N_5731,N_4001,N_4912);
nand U5732 (N_5732,N_4857,N_4226);
or U5733 (N_5733,N_4831,N_4072);
and U5734 (N_5734,N_4549,N_4475);
and U5735 (N_5735,N_3971,N_4366);
nor U5736 (N_5736,N_3822,N_4038);
or U5737 (N_5737,N_3871,N_4913);
nand U5738 (N_5738,N_4096,N_4247);
nor U5739 (N_5739,N_4884,N_4110);
and U5740 (N_5740,N_4957,N_4520);
xnor U5741 (N_5741,N_4345,N_4833);
or U5742 (N_5742,N_4480,N_4066);
or U5743 (N_5743,N_4898,N_4883);
xnor U5744 (N_5744,N_3988,N_4409);
and U5745 (N_5745,N_4695,N_4386);
xor U5746 (N_5746,N_4595,N_4909);
nor U5747 (N_5747,N_4516,N_4961);
or U5748 (N_5748,N_4287,N_4728);
nor U5749 (N_5749,N_4635,N_3934);
nor U5750 (N_5750,N_4734,N_4434);
or U5751 (N_5751,N_4949,N_4680);
and U5752 (N_5752,N_4124,N_3877);
or U5753 (N_5753,N_4981,N_4504);
nand U5754 (N_5754,N_4006,N_4961);
nand U5755 (N_5755,N_4837,N_4718);
or U5756 (N_5756,N_4924,N_4297);
xor U5757 (N_5757,N_4349,N_4328);
or U5758 (N_5758,N_3931,N_4181);
and U5759 (N_5759,N_4117,N_4794);
xor U5760 (N_5760,N_4236,N_4828);
xor U5761 (N_5761,N_4412,N_4754);
xnor U5762 (N_5762,N_4509,N_3757);
nor U5763 (N_5763,N_4673,N_4581);
or U5764 (N_5764,N_3883,N_4224);
nor U5765 (N_5765,N_4755,N_4081);
xnor U5766 (N_5766,N_4075,N_4951);
nor U5767 (N_5767,N_4514,N_4224);
or U5768 (N_5768,N_4052,N_3843);
and U5769 (N_5769,N_4117,N_4046);
xor U5770 (N_5770,N_4198,N_3998);
xor U5771 (N_5771,N_3871,N_4138);
or U5772 (N_5772,N_4101,N_4191);
nand U5773 (N_5773,N_4992,N_3977);
nor U5774 (N_5774,N_4698,N_3812);
or U5775 (N_5775,N_4791,N_4232);
xnor U5776 (N_5776,N_4903,N_4932);
xor U5777 (N_5777,N_4777,N_4057);
xor U5778 (N_5778,N_4109,N_4280);
nand U5779 (N_5779,N_3845,N_4190);
and U5780 (N_5780,N_4605,N_4746);
or U5781 (N_5781,N_4273,N_4700);
or U5782 (N_5782,N_4806,N_4468);
and U5783 (N_5783,N_4336,N_4961);
nor U5784 (N_5784,N_4385,N_3912);
xnor U5785 (N_5785,N_3753,N_4273);
xnor U5786 (N_5786,N_4978,N_4689);
nand U5787 (N_5787,N_3962,N_4605);
and U5788 (N_5788,N_4799,N_4261);
nor U5789 (N_5789,N_4474,N_4215);
or U5790 (N_5790,N_4822,N_3900);
and U5791 (N_5791,N_4644,N_4349);
xnor U5792 (N_5792,N_4587,N_4169);
and U5793 (N_5793,N_4802,N_4949);
xor U5794 (N_5794,N_4677,N_4530);
or U5795 (N_5795,N_4693,N_4660);
or U5796 (N_5796,N_4501,N_3918);
nand U5797 (N_5797,N_4575,N_4998);
and U5798 (N_5798,N_3779,N_4563);
nor U5799 (N_5799,N_4928,N_4328);
nand U5800 (N_5800,N_4942,N_4922);
xnor U5801 (N_5801,N_3893,N_4698);
and U5802 (N_5802,N_4086,N_4593);
xnor U5803 (N_5803,N_4500,N_3923);
nor U5804 (N_5804,N_4786,N_3758);
xnor U5805 (N_5805,N_4083,N_4210);
nand U5806 (N_5806,N_4431,N_4597);
xnor U5807 (N_5807,N_4220,N_3817);
and U5808 (N_5808,N_4344,N_4888);
xnor U5809 (N_5809,N_4923,N_4263);
and U5810 (N_5810,N_4908,N_3750);
nand U5811 (N_5811,N_4355,N_3842);
nor U5812 (N_5812,N_4049,N_4391);
nand U5813 (N_5813,N_4487,N_4229);
and U5814 (N_5814,N_4007,N_3777);
nand U5815 (N_5815,N_4327,N_3801);
nand U5816 (N_5816,N_4699,N_4174);
or U5817 (N_5817,N_4928,N_4046);
nor U5818 (N_5818,N_4641,N_4650);
or U5819 (N_5819,N_3901,N_3916);
and U5820 (N_5820,N_4660,N_3965);
or U5821 (N_5821,N_4482,N_4880);
nor U5822 (N_5822,N_4109,N_3855);
and U5823 (N_5823,N_4155,N_4925);
or U5824 (N_5824,N_4093,N_4788);
and U5825 (N_5825,N_4602,N_4725);
nand U5826 (N_5826,N_4464,N_4139);
xor U5827 (N_5827,N_4032,N_4309);
or U5828 (N_5828,N_4020,N_4964);
and U5829 (N_5829,N_4699,N_4026);
xor U5830 (N_5830,N_4927,N_4283);
nor U5831 (N_5831,N_4666,N_4403);
and U5832 (N_5832,N_3786,N_4467);
xor U5833 (N_5833,N_3854,N_4442);
nor U5834 (N_5834,N_4809,N_3955);
and U5835 (N_5835,N_4059,N_4249);
nor U5836 (N_5836,N_4679,N_3944);
xnor U5837 (N_5837,N_4112,N_4733);
nand U5838 (N_5838,N_4459,N_4666);
or U5839 (N_5839,N_4167,N_4520);
and U5840 (N_5840,N_4700,N_3795);
or U5841 (N_5841,N_3892,N_3815);
and U5842 (N_5842,N_4770,N_3815);
and U5843 (N_5843,N_3970,N_4967);
nand U5844 (N_5844,N_4742,N_4942);
or U5845 (N_5845,N_4976,N_3849);
nor U5846 (N_5846,N_4718,N_4948);
xor U5847 (N_5847,N_4156,N_3760);
nor U5848 (N_5848,N_4944,N_4147);
nand U5849 (N_5849,N_3904,N_3881);
nand U5850 (N_5850,N_4555,N_3979);
nor U5851 (N_5851,N_4667,N_3887);
nor U5852 (N_5852,N_4080,N_4078);
xor U5853 (N_5853,N_3877,N_4812);
and U5854 (N_5854,N_4858,N_4225);
nand U5855 (N_5855,N_4323,N_3802);
nand U5856 (N_5856,N_3804,N_4745);
nand U5857 (N_5857,N_4688,N_4513);
xnor U5858 (N_5858,N_4136,N_4750);
nand U5859 (N_5859,N_4352,N_4949);
nand U5860 (N_5860,N_4619,N_3902);
and U5861 (N_5861,N_4085,N_3793);
xnor U5862 (N_5862,N_3911,N_4963);
nand U5863 (N_5863,N_4659,N_4277);
nor U5864 (N_5864,N_4290,N_4621);
nor U5865 (N_5865,N_3857,N_4725);
or U5866 (N_5866,N_3882,N_3860);
or U5867 (N_5867,N_4299,N_4565);
nand U5868 (N_5868,N_4284,N_4247);
and U5869 (N_5869,N_4693,N_4027);
and U5870 (N_5870,N_3897,N_4541);
nand U5871 (N_5871,N_4846,N_3973);
xnor U5872 (N_5872,N_3890,N_4096);
xnor U5873 (N_5873,N_4516,N_4333);
nor U5874 (N_5874,N_4246,N_4623);
nor U5875 (N_5875,N_4372,N_4633);
and U5876 (N_5876,N_4419,N_4955);
or U5877 (N_5877,N_4650,N_4723);
nor U5878 (N_5878,N_4190,N_4789);
nor U5879 (N_5879,N_4757,N_3766);
nor U5880 (N_5880,N_4897,N_4709);
and U5881 (N_5881,N_4239,N_4595);
xnor U5882 (N_5882,N_4270,N_4766);
nor U5883 (N_5883,N_4078,N_4184);
nand U5884 (N_5884,N_4802,N_4761);
nand U5885 (N_5885,N_4476,N_4668);
and U5886 (N_5886,N_4065,N_4948);
nand U5887 (N_5887,N_4049,N_4333);
xnor U5888 (N_5888,N_4248,N_4204);
nor U5889 (N_5889,N_4709,N_4484);
and U5890 (N_5890,N_4135,N_4540);
nor U5891 (N_5891,N_4722,N_4679);
or U5892 (N_5892,N_4300,N_4238);
or U5893 (N_5893,N_4965,N_4499);
nand U5894 (N_5894,N_4169,N_4943);
nand U5895 (N_5895,N_4516,N_3897);
xor U5896 (N_5896,N_4581,N_4331);
nand U5897 (N_5897,N_3937,N_3934);
or U5898 (N_5898,N_4311,N_4524);
nand U5899 (N_5899,N_4677,N_4906);
or U5900 (N_5900,N_4783,N_4366);
xor U5901 (N_5901,N_4673,N_4762);
and U5902 (N_5902,N_4594,N_4404);
and U5903 (N_5903,N_4997,N_3776);
and U5904 (N_5904,N_3761,N_4928);
nand U5905 (N_5905,N_4798,N_4125);
xor U5906 (N_5906,N_4371,N_3968);
nand U5907 (N_5907,N_4487,N_4483);
or U5908 (N_5908,N_4604,N_4283);
xnor U5909 (N_5909,N_4874,N_4889);
nand U5910 (N_5910,N_3870,N_4708);
xor U5911 (N_5911,N_4475,N_3906);
and U5912 (N_5912,N_4427,N_4598);
xnor U5913 (N_5913,N_4312,N_4248);
nor U5914 (N_5914,N_4629,N_4901);
or U5915 (N_5915,N_4961,N_4618);
nand U5916 (N_5916,N_4898,N_4834);
or U5917 (N_5917,N_4811,N_4329);
or U5918 (N_5918,N_4504,N_3863);
xnor U5919 (N_5919,N_4528,N_3760);
or U5920 (N_5920,N_3876,N_3874);
nand U5921 (N_5921,N_4062,N_4363);
or U5922 (N_5922,N_4552,N_4660);
or U5923 (N_5923,N_4899,N_4990);
and U5924 (N_5924,N_4467,N_3863);
xor U5925 (N_5925,N_4367,N_4578);
or U5926 (N_5926,N_3996,N_3852);
xor U5927 (N_5927,N_3993,N_4090);
and U5928 (N_5928,N_4606,N_3812);
or U5929 (N_5929,N_4266,N_3999);
and U5930 (N_5930,N_4585,N_4499);
nor U5931 (N_5931,N_4145,N_4590);
nor U5932 (N_5932,N_4862,N_4498);
and U5933 (N_5933,N_3754,N_4897);
nor U5934 (N_5934,N_4859,N_4527);
and U5935 (N_5935,N_4599,N_3869);
and U5936 (N_5936,N_4258,N_4912);
nand U5937 (N_5937,N_4863,N_3939);
nor U5938 (N_5938,N_4509,N_4399);
and U5939 (N_5939,N_3992,N_3939);
nor U5940 (N_5940,N_4507,N_4404);
xor U5941 (N_5941,N_4912,N_4613);
nand U5942 (N_5942,N_4099,N_4859);
nand U5943 (N_5943,N_4521,N_4811);
xnor U5944 (N_5944,N_4474,N_4944);
or U5945 (N_5945,N_4108,N_4678);
nand U5946 (N_5946,N_4390,N_4375);
nand U5947 (N_5947,N_4138,N_4444);
xnor U5948 (N_5948,N_4803,N_4981);
nor U5949 (N_5949,N_4988,N_4006);
or U5950 (N_5950,N_4960,N_4704);
xor U5951 (N_5951,N_4901,N_3775);
nor U5952 (N_5952,N_4817,N_4127);
xnor U5953 (N_5953,N_4627,N_4115);
nand U5954 (N_5954,N_4271,N_4763);
xor U5955 (N_5955,N_4613,N_4483);
or U5956 (N_5956,N_4859,N_4759);
or U5957 (N_5957,N_4512,N_4374);
or U5958 (N_5958,N_4155,N_4450);
xnor U5959 (N_5959,N_4311,N_4610);
xor U5960 (N_5960,N_4234,N_4357);
xnor U5961 (N_5961,N_4850,N_4699);
or U5962 (N_5962,N_4694,N_4357);
xnor U5963 (N_5963,N_4189,N_4632);
nor U5964 (N_5964,N_4007,N_4479);
nand U5965 (N_5965,N_4773,N_4126);
and U5966 (N_5966,N_4721,N_4702);
nor U5967 (N_5967,N_4491,N_3764);
and U5968 (N_5968,N_4257,N_3787);
nand U5969 (N_5969,N_4234,N_3831);
nor U5970 (N_5970,N_4747,N_4807);
nand U5971 (N_5971,N_4063,N_4830);
or U5972 (N_5972,N_4526,N_4254);
or U5973 (N_5973,N_4789,N_4225);
nor U5974 (N_5974,N_4186,N_4791);
nand U5975 (N_5975,N_4664,N_4270);
or U5976 (N_5976,N_4682,N_4798);
nand U5977 (N_5977,N_4440,N_3829);
nor U5978 (N_5978,N_4454,N_4861);
and U5979 (N_5979,N_4104,N_4530);
xnor U5980 (N_5980,N_4910,N_4683);
nor U5981 (N_5981,N_4845,N_4736);
or U5982 (N_5982,N_4577,N_4192);
and U5983 (N_5983,N_3823,N_4458);
nor U5984 (N_5984,N_4045,N_3942);
and U5985 (N_5985,N_3933,N_4247);
nand U5986 (N_5986,N_4896,N_4573);
or U5987 (N_5987,N_4849,N_3826);
and U5988 (N_5988,N_4481,N_4854);
xnor U5989 (N_5989,N_4557,N_3806);
xor U5990 (N_5990,N_4991,N_4655);
xnor U5991 (N_5991,N_4866,N_3820);
nor U5992 (N_5992,N_4873,N_4474);
xnor U5993 (N_5993,N_4761,N_4451);
and U5994 (N_5994,N_4990,N_3973);
and U5995 (N_5995,N_4551,N_4836);
nand U5996 (N_5996,N_4903,N_4939);
or U5997 (N_5997,N_4916,N_4441);
nand U5998 (N_5998,N_4300,N_4032);
and U5999 (N_5999,N_4452,N_4347);
nand U6000 (N_6000,N_4029,N_4948);
or U6001 (N_6001,N_4627,N_4318);
xnor U6002 (N_6002,N_4764,N_4950);
or U6003 (N_6003,N_4918,N_4510);
nand U6004 (N_6004,N_4456,N_4789);
and U6005 (N_6005,N_4606,N_3817);
or U6006 (N_6006,N_4209,N_3861);
nor U6007 (N_6007,N_4185,N_4145);
nand U6008 (N_6008,N_4867,N_4340);
xnor U6009 (N_6009,N_4848,N_4266);
or U6010 (N_6010,N_4571,N_4986);
nand U6011 (N_6011,N_4237,N_3753);
and U6012 (N_6012,N_4690,N_3883);
and U6013 (N_6013,N_4782,N_4909);
nor U6014 (N_6014,N_4558,N_4305);
and U6015 (N_6015,N_3895,N_4530);
xor U6016 (N_6016,N_4183,N_4241);
xor U6017 (N_6017,N_4020,N_3770);
and U6018 (N_6018,N_4127,N_4747);
and U6019 (N_6019,N_4760,N_4066);
or U6020 (N_6020,N_4499,N_4145);
or U6021 (N_6021,N_4343,N_4209);
nor U6022 (N_6022,N_4574,N_3818);
or U6023 (N_6023,N_4362,N_4802);
nor U6024 (N_6024,N_4706,N_4232);
xnor U6025 (N_6025,N_4222,N_4220);
nor U6026 (N_6026,N_4999,N_4010);
or U6027 (N_6027,N_3851,N_4663);
nand U6028 (N_6028,N_4798,N_4614);
xor U6029 (N_6029,N_4235,N_4897);
or U6030 (N_6030,N_4436,N_4616);
and U6031 (N_6031,N_4463,N_3898);
nor U6032 (N_6032,N_4548,N_4533);
nand U6033 (N_6033,N_4288,N_4579);
nor U6034 (N_6034,N_4181,N_3792);
nand U6035 (N_6035,N_3906,N_4952);
nor U6036 (N_6036,N_3801,N_4170);
or U6037 (N_6037,N_4578,N_4256);
xor U6038 (N_6038,N_4011,N_4991);
or U6039 (N_6039,N_4329,N_4718);
nor U6040 (N_6040,N_4462,N_4490);
xnor U6041 (N_6041,N_4253,N_4758);
nand U6042 (N_6042,N_4532,N_3900);
nand U6043 (N_6043,N_4769,N_4615);
and U6044 (N_6044,N_4447,N_4893);
nor U6045 (N_6045,N_4332,N_4882);
and U6046 (N_6046,N_4650,N_4881);
and U6047 (N_6047,N_4923,N_4688);
and U6048 (N_6048,N_4004,N_3848);
nand U6049 (N_6049,N_4138,N_4455);
or U6050 (N_6050,N_3965,N_4981);
and U6051 (N_6051,N_4286,N_4745);
or U6052 (N_6052,N_4299,N_4650);
nand U6053 (N_6053,N_4804,N_4512);
or U6054 (N_6054,N_4357,N_4245);
or U6055 (N_6055,N_3780,N_4458);
nand U6056 (N_6056,N_4616,N_4682);
nand U6057 (N_6057,N_4866,N_3858);
or U6058 (N_6058,N_4155,N_3909);
and U6059 (N_6059,N_4803,N_3828);
nor U6060 (N_6060,N_3950,N_4550);
or U6061 (N_6061,N_4852,N_4005);
nor U6062 (N_6062,N_4255,N_4402);
and U6063 (N_6063,N_4123,N_4979);
nor U6064 (N_6064,N_3822,N_3795);
nand U6065 (N_6065,N_4218,N_3992);
xnor U6066 (N_6066,N_4037,N_3923);
and U6067 (N_6067,N_4737,N_4025);
nor U6068 (N_6068,N_4341,N_4127);
nor U6069 (N_6069,N_4900,N_4793);
and U6070 (N_6070,N_4937,N_3906);
xnor U6071 (N_6071,N_4200,N_4095);
nor U6072 (N_6072,N_4859,N_3851);
xnor U6073 (N_6073,N_4529,N_3786);
nor U6074 (N_6074,N_4567,N_4338);
nor U6075 (N_6075,N_4182,N_3986);
and U6076 (N_6076,N_4416,N_4197);
xor U6077 (N_6077,N_4276,N_4013);
or U6078 (N_6078,N_4122,N_4159);
and U6079 (N_6079,N_4574,N_4537);
nor U6080 (N_6080,N_4889,N_4333);
xor U6081 (N_6081,N_4989,N_4088);
nor U6082 (N_6082,N_4400,N_4969);
nor U6083 (N_6083,N_3791,N_4347);
xor U6084 (N_6084,N_3985,N_4496);
and U6085 (N_6085,N_4409,N_4086);
or U6086 (N_6086,N_3797,N_4748);
nor U6087 (N_6087,N_4798,N_4622);
and U6088 (N_6088,N_4312,N_4283);
or U6089 (N_6089,N_3882,N_4844);
or U6090 (N_6090,N_4111,N_4519);
nand U6091 (N_6091,N_4931,N_3851);
and U6092 (N_6092,N_4371,N_4669);
nor U6093 (N_6093,N_3945,N_4989);
xor U6094 (N_6094,N_4972,N_3753);
nand U6095 (N_6095,N_4467,N_3894);
and U6096 (N_6096,N_4078,N_4848);
nor U6097 (N_6097,N_4647,N_4817);
xnor U6098 (N_6098,N_4224,N_4503);
and U6099 (N_6099,N_4931,N_3907);
xor U6100 (N_6100,N_3810,N_4637);
nor U6101 (N_6101,N_4226,N_4855);
nand U6102 (N_6102,N_4051,N_3902);
and U6103 (N_6103,N_3991,N_4035);
nand U6104 (N_6104,N_4074,N_4941);
nor U6105 (N_6105,N_4176,N_4491);
nor U6106 (N_6106,N_4475,N_3814);
nand U6107 (N_6107,N_3763,N_3815);
and U6108 (N_6108,N_4539,N_4750);
nand U6109 (N_6109,N_4608,N_4135);
nor U6110 (N_6110,N_4958,N_3804);
xor U6111 (N_6111,N_4064,N_4187);
nor U6112 (N_6112,N_4871,N_4489);
xor U6113 (N_6113,N_4919,N_4807);
nor U6114 (N_6114,N_3874,N_3856);
nor U6115 (N_6115,N_4806,N_4910);
xor U6116 (N_6116,N_4342,N_3765);
and U6117 (N_6117,N_4821,N_4839);
and U6118 (N_6118,N_4473,N_4023);
xnor U6119 (N_6119,N_4913,N_4224);
or U6120 (N_6120,N_3800,N_4770);
or U6121 (N_6121,N_4561,N_3982);
xnor U6122 (N_6122,N_3816,N_4503);
nand U6123 (N_6123,N_4179,N_4610);
nor U6124 (N_6124,N_4999,N_3852);
xnor U6125 (N_6125,N_3993,N_4545);
or U6126 (N_6126,N_4995,N_4208);
xor U6127 (N_6127,N_3853,N_4341);
nor U6128 (N_6128,N_4216,N_3905);
xnor U6129 (N_6129,N_4925,N_4354);
or U6130 (N_6130,N_3817,N_4573);
nor U6131 (N_6131,N_3881,N_4416);
nor U6132 (N_6132,N_3922,N_4393);
or U6133 (N_6133,N_4199,N_4133);
nor U6134 (N_6134,N_3811,N_4464);
xor U6135 (N_6135,N_4064,N_4228);
and U6136 (N_6136,N_3871,N_4751);
nor U6137 (N_6137,N_4623,N_4421);
xnor U6138 (N_6138,N_4689,N_3788);
and U6139 (N_6139,N_4260,N_4163);
or U6140 (N_6140,N_4000,N_4614);
nor U6141 (N_6141,N_3879,N_4237);
and U6142 (N_6142,N_3952,N_4556);
nor U6143 (N_6143,N_4547,N_3943);
nand U6144 (N_6144,N_3895,N_3766);
nor U6145 (N_6145,N_3860,N_4434);
and U6146 (N_6146,N_4005,N_3771);
nor U6147 (N_6147,N_3941,N_4737);
or U6148 (N_6148,N_4914,N_4934);
or U6149 (N_6149,N_3815,N_3864);
nor U6150 (N_6150,N_4393,N_4553);
nand U6151 (N_6151,N_3810,N_4765);
xor U6152 (N_6152,N_4875,N_4161);
or U6153 (N_6153,N_3920,N_4102);
nor U6154 (N_6154,N_4323,N_4266);
and U6155 (N_6155,N_4455,N_4027);
nand U6156 (N_6156,N_4004,N_4907);
nand U6157 (N_6157,N_4743,N_4965);
nor U6158 (N_6158,N_4807,N_4121);
nor U6159 (N_6159,N_4776,N_4750);
xor U6160 (N_6160,N_4688,N_4088);
nor U6161 (N_6161,N_4915,N_4285);
or U6162 (N_6162,N_4210,N_4524);
or U6163 (N_6163,N_4685,N_3816);
nor U6164 (N_6164,N_4552,N_4692);
nor U6165 (N_6165,N_4160,N_4777);
nand U6166 (N_6166,N_4818,N_4875);
nor U6167 (N_6167,N_4583,N_4239);
and U6168 (N_6168,N_3825,N_4668);
or U6169 (N_6169,N_4744,N_3902);
and U6170 (N_6170,N_3837,N_4367);
nand U6171 (N_6171,N_4403,N_4004);
nand U6172 (N_6172,N_4526,N_4767);
xor U6173 (N_6173,N_4129,N_4408);
nand U6174 (N_6174,N_3776,N_3813);
nand U6175 (N_6175,N_4291,N_4767);
nand U6176 (N_6176,N_4793,N_3985);
nor U6177 (N_6177,N_4717,N_4473);
or U6178 (N_6178,N_4150,N_4310);
or U6179 (N_6179,N_4008,N_4543);
nand U6180 (N_6180,N_4854,N_4120);
and U6181 (N_6181,N_4060,N_3933);
or U6182 (N_6182,N_3837,N_4968);
nand U6183 (N_6183,N_4780,N_4166);
nor U6184 (N_6184,N_4992,N_4169);
nand U6185 (N_6185,N_4494,N_4117);
and U6186 (N_6186,N_4512,N_4504);
nand U6187 (N_6187,N_3970,N_4572);
or U6188 (N_6188,N_4483,N_4548);
nor U6189 (N_6189,N_3797,N_4891);
nand U6190 (N_6190,N_4874,N_4315);
and U6191 (N_6191,N_4478,N_4515);
xnor U6192 (N_6192,N_3775,N_4171);
nor U6193 (N_6193,N_4193,N_4130);
nor U6194 (N_6194,N_4256,N_3976);
and U6195 (N_6195,N_3770,N_4802);
and U6196 (N_6196,N_4110,N_4444);
nor U6197 (N_6197,N_4834,N_4948);
nand U6198 (N_6198,N_4334,N_4065);
xor U6199 (N_6199,N_4177,N_4570);
xor U6200 (N_6200,N_4002,N_4261);
xnor U6201 (N_6201,N_3837,N_4361);
xnor U6202 (N_6202,N_3948,N_4994);
nor U6203 (N_6203,N_4399,N_4719);
and U6204 (N_6204,N_4590,N_4822);
nor U6205 (N_6205,N_4145,N_4271);
and U6206 (N_6206,N_4673,N_4217);
nand U6207 (N_6207,N_4680,N_3997);
or U6208 (N_6208,N_4056,N_4009);
and U6209 (N_6209,N_4760,N_4681);
and U6210 (N_6210,N_4271,N_4404);
nand U6211 (N_6211,N_3865,N_4960);
xor U6212 (N_6212,N_4211,N_4660);
nor U6213 (N_6213,N_4632,N_3921);
or U6214 (N_6214,N_4952,N_4612);
or U6215 (N_6215,N_4400,N_4681);
nor U6216 (N_6216,N_4163,N_3811);
xnor U6217 (N_6217,N_4539,N_3799);
nand U6218 (N_6218,N_4596,N_4810);
nand U6219 (N_6219,N_4534,N_4298);
xnor U6220 (N_6220,N_3910,N_4985);
nand U6221 (N_6221,N_4497,N_3825);
nand U6222 (N_6222,N_3847,N_4578);
and U6223 (N_6223,N_4490,N_3805);
xor U6224 (N_6224,N_3813,N_4632);
nand U6225 (N_6225,N_4309,N_3852);
xor U6226 (N_6226,N_4484,N_4235);
nand U6227 (N_6227,N_4686,N_3962);
nand U6228 (N_6228,N_4214,N_3993);
nor U6229 (N_6229,N_4266,N_4146);
or U6230 (N_6230,N_3867,N_4251);
or U6231 (N_6231,N_4842,N_4039);
nand U6232 (N_6232,N_4955,N_4361);
xnor U6233 (N_6233,N_4839,N_4382);
or U6234 (N_6234,N_4803,N_4795);
or U6235 (N_6235,N_3966,N_4656);
and U6236 (N_6236,N_4128,N_4218);
nand U6237 (N_6237,N_4758,N_4056);
xnor U6238 (N_6238,N_4785,N_3992);
xor U6239 (N_6239,N_4223,N_4513);
and U6240 (N_6240,N_4487,N_4476);
nor U6241 (N_6241,N_4131,N_4765);
and U6242 (N_6242,N_3767,N_4732);
or U6243 (N_6243,N_3959,N_4382);
nand U6244 (N_6244,N_4409,N_4775);
nand U6245 (N_6245,N_4860,N_3981);
or U6246 (N_6246,N_4902,N_4614);
and U6247 (N_6247,N_4470,N_4795);
and U6248 (N_6248,N_3816,N_4408);
or U6249 (N_6249,N_4989,N_4730);
nor U6250 (N_6250,N_6147,N_5199);
nand U6251 (N_6251,N_5882,N_5796);
nor U6252 (N_6252,N_5202,N_5488);
xnor U6253 (N_6253,N_5910,N_5980);
nand U6254 (N_6254,N_5175,N_5942);
xnor U6255 (N_6255,N_5244,N_5286);
nand U6256 (N_6256,N_5473,N_5191);
and U6257 (N_6257,N_6041,N_5737);
and U6258 (N_6258,N_5059,N_6005);
nor U6259 (N_6259,N_5100,N_5197);
xnor U6260 (N_6260,N_5109,N_6039);
xor U6261 (N_6261,N_5088,N_5502);
and U6262 (N_6262,N_5990,N_5805);
or U6263 (N_6263,N_5659,N_6053);
nand U6264 (N_6264,N_5650,N_6152);
and U6265 (N_6265,N_5628,N_5418);
or U6266 (N_6266,N_6232,N_5490);
nor U6267 (N_6267,N_5698,N_5128);
or U6268 (N_6268,N_5417,N_5551);
nand U6269 (N_6269,N_5918,N_6081);
and U6270 (N_6270,N_5376,N_5930);
and U6271 (N_6271,N_5086,N_5213);
nand U6272 (N_6272,N_5791,N_5906);
nand U6273 (N_6273,N_5851,N_5187);
xor U6274 (N_6274,N_5716,N_6032);
and U6275 (N_6275,N_5093,N_5750);
or U6276 (N_6276,N_6000,N_5526);
nand U6277 (N_6277,N_5949,N_5630);
nand U6278 (N_6278,N_5255,N_5669);
or U6279 (N_6279,N_5766,N_6084);
or U6280 (N_6280,N_5829,N_5308);
nand U6281 (N_6281,N_6087,N_5617);
nor U6282 (N_6282,N_5683,N_5374);
nor U6283 (N_6283,N_5578,N_5470);
xnor U6284 (N_6284,N_5641,N_5472);
and U6285 (N_6285,N_5667,N_5499);
nand U6286 (N_6286,N_5133,N_5728);
nor U6287 (N_6287,N_5537,N_5642);
or U6288 (N_6288,N_5858,N_5575);
xnor U6289 (N_6289,N_5733,N_5127);
xor U6290 (N_6290,N_6141,N_5515);
xor U6291 (N_6291,N_5184,N_5715);
nor U6292 (N_6292,N_5913,N_5973);
xor U6293 (N_6293,N_5707,N_6192);
nand U6294 (N_6294,N_5168,N_5269);
and U6295 (N_6295,N_6221,N_5521);
or U6296 (N_6296,N_5223,N_5686);
or U6297 (N_6297,N_6091,N_5289);
xor U6298 (N_6298,N_5640,N_5006);
nand U6299 (N_6299,N_5020,N_5662);
xnor U6300 (N_6300,N_5013,N_5850);
nor U6301 (N_6301,N_5482,N_5562);
xor U6302 (N_6302,N_5649,N_5679);
and U6303 (N_6303,N_5305,N_5954);
xnor U6304 (N_6304,N_5206,N_5964);
nand U6305 (N_6305,N_5671,N_5437);
and U6306 (N_6306,N_6101,N_5345);
or U6307 (N_6307,N_5124,N_5183);
or U6308 (N_6308,N_5518,N_5262);
and U6309 (N_6309,N_5752,N_6003);
xor U6310 (N_6310,N_6138,N_6227);
or U6311 (N_6311,N_5844,N_5756);
nor U6312 (N_6312,N_5665,N_5448);
nor U6313 (N_6313,N_5167,N_5280);
xnor U6314 (N_6314,N_6212,N_6204);
nand U6315 (N_6315,N_6109,N_5123);
nand U6316 (N_6316,N_5384,N_5445);
nand U6317 (N_6317,N_5792,N_5517);
and U6318 (N_6318,N_6054,N_6052);
nor U6319 (N_6319,N_5081,N_6049);
or U6320 (N_6320,N_5079,N_6243);
nand U6321 (N_6321,N_5297,N_5090);
or U6322 (N_6322,N_5390,N_5357);
nand U6323 (N_6323,N_5238,N_6067);
nor U6324 (N_6324,N_5353,N_5233);
xor U6325 (N_6325,N_5475,N_6133);
nor U6326 (N_6326,N_5877,N_6105);
or U6327 (N_6327,N_6010,N_5443);
nand U6328 (N_6328,N_5044,N_6045);
and U6329 (N_6329,N_5959,N_6124);
nor U6330 (N_6330,N_5739,N_5977);
xor U6331 (N_6331,N_6198,N_5565);
nor U6332 (N_6332,N_5346,N_6034);
xnor U6333 (N_6333,N_5343,N_5011);
or U6334 (N_6334,N_6188,N_5666);
or U6335 (N_6335,N_5697,N_5434);
or U6336 (N_6336,N_5382,N_5997);
nor U6337 (N_6337,N_5950,N_5180);
xnor U6338 (N_6338,N_6040,N_5788);
xnor U6339 (N_6339,N_5208,N_5724);
xnor U6340 (N_6340,N_6161,N_6072);
xor U6341 (N_6341,N_5420,N_5084);
and U6342 (N_6342,N_5531,N_5073);
nor U6343 (N_6343,N_5237,N_5111);
xor U6344 (N_6344,N_5657,N_5317);
and U6345 (N_6345,N_5461,N_5224);
nor U6346 (N_6346,N_5933,N_5916);
nand U6347 (N_6347,N_5115,N_5614);
nand U6348 (N_6348,N_5102,N_5141);
and U6349 (N_6349,N_6136,N_5035);
or U6350 (N_6350,N_6203,N_5275);
xnor U6351 (N_6351,N_5825,N_5572);
nand U6352 (N_6352,N_5622,N_5075);
nand U6353 (N_6353,N_5188,N_5032);
xor U6354 (N_6354,N_5014,N_5501);
and U6355 (N_6355,N_5156,N_5591);
xnor U6356 (N_6356,N_5982,N_6128);
or U6357 (N_6357,N_5594,N_6144);
xor U6358 (N_6358,N_6015,N_5999);
nand U6359 (N_6359,N_6107,N_5493);
or U6360 (N_6360,N_5822,N_5413);
or U6361 (N_6361,N_5462,N_5178);
and U6362 (N_6362,N_5896,N_5777);
xor U6363 (N_6363,N_6169,N_6083);
or U6364 (N_6364,N_5052,N_5423);
nand U6365 (N_6365,N_5498,N_5476);
and U6366 (N_6366,N_6085,N_5046);
nand U6367 (N_6367,N_5672,N_5455);
xor U6368 (N_6368,N_5266,N_5547);
xor U6369 (N_6369,N_5027,N_5638);
xnor U6370 (N_6370,N_5512,N_5323);
or U6371 (N_6371,N_5467,N_5542);
nand U6372 (N_6372,N_5878,N_6194);
xor U6373 (N_6373,N_5385,N_5500);
and U6374 (N_6374,N_5532,N_5194);
nand U6375 (N_6375,N_5313,N_5159);
nand U6376 (N_6376,N_6055,N_5274);
nor U6377 (N_6377,N_6125,N_5583);
xnor U6378 (N_6378,N_6095,N_6234);
nor U6379 (N_6379,N_5963,N_6225);
and U6380 (N_6380,N_5938,N_5969);
nor U6381 (N_6381,N_5053,N_5925);
or U6382 (N_6382,N_5377,N_5061);
nor U6383 (N_6383,N_5908,N_5145);
nor U6384 (N_6384,N_5058,N_5104);
nand U6385 (N_6385,N_5380,N_5107);
nand U6386 (N_6386,N_5051,N_5734);
and U6387 (N_6387,N_6193,N_5464);
and U6388 (N_6388,N_5827,N_5338);
nand U6389 (N_6389,N_5398,N_5173);
or U6390 (N_6390,N_5264,N_5060);
and U6391 (N_6391,N_5272,N_5391);
nor U6392 (N_6392,N_6209,N_5181);
or U6393 (N_6393,N_6154,N_5101);
nand U6394 (N_6394,N_5694,N_6071);
and U6395 (N_6395,N_5875,N_5099);
nand U6396 (N_6396,N_5745,N_5900);
nand U6397 (N_6397,N_5821,N_5163);
and U6398 (N_6398,N_5587,N_6143);
and U6399 (N_6399,N_5782,N_5325);
or U6400 (N_6400,N_5207,N_6206);
or U6401 (N_6401,N_5215,N_5430);
nor U6402 (N_6402,N_5684,N_5336);
nand U6403 (N_6403,N_5172,N_5496);
xnor U6404 (N_6404,N_5431,N_5826);
xor U6405 (N_6405,N_5072,N_6146);
xor U6406 (N_6406,N_5477,N_5373);
nand U6407 (N_6407,N_5403,N_5301);
or U6408 (N_6408,N_5130,N_5946);
xor U6409 (N_6409,N_5371,N_5656);
and U6410 (N_6410,N_5597,N_5315);
nor U6411 (N_6411,N_5593,N_5911);
or U6412 (N_6412,N_6007,N_6176);
nor U6413 (N_6413,N_5541,N_5419);
nand U6414 (N_6414,N_6102,N_5263);
nand U6415 (N_6415,N_5654,N_6199);
nand U6416 (N_6416,N_5394,N_5146);
xor U6417 (N_6417,N_5387,N_5375);
xor U6418 (N_6418,N_5732,N_5355);
nand U6419 (N_6419,N_5234,N_6082);
and U6420 (N_6420,N_5625,N_5389);
nor U6421 (N_6421,N_6051,N_6249);
nand U6422 (N_6422,N_5564,N_6175);
xnor U6423 (N_6423,N_6189,N_6111);
nand U6424 (N_6424,N_5074,N_5432);
nand U6425 (N_6425,N_6150,N_6057);
nor U6426 (N_6426,N_5801,N_5504);
nor U6427 (N_6427,N_5474,N_5205);
nand U6428 (N_6428,N_5189,N_5953);
and U6429 (N_6429,N_5056,N_6219);
or U6430 (N_6430,N_5701,N_6205);
nor U6431 (N_6431,N_6190,N_6118);
nand U6432 (N_6432,N_5571,N_6166);
xnor U6433 (N_6433,N_5383,N_5256);
nand U6434 (N_6434,N_5116,N_5247);
nor U6435 (N_6435,N_5307,N_5129);
nand U6436 (N_6436,N_5018,N_5807);
or U6437 (N_6437,N_5726,N_5166);
nor U6438 (N_6438,N_5704,N_6173);
nor U6439 (N_6439,N_5566,N_5426);
or U6440 (N_6440,N_5246,N_5700);
xnor U6441 (N_6441,N_5555,N_5548);
or U6442 (N_6442,N_5958,N_5160);
nand U6443 (N_6443,N_5868,N_5561);
nor U6444 (N_6444,N_5103,N_6079);
and U6445 (N_6445,N_5261,N_5321);
nand U6446 (N_6446,N_5012,N_5717);
nand U6447 (N_6447,N_5795,N_5125);
xnor U6448 (N_6448,N_5652,N_5438);
nor U6449 (N_6449,N_5076,N_5457);
xnor U6450 (N_6450,N_5753,N_5161);
nor U6451 (N_6451,N_6020,N_5574);
xor U6452 (N_6452,N_6027,N_5507);
or U6453 (N_6453,N_5558,N_5968);
or U6454 (N_6454,N_5624,N_5019);
nor U6455 (N_6455,N_5023,N_5522);
nor U6456 (N_6456,N_5303,N_5055);
or U6457 (N_6457,N_5809,N_6037);
or U6458 (N_6458,N_6122,N_5509);
xnor U6459 (N_6459,N_5126,N_5573);
xor U6460 (N_6460,N_5468,N_6035);
or U6461 (N_6461,N_6014,N_5190);
or U6462 (N_6462,N_6047,N_5031);
and U6463 (N_6463,N_5370,N_6202);
nor U6464 (N_6464,N_5550,N_6210);
nand U6465 (N_6465,N_5563,N_6145);
and U6466 (N_6466,N_5143,N_5904);
nor U6467 (N_6467,N_6117,N_6215);
or U6468 (N_6468,N_5038,N_5216);
and U6469 (N_6469,N_5632,N_5048);
or U6470 (N_6470,N_5281,N_5861);
nor U6471 (N_6471,N_5252,N_5395);
nand U6472 (N_6472,N_5460,N_5818);
nor U6473 (N_6473,N_6213,N_5581);
or U6474 (N_6474,N_5714,N_5556);
and U6475 (N_6475,N_5872,N_5901);
nand U6476 (N_6476,N_5322,N_5582);
and U6477 (N_6477,N_6038,N_6123);
nor U6478 (N_6478,N_5740,N_5506);
nand U6479 (N_6479,N_5298,N_5170);
nor U6480 (N_6480,N_5951,N_5863);
nor U6481 (N_6481,N_5235,N_6247);
and U6482 (N_6482,N_5781,N_5560);
xnor U6483 (N_6483,N_5691,N_5042);
or U6484 (N_6484,N_6248,N_5520);
or U6485 (N_6485,N_5559,N_5282);
nor U6486 (N_6486,N_5152,N_5203);
or U6487 (N_6487,N_5033,N_5983);
nand U6488 (N_6488,N_5505,N_5530);
and U6489 (N_6489,N_6228,N_5940);
nand U6490 (N_6490,N_5293,N_5804);
and U6491 (N_6491,N_5670,N_6241);
or U6492 (N_6492,N_6028,N_5705);
nand U6493 (N_6493,N_5544,N_5962);
and U6494 (N_6494,N_5250,N_5318);
nor U6495 (N_6495,N_5794,N_5535);
nor U6496 (N_6496,N_5253,N_5491);
xor U6497 (N_6497,N_5956,N_5897);
and U6498 (N_6498,N_5119,N_5689);
and U6499 (N_6499,N_6030,N_6177);
or U6500 (N_6500,N_5273,N_5957);
nand U6501 (N_6501,N_5337,N_6093);
or U6502 (N_6502,N_5779,N_6024);
xor U6503 (N_6503,N_5598,N_5121);
and U6504 (N_6504,N_5955,N_5618);
or U6505 (N_6505,N_5586,N_6131);
or U6506 (N_6506,N_5142,N_5139);
xnor U6507 (N_6507,N_5894,N_5041);
xnor U6508 (N_6508,N_5828,N_5135);
xor U6509 (N_6509,N_5113,N_5211);
and U6510 (N_6510,N_5935,N_5040);
nor U6511 (N_6511,N_5352,N_5711);
and U6512 (N_6512,N_5446,N_5162);
or U6513 (N_6513,N_5047,N_6006);
nor U6514 (N_6514,N_5816,N_5703);
nor U6515 (N_6515,N_5533,N_5481);
nor U6516 (N_6516,N_5960,N_5007);
nor U6517 (N_6517,N_5616,N_5106);
and U6518 (N_6518,N_6086,N_5010);
nor U6519 (N_6519,N_5415,N_6069);
and U6520 (N_6520,N_5105,N_5772);
xnor U6521 (N_6521,N_5839,N_5865);
nand U6522 (N_6522,N_6226,N_5629);
nand U6523 (N_6523,N_5379,N_5880);
nor U6524 (N_6524,N_5721,N_5834);
or U6525 (N_6525,N_5277,N_5165);
and U6526 (N_6526,N_5751,N_5429);
xnor U6527 (N_6527,N_5069,N_6075);
nand U6528 (N_6528,N_5433,N_5903);
and U6529 (N_6529,N_5201,N_5929);
nand U6530 (N_6530,N_5236,N_6004);
nand U6531 (N_6531,N_5319,N_6246);
nand U6532 (N_6532,N_6151,N_5039);
nor U6533 (N_6533,N_5987,N_5242);
nand U6534 (N_6534,N_5015,N_5569);
or U6535 (N_6535,N_5265,N_6172);
nand U6536 (N_6536,N_6050,N_5089);
nand U6537 (N_6537,N_5458,N_5970);
nor U6538 (N_6538,N_5890,N_6181);
or U6539 (N_6539,N_5579,N_5984);
nand U6540 (N_6540,N_6155,N_5747);
nor U6541 (N_6541,N_6160,N_5769);
nor U6542 (N_6542,N_5932,N_5595);
nand U6543 (N_6543,N_5147,N_5278);
nand U6544 (N_6544,N_5644,N_5049);
or U6545 (N_6545,N_5552,N_5514);
or U6546 (N_6546,N_5611,N_5978);
nor U6547 (N_6547,N_6036,N_5661);
or U6548 (N_6548,N_5568,N_6073);
or U6549 (N_6549,N_5299,N_5225);
or U6550 (N_6550,N_5939,N_6167);
and U6551 (N_6551,N_5866,N_6217);
nor U6552 (N_6552,N_5407,N_5787);
nor U6553 (N_6553,N_5832,N_5295);
nand U6554 (N_6554,N_5812,N_5722);
and U6555 (N_6555,N_5214,N_5241);
and U6556 (N_6556,N_6171,N_5754);
nand U6557 (N_6557,N_5898,N_5838);
or U6558 (N_6558,N_5174,N_5022);
and U6559 (N_6559,N_5186,N_5068);
or U6560 (N_6560,N_5171,N_5848);
nor U6561 (N_6561,N_5945,N_5372);
or U6562 (N_6562,N_5204,N_5378);
xnor U6563 (N_6563,N_5647,N_5185);
xnor U6564 (N_6564,N_5120,N_5329);
or U6565 (N_6565,N_5158,N_6218);
or U6566 (N_6566,N_5399,N_5879);
and U6567 (N_6567,N_5590,N_5677);
or U6568 (N_6568,N_5483,N_5356);
and U6569 (N_6569,N_5292,N_6008);
or U6570 (N_6570,N_5621,N_5856);
nor U6571 (N_6571,N_5258,N_6236);
and U6572 (N_6572,N_5988,N_5545);
nand U6573 (N_6573,N_5347,N_5284);
xnor U6574 (N_6574,N_5678,N_5094);
nor U6575 (N_6575,N_5967,N_5360);
nand U6576 (N_6576,N_5132,N_5316);
xor U6577 (N_6577,N_6002,N_5341);
xor U6578 (N_6578,N_5546,N_5744);
nand U6579 (N_6579,N_6207,N_6099);
and U6580 (N_6580,N_5895,N_5131);
and U6581 (N_6581,N_6021,N_5260);
xnor U6582 (N_6582,N_5909,N_5695);
nand U6583 (N_6583,N_5915,N_5064);
nand U6584 (N_6584,N_5524,N_5326);
nor U6585 (N_6585,N_5806,N_5924);
and U6586 (N_6586,N_6022,N_5408);
and U6587 (N_6587,N_5192,N_5869);
nor U6588 (N_6588,N_5485,N_6018);
xor U6589 (N_6589,N_5674,N_5422);
or U6590 (N_6590,N_5681,N_5034);
and U6591 (N_6591,N_5912,N_5062);
nand U6592 (N_6592,N_5444,N_5610);
or U6593 (N_6593,N_5921,N_5279);
nand U6594 (N_6594,N_5251,N_5853);
nand U6595 (N_6595,N_5029,N_6078);
and U6596 (N_6596,N_5577,N_5815);
and U6597 (N_6597,N_5270,N_5442);
nand U6598 (N_6598,N_5534,N_5736);
xor U6599 (N_6599,N_6009,N_5157);
and U6600 (N_6600,N_5523,N_5396);
and U6601 (N_6601,N_5486,N_5592);
and U6602 (N_6602,N_6238,N_5096);
nor U6603 (N_6603,N_5045,N_6180);
or U6604 (N_6604,N_5823,N_5465);
nand U6605 (N_6605,N_5288,N_5397);
or U6606 (N_6606,N_5786,N_5584);
xnor U6607 (N_6607,N_5009,N_5862);
nor U6608 (N_6608,N_5845,N_5966);
and U6609 (N_6609,N_5995,N_6183);
xnor U6610 (N_6610,N_5176,N_5169);
or U6611 (N_6611,N_5527,N_6056);
or U6612 (N_6612,N_5008,N_5095);
and U6613 (N_6613,N_6080,N_5016);
and U6614 (N_6614,N_5765,N_5257);
xor U6615 (N_6615,N_5785,N_5092);
or U6616 (N_6616,N_5841,N_5543);
xnor U6617 (N_6617,N_6119,N_5363);
nor U6618 (N_6618,N_6163,N_5003);
nand U6619 (N_6619,N_5842,N_5585);
nor U6620 (N_6620,N_5428,N_5540);
nand U6621 (N_6621,N_5302,N_5221);
and U6622 (N_6622,N_5344,N_5881);
xnor U6623 (N_6623,N_5510,N_5164);
xnor U6624 (N_6624,N_5080,N_5330);
nor U6625 (N_6625,N_5934,N_5919);
and U6626 (N_6626,N_6096,N_5944);
and U6627 (N_6627,N_5004,N_5404);
nand U6628 (N_6628,N_5349,N_5054);
xor U6629 (N_6629,N_5369,N_5602);
or U6630 (N_6630,N_5601,N_5495);
or U6631 (N_6631,N_5713,N_5928);
and U6632 (N_6632,N_5761,N_5692);
nand U6633 (N_6633,N_5831,N_5494);
and U6634 (N_6634,N_5658,N_5864);
or U6635 (N_6635,N_5757,N_5409);
or U6636 (N_6636,N_6017,N_5226);
nand U6637 (N_6637,N_5808,N_5400);
or U6638 (N_6638,N_5361,N_5220);
xnor U6639 (N_6639,N_5513,N_5209);
nand U6640 (N_6640,N_5972,N_5440);
or U6641 (N_6641,N_5604,N_6235);
and U6642 (N_6642,N_6013,N_6089);
or U6643 (N_6643,N_5367,N_5835);
or U6644 (N_6644,N_5730,N_5706);
nor U6645 (N_6645,N_5085,N_5771);
nor U6646 (N_6646,N_5889,N_6106);
nand U6647 (N_6647,N_5452,N_5870);
nand U6648 (N_6648,N_5025,N_5368);
and U6649 (N_6649,N_5873,N_5976);
nand U6650 (N_6650,N_5327,N_5331);
nor U6651 (N_6651,N_6130,N_6059);
and U6652 (N_6652,N_5451,N_5436);
nand U6653 (N_6653,N_5230,N_5758);
xor U6654 (N_6654,N_5259,N_5480);
xor U6655 (N_6655,N_5425,N_6113);
nor U6656 (N_6656,N_5249,N_6110);
or U6657 (N_6657,N_5603,N_6242);
nor U6658 (N_6658,N_5857,N_5114);
nor U6659 (N_6659,N_5626,N_5000);
nor U6660 (N_6660,N_5294,N_5859);
and U6661 (N_6661,N_5673,N_6162);
nor U6662 (N_6662,N_5899,N_5516);
xor U6663 (N_6663,N_6090,N_5267);
and U6664 (N_6664,N_5210,N_5810);
or U6665 (N_6665,N_5005,N_6126);
and U6666 (N_6666,N_5497,N_5291);
or U6667 (N_6667,N_5557,N_5239);
nor U6668 (N_6668,N_5466,N_5767);
nand U6669 (N_6669,N_5979,N_6100);
or U6670 (N_6670,N_5763,N_5675);
nand U6671 (N_6671,N_5748,N_6063);
nor U6672 (N_6672,N_5986,N_6200);
or U6673 (N_6673,N_5710,N_5636);
nand U6674 (N_6674,N_5854,N_5914);
and U6675 (N_6675,N_5198,N_5097);
nand U6676 (N_6676,N_5248,N_5800);
nand U6677 (N_6677,N_6157,N_5177);
and U6678 (N_6678,N_5920,N_6062);
xor U6679 (N_6679,N_5364,N_5655);
xnor U6680 (N_6680,N_6098,N_5580);
or U6681 (N_6681,N_5676,N_5087);
xnor U6682 (N_6682,N_5334,N_5975);
nand U6683 (N_6683,N_5471,N_5685);
nor U6684 (N_6684,N_5609,N_5682);
xor U6685 (N_6685,N_6042,N_5340);
xnor U6686 (N_6686,N_6239,N_5833);
and U6687 (N_6687,N_5876,N_6223);
nand U6688 (N_6688,N_5797,N_5511);
xnor U6689 (N_6689,N_5450,N_5439);
and U6690 (N_6690,N_5410,N_6142);
nand U6691 (N_6691,N_5342,N_5359);
nor U6692 (N_6692,N_5339,N_5615);
nor U6693 (N_6693,N_6158,N_6139);
and U6694 (N_6694,N_5793,N_6011);
and U6695 (N_6695,N_5830,N_5599);
xnor U6696 (N_6696,N_5843,N_5122);
or U6697 (N_6697,N_5783,N_5002);
or U6698 (N_6698,N_5118,N_6134);
nand U6699 (N_6699,N_5709,N_6023);
nand U6700 (N_6700,N_5243,N_5077);
nand U6701 (N_6701,N_5567,N_6127);
and U6702 (N_6702,N_6120,N_5276);
nor U6703 (N_6703,N_6060,N_6088);
xnor U6704 (N_6704,N_5028,N_5348);
xnor U6705 (N_6705,N_6135,N_5653);
nor U6706 (N_6706,N_5926,N_5441);
and U6707 (N_6707,N_5287,N_5193);
and U6708 (N_6708,N_5487,N_5196);
or U6709 (N_6709,N_6132,N_5043);
nor U6710 (N_6710,N_5469,N_5905);
nand U6711 (N_6711,N_6097,N_5140);
nand U6712 (N_6712,N_6103,N_5775);
nand U6713 (N_6713,N_5971,N_5774);
or U6714 (N_6714,N_5296,N_5320);
xor U6715 (N_6715,N_5227,N_6222);
xor U6716 (N_6716,N_5633,N_5778);
and U6717 (N_6717,N_5749,N_5553);
nor U6718 (N_6718,N_5708,N_5082);
nand U6719 (N_6719,N_5155,N_5729);
nor U6720 (N_6720,N_5232,N_5608);
xor U6721 (N_6721,N_6140,N_5917);
nor U6722 (N_6722,N_5388,N_5727);
nand U6723 (N_6723,N_5643,N_5941);
nor U6724 (N_6724,N_5902,N_5290);
xnor U6725 (N_6725,N_5151,N_5134);
xnor U6726 (N_6726,N_5071,N_5021);
nand U6727 (N_6727,N_5217,N_6245);
or U6728 (N_6728,N_5627,N_5936);
nand U6729 (N_6729,N_5350,N_5416);
xor U6730 (N_6730,N_5885,N_5952);
or U6731 (N_6731,N_5663,N_5366);
or U6732 (N_6732,N_5712,N_6197);
xor U6733 (N_6733,N_5182,N_6092);
xnor U6734 (N_6734,N_6240,N_5057);
nand U6735 (N_6735,N_6025,N_5600);
or U6736 (N_6736,N_5743,N_5820);
nor U6737 (N_6737,N_5731,N_5228);
nor U6738 (N_6738,N_5718,N_5639);
or U6739 (N_6739,N_5631,N_6019);
and U6740 (N_6740,N_5884,N_5735);
xor U6741 (N_6741,N_5847,N_5351);
and U6742 (N_6742,N_5525,N_5268);
nor U6743 (N_6743,N_5994,N_5738);
or U6744 (N_6744,N_5519,N_5755);
nand U6745 (N_6745,N_6244,N_6104);
or U6746 (N_6746,N_5961,N_5271);
nor U6747 (N_6747,N_5283,N_5947);
xnor U6748 (N_6748,N_5803,N_5992);
nor U6749 (N_6749,N_5314,N_5720);
and U6750 (N_6750,N_5484,N_6156);
nand U6751 (N_6751,N_5137,N_5402);
and U6752 (N_6752,N_5867,N_5874);
nor U6753 (N_6753,N_5696,N_5001);
xor U6754 (N_6754,N_5846,N_5931);
nor U6755 (N_6755,N_5887,N_5179);
xnor U6756 (N_6756,N_5381,N_6224);
nand U6757 (N_6757,N_5993,N_5050);
or U6758 (N_6758,N_5646,N_5989);
nand U6759 (N_6759,N_6187,N_6211);
nor U6760 (N_6760,N_5576,N_5549);
nand U6761 (N_6761,N_5229,N_6184);
xor U6762 (N_6762,N_5798,N_5453);
nand U6763 (N_6763,N_6214,N_5067);
xnor U6764 (N_6764,N_5892,N_5463);
nor U6765 (N_6765,N_6148,N_5883);
nand U6766 (N_6766,N_5855,N_5746);
and U6767 (N_6767,N_5725,N_6077);
nand U6768 (N_6768,N_5240,N_5362);
nand U6769 (N_6769,N_5742,N_6129);
xor U6770 (N_6770,N_6208,N_6048);
and U6771 (N_6771,N_5424,N_5017);
nor U6772 (N_6772,N_5651,N_5871);
nand U6773 (N_6773,N_5922,N_6001);
and U6774 (N_6774,N_5780,N_5817);
or U6775 (N_6775,N_5195,N_5414);
xor U6776 (N_6776,N_5648,N_5588);
and U6777 (N_6777,N_5606,N_6170);
or U6778 (N_6778,N_6066,N_5923);
and U6779 (N_6779,N_5539,N_5245);
or U6780 (N_6780,N_6029,N_6229);
nor U6781 (N_6781,N_5112,N_6182);
nand U6782 (N_6782,N_5699,N_6230);
or U6783 (N_6783,N_5741,N_5776);
and U6784 (N_6784,N_5148,N_5554);
or U6785 (N_6785,N_5063,N_5219);
nor U6786 (N_6786,N_5943,N_5702);
xnor U6787 (N_6787,N_6149,N_5770);
and U6788 (N_6788,N_5098,N_5401);
or U6789 (N_6789,N_5144,N_6216);
and U6790 (N_6790,N_5386,N_5406);
and U6791 (N_6791,N_6121,N_6179);
xor U6792 (N_6792,N_5529,N_5764);
or U6793 (N_6793,N_5891,N_5138);
xor U6794 (N_6794,N_5311,N_5405);
nor U6795 (N_6795,N_5538,N_6220);
or U6796 (N_6796,N_5635,N_6046);
and U6797 (N_6797,N_5304,N_5723);
nand U6798 (N_6798,N_6168,N_6061);
nor U6799 (N_6799,N_6174,N_5149);
nor U6800 (N_6800,N_5596,N_5108);
nand U6801 (N_6801,N_5802,N_5066);
or U6802 (N_6802,N_5285,N_6076);
nand U6803 (N_6803,N_5836,N_5354);
and U6804 (N_6804,N_5768,N_6191);
or U6805 (N_6805,N_5150,N_6112);
xor U6806 (N_6806,N_6164,N_5623);
xor U6807 (N_6807,N_6033,N_5840);
and U6808 (N_6808,N_6185,N_5790);
xor U6809 (N_6809,N_5328,N_5492);
or U6810 (N_6810,N_5849,N_5024);
nor U6811 (N_6811,N_5306,N_5037);
nand U6812 (N_6812,N_5435,N_5784);
and U6813 (N_6813,N_5412,N_5937);
and U6814 (N_6814,N_5688,N_5503);
and U6815 (N_6815,N_5965,N_5760);
and U6816 (N_6816,N_5254,N_5411);
nand U6817 (N_6817,N_6233,N_5026);
nor U6818 (N_6818,N_6043,N_6012);
xor U6819 (N_6819,N_5218,N_5660);
nand U6820 (N_6820,N_5222,N_5907);
and U6821 (N_6821,N_6026,N_5200);
or U6822 (N_6822,N_6186,N_5212);
xor U6823 (N_6823,N_5637,N_6159);
nand U6824 (N_6824,N_5333,N_5773);
or U6825 (N_6825,N_6058,N_5981);
and U6826 (N_6826,N_5091,N_5619);
xor U6827 (N_6827,N_6068,N_5065);
xor U6828 (N_6828,N_5837,N_5948);
nand U6829 (N_6829,N_5693,N_5393);
or U6830 (N_6830,N_5814,N_6201);
or U6831 (N_6831,N_5759,N_5309);
or U6832 (N_6832,N_5083,N_6153);
xnor U6833 (N_6833,N_5886,N_5136);
xor U6834 (N_6834,N_5852,N_5070);
nand U6835 (N_6835,N_5335,N_6070);
or U6836 (N_6836,N_5974,N_5449);
or U6837 (N_6837,N_5421,N_5680);
and U6838 (N_6838,N_5719,N_5030);
or U6839 (N_6839,N_6116,N_5813);
and U6840 (N_6840,N_6074,N_5998);
or U6841 (N_6841,N_6064,N_5620);
nor U6842 (N_6842,N_5570,N_5427);
xnor U6843 (N_6843,N_5536,N_5888);
xor U6844 (N_6844,N_6195,N_5811);
and U6845 (N_6845,N_5365,N_5985);
nor U6846 (N_6846,N_5860,N_5154);
nor U6847 (N_6847,N_5528,N_5459);
and U6848 (N_6848,N_5447,N_5690);
nor U6849 (N_6849,N_5454,N_5893);
or U6850 (N_6850,N_5762,N_5612);
xnor U6851 (N_6851,N_5605,N_5589);
or U6852 (N_6852,N_5996,N_5645);
or U6853 (N_6853,N_5324,N_5819);
or U6854 (N_6854,N_6196,N_6108);
nor U6855 (N_6855,N_6094,N_6016);
nand U6856 (N_6856,N_5456,N_5634);
xor U6857 (N_6857,N_5991,N_5312);
nand U6858 (N_6858,N_6114,N_6231);
and U6859 (N_6859,N_5607,N_5310);
nor U6860 (N_6860,N_6115,N_6137);
and U6861 (N_6861,N_5508,N_5478);
or U6862 (N_6862,N_6237,N_5927);
and U6863 (N_6863,N_5799,N_5036);
nand U6864 (N_6864,N_5687,N_5824);
or U6865 (N_6865,N_6178,N_5110);
and U6866 (N_6866,N_5479,N_5117);
nor U6867 (N_6867,N_5300,N_5613);
or U6868 (N_6868,N_5664,N_5668);
or U6869 (N_6869,N_5078,N_5789);
or U6870 (N_6870,N_6065,N_5153);
xnor U6871 (N_6871,N_6165,N_5489);
xor U6872 (N_6872,N_5231,N_5392);
nor U6873 (N_6873,N_6044,N_5358);
or U6874 (N_6874,N_5332,N_6031);
nand U6875 (N_6875,N_5529,N_5397);
and U6876 (N_6876,N_5699,N_5297);
nand U6877 (N_6877,N_5121,N_5930);
or U6878 (N_6878,N_5145,N_5122);
and U6879 (N_6879,N_6117,N_5382);
xor U6880 (N_6880,N_6053,N_5735);
nor U6881 (N_6881,N_5754,N_5663);
xor U6882 (N_6882,N_5614,N_6071);
and U6883 (N_6883,N_5443,N_5576);
or U6884 (N_6884,N_5081,N_5806);
or U6885 (N_6885,N_5739,N_5134);
xnor U6886 (N_6886,N_5047,N_5315);
nor U6887 (N_6887,N_5806,N_5743);
or U6888 (N_6888,N_6090,N_5595);
nor U6889 (N_6889,N_5535,N_6175);
nand U6890 (N_6890,N_5850,N_6073);
xnor U6891 (N_6891,N_5624,N_6014);
or U6892 (N_6892,N_5732,N_6048);
nor U6893 (N_6893,N_5947,N_5275);
or U6894 (N_6894,N_5716,N_6231);
and U6895 (N_6895,N_5709,N_5613);
xnor U6896 (N_6896,N_5870,N_5383);
and U6897 (N_6897,N_5029,N_6022);
nand U6898 (N_6898,N_6006,N_5100);
nor U6899 (N_6899,N_5512,N_5575);
or U6900 (N_6900,N_5265,N_5383);
nand U6901 (N_6901,N_5689,N_6018);
xor U6902 (N_6902,N_6102,N_5359);
and U6903 (N_6903,N_5058,N_6183);
and U6904 (N_6904,N_6169,N_5084);
nand U6905 (N_6905,N_5441,N_5603);
xor U6906 (N_6906,N_5854,N_5262);
xnor U6907 (N_6907,N_6030,N_5004);
nor U6908 (N_6908,N_5632,N_5060);
nand U6909 (N_6909,N_5483,N_5163);
nand U6910 (N_6910,N_5938,N_5227);
nor U6911 (N_6911,N_5186,N_6018);
nor U6912 (N_6912,N_6003,N_5155);
nand U6913 (N_6913,N_5326,N_5102);
xor U6914 (N_6914,N_5653,N_5740);
xnor U6915 (N_6915,N_5229,N_5874);
nand U6916 (N_6916,N_5602,N_5165);
and U6917 (N_6917,N_5345,N_5030);
or U6918 (N_6918,N_5330,N_5404);
nor U6919 (N_6919,N_5151,N_5947);
nand U6920 (N_6920,N_5577,N_5420);
nor U6921 (N_6921,N_5969,N_5319);
nor U6922 (N_6922,N_6247,N_5862);
and U6923 (N_6923,N_5903,N_5200);
or U6924 (N_6924,N_5916,N_5653);
and U6925 (N_6925,N_5878,N_5271);
nand U6926 (N_6926,N_6156,N_5553);
nand U6927 (N_6927,N_5624,N_5302);
or U6928 (N_6928,N_6070,N_5606);
and U6929 (N_6929,N_5654,N_5512);
nand U6930 (N_6930,N_5140,N_5779);
or U6931 (N_6931,N_5612,N_5275);
xor U6932 (N_6932,N_6230,N_5581);
xor U6933 (N_6933,N_5563,N_5143);
and U6934 (N_6934,N_5359,N_5126);
xnor U6935 (N_6935,N_5901,N_5204);
nand U6936 (N_6936,N_5102,N_6094);
xnor U6937 (N_6937,N_5161,N_6049);
or U6938 (N_6938,N_6219,N_5955);
or U6939 (N_6939,N_6060,N_5716);
nor U6940 (N_6940,N_5416,N_6235);
nand U6941 (N_6941,N_6089,N_5231);
nor U6942 (N_6942,N_5565,N_5535);
xnor U6943 (N_6943,N_5164,N_5524);
or U6944 (N_6944,N_6134,N_5662);
or U6945 (N_6945,N_5678,N_5211);
nand U6946 (N_6946,N_5967,N_5328);
nand U6947 (N_6947,N_5824,N_5636);
and U6948 (N_6948,N_5349,N_5972);
nand U6949 (N_6949,N_5876,N_6103);
nand U6950 (N_6950,N_5183,N_6138);
nor U6951 (N_6951,N_5248,N_5941);
nand U6952 (N_6952,N_5678,N_5099);
or U6953 (N_6953,N_5814,N_5044);
or U6954 (N_6954,N_5022,N_5498);
and U6955 (N_6955,N_5150,N_5315);
xor U6956 (N_6956,N_5900,N_5419);
nor U6957 (N_6957,N_5600,N_5952);
xnor U6958 (N_6958,N_6112,N_5531);
and U6959 (N_6959,N_5074,N_5364);
xnor U6960 (N_6960,N_6241,N_5918);
nand U6961 (N_6961,N_6203,N_5927);
or U6962 (N_6962,N_5462,N_5846);
nor U6963 (N_6963,N_6188,N_6235);
nand U6964 (N_6964,N_5273,N_5715);
nor U6965 (N_6965,N_5276,N_5292);
nand U6966 (N_6966,N_5779,N_5415);
or U6967 (N_6967,N_5964,N_5367);
or U6968 (N_6968,N_5487,N_5756);
and U6969 (N_6969,N_6012,N_5315);
xnor U6970 (N_6970,N_5160,N_5247);
xnor U6971 (N_6971,N_5907,N_5932);
or U6972 (N_6972,N_6184,N_5812);
and U6973 (N_6973,N_5799,N_5090);
xnor U6974 (N_6974,N_5267,N_5768);
or U6975 (N_6975,N_5568,N_6225);
xor U6976 (N_6976,N_6179,N_5188);
nor U6977 (N_6977,N_5288,N_5302);
or U6978 (N_6978,N_5873,N_5102);
xnor U6979 (N_6979,N_5892,N_5880);
and U6980 (N_6980,N_5382,N_5316);
nor U6981 (N_6981,N_5250,N_5314);
nand U6982 (N_6982,N_5555,N_5997);
or U6983 (N_6983,N_5396,N_5633);
nor U6984 (N_6984,N_5518,N_6212);
nand U6985 (N_6985,N_5981,N_5615);
xnor U6986 (N_6986,N_5497,N_5117);
nand U6987 (N_6987,N_6045,N_5669);
nand U6988 (N_6988,N_5753,N_5755);
nand U6989 (N_6989,N_5893,N_5400);
nor U6990 (N_6990,N_5602,N_5848);
or U6991 (N_6991,N_5815,N_5135);
and U6992 (N_6992,N_6029,N_5359);
xnor U6993 (N_6993,N_5243,N_6055);
and U6994 (N_6994,N_6243,N_5724);
and U6995 (N_6995,N_6182,N_5991);
or U6996 (N_6996,N_5685,N_5275);
nor U6997 (N_6997,N_5201,N_5351);
nand U6998 (N_6998,N_5258,N_5308);
or U6999 (N_6999,N_5313,N_5903);
nor U7000 (N_7000,N_5549,N_6094);
and U7001 (N_7001,N_5917,N_6091);
or U7002 (N_7002,N_5063,N_5166);
nor U7003 (N_7003,N_5568,N_6015);
nor U7004 (N_7004,N_6111,N_5786);
xnor U7005 (N_7005,N_5997,N_5885);
xor U7006 (N_7006,N_6089,N_6164);
nand U7007 (N_7007,N_5446,N_5626);
nand U7008 (N_7008,N_6012,N_5241);
nor U7009 (N_7009,N_5983,N_5319);
nand U7010 (N_7010,N_5077,N_5994);
nand U7011 (N_7011,N_5260,N_5634);
or U7012 (N_7012,N_5809,N_6204);
or U7013 (N_7013,N_6188,N_5160);
and U7014 (N_7014,N_5984,N_5003);
or U7015 (N_7015,N_5642,N_5313);
and U7016 (N_7016,N_5356,N_5655);
nand U7017 (N_7017,N_5622,N_5557);
nand U7018 (N_7018,N_5895,N_5856);
xnor U7019 (N_7019,N_5032,N_5945);
xor U7020 (N_7020,N_5325,N_5716);
and U7021 (N_7021,N_5670,N_5863);
or U7022 (N_7022,N_5063,N_6243);
and U7023 (N_7023,N_5185,N_5260);
xnor U7024 (N_7024,N_5512,N_5091);
nor U7025 (N_7025,N_5750,N_5463);
nand U7026 (N_7026,N_5670,N_5106);
nand U7027 (N_7027,N_6033,N_5278);
nand U7028 (N_7028,N_5456,N_5405);
nor U7029 (N_7029,N_5581,N_5622);
xnor U7030 (N_7030,N_5452,N_5511);
and U7031 (N_7031,N_5001,N_6228);
nor U7032 (N_7032,N_6143,N_5502);
and U7033 (N_7033,N_6090,N_5766);
or U7034 (N_7034,N_5119,N_5609);
nand U7035 (N_7035,N_5317,N_5868);
xnor U7036 (N_7036,N_6234,N_5600);
xnor U7037 (N_7037,N_5868,N_5004);
xor U7038 (N_7038,N_5867,N_6020);
nor U7039 (N_7039,N_5190,N_5716);
nor U7040 (N_7040,N_5674,N_6008);
nor U7041 (N_7041,N_5619,N_6006);
nor U7042 (N_7042,N_5355,N_5049);
nand U7043 (N_7043,N_6073,N_5088);
or U7044 (N_7044,N_6122,N_5226);
nor U7045 (N_7045,N_5896,N_5026);
nor U7046 (N_7046,N_5747,N_6238);
nand U7047 (N_7047,N_5088,N_5320);
or U7048 (N_7048,N_5993,N_5708);
nand U7049 (N_7049,N_6016,N_5944);
nor U7050 (N_7050,N_5807,N_5236);
xnor U7051 (N_7051,N_5344,N_5323);
nor U7052 (N_7052,N_5464,N_5242);
or U7053 (N_7053,N_6020,N_6001);
xnor U7054 (N_7054,N_5346,N_6012);
xnor U7055 (N_7055,N_5354,N_5582);
and U7056 (N_7056,N_5476,N_5229);
nor U7057 (N_7057,N_5566,N_5635);
nand U7058 (N_7058,N_5972,N_5011);
and U7059 (N_7059,N_5389,N_5643);
or U7060 (N_7060,N_5619,N_6241);
and U7061 (N_7061,N_5261,N_5279);
and U7062 (N_7062,N_5890,N_5029);
nand U7063 (N_7063,N_6192,N_5202);
and U7064 (N_7064,N_5612,N_6117);
nor U7065 (N_7065,N_5425,N_5275);
xnor U7066 (N_7066,N_5069,N_5542);
and U7067 (N_7067,N_5410,N_6005);
or U7068 (N_7068,N_5231,N_5741);
nor U7069 (N_7069,N_5013,N_5119);
xor U7070 (N_7070,N_5606,N_5055);
xnor U7071 (N_7071,N_5881,N_6219);
or U7072 (N_7072,N_5741,N_5396);
nand U7073 (N_7073,N_6072,N_5606);
xnor U7074 (N_7074,N_6104,N_5443);
xnor U7075 (N_7075,N_5122,N_6130);
nor U7076 (N_7076,N_5020,N_5173);
and U7077 (N_7077,N_5574,N_5653);
nand U7078 (N_7078,N_5712,N_5496);
nand U7079 (N_7079,N_5078,N_6239);
and U7080 (N_7080,N_5859,N_5190);
nor U7081 (N_7081,N_5711,N_5257);
and U7082 (N_7082,N_6035,N_5010);
nand U7083 (N_7083,N_5656,N_5825);
and U7084 (N_7084,N_5512,N_5146);
or U7085 (N_7085,N_5592,N_5757);
or U7086 (N_7086,N_6085,N_5788);
and U7087 (N_7087,N_5258,N_6132);
and U7088 (N_7088,N_5060,N_5497);
and U7089 (N_7089,N_5502,N_5724);
and U7090 (N_7090,N_6120,N_6140);
and U7091 (N_7091,N_5857,N_5029);
nand U7092 (N_7092,N_5928,N_5204);
and U7093 (N_7093,N_5911,N_6062);
xnor U7094 (N_7094,N_5712,N_5898);
nor U7095 (N_7095,N_5638,N_5648);
xor U7096 (N_7096,N_5876,N_5673);
nor U7097 (N_7097,N_6042,N_6245);
nor U7098 (N_7098,N_5519,N_5917);
nand U7099 (N_7099,N_5791,N_5877);
nand U7100 (N_7100,N_5849,N_5704);
nor U7101 (N_7101,N_5889,N_5962);
xor U7102 (N_7102,N_6009,N_6008);
or U7103 (N_7103,N_5948,N_5993);
or U7104 (N_7104,N_5130,N_5214);
xnor U7105 (N_7105,N_5179,N_5306);
xor U7106 (N_7106,N_5887,N_6144);
nor U7107 (N_7107,N_6077,N_5928);
and U7108 (N_7108,N_5312,N_5397);
and U7109 (N_7109,N_5698,N_5536);
and U7110 (N_7110,N_6188,N_5242);
nor U7111 (N_7111,N_6074,N_5352);
and U7112 (N_7112,N_5212,N_5363);
and U7113 (N_7113,N_5719,N_5176);
or U7114 (N_7114,N_5061,N_5923);
and U7115 (N_7115,N_5964,N_6144);
nand U7116 (N_7116,N_5477,N_5005);
nand U7117 (N_7117,N_6074,N_5325);
and U7118 (N_7118,N_6060,N_5424);
and U7119 (N_7119,N_5509,N_5889);
or U7120 (N_7120,N_5603,N_5986);
nand U7121 (N_7121,N_5196,N_6088);
nor U7122 (N_7122,N_5792,N_5590);
nor U7123 (N_7123,N_6160,N_5536);
and U7124 (N_7124,N_5223,N_5698);
xor U7125 (N_7125,N_5414,N_5029);
and U7126 (N_7126,N_5787,N_5602);
nor U7127 (N_7127,N_5044,N_5889);
nand U7128 (N_7128,N_5105,N_6078);
nor U7129 (N_7129,N_5614,N_5351);
and U7130 (N_7130,N_5022,N_5659);
or U7131 (N_7131,N_5789,N_5454);
xor U7132 (N_7132,N_5416,N_5965);
or U7133 (N_7133,N_6248,N_6219);
and U7134 (N_7134,N_6125,N_5203);
or U7135 (N_7135,N_5210,N_6148);
and U7136 (N_7136,N_5579,N_6198);
or U7137 (N_7137,N_5815,N_5589);
and U7138 (N_7138,N_5265,N_5650);
nand U7139 (N_7139,N_5561,N_5865);
and U7140 (N_7140,N_5897,N_5154);
xnor U7141 (N_7141,N_5121,N_5856);
nand U7142 (N_7142,N_5052,N_5213);
nor U7143 (N_7143,N_5631,N_5643);
nand U7144 (N_7144,N_5873,N_5938);
and U7145 (N_7145,N_6139,N_5007);
nor U7146 (N_7146,N_5703,N_5546);
xor U7147 (N_7147,N_5277,N_5968);
xor U7148 (N_7148,N_5566,N_5877);
xor U7149 (N_7149,N_5189,N_5108);
xnor U7150 (N_7150,N_5432,N_5298);
and U7151 (N_7151,N_6035,N_5535);
or U7152 (N_7152,N_5409,N_5077);
nor U7153 (N_7153,N_5030,N_5737);
or U7154 (N_7154,N_5219,N_5501);
or U7155 (N_7155,N_5625,N_5794);
and U7156 (N_7156,N_6185,N_6195);
or U7157 (N_7157,N_5857,N_5147);
nand U7158 (N_7158,N_5761,N_5249);
nor U7159 (N_7159,N_5387,N_5501);
nor U7160 (N_7160,N_5407,N_6223);
nor U7161 (N_7161,N_5649,N_5141);
or U7162 (N_7162,N_5425,N_5069);
xnor U7163 (N_7163,N_5063,N_5179);
nand U7164 (N_7164,N_5438,N_5666);
and U7165 (N_7165,N_6200,N_5583);
and U7166 (N_7166,N_5461,N_5814);
and U7167 (N_7167,N_6131,N_5766);
or U7168 (N_7168,N_5161,N_5261);
nand U7169 (N_7169,N_5987,N_5860);
and U7170 (N_7170,N_5271,N_5514);
xor U7171 (N_7171,N_5572,N_5668);
or U7172 (N_7172,N_5894,N_5645);
nand U7173 (N_7173,N_5076,N_6158);
nor U7174 (N_7174,N_5342,N_6098);
or U7175 (N_7175,N_5629,N_5856);
or U7176 (N_7176,N_5297,N_5844);
nor U7177 (N_7177,N_5519,N_5089);
nand U7178 (N_7178,N_5854,N_5794);
nand U7179 (N_7179,N_6194,N_5821);
nand U7180 (N_7180,N_5130,N_5965);
or U7181 (N_7181,N_5901,N_6105);
nor U7182 (N_7182,N_5089,N_5999);
nor U7183 (N_7183,N_5870,N_5744);
nand U7184 (N_7184,N_5999,N_5133);
nand U7185 (N_7185,N_5725,N_5193);
nand U7186 (N_7186,N_5802,N_6141);
nor U7187 (N_7187,N_6087,N_5538);
xnor U7188 (N_7188,N_5067,N_5611);
and U7189 (N_7189,N_5664,N_5684);
nor U7190 (N_7190,N_6092,N_6108);
nand U7191 (N_7191,N_6201,N_5737);
nand U7192 (N_7192,N_5120,N_5537);
nand U7193 (N_7193,N_5513,N_5002);
and U7194 (N_7194,N_5525,N_5732);
nand U7195 (N_7195,N_5489,N_6102);
or U7196 (N_7196,N_5615,N_5516);
or U7197 (N_7197,N_5986,N_5968);
xnor U7198 (N_7198,N_6007,N_5548);
nand U7199 (N_7199,N_5437,N_5506);
xnor U7200 (N_7200,N_5654,N_5341);
xor U7201 (N_7201,N_6179,N_5385);
or U7202 (N_7202,N_6025,N_5321);
and U7203 (N_7203,N_5446,N_6114);
and U7204 (N_7204,N_5996,N_5288);
nand U7205 (N_7205,N_5941,N_5704);
xor U7206 (N_7206,N_5006,N_5269);
nand U7207 (N_7207,N_6157,N_5891);
nor U7208 (N_7208,N_5972,N_5351);
xor U7209 (N_7209,N_6083,N_5746);
xnor U7210 (N_7210,N_5453,N_6105);
xor U7211 (N_7211,N_5997,N_5563);
xnor U7212 (N_7212,N_6189,N_6092);
nor U7213 (N_7213,N_5622,N_5133);
and U7214 (N_7214,N_6037,N_5310);
nor U7215 (N_7215,N_5093,N_5432);
xor U7216 (N_7216,N_5979,N_6210);
xor U7217 (N_7217,N_6106,N_5461);
xnor U7218 (N_7218,N_6159,N_5860);
nand U7219 (N_7219,N_6159,N_6120);
and U7220 (N_7220,N_5338,N_5193);
nand U7221 (N_7221,N_6070,N_5561);
or U7222 (N_7222,N_5020,N_5548);
and U7223 (N_7223,N_5722,N_5011);
nand U7224 (N_7224,N_6169,N_5431);
nor U7225 (N_7225,N_5588,N_5493);
or U7226 (N_7226,N_6031,N_5000);
nand U7227 (N_7227,N_5985,N_5729);
xnor U7228 (N_7228,N_5016,N_5493);
xor U7229 (N_7229,N_6174,N_6089);
or U7230 (N_7230,N_6059,N_5323);
and U7231 (N_7231,N_5336,N_6119);
nor U7232 (N_7232,N_6206,N_6249);
and U7233 (N_7233,N_5260,N_5728);
xor U7234 (N_7234,N_5624,N_5362);
or U7235 (N_7235,N_5787,N_6123);
nand U7236 (N_7236,N_5380,N_5095);
nand U7237 (N_7237,N_6178,N_5247);
or U7238 (N_7238,N_6152,N_5744);
xor U7239 (N_7239,N_5579,N_5629);
and U7240 (N_7240,N_5812,N_5467);
or U7241 (N_7241,N_5138,N_5160);
or U7242 (N_7242,N_5056,N_5421);
and U7243 (N_7243,N_5025,N_5002);
nand U7244 (N_7244,N_5026,N_5800);
nand U7245 (N_7245,N_5931,N_5370);
and U7246 (N_7246,N_5144,N_5618);
xnor U7247 (N_7247,N_5979,N_6038);
xnor U7248 (N_7248,N_6229,N_5638);
or U7249 (N_7249,N_5063,N_6175);
and U7250 (N_7250,N_5475,N_5177);
or U7251 (N_7251,N_5433,N_6224);
xnor U7252 (N_7252,N_5150,N_5577);
nand U7253 (N_7253,N_5605,N_5397);
xor U7254 (N_7254,N_5614,N_5665);
nor U7255 (N_7255,N_5803,N_5106);
and U7256 (N_7256,N_5229,N_5834);
xor U7257 (N_7257,N_5825,N_5548);
nor U7258 (N_7258,N_6030,N_5750);
or U7259 (N_7259,N_5976,N_5999);
nand U7260 (N_7260,N_5157,N_5854);
or U7261 (N_7261,N_6127,N_5188);
or U7262 (N_7262,N_5390,N_5349);
and U7263 (N_7263,N_5320,N_5130);
nor U7264 (N_7264,N_6039,N_5252);
xor U7265 (N_7265,N_5610,N_5945);
and U7266 (N_7266,N_6133,N_5329);
nor U7267 (N_7267,N_5485,N_5082);
or U7268 (N_7268,N_6154,N_5110);
nand U7269 (N_7269,N_5908,N_6236);
nand U7270 (N_7270,N_5117,N_5741);
nor U7271 (N_7271,N_5610,N_6232);
or U7272 (N_7272,N_5378,N_6000);
or U7273 (N_7273,N_5853,N_5392);
nor U7274 (N_7274,N_5658,N_5081);
xnor U7275 (N_7275,N_6012,N_5238);
xor U7276 (N_7276,N_5119,N_5931);
nand U7277 (N_7277,N_5344,N_5090);
nor U7278 (N_7278,N_5154,N_5582);
nor U7279 (N_7279,N_5130,N_6105);
and U7280 (N_7280,N_6048,N_5860);
nor U7281 (N_7281,N_5943,N_5868);
and U7282 (N_7282,N_5924,N_6038);
nor U7283 (N_7283,N_6009,N_6204);
nand U7284 (N_7284,N_5249,N_6137);
nor U7285 (N_7285,N_5070,N_5318);
nand U7286 (N_7286,N_6201,N_5830);
nand U7287 (N_7287,N_5961,N_5228);
nor U7288 (N_7288,N_5027,N_6048);
nor U7289 (N_7289,N_5584,N_5516);
and U7290 (N_7290,N_5134,N_5061);
nor U7291 (N_7291,N_5608,N_5923);
and U7292 (N_7292,N_6235,N_6161);
and U7293 (N_7293,N_6034,N_5627);
nand U7294 (N_7294,N_6093,N_5787);
nor U7295 (N_7295,N_5601,N_5563);
and U7296 (N_7296,N_5591,N_6216);
nor U7297 (N_7297,N_5888,N_5959);
and U7298 (N_7298,N_5623,N_5699);
and U7299 (N_7299,N_6166,N_5319);
nor U7300 (N_7300,N_5180,N_5052);
nand U7301 (N_7301,N_5706,N_5828);
and U7302 (N_7302,N_5458,N_5951);
nor U7303 (N_7303,N_5623,N_5229);
nor U7304 (N_7304,N_5835,N_5651);
or U7305 (N_7305,N_5749,N_5900);
nand U7306 (N_7306,N_5079,N_5088);
xor U7307 (N_7307,N_5849,N_5753);
or U7308 (N_7308,N_5855,N_5231);
xnor U7309 (N_7309,N_5728,N_5359);
nand U7310 (N_7310,N_6172,N_6171);
and U7311 (N_7311,N_5982,N_6163);
and U7312 (N_7312,N_5861,N_5535);
and U7313 (N_7313,N_5978,N_6152);
and U7314 (N_7314,N_5289,N_5551);
xor U7315 (N_7315,N_5176,N_5453);
or U7316 (N_7316,N_5906,N_6104);
xnor U7317 (N_7317,N_6215,N_5612);
and U7318 (N_7318,N_6238,N_5988);
and U7319 (N_7319,N_5441,N_5670);
and U7320 (N_7320,N_6236,N_5157);
xnor U7321 (N_7321,N_5193,N_6013);
nand U7322 (N_7322,N_5811,N_5247);
or U7323 (N_7323,N_5799,N_5592);
or U7324 (N_7324,N_5352,N_5186);
nand U7325 (N_7325,N_5816,N_6132);
nand U7326 (N_7326,N_5824,N_5311);
nor U7327 (N_7327,N_5701,N_5918);
and U7328 (N_7328,N_5770,N_6043);
nand U7329 (N_7329,N_5874,N_5187);
and U7330 (N_7330,N_5618,N_5218);
or U7331 (N_7331,N_5447,N_6140);
nor U7332 (N_7332,N_5135,N_5655);
nor U7333 (N_7333,N_5077,N_5272);
nor U7334 (N_7334,N_5135,N_6138);
xor U7335 (N_7335,N_5701,N_6112);
xor U7336 (N_7336,N_5885,N_5959);
nand U7337 (N_7337,N_5614,N_6060);
and U7338 (N_7338,N_5293,N_5682);
or U7339 (N_7339,N_6105,N_5180);
nor U7340 (N_7340,N_6086,N_5076);
nor U7341 (N_7341,N_6176,N_5662);
nand U7342 (N_7342,N_5639,N_5662);
nor U7343 (N_7343,N_6025,N_5361);
and U7344 (N_7344,N_6215,N_6050);
or U7345 (N_7345,N_5797,N_5920);
nor U7346 (N_7346,N_5508,N_5868);
nand U7347 (N_7347,N_5370,N_5036);
or U7348 (N_7348,N_5936,N_5647);
nand U7349 (N_7349,N_5706,N_5908);
nand U7350 (N_7350,N_5560,N_5664);
or U7351 (N_7351,N_6133,N_5944);
and U7352 (N_7352,N_5597,N_5545);
nor U7353 (N_7353,N_6150,N_5196);
or U7354 (N_7354,N_5706,N_5729);
or U7355 (N_7355,N_5693,N_5163);
and U7356 (N_7356,N_6090,N_5204);
nor U7357 (N_7357,N_5479,N_5486);
and U7358 (N_7358,N_5347,N_5916);
nand U7359 (N_7359,N_5674,N_5339);
nor U7360 (N_7360,N_5566,N_6023);
nor U7361 (N_7361,N_5511,N_5831);
or U7362 (N_7362,N_5350,N_6202);
nand U7363 (N_7363,N_5347,N_5843);
xor U7364 (N_7364,N_5257,N_5532);
xor U7365 (N_7365,N_5408,N_6194);
or U7366 (N_7366,N_6183,N_5446);
nor U7367 (N_7367,N_5016,N_5961);
nand U7368 (N_7368,N_5456,N_5166);
xor U7369 (N_7369,N_5626,N_6153);
xor U7370 (N_7370,N_5140,N_6039);
nand U7371 (N_7371,N_5243,N_5822);
and U7372 (N_7372,N_5866,N_6030);
nor U7373 (N_7373,N_5073,N_5642);
or U7374 (N_7374,N_5758,N_5685);
and U7375 (N_7375,N_5908,N_5959);
nor U7376 (N_7376,N_5526,N_5713);
and U7377 (N_7377,N_5870,N_5038);
nor U7378 (N_7378,N_5957,N_6241);
nor U7379 (N_7379,N_5915,N_5215);
xor U7380 (N_7380,N_5171,N_5798);
xnor U7381 (N_7381,N_6233,N_5018);
and U7382 (N_7382,N_5332,N_5257);
or U7383 (N_7383,N_5844,N_5528);
or U7384 (N_7384,N_5811,N_5329);
xnor U7385 (N_7385,N_5006,N_5147);
and U7386 (N_7386,N_5204,N_5241);
xnor U7387 (N_7387,N_5386,N_5311);
xor U7388 (N_7388,N_5844,N_5283);
and U7389 (N_7389,N_5664,N_5786);
nand U7390 (N_7390,N_6182,N_5748);
xnor U7391 (N_7391,N_5184,N_5459);
or U7392 (N_7392,N_5174,N_5865);
nor U7393 (N_7393,N_5486,N_6224);
and U7394 (N_7394,N_5045,N_5617);
xor U7395 (N_7395,N_6201,N_6099);
nor U7396 (N_7396,N_5646,N_5011);
or U7397 (N_7397,N_6072,N_5358);
xor U7398 (N_7398,N_5863,N_5184);
nor U7399 (N_7399,N_5011,N_5850);
nor U7400 (N_7400,N_5609,N_6165);
nor U7401 (N_7401,N_5630,N_6098);
and U7402 (N_7402,N_5271,N_6026);
nor U7403 (N_7403,N_5225,N_5924);
or U7404 (N_7404,N_5060,N_5935);
nor U7405 (N_7405,N_6215,N_5608);
nand U7406 (N_7406,N_6016,N_5356);
and U7407 (N_7407,N_5738,N_5204);
and U7408 (N_7408,N_6045,N_5236);
nand U7409 (N_7409,N_6194,N_5540);
nand U7410 (N_7410,N_5872,N_5371);
xnor U7411 (N_7411,N_5285,N_5935);
nand U7412 (N_7412,N_5569,N_6201);
nor U7413 (N_7413,N_6017,N_6193);
and U7414 (N_7414,N_5409,N_5046);
and U7415 (N_7415,N_5077,N_5804);
or U7416 (N_7416,N_5232,N_5078);
nor U7417 (N_7417,N_5457,N_5769);
or U7418 (N_7418,N_5622,N_6228);
nand U7419 (N_7419,N_5962,N_5270);
xnor U7420 (N_7420,N_5379,N_5582);
or U7421 (N_7421,N_5421,N_5252);
or U7422 (N_7422,N_5865,N_5825);
and U7423 (N_7423,N_5472,N_5945);
xor U7424 (N_7424,N_5929,N_5454);
or U7425 (N_7425,N_5472,N_6031);
nor U7426 (N_7426,N_5170,N_5270);
or U7427 (N_7427,N_5096,N_5837);
nand U7428 (N_7428,N_5029,N_6102);
xor U7429 (N_7429,N_5769,N_5122);
xnor U7430 (N_7430,N_5645,N_6122);
xnor U7431 (N_7431,N_5848,N_5045);
nand U7432 (N_7432,N_5621,N_5536);
and U7433 (N_7433,N_5398,N_5654);
nand U7434 (N_7434,N_5742,N_5833);
or U7435 (N_7435,N_6163,N_5319);
nor U7436 (N_7436,N_5378,N_6207);
and U7437 (N_7437,N_5147,N_5362);
nand U7438 (N_7438,N_5165,N_5716);
nor U7439 (N_7439,N_5531,N_5948);
or U7440 (N_7440,N_5921,N_5317);
nor U7441 (N_7441,N_5022,N_5809);
xor U7442 (N_7442,N_5562,N_5399);
or U7443 (N_7443,N_5429,N_6027);
nand U7444 (N_7444,N_5379,N_5415);
and U7445 (N_7445,N_6243,N_6222);
nor U7446 (N_7446,N_6188,N_5151);
and U7447 (N_7447,N_5706,N_5980);
and U7448 (N_7448,N_5730,N_5152);
or U7449 (N_7449,N_5252,N_6049);
and U7450 (N_7450,N_5623,N_5703);
and U7451 (N_7451,N_5892,N_5333);
or U7452 (N_7452,N_5615,N_5475);
and U7453 (N_7453,N_6205,N_5733);
and U7454 (N_7454,N_5962,N_6028);
nor U7455 (N_7455,N_6083,N_5379);
xnor U7456 (N_7456,N_5848,N_5316);
nor U7457 (N_7457,N_5832,N_6161);
xor U7458 (N_7458,N_5828,N_5561);
nand U7459 (N_7459,N_5491,N_6187);
or U7460 (N_7460,N_5375,N_5412);
nand U7461 (N_7461,N_5002,N_5921);
nor U7462 (N_7462,N_5049,N_6155);
and U7463 (N_7463,N_6107,N_5170);
and U7464 (N_7464,N_5096,N_5556);
nand U7465 (N_7465,N_5358,N_5047);
xor U7466 (N_7466,N_6229,N_5755);
or U7467 (N_7467,N_5849,N_5066);
nor U7468 (N_7468,N_5503,N_5793);
and U7469 (N_7469,N_6144,N_5202);
or U7470 (N_7470,N_5023,N_6249);
and U7471 (N_7471,N_6154,N_5308);
xor U7472 (N_7472,N_5789,N_6034);
or U7473 (N_7473,N_5753,N_5637);
nand U7474 (N_7474,N_6183,N_5220);
or U7475 (N_7475,N_5583,N_5623);
nand U7476 (N_7476,N_6061,N_6097);
xnor U7477 (N_7477,N_5539,N_6093);
nand U7478 (N_7478,N_5531,N_5936);
and U7479 (N_7479,N_5608,N_5745);
nand U7480 (N_7480,N_5620,N_5973);
nor U7481 (N_7481,N_5228,N_5002);
nor U7482 (N_7482,N_5189,N_6076);
xor U7483 (N_7483,N_6068,N_5360);
xor U7484 (N_7484,N_5241,N_5484);
and U7485 (N_7485,N_5326,N_5407);
xor U7486 (N_7486,N_5809,N_5859);
xnor U7487 (N_7487,N_5352,N_5966);
nand U7488 (N_7488,N_5947,N_5345);
nand U7489 (N_7489,N_6122,N_5895);
xor U7490 (N_7490,N_5482,N_6000);
or U7491 (N_7491,N_5189,N_5643);
and U7492 (N_7492,N_5315,N_5421);
and U7493 (N_7493,N_5631,N_6203);
nor U7494 (N_7494,N_5584,N_5462);
xnor U7495 (N_7495,N_5776,N_5788);
xor U7496 (N_7496,N_5702,N_5758);
xor U7497 (N_7497,N_5409,N_5870);
nor U7498 (N_7498,N_5798,N_5124);
nand U7499 (N_7499,N_5646,N_6035);
nor U7500 (N_7500,N_6681,N_6841);
nor U7501 (N_7501,N_6293,N_6898);
nor U7502 (N_7502,N_7398,N_6676);
and U7503 (N_7503,N_6949,N_6272);
and U7504 (N_7504,N_6350,N_6974);
or U7505 (N_7505,N_7208,N_6426);
xnor U7506 (N_7506,N_6634,N_6734);
xnor U7507 (N_7507,N_6398,N_7069);
and U7508 (N_7508,N_6325,N_6786);
or U7509 (N_7509,N_7475,N_7345);
nand U7510 (N_7510,N_6502,N_6929);
nor U7511 (N_7511,N_6274,N_6557);
and U7512 (N_7512,N_7034,N_6416);
xor U7513 (N_7513,N_6935,N_7369);
nor U7514 (N_7514,N_7453,N_7057);
nor U7515 (N_7515,N_7048,N_6905);
nand U7516 (N_7516,N_7065,N_6952);
xor U7517 (N_7517,N_6652,N_6304);
and U7518 (N_7518,N_6743,N_6998);
nand U7519 (N_7519,N_7148,N_7128);
nand U7520 (N_7520,N_6533,N_7095);
and U7521 (N_7521,N_7364,N_6314);
or U7522 (N_7522,N_6486,N_6447);
nor U7523 (N_7523,N_6461,N_6883);
and U7524 (N_7524,N_6972,N_7330);
nor U7525 (N_7525,N_6732,N_7438);
xnor U7526 (N_7526,N_6712,N_6751);
nor U7527 (N_7527,N_7221,N_6363);
and U7528 (N_7528,N_7104,N_6637);
xor U7529 (N_7529,N_6537,N_6921);
nor U7530 (N_7530,N_7219,N_7411);
nand U7531 (N_7531,N_6779,N_6451);
or U7532 (N_7532,N_6810,N_6744);
xnor U7533 (N_7533,N_6323,N_7175);
and U7534 (N_7534,N_7180,N_7483);
nor U7535 (N_7535,N_6377,N_6835);
nor U7536 (N_7536,N_6903,N_7185);
or U7537 (N_7537,N_6500,N_6573);
nand U7538 (N_7538,N_7113,N_7135);
or U7539 (N_7539,N_6780,N_7010);
nand U7540 (N_7540,N_7316,N_6704);
or U7541 (N_7541,N_6483,N_6262);
xnor U7542 (N_7542,N_6540,N_6402);
or U7543 (N_7543,N_6672,N_6971);
and U7544 (N_7544,N_6446,N_6899);
or U7545 (N_7545,N_6508,N_7380);
xor U7546 (N_7546,N_7144,N_7233);
nor U7547 (N_7547,N_6651,N_6376);
nor U7548 (N_7548,N_7377,N_6911);
and U7549 (N_7549,N_7348,N_6940);
nor U7550 (N_7550,N_7414,N_7226);
and U7551 (N_7551,N_6658,N_7045);
nand U7552 (N_7552,N_6526,N_6916);
or U7553 (N_7553,N_6393,N_6352);
and U7554 (N_7554,N_6963,N_6875);
xnor U7555 (N_7555,N_6589,N_6284);
nand U7556 (N_7556,N_6542,N_6730);
nand U7557 (N_7557,N_6296,N_7047);
nand U7558 (N_7558,N_6413,N_6522);
nor U7559 (N_7559,N_6607,N_6546);
nand U7560 (N_7560,N_6336,N_7477);
and U7561 (N_7561,N_6696,N_6485);
nor U7562 (N_7562,N_6392,N_7147);
xor U7563 (N_7563,N_6709,N_6406);
nand U7564 (N_7564,N_7202,N_6938);
and U7565 (N_7565,N_6547,N_6654);
or U7566 (N_7566,N_6509,N_6669);
xnor U7567 (N_7567,N_7370,N_7053);
and U7568 (N_7568,N_6846,N_6816);
nand U7569 (N_7569,N_6726,N_7440);
or U7570 (N_7570,N_6884,N_6452);
nor U7571 (N_7571,N_6610,N_7066);
and U7572 (N_7572,N_7344,N_7466);
and U7573 (N_7573,N_7012,N_7030);
xnor U7574 (N_7574,N_6682,N_7179);
xor U7575 (N_7575,N_6567,N_6317);
xnor U7576 (N_7576,N_6869,N_6775);
nand U7577 (N_7577,N_7035,N_7319);
and U7578 (N_7578,N_6995,N_6324);
nand U7579 (N_7579,N_6687,N_7323);
nand U7580 (N_7580,N_6424,N_6806);
or U7581 (N_7581,N_6504,N_6927);
and U7582 (N_7582,N_6563,N_6435);
or U7583 (N_7583,N_6467,N_7365);
nand U7584 (N_7584,N_7176,N_7161);
nand U7585 (N_7585,N_7401,N_7336);
nor U7586 (N_7586,N_7020,N_7082);
nand U7587 (N_7587,N_6805,N_6784);
and U7588 (N_7588,N_6878,N_7172);
xnor U7589 (N_7589,N_6590,N_6405);
and U7590 (N_7590,N_7357,N_7286);
nand U7591 (N_7591,N_6608,N_7402);
and U7592 (N_7592,N_6621,N_6997);
or U7593 (N_7593,N_6720,N_6866);
or U7594 (N_7594,N_6842,N_6962);
xnor U7595 (N_7595,N_6561,N_7284);
nor U7596 (N_7596,N_7397,N_6966);
nor U7597 (N_7597,N_7278,N_7299);
xor U7598 (N_7598,N_7085,N_7156);
or U7599 (N_7599,N_7014,N_6694);
xnor U7600 (N_7600,N_6993,N_7427);
nor U7601 (N_7601,N_6689,N_6260);
xnor U7602 (N_7602,N_7404,N_7400);
nor U7603 (N_7603,N_6987,N_7109);
nand U7604 (N_7604,N_7367,N_7498);
xor U7605 (N_7605,N_6517,N_6626);
nand U7606 (N_7606,N_6353,N_6341);
xnor U7607 (N_7607,N_7274,N_6450);
xor U7608 (N_7608,N_7496,N_6579);
xnor U7609 (N_7609,N_7435,N_6867);
nor U7610 (N_7610,N_6301,N_7416);
nor U7611 (N_7611,N_6918,N_6267);
and U7612 (N_7612,N_6415,N_7324);
nor U7613 (N_7613,N_6699,N_7228);
xor U7614 (N_7614,N_6263,N_6489);
or U7615 (N_7615,N_6339,N_6576);
and U7616 (N_7616,N_6438,N_7140);
or U7617 (N_7617,N_6913,N_6714);
xnor U7618 (N_7618,N_7386,N_7242);
nand U7619 (N_7619,N_6520,N_7063);
nand U7620 (N_7620,N_6470,N_6876);
nand U7621 (N_7621,N_6664,N_6365);
or U7622 (N_7622,N_6457,N_6863);
nand U7623 (N_7623,N_6641,N_7118);
and U7624 (N_7624,N_6719,N_6308);
or U7625 (N_7625,N_7258,N_6678);
nor U7626 (N_7626,N_6854,N_6991);
nand U7627 (N_7627,N_6978,N_7351);
nand U7628 (N_7628,N_7216,N_7042);
and U7629 (N_7629,N_6462,N_7004);
nor U7630 (N_7630,N_6787,N_7259);
nand U7631 (N_7631,N_6348,N_7439);
xor U7632 (N_7632,N_6748,N_6773);
nand U7633 (N_7633,N_7194,N_6311);
xor U7634 (N_7634,N_6631,N_6739);
and U7635 (N_7635,N_6662,N_6410);
nand U7636 (N_7636,N_7252,N_6443);
and U7637 (N_7637,N_6364,N_7317);
nand U7638 (N_7638,N_6812,N_6275);
nand U7639 (N_7639,N_7360,N_6697);
nand U7640 (N_7640,N_6737,N_7461);
xor U7641 (N_7641,N_6615,N_7268);
and U7642 (N_7642,N_7346,N_7025);
nand U7643 (N_7643,N_7335,N_7153);
nand U7644 (N_7644,N_6924,N_6956);
nor U7645 (N_7645,N_6320,N_6493);
or U7646 (N_7646,N_6853,N_6513);
or U7647 (N_7647,N_7120,N_6831);
nand U7648 (N_7648,N_6278,N_6407);
xnor U7649 (N_7649,N_7124,N_7467);
xor U7650 (N_7650,N_7392,N_7298);
or U7651 (N_7651,N_6635,N_6487);
and U7652 (N_7652,N_6767,N_6342);
nand U7653 (N_7653,N_6827,N_7205);
nor U7654 (N_7654,N_6616,N_6516);
nor U7655 (N_7655,N_7409,N_6727);
nor U7656 (N_7656,N_7471,N_7184);
nand U7657 (N_7657,N_6919,N_6448);
or U7658 (N_7658,N_7366,N_7111);
and U7659 (N_7659,N_6644,N_6981);
or U7660 (N_7660,N_6813,N_6915);
and U7661 (N_7661,N_6596,N_6569);
nor U7662 (N_7662,N_7302,N_6926);
nand U7663 (N_7663,N_6809,N_6481);
nor U7664 (N_7664,N_7432,N_6514);
and U7665 (N_7665,N_6477,N_7381);
nor U7666 (N_7666,N_6575,N_6560);
xor U7667 (N_7667,N_6396,N_6670);
xnor U7668 (N_7668,N_7385,N_6459);
and U7669 (N_7669,N_6894,N_6543);
and U7670 (N_7670,N_7350,N_7455);
xnor U7671 (N_7671,N_6584,N_6335);
xor U7672 (N_7672,N_6280,N_6856);
xor U7673 (N_7673,N_6553,N_6791);
or U7674 (N_7674,N_6925,N_7145);
nor U7675 (N_7675,N_7157,N_7277);
and U7676 (N_7676,N_6307,N_6361);
xnor U7677 (N_7677,N_6414,N_7245);
and U7678 (N_7678,N_6490,N_7015);
nor U7679 (N_7679,N_6985,N_6800);
or U7680 (N_7680,N_7134,N_7378);
nor U7681 (N_7681,N_7230,N_6781);
and U7682 (N_7682,N_7307,N_7193);
xnor U7683 (N_7683,N_7026,N_6713);
and U7684 (N_7684,N_6653,N_6265);
nand U7685 (N_7685,N_7059,N_6758);
and U7686 (N_7686,N_7490,N_7169);
or U7687 (N_7687,N_6783,N_7248);
or U7688 (N_7688,N_6454,N_6491);
or U7689 (N_7689,N_7072,N_7342);
xor U7690 (N_7690,N_7141,N_7390);
and U7691 (N_7691,N_6578,N_7181);
nand U7692 (N_7692,N_6297,N_7162);
or U7693 (N_7693,N_7333,N_6499);
and U7694 (N_7694,N_7368,N_7224);
xnor U7695 (N_7695,N_6735,N_6683);
nor U7696 (N_7696,N_7071,N_6897);
nand U7697 (N_7697,N_7287,N_6507);
and U7698 (N_7698,N_7343,N_7146);
or U7699 (N_7699,N_6439,N_7472);
xor U7700 (N_7700,N_6718,N_6945);
and U7701 (N_7701,N_6292,N_7003);
and U7702 (N_7702,N_7173,N_6506);
and U7703 (N_7703,N_6908,N_6917);
and U7704 (N_7704,N_7158,N_7257);
and U7705 (N_7705,N_7160,N_6822);
nand U7706 (N_7706,N_6871,N_7174);
and U7707 (N_7707,N_6371,N_6256);
and U7708 (N_7708,N_6288,N_6999);
nand U7709 (N_7709,N_6281,N_6638);
nand U7710 (N_7710,N_6961,N_6649);
and U7711 (N_7711,N_6347,N_7002);
xnor U7712 (N_7712,N_6552,N_7499);
nor U7713 (N_7713,N_7149,N_7449);
or U7714 (N_7714,N_7070,N_7426);
and U7715 (N_7715,N_6693,N_7288);
xor U7716 (N_7716,N_6826,N_7339);
nand U7717 (N_7717,N_6989,N_6891);
or U7718 (N_7718,N_7254,N_6928);
xnor U7719 (N_7719,N_6702,N_6852);
nand U7720 (N_7720,N_7285,N_7321);
or U7721 (N_7721,N_7131,N_6289);
nand U7722 (N_7722,N_6904,N_7136);
xnor U7723 (N_7723,N_6515,N_7265);
nor U7724 (N_7724,N_7138,N_6839);
xor U7725 (N_7725,N_6948,N_7340);
nand U7726 (N_7726,N_7039,N_7328);
or U7727 (N_7727,N_7320,N_7276);
and U7728 (N_7728,N_7130,N_7347);
or U7729 (N_7729,N_7044,N_6770);
or U7730 (N_7730,N_6630,N_6474);
nand U7731 (N_7731,N_7283,N_7001);
nor U7732 (N_7732,N_7210,N_7253);
nor U7733 (N_7733,N_7054,N_7083);
nor U7734 (N_7734,N_7052,N_7318);
nand U7735 (N_7735,N_6302,N_7207);
and U7736 (N_7736,N_6355,N_7204);
xnor U7737 (N_7737,N_6532,N_7217);
and U7738 (N_7738,N_6759,N_6668);
nor U7739 (N_7739,N_7206,N_7356);
nand U7740 (N_7740,N_6471,N_7363);
nand U7741 (N_7741,N_7308,N_6837);
nand U7742 (N_7742,N_7456,N_7215);
or U7743 (N_7743,N_6583,N_7101);
xnor U7744 (N_7744,N_7244,N_6711);
xor U7745 (N_7745,N_7355,N_6251);
nand U7746 (N_7746,N_6482,N_6738);
nor U7747 (N_7747,N_7457,N_6257);
nor U7748 (N_7748,N_7213,N_7338);
xnor U7749 (N_7749,N_6980,N_7227);
xnor U7750 (N_7750,N_6661,N_6671);
nor U7751 (N_7751,N_6266,N_6434);
nor U7752 (N_7752,N_6437,N_7168);
or U7753 (N_7753,N_6970,N_7068);
nand U7754 (N_7754,N_6521,N_7163);
and U7755 (N_7755,N_7186,N_6923);
nor U7756 (N_7756,N_7463,N_6544);
xnor U7757 (N_7757,N_6665,N_7275);
xnor U7758 (N_7758,N_7073,N_7492);
nand U7759 (N_7759,N_6942,N_7023);
and U7760 (N_7760,N_6975,N_7271);
xor U7761 (N_7761,N_6657,N_6494);
and U7762 (N_7762,N_6378,N_7470);
xnor U7763 (N_7763,N_7127,N_7129);
or U7764 (N_7764,N_6357,N_6954);
and U7765 (N_7765,N_6395,N_7087);
xor U7766 (N_7766,N_6534,N_7451);
nor U7767 (N_7767,N_6977,N_7376);
xor U7768 (N_7768,N_6893,N_6967);
xor U7769 (N_7769,N_6785,N_6880);
and U7770 (N_7770,N_6536,N_7099);
xnor U7771 (N_7771,N_6740,N_6648);
xnor U7772 (N_7772,N_6259,N_6855);
nor U7773 (N_7773,N_6725,N_7266);
xnor U7774 (N_7774,N_6582,N_7081);
or U7775 (N_7775,N_6468,N_6715);
or U7776 (N_7776,N_6306,N_6969);
or U7777 (N_7777,N_6707,N_6890);
xor U7778 (N_7778,N_7300,N_7491);
nand U7779 (N_7779,N_7079,N_6602);
or U7780 (N_7780,N_7291,N_6294);
and U7781 (N_7781,N_7112,N_7132);
xor U7782 (N_7782,N_6922,N_6555);
nor U7783 (N_7783,N_6287,N_7262);
or U7784 (N_7784,N_6619,N_6811);
nand U7785 (N_7785,N_7166,N_6895);
nand U7786 (N_7786,N_6310,N_6749);
nand U7787 (N_7787,N_7116,N_6959);
nand U7788 (N_7788,N_7263,N_6425);
and U7789 (N_7789,N_6369,N_6503);
or U7790 (N_7790,N_7220,N_7407);
and U7791 (N_7791,N_6828,N_7315);
and U7792 (N_7792,N_7088,N_6679);
nand U7793 (N_7793,N_6529,N_7322);
or U7794 (N_7794,N_6762,N_6777);
and U7795 (N_7795,N_6313,N_6585);
and U7796 (N_7796,N_7337,N_6857);
nand U7797 (N_7797,N_7165,N_7021);
nor U7798 (N_7798,N_6606,N_6271);
and U7799 (N_7799,N_6586,N_6303);
nand U7800 (N_7800,N_6383,N_6497);
nand U7801 (N_7801,N_6690,N_7009);
nand U7802 (N_7802,N_6958,N_7249);
nor U7803 (N_7803,N_6801,N_7445);
nand U7804 (N_7804,N_6545,N_6754);
nor U7805 (N_7805,N_7097,N_6939);
xor U7806 (N_7806,N_7067,N_6273);
nand U7807 (N_7807,N_6464,N_6799);
or U7808 (N_7808,N_7016,N_6283);
or U7809 (N_7809,N_6539,N_7279);
xor U7810 (N_7810,N_7353,N_6535);
xor U7811 (N_7811,N_7326,N_7024);
xor U7812 (N_7812,N_7464,N_6830);
and U7813 (N_7813,N_6473,N_6556);
xor U7814 (N_7814,N_6488,N_6788);
nor U7815 (N_7815,N_6327,N_6742);
nor U7816 (N_7816,N_7479,N_7029);
nor U7817 (N_7817,N_6331,N_6609);
nand U7818 (N_7818,N_6382,N_6733);
or U7819 (N_7819,N_7062,N_7056);
xor U7820 (N_7820,N_6312,N_7311);
and U7821 (N_7821,N_6408,N_6695);
nor U7822 (N_7822,N_7243,N_7159);
or U7823 (N_7823,N_6337,N_6409);
nand U7824 (N_7824,N_6255,N_6870);
or U7825 (N_7825,N_7028,N_6479);
nor U7826 (N_7826,N_6269,N_7123);
and U7827 (N_7827,N_6844,N_7334);
or U7828 (N_7828,N_6953,N_7151);
and U7829 (N_7829,N_6627,N_6458);
and U7830 (N_7830,N_7305,N_6701);
nand U7831 (N_7831,N_6492,N_6322);
xnor U7832 (N_7832,N_7005,N_6528);
xnor U7833 (N_7833,N_7375,N_6817);
or U7834 (N_7834,N_7481,N_7078);
xnor U7835 (N_7835,N_6444,N_7484);
xnor U7836 (N_7836,N_6937,N_7294);
nor U7837 (N_7837,N_7006,N_6531);
nor U7838 (N_7838,N_6976,N_6973);
nand U7839 (N_7839,N_6356,N_6882);
xnor U7840 (N_7840,N_6650,N_7108);
and U7841 (N_7841,N_6753,N_6527);
and U7842 (N_7842,N_7421,N_6333);
and U7843 (N_7843,N_6403,N_7306);
nand U7844 (N_7844,N_6418,N_7459);
and U7845 (N_7845,N_7177,N_7032);
xnor U7846 (N_7846,N_6614,N_6698);
nand U7847 (N_7847,N_7237,N_6309);
nor U7848 (N_7848,N_7256,N_7359);
nand U7849 (N_7849,N_7027,N_7289);
nor U7850 (N_7850,N_6815,N_6765);
xnor U7851 (N_7851,N_6512,N_6932);
or U7852 (N_7852,N_7329,N_6746);
nor U7853 (N_7853,N_6564,N_7013);
nand U7854 (N_7854,N_6673,N_6794);
or U7855 (N_7855,N_6776,N_6909);
and U7856 (N_7856,N_7121,N_6814);
xnor U7857 (N_7857,N_6797,N_6571);
nand U7858 (N_7858,N_7443,N_7474);
and U7859 (N_7859,N_7094,N_6549);
nand U7860 (N_7860,N_6505,N_6605);
and U7861 (N_7861,N_6326,N_6793);
xnor U7862 (N_7862,N_6404,N_6321);
xor U7863 (N_7863,N_6421,N_6642);
xor U7864 (N_7864,N_7164,N_7198);
or U7865 (N_7865,N_7431,N_7423);
xnor U7866 (N_7866,N_6947,N_6285);
nor U7867 (N_7867,N_7225,N_7465);
and U7868 (N_7868,N_6343,N_6384);
and U7869 (N_7869,N_6286,N_7497);
nand U7870 (N_7870,N_6849,N_7086);
nor U7871 (N_7871,N_6778,N_7191);
xnor U7872 (N_7872,N_6807,N_6675);
nand U7873 (N_7873,N_6722,N_6595);
xnor U7874 (N_7874,N_7267,N_6752);
xor U7875 (N_7875,N_7417,N_6588);
and U7876 (N_7876,N_7077,N_6340);
or U7877 (N_7877,N_6562,N_6756);
nor U7878 (N_7878,N_7406,N_6769);
xnor U7879 (N_7879,N_6618,N_7061);
nor U7880 (N_7880,N_6747,N_6423);
xor U7881 (N_7881,N_7246,N_7152);
or U7882 (N_7882,N_7234,N_6864);
and U7883 (N_7883,N_7040,N_6677);
and U7884 (N_7884,N_7117,N_6572);
xor U7885 (N_7885,N_6836,N_7485);
and U7886 (N_7886,N_6881,N_6757);
nor U7887 (N_7887,N_6463,N_7167);
or U7888 (N_7888,N_6795,N_6933);
xor U7889 (N_7889,N_6684,N_6299);
nand U7890 (N_7890,N_6934,N_7084);
and U7891 (N_7891,N_6655,N_6349);
nor U7892 (N_7892,N_6873,N_6375);
and U7893 (N_7893,N_6790,N_6253);
or U7894 (N_7894,N_6982,N_6736);
and U7895 (N_7895,N_6436,N_7241);
nand U7896 (N_7896,N_6600,N_6632);
nand U7897 (N_7897,N_6859,N_7436);
nor U7898 (N_7898,N_6660,N_6766);
or U7899 (N_7899,N_6902,N_6374);
and U7900 (N_7900,N_6441,N_7495);
and U7901 (N_7901,N_6832,N_7211);
xnor U7902 (N_7902,N_6510,N_6329);
nor U7903 (N_7903,N_6834,N_6388);
nor U7904 (N_7904,N_7110,N_6354);
nand U7905 (N_7905,N_6495,N_6291);
xnor U7906 (N_7906,N_7125,N_6772);
nor U7907 (N_7907,N_7058,N_7096);
nor U7908 (N_7908,N_6358,N_6745);
nand U7909 (N_7909,N_6565,N_6829);
and U7910 (N_7910,N_7212,N_7214);
nor U7911 (N_7911,N_6680,N_6700);
xnor U7912 (N_7912,N_6957,N_7430);
nand U7913 (N_7913,N_7038,N_6639);
nor U7914 (N_7914,N_6886,N_6659);
nor U7915 (N_7915,N_7396,N_6819);
and U7916 (N_7916,N_7037,N_6420);
and U7917 (N_7917,N_7049,N_6433);
nor U7918 (N_7918,N_6907,N_7458);
nor U7919 (N_7919,N_7280,N_6782);
or U7920 (N_7920,N_7428,N_6910);
nand U7921 (N_7921,N_6647,N_7195);
nand U7922 (N_7922,N_7296,N_6686);
xor U7923 (N_7923,N_6319,N_6599);
xnor U7924 (N_7924,N_7126,N_6798);
nor U7925 (N_7925,N_7420,N_6900);
xnor U7926 (N_7926,N_7142,N_6877);
and U7927 (N_7927,N_7192,N_6611);
and U7928 (N_7928,N_7405,N_6628);
xnor U7929 (N_7929,N_6721,N_7255);
nor U7930 (N_7930,N_7229,N_7238);
xnor U7931 (N_7931,N_7310,N_7442);
nor U7932 (N_7932,N_7133,N_7064);
and U7933 (N_7933,N_7408,N_6428);
xnor U7934 (N_7934,N_7240,N_6845);
xor U7935 (N_7935,N_7482,N_7388);
xor U7936 (N_7936,N_6268,N_7107);
or U7937 (N_7937,N_6295,N_6594);
or U7938 (N_7938,N_7199,N_7489);
and U7939 (N_7939,N_7115,N_6808);
nor U7940 (N_7940,N_6518,N_6625);
nand U7941 (N_7941,N_7270,N_6861);
and U7942 (N_7942,N_6362,N_7494);
xor U7943 (N_7943,N_6601,N_6417);
or U7944 (N_7944,N_7476,N_7422);
nor U7945 (N_7945,N_6351,N_7410);
nor U7946 (N_7946,N_7017,N_6768);
or U7947 (N_7947,N_6685,N_6858);
and U7948 (N_7948,N_7170,N_7383);
nand U7949 (N_7949,N_6366,N_7473);
nor U7950 (N_7950,N_6710,N_7281);
and U7951 (N_7951,N_6906,N_6568);
nor U7952 (N_7952,N_6663,N_6604);
nor U7953 (N_7953,N_6442,N_6796);
xnor U7954 (N_7954,N_7074,N_6723);
or U7955 (N_7955,N_6760,N_7209);
nor U7956 (N_7956,N_6896,N_7060);
nand U7957 (N_7957,N_7137,N_6332);
xnor U7958 (N_7958,N_7041,N_6623);
and U7959 (N_7959,N_7187,N_6823);
and U7960 (N_7960,N_7196,N_7327);
xnor U7961 (N_7961,N_7332,N_6612);
and U7962 (N_7962,N_7203,N_7478);
nor U7963 (N_7963,N_7106,N_6465);
nand U7964 (N_7964,N_6636,N_6430);
and U7965 (N_7965,N_6551,N_6381);
xor U7966 (N_7966,N_6617,N_6821);
and U7967 (N_7967,N_6764,N_6334);
or U7968 (N_7968,N_7293,N_7139);
xnor U7969 (N_7969,N_7269,N_6724);
nor U7970 (N_7970,N_7018,N_6419);
and U7971 (N_7971,N_6580,N_6789);
xnor U7972 (N_7972,N_6988,N_7387);
nor U7973 (N_7973,N_6622,N_7309);
xor U7974 (N_7974,N_6692,N_7358);
or U7975 (N_7975,N_6761,N_7119);
and U7976 (N_7976,N_6960,N_6305);
nand U7977 (N_7977,N_7122,N_6755);
and U7978 (N_7978,N_6771,N_6252);
and U7979 (N_7979,N_6951,N_6792);
nand U7980 (N_7980,N_6472,N_6865);
or U7981 (N_7981,N_7092,N_6843);
or U7982 (N_7982,N_6538,N_6386);
xor U7983 (N_7983,N_7000,N_7349);
and U7984 (N_7984,N_6346,N_7182);
or U7985 (N_7985,N_6731,N_6597);
nand U7986 (N_7986,N_6401,N_7362);
nor U7987 (N_7987,N_7183,N_6432);
or U7988 (N_7988,N_6892,N_6277);
nor U7989 (N_7989,N_6559,N_6717);
xor U7990 (N_7990,N_7091,N_6888);
or U7991 (N_7991,N_6691,N_6548);
xnor U7992 (N_7992,N_6577,N_7452);
nand U7993 (N_7993,N_7239,N_6901);
xnor U7994 (N_7994,N_7448,N_7273);
nor U7995 (N_7995,N_6554,N_6936);
nand U7996 (N_7996,N_7011,N_6345);
nor U7997 (N_7997,N_7098,N_7022);
nor U7998 (N_7998,N_7372,N_6920);
xnor U7999 (N_7999,N_7301,N_7080);
or U8000 (N_8000,N_7419,N_7303);
xor U8001 (N_8001,N_6399,N_6412);
nand U8002 (N_8002,N_7250,N_7007);
xnor U8003 (N_8003,N_6656,N_6429);
or U8004 (N_8004,N_6541,N_6391);
and U8005 (N_8005,N_6804,N_6645);
xor U8006 (N_8006,N_6422,N_6833);
and U8007 (N_8007,N_7260,N_7075);
xor U8008 (N_8008,N_7469,N_7462);
and U8009 (N_8009,N_6818,N_7008);
or U8010 (N_8010,N_7292,N_6624);
or U8011 (N_8011,N_6592,N_7076);
or U8012 (N_8012,N_6629,N_6965);
xnor U8013 (N_8013,N_6848,N_7031);
nor U8014 (N_8014,N_6613,N_6368);
nand U8015 (N_8015,N_7222,N_7487);
and U8016 (N_8016,N_6943,N_6431);
or U8017 (N_8017,N_7354,N_6992);
nor U8018 (N_8018,N_6276,N_6344);
or U8019 (N_8019,N_6674,N_6498);
nand U8020 (N_8020,N_7437,N_6282);
and U8021 (N_8021,N_7403,N_6633);
and U8022 (N_8022,N_6703,N_6370);
nand U8023 (N_8023,N_6390,N_6480);
and U8024 (N_8024,N_6254,N_6587);
and U8025 (N_8025,N_6328,N_7189);
nor U8026 (N_8026,N_6258,N_7261);
or U8027 (N_8027,N_6496,N_6372);
nor U8028 (N_8028,N_7413,N_6868);
or U8029 (N_8029,N_6440,N_7236);
nand U8030 (N_8030,N_7036,N_7190);
nor U8031 (N_8031,N_7295,N_6367);
and U8032 (N_8032,N_6968,N_7418);
nand U8033 (N_8033,N_6300,N_6469);
and U8034 (N_8034,N_7231,N_7460);
and U8035 (N_8035,N_6941,N_6824);
and U8036 (N_8036,N_6708,N_6990);
nand U8037 (N_8037,N_6946,N_6449);
xnor U8038 (N_8038,N_6774,N_6593);
or U8039 (N_8039,N_6387,N_6729);
and U8040 (N_8040,N_6874,N_7188);
xnor U8041 (N_8041,N_6298,N_6574);
nand U8042 (N_8042,N_7391,N_6840);
xor U8043 (N_8043,N_7331,N_7447);
and U8044 (N_8044,N_6850,N_7399);
nand U8045 (N_8045,N_6373,N_6741);
and U8046 (N_8046,N_6728,N_6290);
nor U8047 (N_8047,N_6820,N_7446);
nand U8048 (N_8048,N_7312,N_6984);
or U8049 (N_8049,N_7379,N_7223);
nor U8050 (N_8050,N_7314,N_7200);
or U8051 (N_8051,N_7382,N_6250);
and U8052 (N_8052,N_6558,N_6466);
nor U8053 (N_8053,N_6887,N_6385);
nor U8054 (N_8054,N_6261,N_6851);
nand U8055 (N_8055,N_6803,N_7493);
nor U8056 (N_8056,N_6872,N_6640);
and U8057 (N_8057,N_7043,N_6996);
nand U8058 (N_8058,N_6994,N_6860);
or U8059 (N_8059,N_7434,N_6270);
or U8060 (N_8060,N_7425,N_6838);
nor U8061 (N_8061,N_6931,N_6667);
nor U8062 (N_8062,N_6705,N_7093);
nand U8063 (N_8063,N_6360,N_7050);
xor U8064 (N_8064,N_6979,N_6598);
or U8065 (N_8065,N_7272,N_6523);
xor U8066 (N_8066,N_7290,N_7178);
nor U8067 (N_8067,N_6646,N_7105);
or U8068 (N_8068,N_6318,N_7374);
or U8069 (N_8069,N_7450,N_6847);
nand U8070 (N_8070,N_6986,N_6944);
nor U8071 (N_8071,N_6950,N_6511);
or U8072 (N_8072,N_7384,N_7201);
or U8073 (N_8073,N_7415,N_7171);
nor U8074 (N_8074,N_7264,N_6930);
xor U8075 (N_8075,N_6581,N_7247);
nand U8076 (N_8076,N_7089,N_7197);
and U8077 (N_8077,N_7304,N_6802);
or U8078 (N_8078,N_6964,N_7486);
nand U8079 (N_8079,N_7412,N_6359);
and U8080 (N_8080,N_7055,N_6889);
nor U8081 (N_8081,N_6912,N_6862);
and U8082 (N_8082,N_6456,N_7100);
nand U8083 (N_8083,N_6688,N_7429);
and U8084 (N_8084,N_6879,N_6566);
or U8085 (N_8085,N_7102,N_6453);
or U8086 (N_8086,N_6914,N_7395);
nor U8087 (N_8087,N_7361,N_6394);
or U8088 (N_8088,N_6643,N_7394);
xor U8089 (N_8089,N_6484,N_7232);
and U8090 (N_8090,N_7488,N_6524);
and U8091 (N_8091,N_7235,N_7480);
or U8092 (N_8092,N_6389,N_6264);
nor U8093 (N_8093,N_7297,N_6460);
nor U8094 (N_8094,N_6445,N_6411);
and U8095 (N_8095,N_6666,N_6478);
nand U8096 (N_8096,N_7150,N_6379);
or U8097 (N_8097,N_7046,N_7051);
nor U8098 (N_8098,N_6475,N_6501);
or U8099 (N_8099,N_6476,N_6716);
and U8100 (N_8100,N_6397,N_7393);
xnor U8101 (N_8101,N_6620,N_6570);
nand U8102 (N_8102,N_6525,N_6316);
nor U8103 (N_8103,N_7352,N_6591);
nand U8104 (N_8104,N_7218,N_7103);
or U8105 (N_8105,N_7114,N_7341);
and U8106 (N_8106,N_6603,N_6550);
xnor U8107 (N_8107,N_6530,N_6400);
nand U8108 (N_8108,N_6825,N_7155);
nor U8109 (N_8109,N_7444,N_7019);
nand U8110 (N_8110,N_6338,N_7433);
xnor U8111 (N_8111,N_6455,N_6763);
or U8112 (N_8112,N_6315,N_7325);
or U8113 (N_8113,N_6983,N_7424);
or U8114 (N_8114,N_6706,N_7468);
or U8115 (N_8115,N_7371,N_6330);
nand U8116 (N_8116,N_7251,N_6279);
xor U8117 (N_8117,N_7282,N_7154);
xnor U8118 (N_8118,N_7143,N_7090);
nand U8119 (N_8119,N_6750,N_6427);
and U8120 (N_8120,N_7441,N_7033);
nor U8121 (N_8121,N_6885,N_7389);
nand U8122 (N_8122,N_6519,N_6380);
nor U8123 (N_8123,N_6955,N_7454);
or U8124 (N_8124,N_7313,N_7373);
nand U8125 (N_8125,N_6417,N_7250);
or U8126 (N_8126,N_6284,N_7290);
xor U8127 (N_8127,N_7060,N_6748);
xor U8128 (N_8128,N_6829,N_6630);
xnor U8129 (N_8129,N_6769,N_6323);
and U8130 (N_8130,N_7309,N_6927);
xor U8131 (N_8131,N_6953,N_7195);
or U8132 (N_8132,N_6930,N_6847);
xor U8133 (N_8133,N_7463,N_6754);
nor U8134 (N_8134,N_7349,N_6752);
or U8135 (N_8135,N_7234,N_6267);
or U8136 (N_8136,N_7400,N_7484);
or U8137 (N_8137,N_6456,N_7395);
and U8138 (N_8138,N_6988,N_6585);
and U8139 (N_8139,N_6677,N_6690);
nor U8140 (N_8140,N_7454,N_7276);
or U8141 (N_8141,N_6724,N_6972);
or U8142 (N_8142,N_6737,N_6999);
nor U8143 (N_8143,N_6462,N_6804);
or U8144 (N_8144,N_6482,N_6419);
xor U8145 (N_8145,N_7417,N_6587);
nand U8146 (N_8146,N_7101,N_6917);
and U8147 (N_8147,N_7404,N_7148);
nor U8148 (N_8148,N_7201,N_6986);
and U8149 (N_8149,N_6884,N_6405);
and U8150 (N_8150,N_6552,N_6420);
nand U8151 (N_8151,N_7362,N_7417);
nor U8152 (N_8152,N_6790,N_7397);
or U8153 (N_8153,N_7133,N_6824);
and U8154 (N_8154,N_6651,N_6732);
xnor U8155 (N_8155,N_6680,N_6796);
xnor U8156 (N_8156,N_7387,N_6550);
nand U8157 (N_8157,N_6395,N_6968);
nor U8158 (N_8158,N_6480,N_6271);
xnor U8159 (N_8159,N_6341,N_6955);
or U8160 (N_8160,N_6369,N_6316);
nor U8161 (N_8161,N_6637,N_7303);
nand U8162 (N_8162,N_7353,N_7028);
and U8163 (N_8163,N_7286,N_6313);
xnor U8164 (N_8164,N_6395,N_6633);
xnor U8165 (N_8165,N_6850,N_6276);
xnor U8166 (N_8166,N_6651,N_7227);
nor U8167 (N_8167,N_7063,N_7154);
and U8168 (N_8168,N_7185,N_7155);
and U8169 (N_8169,N_7109,N_6394);
and U8170 (N_8170,N_6250,N_6695);
xnor U8171 (N_8171,N_6497,N_7007);
nor U8172 (N_8172,N_7473,N_6795);
xnor U8173 (N_8173,N_7433,N_7435);
and U8174 (N_8174,N_6362,N_6792);
or U8175 (N_8175,N_6681,N_7364);
or U8176 (N_8176,N_7372,N_6293);
or U8177 (N_8177,N_6845,N_6629);
and U8178 (N_8178,N_6714,N_6369);
nor U8179 (N_8179,N_6458,N_6466);
xor U8180 (N_8180,N_6400,N_6890);
nand U8181 (N_8181,N_7241,N_6844);
or U8182 (N_8182,N_6497,N_7446);
nand U8183 (N_8183,N_6652,N_6390);
xor U8184 (N_8184,N_7111,N_6488);
nand U8185 (N_8185,N_6611,N_6319);
nor U8186 (N_8186,N_6376,N_6755);
xnor U8187 (N_8187,N_6990,N_6671);
or U8188 (N_8188,N_6929,N_7212);
nor U8189 (N_8189,N_6294,N_7269);
and U8190 (N_8190,N_6915,N_6897);
nand U8191 (N_8191,N_6659,N_6898);
nand U8192 (N_8192,N_6770,N_7055);
nor U8193 (N_8193,N_6651,N_7448);
or U8194 (N_8194,N_6283,N_7055);
nand U8195 (N_8195,N_7280,N_7209);
and U8196 (N_8196,N_6405,N_7137);
nand U8197 (N_8197,N_7297,N_6779);
or U8198 (N_8198,N_7390,N_6426);
nand U8199 (N_8199,N_7467,N_6771);
or U8200 (N_8200,N_6863,N_7099);
nand U8201 (N_8201,N_6357,N_6504);
nor U8202 (N_8202,N_7299,N_7105);
or U8203 (N_8203,N_7388,N_7109);
or U8204 (N_8204,N_6773,N_6498);
nand U8205 (N_8205,N_7434,N_6645);
nand U8206 (N_8206,N_7403,N_6623);
nand U8207 (N_8207,N_7212,N_6655);
xor U8208 (N_8208,N_6409,N_6548);
nand U8209 (N_8209,N_6506,N_6396);
nand U8210 (N_8210,N_6407,N_7364);
or U8211 (N_8211,N_6469,N_6950);
xor U8212 (N_8212,N_7227,N_6617);
xnor U8213 (N_8213,N_7361,N_7380);
and U8214 (N_8214,N_7369,N_6674);
or U8215 (N_8215,N_7124,N_7369);
nand U8216 (N_8216,N_7370,N_7063);
xor U8217 (N_8217,N_6471,N_6296);
and U8218 (N_8218,N_7238,N_6328);
and U8219 (N_8219,N_7179,N_6908);
xor U8220 (N_8220,N_6481,N_6917);
or U8221 (N_8221,N_6828,N_7489);
nand U8222 (N_8222,N_7141,N_6853);
and U8223 (N_8223,N_6969,N_7078);
nor U8224 (N_8224,N_7365,N_6740);
or U8225 (N_8225,N_6699,N_7059);
nor U8226 (N_8226,N_7274,N_6378);
nand U8227 (N_8227,N_6366,N_7271);
nor U8228 (N_8228,N_6790,N_7072);
xnor U8229 (N_8229,N_6337,N_6941);
nand U8230 (N_8230,N_6794,N_6828);
xnor U8231 (N_8231,N_6911,N_7049);
or U8232 (N_8232,N_7482,N_6451);
xor U8233 (N_8233,N_6619,N_6282);
and U8234 (N_8234,N_7484,N_6932);
and U8235 (N_8235,N_6996,N_6475);
nor U8236 (N_8236,N_7422,N_6905);
and U8237 (N_8237,N_6706,N_6636);
and U8238 (N_8238,N_7050,N_6436);
nand U8239 (N_8239,N_6389,N_6400);
xnor U8240 (N_8240,N_7172,N_6717);
xor U8241 (N_8241,N_6890,N_6555);
or U8242 (N_8242,N_6591,N_7156);
nand U8243 (N_8243,N_6861,N_6630);
and U8244 (N_8244,N_6383,N_7149);
nor U8245 (N_8245,N_7424,N_7480);
or U8246 (N_8246,N_6660,N_6827);
or U8247 (N_8247,N_6623,N_6633);
xor U8248 (N_8248,N_6787,N_6579);
or U8249 (N_8249,N_6434,N_7121);
nor U8250 (N_8250,N_6671,N_6853);
xor U8251 (N_8251,N_6538,N_6505);
nand U8252 (N_8252,N_6835,N_7352);
nor U8253 (N_8253,N_6417,N_7285);
nor U8254 (N_8254,N_6949,N_6880);
xnor U8255 (N_8255,N_7332,N_6750);
nor U8256 (N_8256,N_6798,N_7070);
nor U8257 (N_8257,N_7422,N_7325);
or U8258 (N_8258,N_6336,N_6375);
nand U8259 (N_8259,N_7368,N_6922);
and U8260 (N_8260,N_6901,N_6889);
and U8261 (N_8261,N_7347,N_6528);
and U8262 (N_8262,N_7092,N_6847);
xnor U8263 (N_8263,N_7471,N_6920);
or U8264 (N_8264,N_6968,N_7121);
and U8265 (N_8265,N_7372,N_6931);
nor U8266 (N_8266,N_7379,N_7456);
xnor U8267 (N_8267,N_6948,N_6577);
xnor U8268 (N_8268,N_6253,N_6839);
xnor U8269 (N_8269,N_7308,N_6368);
nor U8270 (N_8270,N_7272,N_7299);
and U8271 (N_8271,N_6607,N_6256);
nor U8272 (N_8272,N_7415,N_6819);
and U8273 (N_8273,N_6407,N_6429);
xnor U8274 (N_8274,N_7025,N_6460);
xor U8275 (N_8275,N_7496,N_6318);
nor U8276 (N_8276,N_7477,N_7134);
or U8277 (N_8277,N_7226,N_6435);
nor U8278 (N_8278,N_6734,N_6771);
nand U8279 (N_8279,N_7350,N_7281);
or U8280 (N_8280,N_6820,N_6977);
nor U8281 (N_8281,N_7433,N_7097);
xnor U8282 (N_8282,N_6871,N_7158);
or U8283 (N_8283,N_7477,N_6470);
or U8284 (N_8284,N_6563,N_6565);
nor U8285 (N_8285,N_6518,N_6312);
xor U8286 (N_8286,N_6669,N_6813);
nor U8287 (N_8287,N_7478,N_6304);
nor U8288 (N_8288,N_6912,N_7433);
and U8289 (N_8289,N_7332,N_6496);
and U8290 (N_8290,N_6853,N_7417);
and U8291 (N_8291,N_6962,N_6369);
nor U8292 (N_8292,N_7404,N_7058);
and U8293 (N_8293,N_7169,N_6590);
nor U8294 (N_8294,N_6707,N_7341);
and U8295 (N_8295,N_6492,N_7422);
nor U8296 (N_8296,N_6884,N_7124);
nor U8297 (N_8297,N_6728,N_6301);
nor U8298 (N_8298,N_6999,N_6652);
nand U8299 (N_8299,N_6466,N_6268);
xor U8300 (N_8300,N_6299,N_7068);
or U8301 (N_8301,N_7451,N_6618);
nand U8302 (N_8302,N_6940,N_7168);
xnor U8303 (N_8303,N_7335,N_6829);
or U8304 (N_8304,N_6695,N_7421);
nor U8305 (N_8305,N_7337,N_7325);
nand U8306 (N_8306,N_6700,N_6547);
xor U8307 (N_8307,N_6453,N_6760);
or U8308 (N_8308,N_7499,N_7133);
xor U8309 (N_8309,N_7161,N_6670);
or U8310 (N_8310,N_6279,N_6879);
or U8311 (N_8311,N_6936,N_6881);
xnor U8312 (N_8312,N_7033,N_6543);
xor U8313 (N_8313,N_6697,N_6952);
xor U8314 (N_8314,N_7411,N_6709);
xnor U8315 (N_8315,N_6328,N_6973);
and U8316 (N_8316,N_6708,N_7322);
nor U8317 (N_8317,N_6989,N_7324);
or U8318 (N_8318,N_6323,N_6338);
and U8319 (N_8319,N_6449,N_6663);
xnor U8320 (N_8320,N_6951,N_6609);
and U8321 (N_8321,N_6809,N_6495);
nand U8322 (N_8322,N_7030,N_7470);
nand U8323 (N_8323,N_7480,N_6640);
nand U8324 (N_8324,N_6631,N_7045);
xnor U8325 (N_8325,N_7425,N_6304);
or U8326 (N_8326,N_6338,N_6324);
or U8327 (N_8327,N_7141,N_7351);
xor U8328 (N_8328,N_7298,N_6836);
nor U8329 (N_8329,N_7344,N_7016);
and U8330 (N_8330,N_7369,N_7401);
and U8331 (N_8331,N_6602,N_7104);
nor U8332 (N_8332,N_7421,N_7026);
and U8333 (N_8333,N_6296,N_6656);
or U8334 (N_8334,N_7434,N_7204);
and U8335 (N_8335,N_7241,N_7345);
or U8336 (N_8336,N_6494,N_7384);
xnor U8337 (N_8337,N_6821,N_7073);
nor U8338 (N_8338,N_7214,N_6407);
xor U8339 (N_8339,N_6272,N_7097);
or U8340 (N_8340,N_6556,N_6407);
and U8341 (N_8341,N_7242,N_6559);
or U8342 (N_8342,N_7307,N_7003);
xor U8343 (N_8343,N_7009,N_7217);
or U8344 (N_8344,N_7316,N_6969);
or U8345 (N_8345,N_6752,N_6955);
xnor U8346 (N_8346,N_7316,N_6655);
nor U8347 (N_8347,N_6805,N_6859);
xnor U8348 (N_8348,N_7208,N_6863);
or U8349 (N_8349,N_6441,N_6583);
and U8350 (N_8350,N_6536,N_7042);
nand U8351 (N_8351,N_7242,N_6928);
nand U8352 (N_8352,N_7075,N_6508);
or U8353 (N_8353,N_6690,N_6881);
nand U8354 (N_8354,N_7167,N_6559);
and U8355 (N_8355,N_6378,N_7099);
and U8356 (N_8356,N_6702,N_7383);
xnor U8357 (N_8357,N_7411,N_6551);
or U8358 (N_8358,N_6634,N_6295);
or U8359 (N_8359,N_6861,N_6913);
xor U8360 (N_8360,N_6572,N_6356);
nor U8361 (N_8361,N_7256,N_6652);
nor U8362 (N_8362,N_7449,N_6948);
and U8363 (N_8363,N_6797,N_7370);
and U8364 (N_8364,N_6628,N_7200);
nor U8365 (N_8365,N_6778,N_6353);
xnor U8366 (N_8366,N_6568,N_7061);
xor U8367 (N_8367,N_6857,N_7099);
nand U8368 (N_8368,N_7452,N_6358);
and U8369 (N_8369,N_7030,N_7468);
nand U8370 (N_8370,N_6868,N_6851);
xnor U8371 (N_8371,N_6319,N_6725);
xnor U8372 (N_8372,N_6780,N_7350);
or U8373 (N_8373,N_6686,N_6255);
or U8374 (N_8374,N_7239,N_6330);
nand U8375 (N_8375,N_6536,N_7494);
nor U8376 (N_8376,N_6269,N_6407);
xor U8377 (N_8377,N_6775,N_6407);
nor U8378 (N_8378,N_6299,N_6758);
xor U8379 (N_8379,N_7456,N_7407);
nor U8380 (N_8380,N_6999,N_6874);
or U8381 (N_8381,N_7192,N_6686);
xnor U8382 (N_8382,N_7051,N_7183);
and U8383 (N_8383,N_6641,N_7075);
and U8384 (N_8384,N_6912,N_7289);
and U8385 (N_8385,N_6978,N_7112);
xnor U8386 (N_8386,N_6349,N_6770);
and U8387 (N_8387,N_6749,N_6797);
and U8388 (N_8388,N_6509,N_7106);
and U8389 (N_8389,N_6611,N_6645);
or U8390 (N_8390,N_7059,N_6251);
or U8391 (N_8391,N_6381,N_6334);
nor U8392 (N_8392,N_7440,N_7118);
xor U8393 (N_8393,N_7233,N_6533);
nand U8394 (N_8394,N_6497,N_6278);
or U8395 (N_8395,N_6529,N_7006);
and U8396 (N_8396,N_6510,N_7165);
or U8397 (N_8397,N_6464,N_7105);
nand U8398 (N_8398,N_6990,N_6793);
and U8399 (N_8399,N_6929,N_7423);
and U8400 (N_8400,N_7403,N_6337);
nor U8401 (N_8401,N_7018,N_7392);
nor U8402 (N_8402,N_7362,N_7249);
nand U8403 (N_8403,N_7240,N_6683);
xnor U8404 (N_8404,N_7214,N_7412);
xnor U8405 (N_8405,N_6653,N_6429);
or U8406 (N_8406,N_7432,N_6890);
xnor U8407 (N_8407,N_6426,N_6462);
and U8408 (N_8408,N_6764,N_6305);
nand U8409 (N_8409,N_7141,N_6539);
nand U8410 (N_8410,N_6743,N_6286);
and U8411 (N_8411,N_6961,N_6512);
nor U8412 (N_8412,N_6441,N_6467);
nand U8413 (N_8413,N_6939,N_6997);
or U8414 (N_8414,N_7388,N_6400);
nand U8415 (N_8415,N_7324,N_7077);
xor U8416 (N_8416,N_6561,N_7041);
or U8417 (N_8417,N_6433,N_6432);
xor U8418 (N_8418,N_7446,N_7200);
xor U8419 (N_8419,N_7169,N_7485);
and U8420 (N_8420,N_7448,N_6510);
and U8421 (N_8421,N_7458,N_6389);
nand U8422 (N_8422,N_7178,N_7291);
nor U8423 (N_8423,N_7140,N_6463);
or U8424 (N_8424,N_7122,N_6749);
and U8425 (N_8425,N_7410,N_7141);
or U8426 (N_8426,N_6724,N_6956);
or U8427 (N_8427,N_6605,N_6627);
nand U8428 (N_8428,N_7013,N_7305);
and U8429 (N_8429,N_6802,N_6357);
and U8430 (N_8430,N_6489,N_6257);
nor U8431 (N_8431,N_6824,N_6308);
and U8432 (N_8432,N_6778,N_7184);
xor U8433 (N_8433,N_6572,N_7480);
nand U8434 (N_8434,N_6854,N_6559);
nor U8435 (N_8435,N_7304,N_7109);
nor U8436 (N_8436,N_6456,N_7249);
nand U8437 (N_8437,N_7356,N_6290);
nand U8438 (N_8438,N_6371,N_6499);
nand U8439 (N_8439,N_7009,N_6720);
and U8440 (N_8440,N_6711,N_6974);
nor U8441 (N_8441,N_7495,N_6514);
and U8442 (N_8442,N_6847,N_6483);
or U8443 (N_8443,N_6980,N_7266);
nor U8444 (N_8444,N_7091,N_6259);
or U8445 (N_8445,N_6625,N_7466);
nor U8446 (N_8446,N_7250,N_7011);
nor U8447 (N_8447,N_7031,N_6369);
xnor U8448 (N_8448,N_6722,N_6293);
xnor U8449 (N_8449,N_6940,N_7431);
nor U8450 (N_8450,N_6368,N_6590);
nor U8451 (N_8451,N_6976,N_6788);
or U8452 (N_8452,N_6485,N_7034);
nand U8453 (N_8453,N_6572,N_6723);
nand U8454 (N_8454,N_7316,N_6589);
xnor U8455 (N_8455,N_7477,N_6398);
and U8456 (N_8456,N_6646,N_6597);
and U8457 (N_8457,N_6865,N_7240);
xor U8458 (N_8458,N_7163,N_6610);
or U8459 (N_8459,N_7342,N_6940);
nor U8460 (N_8460,N_7248,N_7452);
or U8461 (N_8461,N_6623,N_7367);
or U8462 (N_8462,N_7413,N_6892);
or U8463 (N_8463,N_6381,N_7287);
nand U8464 (N_8464,N_6941,N_7459);
or U8465 (N_8465,N_6662,N_7202);
and U8466 (N_8466,N_7443,N_6448);
or U8467 (N_8467,N_6488,N_6480);
or U8468 (N_8468,N_7331,N_6555);
nand U8469 (N_8469,N_7475,N_7372);
or U8470 (N_8470,N_7152,N_6474);
or U8471 (N_8471,N_6607,N_6944);
or U8472 (N_8472,N_7059,N_6720);
or U8473 (N_8473,N_6870,N_7058);
nand U8474 (N_8474,N_6318,N_6943);
and U8475 (N_8475,N_6606,N_6441);
and U8476 (N_8476,N_7031,N_6315);
xor U8477 (N_8477,N_7091,N_6841);
xnor U8478 (N_8478,N_7330,N_7179);
nor U8479 (N_8479,N_6832,N_7333);
nor U8480 (N_8480,N_7423,N_7264);
and U8481 (N_8481,N_7098,N_7017);
nor U8482 (N_8482,N_6814,N_7432);
and U8483 (N_8483,N_6477,N_7055);
and U8484 (N_8484,N_6391,N_6502);
and U8485 (N_8485,N_6594,N_7292);
nor U8486 (N_8486,N_7402,N_6930);
xnor U8487 (N_8487,N_6651,N_7489);
or U8488 (N_8488,N_7051,N_6655);
nor U8489 (N_8489,N_6524,N_6435);
xor U8490 (N_8490,N_6789,N_7122);
and U8491 (N_8491,N_7060,N_7422);
xnor U8492 (N_8492,N_7471,N_7123);
xor U8493 (N_8493,N_7027,N_7313);
or U8494 (N_8494,N_6793,N_6401);
xnor U8495 (N_8495,N_6592,N_6740);
xnor U8496 (N_8496,N_7422,N_7406);
and U8497 (N_8497,N_6768,N_6625);
or U8498 (N_8498,N_6282,N_7451);
nand U8499 (N_8499,N_7495,N_7017);
and U8500 (N_8500,N_7370,N_6609);
nor U8501 (N_8501,N_6628,N_6478);
or U8502 (N_8502,N_7280,N_7232);
and U8503 (N_8503,N_7267,N_6376);
or U8504 (N_8504,N_7198,N_6761);
and U8505 (N_8505,N_6350,N_7381);
xnor U8506 (N_8506,N_7055,N_6623);
xnor U8507 (N_8507,N_6685,N_6956);
and U8508 (N_8508,N_6578,N_7076);
nand U8509 (N_8509,N_7115,N_6611);
and U8510 (N_8510,N_7425,N_6432);
and U8511 (N_8511,N_7008,N_6872);
and U8512 (N_8512,N_7333,N_7335);
nor U8513 (N_8513,N_6611,N_6736);
xor U8514 (N_8514,N_6853,N_6662);
nand U8515 (N_8515,N_6267,N_6549);
and U8516 (N_8516,N_7087,N_6535);
nand U8517 (N_8517,N_6876,N_6603);
nor U8518 (N_8518,N_7307,N_7390);
and U8519 (N_8519,N_7349,N_6405);
or U8520 (N_8520,N_7008,N_7436);
xnor U8521 (N_8521,N_7199,N_6465);
xnor U8522 (N_8522,N_6434,N_6334);
and U8523 (N_8523,N_7181,N_7259);
or U8524 (N_8524,N_7329,N_6676);
or U8525 (N_8525,N_6661,N_6322);
xor U8526 (N_8526,N_6493,N_7225);
nand U8527 (N_8527,N_7225,N_6533);
and U8528 (N_8528,N_7293,N_7301);
and U8529 (N_8529,N_7078,N_7396);
nand U8530 (N_8530,N_7000,N_7061);
xor U8531 (N_8531,N_7186,N_7408);
and U8532 (N_8532,N_7002,N_6699);
or U8533 (N_8533,N_7286,N_6858);
nand U8534 (N_8534,N_7334,N_6744);
and U8535 (N_8535,N_6337,N_7036);
or U8536 (N_8536,N_7272,N_6417);
or U8537 (N_8537,N_6414,N_7289);
nand U8538 (N_8538,N_6534,N_7009);
nor U8539 (N_8539,N_6914,N_6862);
nor U8540 (N_8540,N_6611,N_6629);
nor U8541 (N_8541,N_7224,N_6606);
or U8542 (N_8542,N_6903,N_6358);
nand U8543 (N_8543,N_7199,N_7371);
xnor U8544 (N_8544,N_6511,N_6741);
and U8545 (N_8545,N_6889,N_7200);
and U8546 (N_8546,N_7454,N_7474);
or U8547 (N_8547,N_7468,N_6966);
xor U8548 (N_8548,N_6720,N_6726);
or U8549 (N_8549,N_7108,N_6934);
or U8550 (N_8550,N_6647,N_6594);
nor U8551 (N_8551,N_6476,N_7319);
nand U8552 (N_8552,N_7487,N_6308);
xnor U8553 (N_8553,N_6506,N_7094);
nor U8554 (N_8554,N_7182,N_6749);
nand U8555 (N_8555,N_6790,N_6669);
xor U8556 (N_8556,N_7159,N_6490);
or U8557 (N_8557,N_6668,N_7423);
xnor U8558 (N_8558,N_7112,N_6426);
or U8559 (N_8559,N_6293,N_6302);
nand U8560 (N_8560,N_6430,N_6631);
nor U8561 (N_8561,N_7159,N_6681);
and U8562 (N_8562,N_7187,N_6491);
or U8563 (N_8563,N_6849,N_6861);
and U8564 (N_8564,N_6281,N_6886);
nor U8565 (N_8565,N_6453,N_6336);
or U8566 (N_8566,N_6310,N_7199);
nor U8567 (N_8567,N_6928,N_7246);
nor U8568 (N_8568,N_6996,N_6990);
or U8569 (N_8569,N_6383,N_7200);
xnor U8570 (N_8570,N_6439,N_7223);
or U8571 (N_8571,N_7457,N_6832);
nor U8572 (N_8572,N_7221,N_6681);
and U8573 (N_8573,N_6942,N_6851);
or U8574 (N_8574,N_6576,N_6693);
nor U8575 (N_8575,N_7299,N_6343);
nor U8576 (N_8576,N_6337,N_6860);
nand U8577 (N_8577,N_6441,N_6683);
xnor U8578 (N_8578,N_7104,N_6346);
or U8579 (N_8579,N_6662,N_7284);
and U8580 (N_8580,N_6783,N_7383);
or U8581 (N_8581,N_7267,N_6974);
nand U8582 (N_8582,N_6332,N_6702);
nand U8583 (N_8583,N_7399,N_6260);
and U8584 (N_8584,N_7322,N_6622);
xnor U8585 (N_8585,N_6703,N_6613);
and U8586 (N_8586,N_6349,N_6995);
and U8587 (N_8587,N_6929,N_7493);
nor U8588 (N_8588,N_6787,N_7450);
nor U8589 (N_8589,N_7208,N_6649);
nand U8590 (N_8590,N_7443,N_6567);
nor U8591 (N_8591,N_6339,N_7027);
nand U8592 (N_8592,N_7381,N_7251);
or U8593 (N_8593,N_7453,N_7202);
nor U8594 (N_8594,N_7305,N_6817);
nand U8595 (N_8595,N_7407,N_7483);
nand U8596 (N_8596,N_7315,N_7382);
or U8597 (N_8597,N_6410,N_6512);
xnor U8598 (N_8598,N_6619,N_7188);
nand U8599 (N_8599,N_6472,N_7013);
and U8600 (N_8600,N_6864,N_7051);
nand U8601 (N_8601,N_6315,N_7483);
or U8602 (N_8602,N_6757,N_7311);
or U8603 (N_8603,N_6955,N_7085);
xnor U8604 (N_8604,N_6385,N_6638);
and U8605 (N_8605,N_7210,N_7291);
nand U8606 (N_8606,N_6577,N_6767);
and U8607 (N_8607,N_7031,N_6645);
nand U8608 (N_8608,N_6977,N_6333);
nor U8609 (N_8609,N_6572,N_6331);
and U8610 (N_8610,N_6354,N_7041);
nand U8611 (N_8611,N_7075,N_7384);
nand U8612 (N_8612,N_6606,N_7168);
nor U8613 (N_8613,N_7166,N_6939);
xnor U8614 (N_8614,N_6563,N_7282);
xnor U8615 (N_8615,N_6797,N_6610);
xor U8616 (N_8616,N_7499,N_6690);
or U8617 (N_8617,N_6848,N_6850);
or U8618 (N_8618,N_7104,N_7289);
or U8619 (N_8619,N_6408,N_7436);
xor U8620 (N_8620,N_6903,N_6652);
xor U8621 (N_8621,N_7395,N_7457);
xor U8622 (N_8622,N_6281,N_6816);
or U8623 (N_8623,N_6432,N_6463);
and U8624 (N_8624,N_6506,N_7471);
xor U8625 (N_8625,N_6846,N_6598);
and U8626 (N_8626,N_7338,N_6301);
nand U8627 (N_8627,N_6776,N_6570);
and U8628 (N_8628,N_7284,N_6439);
or U8629 (N_8629,N_6310,N_6639);
or U8630 (N_8630,N_7412,N_6793);
and U8631 (N_8631,N_6812,N_6331);
or U8632 (N_8632,N_6911,N_6496);
xor U8633 (N_8633,N_6486,N_6572);
nor U8634 (N_8634,N_6678,N_7484);
nor U8635 (N_8635,N_6863,N_7313);
or U8636 (N_8636,N_7165,N_6419);
xnor U8637 (N_8637,N_7467,N_6361);
or U8638 (N_8638,N_7470,N_6937);
and U8639 (N_8639,N_6956,N_6728);
xnor U8640 (N_8640,N_6593,N_6375);
xnor U8641 (N_8641,N_6440,N_7023);
nand U8642 (N_8642,N_6331,N_6946);
and U8643 (N_8643,N_6515,N_7445);
or U8644 (N_8644,N_7097,N_6925);
nor U8645 (N_8645,N_6583,N_6434);
xor U8646 (N_8646,N_7129,N_7362);
nand U8647 (N_8647,N_6847,N_6334);
xor U8648 (N_8648,N_7399,N_6445);
nand U8649 (N_8649,N_6421,N_6996);
and U8650 (N_8650,N_7394,N_7170);
and U8651 (N_8651,N_6651,N_6809);
and U8652 (N_8652,N_6898,N_6799);
nor U8653 (N_8653,N_6588,N_6896);
nand U8654 (N_8654,N_6337,N_6398);
nand U8655 (N_8655,N_6970,N_7381);
nand U8656 (N_8656,N_6380,N_6539);
or U8657 (N_8657,N_7487,N_7239);
xor U8658 (N_8658,N_7335,N_6704);
xnor U8659 (N_8659,N_6741,N_7094);
xnor U8660 (N_8660,N_7437,N_7317);
or U8661 (N_8661,N_6661,N_7463);
xor U8662 (N_8662,N_6562,N_7360);
nor U8663 (N_8663,N_7497,N_6997);
nor U8664 (N_8664,N_6870,N_6583);
and U8665 (N_8665,N_7406,N_7281);
nor U8666 (N_8666,N_6980,N_6476);
nand U8667 (N_8667,N_6960,N_7187);
or U8668 (N_8668,N_7084,N_6250);
xnor U8669 (N_8669,N_7476,N_6855);
or U8670 (N_8670,N_6641,N_6618);
nor U8671 (N_8671,N_6693,N_7453);
nor U8672 (N_8672,N_6885,N_6777);
and U8673 (N_8673,N_7267,N_7239);
or U8674 (N_8674,N_6853,N_6426);
nand U8675 (N_8675,N_7125,N_6728);
xnor U8676 (N_8676,N_6475,N_6812);
nand U8677 (N_8677,N_7203,N_6500);
nand U8678 (N_8678,N_6541,N_7332);
and U8679 (N_8679,N_6985,N_6567);
nor U8680 (N_8680,N_6612,N_7098);
and U8681 (N_8681,N_7431,N_6454);
xor U8682 (N_8682,N_6784,N_7140);
or U8683 (N_8683,N_6804,N_6475);
and U8684 (N_8684,N_6961,N_6640);
or U8685 (N_8685,N_7485,N_6898);
nand U8686 (N_8686,N_6920,N_7418);
xor U8687 (N_8687,N_6437,N_6732);
nor U8688 (N_8688,N_6700,N_6934);
or U8689 (N_8689,N_6825,N_6362);
xor U8690 (N_8690,N_6938,N_6656);
nand U8691 (N_8691,N_7343,N_6341);
or U8692 (N_8692,N_6479,N_6444);
nor U8693 (N_8693,N_7116,N_7029);
xor U8694 (N_8694,N_7080,N_6720);
or U8695 (N_8695,N_6505,N_6275);
nand U8696 (N_8696,N_7458,N_6697);
xor U8697 (N_8697,N_7309,N_6775);
or U8698 (N_8698,N_6498,N_6747);
nor U8699 (N_8699,N_7337,N_6810);
or U8700 (N_8700,N_6516,N_7241);
nand U8701 (N_8701,N_6829,N_7240);
nand U8702 (N_8702,N_7344,N_6833);
xor U8703 (N_8703,N_7426,N_6433);
nor U8704 (N_8704,N_7445,N_6767);
and U8705 (N_8705,N_7305,N_7096);
and U8706 (N_8706,N_6370,N_6782);
xor U8707 (N_8707,N_6424,N_6378);
and U8708 (N_8708,N_6730,N_6427);
nand U8709 (N_8709,N_7426,N_6600);
nor U8710 (N_8710,N_6377,N_6750);
or U8711 (N_8711,N_7434,N_6836);
xnor U8712 (N_8712,N_7080,N_6613);
or U8713 (N_8713,N_7447,N_7039);
and U8714 (N_8714,N_6713,N_6577);
nand U8715 (N_8715,N_7415,N_7426);
and U8716 (N_8716,N_7066,N_7238);
xor U8717 (N_8717,N_7153,N_7435);
or U8718 (N_8718,N_6316,N_6277);
xnor U8719 (N_8719,N_7278,N_7295);
or U8720 (N_8720,N_7041,N_7140);
nor U8721 (N_8721,N_7118,N_7356);
or U8722 (N_8722,N_6999,N_6309);
or U8723 (N_8723,N_6538,N_6832);
nor U8724 (N_8724,N_7499,N_7101);
and U8725 (N_8725,N_6841,N_6628);
or U8726 (N_8726,N_6391,N_6787);
or U8727 (N_8727,N_7358,N_6958);
nand U8728 (N_8728,N_6835,N_6330);
or U8729 (N_8729,N_6586,N_6426);
and U8730 (N_8730,N_6311,N_7122);
and U8731 (N_8731,N_7463,N_7464);
xor U8732 (N_8732,N_6887,N_6953);
and U8733 (N_8733,N_7292,N_7043);
xnor U8734 (N_8734,N_6574,N_6470);
or U8735 (N_8735,N_7359,N_6640);
and U8736 (N_8736,N_7430,N_6689);
nand U8737 (N_8737,N_7395,N_6369);
nand U8738 (N_8738,N_7148,N_6690);
or U8739 (N_8739,N_7184,N_6264);
or U8740 (N_8740,N_7078,N_6320);
and U8741 (N_8741,N_6957,N_6881);
or U8742 (N_8742,N_7076,N_6620);
xnor U8743 (N_8743,N_6974,N_7350);
and U8744 (N_8744,N_6470,N_7419);
nand U8745 (N_8745,N_7431,N_6469);
nor U8746 (N_8746,N_7283,N_7335);
or U8747 (N_8747,N_6552,N_6975);
nand U8748 (N_8748,N_7054,N_6878);
and U8749 (N_8749,N_6796,N_6325);
nand U8750 (N_8750,N_7688,N_8113);
nor U8751 (N_8751,N_8746,N_8524);
nand U8752 (N_8752,N_8387,N_8470);
xor U8753 (N_8753,N_8529,N_8189);
nand U8754 (N_8754,N_7666,N_8336);
nand U8755 (N_8755,N_8303,N_8504);
nor U8756 (N_8756,N_8543,N_7903);
nand U8757 (N_8757,N_8466,N_8196);
xor U8758 (N_8758,N_8489,N_7714);
and U8759 (N_8759,N_8660,N_8555);
or U8760 (N_8760,N_7799,N_8464);
and U8761 (N_8761,N_8241,N_8662);
nor U8762 (N_8762,N_8256,N_7588);
nor U8763 (N_8763,N_8187,N_8618);
nor U8764 (N_8764,N_7732,N_8418);
xor U8765 (N_8765,N_8063,N_8348);
and U8766 (N_8766,N_7633,N_8652);
xnor U8767 (N_8767,N_8337,N_8683);
and U8768 (N_8768,N_8086,N_8133);
xor U8769 (N_8769,N_8078,N_7820);
and U8770 (N_8770,N_8526,N_7758);
or U8771 (N_8771,N_8162,N_8095);
nor U8772 (N_8772,N_8321,N_7505);
xnor U8773 (N_8773,N_8048,N_7961);
or U8774 (N_8774,N_7899,N_8075);
or U8775 (N_8775,N_8147,N_8592);
nand U8776 (N_8776,N_7625,N_7509);
nand U8777 (N_8777,N_7719,N_8460);
xor U8778 (N_8778,N_7839,N_7811);
nand U8779 (N_8779,N_7773,N_7819);
and U8780 (N_8780,N_7703,N_8422);
nand U8781 (N_8781,N_8567,N_8476);
and U8782 (N_8782,N_7927,N_7574);
and U8783 (N_8783,N_8545,N_8277);
nand U8784 (N_8784,N_8223,N_8663);
or U8785 (N_8785,N_7868,N_7896);
nand U8786 (N_8786,N_7947,N_7645);
nor U8787 (N_8787,N_8602,N_8339);
nor U8788 (N_8788,N_8508,N_7988);
nand U8789 (N_8789,N_8289,N_7965);
and U8790 (N_8790,N_7523,N_7715);
nor U8791 (N_8791,N_8010,N_7668);
nor U8792 (N_8792,N_8395,N_8428);
nor U8793 (N_8793,N_8064,N_8347);
nor U8794 (N_8794,N_8188,N_8326);
nand U8795 (N_8795,N_7849,N_8116);
and U8796 (N_8796,N_7545,N_8722);
or U8797 (N_8797,N_7829,N_8157);
xor U8798 (N_8798,N_7952,N_8194);
xnor U8799 (N_8799,N_8186,N_7731);
or U8800 (N_8800,N_7838,N_7913);
nor U8801 (N_8801,N_8017,N_8364);
xor U8802 (N_8802,N_8169,N_7759);
or U8803 (N_8803,N_8546,N_8203);
xor U8804 (N_8804,N_8222,N_7966);
or U8805 (N_8805,N_7806,N_7689);
xnor U8806 (N_8806,N_8741,N_8003);
nand U8807 (N_8807,N_8340,N_8153);
or U8808 (N_8808,N_8518,N_7904);
nand U8809 (N_8809,N_8324,N_8624);
or U8810 (N_8810,N_8513,N_7590);
and U8811 (N_8811,N_8570,N_8512);
xnor U8812 (N_8812,N_8502,N_8425);
and U8813 (N_8813,N_7814,N_8630);
nand U8814 (N_8814,N_8184,N_8376);
xor U8815 (N_8815,N_7608,N_8148);
nor U8816 (N_8816,N_8439,N_8060);
nand U8817 (N_8817,N_7857,N_8329);
nor U8818 (N_8818,N_8552,N_8551);
nor U8819 (N_8819,N_7748,N_8354);
or U8820 (N_8820,N_8454,N_8380);
or U8821 (N_8821,N_8608,N_8150);
or U8822 (N_8822,N_8311,N_8572);
nor U8823 (N_8823,N_8028,N_8485);
or U8824 (N_8824,N_8463,N_8441);
and U8825 (N_8825,N_8645,N_7907);
nor U8826 (N_8826,N_7976,N_7746);
nand U8827 (N_8827,N_7848,N_8007);
nor U8828 (N_8828,N_8357,N_8604);
nand U8829 (N_8829,N_7978,N_8295);
nand U8830 (N_8830,N_8175,N_7793);
or U8831 (N_8831,N_7824,N_8469);
and U8832 (N_8832,N_7716,N_8310);
nor U8833 (N_8833,N_7891,N_7541);
or U8834 (N_8834,N_8414,N_7805);
nor U8835 (N_8835,N_7835,N_7556);
nand U8836 (N_8836,N_8688,N_7999);
nand U8837 (N_8837,N_7932,N_7885);
and U8838 (N_8838,N_7971,N_8548);
nand U8839 (N_8839,N_8163,N_7612);
nor U8840 (N_8840,N_8655,N_8675);
xor U8841 (N_8841,N_7882,N_8609);
and U8842 (N_8842,N_8250,N_8114);
nand U8843 (N_8843,N_7677,N_8069);
nor U8844 (N_8844,N_8043,N_8294);
and U8845 (N_8845,N_8573,N_7636);
nand U8846 (N_8846,N_7985,N_7935);
xor U8847 (N_8847,N_7524,N_8495);
nor U8848 (N_8848,N_8005,N_7513);
nor U8849 (N_8849,N_7867,N_7699);
or U8850 (N_8850,N_8192,N_7775);
nor U8851 (N_8851,N_7836,N_8229);
and U8852 (N_8852,N_8083,N_7963);
nand U8853 (N_8853,N_7660,N_7841);
xnor U8854 (N_8854,N_8183,N_7765);
nor U8855 (N_8855,N_7621,N_7946);
xnor U8856 (N_8856,N_7776,N_7847);
or U8857 (N_8857,N_8238,N_8651);
nor U8858 (N_8858,N_8103,N_8316);
nor U8859 (N_8859,N_7506,N_8656);
nor U8860 (N_8860,N_8381,N_8047);
or U8861 (N_8861,N_7928,N_8450);
and U8862 (N_8862,N_8059,N_8534);
or U8863 (N_8863,N_8230,N_7661);
nand U8864 (N_8864,N_8459,N_8491);
nand U8865 (N_8865,N_8237,N_8542);
and U8866 (N_8866,N_8653,N_8676);
or U8867 (N_8867,N_7603,N_7628);
xnor U8868 (N_8868,N_7834,N_7830);
nand U8869 (N_8869,N_8701,N_7649);
and U8870 (N_8870,N_8374,N_8699);
xor U8871 (N_8871,N_8506,N_7914);
nor U8872 (N_8872,N_7873,N_8168);
and U8873 (N_8873,N_8525,N_8115);
and U8874 (N_8874,N_7630,N_8536);
nor U8875 (N_8875,N_7831,N_8367);
or U8876 (N_8876,N_8234,N_8023);
or U8877 (N_8877,N_8293,N_8700);
xnor U8878 (N_8878,N_8094,N_8679);
nand U8879 (N_8879,N_8343,N_7722);
or U8880 (N_8880,N_8338,N_7727);
nand U8881 (N_8881,N_7774,N_8711);
nand U8882 (N_8882,N_7926,N_7990);
or U8883 (N_8883,N_7631,N_8145);
nor U8884 (N_8884,N_8334,N_8671);
xnor U8885 (N_8885,N_8008,N_8360);
nand U8886 (N_8886,N_7723,N_8472);
nor U8887 (N_8887,N_7797,N_8614);
nor U8888 (N_8888,N_8386,N_7655);
nor U8889 (N_8889,N_7557,N_8549);
xor U8890 (N_8890,N_8582,N_7742);
or U8891 (N_8891,N_8102,N_8134);
or U8892 (N_8892,N_8280,N_7972);
xor U8893 (N_8893,N_8680,N_8693);
xor U8894 (N_8894,N_7786,N_7718);
nand U8895 (N_8895,N_7702,N_8452);
xor U8896 (N_8896,N_8071,N_8607);
or U8897 (N_8897,N_7500,N_7665);
and U8898 (N_8898,N_8649,N_8268);
or U8899 (N_8899,N_8461,N_8319);
nand U8900 (N_8900,N_8687,N_7686);
nor U8901 (N_8901,N_7578,N_8279);
nor U8902 (N_8902,N_8274,N_7547);
nand U8903 (N_8903,N_8253,N_7683);
and U8904 (N_8904,N_7510,N_8097);
or U8905 (N_8905,N_8317,N_8217);
and U8906 (N_8906,N_8022,N_7890);
or U8907 (N_8907,N_8120,N_8053);
or U8908 (N_8908,N_7991,N_8174);
and U8909 (N_8909,N_8382,N_8181);
nand U8910 (N_8910,N_7512,N_7568);
and U8911 (N_8911,N_8409,N_8715);
nand U8912 (N_8912,N_8080,N_7794);
or U8913 (N_8913,N_8696,N_8718);
or U8914 (N_8914,N_8691,N_7530);
or U8915 (N_8915,N_7700,N_8642);
nand U8916 (N_8916,N_7817,N_8226);
nand U8917 (N_8917,N_8666,N_7583);
xor U8918 (N_8918,N_8659,N_7733);
nor U8919 (N_8919,N_8131,N_7606);
and U8920 (N_8920,N_8308,N_8510);
nand U8921 (N_8921,N_7930,N_8532);
xnor U8922 (N_8922,N_8569,N_7860);
nor U8923 (N_8923,N_7651,N_8503);
xnor U8924 (N_8924,N_7987,N_7949);
or U8925 (N_8925,N_8323,N_8039);
or U8926 (N_8926,N_7535,N_8559);
or U8927 (N_8927,N_8202,N_8352);
and U8928 (N_8928,N_8623,N_7771);
nor U8929 (N_8929,N_7735,N_7642);
nand U8930 (N_8930,N_8378,N_8051);
xnor U8931 (N_8931,N_8541,N_7532);
or U8932 (N_8932,N_8037,N_7669);
and U8933 (N_8933,N_7975,N_8458);
and U8934 (N_8934,N_7560,N_8389);
or U8935 (N_8935,N_7923,N_7752);
xnor U8936 (N_8936,N_8456,N_8578);
and U8937 (N_8937,N_7878,N_8695);
or U8938 (N_8938,N_8499,N_7825);
and U8939 (N_8939,N_7865,N_8694);
nor U8940 (N_8940,N_8304,N_7508);
xor U8941 (N_8941,N_8090,N_8739);
xnor U8942 (N_8942,N_8365,N_7922);
nand U8943 (N_8943,N_7717,N_7537);
nand U8944 (N_8944,N_7569,N_8706);
nor U8945 (N_8945,N_7581,N_8014);
and U8946 (N_8946,N_8519,N_8285);
and U8947 (N_8947,N_8180,N_8550);
nor U8948 (N_8948,N_7682,N_8435);
and U8949 (N_8949,N_8408,N_8533);
nor U8950 (N_8950,N_7837,N_7840);
nand U8951 (N_8951,N_8021,N_7821);
xnor U8952 (N_8952,N_7685,N_7692);
nor U8953 (N_8953,N_8266,N_7983);
or U8954 (N_8954,N_8528,N_8099);
and U8955 (N_8955,N_8209,N_8032);
or U8956 (N_8956,N_7909,N_7981);
or U8957 (N_8957,N_8346,N_7720);
and U8958 (N_8958,N_7519,N_7802);
nand U8959 (N_8959,N_7626,N_8641);
xnor U8960 (N_8960,N_7772,N_7851);
nand U8961 (N_8961,N_7609,N_7943);
nand U8962 (N_8962,N_8646,N_8644);
and U8963 (N_8963,N_7667,N_7889);
nor U8964 (N_8964,N_7536,N_7933);
nor U8965 (N_8965,N_7542,N_7833);
or U8966 (N_8966,N_8149,N_7577);
or U8967 (N_8967,N_7763,N_7747);
or U8968 (N_8968,N_7529,N_8391);
nand U8969 (N_8969,N_8027,N_7623);
and U8970 (N_8970,N_8333,N_8611);
and U8971 (N_8971,N_8605,N_7595);
or U8972 (N_8972,N_7740,N_7599);
nand U8973 (N_8973,N_8584,N_7950);
nand U8974 (N_8974,N_8400,N_8399);
nor U8975 (N_8975,N_8024,N_7916);
nand U8976 (N_8976,N_8061,N_8154);
and U8977 (N_8977,N_8057,N_8239);
nand U8978 (N_8978,N_7571,N_8554);
xnor U8979 (N_8979,N_8588,N_8708);
or U8980 (N_8980,N_7613,N_7969);
or U8981 (N_8981,N_8235,N_8204);
or U8982 (N_8982,N_7711,N_7974);
or U8983 (N_8983,N_7902,N_7812);
or U8984 (N_8984,N_8073,N_7673);
xor U8985 (N_8985,N_7934,N_8105);
nand U8986 (N_8986,N_7610,N_8233);
and U8987 (N_8987,N_8451,N_8509);
nand U8988 (N_8988,N_8366,N_7550);
or U8989 (N_8989,N_7596,N_8232);
and U8990 (N_8990,N_8433,N_7931);
or U8991 (N_8991,N_8521,N_8434);
or U8992 (N_8992,N_7687,N_7526);
or U8993 (N_8993,N_8088,N_7944);
and U8994 (N_8994,N_7910,N_8001);
xnor U8995 (N_8995,N_8544,N_7770);
nor U8996 (N_8996,N_8138,N_8132);
and U8997 (N_8997,N_7887,N_7901);
xor U8998 (N_8998,N_8261,N_8299);
nor U8999 (N_8999,N_8026,N_8698);
nor U9000 (N_9000,N_8568,N_7850);
xor U9001 (N_9001,N_7982,N_7518);
nor U9002 (N_9002,N_7869,N_7852);
nand U9003 (N_9003,N_7657,N_8595);
xnor U9004 (N_9004,N_8212,N_8396);
nor U9005 (N_9005,N_8394,N_8634);
nand U9006 (N_9006,N_8298,N_8457);
nand U9007 (N_9007,N_7604,N_8488);
nor U9008 (N_9008,N_7632,N_8054);
and U9009 (N_9009,N_8328,N_8004);
nand U9010 (N_9010,N_8580,N_8446);
xor U9011 (N_9011,N_8402,N_7984);
xnor U9012 (N_9012,N_8585,N_7582);
nand U9013 (N_9013,N_7784,N_7664);
and U9014 (N_9014,N_8437,N_8723);
xnor U9015 (N_9015,N_7807,N_7548);
nand U9016 (N_9016,N_7941,N_8633);
nand U9017 (N_9017,N_8717,N_8193);
nor U9018 (N_9018,N_8487,N_8537);
nor U9019 (N_9019,N_8709,N_7729);
and U9020 (N_9020,N_8377,N_8330);
and U9021 (N_9021,N_8412,N_7674);
or U9022 (N_9022,N_7895,N_8142);
nor U9023 (N_9023,N_7912,N_8052);
xnor U9024 (N_9024,N_8426,N_7622);
or U9025 (N_9025,N_8140,N_8714);
xnor U9026 (N_9026,N_7921,N_8379);
nor U9027 (N_9027,N_7945,N_8164);
or U9028 (N_9028,N_8036,N_8496);
or U9029 (N_9029,N_8689,N_8690);
xnor U9030 (N_9030,N_7955,N_8242);
and U9031 (N_9031,N_8144,N_8259);
nor U9032 (N_9032,N_7862,N_7940);
or U9033 (N_9033,N_7875,N_8015);
nor U9034 (N_9034,N_7798,N_8190);
or U9035 (N_9035,N_7705,N_8109);
nand U9036 (N_9036,N_7566,N_8678);
or U9037 (N_9037,N_7757,N_8411);
xnor U9038 (N_9038,N_8031,N_7691);
xnor U9039 (N_9039,N_8287,N_8449);
nand U9040 (N_9040,N_7654,N_8087);
and U9041 (N_9041,N_8249,N_8341);
or U9042 (N_9042,N_8535,N_8221);
or U9043 (N_9043,N_8597,N_8076);
nor U9044 (N_9044,N_8166,N_8284);
nor U9045 (N_9045,N_8020,N_7652);
xor U9046 (N_9046,N_8443,N_7874);
and U9047 (N_9047,N_8269,N_7809);
xor U9048 (N_9048,N_8273,N_7618);
nor U9049 (N_9049,N_8483,N_8479);
and U9050 (N_9050,N_8553,N_7501);
nand U9051 (N_9051,N_8123,N_8514);
nand U9052 (N_9052,N_7905,N_7779);
nor U9053 (N_9053,N_8351,N_8098);
nor U9054 (N_9054,N_8161,N_7639);
xnor U9055 (N_9055,N_8122,N_8356);
nand U9056 (N_9056,N_8079,N_8359);
and U9057 (N_9057,N_8719,N_7832);
and U9058 (N_9058,N_8306,N_8478);
xor U9059 (N_9059,N_7602,N_8282);
and U9060 (N_9060,N_8598,N_8658);
nor U9061 (N_9061,N_8564,N_8267);
and U9062 (N_9062,N_7866,N_7813);
and U9063 (N_9063,N_8068,N_8118);
nor U9064 (N_9064,N_8639,N_8480);
or U9065 (N_9065,N_7521,N_7533);
or U9066 (N_9066,N_8093,N_7822);
xnor U9067 (N_9067,N_7884,N_8225);
nand U9068 (N_9068,N_8013,N_8558);
and U9069 (N_9069,N_8160,N_8342);
or U9070 (N_9070,N_8523,N_8601);
or U9071 (N_9071,N_8596,N_8254);
and U9072 (N_9072,N_8406,N_8141);
and U9073 (N_9073,N_7531,N_7743);
and U9074 (N_9074,N_8170,N_8471);
xor U9075 (N_9075,N_8576,N_8072);
nor U9076 (N_9076,N_8029,N_8107);
nor U9077 (N_9077,N_7561,N_8587);
and U9078 (N_9078,N_7540,N_8600);
xor U9079 (N_9079,N_8628,N_7894);
nor U9080 (N_9080,N_7650,N_7724);
or U9081 (N_9081,N_7803,N_8643);
and U9082 (N_9082,N_8302,N_8668);
nor U9083 (N_9083,N_7515,N_8673);
nand U9084 (N_9084,N_7730,N_8627);
and U9085 (N_9085,N_7964,N_8345);
nor U9086 (N_9086,N_8527,N_7788);
nor U9087 (N_9087,N_8473,N_8165);
nand U9088 (N_9088,N_8650,N_8501);
or U9089 (N_9089,N_8091,N_7783);
or U9090 (N_9090,N_8415,N_7695);
xor U9091 (N_9091,N_8677,N_7953);
and U9092 (N_9092,N_8251,N_8156);
nor U9093 (N_9093,N_7843,N_8146);
nand U9094 (N_9094,N_7768,N_7614);
nand U9095 (N_9095,N_7995,N_8125);
and U9096 (N_9096,N_7883,N_8665);
nor U9097 (N_9097,N_8176,N_7973);
nand U9098 (N_9098,N_8286,N_8388);
xor U9099 (N_9099,N_7967,N_7681);
nor U9100 (N_9100,N_8724,N_8486);
nor U9101 (N_9101,N_8240,N_8368);
or U9102 (N_9102,N_7565,N_7968);
nand U9103 (N_9103,N_8583,N_7777);
xor U9104 (N_9104,N_8208,N_8127);
or U9105 (N_9105,N_8197,N_8331);
or U9106 (N_9106,N_7787,N_7977);
nor U9107 (N_9107,N_7864,N_8077);
or U9108 (N_9108,N_8151,N_8228);
nand U9109 (N_9109,N_8562,N_7637);
nor U9110 (N_9110,N_8561,N_7801);
or U9111 (N_9111,N_8255,N_8297);
and U9112 (N_9112,N_8684,N_7853);
nor U9113 (N_9113,N_7906,N_8124);
and U9114 (N_9114,N_8016,N_7888);
nand U9115 (N_9115,N_8500,N_8704);
nor U9116 (N_9116,N_7816,N_8729);
nor U9117 (N_9117,N_8565,N_7791);
nand U9118 (N_9118,N_7611,N_7552);
xnor U9119 (N_9119,N_8713,N_8742);
or U9120 (N_9120,N_8231,N_8637);
nor U9121 (N_9121,N_7992,N_8421);
and U9122 (N_9122,N_7620,N_8246);
nand U9123 (N_9123,N_8350,N_8465);
nand U9124 (N_9124,N_7886,N_8200);
or U9125 (N_9125,N_7881,N_7517);
nand U9126 (N_9126,N_7781,N_8405);
nor U9127 (N_9127,N_8030,N_7855);
or U9128 (N_9128,N_7744,N_8362);
nor U9129 (N_9129,N_8258,N_7607);
nand U9130 (N_9130,N_8272,N_8606);
or U9131 (N_9131,N_8292,N_7854);
xor U9132 (N_9132,N_8332,N_7929);
xor U9133 (N_9133,N_7948,N_8593);
nand U9134 (N_9134,N_7994,N_7710);
nor U9135 (N_9135,N_8011,N_7551);
and U9136 (N_9136,N_7584,N_8248);
xnor U9137 (N_9137,N_7956,N_8427);
nand U9138 (N_9138,N_7647,N_7725);
nor U9139 (N_9139,N_8590,N_8490);
and U9140 (N_9140,N_8737,N_7876);
or U9141 (N_9141,N_8516,N_7564);
nor U9142 (N_9142,N_7616,N_7586);
or U9143 (N_9143,N_8511,N_7957);
xnor U9144 (N_9144,N_8372,N_8625);
and U9145 (N_9145,N_8135,N_8444);
nand U9146 (N_9146,N_8557,N_7958);
xnor U9147 (N_9147,N_8358,N_7514);
nor U9148 (N_9148,N_8577,N_7919);
nor U9149 (N_9149,N_8620,N_8686);
xor U9150 (N_9150,N_7589,N_7576);
nand U9151 (N_9151,N_7960,N_7741);
xnor U9152 (N_9152,N_8111,N_8661);
and U9153 (N_9153,N_8244,N_7549);
and U9154 (N_9154,N_8455,N_7738);
nand U9155 (N_9155,N_8617,N_8738);
or U9156 (N_9156,N_8104,N_7562);
or U9157 (N_9157,N_8000,N_7755);
or U9158 (N_9158,N_8615,N_8089);
xnor U9159 (N_9159,N_8445,N_8494);
and U9160 (N_9160,N_8171,N_7892);
nor U9161 (N_9161,N_8591,N_7917);
xor U9162 (N_9162,N_8664,N_7936);
and U9163 (N_9163,N_8301,N_8440);
and U9164 (N_9164,N_8172,N_8305);
nor U9165 (N_9165,N_8227,N_8058);
nand U9166 (N_9166,N_8447,N_7846);
or U9167 (N_9167,N_8744,N_8220);
nand U9168 (N_9168,N_7749,N_7646);
xor U9169 (N_9169,N_8370,N_8419);
or U9170 (N_9170,N_8081,N_8397);
nand U9171 (N_9171,N_7638,N_8199);
xnor U9172 (N_9172,N_7546,N_7684);
and U9173 (N_9173,N_7736,N_7827);
nand U9174 (N_9174,N_8626,N_7810);
and U9175 (N_9175,N_8622,N_8117);
nand U9176 (N_9176,N_8074,N_7893);
xor U9177 (N_9177,N_8100,N_7962);
xor U9178 (N_9178,N_7789,N_8672);
nor U9179 (N_9179,N_8278,N_7754);
nor U9180 (N_9180,N_7558,N_8385);
or U9181 (N_9181,N_8106,N_8401);
nand U9182 (N_9182,N_7572,N_8477);
or U9183 (N_9183,N_8312,N_8355);
xor U9184 (N_9184,N_7575,N_8575);
nand U9185 (N_9185,N_8291,N_8264);
or U9186 (N_9186,N_8727,N_7503);
nor U9187 (N_9187,N_7567,N_8670);
nor U9188 (N_9188,N_8353,N_7823);
xor U9189 (N_9189,N_8314,N_8056);
or U9190 (N_9190,N_8185,N_8398);
and U9191 (N_9191,N_7863,N_8685);
and U9192 (N_9192,N_7861,N_7538);
nor U9193 (N_9193,N_7998,N_7653);
xnor U9194 (N_9194,N_8726,N_8647);
nand U9195 (N_9195,N_8619,N_8621);
nor U9196 (N_9196,N_7959,N_8044);
nand U9197 (N_9197,N_7658,N_7585);
nand U9198 (N_9198,N_8531,N_8632);
and U9199 (N_9199,N_7698,N_7709);
and U9200 (N_9200,N_8566,N_8612);
nand U9201 (N_9201,N_8474,N_8179);
or U9202 (N_9202,N_8467,N_8050);
nor U9203 (N_9203,N_8296,N_7790);
or U9204 (N_9204,N_8236,N_8252);
or U9205 (N_9205,N_7897,N_7663);
and U9206 (N_9206,N_8482,N_7563);
xnor U9207 (N_9207,N_8375,N_7726);
xnor U9208 (N_9208,N_8126,N_8344);
or U9209 (N_9209,N_8315,N_7764);
xnor U9210 (N_9210,N_7871,N_7721);
nand U9211 (N_9211,N_7766,N_8636);
and U9212 (N_9212,N_8390,N_8167);
xor U9213 (N_9213,N_8198,N_8707);
xnor U9214 (N_9214,N_8009,N_7615);
nor U9215 (N_9215,N_7516,N_8430);
or U9216 (N_9216,N_8307,N_7782);
nor U9217 (N_9217,N_8498,N_7527);
and U9218 (N_9218,N_7690,N_8505);
or U9219 (N_9219,N_7760,N_7641);
nor U9220 (N_9220,N_7920,N_8139);
nor U9221 (N_9221,N_7600,N_7591);
and U9222 (N_9222,N_8335,N_8173);
and U9223 (N_9223,N_7761,N_7511);
or U9224 (N_9224,N_8322,N_8436);
nor U9225 (N_9225,N_8309,N_7767);
or U9226 (N_9226,N_8635,N_8654);
nor U9227 (N_9227,N_7970,N_8349);
xnor U9228 (N_9228,N_7915,N_8734);
nor U9229 (N_9229,N_8327,N_8018);
and U9230 (N_9230,N_8431,N_7826);
nand U9231 (N_9231,N_8096,N_8067);
xnor U9232 (N_9232,N_8539,N_8520);
xnor U9233 (N_9233,N_8159,N_7543);
nor U9234 (N_9234,N_8424,N_8206);
or U9235 (N_9235,N_8556,N_8697);
nand U9236 (N_9236,N_8092,N_7679);
and U9237 (N_9237,N_7696,N_8262);
or U9238 (N_9238,N_7627,N_8260);
nand U9239 (N_9239,N_8112,N_7594);
and U9240 (N_9240,N_8288,N_7842);
nor U9241 (N_9241,N_8731,N_8213);
nand U9242 (N_9242,N_8712,N_7708);
or U9243 (N_9243,N_7938,N_8207);
and U9244 (N_9244,N_8579,N_7553);
and U9245 (N_9245,N_8034,N_7937);
nor U9246 (N_9246,N_7751,N_7648);
and U9247 (N_9247,N_8733,N_8263);
nor U9248 (N_9248,N_7644,N_7844);
xnor U9249 (N_9249,N_8245,N_7911);
nor U9250 (N_9250,N_8152,N_7544);
and U9251 (N_9251,N_7656,N_8692);
and U9252 (N_9252,N_7670,N_8038);
or U9253 (N_9253,N_8178,N_7745);
or U9254 (N_9254,N_8507,N_8747);
or U9255 (N_9255,N_8101,N_7507);
and U9256 (N_9256,N_8610,N_8129);
nor U9257 (N_9257,N_8070,N_7942);
nor U9258 (N_9258,N_8736,N_7845);
nor U9259 (N_9259,N_8404,N_8035);
nor U9260 (N_9260,N_7734,N_8128);
or U9261 (N_9261,N_7593,N_8210);
xor U9262 (N_9262,N_8682,N_7858);
nand U9263 (N_9263,N_8417,N_8725);
nor U9264 (N_9264,N_7634,N_8085);
and U9265 (N_9265,N_7753,N_7697);
xor U9266 (N_9266,N_8224,N_8042);
or U9267 (N_9267,N_8283,N_7671);
or U9268 (N_9268,N_7939,N_8247);
nand U9269 (N_9269,N_7900,N_7554);
xnor U9270 (N_9270,N_8361,N_8110);
xnor U9271 (N_9271,N_8219,N_8538);
xor U9272 (N_9272,N_8205,N_7780);
xnor U9273 (N_9273,N_8631,N_8448);
nor U9274 (N_9274,N_8383,N_7597);
nor U9275 (N_9275,N_8121,N_7678);
nor U9276 (N_9276,N_8363,N_7778);
nand U9277 (N_9277,N_8462,N_8540);
or U9278 (N_9278,N_7587,N_7756);
nand U9279 (N_9279,N_8530,N_8720);
nand U9280 (N_9280,N_8702,N_8748);
nand U9281 (N_9281,N_8413,N_8594);
nor U9282 (N_9282,N_8416,N_8453);
nor U9283 (N_9283,N_8517,N_8581);
nand U9284 (N_9284,N_7573,N_7712);
nor U9285 (N_9285,N_8410,N_7818);
or U9286 (N_9286,N_8045,N_8740);
nor U9287 (N_9287,N_7624,N_8033);
xor U9288 (N_9288,N_8468,N_8603);
or U9289 (N_9289,N_8320,N_7737);
or U9290 (N_9290,N_8191,N_8055);
and U9291 (N_9291,N_7707,N_7672);
nor U9292 (N_9292,N_8019,N_8384);
or U9293 (N_9293,N_8393,N_8155);
nand U9294 (N_9294,N_7877,N_8730);
xnor U9295 (N_9295,N_7520,N_8586);
and U9296 (N_9296,N_8493,N_8589);
or U9297 (N_9297,N_8130,N_8728);
nor U9298 (N_9298,N_7640,N_8216);
nand U9299 (N_9299,N_8710,N_8484);
or U9300 (N_9300,N_8215,N_8137);
xnor U9301 (N_9301,N_8182,N_8640);
and U9302 (N_9302,N_7898,N_7792);
xor U9303 (N_9303,N_8522,N_8732);
nor U9304 (N_9304,N_8371,N_8749);
nor U9305 (N_9305,N_7872,N_7539);
nand U9306 (N_9306,N_7769,N_8177);
nor U9307 (N_9307,N_8325,N_7951);
nand U9308 (N_9308,N_8300,N_8667);
or U9309 (N_9309,N_8002,N_8012);
nand U9310 (N_9310,N_7986,N_8657);
or U9311 (N_9311,N_7924,N_8669);
and U9312 (N_9312,N_8265,N_7598);
xor U9313 (N_9313,N_7856,N_7739);
nand U9314 (N_9314,N_7570,N_7925);
xnor U9315 (N_9315,N_7918,N_8290);
and U9316 (N_9316,N_7980,N_8703);
xnor U9317 (N_9317,N_8571,N_7979);
and U9318 (N_9318,N_8049,N_8211);
nor U9319 (N_9319,N_7559,N_7676);
nor U9320 (N_9320,N_7601,N_8438);
or U9321 (N_9321,N_8475,N_8082);
or U9322 (N_9322,N_7504,N_7605);
nand U9323 (N_9323,N_7993,N_7796);
nor U9324 (N_9324,N_7795,N_8481);
or U9325 (N_9325,N_8369,N_8407);
nand U9326 (N_9326,N_8629,N_8423);
or U9327 (N_9327,N_7706,N_7680);
xnor U9328 (N_9328,N_7659,N_8257);
nor U9329 (N_9329,N_8270,N_7643);
nor U9330 (N_9330,N_8681,N_8432);
and U9331 (N_9331,N_7713,N_7694);
nor U9332 (N_9332,N_8442,N_7629);
or U9333 (N_9333,N_8403,N_8716);
or U9334 (N_9334,N_7619,N_8062);
or U9335 (N_9335,N_8136,N_7762);
xnor U9336 (N_9336,N_8025,N_8648);
nor U9337 (N_9337,N_8281,N_7635);
and U9338 (N_9338,N_7693,N_7579);
and U9339 (N_9339,N_8084,N_8613);
and U9340 (N_9340,N_7879,N_8574);
xnor U9341 (N_9341,N_8560,N_7828);
and U9342 (N_9342,N_8745,N_8547);
and U9343 (N_9343,N_8318,N_7815);
nor U9344 (N_9344,N_7785,N_8313);
nor U9345 (N_9345,N_8373,N_8243);
or U9346 (N_9346,N_8515,N_8638);
nand U9347 (N_9347,N_8563,N_7908);
nor U9348 (N_9348,N_8158,N_7996);
and U9349 (N_9349,N_8143,N_8040);
xor U9350 (N_9350,N_7870,N_7502);
xor U9351 (N_9351,N_8497,N_7989);
xor U9352 (N_9352,N_8041,N_7534);
nand U9353 (N_9353,N_7662,N_7592);
nor U9354 (N_9354,N_8108,N_8275);
or U9355 (N_9355,N_7750,N_8492);
xnor U9356 (N_9356,N_7997,N_8616);
nand U9357 (N_9357,N_8065,N_7804);
nand U9358 (N_9358,N_8599,N_8420);
xor U9359 (N_9359,N_8674,N_7808);
or U9360 (N_9360,N_8721,N_8006);
or U9361 (N_9361,N_7728,N_7555);
nand U9362 (N_9362,N_8195,N_8046);
nand U9363 (N_9363,N_7704,N_8119);
or U9364 (N_9364,N_7675,N_7528);
and U9365 (N_9365,N_8218,N_8214);
nand U9366 (N_9366,N_8276,N_7701);
or U9367 (N_9367,N_8429,N_7859);
nor U9368 (N_9368,N_7880,N_7522);
xor U9369 (N_9369,N_7800,N_8392);
or U9370 (N_9370,N_7580,N_8066);
nand U9371 (N_9371,N_8271,N_8201);
nor U9372 (N_9372,N_8735,N_7525);
nor U9373 (N_9373,N_8743,N_7617);
and U9374 (N_9374,N_8705,N_7954);
nor U9375 (N_9375,N_8363,N_8625);
nor U9376 (N_9376,N_8240,N_8096);
nand U9377 (N_9377,N_8642,N_7500);
xor U9378 (N_9378,N_8446,N_8314);
nand U9379 (N_9379,N_8339,N_7699);
xnor U9380 (N_9380,N_7929,N_8543);
nor U9381 (N_9381,N_7523,N_8400);
xnor U9382 (N_9382,N_8166,N_7712);
nor U9383 (N_9383,N_7922,N_7926);
and U9384 (N_9384,N_8515,N_8710);
xnor U9385 (N_9385,N_8672,N_8617);
nand U9386 (N_9386,N_7707,N_7788);
and U9387 (N_9387,N_8505,N_7683);
nand U9388 (N_9388,N_8012,N_7586);
and U9389 (N_9389,N_7598,N_8043);
and U9390 (N_9390,N_7734,N_7587);
nand U9391 (N_9391,N_8614,N_7624);
nand U9392 (N_9392,N_8634,N_8590);
xnor U9393 (N_9393,N_8332,N_8268);
and U9394 (N_9394,N_8519,N_8218);
or U9395 (N_9395,N_8322,N_8026);
xnor U9396 (N_9396,N_7821,N_7916);
nor U9397 (N_9397,N_7893,N_8624);
nand U9398 (N_9398,N_7566,N_7766);
nor U9399 (N_9399,N_8208,N_7954);
and U9400 (N_9400,N_7935,N_8545);
and U9401 (N_9401,N_7568,N_8306);
or U9402 (N_9402,N_7688,N_7946);
and U9403 (N_9403,N_8281,N_7760);
or U9404 (N_9404,N_8396,N_7570);
or U9405 (N_9405,N_8208,N_8311);
nor U9406 (N_9406,N_8205,N_8398);
xnor U9407 (N_9407,N_7706,N_7625);
nor U9408 (N_9408,N_7740,N_8553);
or U9409 (N_9409,N_7918,N_8062);
nor U9410 (N_9410,N_7666,N_7849);
or U9411 (N_9411,N_8729,N_8645);
nand U9412 (N_9412,N_7760,N_8263);
xor U9413 (N_9413,N_8384,N_8294);
and U9414 (N_9414,N_8211,N_7624);
and U9415 (N_9415,N_8745,N_8156);
nand U9416 (N_9416,N_7625,N_7927);
nor U9417 (N_9417,N_7757,N_8557);
nor U9418 (N_9418,N_8341,N_7784);
nor U9419 (N_9419,N_8250,N_7819);
nand U9420 (N_9420,N_8436,N_7900);
and U9421 (N_9421,N_7909,N_7962);
xor U9422 (N_9422,N_8291,N_8627);
and U9423 (N_9423,N_8023,N_8346);
and U9424 (N_9424,N_8701,N_8548);
or U9425 (N_9425,N_8666,N_7819);
and U9426 (N_9426,N_8040,N_7699);
xnor U9427 (N_9427,N_8552,N_8331);
nor U9428 (N_9428,N_7878,N_8336);
or U9429 (N_9429,N_8400,N_7803);
or U9430 (N_9430,N_7534,N_8669);
xor U9431 (N_9431,N_7774,N_7927);
nor U9432 (N_9432,N_8303,N_8301);
nand U9433 (N_9433,N_8404,N_7529);
and U9434 (N_9434,N_7782,N_8006);
nand U9435 (N_9435,N_8314,N_8321);
xnor U9436 (N_9436,N_7605,N_8551);
nor U9437 (N_9437,N_8005,N_7676);
xor U9438 (N_9438,N_8693,N_8179);
xor U9439 (N_9439,N_8624,N_7926);
nand U9440 (N_9440,N_8024,N_7643);
nand U9441 (N_9441,N_7929,N_8190);
nor U9442 (N_9442,N_7755,N_7510);
nor U9443 (N_9443,N_8670,N_8109);
nand U9444 (N_9444,N_8314,N_7993);
xor U9445 (N_9445,N_7609,N_8634);
nor U9446 (N_9446,N_7679,N_8309);
or U9447 (N_9447,N_8662,N_8052);
nor U9448 (N_9448,N_7883,N_7668);
nand U9449 (N_9449,N_7712,N_7637);
or U9450 (N_9450,N_7732,N_8140);
and U9451 (N_9451,N_8714,N_8698);
nand U9452 (N_9452,N_7768,N_7585);
nand U9453 (N_9453,N_7865,N_8439);
nor U9454 (N_9454,N_8736,N_7906);
nand U9455 (N_9455,N_8657,N_7525);
xnor U9456 (N_9456,N_7821,N_7972);
and U9457 (N_9457,N_7996,N_8708);
or U9458 (N_9458,N_7854,N_7739);
nand U9459 (N_9459,N_8598,N_7610);
nor U9460 (N_9460,N_8182,N_7550);
nand U9461 (N_9461,N_8695,N_8423);
nor U9462 (N_9462,N_8174,N_7946);
nor U9463 (N_9463,N_8616,N_7805);
xor U9464 (N_9464,N_8668,N_8316);
and U9465 (N_9465,N_8266,N_8564);
nand U9466 (N_9466,N_7741,N_8062);
nor U9467 (N_9467,N_8396,N_7516);
and U9468 (N_9468,N_8370,N_8155);
nand U9469 (N_9469,N_8365,N_8290);
and U9470 (N_9470,N_8730,N_8269);
xnor U9471 (N_9471,N_8550,N_7527);
or U9472 (N_9472,N_8035,N_8175);
and U9473 (N_9473,N_8516,N_8001);
or U9474 (N_9474,N_8058,N_7936);
xor U9475 (N_9475,N_7943,N_8684);
and U9476 (N_9476,N_8242,N_8582);
nor U9477 (N_9477,N_7816,N_7935);
nor U9478 (N_9478,N_8585,N_7611);
nand U9479 (N_9479,N_8277,N_8235);
and U9480 (N_9480,N_8359,N_7741);
and U9481 (N_9481,N_8686,N_8184);
nor U9482 (N_9482,N_7937,N_8640);
nor U9483 (N_9483,N_7623,N_7598);
nor U9484 (N_9484,N_7792,N_8111);
xor U9485 (N_9485,N_7830,N_7643);
xnor U9486 (N_9486,N_7741,N_8378);
and U9487 (N_9487,N_8045,N_8181);
nand U9488 (N_9488,N_7749,N_8035);
or U9489 (N_9489,N_8056,N_8568);
nor U9490 (N_9490,N_7501,N_8683);
nor U9491 (N_9491,N_7991,N_7768);
or U9492 (N_9492,N_7734,N_7506);
nor U9493 (N_9493,N_8633,N_7959);
nor U9494 (N_9494,N_8357,N_7805);
xor U9495 (N_9495,N_8119,N_7791);
xnor U9496 (N_9496,N_8165,N_7791);
and U9497 (N_9497,N_8653,N_8449);
nand U9498 (N_9498,N_7799,N_7694);
and U9499 (N_9499,N_7561,N_7731);
or U9500 (N_9500,N_7753,N_7651);
and U9501 (N_9501,N_8389,N_8493);
xnor U9502 (N_9502,N_7505,N_8005);
or U9503 (N_9503,N_8480,N_8578);
xnor U9504 (N_9504,N_8618,N_7505);
nor U9505 (N_9505,N_7898,N_8265);
xor U9506 (N_9506,N_7983,N_8101);
xnor U9507 (N_9507,N_8416,N_8665);
or U9508 (N_9508,N_8591,N_8125);
nand U9509 (N_9509,N_7681,N_7936);
xnor U9510 (N_9510,N_7550,N_8509);
nor U9511 (N_9511,N_8601,N_7789);
nor U9512 (N_9512,N_7775,N_7550);
or U9513 (N_9513,N_8352,N_8386);
or U9514 (N_9514,N_8027,N_8336);
or U9515 (N_9515,N_8420,N_7795);
xor U9516 (N_9516,N_7580,N_7837);
or U9517 (N_9517,N_7888,N_7999);
and U9518 (N_9518,N_8204,N_8358);
or U9519 (N_9519,N_8602,N_8347);
xor U9520 (N_9520,N_8003,N_8546);
or U9521 (N_9521,N_7990,N_8376);
nor U9522 (N_9522,N_8736,N_7582);
or U9523 (N_9523,N_8183,N_8525);
or U9524 (N_9524,N_8163,N_8062);
and U9525 (N_9525,N_7649,N_7676);
nor U9526 (N_9526,N_8518,N_7982);
xor U9527 (N_9527,N_8110,N_7669);
nand U9528 (N_9528,N_7658,N_8146);
or U9529 (N_9529,N_7864,N_8541);
nand U9530 (N_9530,N_8587,N_8135);
nand U9531 (N_9531,N_7780,N_8409);
nor U9532 (N_9532,N_7959,N_8205);
and U9533 (N_9533,N_7580,N_8437);
and U9534 (N_9534,N_8098,N_8470);
or U9535 (N_9535,N_7655,N_7625);
nor U9536 (N_9536,N_7704,N_7772);
and U9537 (N_9537,N_8604,N_8406);
nor U9538 (N_9538,N_8220,N_7805);
and U9539 (N_9539,N_7821,N_8399);
nor U9540 (N_9540,N_8163,N_8126);
nand U9541 (N_9541,N_7627,N_8484);
xnor U9542 (N_9542,N_8038,N_7509);
xnor U9543 (N_9543,N_8567,N_8036);
xor U9544 (N_9544,N_7729,N_7816);
and U9545 (N_9545,N_8718,N_8228);
nand U9546 (N_9546,N_8114,N_8492);
xor U9547 (N_9547,N_8204,N_8539);
nor U9548 (N_9548,N_8295,N_8475);
nand U9549 (N_9549,N_7756,N_7878);
nand U9550 (N_9550,N_8381,N_8622);
nor U9551 (N_9551,N_7548,N_7506);
and U9552 (N_9552,N_8589,N_8041);
and U9553 (N_9553,N_7922,N_7818);
xor U9554 (N_9554,N_8575,N_8325);
and U9555 (N_9555,N_7866,N_7597);
nand U9556 (N_9556,N_7754,N_8516);
nand U9557 (N_9557,N_7571,N_8447);
and U9558 (N_9558,N_7817,N_7847);
xnor U9559 (N_9559,N_8402,N_8534);
or U9560 (N_9560,N_8003,N_8271);
and U9561 (N_9561,N_8572,N_8208);
nor U9562 (N_9562,N_8648,N_8571);
or U9563 (N_9563,N_7668,N_8181);
or U9564 (N_9564,N_8605,N_8499);
and U9565 (N_9565,N_7977,N_7790);
nor U9566 (N_9566,N_8133,N_8743);
xor U9567 (N_9567,N_7663,N_8175);
nand U9568 (N_9568,N_8049,N_8637);
nand U9569 (N_9569,N_8376,N_8316);
xnor U9570 (N_9570,N_8023,N_8030);
or U9571 (N_9571,N_7995,N_7678);
and U9572 (N_9572,N_8539,N_7577);
or U9573 (N_9573,N_8404,N_8004);
xnor U9574 (N_9574,N_8405,N_7887);
nor U9575 (N_9575,N_8588,N_7615);
and U9576 (N_9576,N_7512,N_8193);
and U9577 (N_9577,N_7609,N_7822);
and U9578 (N_9578,N_7857,N_7819);
or U9579 (N_9579,N_7603,N_7878);
or U9580 (N_9580,N_7897,N_7990);
xor U9581 (N_9581,N_7746,N_8252);
nand U9582 (N_9582,N_7922,N_8380);
xnor U9583 (N_9583,N_8072,N_8211);
nor U9584 (N_9584,N_8736,N_7782);
nor U9585 (N_9585,N_8034,N_7824);
and U9586 (N_9586,N_7935,N_8401);
or U9587 (N_9587,N_7949,N_7918);
nor U9588 (N_9588,N_7761,N_7650);
nor U9589 (N_9589,N_8509,N_7753);
or U9590 (N_9590,N_7984,N_8288);
or U9591 (N_9591,N_8096,N_7643);
nand U9592 (N_9592,N_7753,N_8259);
and U9593 (N_9593,N_8740,N_8712);
nand U9594 (N_9594,N_8160,N_7821);
xnor U9595 (N_9595,N_7971,N_7730);
and U9596 (N_9596,N_7967,N_8027);
xnor U9597 (N_9597,N_8093,N_8099);
nand U9598 (N_9598,N_7813,N_7527);
or U9599 (N_9599,N_8605,N_8510);
and U9600 (N_9600,N_8439,N_8626);
xnor U9601 (N_9601,N_8626,N_8504);
and U9602 (N_9602,N_8203,N_8223);
and U9603 (N_9603,N_8560,N_7922);
xor U9604 (N_9604,N_8304,N_7906);
xnor U9605 (N_9605,N_8426,N_7833);
and U9606 (N_9606,N_8143,N_8620);
nand U9607 (N_9607,N_8666,N_8515);
and U9608 (N_9608,N_7916,N_8521);
nor U9609 (N_9609,N_8737,N_8161);
xor U9610 (N_9610,N_7717,N_8730);
or U9611 (N_9611,N_8178,N_7979);
xnor U9612 (N_9612,N_8429,N_8218);
and U9613 (N_9613,N_8692,N_8195);
nand U9614 (N_9614,N_8641,N_7954);
and U9615 (N_9615,N_8150,N_7507);
nand U9616 (N_9616,N_7958,N_8030);
and U9617 (N_9617,N_8399,N_7953);
nand U9618 (N_9618,N_7964,N_8282);
or U9619 (N_9619,N_8544,N_8474);
nand U9620 (N_9620,N_7910,N_7648);
and U9621 (N_9621,N_7674,N_8136);
and U9622 (N_9622,N_7613,N_7930);
nor U9623 (N_9623,N_8172,N_7980);
nand U9624 (N_9624,N_8077,N_8237);
nand U9625 (N_9625,N_7677,N_7665);
xnor U9626 (N_9626,N_8594,N_7725);
xor U9627 (N_9627,N_8644,N_7701);
or U9628 (N_9628,N_8435,N_8726);
nand U9629 (N_9629,N_7680,N_8409);
or U9630 (N_9630,N_8124,N_8746);
nand U9631 (N_9631,N_8654,N_7906);
nor U9632 (N_9632,N_8618,N_7664);
and U9633 (N_9633,N_8478,N_7671);
xnor U9634 (N_9634,N_8269,N_8040);
xor U9635 (N_9635,N_8161,N_8079);
nor U9636 (N_9636,N_8501,N_7805);
or U9637 (N_9637,N_8732,N_8279);
nor U9638 (N_9638,N_8159,N_8428);
and U9639 (N_9639,N_8609,N_7962);
or U9640 (N_9640,N_8657,N_7674);
xor U9641 (N_9641,N_8226,N_8289);
xor U9642 (N_9642,N_7629,N_7858);
xor U9643 (N_9643,N_8518,N_7702);
and U9644 (N_9644,N_7735,N_8724);
xor U9645 (N_9645,N_8612,N_7609);
nor U9646 (N_9646,N_8240,N_7741);
and U9647 (N_9647,N_8638,N_8358);
xor U9648 (N_9648,N_8112,N_8576);
or U9649 (N_9649,N_8005,N_8374);
nand U9650 (N_9650,N_8449,N_8576);
nand U9651 (N_9651,N_8464,N_8579);
and U9652 (N_9652,N_7527,N_8344);
nand U9653 (N_9653,N_8516,N_7501);
and U9654 (N_9654,N_7658,N_8445);
and U9655 (N_9655,N_8128,N_8710);
and U9656 (N_9656,N_7544,N_8688);
xor U9657 (N_9657,N_8407,N_7609);
and U9658 (N_9658,N_8354,N_8062);
and U9659 (N_9659,N_7703,N_8492);
nor U9660 (N_9660,N_7985,N_8034);
xor U9661 (N_9661,N_7971,N_7988);
nand U9662 (N_9662,N_7616,N_7672);
xor U9663 (N_9663,N_7529,N_7909);
xnor U9664 (N_9664,N_8380,N_8069);
and U9665 (N_9665,N_8059,N_8217);
or U9666 (N_9666,N_7565,N_8413);
or U9667 (N_9667,N_7737,N_8284);
nand U9668 (N_9668,N_7818,N_8319);
or U9669 (N_9669,N_8541,N_7999);
xor U9670 (N_9670,N_7978,N_7975);
nor U9671 (N_9671,N_7618,N_8591);
and U9672 (N_9672,N_8562,N_8210);
nor U9673 (N_9673,N_7519,N_8209);
nand U9674 (N_9674,N_7977,N_8133);
or U9675 (N_9675,N_8064,N_7809);
xnor U9676 (N_9676,N_7548,N_8183);
nor U9677 (N_9677,N_8675,N_8579);
xnor U9678 (N_9678,N_7808,N_7870);
xor U9679 (N_9679,N_8271,N_8086);
nor U9680 (N_9680,N_7949,N_7786);
xor U9681 (N_9681,N_8120,N_8413);
xnor U9682 (N_9682,N_7919,N_8478);
or U9683 (N_9683,N_8497,N_8369);
nand U9684 (N_9684,N_8056,N_7863);
xnor U9685 (N_9685,N_8355,N_7681);
xnor U9686 (N_9686,N_8574,N_7900);
and U9687 (N_9687,N_8204,N_7696);
nand U9688 (N_9688,N_8531,N_8623);
nand U9689 (N_9689,N_7625,N_8448);
and U9690 (N_9690,N_8609,N_8240);
nand U9691 (N_9691,N_8530,N_8039);
nor U9692 (N_9692,N_7994,N_7526);
and U9693 (N_9693,N_8401,N_7601);
xnor U9694 (N_9694,N_8149,N_8250);
nor U9695 (N_9695,N_8639,N_7810);
nor U9696 (N_9696,N_7928,N_8265);
or U9697 (N_9697,N_7670,N_7651);
nor U9698 (N_9698,N_7924,N_8389);
xor U9699 (N_9699,N_8357,N_8460);
nand U9700 (N_9700,N_8370,N_8683);
nor U9701 (N_9701,N_8138,N_7891);
nand U9702 (N_9702,N_8501,N_8168);
xor U9703 (N_9703,N_7908,N_7735);
xor U9704 (N_9704,N_8313,N_7875);
nand U9705 (N_9705,N_8450,N_8219);
and U9706 (N_9706,N_8383,N_8643);
nand U9707 (N_9707,N_8508,N_7646);
nor U9708 (N_9708,N_7897,N_8387);
nand U9709 (N_9709,N_8364,N_8323);
or U9710 (N_9710,N_8744,N_8112);
nand U9711 (N_9711,N_8351,N_7595);
and U9712 (N_9712,N_8499,N_8410);
and U9713 (N_9713,N_8727,N_7506);
xor U9714 (N_9714,N_8599,N_7816);
nor U9715 (N_9715,N_7520,N_7919);
nand U9716 (N_9716,N_8383,N_7742);
nand U9717 (N_9717,N_7931,N_8150);
and U9718 (N_9718,N_8415,N_7952);
or U9719 (N_9719,N_7803,N_7559);
xnor U9720 (N_9720,N_8238,N_8383);
nor U9721 (N_9721,N_7689,N_8632);
xnor U9722 (N_9722,N_7657,N_7845);
or U9723 (N_9723,N_7541,N_8445);
nor U9724 (N_9724,N_8389,N_7758);
nand U9725 (N_9725,N_7712,N_8263);
or U9726 (N_9726,N_8357,N_8625);
or U9727 (N_9727,N_7595,N_7740);
and U9728 (N_9728,N_7985,N_8260);
and U9729 (N_9729,N_7954,N_7792);
and U9730 (N_9730,N_7716,N_7511);
xnor U9731 (N_9731,N_8726,N_7935);
and U9732 (N_9732,N_7537,N_7733);
xor U9733 (N_9733,N_7947,N_8671);
nand U9734 (N_9734,N_8610,N_8533);
xor U9735 (N_9735,N_8447,N_8650);
xnor U9736 (N_9736,N_8325,N_7770);
nor U9737 (N_9737,N_8483,N_8724);
or U9738 (N_9738,N_7574,N_8136);
and U9739 (N_9739,N_8016,N_7633);
nand U9740 (N_9740,N_8377,N_8356);
nor U9741 (N_9741,N_8523,N_7591);
nand U9742 (N_9742,N_7945,N_8175);
nor U9743 (N_9743,N_8124,N_8333);
and U9744 (N_9744,N_7575,N_8179);
and U9745 (N_9745,N_7807,N_7821);
nand U9746 (N_9746,N_8643,N_8335);
and U9747 (N_9747,N_8733,N_8381);
nand U9748 (N_9748,N_8699,N_7703);
xnor U9749 (N_9749,N_8409,N_8226);
nor U9750 (N_9750,N_7526,N_8186);
and U9751 (N_9751,N_8215,N_8021);
and U9752 (N_9752,N_7691,N_8584);
or U9753 (N_9753,N_7713,N_7522);
xnor U9754 (N_9754,N_8735,N_7940);
and U9755 (N_9755,N_8307,N_8517);
nand U9756 (N_9756,N_7676,N_7547);
or U9757 (N_9757,N_8472,N_7772);
or U9758 (N_9758,N_8618,N_7662);
and U9759 (N_9759,N_8335,N_8239);
xor U9760 (N_9760,N_7883,N_8096);
xor U9761 (N_9761,N_8177,N_8059);
xor U9762 (N_9762,N_7610,N_7852);
or U9763 (N_9763,N_8303,N_8003);
and U9764 (N_9764,N_8678,N_7760);
nand U9765 (N_9765,N_7846,N_8592);
nor U9766 (N_9766,N_8096,N_8051);
and U9767 (N_9767,N_7847,N_8205);
or U9768 (N_9768,N_8724,N_8540);
or U9769 (N_9769,N_7929,N_7746);
or U9770 (N_9770,N_8620,N_7959);
xnor U9771 (N_9771,N_8276,N_8740);
nor U9772 (N_9772,N_8695,N_8224);
nand U9773 (N_9773,N_8432,N_8151);
and U9774 (N_9774,N_8607,N_8095);
or U9775 (N_9775,N_8107,N_7856);
or U9776 (N_9776,N_8608,N_8104);
xor U9777 (N_9777,N_8058,N_8365);
and U9778 (N_9778,N_8357,N_7872);
nand U9779 (N_9779,N_8609,N_8061);
xor U9780 (N_9780,N_8444,N_7835);
or U9781 (N_9781,N_8587,N_8170);
and U9782 (N_9782,N_8354,N_8497);
nor U9783 (N_9783,N_8023,N_8063);
nand U9784 (N_9784,N_7825,N_8355);
nand U9785 (N_9785,N_8452,N_8426);
nor U9786 (N_9786,N_8437,N_8258);
and U9787 (N_9787,N_8551,N_7694);
xnor U9788 (N_9788,N_8688,N_7857);
and U9789 (N_9789,N_7804,N_7807);
xnor U9790 (N_9790,N_8358,N_8608);
and U9791 (N_9791,N_7987,N_8350);
nand U9792 (N_9792,N_8419,N_8277);
nor U9793 (N_9793,N_8242,N_7537);
nor U9794 (N_9794,N_8023,N_8581);
and U9795 (N_9795,N_7736,N_7615);
or U9796 (N_9796,N_7542,N_8012);
or U9797 (N_9797,N_8114,N_8363);
and U9798 (N_9798,N_8223,N_7929);
nor U9799 (N_9799,N_7998,N_8671);
nand U9800 (N_9800,N_7993,N_7655);
nand U9801 (N_9801,N_8343,N_8064);
and U9802 (N_9802,N_7882,N_8318);
xnor U9803 (N_9803,N_8422,N_7980);
nand U9804 (N_9804,N_7996,N_8299);
and U9805 (N_9805,N_7598,N_8167);
nand U9806 (N_9806,N_8100,N_8169);
nand U9807 (N_9807,N_8134,N_8537);
xor U9808 (N_9808,N_8356,N_8126);
xor U9809 (N_9809,N_7708,N_8272);
or U9810 (N_9810,N_8336,N_7742);
or U9811 (N_9811,N_8594,N_7676);
nand U9812 (N_9812,N_8673,N_8506);
nor U9813 (N_9813,N_7614,N_8200);
nand U9814 (N_9814,N_8255,N_8632);
nor U9815 (N_9815,N_8497,N_8344);
xnor U9816 (N_9816,N_7901,N_8510);
and U9817 (N_9817,N_7654,N_7532);
and U9818 (N_9818,N_8402,N_8114);
nor U9819 (N_9819,N_8610,N_8586);
or U9820 (N_9820,N_8630,N_8129);
nor U9821 (N_9821,N_7654,N_8215);
nor U9822 (N_9822,N_8191,N_7657);
xor U9823 (N_9823,N_7982,N_7984);
nand U9824 (N_9824,N_7547,N_7659);
nand U9825 (N_9825,N_8662,N_8350);
xor U9826 (N_9826,N_8294,N_8195);
nand U9827 (N_9827,N_7745,N_8136);
or U9828 (N_9828,N_8716,N_8621);
or U9829 (N_9829,N_8706,N_8549);
nor U9830 (N_9830,N_8051,N_8622);
nor U9831 (N_9831,N_7825,N_8655);
nand U9832 (N_9832,N_8496,N_8096);
and U9833 (N_9833,N_8099,N_8186);
or U9834 (N_9834,N_7793,N_7781);
and U9835 (N_9835,N_7852,N_8153);
xor U9836 (N_9836,N_8465,N_7670);
nand U9837 (N_9837,N_8642,N_8109);
nor U9838 (N_9838,N_8748,N_7773);
xor U9839 (N_9839,N_8016,N_8724);
nand U9840 (N_9840,N_7597,N_8085);
nor U9841 (N_9841,N_8452,N_8019);
and U9842 (N_9842,N_8136,N_7962);
and U9843 (N_9843,N_8689,N_7710);
and U9844 (N_9844,N_8619,N_8210);
nand U9845 (N_9845,N_7513,N_7725);
or U9846 (N_9846,N_8721,N_8035);
nor U9847 (N_9847,N_8330,N_7536);
nor U9848 (N_9848,N_8625,N_7902);
nand U9849 (N_9849,N_8448,N_8730);
xnor U9850 (N_9850,N_7753,N_8461);
or U9851 (N_9851,N_7706,N_8647);
xor U9852 (N_9852,N_7688,N_8487);
nand U9853 (N_9853,N_8475,N_8568);
or U9854 (N_9854,N_7884,N_7902);
nand U9855 (N_9855,N_8748,N_8604);
xor U9856 (N_9856,N_7842,N_7825);
or U9857 (N_9857,N_8093,N_8615);
and U9858 (N_9858,N_8437,N_7981);
nor U9859 (N_9859,N_8733,N_7583);
nor U9860 (N_9860,N_7845,N_8009);
nor U9861 (N_9861,N_8408,N_8232);
xor U9862 (N_9862,N_7612,N_8440);
and U9863 (N_9863,N_7894,N_8365);
nor U9864 (N_9864,N_8614,N_7619);
nand U9865 (N_9865,N_8567,N_8692);
or U9866 (N_9866,N_8555,N_8472);
nand U9867 (N_9867,N_8189,N_8052);
nor U9868 (N_9868,N_8656,N_7746);
or U9869 (N_9869,N_8397,N_8003);
and U9870 (N_9870,N_7912,N_8174);
xor U9871 (N_9871,N_8633,N_8659);
xor U9872 (N_9872,N_8358,N_8216);
or U9873 (N_9873,N_7882,N_8571);
or U9874 (N_9874,N_7951,N_8317);
or U9875 (N_9875,N_8011,N_8739);
xnor U9876 (N_9876,N_7563,N_8737);
nand U9877 (N_9877,N_8721,N_7668);
and U9878 (N_9878,N_8506,N_8344);
nand U9879 (N_9879,N_7966,N_8624);
xor U9880 (N_9880,N_8054,N_7725);
nand U9881 (N_9881,N_8483,N_8603);
or U9882 (N_9882,N_8544,N_8397);
nand U9883 (N_9883,N_7989,N_8092);
or U9884 (N_9884,N_8373,N_7836);
and U9885 (N_9885,N_8674,N_8400);
or U9886 (N_9886,N_8140,N_8647);
or U9887 (N_9887,N_7554,N_7543);
and U9888 (N_9888,N_8694,N_8489);
nand U9889 (N_9889,N_7841,N_8250);
xor U9890 (N_9890,N_7871,N_8508);
or U9891 (N_9891,N_8014,N_8099);
xor U9892 (N_9892,N_8360,N_8322);
nand U9893 (N_9893,N_8120,N_7615);
xnor U9894 (N_9894,N_7721,N_8232);
or U9895 (N_9895,N_8679,N_8516);
xor U9896 (N_9896,N_7512,N_8543);
xnor U9897 (N_9897,N_8044,N_7666);
or U9898 (N_9898,N_7671,N_7850);
and U9899 (N_9899,N_8100,N_8070);
and U9900 (N_9900,N_8583,N_7816);
and U9901 (N_9901,N_7779,N_7920);
or U9902 (N_9902,N_8700,N_8322);
and U9903 (N_9903,N_8266,N_8357);
nor U9904 (N_9904,N_8117,N_7517);
and U9905 (N_9905,N_8535,N_8433);
nand U9906 (N_9906,N_8066,N_8461);
and U9907 (N_9907,N_8468,N_7583);
nor U9908 (N_9908,N_8342,N_8411);
nor U9909 (N_9909,N_7903,N_7969);
nand U9910 (N_9910,N_7865,N_8175);
or U9911 (N_9911,N_7859,N_8423);
and U9912 (N_9912,N_8078,N_8214);
nor U9913 (N_9913,N_7925,N_8451);
nand U9914 (N_9914,N_8721,N_8073);
nor U9915 (N_9915,N_8740,N_8113);
xor U9916 (N_9916,N_8177,N_7597);
nor U9917 (N_9917,N_8153,N_7664);
and U9918 (N_9918,N_8422,N_7644);
and U9919 (N_9919,N_7789,N_7578);
or U9920 (N_9920,N_7812,N_8373);
nor U9921 (N_9921,N_7987,N_8670);
nor U9922 (N_9922,N_8298,N_8213);
and U9923 (N_9923,N_8694,N_8660);
nor U9924 (N_9924,N_7971,N_8376);
and U9925 (N_9925,N_7934,N_8276);
and U9926 (N_9926,N_8228,N_7655);
nand U9927 (N_9927,N_7531,N_7660);
or U9928 (N_9928,N_8037,N_8534);
nand U9929 (N_9929,N_8032,N_8044);
and U9930 (N_9930,N_8091,N_8502);
nor U9931 (N_9931,N_8200,N_8051);
nand U9932 (N_9932,N_7717,N_8058);
xor U9933 (N_9933,N_7699,N_8170);
nand U9934 (N_9934,N_7772,N_7675);
nor U9935 (N_9935,N_8043,N_8559);
nor U9936 (N_9936,N_8305,N_7970);
xor U9937 (N_9937,N_8096,N_7930);
or U9938 (N_9938,N_8173,N_7983);
nand U9939 (N_9939,N_8596,N_7591);
xnor U9940 (N_9940,N_8477,N_8685);
and U9941 (N_9941,N_8581,N_8661);
xor U9942 (N_9942,N_7893,N_8672);
and U9943 (N_9943,N_7833,N_7522);
and U9944 (N_9944,N_7537,N_8532);
or U9945 (N_9945,N_7780,N_8162);
and U9946 (N_9946,N_7603,N_8379);
and U9947 (N_9947,N_7729,N_8623);
nand U9948 (N_9948,N_8125,N_7537);
nand U9949 (N_9949,N_7717,N_8153);
xnor U9950 (N_9950,N_7796,N_8585);
nand U9951 (N_9951,N_8110,N_7831);
and U9952 (N_9952,N_8450,N_7588);
xnor U9953 (N_9953,N_8134,N_8254);
or U9954 (N_9954,N_7963,N_8512);
or U9955 (N_9955,N_8188,N_7886);
and U9956 (N_9956,N_7947,N_7691);
nand U9957 (N_9957,N_8641,N_7655);
xnor U9958 (N_9958,N_8671,N_8499);
or U9959 (N_9959,N_7590,N_7862);
nor U9960 (N_9960,N_8447,N_8500);
and U9961 (N_9961,N_7552,N_7954);
nor U9962 (N_9962,N_8505,N_8305);
and U9963 (N_9963,N_7673,N_7927);
or U9964 (N_9964,N_7832,N_7593);
or U9965 (N_9965,N_8166,N_7737);
xnor U9966 (N_9966,N_7683,N_7995);
nand U9967 (N_9967,N_7689,N_7669);
xor U9968 (N_9968,N_7612,N_8049);
nor U9969 (N_9969,N_8246,N_8341);
nand U9970 (N_9970,N_7966,N_8406);
nor U9971 (N_9971,N_8659,N_8717);
and U9972 (N_9972,N_7742,N_8562);
and U9973 (N_9973,N_8182,N_7615);
nand U9974 (N_9974,N_7651,N_8500);
or U9975 (N_9975,N_8680,N_7908);
and U9976 (N_9976,N_8055,N_7546);
nand U9977 (N_9977,N_7794,N_7521);
or U9978 (N_9978,N_7846,N_7766);
and U9979 (N_9979,N_7512,N_7673);
xor U9980 (N_9980,N_7714,N_7799);
or U9981 (N_9981,N_8552,N_8106);
and U9982 (N_9982,N_7687,N_8327);
nand U9983 (N_9983,N_7841,N_8682);
xor U9984 (N_9984,N_8087,N_7956);
or U9985 (N_9985,N_8606,N_7639);
xor U9986 (N_9986,N_7774,N_8692);
or U9987 (N_9987,N_8177,N_8610);
xor U9988 (N_9988,N_8036,N_7609);
and U9989 (N_9989,N_8497,N_8561);
xor U9990 (N_9990,N_8198,N_7824);
nor U9991 (N_9991,N_7920,N_7765);
nand U9992 (N_9992,N_7980,N_8418);
nand U9993 (N_9993,N_8306,N_8106);
and U9994 (N_9994,N_7975,N_8565);
or U9995 (N_9995,N_7759,N_8014);
or U9996 (N_9996,N_8166,N_8303);
and U9997 (N_9997,N_8277,N_8254);
nand U9998 (N_9998,N_7875,N_7878);
or U9999 (N_9999,N_8591,N_8382);
and U10000 (N_10000,N_9856,N_8946);
and U10001 (N_10001,N_9361,N_9189);
nand U10002 (N_10002,N_9779,N_8943);
and U10003 (N_10003,N_9332,N_9049);
nand U10004 (N_10004,N_9430,N_9754);
nor U10005 (N_10005,N_8923,N_9264);
or U10006 (N_10006,N_9493,N_9663);
and U10007 (N_10007,N_8964,N_9561);
or U10008 (N_10008,N_9733,N_9146);
or U10009 (N_10009,N_8905,N_8882);
nor U10010 (N_10010,N_9028,N_9594);
and U10011 (N_10011,N_8957,N_9042);
nor U10012 (N_10012,N_9622,N_9232);
nand U10013 (N_10013,N_9897,N_9983);
nand U10014 (N_10014,N_9180,N_9112);
xnor U10015 (N_10015,N_9885,N_9477);
or U10016 (N_10016,N_8908,N_9684);
or U10017 (N_10017,N_9910,N_8936);
xor U10018 (N_10018,N_9081,N_9826);
or U10019 (N_10019,N_9389,N_9970);
nor U10020 (N_10020,N_8968,N_9035);
nand U10021 (N_10021,N_9420,N_9019);
nand U10022 (N_10022,N_9410,N_8807);
xor U10023 (N_10023,N_8953,N_8907);
nor U10024 (N_10024,N_9796,N_8871);
nor U10025 (N_10025,N_9501,N_9708);
nor U10026 (N_10026,N_9356,N_8757);
xor U10027 (N_10027,N_9539,N_9080);
xor U10028 (N_10028,N_9169,N_9216);
nand U10029 (N_10029,N_8920,N_9737);
or U10030 (N_10030,N_9235,N_9564);
and U10031 (N_10031,N_9238,N_9914);
xor U10032 (N_10032,N_9443,N_8862);
nand U10033 (N_10033,N_8759,N_9311);
and U10034 (N_10034,N_9157,N_9660);
and U10035 (N_10035,N_9368,N_9106);
nand U10036 (N_10036,N_9740,N_9706);
nor U10037 (N_10037,N_9800,N_9482);
or U10038 (N_10038,N_9436,N_9251);
and U10039 (N_10039,N_9467,N_8947);
and U10040 (N_10040,N_8951,N_9718);
nand U10041 (N_10041,N_9058,N_9476);
and U10042 (N_10042,N_8805,N_8795);
nor U10043 (N_10043,N_9385,N_9269);
or U10044 (N_10044,N_9405,N_9666);
nor U10045 (N_10045,N_9346,N_8984);
or U10046 (N_10046,N_8995,N_8952);
xor U10047 (N_10047,N_9761,N_9426);
and U10048 (N_10048,N_8962,N_9858);
nor U10049 (N_10049,N_8806,N_9782);
or U10050 (N_10050,N_9215,N_9571);
and U10051 (N_10051,N_9535,N_9509);
and U10052 (N_10052,N_9089,N_9766);
nor U10053 (N_10053,N_9808,N_9619);
and U10054 (N_10054,N_9620,N_9004);
nor U10055 (N_10055,N_8988,N_9876);
nor U10056 (N_10056,N_8863,N_9669);
xnor U10057 (N_10057,N_9519,N_9769);
and U10058 (N_10058,N_9022,N_8776);
nand U10059 (N_10059,N_9875,N_9044);
or U10060 (N_10060,N_9202,N_9905);
nand U10061 (N_10061,N_8950,N_8876);
nor U10062 (N_10062,N_9812,N_8883);
or U10063 (N_10063,N_9616,N_9580);
nand U10064 (N_10064,N_9674,N_9111);
nor U10065 (N_10065,N_8755,N_8775);
or U10066 (N_10066,N_9199,N_8915);
nand U10067 (N_10067,N_9387,N_9374);
and U10068 (N_10068,N_9141,N_9802);
nor U10069 (N_10069,N_9661,N_9600);
or U10070 (N_10070,N_9825,N_9234);
and U10071 (N_10071,N_8985,N_9143);
or U10072 (N_10072,N_9518,N_9750);
nand U10073 (N_10073,N_8855,N_9562);
nand U10074 (N_10074,N_9348,N_9790);
and U10075 (N_10075,N_9760,N_9791);
xor U10076 (N_10076,N_9813,N_9176);
and U10077 (N_10077,N_9915,N_9391);
and U10078 (N_10078,N_9676,N_9188);
nand U10079 (N_10079,N_9354,N_8769);
or U10080 (N_10080,N_9423,N_9555);
nand U10081 (N_10081,N_8924,N_9916);
nor U10082 (N_10082,N_9989,N_9634);
or U10083 (N_10083,N_9609,N_9225);
nand U10084 (N_10084,N_9957,N_8999);
nand U10085 (N_10085,N_9558,N_8994);
and U10086 (N_10086,N_9161,N_9831);
or U10087 (N_10087,N_8892,N_9413);
and U10088 (N_10088,N_9147,N_9378);
or U10089 (N_10089,N_8982,N_9290);
or U10090 (N_10090,N_9054,N_9455);
nor U10091 (N_10091,N_9881,N_9966);
nor U10092 (N_10092,N_9972,N_9456);
and U10093 (N_10093,N_9187,N_9593);
nor U10094 (N_10094,N_8828,N_8827);
or U10095 (N_10095,N_9138,N_9412);
nor U10096 (N_10096,N_9742,N_9277);
nor U10097 (N_10097,N_9317,N_9590);
nor U10098 (N_10098,N_9649,N_9442);
and U10099 (N_10099,N_9282,N_9383);
nand U10100 (N_10100,N_9960,N_9931);
or U10101 (N_10101,N_9712,N_9308);
and U10102 (N_10102,N_9369,N_9065);
nand U10103 (N_10103,N_9386,N_9909);
and U10104 (N_10104,N_9472,N_9011);
and U10105 (N_10105,N_9091,N_9878);
nand U10106 (N_10106,N_9118,N_9337);
nor U10107 (N_10107,N_9792,N_9101);
nand U10108 (N_10108,N_9345,N_8959);
xnor U10109 (N_10109,N_8851,N_9009);
nor U10110 (N_10110,N_9324,N_9441);
xnor U10111 (N_10111,N_8991,N_9110);
and U10112 (N_10112,N_9736,N_9124);
nand U10113 (N_10113,N_8928,N_8812);
nor U10114 (N_10114,N_9667,N_9911);
xor U10115 (N_10115,N_9437,N_9727);
and U10116 (N_10116,N_8937,N_9016);
nand U10117 (N_10117,N_9206,N_9228);
or U10118 (N_10118,N_9135,N_9945);
nand U10119 (N_10119,N_9191,N_8902);
or U10120 (N_10120,N_9048,N_9670);
or U10121 (N_10121,N_9172,N_9953);
nor U10122 (N_10122,N_9104,N_9848);
nor U10123 (N_10123,N_9523,N_8773);
nor U10124 (N_10124,N_9056,N_8949);
and U10125 (N_10125,N_8867,N_9505);
and U10126 (N_10126,N_9133,N_8872);
or U10127 (N_10127,N_9087,N_9250);
nand U10128 (N_10128,N_9963,N_9353);
or U10129 (N_10129,N_8890,N_9064);
nor U10130 (N_10130,N_9891,N_9700);
nand U10131 (N_10131,N_9578,N_9732);
or U10132 (N_10132,N_8939,N_8824);
nor U10133 (N_10133,N_9845,N_9409);
and U10134 (N_10134,N_8992,N_9190);
or U10135 (N_10135,N_9956,N_9279);
nor U10136 (N_10136,N_9063,N_9565);
nand U10137 (N_10137,N_8869,N_9928);
nor U10138 (N_10138,N_9842,N_9057);
xor U10139 (N_10139,N_9302,N_9168);
or U10140 (N_10140,N_8954,N_9462);
and U10141 (N_10141,N_9803,N_8986);
or U10142 (N_10142,N_9388,N_9278);
and U10143 (N_10143,N_8932,N_9086);
nand U10144 (N_10144,N_8843,N_9165);
and U10145 (N_10145,N_9984,N_9993);
nand U10146 (N_10146,N_9635,N_9958);
nand U10147 (N_10147,N_9839,N_8958);
or U10148 (N_10148,N_9287,N_9834);
nand U10149 (N_10149,N_9998,N_9285);
nor U10150 (N_10150,N_9399,N_9887);
xnor U10151 (N_10151,N_9488,N_9651);
or U10152 (N_10152,N_9005,N_9039);
or U10153 (N_10153,N_9544,N_8831);
nor U10154 (N_10154,N_8891,N_9673);
xor U10155 (N_10155,N_9381,N_9284);
nand U10156 (N_10156,N_9312,N_8866);
nand U10157 (N_10157,N_9703,N_8990);
nand U10158 (N_10158,N_8938,N_9241);
nand U10159 (N_10159,N_8844,N_8976);
nor U10160 (N_10160,N_9866,N_9077);
or U10161 (N_10161,N_9257,N_9650);
xor U10162 (N_10162,N_8916,N_8931);
nor U10163 (N_10163,N_9880,N_9721);
and U10164 (N_10164,N_9854,N_9390);
or U10165 (N_10165,N_9321,N_9605);
or U10166 (N_10166,N_9171,N_9836);
and U10167 (N_10167,N_9946,N_9526);
xnor U10168 (N_10168,N_8787,N_9102);
nand U10169 (N_10169,N_9444,N_9006);
nor U10170 (N_10170,N_9396,N_9474);
or U10171 (N_10171,N_9731,N_8822);
and U10172 (N_10172,N_8761,N_9184);
nand U10173 (N_10173,N_8980,N_9608);
or U10174 (N_10174,N_9799,N_9490);
xor U10175 (N_10175,N_9314,N_9645);
and U10176 (N_10176,N_9358,N_9429);
or U10177 (N_10177,N_8912,N_9955);
nand U10178 (N_10178,N_9496,N_9258);
nand U10179 (N_10179,N_9768,N_9092);
nand U10180 (N_10180,N_9491,N_9751);
nand U10181 (N_10181,N_8978,N_8893);
and U10182 (N_10182,N_9116,N_8799);
and U10183 (N_10183,N_9355,N_9267);
and U10184 (N_10184,N_9581,N_9136);
or U10185 (N_10185,N_9722,N_9806);
nor U10186 (N_10186,N_9626,N_9394);
nor U10187 (N_10187,N_8821,N_9599);
or U10188 (N_10188,N_9236,N_9170);
or U10189 (N_10189,N_9631,N_9985);
and U10190 (N_10190,N_8911,N_9967);
xor U10191 (N_10191,N_9687,N_9363);
and U10192 (N_10192,N_9705,N_9300);
and U10193 (N_10193,N_9741,N_9400);
nand U10194 (N_10194,N_9192,N_9772);
and U10195 (N_10195,N_9130,N_9018);
and U10196 (N_10196,N_9654,N_9852);
and U10197 (N_10197,N_9720,N_8913);
nand U10198 (N_10198,N_9893,N_9506);
xnor U10199 (N_10199,N_9589,N_9568);
xor U10200 (N_10200,N_9922,N_9725);
or U10201 (N_10201,N_9197,N_9465);
or U10202 (N_10202,N_9884,N_9224);
and U10203 (N_10203,N_9890,N_9752);
and U10204 (N_10204,N_9747,N_9869);
xor U10205 (N_10205,N_9560,N_9194);
nor U10206 (N_10206,N_9757,N_9694);
nor U10207 (N_10207,N_8922,N_9053);
or U10208 (N_10208,N_9440,N_9533);
or U10209 (N_10209,N_9098,N_9809);
and U10210 (N_10210,N_9129,N_8861);
and U10211 (N_10211,N_8974,N_9811);
xor U10212 (N_10212,N_9883,N_9601);
and U10213 (N_10213,N_8750,N_9699);
or U10214 (N_10214,N_9729,N_9299);
nand U10215 (N_10215,N_9331,N_9029);
and U10216 (N_10216,N_9280,N_9272);
nand U10217 (N_10217,N_9096,N_9941);
nor U10218 (N_10218,N_9913,N_9596);
xor U10219 (N_10219,N_9713,N_9587);
xor U10220 (N_10220,N_9829,N_9662);
nor U10221 (N_10221,N_8778,N_9934);
nor U10222 (N_10222,N_9336,N_9524);
nor U10223 (N_10223,N_9397,N_9043);
xnor U10224 (N_10224,N_8839,N_9657);
or U10225 (N_10225,N_9326,N_9344);
xnor U10226 (N_10226,N_9586,N_8766);
nor U10227 (N_10227,N_9155,N_9602);
and U10228 (N_10228,N_9283,N_9748);
or U10229 (N_10229,N_9621,N_9027);
or U10230 (N_10230,N_9182,N_9156);
nor U10231 (N_10231,N_8804,N_9648);
or U10232 (N_10232,N_9497,N_9855);
nand U10233 (N_10233,N_9514,N_8772);
nand U10234 (N_10234,N_9338,N_9319);
nand U10235 (N_10235,N_9384,N_8850);
nor U10236 (N_10236,N_9347,N_9370);
or U10237 (N_10237,N_9117,N_8792);
and U10238 (N_10238,N_8783,N_9849);
nand U10239 (N_10239,N_9214,N_9487);
or U10240 (N_10240,N_9060,N_8845);
xnor U10241 (N_10241,N_8878,N_9068);
nor U10242 (N_10242,N_9286,N_9313);
nor U10243 (N_10243,N_9017,N_8789);
or U10244 (N_10244,N_9781,N_8971);
and U10245 (N_10245,N_9263,N_8918);
and U10246 (N_10246,N_9398,N_8823);
and U10247 (N_10247,N_9230,N_9209);
and U10248 (N_10248,N_9499,N_9980);
nand U10249 (N_10249,N_9614,N_9142);
xor U10250 (N_10250,N_8816,N_9502);
nor U10251 (N_10251,N_8790,N_9002);
nor U10252 (N_10252,N_9219,N_9656);
or U10253 (N_10253,N_8934,N_8836);
and U10254 (N_10254,N_9647,N_8830);
nor U10255 (N_10255,N_9861,N_9296);
or U10256 (N_10256,N_9690,N_8960);
xnor U10257 (N_10257,N_9968,N_9828);
nor U10258 (N_10258,N_9515,N_9419);
or U10259 (N_10259,N_9469,N_9083);
nand U10260 (N_10260,N_9366,N_9173);
nand U10261 (N_10261,N_9585,N_8870);
xnor U10262 (N_10262,N_9888,N_9239);
and U10263 (N_10263,N_9333,N_9498);
or U10264 (N_10264,N_9689,N_9335);
or U10265 (N_10265,N_9525,N_8925);
nand U10266 (N_10266,N_8865,N_9582);
nand U10267 (N_10267,N_9521,N_9433);
and U10268 (N_10268,N_9222,N_8780);
and U10269 (N_10269,N_9807,N_9638);
or U10270 (N_10270,N_8930,N_9925);
nor U10271 (N_10271,N_8852,N_9072);
or U10272 (N_10272,N_8966,N_8849);
nor U10273 (N_10273,N_8903,N_9059);
xor U10274 (N_10274,N_9912,N_9898);
nor U10275 (N_10275,N_9427,N_9853);
and U10276 (N_10276,N_9964,N_9046);
or U10277 (N_10277,N_9652,N_8972);
xnor U10278 (N_10278,N_8965,N_9863);
or U10279 (N_10279,N_9001,N_9052);
nand U10280 (N_10280,N_9554,N_8899);
xnor U10281 (N_10281,N_9458,N_8975);
and U10282 (N_10282,N_9728,N_9947);
and U10283 (N_10283,N_8888,N_9550);
and U10284 (N_10284,N_8967,N_9756);
or U10285 (N_10285,N_9045,N_9952);
xnor U10286 (N_10286,N_9896,N_9357);
or U10287 (N_10287,N_9907,N_9714);
nand U10288 (N_10288,N_9198,N_9873);
xor U10289 (N_10289,N_8808,N_9613);
nand U10290 (N_10290,N_8765,N_8791);
and U10291 (N_10291,N_9801,N_9918);
nor U10292 (N_10292,N_9901,N_8997);
and U10293 (N_10293,N_8896,N_9903);
and U10294 (N_10294,N_9658,N_9109);
and U10295 (N_10295,N_9719,N_9724);
nand U10296 (N_10296,N_9208,N_9457);
nor U10297 (N_10297,N_9070,N_8901);
xnor U10298 (N_10298,N_9938,N_9921);
xnor U10299 (N_10299,N_9233,N_8837);
or U10300 (N_10300,N_9342,N_9862);
xor U10301 (N_10301,N_9664,N_9261);
nor U10302 (N_10302,N_9451,N_8763);
and U10303 (N_10303,N_9382,N_9681);
and U10304 (N_10304,N_9851,N_9305);
or U10305 (N_10305,N_9987,N_8874);
xor U10306 (N_10306,N_9951,N_9692);
nand U10307 (N_10307,N_9598,N_9449);
nand U10308 (N_10308,N_9328,N_9906);
and U10309 (N_10309,N_8818,N_9997);
xor U10310 (N_10310,N_9776,N_9735);
and U10311 (N_10311,N_9365,N_9579);
nor U10312 (N_10312,N_9961,N_8961);
nand U10313 (N_10313,N_9838,N_9623);
nor U10314 (N_10314,N_8770,N_9541);
xor U10315 (N_10315,N_9144,N_8797);
nor U10316 (N_10316,N_9886,N_9431);
nor U10317 (N_10317,N_9798,N_9734);
nor U10318 (N_10318,N_9618,N_9084);
nor U10319 (N_10319,N_9577,N_9995);
nand U10320 (N_10320,N_9453,N_9773);
nand U10321 (N_10321,N_9847,N_9341);
and U10322 (N_10322,N_8963,N_9683);
xnor U10323 (N_10323,N_9537,N_9289);
or U10324 (N_10324,N_9411,N_9872);
xor U10325 (N_10325,N_8929,N_9291);
xnor U10326 (N_10326,N_8857,N_8764);
nand U10327 (N_10327,N_9085,N_9307);
xnor U10328 (N_10328,N_9023,N_9977);
and U10329 (N_10329,N_9034,N_9227);
or U10330 (N_10330,N_9538,N_9148);
and U10331 (N_10331,N_9920,N_8801);
or U10332 (N_10332,N_9330,N_9762);
and U10333 (N_10333,N_8989,N_9041);
and U10334 (N_10334,N_8811,N_9013);
or U10335 (N_10335,N_9529,N_8970);
nand U10336 (N_10336,N_9857,N_9573);
or U10337 (N_10337,N_9764,N_9971);
nand U10338 (N_10338,N_9758,N_9014);
nor U10339 (N_10339,N_8942,N_9007);
or U10340 (N_10340,N_9510,N_8877);
xor U10341 (N_10341,N_9817,N_9755);
or U10342 (N_10342,N_9607,N_9774);
and U10343 (N_10343,N_9882,N_9484);
and U10344 (N_10344,N_9371,N_9037);
xor U10345 (N_10345,N_9047,N_9545);
and U10346 (N_10346,N_9819,N_8868);
and U10347 (N_10347,N_8983,N_8881);
and U10348 (N_10348,N_9534,N_9500);
xor U10349 (N_10349,N_9994,N_9243);
or U10350 (N_10350,N_9164,N_9273);
xnor U10351 (N_10351,N_8904,N_9536);
and U10352 (N_10352,N_8898,N_9785);
nor U10353 (N_10353,N_9376,N_9435);
or U10354 (N_10354,N_9074,N_9702);
nand U10355 (N_10355,N_9375,N_9868);
and U10356 (N_10356,N_8835,N_9973);
nor U10357 (N_10357,N_9789,N_8873);
and U10358 (N_10358,N_8885,N_9540);
nand U10359 (N_10359,N_9818,N_9902);
nor U10360 (N_10360,N_9158,N_9434);
xor U10361 (N_10361,N_9351,N_9942);
xnor U10362 (N_10362,N_9404,N_9069);
or U10363 (N_10363,N_8879,N_9615);
nand U10364 (N_10364,N_9867,N_9840);
nor U10365 (N_10365,N_9094,N_9894);
nand U10366 (N_10366,N_9193,N_9489);
nand U10367 (N_10367,N_9270,N_8981);
nand U10368 (N_10368,N_9175,N_9483);
and U10369 (N_10369,N_9183,N_8841);
xnor U10370 (N_10370,N_9804,N_9644);
nand U10371 (N_10371,N_9119,N_9606);
nand U10372 (N_10372,N_8771,N_9295);
nor U10373 (N_10373,N_9528,N_9557);
xor U10374 (N_10374,N_9162,N_9716);
or U10375 (N_10375,N_9167,N_9140);
xnor U10376 (N_10376,N_9822,N_9242);
or U10377 (N_10377,N_9895,N_8940);
and U10378 (N_10378,N_9900,N_9749);
or U10379 (N_10379,N_9646,N_9595);
nand U10380 (N_10380,N_9334,N_9108);
or U10381 (N_10381,N_9309,N_9643);
nor U10382 (N_10382,N_9088,N_9260);
and U10383 (N_10383,N_9432,N_9563);
xor U10384 (N_10384,N_9950,N_9195);
and U10385 (N_10385,N_8785,N_8996);
and U10386 (N_10386,N_9244,N_9120);
nand U10387 (N_10387,N_9686,N_9697);
xnor U10388 (N_10388,N_9292,N_9680);
xor U10389 (N_10389,N_9349,N_9255);
or U10390 (N_10390,N_9262,N_9710);
and U10391 (N_10391,N_9556,N_8754);
and U10392 (N_10392,N_9293,N_9870);
or U10393 (N_10393,N_9943,N_8756);
xnor U10394 (N_10394,N_9949,N_9767);
or U10395 (N_10395,N_9276,N_9205);
and U10396 (N_10396,N_9632,N_8784);
nor U10397 (N_10397,N_9665,N_9929);
nand U10398 (N_10398,N_9899,N_9207);
or U10399 (N_10399,N_9253,N_9816);
or U10400 (N_10400,N_8864,N_9030);
nor U10401 (N_10401,N_9924,N_9154);
and U10402 (N_10402,N_9424,N_9297);
nor U10403 (N_10403,N_9461,N_9055);
xnor U10404 (N_10404,N_9275,N_9329);
nand U10405 (N_10405,N_8820,N_9325);
nand U10406 (N_10406,N_9303,N_8889);
nor U10407 (N_10407,N_9380,N_9935);
xor U10408 (N_10408,N_9360,N_8969);
or U10409 (N_10409,N_9576,N_9186);
and U10410 (N_10410,N_9990,N_9097);
and U10411 (N_10411,N_8895,N_9036);
or U10412 (N_10412,N_8767,N_9777);
or U10413 (N_10413,N_9012,N_9495);
and U10414 (N_10414,N_9475,N_8900);
xor U10415 (N_10415,N_9723,N_9628);
and U10416 (N_10416,N_9231,N_9226);
and U10417 (N_10417,N_8897,N_9439);
nand U10418 (N_10418,N_9463,N_9551);
or U10419 (N_10419,N_9421,N_9259);
or U10420 (N_10420,N_9693,N_9408);
nand U10421 (N_10421,N_9210,N_8926);
xor U10422 (N_10422,N_8979,N_9402);
nor U10423 (N_10423,N_8848,N_9864);
nor U10424 (N_10424,N_9927,N_9221);
or U10425 (N_10425,N_9999,N_8793);
or U10426 (N_10426,N_9322,N_9832);
xnor U10427 (N_10427,N_9917,N_9494);
nand U10428 (N_10428,N_9076,N_9316);
xor U10429 (N_10429,N_8752,N_9522);
or U10430 (N_10430,N_8786,N_9611);
nand U10431 (N_10431,N_9425,N_9552);
or U10432 (N_10432,N_9079,N_8800);
and U10433 (N_10433,N_9352,N_9592);
and U10434 (N_10434,N_9151,N_9266);
and U10435 (N_10435,N_9218,N_9470);
nor U10436 (N_10436,N_9038,N_8875);
nor U10437 (N_10437,N_9637,N_9617);
nand U10438 (N_10438,N_8796,N_9181);
xnor U10439 (N_10439,N_9377,N_9824);
nand U10440 (N_10440,N_9520,N_9254);
nor U10441 (N_10441,N_8826,N_9978);
and U10442 (N_10442,N_9678,N_9020);
nor U10443 (N_10443,N_9629,N_9268);
or U10444 (N_10444,N_9603,N_9583);
nand U10445 (N_10445,N_9671,N_9464);
and U10446 (N_10446,N_9471,N_8860);
nand U10447 (N_10447,N_9711,N_8933);
nand U10448 (N_10448,N_9185,N_9416);
xor U10449 (N_10449,N_9948,N_9149);
or U10450 (N_10450,N_9530,N_9446);
or U10451 (N_10451,N_9659,N_9575);
or U10452 (N_10452,N_9753,N_9159);
nand U10453 (N_10453,N_9770,N_9696);
xor U10454 (N_10454,N_8798,N_9889);
nand U10455 (N_10455,N_9062,N_9937);
or U10456 (N_10456,N_9107,N_8779);
or U10457 (N_10457,N_9392,N_9531);
nand U10458 (N_10458,N_9339,N_8894);
nand U10459 (N_10459,N_9996,N_9821);
nor U10460 (N_10460,N_9771,N_9981);
or U10461 (N_10461,N_9406,N_8803);
xnor U10462 (N_10462,N_9468,N_9679);
nand U10463 (N_10463,N_9220,N_9031);
xor U10464 (N_10464,N_9163,N_9672);
or U10465 (N_10465,N_9032,N_8819);
or U10466 (N_10466,N_8914,N_8993);
nor U10467 (N_10467,N_9639,N_9125);
and U10468 (N_10468,N_9549,N_9067);
nor U10469 (N_10469,N_8842,N_9962);
nand U10470 (N_10470,N_9403,N_9100);
or U10471 (N_10471,N_9860,N_9932);
nand U10472 (N_10472,N_9548,N_8884);
nand U10473 (N_10473,N_9763,N_9203);
xnor U10474 (N_10474,N_9513,N_9256);
nor U10475 (N_10475,N_9340,N_8753);
or U10476 (N_10476,N_9991,N_9688);
nor U10477 (N_10477,N_9940,N_9139);
xor U10478 (N_10478,N_8760,N_9833);
or U10479 (N_10479,N_9015,N_9746);
nand U10480 (N_10480,N_9126,N_8834);
or U10481 (N_10481,N_9407,N_9936);
nor U10482 (N_10482,N_9445,N_9372);
or U10483 (N_10483,N_9675,N_9788);
nand U10484 (N_10484,N_8987,N_9252);
xnor U10485 (N_10485,N_9304,N_9908);
or U10486 (N_10486,N_8794,N_9553);
xnor U10487 (N_10487,N_8880,N_9780);
nand U10488 (N_10488,N_9479,N_8774);
xor U10489 (N_10489,N_9415,N_8777);
nor U10490 (N_10490,N_9919,N_9315);
nand U10491 (N_10491,N_9212,N_8856);
nand U10492 (N_10492,N_9507,N_9301);
xor U10493 (N_10493,N_8919,N_8768);
and U10494 (N_10494,N_9122,N_9024);
and U10495 (N_10495,N_9265,N_8906);
and U10496 (N_10496,N_9153,N_9177);
nor U10497 (N_10497,N_9633,N_9926);
nand U10498 (N_10498,N_9213,N_9466);
or U10499 (N_10499,N_9401,N_9892);
and U10500 (N_10500,N_8927,N_9066);
nor U10501 (N_10501,N_9765,N_9527);
xnor U10502 (N_10502,N_9944,N_9604);
xnor U10503 (N_10503,N_9217,N_9584);
nor U10504 (N_10504,N_9532,N_9040);
and U10505 (N_10505,N_9492,N_8762);
nand U10506 (N_10506,N_9438,N_9414);
and U10507 (N_10507,N_9841,N_9008);
nor U10508 (N_10508,N_9115,N_9827);
or U10509 (N_10509,N_8758,N_9879);
and U10510 (N_10510,N_9503,N_9709);
or U10511 (N_10511,N_9744,N_8847);
nand U10512 (N_10512,N_9965,N_9923);
nand U10513 (N_10513,N_8977,N_9200);
and U10514 (N_10514,N_9701,N_9240);
xor U10515 (N_10515,N_9640,N_9178);
and U10516 (N_10516,N_9123,N_9570);
nor U10517 (N_10517,N_9274,N_9196);
nor U10518 (N_10518,N_9174,N_9704);
xnor U10519 (N_10519,N_9846,N_9850);
nand U10520 (N_10520,N_9298,N_9954);
nor U10521 (N_10521,N_9452,N_9715);
nor U10522 (N_10522,N_8817,N_9597);
or U10523 (N_10523,N_8948,N_9547);
nor U10524 (N_10524,N_9075,N_9237);
xnor U10525 (N_10525,N_8941,N_8802);
xor U10526 (N_10526,N_9745,N_9327);
and U10527 (N_10527,N_9320,N_9450);
or U10528 (N_10528,N_9114,N_9512);
nand U10529 (N_10529,N_9569,N_9294);
nor U10530 (N_10530,N_9061,N_9979);
or U10531 (N_10531,N_8853,N_9473);
or U10532 (N_10532,N_9417,N_9033);
or U10533 (N_10533,N_9775,N_8810);
or U10534 (N_10534,N_9201,N_9976);
or U10535 (N_10535,N_9815,N_9641);
nand U10536 (N_10536,N_9343,N_9787);
xor U10537 (N_10537,N_9318,N_9682);
or U10538 (N_10538,N_8833,N_8935);
or U10539 (N_10539,N_9837,N_9223);
nand U10540 (N_10540,N_9516,N_9636);
xnor U10541 (N_10541,N_9778,N_9843);
nand U10542 (N_10542,N_9795,N_9668);
nor U10543 (N_10543,N_9362,N_9395);
nor U10544 (N_10544,N_9051,N_9653);
xor U10545 (N_10545,N_9447,N_9743);
xnor U10546 (N_10546,N_9992,N_9359);
and U10547 (N_10547,N_9003,N_9695);
xor U10548 (N_10548,N_9160,N_9630);
xor U10549 (N_10549,N_9026,N_8909);
nand U10550 (N_10550,N_9572,N_9786);
nand U10551 (N_10551,N_8846,N_8858);
xnor U10552 (N_10552,N_8998,N_9784);
xnor U10553 (N_10553,N_9152,N_9871);
nand U10554 (N_10554,N_9759,N_9610);
and U10555 (N_10555,N_8917,N_9103);
or U10556 (N_10556,N_9418,N_8751);
or U10557 (N_10557,N_9211,N_8782);
xor U10558 (N_10558,N_9739,N_9350);
or U10559 (N_10559,N_9933,N_9717);
nand U10560 (N_10560,N_9454,N_9010);
xnor U10561 (N_10561,N_9379,N_9877);
and U10562 (N_10562,N_8825,N_8921);
or U10563 (N_10563,N_9127,N_9559);
and U10564 (N_10564,N_9288,N_9591);
or U10565 (N_10565,N_8886,N_9364);
nand U10566 (N_10566,N_8956,N_9021);
nand U10567 (N_10567,N_8973,N_9000);
and U10568 (N_10568,N_8809,N_9810);
nor U10569 (N_10569,N_8832,N_9930);
xnor U10570 (N_10570,N_9959,N_9204);
nor U10571 (N_10571,N_9134,N_9508);
xnor U10572 (N_10572,N_9820,N_9073);
or U10573 (N_10573,N_9835,N_9655);
and U10574 (N_10574,N_9166,N_9738);
and U10575 (N_10575,N_9974,N_9546);
nor U10576 (N_10576,N_9137,N_9367);
nor U10577 (N_10577,N_9306,N_9793);
xor U10578 (N_10578,N_9099,N_9128);
xnor U10579 (N_10579,N_9517,N_9797);
or U10580 (N_10580,N_9574,N_9566);
and U10581 (N_10581,N_9691,N_9105);
and U10582 (N_10582,N_8829,N_9511);
and U10583 (N_10583,N_8945,N_9131);
nand U10584 (N_10584,N_9707,N_9904);
xnor U10585 (N_10585,N_8815,N_9642);
nor U10586 (N_10586,N_9612,N_9844);
and U10587 (N_10587,N_9422,N_9480);
nand U10588 (N_10588,N_9247,N_9050);
and U10589 (N_10589,N_9179,N_9459);
xnor U10590 (N_10590,N_9783,N_9246);
or U10591 (N_10591,N_9393,N_9988);
nand U10592 (N_10592,N_9874,N_9248);
and U10593 (N_10593,N_9969,N_9830);
and U10594 (N_10594,N_9460,N_9121);
or U10595 (N_10595,N_9090,N_8944);
and U10596 (N_10596,N_9428,N_9939);
and U10597 (N_10597,N_8838,N_9095);
or U10598 (N_10598,N_8840,N_9865);
nor U10599 (N_10599,N_9485,N_9271);
and U10600 (N_10600,N_9310,N_9627);
and U10601 (N_10601,N_9245,N_9093);
or U10602 (N_10602,N_8781,N_9448);
xnor U10603 (N_10603,N_9281,N_8854);
nor U10604 (N_10604,N_9986,N_8788);
nor U10605 (N_10605,N_9975,N_9132);
or U10606 (N_10606,N_9543,N_9814);
xnor U10607 (N_10607,N_8814,N_9730);
nand U10608 (N_10608,N_9794,N_9150);
nand U10609 (N_10609,N_9677,N_9373);
xor U10610 (N_10610,N_9078,N_9625);
or U10611 (N_10611,N_8887,N_9823);
and U10612 (N_10612,N_9982,N_8955);
nand U10613 (N_10613,N_9726,N_9624);
xor U10614 (N_10614,N_8813,N_9082);
or U10615 (N_10615,N_9486,N_9071);
and U10616 (N_10616,N_8859,N_9542);
xnor U10617 (N_10617,N_9145,N_9805);
nand U10618 (N_10618,N_9567,N_9859);
or U10619 (N_10619,N_9685,N_9025);
nor U10620 (N_10620,N_9698,N_8910);
xor U10621 (N_10621,N_9588,N_9481);
xnor U10622 (N_10622,N_9229,N_9323);
and U10623 (N_10623,N_9249,N_9478);
and U10624 (N_10624,N_9504,N_9113);
nand U10625 (N_10625,N_8846,N_8929);
or U10626 (N_10626,N_9537,N_9368);
nand U10627 (N_10627,N_9107,N_9281);
or U10628 (N_10628,N_9976,N_8944);
xnor U10629 (N_10629,N_9497,N_9300);
and U10630 (N_10630,N_8788,N_9303);
and U10631 (N_10631,N_8767,N_9478);
and U10632 (N_10632,N_9622,N_9323);
xor U10633 (N_10633,N_8848,N_9702);
and U10634 (N_10634,N_8784,N_9854);
or U10635 (N_10635,N_8770,N_9386);
nand U10636 (N_10636,N_9431,N_9940);
xnor U10637 (N_10637,N_9178,N_9331);
nand U10638 (N_10638,N_9729,N_9781);
and U10639 (N_10639,N_8890,N_8877);
nand U10640 (N_10640,N_8978,N_8841);
xor U10641 (N_10641,N_9552,N_9123);
nand U10642 (N_10642,N_9333,N_9600);
nand U10643 (N_10643,N_9856,N_9102);
and U10644 (N_10644,N_9445,N_8750);
nand U10645 (N_10645,N_9712,N_9984);
xnor U10646 (N_10646,N_9681,N_9732);
nor U10647 (N_10647,N_9678,N_9907);
and U10648 (N_10648,N_9821,N_9856);
nand U10649 (N_10649,N_9285,N_9626);
nand U10650 (N_10650,N_9605,N_9341);
nand U10651 (N_10651,N_8939,N_9841);
and U10652 (N_10652,N_9797,N_9237);
or U10653 (N_10653,N_9918,N_9084);
and U10654 (N_10654,N_9057,N_9825);
nor U10655 (N_10655,N_8801,N_9648);
xnor U10656 (N_10656,N_9886,N_8824);
and U10657 (N_10657,N_9511,N_9569);
xor U10658 (N_10658,N_9478,N_9577);
nand U10659 (N_10659,N_9449,N_9869);
nand U10660 (N_10660,N_9597,N_8863);
and U10661 (N_10661,N_8856,N_9163);
nand U10662 (N_10662,N_8924,N_9373);
xnor U10663 (N_10663,N_9271,N_9648);
or U10664 (N_10664,N_9301,N_8953);
nand U10665 (N_10665,N_9860,N_9110);
or U10666 (N_10666,N_9527,N_9644);
and U10667 (N_10667,N_9398,N_9433);
nor U10668 (N_10668,N_9082,N_9001);
xnor U10669 (N_10669,N_9763,N_9678);
and U10670 (N_10670,N_8958,N_9720);
xnor U10671 (N_10671,N_9701,N_9699);
nand U10672 (N_10672,N_9843,N_9812);
nand U10673 (N_10673,N_8799,N_9351);
nand U10674 (N_10674,N_8828,N_8976);
xnor U10675 (N_10675,N_8945,N_8973);
or U10676 (N_10676,N_9514,N_9864);
or U10677 (N_10677,N_9067,N_9070);
or U10678 (N_10678,N_8852,N_9606);
or U10679 (N_10679,N_9473,N_9358);
xnor U10680 (N_10680,N_9601,N_8993);
or U10681 (N_10681,N_9508,N_9109);
or U10682 (N_10682,N_9210,N_9225);
nor U10683 (N_10683,N_9775,N_9425);
or U10684 (N_10684,N_9284,N_8914);
and U10685 (N_10685,N_9880,N_9295);
xnor U10686 (N_10686,N_9834,N_9344);
nor U10687 (N_10687,N_9085,N_9012);
or U10688 (N_10688,N_8837,N_9512);
and U10689 (N_10689,N_9596,N_9882);
or U10690 (N_10690,N_9693,N_9013);
or U10691 (N_10691,N_9812,N_9291);
nor U10692 (N_10692,N_9084,N_9490);
and U10693 (N_10693,N_8962,N_9510);
or U10694 (N_10694,N_9912,N_9712);
nand U10695 (N_10695,N_9299,N_8835);
xnor U10696 (N_10696,N_9100,N_9476);
xor U10697 (N_10697,N_9722,N_9094);
or U10698 (N_10698,N_9516,N_9880);
or U10699 (N_10699,N_9000,N_8888);
and U10700 (N_10700,N_9847,N_8939);
nor U10701 (N_10701,N_9737,N_8795);
nor U10702 (N_10702,N_8929,N_8927);
xor U10703 (N_10703,N_8913,N_9194);
xnor U10704 (N_10704,N_8829,N_9334);
xor U10705 (N_10705,N_9338,N_9361);
or U10706 (N_10706,N_9998,N_9231);
nand U10707 (N_10707,N_9949,N_9035);
nor U10708 (N_10708,N_9297,N_9374);
nor U10709 (N_10709,N_9743,N_9320);
or U10710 (N_10710,N_9084,N_9156);
and U10711 (N_10711,N_8978,N_9425);
and U10712 (N_10712,N_9501,N_9056);
xnor U10713 (N_10713,N_9272,N_9311);
nand U10714 (N_10714,N_8778,N_9061);
xnor U10715 (N_10715,N_9063,N_9732);
and U10716 (N_10716,N_8996,N_8825);
nor U10717 (N_10717,N_9862,N_9642);
xor U10718 (N_10718,N_9861,N_9074);
nor U10719 (N_10719,N_9451,N_9049);
xor U10720 (N_10720,N_9938,N_9508);
and U10721 (N_10721,N_9008,N_9103);
nand U10722 (N_10722,N_9292,N_9393);
and U10723 (N_10723,N_9272,N_9888);
or U10724 (N_10724,N_8821,N_9910);
or U10725 (N_10725,N_9773,N_9836);
xnor U10726 (N_10726,N_9118,N_9105);
and U10727 (N_10727,N_9557,N_9814);
or U10728 (N_10728,N_9004,N_9922);
and U10729 (N_10729,N_9473,N_9398);
xor U10730 (N_10730,N_9176,N_9074);
nand U10731 (N_10731,N_9392,N_9180);
xnor U10732 (N_10732,N_9541,N_9190);
or U10733 (N_10733,N_9750,N_9621);
nor U10734 (N_10734,N_9842,N_9689);
and U10735 (N_10735,N_9523,N_8940);
nand U10736 (N_10736,N_9687,N_9328);
nor U10737 (N_10737,N_9238,N_9359);
and U10738 (N_10738,N_9617,N_9373);
nand U10739 (N_10739,N_9435,N_9585);
or U10740 (N_10740,N_9321,N_9150);
and U10741 (N_10741,N_9443,N_9287);
or U10742 (N_10742,N_8830,N_9105);
and U10743 (N_10743,N_9005,N_8770);
nand U10744 (N_10744,N_8796,N_9414);
xnor U10745 (N_10745,N_9176,N_9936);
xnor U10746 (N_10746,N_9539,N_9534);
or U10747 (N_10747,N_9407,N_9708);
nor U10748 (N_10748,N_8916,N_9290);
and U10749 (N_10749,N_9430,N_9058);
or U10750 (N_10750,N_9232,N_9533);
or U10751 (N_10751,N_9205,N_9982);
or U10752 (N_10752,N_9847,N_9137);
or U10753 (N_10753,N_9331,N_9513);
nor U10754 (N_10754,N_9469,N_9453);
nand U10755 (N_10755,N_9586,N_9060);
nor U10756 (N_10756,N_8791,N_9154);
nand U10757 (N_10757,N_8793,N_9195);
or U10758 (N_10758,N_9385,N_9168);
xor U10759 (N_10759,N_9274,N_8802);
nor U10760 (N_10760,N_9977,N_9231);
or U10761 (N_10761,N_9791,N_8856);
xor U10762 (N_10762,N_8944,N_9427);
and U10763 (N_10763,N_9012,N_9894);
and U10764 (N_10764,N_9131,N_9573);
nor U10765 (N_10765,N_9492,N_8929);
xor U10766 (N_10766,N_9704,N_8817);
nor U10767 (N_10767,N_9114,N_9459);
nand U10768 (N_10768,N_8794,N_8784);
nand U10769 (N_10769,N_9454,N_9571);
nor U10770 (N_10770,N_8913,N_9697);
or U10771 (N_10771,N_9506,N_9345);
or U10772 (N_10772,N_8984,N_9227);
or U10773 (N_10773,N_9305,N_9939);
nor U10774 (N_10774,N_8821,N_9262);
nor U10775 (N_10775,N_9944,N_9129);
and U10776 (N_10776,N_9247,N_9460);
and U10777 (N_10777,N_9791,N_9057);
nand U10778 (N_10778,N_9402,N_9551);
or U10779 (N_10779,N_9794,N_9406);
xnor U10780 (N_10780,N_8873,N_8917);
nand U10781 (N_10781,N_9376,N_9550);
and U10782 (N_10782,N_8959,N_8824);
xor U10783 (N_10783,N_9339,N_9563);
nor U10784 (N_10784,N_9527,N_9946);
nand U10785 (N_10785,N_9300,N_8800);
xor U10786 (N_10786,N_8938,N_8817);
or U10787 (N_10787,N_9682,N_9189);
nor U10788 (N_10788,N_9434,N_9285);
and U10789 (N_10789,N_8976,N_9730);
xnor U10790 (N_10790,N_9526,N_9300);
or U10791 (N_10791,N_9903,N_9620);
and U10792 (N_10792,N_8948,N_9534);
nor U10793 (N_10793,N_9633,N_9111);
nor U10794 (N_10794,N_9745,N_9728);
nor U10795 (N_10795,N_9089,N_9050);
and U10796 (N_10796,N_9175,N_8872);
and U10797 (N_10797,N_9745,N_9297);
nor U10798 (N_10798,N_9704,N_8795);
xnor U10799 (N_10799,N_9147,N_9893);
nand U10800 (N_10800,N_9280,N_8961);
nand U10801 (N_10801,N_9761,N_8921);
and U10802 (N_10802,N_9641,N_9464);
or U10803 (N_10803,N_9560,N_9048);
nor U10804 (N_10804,N_9022,N_9172);
nor U10805 (N_10805,N_9374,N_9553);
or U10806 (N_10806,N_9129,N_9863);
and U10807 (N_10807,N_9802,N_9331);
and U10808 (N_10808,N_9949,N_9066);
nor U10809 (N_10809,N_8934,N_8883);
nor U10810 (N_10810,N_9806,N_9641);
nor U10811 (N_10811,N_9273,N_9184);
nor U10812 (N_10812,N_9739,N_9296);
nand U10813 (N_10813,N_8761,N_9445);
nand U10814 (N_10814,N_8949,N_9282);
or U10815 (N_10815,N_9090,N_8892);
nand U10816 (N_10816,N_8772,N_9888);
and U10817 (N_10817,N_9744,N_8913);
nand U10818 (N_10818,N_9189,N_9004);
nand U10819 (N_10819,N_9450,N_9188);
or U10820 (N_10820,N_9414,N_9949);
nor U10821 (N_10821,N_8870,N_9186);
or U10822 (N_10822,N_9069,N_9816);
nor U10823 (N_10823,N_9971,N_9354);
or U10824 (N_10824,N_8763,N_9682);
nand U10825 (N_10825,N_9905,N_9085);
and U10826 (N_10826,N_9819,N_9163);
and U10827 (N_10827,N_9922,N_8824);
nand U10828 (N_10828,N_9191,N_9918);
and U10829 (N_10829,N_9482,N_9224);
nor U10830 (N_10830,N_9228,N_9638);
nand U10831 (N_10831,N_9779,N_9657);
or U10832 (N_10832,N_9658,N_9416);
and U10833 (N_10833,N_9616,N_9900);
and U10834 (N_10834,N_9062,N_9947);
or U10835 (N_10835,N_9907,N_9847);
or U10836 (N_10836,N_8862,N_9611);
nor U10837 (N_10837,N_8788,N_9454);
xor U10838 (N_10838,N_8843,N_8952);
nand U10839 (N_10839,N_9790,N_9686);
nand U10840 (N_10840,N_9947,N_9792);
nor U10841 (N_10841,N_9767,N_9271);
or U10842 (N_10842,N_9136,N_8780);
and U10843 (N_10843,N_9113,N_9941);
nor U10844 (N_10844,N_9988,N_9589);
xor U10845 (N_10845,N_9916,N_9509);
or U10846 (N_10846,N_9686,N_9010);
nor U10847 (N_10847,N_9719,N_9218);
or U10848 (N_10848,N_9317,N_8916);
nand U10849 (N_10849,N_9043,N_9895);
or U10850 (N_10850,N_9651,N_9977);
nor U10851 (N_10851,N_9333,N_9803);
nand U10852 (N_10852,N_9589,N_9978);
and U10853 (N_10853,N_9305,N_8920);
xor U10854 (N_10854,N_8805,N_9065);
and U10855 (N_10855,N_9200,N_9959);
and U10856 (N_10856,N_9689,N_9188);
xor U10857 (N_10857,N_9346,N_9451);
nor U10858 (N_10858,N_9803,N_9442);
nor U10859 (N_10859,N_9748,N_9345);
nand U10860 (N_10860,N_9061,N_8997);
nor U10861 (N_10861,N_8877,N_8778);
nor U10862 (N_10862,N_8941,N_9261);
or U10863 (N_10863,N_9463,N_9445);
xnor U10864 (N_10864,N_9568,N_9670);
nand U10865 (N_10865,N_9013,N_9870);
xnor U10866 (N_10866,N_9938,N_8955);
xnor U10867 (N_10867,N_9587,N_9187);
xnor U10868 (N_10868,N_8799,N_9452);
nor U10869 (N_10869,N_8827,N_9012);
nor U10870 (N_10870,N_9605,N_8876);
or U10871 (N_10871,N_9626,N_9936);
nand U10872 (N_10872,N_9746,N_9193);
or U10873 (N_10873,N_9380,N_9015);
and U10874 (N_10874,N_9279,N_8937);
nor U10875 (N_10875,N_9339,N_9500);
nor U10876 (N_10876,N_9469,N_8999);
nor U10877 (N_10877,N_9610,N_9972);
xnor U10878 (N_10878,N_9985,N_9220);
and U10879 (N_10879,N_9918,N_8841);
nand U10880 (N_10880,N_9362,N_8862);
xnor U10881 (N_10881,N_8864,N_9144);
and U10882 (N_10882,N_9836,N_9871);
nand U10883 (N_10883,N_9055,N_9341);
and U10884 (N_10884,N_9078,N_9682);
and U10885 (N_10885,N_8825,N_9309);
xnor U10886 (N_10886,N_9136,N_8833);
or U10887 (N_10887,N_9869,N_9222);
or U10888 (N_10888,N_9485,N_9314);
and U10889 (N_10889,N_9794,N_9927);
xor U10890 (N_10890,N_9788,N_9650);
nor U10891 (N_10891,N_9832,N_9617);
or U10892 (N_10892,N_9310,N_9364);
xor U10893 (N_10893,N_9036,N_9747);
nor U10894 (N_10894,N_9695,N_9873);
xnor U10895 (N_10895,N_9426,N_9515);
nand U10896 (N_10896,N_9339,N_9631);
nand U10897 (N_10897,N_9442,N_9508);
nand U10898 (N_10898,N_9623,N_9398);
nor U10899 (N_10899,N_9093,N_9660);
xnor U10900 (N_10900,N_9406,N_9233);
xor U10901 (N_10901,N_8957,N_9050);
nand U10902 (N_10902,N_9760,N_9939);
xor U10903 (N_10903,N_9443,N_9424);
or U10904 (N_10904,N_9591,N_8858);
nand U10905 (N_10905,N_9167,N_9360);
and U10906 (N_10906,N_9323,N_8763);
and U10907 (N_10907,N_9047,N_9903);
nor U10908 (N_10908,N_9267,N_9553);
and U10909 (N_10909,N_9293,N_9449);
xor U10910 (N_10910,N_9660,N_9755);
nand U10911 (N_10911,N_9353,N_8986);
xnor U10912 (N_10912,N_9709,N_9483);
or U10913 (N_10913,N_8956,N_9225);
nand U10914 (N_10914,N_9089,N_9276);
or U10915 (N_10915,N_9482,N_8928);
nor U10916 (N_10916,N_8841,N_9761);
xnor U10917 (N_10917,N_8755,N_9313);
nor U10918 (N_10918,N_9222,N_8822);
nor U10919 (N_10919,N_8804,N_9029);
nand U10920 (N_10920,N_9219,N_9652);
and U10921 (N_10921,N_9399,N_8960);
xor U10922 (N_10922,N_8869,N_9915);
and U10923 (N_10923,N_9887,N_9927);
or U10924 (N_10924,N_9704,N_9261);
xor U10925 (N_10925,N_9168,N_9010);
or U10926 (N_10926,N_9863,N_9481);
and U10927 (N_10927,N_8818,N_8874);
nand U10928 (N_10928,N_9425,N_8940);
nor U10929 (N_10929,N_9689,N_9953);
nand U10930 (N_10930,N_9931,N_9834);
nand U10931 (N_10931,N_9882,N_9766);
nand U10932 (N_10932,N_9273,N_9103);
nor U10933 (N_10933,N_9495,N_9870);
or U10934 (N_10934,N_9722,N_9671);
and U10935 (N_10935,N_9057,N_9871);
xnor U10936 (N_10936,N_8900,N_9830);
or U10937 (N_10937,N_9678,N_9768);
nand U10938 (N_10938,N_9116,N_8884);
nor U10939 (N_10939,N_9043,N_9135);
xnor U10940 (N_10940,N_8855,N_8874);
xor U10941 (N_10941,N_9750,N_9821);
nor U10942 (N_10942,N_9261,N_9730);
nor U10943 (N_10943,N_9416,N_9150);
xor U10944 (N_10944,N_9678,N_9255);
and U10945 (N_10945,N_9588,N_8926);
xnor U10946 (N_10946,N_9751,N_9781);
or U10947 (N_10947,N_8907,N_8811);
xnor U10948 (N_10948,N_9853,N_8954);
xor U10949 (N_10949,N_9435,N_9324);
nor U10950 (N_10950,N_9073,N_9205);
and U10951 (N_10951,N_8873,N_9486);
xor U10952 (N_10952,N_9209,N_9062);
xor U10953 (N_10953,N_9838,N_9785);
nor U10954 (N_10954,N_9814,N_9714);
or U10955 (N_10955,N_9875,N_9131);
and U10956 (N_10956,N_9784,N_9235);
and U10957 (N_10957,N_9489,N_8840);
and U10958 (N_10958,N_9347,N_9105);
nand U10959 (N_10959,N_9882,N_9138);
nor U10960 (N_10960,N_9685,N_9167);
nor U10961 (N_10961,N_9634,N_9834);
nand U10962 (N_10962,N_9722,N_9246);
or U10963 (N_10963,N_9609,N_9719);
and U10964 (N_10964,N_9776,N_9075);
or U10965 (N_10965,N_8798,N_9367);
or U10966 (N_10966,N_9933,N_9011);
nand U10967 (N_10967,N_9109,N_9421);
nor U10968 (N_10968,N_9832,N_9113);
nand U10969 (N_10969,N_9038,N_9005);
nor U10970 (N_10970,N_9978,N_9411);
nor U10971 (N_10971,N_9424,N_9304);
or U10972 (N_10972,N_9200,N_8771);
xor U10973 (N_10973,N_8858,N_8797);
nor U10974 (N_10974,N_9128,N_9522);
nand U10975 (N_10975,N_9217,N_9453);
nor U10976 (N_10976,N_8911,N_8789);
and U10977 (N_10977,N_9380,N_8757);
and U10978 (N_10978,N_8760,N_8910);
nand U10979 (N_10979,N_8835,N_9559);
nand U10980 (N_10980,N_9160,N_8763);
nand U10981 (N_10981,N_9885,N_9861);
and U10982 (N_10982,N_9922,N_9241);
xor U10983 (N_10983,N_9074,N_9661);
or U10984 (N_10984,N_8805,N_9342);
nor U10985 (N_10985,N_9323,N_9837);
and U10986 (N_10986,N_9743,N_9335);
nand U10987 (N_10987,N_9025,N_8879);
xor U10988 (N_10988,N_8833,N_9144);
nor U10989 (N_10989,N_9864,N_9142);
and U10990 (N_10990,N_9980,N_9884);
xnor U10991 (N_10991,N_8945,N_9544);
nor U10992 (N_10992,N_8866,N_8889);
and U10993 (N_10993,N_8934,N_9926);
or U10994 (N_10994,N_9818,N_9125);
and U10995 (N_10995,N_8893,N_9716);
and U10996 (N_10996,N_8942,N_9492);
xnor U10997 (N_10997,N_9761,N_9529);
nor U10998 (N_10998,N_8907,N_9462);
or U10999 (N_10999,N_9805,N_9245);
nand U11000 (N_11000,N_9907,N_9276);
xor U11001 (N_11001,N_9697,N_9674);
nor U11002 (N_11002,N_9662,N_8808);
nand U11003 (N_11003,N_8965,N_9203);
and U11004 (N_11004,N_9181,N_9718);
xnor U11005 (N_11005,N_9174,N_9581);
or U11006 (N_11006,N_9268,N_9384);
or U11007 (N_11007,N_8998,N_9931);
or U11008 (N_11008,N_9190,N_9065);
nor U11009 (N_11009,N_8995,N_9256);
nand U11010 (N_11010,N_9495,N_9407);
and U11011 (N_11011,N_8845,N_8885);
xor U11012 (N_11012,N_8968,N_9140);
and U11013 (N_11013,N_9214,N_9285);
nand U11014 (N_11014,N_9443,N_9311);
nand U11015 (N_11015,N_9946,N_9125);
xnor U11016 (N_11016,N_9591,N_9293);
nand U11017 (N_11017,N_8802,N_9760);
or U11018 (N_11018,N_9620,N_9483);
and U11019 (N_11019,N_9349,N_9360);
nor U11020 (N_11020,N_9581,N_9371);
or U11021 (N_11021,N_9682,N_8986);
and U11022 (N_11022,N_9881,N_9143);
nand U11023 (N_11023,N_9481,N_9202);
nor U11024 (N_11024,N_8960,N_9538);
or U11025 (N_11025,N_9563,N_9239);
and U11026 (N_11026,N_8937,N_9471);
nand U11027 (N_11027,N_8770,N_9082);
nor U11028 (N_11028,N_9916,N_8949);
xor U11029 (N_11029,N_9611,N_9232);
and U11030 (N_11030,N_8863,N_8903);
or U11031 (N_11031,N_9491,N_9677);
nor U11032 (N_11032,N_9920,N_8970);
or U11033 (N_11033,N_9683,N_9381);
and U11034 (N_11034,N_9984,N_9768);
nand U11035 (N_11035,N_9703,N_9776);
nand U11036 (N_11036,N_8832,N_8952);
xnor U11037 (N_11037,N_9604,N_8829);
xor U11038 (N_11038,N_9864,N_9959);
or U11039 (N_11039,N_9485,N_9067);
xnor U11040 (N_11040,N_8919,N_9642);
nor U11041 (N_11041,N_9905,N_9032);
and U11042 (N_11042,N_9594,N_9277);
or U11043 (N_11043,N_9063,N_9939);
or U11044 (N_11044,N_8791,N_9894);
and U11045 (N_11045,N_9622,N_9755);
or U11046 (N_11046,N_9770,N_9724);
nor U11047 (N_11047,N_9400,N_9384);
and U11048 (N_11048,N_9027,N_8922);
or U11049 (N_11049,N_9261,N_9101);
xor U11050 (N_11050,N_9466,N_9283);
or U11051 (N_11051,N_9543,N_9361);
and U11052 (N_11052,N_9064,N_8852);
and U11053 (N_11053,N_9001,N_9351);
nor U11054 (N_11054,N_9891,N_9474);
or U11055 (N_11055,N_8981,N_9060);
and U11056 (N_11056,N_9549,N_9527);
or U11057 (N_11057,N_9029,N_9489);
xnor U11058 (N_11058,N_9574,N_9606);
or U11059 (N_11059,N_9758,N_9131);
nor U11060 (N_11060,N_9345,N_8872);
nor U11061 (N_11061,N_9058,N_9371);
xnor U11062 (N_11062,N_9015,N_9160);
nand U11063 (N_11063,N_9754,N_9120);
xnor U11064 (N_11064,N_8880,N_8998);
nand U11065 (N_11065,N_9437,N_9709);
nor U11066 (N_11066,N_9543,N_8769);
or U11067 (N_11067,N_9231,N_9085);
and U11068 (N_11068,N_9116,N_8919);
nand U11069 (N_11069,N_8810,N_9449);
xnor U11070 (N_11070,N_9902,N_9429);
or U11071 (N_11071,N_9207,N_9253);
nand U11072 (N_11072,N_9440,N_8838);
nor U11073 (N_11073,N_9817,N_9793);
or U11074 (N_11074,N_9154,N_9098);
xnor U11075 (N_11075,N_9115,N_8764);
nor U11076 (N_11076,N_9954,N_9210);
nor U11077 (N_11077,N_9448,N_9017);
nor U11078 (N_11078,N_9665,N_9510);
and U11079 (N_11079,N_9354,N_8752);
xnor U11080 (N_11080,N_9549,N_9052);
nand U11081 (N_11081,N_9485,N_9747);
nor U11082 (N_11082,N_9486,N_9982);
and U11083 (N_11083,N_9288,N_9627);
xor U11084 (N_11084,N_9246,N_8820);
nand U11085 (N_11085,N_9450,N_8865);
xor U11086 (N_11086,N_9038,N_9966);
and U11087 (N_11087,N_9102,N_9606);
or U11088 (N_11088,N_9484,N_9391);
or U11089 (N_11089,N_9011,N_9834);
xor U11090 (N_11090,N_9739,N_9270);
and U11091 (N_11091,N_8810,N_8890);
nand U11092 (N_11092,N_9600,N_9301);
or U11093 (N_11093,N_8843,N_8828);
xnor U11094 (N_11094,N_9850,N_9782);
or U11095 (N_11095,N_9730,N_9130);
nand U11096 (N_11096,N_9167,N_9485);
and U11097 (N_11097,N_8924,N_9375);
xnor U11098 (N_11098,N_8760,N_9219);
nand U11099 (N_11099,N_9883,N_9809);
nand U11100 (N_11100,N_9199,N_8973);
nor U11101 (N_11101,N_9667,N_9672);
xnor U11102 (N_11102,N_9600,N_9879);
xor U11103 (N_11103,N_9711,N_9126);
xnor U11104 (N_11104,N_9941,N_9153);
nand U11105 (N_11105,N_8763,N_9796);
or U11106 (N_11106,N_9706,N_8901);
xor U11107 (N_11107,N_8978,N_9057);
and U11108 (N_11108,N_8970,N_8949);
and U11109 (N_11109,N_9794,N_9976);
nand U11110 (N_11110,N_8841,N_9606);
or U11111 (N_11111,N_9207,N_9654);
nor U11112 (N_11112,N_9464,N_9612);
nand U11113 (N_11113,N_8868,N_9190);
nand U11114 (N_11114,N_8888,N_9382);
or U11115 (N_11115,N_9882,N_9294);
nor U11116 (N_11116,N_9830,N_8912);
xnor U11117 (N_11117,N_9955,N_9951);
nand U11118 (N_11118,N_8758,N_9979);
and U11119 (N_11119,N_9870,N_9124);
and U11120 (N_11120,N_9129,N_9394);
or U11121 (N_11121,N_8816,N_9037);
xor U11122 (N_11122,N_8926,N_9653);
nand U11123 (N_11123,N_9757,N_9973);
nor U11124 (N_11124,N_9106,N_9663);
or U11125 (N_11125,N_9461,N_8891);
nand U11126 (N_11126,N_8892,N_9283);
nor U11127 (N_11127,N_8824,N_8863);
or U11128 (N_11128,N_9849,N_9550);
xor U11129 (N_11129,N_9477,N_9114);
xnor U11130 (N_11130,N_9799,N_9097);
nor U11131 (N_11131,N_9458,N_9648);
nor U11132 (N_11132,N_9654,N_9753);
nor U11133 (N_11133,N_8801,N_9096);
xnor U11134 (N_11134,N_9775,N_8764);
or U11135 (N_11135,N_9582,N_9020);
and U11136 (N_11136,N_9919,N_9515);
nand U11137 (N_11137,N_9027,N_9944);
or U11138 (N_11138,N_9171,N_9262);
or U11139 (N_11139,N_8788,N_8963);
xor U11140 (N_11140,N_9018,N_9146);
nand U11141 (N_11141,N_9111,N_9212);
nand U11142 (N_11142,N_9440,N_8912);
nor U11143 (N_11143,N_9801,N_9989);
nand U11144 (N_11144,N_8917,N_9046);
or U11145 (N_11145,N_9383,N_9795);
and U11146 (N_11146,N_9327,N_9910);
nor U11147 (N_11147,N_8852,N_8961);
nor U11148 (N_11148,N_9295,N_9047);
xnor U11149 (N_11149,N_9660,N_9582);
xnor U11150 (N_11150,N_9883,N_9244);
nand U11151 (N_11151,N_9581,N_9463);
or U11152 (N_11152,N_9115,N_8978);
nor U11153 (N_11153,N_8968,N_9317);
nor U11154 (N_11154,N_9178,N_9614);
nor U11155 (N_11155,N_9980,N_9558);
nor U11156 (N_11156,N_9800,N_9914);
nand U11157 (N_11157,N_9773,N_9459);
nor U11158 (N_11158,N_9062,N_9059);
xnor U11159 (N_11159,N_9142,N_8999);
or U11160 (N_11160,N_8988,N_9731);
nand U11161 (N_11161,N_8875,N_9809);
or U11162 (N_11162,N_9542,N_9508);
or U11163 (N_11163,N_9724,N_9409);
nor U11164 (N_11164,N_8765,N_9040);
or U11165 (N_11165,N_9359,N_9041);
nor U11166 (N_11166,N_8950,N_8970);
and U11167 (N_11167,N_8784,N_8944);
xnor U11168 (N_11168,N_9111,N_9659);
xor U11169 (N_11169,N_8791,N_8966);
nand U11170 (N_11170,N_9533,N_9483);
and U11171 (N_11171,N_9823,N_8914);
nor U11172 (N_11172,N_8895,N_8974);
nand U11173 (N_11173,N_9551,N_9011);
xnor U11174 (N_11174,N_9395,N_9538);
or U11175 (N_11175,N_9243,N_9464);
xor U11176 (N_11176,N_9674,N_8910);
xor U11177 (N_11177,N_9770,N_9267);
or U11178 (N_11178,N_9641,N_8959);
and U11179 (N_11179,N_8908,N_8959);
nor U11180 (N_11180,N_9842,N_9228);
xor U11181 (N_11181,N_9296,N_9778);
nand U11182 (N_11182,N_9005,N_9900);
and U11183 (N_11183,N_9611,N_9370);
nor U11184 (N_11184,N_8976,N_9267);
and U11185 (N_11185,N_9916,N_8791);
or U11186 (N_11186,N_8830,N_9137);
xnor U11187 (N_11187,N_9441,N_9835);
nand U11188 (N_11188,N_9970,N_9878);
xnor U11189 (N_11189,N_9275,N_9933);
or U11190 (N_11190,N_8998,N_8950);
and U11191 (N_11191,N_9243,N_9016);
xor U11192 (N_11192,N_9217,N_8858);
nand U11193 (N_11193,N_9958,N_9782);
nor U11194 (N_11194,N_9623,N_9681);
and U11195 (N_11195,N_9209,N_9148);
and U11196 (N_11196,N_9447,N_8788);
nand U11197 (N_11197,N_9106,N_9979);
or U11198 (N_11198,N_9399,N_9463);
xor U11199 (N_11199,N_9222,N_9563);
or U11200 (N_11200,N_8837,N_9279);
xnor U11201 (N_11201,N_8934,N_9250);
xnor U11202 (N_11202,N_8947,N_8934);
xor U11203 (N_11203,N_9148,N_9992);
and U11204 (N_11204,N_8921,N_9019);
or U11205 (N_11205,N_9665,N_9082);
nor U11206 (N_11206,N_9080,N_8758);
xnor U11207 (N_11207,N_9317,N_9436);
nor U11208 (N_11208,N_9198,N_9313);
xnor U11209 (N_11209,N_8919,N_8815);
nand U11210 (N_11210,N_9798,N_8998);
or U11211 (N_11211,N_9475,N_9190);
xnor U11212 (N_11212,N_9708,N_8957);
and U11213 (N_11213,N_8971,N_9966);
and U11214 (N_11214,N_9205,N_9309);
nand U11215 (N_11215,N_9080,N_9986);
nand U11216 (N_11216,N_9930,N_9347);
xnor U11217 (N_11217,N_8803,N_9650);
and U11218 (N_11218,N_9012,N_9534);
or U11219 (N_11219,N_9337,N_9645);
and U11220 (N_11220,N_9569,N_9736);
and U11221 (N_11221,N_9951,N_9813);
xor U11222 (N_11222,N_9472,N_9567);
nor U11223 (N_11223,N_9420,N_9561);
nor U11224 (N_11224,N_9862,N_9751);
or U11225 (N_11225,N_8820,N_8947);
or U11226 (N_11226,N_9791,N_9873);
nor U11227 (N_11227,N_9738,N_9268);
or U11228 (N_11228,N_9105,N_9699);
and U11229 (N_11229,N_9988,N_8907);
or U11230 (N_11230,N_9340,N_9711);
nand U11231 (N_11231,N_8824,N_9323);
and U11232 (N_11232,N_9662,N_9922);
nand U11233 (N_11233,N_9586,N_9390);
or U11234 (N_11234,N_9629,N_9586);
nand U11235 (N_11235,N_9546,N_9585);
and U11236 (N_11236,N_9781,N_9376);
nand U11237 (N_11237,N_9973,N_8923);
nand U11238 (N_11238,N_9022,N_9033);
xor U11239 (N_11239,N_9530,N_9985);
nand U11240 (N_11240,N_9866,N_8816);
and U11241 (N_11241,N_9004,N_9536);
or U11242 (N_11242,N_9268,N_9953);
or U11243 (N_11243,N_9724,N_9218);
or U11244 (N_11244,N_8838,N_9988);
xor U11245 (N_11245,N_9121,N_9515);
xnor U11246 (N_11246,N_9396,N_8901);
nor U11247 (N_11247,N_9568,N_9083);
xor U11248 (N_11248,N_9263,N_9180);
nand U11249 (N_11249,N_9518,N_9212);
nand U11250 (N_11250,N_10197,N_10455);
or U11251 (N_11251,N_10771,N_10140);
and U11252 (N_11252,N_10638,N_10391);
and U11253 (N_11253,N_11223,N_10476);
xnor U11254 (N_11254,N_10873,N_10867);
or U11255 (N_11255,N_11085,N_11058);
xor U11256 (N_11256,N_10023,N_10827);
nor U11257 (N_11257,N_11070,N_10424);
and U11258 (N_11258,N_11066,N_10637);
nor U11259 (N_11259,N_11052,N_10312);
xor U11260 (N_11260,N_10046,N_11235);
xnor U11261 (N_11261,N_10387,N_10869);
nand U11262 (N_11262,N_10672,N_10372);
or U11263 (N_11263,N_10982,N_10325);
nor U11264 (N_11264,N_10803,N_10788);
nor U11265 (N_11265,N_11083,N_10795);
and U11266 (N_11266,N_11116,N_10336);
or U11267 (N_11267,N_10112,N_10700);
and U11268 (N_11268,N_10826,N_10430);
nand U11269 (N_11269,N_10497,N_11055);
xor U11270 (N_11270,N_10825,N_11148);
or U11271 (N_11271,N_10540,N_10519);
or U11272 (N_11272,N_11050,N_10089);
nor U11273 (N_11273,N_10020,N_10151);
or U11274 (N_11274,N_10723,N_10792);
or U11275 (N_11275,N_11152,N_10470);
and U11276 (N_11276,N_11018,N_10431);
and U11277 (N_11277,N_10742,N_10362);
nor U11278 (N_11278,N_10775,N_11047);
xnor U11279 (N_11279,N_11138,N_10852);
nor U11280 (N_11280,N_11035,N_10373);
and U11281 (N_11281,N_10656,N_10056);
nor U11282 (N_11282,N_10279,N_10328);
or U11283 (N_11283,N_10643,N_10975);
nand U11284 (N_11284,N_10908,N_10642);
and U11285 (N_11285,N_11079,N_11180);
or U11286 (N_11286,N_10257,N_10349);
or U11287 (N_11287,N_10084,N_10466);
nand U11288 (N_11288,N_10443,N_10760);
and U11289 (N_11289,N_10664,N_10233);
xor U11290 (N_11290,N_11068,N_10215);
nand U11291 (N_11291,N_10575,N_10761);
nor U11292 (N_11292,N_10845,N_10011);
or U11293 (N_11293,N_10940,N_10207);
and U11294 (N_11294,N_11040,N_10914);
and U11295 (N_11295,N_11041,N_11209);
or U11296 (N_11296,N_10160,N_11100);
or U11297 (N_11297,N_10369,N_10976);
nor U11298 (N_11298,N_11030,N_10404);
nor U11299 (N_11299,N_10150,N_10678);
and U11300 (N_11300,N_10662,N_10807);
nor U11301 (N_11301,N_10117,N_10813);
and U11302 (N_11302,N_11219,N_10456);
xor U11303 (N_11303,N_10350,N_10554);
nand U11304 (N_11304,N_10818,N_10446);
nor U11305 (N_11305,N_10270,N_10861);
xnor U11306 (N_11306,N_10066,N_10314);
or U11307 (N_11307,N_11043,N_10205);
and U11308 (N_11308,N_11194,N_11122);
nor U11309 (N_11309,N_10783,N_10756);
or U11310 (N_11310,N_10037,N_10832);
nand U11311 (N_11311,N_10582,N_10725);
and U11312 (N_11312,N_10418,N_10543);
xor U11313 (N_11313,N_10405,N_10768);
and U11314 (N_11314,N_10401,N_10359);
nand U11315 (N_11315,N_10413,N_10434);
or U11316 (N_11316,N_10625,N_10087);
and U11317 (N_11317,N_10167,N_11182);
or U11318 (N_11318,N_10367,N_10896);
xor U11319 (N_11319,N_10200,N_10267);
or U11320 (N_11320,N_10786,N_10196);
nand U11321 (N_11321,N_10144,N_11073);
and U11322 (N_11322,N_10016,N_10866);
nand U11323 (N_11323,N_10142,N_10546);
and U11324 (N_11324,N_10291,N_10879);
nor U11325 (N_11325,N_11239,N_10882);
or U11326 (N_11326,N_10102,N_10495);
nand U11327 (N_11327,N_10079,N_10222);
or U11328 (N_11328,N_10149,N_10365);
nand U11329 (N_11329,N_10006,N_10030);
nor U11330 (N_11330,N_10473,N_10623);
nor U11331 (N_11331,N_10624,N_10242);
or U11332 (N_11332,N_10542,N_11137);
nand U11333 (N_11333,N_10422,N_10416);
and U11334 (N_11334,N_10534,N_10272);
or U11335 (N_11335,N_10920,N_11130);
and U11336 (N_11336,N_10281,N_10979);
and U11337 (N_11337,N_10703,N_10880);
and U11338 (N_11338,N_10206,N_10518);
nand U11339 (N_11339,N_10123,N_10973);
nand U11340 (N_11340,N_10000,N_10798);
xor U11341 (N_11341,N_11129,N_10351);
xnor U11342 (N_11342,N_11039,N_10185);
nand U11343 (N_11343,N_10647,N_10857);
nand U11344 (N_11344,N_10286,N_10346);
and U11345 (N_11345,N_10584,N_10115);
nor U11346 (N_11346,N_11192,N_10411);
and U11347 (N_11347,N_10989,N_10716);
or U11348 (N_11348,N_11088,N_10746);
and U11349 (N_11349,N_10284,N_11104);
and U11350 (N_11350,N_10382,N_10025);
or U11351 (N_11351,N_11119,N_10441);
xor U11352 (N_11352,N_10461,N_11190);
xor U11353 (N_11353,N_10467,N_11141);
or U11354 (N_11354,N_10577,N_10711);
and U11355 (N_11355,N_10212,N_11062);
xnor U11356 (N_11356,N_11011,N_10189);
xor U11357 (N_11357,N_10528,N_11218);
nand U11358 (N_11358,N_10428,N_10892);
nor U11359 (N_11359,N_10371,N_10343);
and U11360 (N_11360,N_10060,N_11044);
nand U11361 (N_11361,N_10042,N_10425);
or U11362 (N_11362,N_10487,N_10671);
nand U11363 (N_11363,N_10930,N_11005);
and U11364 (N_11364,N_10226,N_11236);
or U11365 (N_11365,N_11102,N_10688);
nand U11366 (N_11366,N_10157,N_10330);
or U11367 (N_11367,N_11206,N_10676);
nor U11368 (N_11368,N_10429,N_10731);
nor U11369 (N_11369,N_10782,N_10718);
nand U11370 (N_11370,N_10258,N_10213);
nor U11371 (N_11371,N_10120,N_11121);
and U11372 (N_11372,N_10093,N_11217);
xnor U11373 (N_11373,N_11074,N_10396);
or U11374 (N_11374,N_10061,N_10100);
or U11375 (N_11375,N_10250,N_10047);
and U11376 (N_11376,N_10837,N_11228);
nand U11377 (N_11377,N_10680,N_11000);
and U11378 (N_11378,N_10763,N_10415);
and U11379 (N_11379,N_10708,N_10663);
xnor U11380 (N_11380,N_10944,N_10444);
nand U11381 (N_11381,N_11127,N_10294);
nand U11382 (N_11382,N_10249,N_10646);
xor U11383 (N_11383,N_11037,N_10915);
nand U11384 (N_11384,N_10210,N_10550);
nor U11385 (N_11385,N_10885,N_10955);
or U11386 (N_11386,N_10757,N_10732);
or U11387 (N_11387,N_10370,N_10218);
nand U11388 (N_11388,N_10306,N_10539);
and U11389 (N_11389,N_11154,N_10627);
nor U11390 (N_11390,N_10881,N_11015);
xor U11391 (N_11391,N_11150,N_10124);
or U11392 (N_11392,N_10427,N_11230);
or U11393 (N_11393,N_10937,N_10406);
nand U11394 (N_11394,N_10521,N_10936);
and U11395 (N_11395,N_10152,N_10987);
and U11396 (N_11396,N_10345,N_10400);
and U11397 (N_11397,N_10465,N_10402);
nand U11398 (N_11398,N_10409,N_10054);
and U11399 (N_11399,N_10863,N_10981);
nand U11400 (N_11400,N_10407,N_11179);
nand U11401 (N_11401,N_10479,N_10116);
and U11402 (N_11402,N_10065,N_10527);
nor U11403 (N_11403,N_10278,N_10552);
nand U11404 (N_11404,N_11022,N_10126);
xor U11405 (N_11405,N_11132,N_11143);
or U11406 (N_11406,N_10209,N_10356);
xor U11407 (N_11407,N_10828,N_11155);
and U11408 (N_11408,N_10526,N_10878);
or U11409 (N_11409,N_10195,N_10352);
and U11410 (N_11410,N_10015,N_10594);
and U11411 (N_11411,N_10490,N_10165);
and U11412 (N_11412,N_10462,N_10502);
and U11413 (N_11413,N_10044,N_10839);
nand U11414 (N_11414,N_11167,N_10288);
or U11415 (N_11415,N_10724,N_10463);
xor U11416 (N_11416,N_10472,N_10793);
and U11417 (N_11417,N_10492,N_11238);
or U11418 (N_11418,N_10018,N_11227);
and U11419 (N_11419,N_10500,N_10655);
nor U11420 (N_11420,N_10318,N_10347);
nand U11421 (N_11421,N_10277,N_10645);
nor U11422 (N_11422,N_11161,N_10097);
nor U11423 (N_11423,N_10603,N_10652);
xor U11424 (N_11424,N_10177,N_10968);
nor U11425 (N_11425,N_11204,N_11147);
or U11426 (N_11426,N_10386,N_11229);
xnor U11427 (N_11427,N_10403,N_10965);
and U11428 (N_11428,N_11195,N_10947);
nor U11429 (N_11429,N_10377,N_10484);
xnor U11430 (N_11430,N_10460,N_10376);
xor U11431 (N_11431,N_10039,N_10769);
nand U11432 (N_11432,N_10851,N_10933);
and U11433 (N_11433,N_11196,N_10544);
or U11434 (N_11434,N_10988,N_10368);
nor U11435 (N_11435,N_10059,N_10545);
nand U11436 (N_11436,N_10145,N_10287);
xnor U11437 (N_11437,N_10875,N_10579);
nand U11438 (N_11438,N_10477,N_10034);
or U11439 (N_11439,N_10560,N_10265);
xor U11440 (N_11440,N_10113,N_10324);
nand U11441 (N_11441,N_10299,N_10618);
xnor U11442 (N_11442,N_10119,N_10191);
nor U11443 (N_11443,N_10040,N_10259);
xor U11444 (N_11444,N_11106,N_10701);
or U11445 (N_11445,N_11065,N_10748);
xor U11446 (N_11446,N_10801,N_10785);
xnor U11447 (N_11447,N_10800,N_10109);
and U11448 (N_11448,N_10053,N_10051);
nor U11449 (N_11449,N_10578,N_10549);
or U11450 (N_11450,N_10841,N_11115);
nand U11451 (N_11451,N_10513,N_11176);
nor U11452 (N_11452,N_10906,N_10326);
nor U11453 (N_11453,N_10078,N_10735);
xnor U11454 (N_11454,N_11247,N_10816);
or U11455 (N_11455,N_10009,N_11232);
nand U11456 (N_11456,N_10354,N_10361);
nor U11457 (N_11457,N_10894,N_10874);
xor U11458 (N_11458,N_10379,N_10236);
nand U11459 (N_11459,N_10335,N_11123);
nor U11460 (N_11460,N_10911,N_11157);
and U11461 (N_11461,N_10969,N_10834);
nor U11462 (N_11462,N_11200,N_10316);
nand U11463 (N_11463,N_10804,N_10055);
or U11464 (N_11464,N_11225,N_10986);
nand U11465 (N_11465,N_10069,N_10175);
xnor U11466 (N_11466,N_10938,N_10694);
and U11467 (N_11467,N_10687,N_10075);
nor U11468 (N_11468,N_11089,N_10166);
or U11469 (N_11469,N_10616,N_10548);
or U11470 (N_11470,N_10946,N_10311);
xnor U11471 (N_11471,N_10012,N_10659);
xor U11472 (N_11472,N_10934,N_10074);
nand U11473 (N_11473,N_10491,N_11101);
xnor U11474 (N_11474,N_10840,N_11210);
and U11475 (N_11475,N_10104,N_10217);
nand U11476 (N_11476,N_10147,N_10192);
nand U11477 (N_11477,N_11215,N_10143);
nor U11478 (N_11478,N_10706,N_10085);
or U11479 (N_11479,N_10949,N_10593);
nor U11480 (N_11480,N_10108,N_10499);
or U11481 (N_11481,N_10759,N_10360);
and U11482 (N_11482,N_10685,N_10410);
and U11483 (N_11483,N_10977,N_10689);
nor U11484 (N_11484,N_10208,N_10329);
or U11485 (N_11485,N_10300,N_10953);
xor U11486 (N_11486,N_10910,N_10547);
and U11487 (N_11487,N_11126,N_11243);
and U11488 (N_11488,N_10905,N_10622);
and U11489 (N_11489,N_10590,N_10961);
xor U11490 (N_11490,N_10134,N_10653);
nand U11491 (N_11491,N_10219,N_10891);
nand U11492 (N_11492,N_10683,N_10812);
nor U11493 (N_11493,N_11033,N_10408);
and U11494 (N_11494,N_10595,N_10179);
xor U11495 (N_11495,N_10833,N_10509);
nand U11496 (N_11496,N_10062,N_10644);
nand U11497 (N_11497,N_10453,N_10844);
and U11498 (N_11498,N_10613,N_10669);
nand U11499 (N_11499,N_10707,N_10159);
and U11500 (N_11500,N_11029,N_10088);
or U11501 (N_11501,N_10187,N_10781);
or U11502 (N_11502,N_10586,N_11197);
and U11503 (N_11503,N_10810,N_10263);
nor U11504 (N_11504,N_11249,N_10138);
xor U11505 (N_11505,N_10570,N_10141);
xor U11506 (N_11506,N_10310,N_10426);
nand U11507 (N_11507,N_10262,N_10237);
nor U11508 (N_11508,N_10156,N_10903);
and U11509 (N_11509,N_10146,N_10870);
nand U11510 (N_11510,N_10727,N_11097);
nor U11511 (N_11511,N_10665,N_10508);
and U11512 (N_11512,N_10736,N_11128);
and U11513 (N_11513,N_10581,N_11096);
or U11514 (N_11514,N_11164,N_10872);
nand U11515 (N_11515,N_10675,N_10071);
and U11516 (N_11516,N_10639,N_10601);
and U11517 (N_11517,N_10805,N_10449);
or U11518 (N_11518,N_11221,N_10384);
nor U11519 (N_11519,N_10538,N_11173);
and U11520 (N_11520,N_10271,N_10564);
xor U11521 (N_11521,N_10983,N_10353);
and U11522 (N_11522,N_11046,N_10510);
or U11523 (N_11523,N_10496,N_10216);
nor U11524 (N_11524,N_10533,N_10650);
nand U11525 (N_11525,N_10133,N_10691);
xnor U11526 (N_11526,N_10433,N_10073);
nor U11527 (N_11527,N_10445,N_10820);
xor U11528 (N_11528,N_11174,N_10302);
and U11529 (N_11529,N_11160,N_11142);
xor U11530 (N_11530,N_10252,N_10733);
nor U11531 (N_11531,N_10559,N_10342);
nor U11532 (N_11532,N_10293,N_11056);
nor U11533 (N_11533,N_11027,N_10997);
and U11534 (N_11534,N_10773,N_10996);
xor U11535 (N_11535,N_11118,N_10323);
xor U11536 (N_11536,N_10823,N_10264);
and U11537 (N_11537,N_10378,N_10715);
and U11538 (N_11538,N_10799,N_10806);
or U11539 (N_11539,N_10363,N_10244);
xor U11540 (N_11540,N_10161,N_10587);
xor U11541 (N_11541,N_10557,N_11092);
and U11542 (N_11542,N_10722,N_10174);
xor U11543 (N_11543,N_10471,N_11188);
xnor U11544 (N_11544,N_10838,N_11017);
and U11545 (N_11545,N_10202,N_10941);
nor U11546 (N_11546,N_10537,N_10829);
nand U11547 (N_11547,N_10058,N_10958);
and U11548 (N_11548,N_10154,N_10963);
or U11549 (N_11549,N_11183,N_10095);
or U11550 (N_11550,N_10610,N_11023);
nor U11551 (N_11551,N_10475,N_10974);
and U11552 (N_11552,N_10243,N_10999);
nand U11553 (N_11553,N_10091,N_11178);
and U11554 (N_11554,N_10331,N_11059);
xnor U11555 (N_11555,N_11103,N_11048);
or U11556 (N_11556,N_10729,N_10511);
nor U11557 (N_11557,N_10515,N_10713);
and U11558 (N_11558,N_10897,N_10574);
and U11559 (N_11559,N_10454,N_11034);
xnor U11560 (N_11560,N_10290,N_10884);
xor U11561 (N_11561,N_10229,N_10067);
nor U11562 (N_11562,N_10366,N_10380);
xnor U11563 (N_11563,N_10423,N_10507);
xor U11564 (N_11564,N_11007,N_10395);
nor U11565 (N_11565,N_10320,N_10419);
xnor U11566 (N_11566,N_11110,N_10033);
or U11567 (N_11567,N_10480,N_10474);
nor U11568 (N_11568,N_10121,N_11010);
xnor U11569 (N_11569,N_11111,N_10576);
and U11570 (N_11570,N_11242,N_10321);
xor U11571 (N_11571,N_10524,N_10494);
nand U11572 (N_11572,N_11199,N_10925);
xor U11573 (N_11573,N_10190,N_10269);
nand U11574 (N_11574,N_10796,N_10155);
nand U11575 (N_11575,N_10929,N_10114);
nor U11576 (N_11576,N_10960,N_10850);
nand U11577 (N_11577,N_11246,N_10596);
nor U11578 (N_11578,N_10348,N_11061);
and U11579 (N_11579,N_10649,N_10978);
nand U11580 (N_11580,N_10274,N_10889);
xnor U11581 (N_11581,N_11078,N_10019);
nand U11582 (N_11582,N_10846,N_10504);
and U11583 (N_11583,N_10754,N_10493);
xnor U11584 (N_11584,N_11248,N_10615);
or U11585 (N_11585,N_10864,N_11014);
nor U11586 (N_11586,N_10086,N_10198);
nor U11587 (N_11587,N_10035,N_10036);
or U11588 (N_11588,N_10612,N_10765);
xnor U11589 (N_11589,N_10442,N_10122);
and U11590 (N_11590,N_10566,N_10822);
and U11591 (N_11591,N_10952,N_10082);
nand U11592 (N_11592,N_11021,N_10355);
xor U11593 (N_11593,N_10333,N_10478);
nor U11594 (N_11594,N_10661,N_10303);
nand U11595 (N_11595,N_10762,N_10186);
or U11596 (N_11596,N_10043,N_10853);
and U11597 (N_11597,N_10717,N_11231);
xnor U11598 (N_11598,N_10483,N_10758);
or U11599 (N_11599,N_10398,N_10931);
nand U11600 (N_11600,N_10130,N_10668);
nand U11601 (N_11601,N_10922,N_11186);
xor U11602 (N_11602,N_10942,N_10090);
or U11603 (N_11603,N_11203,N_10740);
or U11604 (N_11604,N_10261,N_10770);
or U11605 (N_11605,N_11158,N_11208);
and U11606 (N_11606,N_10247,N_11016);
nor U11607 (N_11607,N_10614,N_11189);
nor U11608 (N_11608,N_10606,N_10092);
or U11609 (N_11609,N_10859,N_10211);
and U11610 (N_11610,N_10730,N_10332);
and U11611 (N_11611,N_10592,N_10726);
nor U11612 (N_11612,N_10127,N_10458);
nor U11613 (N_11613,N_10636,N_10240);
and U11614 (N_11614,N_10912,N_10923);
xnor U11615 (N_11615,N_11053,N_10710);
xor U11616 (N_11616,N_11108,N_10917);
xor U11617 (N_11617,N_10181,N_10657);
xnor U11618 (N_11618,N_10180,N_10744);
nand U11619 (N_11619,N_10970,N_11026);
or U11620 (N_11620,N_10038,N_10565);
xor U11621 (N_11621,N_10990,N_10790);
nor U11622 (N_11622,N_10898,N_10225);
xnor U11623 (N_11623,N_10251,N_11187);
nor U11624 (N_11624,N_10635,N_10531);
xnor U11625 (N_11625,N_10420,N_10862);
and U11626 (N_11626,N_10702,N_10985);
and U11627 (N_11627,N_11166,N_10464);
or U11628 (N_11628,N_10232,N_10860);
xnor U11629 (N_11629,N_10337,N_10005);
xnor U11630 (N_11630,N_10132,N_10682);
or U11631 (N_11631,N_10517,N_11184);
nor U11632 (N_11632,N_10695,N_10690);
and U11633 (N_11633,N_10532,N_10600);
and U11634 (N_11634,N_10414,N_11002);
nand U11635 (N_11635,N_10802,N_11072);
or U11636 (N_11636,N_10608,N_10536);
nand U11637 (N_11637,N_10501,N_10957);
nor U11638 (N_11638,N_10573,N_10224);
and U11639 (N_11639,N_10001,N_10516);
nand U11640 (N_11640,N_10745,N_10070);
xor U11641 (N_11641,N_11012,N_11172);
or U11642 (N_11642,N_10569,N_10309);
and U11643 (N_11643,N_10842,N_10909);
nand U11644 (N_11644,N_10003,N_10815);
or U11645 (N_11645,N_10172,N_10966);
xor U11646 (N_11646,N_10292,N_10266);
xnor U11647 (N_11647,N_10855,N_11006);
and U11648 (N_11648,N_10541,N_10628);
or U11649 (N_11649,N_10289,N_10535);
xor U11650 (N_11650,N_10971,N_11087);
xnor U11651 (N_11651,N_10170,N_10887);
nand U11652 (N_11652,N_10945,N_10883);
nand U11653 (N_11653,N_11090,N_10588);
nor U11654 (N_11654,N_10305,N_10072);
nor U11655 (N_11655,N_10617,N_10720);
xnor U11656 (N_11656,N_11114,N_10836);
or U11657 (N_11657,N_10630,N_10993);
and U11658 (N_11658,N_10273,N_11008);
nand U11659 (N_11659,N_10118,N_10948);
nand U11660 (N_11660,N_10027,N_10438);
and U11661 (N_11661,N_10105,N_10245);
nand U11662 (N_11662,N_10469,N_10021);
nand U11663 (N_11663,N_11060,N_10776);
or U11664 (N_11664,N_10611,N_10136);
or U11665 (N_11665,N_10699,N_10609);
nand U11666 (N_11666,N_10194,N_10918);
nor U11667 (N_11667,N_10779,N_10107);
nand U11668 (N_11668,N_10819,N_10101);
nand U11669 (N_11669,N_10629,N_10686);
and U11670 (N_11670,N_11177,N_10809);
or U11671 (N_11671,N_10913,N_10421);
and U11672 (N_11672,N_10709,N_10784);
nand U11673 (N_11673,N_10276,N_10563);
and U11674 (N_11674,N_10241,N_11125);
xnor U11675 (N_11675,N_10670,N_10417);
nor U11676 (N_11676,N_11024,N_10489);
nand U11677 (N_11677,N_10254,N_11082);
and U11678 (N_11678,N_11095,N_10026);
or U11679 (N_11679,N_10094,N_10052);
nand U11680 (N_11680,N_10512,N_11241);
or U11681 (N_11681,N_10280,N_10392);
nor U11682 (N_11682,N_10028,N_10201);
nor U11683 (N_11683,N_10641,N_10571);
and U11684 (N_11684,N_10858,N_10951);
and U11685 (N_11685,N_10103,N_10468);
nor U11686 (N_11686,N_11112,N_10283);
nor U11687 (N_11687,N_10602,N_10317);
xor U11688 (N_11688,N_10375,N_10835);
nor U11689 (N_11689,N_10959,N_10199);
and U11690 (N_11690,N_10849,N_10660);
and U11691 (N_11691,N_10814,N_10824);
xor U11692 (N_11692,N_11144,N_11028);
and U11693 (N_11693,N_10048,N_10248);
and U11694 (N_11694,N_10432,N_11193);
nor U11695 (N_11695,N_10004,N_10296);
nor U11696 (N_11696,N_10871,N_10246);
or U11697 (N_11697,N_10750,N_10227);
nor U11698 (N_11698,N_11057,N_10556);
and U11699 (N_11699,N_10943,N_10488);
nand U11700 (N_11700,N_11067,N_10697);
nor U11701 (N_11701,N_10457,N_11216);
nor U11702 (N_11702,N_10435,N_10153);
and U11703 (N_11703,N_10604,N_10865);
nand U11704 (N_11704,N_10080,N_10388);
nor U11705 (N_11705,N_10385,N_10188);
and U11706 (N_11706,N_11075,N_10752);
nand U11707 (N_11707,N_10921,N_10394);
nand U11708 (N_11708,N_10572,N_10598);
nor U11709 (N_11709,N_10684,N_10916);
nor U11710 (N_11710,N_10412,N_10967);
nor U11711 (N_11711,N_10131,N_10451);
and U11712 (N_11712,N_11051,N_10525);
or U11713 (N_11713,N_10791,N_10529);
nor U11714 (N_11714,N_10505,N_10591);
xor U11715 (N_11715,N_11245,N_11113);
or U11716 (N_11716,N_10739,N_10995);
nand U11717 (N_11717,N_10285,N_11201);
and U11718 (N_11718,N_10313,N_10924);
xor U11719 (N_11719,N_11181,N_10128);
or U11720 (N_11720,N_10939,N_10341);
nand U11721 (N_11721,N_11224,N_10327);
or U11722 (N_11722,N_10282,N_10705);
nor U11723 (N_11723,N_10322,N_10777);
or U11724 (N_11724,N_10597,N_10163);
nor U11725 (N_11725,N_10766,N_10704);
nor U11726 (N_11726,N_10340,N_10962);
xnor U11727 (N_11727,N_10077,N_10902);
nor U11728 (N_11728,N_11149,N_11038);
nor U11729 (N_11729,N_10255,N_10741);
nand U11730 (N_11730,N_10868,N_11153);
xnor U11731 (N_11731,N_10928,N_10831);
nand U11732 (N_11732,N_10171,N_11212);
xnor U11733 (N_11733,N_11198,N_11222);
nor U11734 (N_11734,N_11207,N_10260);
and U11735 (N_11735,N_10935,N_10383);
or U11736 (N_11736,N_10439,N_11107);
xor U11737 (N_11737,N_11049,N_10334);
nor U11738 (N_11738,N_10568,N_10319);
or U11739 (N_11739,N_10008,N_10964);
and U11740 (N_11740,N_10397,N_10956);
nor U11741 (N_11741,N_11244,N_10607);
xor U11742 (N_11742,N_10137,N_10393);
or U11743 (N_11743,N_11213,N_10485);
xor U11744 (N_11744,N_10658,N_10677);
xor U11745 (N_11745,N_10558,N_10692);
nand U11746 (N_11746,N_11159,N_10106);
or U11747 (N_11747,N_10256,N_10486);
nor U11748 (N_11748,N_10932,N_10482);
nor U11749 (N_11749,N_10821,N_10498);
or U11750 (N_11750,N_11025,N_10437);
nor U11751 (N_11751,N_11001,N_10778);
and U11752 (N_11752,N_10843,N_11131);
or U11753 (N_11753,N_10076,N_10553);
nor U11754 (N_11754,N_11205,N_10307);
nor U11755 (N_11755,N_10679,N_10751);
and U11756 (N_11756,N_10998,N_11091);
or U11757 (N_11757,N_10737,N_11009);
and U11758 (N_11758,N_10111,N_10221);
nand U11759 (N_11759,N_10002,N_10007);
xnor U11760 (N_11760,N_10808,N_10774);
nand U11761 (N_11761,N_10619,N_11226);
nand U11762 (N_11762,N_11165,N_10041);
and U11763 (N_11763,N_10551,N_10714);
nand U11764 (N_11764,N_10447,N_10139);
or U11765 (N_11765,N_10031,N_11081);
or U11766 (N_11766,N_10797,N_10178);
or U11767 (N_11767,N_10193,N_10888);
or U11768 (N_11768,N_10235,N_10721);
and U11769 (N_11769,N_10904,N_10626);
xor U11770 (N_11770,N_10900,N_10919);
or U11771 (N_11771,N_10927,N_11042);
and U11772 (N_11772,N_10696,N_10049);
nand U11773 (N_11773,N_10013,N_11175);
nand U11774 (N_11774,N_10135,N_10148);
nand U11775 (N_11775,N_10893,N_10176);
xor U11776 (N_11776,N_10632,N_10877);
nand U11777 (N_11777,N_10164,N_10068);
or U11778 (N_11778,N_11054,N_10204);
and U11779 (N_11779,N_10389,N_10017);
nor U11780 (N_11780,N_10064,N_10399);
xnor U11781 (N_11781,N_11098,N_10358);
or U11782 (N_11782,N_10681,N_10901);
or U11783 (N_11783,N_10275,N_10010);
nor U11784 (N_11784,N_10481,N_10580);
nand U11785 (N_11785,N_10780,N_10344);
or U11786 (N_11786,N_11086,N_10755);
and U11787 (N_11787,N_11168,N_10029);
nor U11788 (N_11788,N_11076,N_11036);
or U11789 (N_11789,N_10228,N_10633);
or U11790 (N_11790,N_10583,N_11080);
nor U11791 (N_11791,N_10253,N_10847);
xnor U11792 (N_11792,N_10712,N_10338);
xnor U11793 (N_11793,N_10315,N_11135);
xor U11794 (N_11794,N_10728,N_10238);
xor U11795 (N_11795,N_10907,N_11214);
or U11796 (N_11796,N_10698,N_10522);
nand U11797 (N_11797,N_11099,N_11170);
or U11798 (N_11798,N_10753,N_10050);
and U11799 (N_11799,N_11140,N_10561);
xor U11800 (N_11800,N_10014,N_11019);
nand U11801 (N_11801,N_10749,N_11063);
nand U11802 (N_11802,N_10585,N_10605);
or U11803 (N_11803,N_10848,N_10231);
nor U11804 (N_11804,N_10984,N_10738);
xnor U11805 (N_11805,N_10886,N_10440);
nor U11806 (N_11806,N_11136,N_10991);
or U11807 (N_11807,N_10162,N_10057);
nor U11808 (N_11808,N_10032,N_11093);
nand U11809 (N_11809,N_10589,N_10390);
nand U11810 (N_11810,N_11003,N_10298);
or U11811 (N_11811,N_11077,N_10743);
xnor U11812 (N_11812,N_10096,N_10523);
nor U11813 (N_11813,N_11071,N_10436);
nor U11814 (N_11814,N_10158,N_10450);
nor U11815 (N_11815,N_11162,N_11020);
nor U11816 (N_11816,N_11084,N_10045);
xor U11817 (N_11817,N_10220,N_11013);
nand U11818 (N_11818,N_10459,N_10183);
xnor U11819 (N_11819,N_10830,N_11069);
or U11820 (N_11820,N_10364,N_10640);
xor U11821 (N_11821,N_11094,N_11133);
and U11822 (N_11822,N_10631,N_11233);
xor U11823 (N_11823,N_10666,N_10452);
and U11824 (N_11824,N_10972,N_10098);
nor U11825 (N_11825,N_10173,N_10125);
or U11826 (N_11826,N_10081,N_11045);
nand U11827 (N_11827,N_11169,N_10381);
nor U11828 (N_11828,N_10530,N_10811);
nand U11829 (N_11829,N_10620,N_11163);
and U11830 (N_11830,N_10268,N_10895);
and U11831 (N_11831,N_10648,N_10223);
or U11832 (N_11832,N_10667,N_10168);
nand U11833 (N_11833,N_10239,N_10110);
or U11834 (N_11834,N_11191,N_10230);
xnor U11835 (N_11835,N_10980,N_10926);
xor U11836 (N_11836,N_11145,N_11004);
or U11837 (N_11837,N_10789,N_10954);
xnor U11838 (N_11838,N_10567,N_11031);
or U11839 (N_11839,N_10129,N_11240);
and U11840 (N_11840,N_11151,N_11117);
xor U11841 (N_11841,N_10992,N_10890);
and U11842 (N_11842,N_11211,N_10599);
xor U11843 (N_11843,N_10203,N_10734);
nor U11844 (N_11844,N_11146,N_10876);
nor U11845 (N_11845,N_11202,N_10182);
nor U11846 (N_11846,N_10214,N_11220);
or U11847 (N_11847,N_10024,N_10674);
nor U11848 (N_11848,N_10297,N_10854);
nand U11849 (N_11849,N_11134,N_10899);
xor U11850 (N_11850,N_10634,N_10767);
or U11851 (N_11851,N_10184,N_10856);
nor U11852 (N_11852,N_10562,N_10994);
or U11853 (N_11853,N_11109,N_10817);
and U11854 (N_11854,N_10794,N_11032);
xnor U11855 (N_11855,N_10787,N_10304);
xnor U11856 (N_11856,N_10621,N_10514);
xnor U11857 (N_11857,N_10339,N_10063);
and U11858 (N_11858,N_10301,N_10764);
and U11859 (N_11859,N_11105,N_11185);
or U11860 (N_11860,N_10357,N_11156);
and U11861 (N_11861,N_11120,N_10295);
or U11862 (N_11862,N_10719,N_10022);
nand U11863 (N_11863,N_10234,N_10555);
nand U11864 (N_11864,N_11064,N_10693);
nand U11865 (N_11865,N_10747,N_10503);
nand U11866 (N_11866,N_10099,N_10308);
xor U11867 (N_11867,N_10520,N_11124);
or U11868 (N_11868,N_10448,N_11139);
nand U11869 (N_11869,N_10506,N_10673);
or U11870 (N_11870,N_10950,N_10772);
or U11871 (N_11871,N_11234,N_10654);
nor U11872 (N_11872,N_10651,N_11171);
nand U11873 (N_11873,N_10374,N_11237);
xnor U11874 (N_11874,N_10083,N_10169);
and U11875 (N_11875,N_10700,N_10113);
xnor U11876 (N_11876,N_10157,N_11000);
nor U11877 (N_11877,N_10635,N_10058);
and U11878 (N_11878,N_10639,N_10593);
and U11879 (N_11879,N_10180,N_11069);
nand U11880 (N_11880,N_11189,N_11013);
and U11881 (N_11881,N_10502,N_10720);
nor U11882 (N_11882,N_10793,N_11231);
nor U11883 (N_11883,N_10620,N_10830);
nand U11884 (N_11884,N_10098,N_10637);
nor U11885 (N_11885,N_10239,N_11078);
nor U11886 (N_11886,N_11228,N_10169);
or U11887 (N_11887,N_10043,N_11188);
nor U11888 (N_11888,N_10455,N_10540);
or U11889 (N_11889,N_11004,N_10569);
xnor U11890 (N_11890,N_10473,N_10877);
xor U11891 (N_11891,N_10712,N_10698);
or U11892 (N_11892,N_11178,N_10264);
or U11893 (N_11893,N_11173,N_10099);
xnor U11894 (N_11894,N_11087,N_11060);
nor U11895 (N_11895,N_11059,N_10139);
and U11896 (N_11896,N_10996,N_10184);
or U11897 (N_11897,N_10495,N_10771);
nand U11898 (N_11898,N_10992,N_10105);
and U11899 (N_11899,N_10580,N_10496);
xor U11900 (N_11900,N_10679,N_10449);
or U11901 (N_11901,N_10514,N_10951);
nor U11902 (N_11902,N_11204,N_10422);
or U11903 (N_11903,N_11167,N_10137);
nand U11904 (N_11904,N_10920,N_11067);
and U11905 (N_11905,N_10017,N_10822);
nor U11906 (N_11906,N_11074,N_10776);
and U11907 (N_11907,N_10068,N_10595);
xor U11908 (N_11908,N_10524,N_10431);
and U11909 (N_11909,N_10346,N_11232);
nor U11910 (N_11910,N_10966,N_10544);
nor U11911 (N_11911,N_10866,N_10994);
nand U11912 (N_11912,N_11074,N_10102);
and U11913 (N_11913,N_11140,N_10878);
nor U11914 (N_11914,N_11081,N_10528);
nand U11915 (N_11915,N_10434,N_10755);
xor U11916 (N_11916,N_10542,N_10648);
or U11917 (N_11917,N_10801,N_11182);
and U11918 (N_11918,N_10107,N_10507);
and U11919 (N_11919,N_10216,N_10143);
xor U11920 (N_11920,N_10787,N_10162);
nand U11921 (N_11921,N_10468,N_10126);
xor U11922 (N_11922,N_10556,N_10101);
nor U11923 (N_11923,N_10889,N_10306);
or U11924 (N_11924,N_11111,N_10189);
nand U11925 (N_11925,N_10689,N_10268);
or U11926 (N_11926,N_10547,N_11154);
nor U11927 (N_11927,N_10528,N_10598);
nor U11928 (N_11928,N_10090,N_10700);
nor U11929 (N_11929,N_10372,N_10568);
and U11930 (N_11930,N_11021,N_11146);
or U11931 (N_11931,N_10371,N_10940);
xor U11932 (N_11932,N_10871,N_10709);
nor U11933 (N_11933,N_10539,N_10440);
nand U11934 (N_11934,N_11126,N_10322);
and U11935 (N_11935,N_10272,N_11021);
xor U11936 (N_11936,N_10825,N_10604);
or U11937 (N_11937,N_11198,N_10566);
and U11938 (N_11938,N_10638,N_10538);
xnor U11939 (N_11939,N_10364,N_10117);
xnor U11940 (N_11940,N_10767,N_11139);
xor U11941 (N_11941,N_10558,N_11037);
nor U11942 (N_11942,N_11122,N_10909);
nand U11943 (N_11943,N_10365,N_10823);
nand U11944 (N_11944,N_10294,N_10137);
and U11945 (N_11945,N_10988,N_10143);
xor U11946 (N_11946,N_10971,N_10970);
or U11947 (N_11947,N_10034,N_10933);
and U11948 (N_11948,N_10447,N_10287);
nor U11949 (N_11949,N_10997,N_10514);
xor U11950 (N_11950,N_10997,N_10758);
or U11951 (N_11951,N_10250,N_10426);
nor U11952 (N_11952,N_10202,N_11020);
nor U11953 (N_11953,N_10913,N_10677);
and U11954 (N_11954,N_10557,N_10492);
nor U11955 (N_11955,N_10910,N_11000);
xor U11956 (N_11956,N_11100,N_10815);
xor U11957 (N_11957,N_10842,N_11034);
or U11958 (N_11958,N_11078,N_10848);
nor U11959 (N_11959,N_10260,N_10646);
nor U11960 (N_11960,N_11058,N_10081);
xnor U11961 (N_11961,N_11043,N_10437);
xnor U11962 (N_11962,N_10305,N_10637);
nor U11963 (N_11963,N_10133,N_10196);
nor U11964 (N_11964,N_10969,N_11232);
and U11965 (N_11965,N_10338,N_10151);
nor U11966 (N_11966,N_11001,N_10669);
nand U11967 (N_11967,N_10659,N_10897);
or U11968 (N_11968,N_10586,N_10854);
xor U11969 (N_11969,N_10273,N_10792);
or U11970 (N_11970,N_10955,N_10153);
or U11971 (N_11971,N_10012,N_10930);
and U11972 (N_11972,N_10097,N_10250);
xnor U11973 (N_11973,N_10696,N_10139);
xor U11974 (N_11974,N_10612,N_10255);
or U11975 (N_11975,N_10843,N_11051);
or U11976 (N_11976,N_11006,N_10853);
or U11977 (N_11977,N_11087,N_10142);
or U11978 (N_11978,N_10199,N_10273);
or U11979 (N_11979,N_10058,N_10213);
and U11980 (N_11980,N_10191,N_10821);
nand U11981 (N_11981,N_10211,N_10356);
nor U11982 (N_11982,N_10260,N_10408);
and U11983 (N_11983,N_11241,N_10076);
nand U11984 (N_11984,N_11063,N_10111);
or U11985 (N_11985,N_11114,N_10767);
nand U11986 (N_11986,N_10541,N_10533);
or U11987 (N_11987,N_10558,N_10998);
and U11988 (N_11988,N_11017,N_10648);
nor U11989 (N_11989,N_10943,N_10482);
nor U11990 (N_11990,N_11116,N_10852);
and U11991 (N_11991,N_11148,N_10734);
nor U11992 (N_11992,N_10160,N_11020);
xor U11993 (N_11993,N_10087,N_11095);
nor U11994 (N_11994,N_10553,N_11236);
xor U11995 (N_11995,N_11182,N_10029);
nor U11996 (N_11996,N_11042,N_10728);
nor U11997 (N_11997,N_10342,N_10410);
or U11998 (N_11998,N_10444,N_11141);
nor U11999 (N_11999,N_10264,N_11004);
nand U12000 (N_12000,N_10133,N_10538);
nand U12001 (N_12001,N_10121,N_10969);
nor U12002 (N_12002,N_10091,N_10627);
nor U12003 (N_12003,N_10690,N_10967);
or U12004 (N_12004,N_10289,N_11160);
nand U12005 (N_12005,N_10694,N_11243);
or U12006 (N_12006,N_10571,N_10739);
nand U12007 (N_12007,N_11009,N_11006);
nor U12008 (N_12008,N_10367,N_10794);
nand U12009 (N_12009,N_10983,N_10976);
or U12010 (N_12010,N_10980,N_10540);
xor U12011 (N_12011,N_11152,N_11025);
and U12012 (N_12012,N_10531,N_11093);
nand U12013 (N_12013,N_10294,N_10619);
or U12014 (N_12014,N_10716,N_10786);
and U12015 (N_12015,N_10404,N_11043);
nor U12016 (N_12016,N_10971,N_10700);
xnor U12017 (N_12017,N_10315,N_10965);
nand U12018 (N_12018,N_10534,N_10735);
and U12019 (N_12019,N_10799,N_10821);
and U12020 (N_12020,N_10281,N_10243);
xnor U12021 (N_12021,N_10628,N_11103);
nor U12022 (N_12022,N_11062,N_10349);
or U12023 (N_12023,N_10341,N_11164);
nand U12024 (N_12024,N_10073,N_11076);
or U12025 (N_12025,N_10170,N_10417);
nand U12026 (N_12026,N_10517,N_10909);
nand U12027 (N_12027,N_10878,N_10733);
and U12028 (N_12028,N_11116,N_10242);
nand U12029 (N_12029,N_11081,N_10859);
xnor U12030 (N_12030,N_11241,N_10245);
xnor U12031 (N_12031,N_10471,N_10516);
nor U12032 (N_12032,N_11209,N_10036);
nor U12033 (N_12033,N_10346,N_10457);
nor U12034 (N_12034,N_11187,N_10801);
xor U12035 (N_12035,N_10138,N_10888);
nand U12036 (N_12036,N_11011,N_10326);
xnor U12037 (N_12037,N_10148,N_11182);
and U12038 (N_12038,N_10225,N_10342);
nor U12039 (N_12039,N_10133,N_10791);
xor U12040 (N_12040,N_10981,N_10846);
or U12041 (N_12041,N_10102,N_11035);
nor U12042 (N_12042,N_11188,N_10511);
nand U12043 (N_12043,N_11097,N_10227);
or U12044 (N_12044,N_10658,N_10155);
xnor U12045 (N_12045,N_10267,N_10791);
and U12046 (N_12046,N_10471,N_10218);
nand U12047 (N_12047,N_10125,N_10427);
or U12048 (N_12048,N_11248,N_10037);
nand U12049 (N_12049,N_10949,N_10242);
and U12050 (N_12050,N_11118,N_11082);
and U12051 (N_12051,N_11103,N_10412);
or U12052 (N_12052,N_10843,N_10899);
or U12053 (N_12053,N_11171,N_10929);
nor U12054 (N_12054,N_11228,N_10205);
or U12055 (N_12055,N_10916,N_11078);
nand U12056 (N_12056,N_10754,N_10391);
or U12057 (N_12057,N_10829,N_10822);
xor U12058 (N_12058,N_10633,N_10419);
or U12059 (N_12059,N_11016,N_11229);
nand U12060 (N_12060,N_10570,N_10557);
nor U12061 (N_12061,N_10260,N_10315);
or U12062 (N_12062,N_10034,N_10129);
nor U12063 (N_12063,N_11140,N_10338);
nand U12064 (N_12064,N_11034,N_10574);
nor U12065 (N_12065,N_10842,N_11145);
and U12066 (N_12066,N_10988,N_10331);
xnor U12067 (N_12067,N_10520,N_10197);
and U12068 (N_12068,N_10083,N_10790);
and U12069 (N_12069,N_11077,N_10884);
and U12070 (N_12070,N_10432,N_10978);
xor U12071 (N_12071,N_10721,N_10995);
and U12072 (N_12072,N_11132,N_10502);
nor U12073 (N_12073,N_10059,N_11035);
and U12074 (N_12074,N_10476,N_10187);
or U12075 (N_12075,N_11112,N_10907);
nand U12076 (N_12076,N_10875,N_10367);
and U12077 (N_12077,N_10337,N_10262);
xnor U12078 (N_12078,N_10952,N_10455);
nand U12079 (N_12079,N_11199,N_10063);
and U12080 (N_12080,N_10606,N_10991);
nand U12081 (N_12081,N_10742,N_10977);
nor U12082 (N_12082,N_10392,N_10662);
xnor U12083 (N_12083,N_10545,N_10183);
or U12084 (N_12084,N_10268,N_10188);
nor U12085 (N_12085,N_11078,N_10738);
nand U12086 (N_12086,N_11186,N_10057);
nor U12087 (N_12087,N_10488,N_11078);
nand U12088 (N_12088,N_10186,N_10697);
xor U12089 (N_12089,N_10309,N_11138);
nand U12090 (N_12090,N_10498,N_10631);
nand U12091 (N_12091,N_10572,N_10165);
xnor U12092 (N_12092,N_11005,N_10997);
xnor U12093 (N_12093,N_10594,N_10003);
and U12094 (N_12094,N_11092,N_10211);
nand U12095 (N_12095,N_10770,N_10219);
and U12096 (N_12096,N_10666,N_11189);
xnor U12097 (N_12097,N_10166,N_10570);
or U12098 (N_12098,N_10508,N_10303);
or U12099 (N_12099,N_10220,N_11014);
and U12100 (N_12100,N_11091,N_10132);
xnor U12101 (N_12101,N_11240,N_11245);
and U12102 (N_12102,N_10303,N_10127);
nor U12103 (N_12103,N_11220,N_10028);
nor U12104 (N_12104,N_10843,N_10453);
nor U12105 (N_12105,N_10663,N_10466);
nand U12106 (N_12106,N_11160,N_10689);
nor U12107 (N_12107,N_11201,N_10347);
xor U12108 (N_12108,N_11018,N_10796);
nor U12109 (N_12109,N_10705,N_11058);
nor U12110 (N_12110,N_10986,N_11208);
nor U12111 (N_12111,N_10703,N_10086);
and U12112 (N_12112,N_10374,N_10511);
or U12113 (N_12113,N_10686,N_10278);
nand U12114 (N_12114,N_11010,N_10740);
nor U12115 (N_12115,N_10118,N_10110);
or U12116 (N_12116,N_11242,N_10074);
and U12117 (N_12117,N_11212,N_10165);
and U12118 (N_12118,N_10428,N_10157);
xnor U12119 (N_12119,N_10106,N_10037);
and U12120 (N_12120,N_10249,N_10431);
or U12121 (N_12121,N_11054,N_10497);
xnor U12122 (N_12122,N_10850,N_11135);
and U12123 (N_12123,N_11084,N_10069);
xnor U12124 (N_12124,N_10631,N_11220);
xor U12125 (N_12125,N_10870,N_11188);
or U12126 (N_12126,N_10401,N_11197);
or U12127 (N_12127,N_10385,N_11213);
nor U12128 (N_12128,N_10906,N_10152);
and U12129 (N_12129,N_10752,N_10041);
nand U12130 (N_12130,N_10405,N_11168);
nor U12131 (N_12131,N_11127,N_10809);
and U12132 (N_12132,N_10986,N_10943);
xor U12133 (N_12133,N_10352,N_10052);
and U12134 (N_12134,N_11175,N_10596);
xor U12135 (N_12135,N_10520,N_10810);
or U12136 (N_12136,N_10878,N_11012);
nor U12137 (N_12137,N_11007,N_10625);
nand U12138 (N_12138,N_11184,N_10922);
nor U12139 (N_12139,N_11240,N_10592);
and U12140 (N_12140,N_11088,N_10733);
xor U12141 (N_12141,N_10523,N_10341);
nand U12142 (N_12142,N_10099,N_10827);
xor U12143 (N_12143,N_10436,N_11203);
nor U12144 (N_12144,N_11230,N_10064);
and U12145 (N_12145,N_10112,N_10295);
or U12146 (N_12146,N_10016,N_10549);
nand U12147 (N_12147,N_11134,N_10900);
nor U12148 (N_12148,N_11057,N_10753);
and U12149 (N_12149,N_11000,N_10061);
and U12150 (N_12150,N_10438,N_10852);
or U12151 (N_12151,N_10450,N_11039);
nand U12152 (N_12152,N_10877,N_10303);
or U12153 (N_12153,N_11132,N_11144);
or U12154 (N_12154,N_10532,N_10143);
and U12155 (N_12155,N_10762,N_11169);
or U12156 (N_12156,N_11025,N_11207);
xor U12157 (N_12157,N_10770,N_10012);
xor U12158 (N_12158,N_10198,N_10304);
nand U12159 (N_12159,N_10360,N_11048);
xor U12160 (N_12160,N_11095,N_11214);
xor U12161 (N_12161,N_10322,N_10275);
and U12162 (N_12162,N_10906,N_10610);
nor U12163 (N_12163,N_11138,N_10470);
or U12164 (N_12164,N_10381,N_11242);
nand U12165 (N_12165,N_11032,N_11125);
nor U12166 (N_12166,N_10106,N_10647);
and U12167 (N_12167,N_11179,N_10104);
xor U12168 (N_12168,N_10246,N_11140);
xor U12169 (N_12169,N_10547,N_11181);
xnor U12170 (N_12170,N_10482,N_10892);
or U12171 (N_12171,N_10430,N_11010);
nand U12172 (N_12172,N_10896,N_10510);
and U12173 (N_12173,N_10425,N_10128);
xnor U12174 (N_12174,N_11015,N_10549);
or U12175 (N_12175,N_10983,N_10764);
xnor U12176 (N_12176,N_10871,N_11025);
and U12177 (N_12177,N_10282,N_11062);
xor U12178 (N_12178,N_10787,N_10645);
and U12179 (N_12179,N_11045,N_10820);
and U12180 (N_12180,N_10201,N_10024);
nor U12181 (N_12181,N_11172,N_10490);
xnor U12182 (N_12182,N_10213,N_10296);
and U12183 (N_12183,N_10483,N_10049);
nor U12184 (N_12184,N_10483,N_10627);
xnor U12185 (N_12185,N_10633,N_10052);
nor U12186 (N_12186,N_10194,N_11193);
or U12187 (N_12187,N_10134,N_10229);
and U12188 (N_12188,N_10635,N_10275);
nor U12189 (N_12189,N_10939,N_10875);
nor U12190 (N_12190,N_10214,N_10179);
nor U12191 (N_12191,N_10881,N_10521);
xor U12192 (N_12192,N_11107,N_10904);
or U12193 (N_12193,N_10071,N_10714);
or U12194 (N_12194,N_10820,N_10515);
xor U12195 (N_12195,N_11177,N_10047);
and U12196 (N_12196,N_10652,N_11130);
and U12197 (N_12197,N_11143,N_10847);
xnor U12198 (N_12198,N_10585,N_10439);
or U12199 (N_12199,N_10272,N_10136);
nor U12200 (N_12200,N_10550,N_10384);
nor U12201 (N_12201,N_10720,N_10243);
nor U12202 (N_12202,N_10693,N_10345);
or U12203 (N_12203,N_10497,N_10390);
xor U12204 (N_12204,N_10974,N_10588);
xnor U12205 (N_12205,N_10910,N_10415);
nor U12206 (N_12206,N_10285,N_10174);
or U12207 (N_12207,N_11084,N_10337);
nand U12208 (N_12208,N_10747,N_10792);
or U12209 (N_12209,N_11221,N_10564);
or U12210 (N_12210,N_10696,N_10942);
or U12211 (N_12211,N_10983,N_10545);
xnor U12212 (N_12212,N_10945,N_10805);
nor U12213 (N_12213,N_10635,N_10479);
and U12214 (N_12214,N_10846,N_10373);
nor U12215 (N_12215,N_10980,N_10527);
and U12216 (N_12216,N_10666,N_10775);
nand U12217 (N_12217,N_10083,N_10545);
xor U12218 (N_12218,N_10315,N_10034);
nor U12219 (N_12219,N_10200,N_10169);
nor U12220 (N_12220,N_10202,N_10456);
xor U12221 (N_12221,N_10004,N_10817);
nand U12222 (N_12222,N_10161,N_11068);
and U12223 (N_12223,N_10983,N_10428);
and U12224 (N_12224,N_10337,N_10446);
nor U12225 (N_12225,N_10326,N_10467);
nor U12226 (N_12226,N_10538,N_10712);
nor U12227 (N_12227,N_10498,N_10632);
and U12228 (N_12228,N_10127,N_10830);
nor U12229 (N_12229,N_10822,N_10880);
and U12230 (N_12230,N_10922,N_10181);
and U12231 (N_12231,N_10780,N_10957);
nor U12232 (N_12232,N_10283,N_10214);
nor U12233 (N_12233,N_10786,N_10009);
nand U12234 (N_12234,N_11058,N_10822);
nand U12235 (N_12235,N_10929,N_10020);
or U12236 (N_12236,N_10782,N_10160);
xor U12237 (N_12237,N_10909,N_10375);
and U12238 (N_12238,N_10067,N_10448);
nand U12239 (N_12239,N_11122,N_10954);
nor U12240 (N_12240,N_10879,N_10647);
xnor U12241 (N_12241,N_10232,N_10975);
nor U12242 (N_12242,N_10296,N_10807);
xnor U12243 (N_12243,N_10053,N_10917);
or U12244 (N_12244,N_10765,N_10354);
and U12245 (N_12245,N_10280,N_10791);
nor U12246 (N_12246,N_11232,N_10471);
or U12247 (N_12247,N_10235,N_11164);
nand U12248 (N_12248,N_10504,N_10763);
and U12249 (N_12249,N_10973,N_10483);
xnor U12250 (N_12250,N_10685,N_10881);
or U12251 (N_12251,N_10747,N_11248);
xor U12252 (N_12252,N_10069,N_10134);
and U12253 (N_12253,N_10595,N_10849);
nand U12254 (N_12254,N_10671,N_10621);
xor U12255 (N_12255,N_10819,N_11069);
or U12256 (N_12256,N_10646,N_11094);
or U12257 (N_12257,N_10505,N_11038);
xnor U12258 (N_12258,N_10644,N_10081);
xnor U12259 (N_12259,N_11035,N_10430);
nand U12260 (N_12260,N_10815,N_10459);
xnor U12261 (N_12261,N_11070,N_10714);
or U12262 (N_12262,N_10960,N_10876);
nor U12263 (N_12263,N_11216,N_11074);
nand U12264 (N_12264,N_10471,N_10207);
and U12265 (N_12265,N_10676,N_10954);
nor U12266 (N_12266,N_11218,N_10218);
or U12267 (N_12267,N_10161,N_10820);
nand U12268 (N_12268,N_11123,N_10552);
nand U12269 (N_12269,N_10381,N_11199);
nor U12270 (N_12270,N_10416,N_11034);
nand U12271 (N_12271,N_11162,N_10917);
and U12272 (N_12272,N_11108,N_10748);
and U12273 (N_12273,N_10240,N_11012);
nor U12274 (N_12274,N_10821,N_10569);
or U12275 (N_12275,N_10468,N_10740);
and U12276 (N_12276,N_10322,N_10319);
and U12277 (N_12277,N_10381,N_11173);
xnor U12278 (N_12278,N_11149,N_11004);
and U12279 (N_12279,N_10937,N_10439);
or U12280 (N_12280,N_10839,N_10362);
nand U12281 (N_12281,N_10713,N_10828);
and U12282 (N_12282,N_10055,N_10820);
nor U12283 (N_12283,N_10750,N_10651);
xnor U12284 (N_12284,N_10120,N_10620);
and U12285 (N_12285,N_10563,N_10708);
or U12286 (N_12286,N_10246,N_10795);
nor U12287 (N_12287,N_10335,N_10992);
nand U12288 (N_12288,N_10966,N_10017);
and U12289 (N_12289,N_10388,N_11203);
xnor U12290 (N_12290,N_10146,N_10477);
nand U12291 (N_12291,N_11076,N_10298);
nor U12292 (N_12292,N_11127,N_10827);
nor U12293 (N_12293,N_10563,N_10440);
or U12294 (N_12294,N_10326,N_11115);
and U12295 (N_12295,N_10481,N_10170);
xor U12296 (N_12296,N_10527,N_11151);
xnor U12297 (N_12297,N_10822,N_10035);
and U12298 (N_12298,N_10895,N_11101);
nor U12299 (N_12299,N_10835,N_10007);
nor U12300 (N_12300,N_10769,N_11096);
xor U12301 (N_12301,N_10059,N_11053);
and U12302 (N_12302,N_10160,N_11068);
nand U12303 (N_12303,N_10933,N_10173);
nor U12304 (N_12304,N_10698,N_10918);
xor U12305 (N_12305,N_10954,N_10337);
nand U12306 (N_12306,N_10642,N_10643);
nor U12307 (N_12307,N_10106,N_10923);
and U12308 (N_12308,N_10838,N_10126);
and U12309 (N_12309,N_10177,N_10088);
nor U12310 (N_12310,N_10836,N_10600);
nand U12311 (N_12311,N_10459,N_11031);
and U12312 (N_12312,N_10653,N_10935);
nand U12313 (N_12313,N_10114,N_10402);
nor U12314 (N_12314,N_10439,N_11118);
nor U12315 (N_12315,N_11126,N_10840);
nor U12316 (N_12316,N_10546,N_10886);
nand U12317 (N_12317,N_10917,N_10760);
xnor U12318 (N_12318,N_10012,N_10933);
or U12319 (N_12319,N_10511,N_10856);
nand U12320 (N_12320,N_10530,N_10578);
xnor U12321 (N_12321,N_11013,N_10436);
xnor U12322 (N_12322,N_11085,N_10686);
and U12323 (N_12323,N_10267,N_10886);
and U12324 (N_12324,N_10776,N_10254);
and U12325 (N_12325,N_11234,N_10209);
nor U12326 (N_12326,N_10684,N_10244);
xor U12327 (N_12327,N_10754,N_10746);
nor U12328 (N_12328,N_10608,N_10846);
nor U12329 (N_12329,N_10745,N_10689);
and U12330 (N_12330,N_10799,N_10310);
or U12331 (N_12331,N_10780,N_10442);
or U12332 (N_12332,N_10995,N_10159);
xor U12333 (N_12333,N_10756,N_10250);
nor U12334 (N_12334,N_10538,N_10788);
nor U12335 (N_12335,N_10288,N_10388);
xor U12336 (N_12336,N_10358,N_10851);
nor U12337 (N_12337,N_11127,N_10938);
or U12338 (N_12338,N_10784,N_10593);
nor U12339 (N_12339,N_10825,N_10183);
nor U12340 (N_12340,N_10900,N_10663);
or U12341 (N_12341,N_10346,N_10544);
or U12342 (N_12342,N_10257,N_10088);
nand U12343 (N_12343,N_11016,N_11146);
nor U12344 (N_12344,N_11041,N_10989);
or U12345 (N_12345,N_10210,N_10797);
and U12346 (N_12346,N_10238,N_10120);
xor U12347 (N_12347,N_10634,N_10925);
or U12348 (N_12348,N_10240,N_10556);
nand U12349 (N_12349,N_10415,N_10474);
or U12350 (N_12350,N_10211,N_10084);
nor U12351 (N_12351,N_10533,N_10725);
and U12352 (N_12352,N_10037,N_10681);
nor U12353 (N_12353,N_10599,N_10937);
nor U12354 (N_12354,N_10297,N_10608);
nor U12355 (N_12355,N_10241,N_10065);
nand U12356 (N_12356,N_10978,N_10280);
nand U12357 (N_12357,N_10517,N_10062);
nor U12358 (N_12358,N_10718,N_10510);
xnor U12359 (N_12359,N_10571,N_11247);
nor U12360 (N_12360,N_11172,N_10342);
xnor U12361 (N_12361,N_10168,N_10607);
nor U12362 (N_12362,N_10393,N_10414);
and U12363 (N_12363,N_10331,N_10494);
and U12364 (N_12364,N_10309,N_10738);
nor U12365 (N_12365,N_10714,N_10250);
or U12366 (N_12366,N_10644,N_10020);
xor U12367 (N_12367,N_10280,N_11152);
nor U12368 (N_12368,N_10321,N_11066);
and U12369 (N_12369,N_11188,N_10575);
and U12370 (N_12370,N_10313,N_10681);
xor U12371 (N_12371,N_10653,N_10615);
nor U12372 (N_12372,N_10976,N_10180);
nand U12373 (N_12373,N_10360,N_10514);
and U12374 (N_12374,N_10500,N_10714);
xor U12375 (N_12375,N_10713,N_10561);
xor U12376 (N_12376,N_11033,N_10986);
nand U12377 (N_12377,N_11082,N_10766);
and U12378 (N_12378,N_10105,N_10430);
nor U12379 (N_12379,N_10519,N_10050);
and U12380 (N_12380,N_10280,N_10966);
nor U12381 (N_12381,N_10043,N_11245);
or U12382 (N_12382,N_10116,N_10110);
or U12383 (N_12383,N_10220,N_10242);
and U12384 (N_12384,N_10281,N_11010);
nor U12385 (N_12385,N_10020,N_10931);
and U12386 (N_12386,N_10520,N_11128);
or U12387 (N_12387,N_10918,N_10673);
xnor U12388 (N_12388,N_10554,N_10488);
and U12389 (N_12389,N_11065,N_10854);
xor U12390 (N_12390,N_10147,N_11103);
and U12391 (N_12391,N_10744,N_11051);
nand U12392 (N_12392,N_10103,N_10277);
xnor U12393 (N_12393,N_10057,N_11170);
and U12394 (N_12394,N_10382,N_10606);
and U12395 (N_12395,N_10518,N_10756);
nand U12396 (N_12396,N_10542,N_10635);
nor U12397 (N_12397,N_10128,N_11245);
nand U12398 (N_12398,N_10102,N_11244);
xor U12399 (N_12399,N_10026,N_11033);
xnor U12400 (N_12400,N_10931,N_10958);
or U12401 (N_12401,N_10680,N_10514);
xnor U12402 (N_12402,N_11157,N_10403);
and U12403 (N_12403,N_11196,N_10814);
xor U12404 (N_12404,N_10421,N_10054);
nor U12405 (N_12405,N_10095,N_10089);
or U12406 (N_12406,N_10759,N_10998);
or U12407 (N_12407,N_10441,N_11233);
nand U12408 (N_12408,N_10480,N_10812);
nor U12409 (N_12409,N_10053,N_11217);
or U12410 (N_12410,N_11151,N_10963);
or U12411 (N_12411,N_10230,N_10376);
and U12412 (N_12412,N_10609,N_10697);
xor U12413 (N_12413,N_10363,N_10837);
or U12414 (N_12414,N_10359,N_10660);
xnor U12415 (N_12415,N_11205,N_11033);
nor U12416 (N_12416,N_10009,N_10264);
nor U12417 (N_12417,N_10988,N_10008);
nand U12418 (N_12418,N_10103,N_10482);
nor U12419 (N_12419,N_10091,N_10903);
xor U12420 (N_12420,N_10651,N_10041);
and U12421 (N_12421,N_10988,N_10180);
nor U12422 (N_12422,N_11244,N_10201);
and U12423 (N_12423,N_10666,N_11079);
and U12424 (N_12424,N_10112,N_11141);
or U12425 (N_12425,N_10872,N_10952);
nor U12426 (N_12426,N_10246,N_10982);
nand U12427 (N_12427,N_10721,N_10133);
xor U12428 (N_12428,N_10496,N_10030);
xor U12429 (N_12429,N_10761,N_11046);
nand U12430 (N_12430,N_10174,N_10121);
nand U12431 (N_12431,N_10916,N_10640);
nand U12432 (N_12432,N_10339,N_10691);
nor U12433 (N_12433,N_10707,N_10435);
nand U12434 (N_12434,N_10519,N_11242);
and U12435 (N_12435,N_11220,N_10736);
nand U12436 (N_12436,N_10137,N_10861);
or U12437 (N_12437,N_10245,N_10486);
or U12438 (N_12438,N_10268,N_11046);
xor U12439 (N_12439,N_11040,N_10226);
and U12440 (N_12440,N_10605,N_10440);
nor U12441 (N_12441,N_10048,N_11091);
nor U12442 (N_12442,N_10739,N_10032);
or U12443 (N_12443,N_11030,N_10363);
nor U12444 (N_12444,N_10447,N_11219);
and U12445 (N_12445,N_10230,N_11004);
or U12446 (N_12446,N_10718,N_10693);
nand U12447 (N_12447,N_11080,N_10476);
xnor U12448 (N_12448,N_10136,N_10860);
nor U12449 (N_12449,N_11180,N_11170);
xnor U12450 (N_12450,N_11168,N_11081);
and U12451 (N_12451,N_10525,N_10379);
nor U12452 (N_12452,N_11179,N_10599);
and U12453 (N_12453,N_11101,N_10391);
or U12454 (N_12454,N_10282,N_10818);
xnor U12455 (N_12455,N_10252,N_10391);
nand U12456 (N_12456,N_10426,N_10051);
nand U12457 (N_12457,N_10034,N_10330);
nand U12458 (N_12458,N_11125,N_10351);
nand U12459 (N_12459,N_11022,N_10737);
nor U12460 (N_12460,N_10703,N_10989);
or U12461 (N_12461,N_11072,N_11158);
and U12462 (N_12462,N_10170,N_10355);
or U12463 (N_12463,N_10545,N_11200);
nor U12464 (N_12464,N_10716,N_10441);
xor U12465 (N_12465,N_10503,N_11086);
and U12466 (N_12466,N_10873,N_10308);
nor U12467 (N_12467,N_10957,N_10753);
or U12468 (N_12468,N_11156,N_11242);
nand U12469 (N_12469,N_11074,N_10599);
nor U12470 (N_12470,N_10013,N_10107);
nor U12471 (N_12471,N_11120,N_10548);
or U12472 (N_12472,N_10932,N_10154);
xor U12473 (N_12473,N_11185,N_10603);
or U12474 (N_12474,N_10621,N_11144);
nand U12475 (N_12475,N_10057,N_11090);
xnor U12476 (N_12476,N_11190,N_10669);
xnor U12477 (N_12477,N_10510,N_10175);
nand U12478 (N_12478,N_11014,N_10776);
xnor U12479 (N_12479,N_10541,N_10296);
xor U12480 (N_12480,N_10705,N_10993);
xor U12481 (N_12481,N_10681,N_10169);
and U12482 (N_12482,N_10913,N_10289);
nor U12483 (N_12483,N_10624,N_10005);
xor U12484 (N_12484,N_11218,N_10469);
xnor U12485 (N_12485,N_10034,N_10067);
nand U12486 (N_12486,N_10289,N_10556);
nor U12487 (N_12487,N_11105,N_10016);
xor U12488 (N_12488,N_11042,N_11223);
xor U12489 (N_12489,N_10732,N_10011);
nand U12490 (N_12490,N_10864,N_10360);
nor U12491 (N_12491,N_10072,N_10010);
and U12492 (N_12492,N_10463,N_10109);
and U12493 (N_12493,N_10357,N_10187);
nor U12494 (N_12494,N_10744,N_10231);
or U12495 (N_12495,N_11042,N_10189);
nand U12496 (N_12496,N_10884,N_10541);
nand U12497 (N_12497,N_10485,N_10157);
nor U12498 (N_12498,N_10374,N_11131);
xor U12499 (N_12499,N_11076,N_10730);
nand U12500 (N_12500,N_11872,N_11923);
nand U12501 (N_12501,N_11540,N_11881);
nand U12502 (N_12502,N_12044,N_11570);
nor U12503 (N_12503,N_12420,N_11632);
nand U12504 (N_12504,N_11522,N_12335);
nand U12505 (N_12505,N_11265,N_12170);
xor U12506 (N_12506,N_11654,N_12314);
nor U12507 (N_12507,N_11481,N_11940);
xor U12508 (N_12508,N_12412,N_11322);
nand U12509 (N_12509,N_12157,N_12297);
nor U12510 (N_12510,N_12180,N_11738);
nor U12511 (N_12511,N_11907,N_11786);
and U12512 (N_12512,N_12199,N_12103);
xor U12513 (N_12513,N_12264,N_11799);
or U12514 (N_12514,N_12267,N_11561);
nand U12515 (N_12515,N_11379,N_11701);
nor U12516 (N_12516,N_11966,N_12194);
nand U12517 (N_12517,N_11502,N_12150);
and U12518 (N_12518,N_11435,N_11480);
xor U12519 (N_12519,N_12275,N_11347);
or U12520 (N_12520,N_12298,N_11539);
xor U12521 (N_12521,N_11696,N_11396);
and U12522 (N_12522,N_12413,N_11357);
and U12523 (N_12523,N_12415,N_12123);
nor U12524 (N_12524,N_11846,N_12059);
and U12525 (N_12525,N_12307,N_12282);
nand U12526 (N_12526,N_12159,N_12033);
nor U12527 (N_12527,N_11600,N_11392);
nor U12528 (N_12528,N_12151,N_11891);
and U12529 (N_12529,N_12001,N_12365);
or U12530 (N_12530,N_11729,N_11721);
nor U12531 (N_12531,N_12014,N_12333);
and U12532 (N_12532,N_11835,N_11301);
xnor U12533 (N_12533,N_11535,N_11732);
nor U12534 (N_12534,N_11817,N_11971);
nor U12535 (N_12535,N_11429,N_11684);
nand U12536 (N_12536,N_12078,N_11767);
and U12537 (N_12537,N_11884,N_12371);
and U12538 (N_12538,N_12010,N_11758);
xnor U12539 (N_12539,N_12056,N_12035);
nand U12540 (N_12540,N_11517,N_11459);
and U12541 (N_12541,N_11713,N_11501);
and U12542 (N_12542,N_11290,N_12337);
or U12543 (N_12543,N_12435,N_11530);
nor U12544 (N_12544,N_12012,N_12254);
xnor U12545 (N_12545,N_11278,N_12479);
xnor U12546 (N_12546,N_11993,N_12030);
nand U12547 (N_12547,N_11267,N_11311);
nor U12548 (N_12548,N_11507,N_11462);
nand U12549 (N_12549,N_12469,N_11682);
xnor U12550 (N_12550,N_12249,N_12156);
nand U12551 (N_12551,N_11860,N_11453);
nand U12552 (N_12552,N_11482,N_12160);
nor U12553 (N_12553,N_12409,N_12467);
nand U12554 (N_12554,N_12009,N_11567);
nand U12555 (N_12555,N_11497,N_11554);
and U12556 (N_12556,N_12101,N_11805);
xor U12557 (N_12557,N_11709,N_12146);
xnor U12558 (N_12558,N_12441,N_11314);
nand U12559 (N_12559,N_11909,N_12223);
and U12560 (N_12560,N_11924,N_12106);
nand U12561 (N_12561,N_11773,N_12179);
nand U12562 (N_12562,N_11927,N_11956);
nor U12563 (N_12563,N_12302,N_11363);
nand U12564 (N_12564,N_11621,N_11663);
nor U12565 (N_12565,N_12144,N_11395);
xor U12566 (N_12566,N_12168,N_11902);
xnor U12567 (N_12567,N_11585,N_12085);
or U12568 (N_12568,N_12212,N_12434);
or U12569 (N_12569,N_11829,N_11740);
nand U12570 (N_12570,N_12060,N_11269);
nand U12571 (N_12571,N_12325,N_11515);
or U12572 (N_12572,N_12155,N_11417);
nand U12573 (N_12573,N_11580,N_11988);
or U12574 (N_12574,N_11910,N_12366);
or U12575 (N_12575,N_11446,N_11270);
xnor U12576 (N_12576,N_12494,N_12131);
xor U12577 (N_12577,N_11808,N_12358);
nand U12578 (N_12578,N_11575,N_11593);
xnor U12579 (N_12579,N_12465,N_12067);
nand U12580 (N_12580,N_11516,N_12000);
or U12581 (N_12581,N_12036,N_12246);
nor U12582 (N_12582,N_11834,N_12100);
nor U12583 (N_12583,N_11430,N_12384);
nor U12584 (N_12584,N_12104,N_12090);
or U12585 (N_12585,N_11411,N_11936);
nor U12586 (N_12586,N_11282,N_12253);
xnor U12587 (N_12587,N_12315,N_12008);
or U12588 (N_12588,N_12174,N_11306);
or U12589 (N_12589,N_11316,N_12236);
xnor U12590 (N_12590,N_11777,N_12427);
nor U12591 (N_12591,N_12062,N_12488);
nor U12592 (N_12592,N_11999,N_12041);
nand U12593 (N_12593,N_11370,N_11707);
nand U12594 (N_12594,N_12079,N_11557);
and U12595 (N_12595,N_11782,N_11486);
or U12596 (N_12596,N_11926,N_11420);
or U12597 (N_12597,N_12265,N_11827);
or U12598 (N_12598,N_11765,N_11665);
or U12599 (N_12599,N_12177,N_11286);
nand U12600 (N_12600,N_11353,N_11399);
or U12601 (N_12601,N_11596,N_12300);
xor U12602 (N_12602,N_12342,N_12122);
and U12603 (N_12603,N_11868,N_12017);
and U12604 (N_12604,N_11636,N_11716);
or U12605 (N_12605,N_12232,N_11293);
nor U12606 (N_12606,N_12225,N_11438);
or U12607 (N_12607,N_11727,N_11785);
or U12608 (N_12608,N_11783,N_12383);
and U12609 (N_12609,N_12181,N_12483);
and U12610 (N_12610,N_11886,N_11376);
nor U12611 (N_12611,N_11662,N_11629);
xnor U12612 (N_12612,N_12252,N_12048);
nand U12613 (N_12613,N_11336,N_11659);
or U12614 (N_12614,N_12098,N_12065);
and U12615 (N_12615,N_11953,N_12481);
and U12616 (N_12616,N_11700,N_11616);
and U12617 (N_12617,N_11869,N_11472);
nand U12618 (N_12618,N_11640,N_11888);
nor U12619 (N_12619,N_12353,N_11615);
or U12620 (N_12620,N_12007,N_11870);
xnor U12621 (N_12621,N_11763,N_12118);
nor U12622 (N_12622,N_11768,N_12096);
and U12623 (N_12623,N_11341,N_12113);
and U12624 (N_12624,N_11813,N_12499);
nand U12625 (N_12625,N_11529,N_11667);
xnor U12626 (N_12626,N_12217,N_11905);
and U12627 (N_12627,N_12140,N_12327);
nand U12628 (N_12628,N_11444,N_12322);
or U12629 (N_12629,N_12206,N_12105);
or U12630 (N_12630,N_11712,N_12152);
nand U12631 (N_12631,N_11979,N_11719);
nand U12632 (N_12632,N_12445,N_12442);
nor U12633 (N_12633,N_12432,N_11352);
and U12634 (N_12634,N_11578,N_11508);
nor U12635 (N_12635,N_11518,N_11441);
nor U12636 (N_12636,N_11449,N_11963);
and U12637 (N_12637,N_11851,N_12373);
xor U12638 (N_12638,N_11724,N_12114);
or U12639 (N_12639,N_11277,N_11503);
or U12640 (N_12640,N_11967,N_12359);
nand U12641 (N_12641,N_11545,N_11349);
xor U12642 (N_12642,N_11769,N_12320);
and U12643 (N_12643,N_11690,N_11405);
xor U12644 (N_12644,N_11258,N_11626);
nor U12645 (N_12645,N_11980,N_12350);
xnor U12646 (N_12646,N_11266,N_11959);
or U12647 (N_12647,N_11549,N_11837);
xnor U12648 (N_12648,N_12295,N_11646);
or U12649 (N_12649,N_11283,N_11833);
or U12650 (N_12650,N_12378,N_12013);
xor U12651 (N_12651,N_11794,N_11468);
nand U12652 (N_12652,N_12002,N_11982);
nor U12653 (N_12653,N_11898,N_11380);
xnor U12654 (N_12654,N_12380,N_11276);
nor U12655 (N_12655,N_12461,N_11630);
or U12656 (N_12656,N_12169,N_11505);
nor U12657 (N_12657,N_11759,N_11873);
xor U12658 (N_12658,N_12074,N_11861);
or U12659 (N_12659,N_12478,N_12063);
xor U12660 (N_12660,N_11698,N_11252);
nand U12661 (N_12661,N_12317,N_11491);
xnor U12662 (N_12662,N_11460,N_11866);
xor U12663 (N_12663,N_12319,N_12278);
nor U12664 (N_12664,N_12258,N_11398);
xor U12665 (N_12665,N_11677,N_12095);
xor U12666 (N_12666,N_11975,N_11487);
xor U12667 (N_12667,N_12238,N_11296);
nand U12668 (N_12668,N_11281,N_11961);
nor U12669 (N_12669,N_11694,N_12287);
or U12670 (N_12670,N_12016,N_12395);
xor U12671 (N_12671,N_12397,N_12487);
and U12672 (N_12672,N_12021,N_12430);
xor U12673 (N_12673,N_12471,N_11431);
xnor U12674 (N_12674,N_11345,N_11594);
or U12675 (N_12675,N_12352,N_11423);
and U12676 (N_12676,N_11402,N_11774);
or U12677 (N_12677,N_11984,N_12042);
nor U12678 (N_12678,N_11974,N_11815);
or U12679 (N_12679,N_11440,N_12326);
xor U12680 (N_12680,N_11302,N_12229);
nand U12681 (N_12681,N_11259,N_12178);
nand U12682 (N_12682,N_11416,N_11744);
nand U12683 (N_12683,N_11401,N_12291);
nor U12684 (N_12684,N_12220,N_11737);
or U12685 (N_12685,N_11915,N_12052);
nand U12686 (N_12686,N_11917,N_11351);
xnor U12687 (N_12687,N_12072,N_12443);
nor U12688 (N_12688,N_11819,N_11770);
or U12689 (N_12689,N_12403,N_12083);
and U12690 (N_12690,N_12490,N_11288);
or U12691 (N_12691,N_12226,N_11775);
and U12692 (N_12692,N_11573,N_12454);
and U12693 (N_12693,N_12200,N_11668);
nand U12694 (N_12694,N_11458,N_12323);
nand U12695 (N_12695,N_11825,N_12474);
nor U12696 (N_12696,N_11928,N_12480);
and U12697 (N_12697,N_11386,N_11525);
and U12698 (N_12698,N_12329,N_12496);
or U12699 (N_12699,N_12354,N_11552);
nor U12700 (N_12700,N_12004,N_11356);
nor U12701 (N_12701,N_12192,N_11367);
nor U12702 (N_12702,N_11736,N_12289);
xor U12703 (N_12703,N_11781,N_11875);
nand U12704 (N_12704,N_12069,N_12316);
xnor U12705 (N_12705,N_12251,N_11368);
or U12706 (N_12706,N_12112,N_12346);
xnor U12707 (N_12707,N_12362,N_11731);
nand U12708 (N_12708,N_12448,N_11317);
or U12709 (N_12709,N_12234,N_12167);
xor U12710 (N_12710,N_11467,N_11421);
xnor U12711 (N_12711,N_12279,N_11796);
xor U12712 (N_12712,N_11921,N_11830);
or U12713 (N_12713,N_11746,N_11795);
and U12714 (N_12714,N_12129,N_11498);
or U12715 (N_12715,N_12215,N_11275);
and U12716 (N_12716,N_12185,N_12293);
and U12717 (N_12717,N_12040,N_11887);
nand U12718 (N_12718,N_12311,N_12050);
nand U12719 (N_12719,N_12489,N_12255);
nand U12720 (N_12720,N_11378,N_11843);
and U12721 (N_12721,N_11653,N_12459);
xnor U12722 (N_12722,N_11673,N_12401);
or U12723 (N_12723,N_12039,N_11894);
nor U12724 (N_12724,N_12141,N_11930);
and U12725 (N_12725,N_11918,N_11279);
nand U12726 (N_12726,N_11251,N_12273);
xor U12727 (N_12727,N_12257,N_11569);
nand U12728 (N_12728,N_11790,N_12093);
or U12729 (N_12729,N_12262,N_11832);
nand U12730 (N_12730,N_11285,N_12283);
or U12731 (N_12731,N_11602,N_11330);
and U12732 (N_12732,N_12472,N_12451);
nand U12733 (N_12733,N_11305,N_11666);
nand U12734 (N_12734,N_11704,N_11849);
nor U12735 (N_12735,N_11315,N_12391);
and U12736 (N_12736,N_11344,N_11893);
and U12737 (N_12737,N_11555,N_11867);
nor U12738 (N_12738,N_11681,N_11726);
xor U12739 (N_12739,N_12306,N_11537);
xor U12740 (N_12740,N_11298,N_12284);
and U12741 (N_12741,N_11513,N_11939);
xnor U12742 (N_12742,N_12055,N_12221);
xor U12743 (N_12743,N_11307,N_11976);
and U12744 (N_12744,N_11526,N_11675);
nor U12745 (N_12745,N_11641,N_11821);
or U12746 (N_12746,N_11261,N_12184);
xor U12747 (N_12747,N_11609,N_11958);
or U12748 (N_12748,N_11346,N_11711);
nand U12749 (N_12749,N_12076,N_11572);
nor U12750 (N_12750,N_11664,N_11280);
nand U12751 (N_12751,N_12020,N_11533);
xor U12752 (N_12752,N_12276,N_12125);
or U12753 (N_12753,N_11735,N_11295);
or U12754 (N_12754,N_12439,N_11824);
xnor U12755 (N_12755,N_12386,N_12368);
and U12756 (N_12756,N_12405,N_11360);
or U12757 (N_12757,N_12071,N_11343);
nand U12758 (N_12758,N_11550,N_11424);
or U12759 (N_12759,N_11553,N_12292);
and U12760 (N_12760,N_12450,N_12025);
or U12761 (N_12761,N_11614,N_12303);
or U12762 (N_12762,N_12037,N_12476);
and U12763 (N_12763,N_11692,N_11433);
nor U12764 (N_12764,N_12449,N_12228);
nand U12765 (N_12765,N_11913,N_12235);
nor U12766 (N_12766,N_12338,N_11257);
nand U12767 (N_12767,N_12374,N_12422);
nor U12768 (N_12768,N_12107,N_11253);
nor U12769 (N_12769,N_11705,N_11509);
nand U12770 (N_12770,N_11916,N_12018);
or U12771 (N_12771,N_12428,N_11787);
xnor U12772 (N_12772,N_11500,N_12193);
nor U12773 (N_12773,N_11685,N_11478);
xnor U12774 (N_12774,N_11457,N_12204);
or U12775 (N_12775,N_11695,N_11826);
nor U12776 (N_12776,N_11865,N_12202);
xor U12777 (N_12777,N_11853,N_12147);
or U12778 (N_12778,N_12187,N_11947);
or U12779 (N_12779,N_12121,N_11670);
nor U12780 (N_12780,N_11359,N_11645);
nand U12781 (N_12781,N_11906,N_11327);
nand U12782 (N_12782,N_12110,N_11941);
and U12783 (N_12783,N_11254,N_11320);
nand U12784 (N_12784,N_11582,N_11328);
nor U12785 (N_12785,N_11605,N_11876);
nor U12786 (N_12786,N_12058,N_12208);
or U12787 (N_12787,N_12334,N_11571);
and U12788 (N_12788,N_11818,N_12134);
nor U12789 (N_12789,N_12046,N_11644);
and U12790 (N_12790,N_11754,N_12089);
nor U12791 (N_12791,N_12308,N_11461);
xor U12792 (N_12792,N_12066,N_11669);
nand U12793 (N_12793,N_11334,N_11960);
or U12794 (N_12794,N_11914,N_11622);
nor U12795 (N_12795,N_12357,N_11426);
or U12796 (N_12796,N_12099,N_11590);
or U12797 (N_12797,N_12266,N_11784);
or U12798 (N_12798,N_12116,N_11772);
xnor U12799 (N_12799,N_11836,N_11776);
xnor U12800 (N_12800,N_12186,N_11403);
or U12801 (N_12801,N_11598,N_11496);
or U12802 (N_12802,N_12064,N_11532);
nor U12803 (N_12803,N_11627,N_12493);
and U12804 (N_12804,N_12305,N_11932);
or U12805 (N_12805,N_12233,N_11452);
xnor U12806 (N_12806,N_11427,N_11948);
and U12807 (N_12807,N_11566,N_11908);
xor U12808 (N_12808,N_12355,N_11450);
or U12809 (N_12809,N_12111,N_11688);
xnor U12810 (N_12810,N_12477,N_12201);
xor U12811 (N_12811,N_11466,N_11400);
or U12812 (N_12812,N_12213,N_11985);
or U12813 (N_12813,N_11374,N_12138);
nand U12814 (N_12814,N_12288,N_12361);
nand U12815 (N_12815,N_12222,N_11965);
xor U12816 (N_12816,N_11633,N_11741);
and U12817 (N_12817,N_12119,N_11862);
or U12818 (N_12818,N_11543,N_12497);
or U12819 (N_12819,N_12117,N_12458);
xnor U12820 (N_12820,N_12363,N_11952);
xnor U12821 (N_12821,N_11548,N_11986);
and U12822 (N_12822,N_12348,N_12456);
and U12823 (N_12823,N_12049,N_11877);
nor U12824 (N_12824,N_12043,N_11895);
and U12825 (N_12825,N_11250,N_11599);
nand U12826 (N_12826,N_12207,N_12047);
and U12827 (N_12827,N_12124,N_11755);
and U12828 (N_12828,N_11384,N_11271);
or U12829 (N_12829,N_12166,N_11514);
or U12830 (N_12830,N_11262,N_11510);
or U12831 (N_12831,N_11992,N_11800);
nor U12832 (N_12832,N_12312,N_11313);
xor U12833 (N_12833,N_11946,N_11848);
nor U12834 (N_12834,N_12195,N_11998);
nor U12835 (N_12835,N_12128,N_11595);
and U12836 (N_12836,N_12163,N_11889);
nand U12837 (N_12837,N_12321,N_11331);
xor U12838 (N_12838,N_11683,N_11631);
and U12839 (N_12839,N_11294,N_11470);
and U12840 (N_12840,N_12299,N_11929);
nand U12841 (N_12841,N_11419,N_11620);
or U12842 (N_12842,N_11495,N_11950);
or U12843 (N_12843,N_11287,N_11981);
nand U12844 (N_12844,N_12349,N_12054);
xor U12845 (N_12845,N_11560,N_12164);
and U12846 (N_12846,N_11977,N_11603);
or U12847 (N_12847,N_11371,N_11676);
nor U12848 (N_12848,N_11814,N_11871);
nand U12849 (N_12849,N_11373,N_11547);
and U12850 (N_12850,N_11272,N_11274);
nand U12851 (N_12851,N_12198,N_11375);
or U12852 (N_12852,N_12224,N_12388);
nand U12853 (N_12853,N_11489,N_12143);
nand U12854 (N_12854,N_11995,N_12081);
and U12855 (N_12855,N_12406,N_12345);
nand U12856 (N_12856,N_11708,N_11439);
nand U12857 (N_12857,N_12399,N_11757);
xnor U12858 (N_12858,N_11604,N_11584);
and U12859 (N_12859,N_11899,N_12250);
or U12860 (N_12860,N_11407,N_12109);
nor U12861 (N_12861,N_12385,N_12424);
or U12862 (N_12862,N_11680,N_11477);
or U12863 (N_12863,N_11479,N_12259);
nor U12864 (N_12864,N_11436,N_11779);
or U12865 (N_12865,N_11568,N_12209);
or U12866 (N_12866,N_11308,N_11937);
and U12867 (N_12867,N_11812,N_12429);
and U12868 (N_12868,N_11855,N_11410);
nor U12869 (N_12869,N_12135,N_11657);
and U12870 (N_12870,N_12084,N_12309);
xnor U12871 (N_12871,N_11404,N_11485);
or U12872 (N_12872,N_12130,N_11583);
or U12873 (N_12873,N_12191,N_12387);
and U12874 (N_12874,N_12402,N_11390);
nand U12875 (N_12875,N_12336,N_11942);
nor U12876 (N_12876,N_12149,N_11945);
xnor U12877 (N_12877,N_11494,N_11310);
or U12878 (N_12878,N_12285,N_12126);
nor U12879 (N_12879,N_12031,N_11706);
or U12880 (N_12880,N_11822,N_11717);
or U12881 (N_12881,N_12230,N_12245);
nand U12882 (N_12882,N_11506,N_11319);
nand U12883 (N_12883,N_11751,N_12390);
or U12884 (N_12884,N_12473,N_12447);
nor U12885 (N_12885,N_11588,N_11422);
and U12886 (N_12886,N_12068,N_11284);
nand U12887 (N_12887,N_12339,N_11660);
xnor U12888 (N_12888,N_11437,N_11970);
and U12889 (N_12889,N_12034,N_12343);
nor U12890 (N_12890,N_11268,N_12281);
and U12891 (N_12891,N_12137,N_12127);
nand U12892 (N_12892,N_12492,N_12457);
xnor U12893 (N_12893,N_11589,N_11989);
and U12894 (N_12894,N_11256,N_11448);
and U12895 (N_12895,N_11739,N_12148);
nor U12896 (N_12896,N_12270,N_11972);
nand U12897 (N_12897,N_11919,N_11810);
or U12898 (N_12898,N_12344,N_12153);
nor U12899 (N_12899,N_12418,N_11389);
nand U12900 (N_12900,N_11393,N_11260);
nor U12901 (N_12901,N_11858,N_12051);
nor U12902 (N_12902,N_11901,N_11303);
and U12903 (N_12903,N_12240,N_11565);
or U12904 (N_12904,N_11304,N_12468);
or U12905 (N_12905,N_11409,N_12197);
nand U12906 (N_12906,N_11839,N_11465);
xnor U12907 (N_12907,N_11576,N_11925);
xor U12908 (N_12908,N_11323,N_11619);
and U12909 (N_12909,N_12057,N_11613);
nand U12910 (N_12910,N_11710,N_11969);
and U12911 (N_12911,N_12028,N_11699);
xnor U12912 (N_12912,N_11647,N_12396);
or U12913 (N_12913,N_12410,N_11753);
and U12914 (N_12914,N_12351,N_11797);
or U12915 (N_12915,N_11512,N_11625);
nand U12916 (N_12916,N_11607,N_12376);
and U12917 (N_12917,N_11809,N_12419);
nor U12918 (N_12918,N_11850,N_12019);
nand U12919 (N_12919,N_11804,N_11394);
xor U12920 (N_12920,N_11354,N_11964);
or U12921 (N_12921,N_11447,N_12214);
and U12922 (N_12922,N_11556,N_11300);
and U12923 (N_12923,N_11689,N_11655);
and U12924 (N_12924,N_11523,N_11483);
nand U12925 (N_12925,N_11324,N_11342);
nand U12926 (N_12926,N_11499,N_11318);
and U12927 (N_12927,N_11333,N_11949);
nor U12928 (N_12928,N_12294,N_12438);
nand U12929 (N_12929,N_12269,N_12003);
or U12930 (N_12930,N_11255,N_12038);
or U12931 (N_12931,N_11364,N_12115);
nor U12932 (N_12932,N_11742,N_11748);
and U12933 (N_12933,N_11475,N_12091);
or U12934 (N_12934,N_11335,N_12132);
xnor U12935 (N_12935,N_11623,N_11355);
xnor U12936 (N_12936,N_11842,N_11760);
and U12937 (N_12937,N_12356,N_11442);
and U12938 (N_12938,N_12022,N_11591);
and U12939 (N_12939,N_12498,N_11551);
nor U12940 (N_12940,N_11703,N_12011);
nor U12941 (N_12941,N_11649,N_11920);
and U12942 (N_12942,N_12176,N_12158);
xor U12943 (N_12943,N_11397,N_11340);
nor U12944 (N_12944,N_12271,N_12218);
nor U12945 (N_12945,N_12304,N_12261);
nand U12946 (N_12946,N_11414,N_11686);
xor U12947 (N_12947,N_11671,N_11954);
xnor U12948 (N_12948,N_12053,N_12411);
or U12949 (N_12949,N_12237,N_11597);
or U12950 (N_12950,N_11885,N_12436);
nand U12951 (N_12951,N_11443,N_11856);
or U12952 (N_12952,N_12061,N_11534);
and U12953 (N_12953,N_12139,N_11951);
nor U12954 (N_12954,N_12075,N_11983);
xor U12955 (N_12955,N_12242,N_11490);
nand U12956 (N_12956,N_12205,N_11878);
or U12957 (N_12957,N_11847,N_11536);
and U12958 (N_12958,N_11361,N_12005);
nand U12959 (N_12959,N_12136,N_12188);
and U12960 (N_12960,N_12394,N_12082);
or U12961 (N_12961,N_11859,N_11382);
and U12962 (N_12962,N_11329,N_12227);
nor U12963 (N_12963,N_11434,N_12444);
nor U12964 (N_12964,N_12086,N_11957);
xor U12965 (N_12965,N_12182,N_11642);
xnor U12966 (N_12966,N_12367,N_11807);
and U12967 (N_12967,N_11743,N_11464);
nor U12968 (N_12968,N_12286,N_11273);
nand U12969 (N_12969,N_12446,N_12133);
xor U12970 (N_12970,N_11788,N_12175);
xor U12971 (N_12971,N_12482,N_11350);
and U12972 (N_12972,N_12340,N_12392);
xnor U12973 (N_12973,N_12372,N_11747);
xor U12974 (N_12974,N_11606,N_11292);
and U12975 (N_12975,N_11801,N_11943);
and U12976 (N_12976,N_11338,N_11321);
nor U12977 (N_12977,N_12389,N_11358);
and U12978 (N_12978,N_11362,N_12260);
xor U12979 (N_12979,N_11634,N_12248);
nand U12980 (N_12980,N_12154,N_12231);
and U12981 (N_12981,N_11728,N_12491);
and U12982 (N_12982,N_11488,N_12382);
and U12983 (N_12983,N_11562,N_11987);
xor U12984 (N_12984,N_11882,N_11493);
xor U12985 (N_12985,N_11864,N_11672);
xor U12986 (N_12986,N_12142,N_11391);
and U12987 (N_12987,N_11381,N_11823);
xor U12988 (N_12988,N_11996,N_11455);
xnor U12989 (N_12989,N_11994,N_12407);
or U12990 (N_12990,N_12370,N_12024);
nor U12991 (N_12991,N_12318,N_11820);
nand U12992 (N_12992,N_12173,N_12080);
nand U12993 (N_12993,N_11387,N_11635);
nand U12994 (N_12994,N_12330,N_11559);
or U12995 (N_12995,N_12190,N_11798);
xor U12996 (N_12996,N_11679,N_12310);
xnor U12997 (N_12997,N_12026,N_11714);
nand U12998 (N_12998,N_12437,N_12455);
and U12999 (N_12999,N_11854,N_11650);
nand U13000 (N_13000,N_11912,N_12421);
and U13001 (N_13001,N_11484,N_12023);
xor U13002 (N_13002,N_11697,N_12277);
xor U13003 (N_13003,N_12045,N_11299);
nor U13004 (N_13004,N_12183,N_12088);
xor U13005 (N_13005,N_12171,N_12097);
and U13006 (N_13006,N_12485,N_11474);
nor U13007 (N_13007,N_11445,N_12189);
nand U13008 (N_13008,N_11564,N_11791);
nor U13009 (N_13009,N_11900,N_11762);
and U13010 (N_13010,N_11406,N_11385);
nand U13011 (N_13011,N_12263,N_11601);
nand U13012 (N_13012,N_11639,N_12463);
and U13013 (N_13013,N_11874,N_12070);
and U13014 (N_13014,N_12375,N_11792);
and U13015 (N_13015,N_11456,N_11750);
or U13016 (N_13016,N_11780,N_11541);
and U13017 (N_13017,N_12162,N_12426);
and U13018 (N_13018,N_12486,N_11451);
nor U13019 (N_13019,N_11643,N_12381);
xnor U13020 (N_13020,N_11931,N_11325);
nor U13021 (N_13021,N_11658,N_12404);
or U13022 (N_13022,N_11715,N_11377);
nor U13023 (N_13023,N_11863,N_12460);
xnor U13024 (N_13024,N_12431,N_11922);
or U13025 (N_13025,N_11938,N_11339);
and U13026 (N_13026,N_12102,N_12216);
and U13027 (N_13027,N_11661,N_11524);
xor U13028 (N_13028,N_11476,N_12203);
xnor U13029 (N_13029,N_11473,N_11463);
nor U13030 (N_13030,N_11693,N_11504);
nand U13031 (N_13031,N_12006,N_11412);
nand U13032 (N_13032,N_11383,N_12360);
nor U13033 (N_13033,N_11366,N_11733);
xnor U13034 (N_13034,N_12347,N_12239);
and U13035 (N_13035,N_11857,N_11766);
xor U13036 (N_13036,N_11520,N_11538);
nand U13037 (N_13037,N_12425,N_12145);
and U13038 (N_13038,N_11544,N_11611);
nor U13039 (N_13039,N_12379,N_11879);
nand U13040 (N_13040,N_11828,N_11592);
and U13041 (N_13041,N_12243,N_12272);
nor U13042 (N_13042,N_11841,N_12464);
nand U13043 (N_13043,N_11723,N_11511);
or U13044 (N_13044,N_11722,N_11806);
xnor U13045 (N_13045,N_11890,N_12196);
and U13046 (N_13046,N_12416,N_11610);
xor U13047 (N_13047,N_11624,N_11312);
nor U13048 (N_13048,N_11574,N_11337);
and U13049 (N_13049,N_12377,N_11844);
nor U13050 (N_13050,N_11531,N_11492);
xor U13051 (N_13051,N_11618,N_11896);
or U13052 (N_13052,N_11816,N_11519);
nor U13053 (N_13053,N_11326,N_12165);
and U13054 (N_13054,N_12400,N_11527);
xnor U13055 (N_13055,N_11309,N_12364);
nor U13056 (N_13056,N_11638,N_12256);
or U13057 (N_13057,N_11652,N_12440);
and U13058 (N_13058,N_11332,N_12280);
nand U13059 (N_13059,N_12301,N_11991);
and U13060 (N_13060,N_11546,N_12172);
or U13061 (N_13061,N_12268,N_11637);
or U13062 (N_13062,N_12274,N_11263);
nor U13063 (N_13063,N_12211,N_11563);
nor U13064 (N_13064,N_11425,N_11725);
xor U13065 (N_13065,N_12369,N_11648);
nor U13066 (N_13066,N_11471,N_12029);
xor U13067 (N_13067,N_12296,N_12393);
nor U13068 (N_13068,N_12433,N_11778);
and U13069 (N_13069,N_12161,N_11745);
nand U13070 (N_13070,N_11892,N_11388);
xor U13071 (N_13071,N_12495,N_11432);
or U13072 (N_13072,N_11978,N_11365);
xor U13073 (N_13073,N_12452,N_12324);
nor U13074 (N_13074,N_11789,N_12219);
and U13075 (N_13075,N_11764,N_11838);
xnor U13076 (N_13076,N_11880,N_11718);
or U13077 (N_13077,N_11955,N_11297);
nand U13078 (N_13078,N_12328,N_11761);
xnor U13079 (N_13079,N_11793,N_11845);
nor U13080 (N_13080,N_11852,N_11883);
nor U13081 (N_13081,N_11730,N_11415);
nand U13082 (N_13082,N_12120,N_12331);
and U13083 (N_13083,N_11811,N_11521);
nor U13084 (N_13084,N_11678,N_12470);
nand U13085 (N_13085,N_11413,N_12094);
nor U13086 (N_13086,N_11628,N_11454);
xor U13087 (N_13087,N_12073,N_12241);
nand U13088 (N_13088,N_11348,N_11944);
nand U13089 (N_13089,N_11997,N_12341);
nor U13090 (N_13090,N_12414,N_11408);
or U13091 (N_13091,N_11749,N_12453);
nand U13092 (N_13092,N_11934,N_12475);
xnor U13093 (N_13093,N_12466,N_11973);
xnor U13094 (N_13094,N_11968,N_12417);
and U13095 (N_13095,N_12108,N_11771);
or U13096 (N_13096,N_11418,N_12015);
nand U13097 (N_13097,N_11702,N_11586);
nor U13098 (N_13098,N_11840,N_11369);
nand U13099 (N_13099,N_11528,N_11558);
xor U13100 (N_13100,N_11264,N_11720);
nor U13101 (N_13101,N_12313,N_11935);
nand U13102 (N_13102,N_11904,N_11933);
or U13103 (N_13103,N_11587,N_12027);
and U13104 (N_13104,N_11752,N_11831);
and U13105 (N_13105,N_11289,N_12247);
nand U13106 (N_13106,N_12462,N_11577);
xnor U13107 (N_13107,N_12244,N_12077);
nor U13108 (N_13108,N_12092,N_12290);
xor U13109 (N_13109,N_11581,N_11656);
nor U13110 (N_13110,N_11579,N_12332);
nand U13111 (N_13111,N_11990,N_11372);
xor U13112 (N_13112,N_11897,N_11674);
xnor U13113 (N_13113,N_11291,N_11962);
nand U13114 (N_13114,N_11756,N_11687);
and U13115 (N_13115,N_11802,N_11612);
or U13116 (N_13116,N_11608,N_12210);
and U13117 (N_13117,N_12423,N_11469);
xnor U13118 (N_13118,N_11428,N_11911);
and U13119 (N_13119,N_12398,N_11803);
xor U13120 (N_13120,N_11651,N_11691);
xnor U13121 (N_13121,N_11903,N_11617);
nor U13122 (N_13122,N_11542,N_12087);
and U13123 (N_13123,N_12032,N_12408);
xnor U13124 (N_13124,N_11734,N_12484);
nand U13125 (N_13125,N_11267,N_11510);
and U13126 (N_13126,N_11333,N_12218);
and U13127 (N_13127,N_11699,N_11886);
or U13128 (N_13128,N_12002,N_11794);
nand U13129 (N_13129,N_11419,N_11879);
or U13130 (N_13130,N_12239,N_12371);
and U13131 (N_13131,N_12248,N_11263);
and U13132 (N_13132,N_11868,N_11321);
and U13133 (N_13133,N_11966,N_11327);
nand U13134 (N_13134,N_12352,N_11392);
nand U13135 (N_13135,N_11856,N_11466);
nand U13136 (N_13136,N_12414,N_11445);
and U13137 (N_13137,N_12330,N_11764);
nor U13138 (N_13138,N_11345,N_11599);
and U13139 (N_13139,N_11680,N_11750);
nand U13140 (N_13140,N_12184,N_11793);
xor U13141 (N_13141,N_11664,N_12084);
nand U13142 (N_13142,N_11689,N_11984);
xnor U13143 (N_13143,N_12179,N_11314);
nor U13144 (N_13144,N_11371,N_11348);
nor U13145 (N_13145,N_12474,N_12052);
and U13146 (N_13146,N_11354,N_12483);
or U13147 (N_13147,N_11326,N_11627);
and U13148 (N_13148,N_12053,N_11490);
or U13149 (N_13149,N_12073,N_12478);
nand U13150 (N_13150,N_12207,N_11648);
xor U13151 (N_13151,N_12441,N_12337);
nand U13152 (N_13152,N_11363,N_11345);
nor U13153 (N_13153,N_11800,N_11852);
nand U13154 (N_13154,N_11629,N_11290);
xnor U13155 (N_13155,N_11985,N_11554);
nor U13156 (N_13156,N_11835,N_12473);
and U13157 (N_13157,N_11320,N_11322);
xor U13158 (N_13158,N_11842,N_12344);
nor U13159 (N_13159,N_12209,N_11794);
and U13160 (N_13160,N_11261,N_11605);
nor U13161 (N_13161,N_11358,N_11877);
xor U13162 (N_13162,N_12006,N_11736);
xnor U13163 (N_13163,N_11699,N_11770);
and U13164 (N_13164,N_11761,N_11455);
and U13165 (N_13165,N_11798,N_11371);
and U13166 (N_13166,N_11494,N_11716);
or U13167 (N_13167,N_11824,N_11880);
and U13168 (N_13168,N_12344,N_12219);
xor U13169 (N_13169,N_11961,N_12084);
nor U13170 (N_13170,N_11699,N_11267);
and U13171 (N_13171,N_11341,N_12135);
or U13172 (N_13172,N_11801,N_12118);
xor U13173 (N_13173,N_12171,N_11947);
nand U13174 (N_13174,N_11686,N_11731);
or U13175 (N_13175,N_11937,N_12468);
nor U13176 (N_13176,N_11712,N_11921);
or U13177 (N_13177,N_12266,N_12485);
nor U13178 (N_13178,N_12360,N_11748);
or U13179 (N_13179,N_12475,N_12138);
nor U13180 (N_13180,N_12431,N_11480);
xor U13181 (N_13181,N_11336,N_11985);
nor U13182 (N_13182,N_12005,N_11567);
xor U13183 (N_13183,N_12414,N_11619);
xnor U13184 (N_13184,N_11941,N_11798);
or U13185 (N_13185,N_11528,N_11582);
and U13186 (N_13186,N_12075,N_11345);
nor U13187 (N_13187,N_11746,N_12030);
or U13188 (N_13188,N_11730,N_11547);
or U13189 (N_13189,N_11364,N_12454);
xnor U13190 (N_13190,N_11398,N_11973);
or U13191 (N_13191,N_11416,N_12334);
xor U13192 (N_13192,N_11452,N_12004);
nor U13193 (N_13193,N_12248,N_12224);
nand U13194 (N_13194,N_11732,N_12326);
nor U13195 (N_13195,N_12282,N_12440);
nor U13196 (N_13196,N_12361,N_12022);
and U13197 (N_13197,N_11370,N_12344);
or U13198 (N_13198,N_12109,N_11483);
nor U13199 (N_13199,N_12445,N_12336);
nor U13200 (N_13200,N_11280,N_12451);
nand U13201 (N_13201,N_12434,N_11987);
nor U13202 (N_13202,N_11286,N_11319);
and U13203 (N_13203,N_12029,N_11530);
xnor U13204 (N_13204,N_12434,N_12229);
xnor U13205 (N_13205,N_12022,N_12299);
nor U13206 (N_13206,N_12063,N_11788);
or U13207 (N_13207,N_11436,N_12063);
xor U13208 (N_13208,N_12473,N_12072);
or U13209 (N_13209,N_12011,N_12057);
or U13210 (N_13210,N_12308,N_11851);
nand U13211 (N_13211,N_12176,N_11279);
or U13212 (N_13212,N_12122,N_11917);
nand U13213 (N_13213,N_11789,N_11880);
or U13214 (N_13214,N_11910,N_11492);
or U13215 (N_13215,N_12248,N_11875);
nor U13216 (N_13216,N_11343,N_11877);
or U13217 (N_13217,N_11321,N_11684);
xor U13218 (N_13218,N_12073,N_12321);
xnor U13219 (N_13219,N_12176,N_12222);
xor U13220 (N_13220,N_12038,N_11373);
xnor U13221 (N_13221,N_12045,N_11862);
xnor U13222 (N_13222,N_11673,N_11676);
and U13223 (N_13223,N_11551,N_12423);
or U13224 (N_13224,N_12408,N_11459);
and U13225 (N_13225,N_11692,N_11998);
xnor U13226 (N_13226,N_11629,N_11798);
and U13227 (N_13227,N_11529,N_12496);
nand U13228 (N_13228,N_11883,N_12402);
nor U13229 (N_13229,N_12427,N_11325);
nor U13230 (N_13230,N_12044,N_11371);
and U13231 (N_13231,N_11722,N_12437);
nor U13232 (N_13232,N_11747,N_11742);
xnor U13233 (N_13233,N_12357,N_12376);
nor U13234 (N_13234,N_12444,N_11876);
nor U13235 (N_13235,N_12014,N_11852);
and U13236 (N_13236,N_11539,N_12369);
nand U13237 (N_13237,N_12231,N_11461);
or U13238 (N_13238,N_11505,N_11419);
or U13239 (N_13239,N_11475,N_12476);
nand U13240 (N_13240,N_11257,N_12057);
nand U13241 (N_13241,N_12209,N_11677);
xor U13242 (N_13242,N_11913,N_11596);
xor U13243 (N_13243,N_11874,N_12371);
nand U13244 (N_13244,N_12003,N_12129);
nand U13245 (N_13245,N_12118,N_11479);
nor U13246 (N_13246,N_11499,N_12240);
nor U13247 (N_13247,N_12383,N_11690);
or U13248 (N_13248,N_12363,N_12399);
nor U13249 (N_13249,N_11292,N_11302);
xnor U13250 (N_13250,N_12354,N_11361);
or U13251 (N_13251,N_12144,N_12254);
nor U13252 (N_13252,N_11388,N_11493);
and U13253 (N_13253,N_11570,N_11632);
nor U13254 (N_13254,N_12030,N_11984);
xor U13255 (N_13255,N_11427,N_12351);
xnor U13256 (N_13256,N_11291,N_11901);
and U13257 (N_13257,N_12318,N_11660);
nand U13258 (N_13258,N_11400,N_11913);
and U13259 (N_13259,N_11782,N_12464);
nor U13260 (N_13260,N_12414,N_11890);
nand U13261 (N_13261,N_12357,N_11421);
nor U13262 (N_13262,N_11545,N_12009);
or U13263 (N_13263,N_11726,N_11575);
nand U13264 (N_13264,N_12066,N_12348);
or U13265 (N_13265,N_12134,N_11495);
and U13266 (N_13266,N_11459,N_11571);
xor U13267 (N_13267,N_11534,N_11405);
or U13268 (N_13268,N_12238,N_11540);
or U13269 (N_13269,N_11823,N_12338);
and U13270 (N_13270,N_12296,N_12242);
or U13271 (N_13271,N_11373,N_11532);
xnor U13272 (N_13272,N_11667,N_11309);
or U13273 (N_13273,N_11362,N_11908);
or U13274 (N_13274,N_11601,N_11508);
xnor U13275 (N_13275,N_11565,N_12428);
nor U13276 (N_13276,N_12119,N_11360);
nand U13277 (N_13277,N_12163,N_12429);
nand U13278 (N_13278,N_12155,N_12388);
or U13279 (N_13279,N_11698,N_11729);
nand U13280 (N_13280,N_11761,N_12276);
and U13281 (N_13281,N_11765,N_11578);
and U13282 (N_13282,N_12320,N_12070);
or U13283 (N_13283,N_12389,N_11902);
xor U13284 (N_13284,N_12481,N_11890);
xnor U13285 (N_13285,N_11268,N_11798);
nor U13286 (N_13286,N_12138,N_11455);
nor U13287 (N_13287,N_11672,N_12348);
and U13288 (N_13288,N_11853,N_11733);
or U13289 (N_13289,N_11796,N_11538);
and U13290 (N_13290,N_11610,N_12141);
or U13291 (N_13291,N_11387,N_12351);
nand U13292 (N_13292,N_11285,N_12118);
or U13293 (N_13293,N_11793,N_12467);
xor U13294 (N_13294,N_11584,N_11883);
or U13295 (N_13295,N_11375,N_12378);
or U13296 (N_13296,N_11326,N_11563);
or U13297 (N_13297,N_12026,N_12261);
nand U13298 (N_13298,N_12391,N_11411);
xor U13299 (N_13299,N_12401,N_12206);
nand U13300 (N_13300,N_12373,N_11778);
xnor U13301 (N_13301,N_11758,N_11267);
nand U13302 (N_13302,N_11357,N_11287);
nand U13303 (N_13303,N_11421,N_12255);
nand U13304 (N_13304,N_12139,N_11366);
and U13305 (N_13305,N_11377,N_11650);
xnor U13306 (N_13306,N_12287,N_12276);
or U13307 (N_13307,N_11653,N_12206);
xor U13308 (N_13308,N_11928,N_11940);
or U13309 (N_13309,N_11301,N_12180);
and U13310 (N_13310,N_12410,N_11989);
nand U13311 (N_13311,N_11620,N_11951);
or U13312 (N_13312,N_11293,N_11591);
nor U13313 (N_13313,N_11844,N_11429);
xor U13314 (N_13314,N_11391,N_12472);
and U13315 (N_13315,N_11979,N_11998);
nand U13316 (N_13316,N_11556,N_11610);
nor U13317 (N_13317,N_12156,N_12324);
or U13318 (N_13318,N_11870,N_11762);
nor U13319 (N_13319,N_12481,N_11647);
or U13320 (N_13320,N_11443,N_11464);
and U13321 (N_13321,N_12374,N_11786);
or U13322 (N_13322,N_12442,N_12456);
and U13323 (N_13323,N_11712,N_11663);
nand U13324 (N_13324,N_11989,N_11862);
and U13325 (N_13325,N_11502,N_12276);
or U13326 (N_13326,N_12270,N_11621);
nand U13327 (N_13327,N_12167,N_11333);
or U13328 (N_13328,N_12454,N_12365);
or U13329 (N_13329,N_11918,N_11904);
nand U13330 (N_13330,N_11845,N_12016);
nor U13331 (N_13331,N_12458,N_11887);
and U13332 (N_13332,N_12167,N_11886);
and U13333 (N_13333,N_12424,N_11641);
or U13334 (N_13334,N_11647,N_12351);
or U13335 (N_13335,N_11264,N_11585);
nand U13336 (N_13336,N_12173,N_11516);
xor U13337 (N_13337,N_12150,N_11507);
xnor U13338 (N_13338,N_11460,N_12083);
or U13339 (N_13339,N_12275,N_12013);
nand U13340 (N_13340,N_12304,N_11697);
xor U13341 (N_13341,N_12266,N_12475);
nor U13342 (N_13342,N_12366,N_11587);
or U13343 (N_13343,N_11550,N_11368);
or U13344 (N_13344,N_12373,N_11343);
nor U13345 (N_13345,N_12401,N_12334);
xor U13346 (N_13346,N_12305,N_12187);
nand U13347 (N_13347,N_11951,N_11725);
nand U13348 (N_13348,N_11819,N_11581);
nand U13349 (N_13349,N_12246,N_12269);
or U13350 (N_13350,N_11720,N_11446);
xnor U13351 (N_13351,N_11826,N_11398);
and U13352 (N_13352,N_11532,N_12462);
and U13353 (N_13353,N_11336,N_12211);
nand U13354 (N_13354,N_11721,N_11596);
and U13355 (N_13355,N_12071,N_12314);
xnor U13356 (N_13356,N_11371,N_11411);
and U13357 (N_13357,N_11676,N_11752);
and U13358 (N_13358,N_11538,N_12251);
nor U13359 (N_13359,N_12145,N_12418);
or U13360 (N_13360,N_11773,N_11616);
xnor U13361 (N_13361,N_11469,N_11378);
or U13362 (N_13362,N_11944,N_11796);
or U13363 (N_13363,N_11341,N_11863);
nand U13364 (N_13364,N_11286,N_11276);
nand U13365 (N_13365,N_12492,N_12292);
xnor U13366 (N_13366,N_11615,N_12294);
and U13367 (N_13367,N_12447,N_12260);
nor U13368 (N_13368,N_11317,N_11471);
xnor U13369 (N_13369,N_12090,N_11680);
nand U13370 (N_13370,N_11759,N_11772);
xor U13371 (N_13371,N_11254,N_11739);
xor U13372 (N_13372,N_11571,N_12313);
nor U13373 (N_13373,N_12489,N_11767);
nor U13374 (N_13374,N_11446,N_12369);
or U13375 (N_13375,N_11553,N_11942);
and U13376 (N_13376,N_11790,N_11906);
or U13377 (N_13377,N_11282,N_12408);
or U13378 (N_13378,N_12063,N_12004);
and U13379 (N_13379,N_11924,N_12100);
or U13380 (N_13380,N_12172,N_11875);
or U13381 (N_13381,N_11841,N_12002);
nor U13382 (N_13382,N_11675,N_11656);
or U13383 (N_13383,N_11407,N_11884);
nand U13384 (N_13384,N_11765,N_11253);
xnor U13385 (N_13385,N_11713,N_11306);
or U13386 (N_13386,N_11628,N_11642);
xor U13387 (N_13387,N_12126,N_11402);
and U13388 (N_13388,N_11760,N_12484);
xor U13389 (N_13389,N_11502,N_12038);
xnor U13390 (N_13390,N_12276,N_12076);
nand U13391 (N_13391,N_12468,N_12029);
nor U13392 (N_13392,N_12423,N_11738);
and U13393 (N_13393,N_11466,N_12227);
or U13394 (N_13394,N_11684,N_11958);
and U13395 (N_13395,N_11525,N_11700);
nand U13396 (N_13396,N_11564,N_11768);
nor U13397 (N_13397,N_11967,N_11294);
nand U13398 (N_13398,N_11600,N_12119);
nor U13399 (N_13399,N_12262,N_11818);
or U13400 (N_13400,N_11842,N_11877);
nor U13401 (N_13401,N_12031,N_12174);
and U13402 (N_13402,N_11466,N_12269);
or U13403 (N_13403,N_12049,N_11991);
nor U13404 (N_13404,N_11835,N_11504);
and U13405 (N_13405,N_11716,N_11813);
xor U13406 (N_13406,N_11305,N_12435);
xor U13407 (N_13407,N_11567,N_11528);
nor U13408 (N_13408,N_12129,N_11351);
nor U13409 (N_13409,N_12422,N_12182);
and U13410 (N_13410,N_12195,N_12221);
and U13411 (N_13411,N_11700,N_11655);
and U13412 (N_13412,N_11457,N_12237);
xor U13413 (N_13413,N_11565,N_12096);
or U13414 (N_13414,N_12070,N_11988);
or U13415 (N_13415,N_12097,N_12053);
xor U13416 (N_13416,N_12090,N_11708);
nor U13417 (N_13417,N_11918,N_11452);
nand U13418 (N_13418,N_11968,N_12210);
nand U13419 (N_13419,N_12164,N_11701);
xnor U13420 (N_13420,N_12364,N_11652);
or U13421 (N_13421,N_11835,N_11552);
or U13422 (N_13422,N_12432,N_11442);
or U13423 (N_13423,N_11770,N_12052);
xor U13424 (N_13424,N_11274,N_11809);
nor U13425 (N_13425,N_11896,N_11476);
and U13426 (N_13426,N_11628,N_12040);
and U13427 (N_13427,N_11983,N_12244);
or U13428 (N_13428,N_11803,N_12274);
nand U13429 (N_13429,N_12413,N_11560);
xnor U13430 (N_13430,N_12108,N_11792);
and U13431 (N_13431,N_12397,N_11973);
and U13432 (N_13432,N_12111,N_11391);
or U13433 (N_13433,N_11636,N_12209);
and U13434 (N_13434,N_12378,N_12389);
or U13435 (N_13435,N_11732,N_11427);
nor U13436 (N_13436,N_11826,N_12475);
xor U13437 (N_13437,N_11555,N_12323);
or U13438 (N_13438,N_11548,N_11606);
or U13439 (N_13439,N_12066,N_11924);
nand U13440 (N_13440,N_11491,N_11742);
nor U13441 (N_13441,N_11732,N_11439);
nor U13442 (N_13442,N_12274,N_12167);
nand U13443 (N_13443,N_12059,N_12280);
nor U13444 (N_13444,N_12424,N_11305);
and U13445 (N_13445,N_12349,N_12070);
and U13446 (N_13446,N_11519,N_11865);
xor U13447 (N_13447,N_12212,N_11995);
xor U13448 (N_13448,N_11867,N_12428);
nor U13449 (N_13449,N_11962,N_12161);
or U13450 (N_13450,N_11291,N_11947);
xor U13451 (N_13451,N_12328,N_12010);
nand U13452 (N_13452,N_11488,N_11268);
xor U13453 (N_13453,N_11864,N_12086);
and U13454 (N_13454,N_11749,N_11739);
and U13455 (N_13455,N_12364,N_12078);
nor U13456 (N_13456,N_12136,N_11604);
nor U13457 (N_13457,N_11598,N_12226);
and U13458 (N_13458,N_12012,N_11872);
and U13459 (N_13459,N_12066,N_11816);
nor U13460 (N_13460,N_11784,N_11880);
and U13461 (N_13461,N_12216,N_12185);
xor U13462 (N_13462,N_11309,N_12208);
xor U13463 (N_13463,N_11482,N_12147);
xnor U13464 (N_13464,N_11584,N_12079);
nand U13465 (N_13465,N_11586,N_12299);
nor U13466 (N_13466,N_11392,N_11548);
xor U13467 (N_13467,N_12147,N_12356);
nand U13468 (N_13468,N_11670,N_11510);
nor U13469 (N_13469,N_11635,N_11319);
nand U13470 (N_13470,N_12200,N_12214);
or U13471 (N_13471,N_11567,N_11394);
or U13472 (N_13472,N_12360,N_11818);
nand U13473 (N_13473,N_12348,N_12179);
and U13474 (N_13474,N_12397,N_11979);
or U13475 (N_13475,N_11685,N_11383);
xor U13476 (N_13476,N_12006,N_12276);
xnor U13477 (N_13477,N_11917,N_11321);
nand U13478 (N_13478,N_12054,N_12146);
xor U13479 (N_13479,N_11933,N_12240);
and U13480 (N_13480,N_12370,N_12190);
or U13481 (N_13481,N_12324,N_11370);
nand U13482 (N_13482,N_12300,N_11974);
xnor U13483 (N_13483,N_12422,N_12261);
xnor U13484 (N_13484,N_11285,N_11261);
nand U13485 (N_13485,N_11372,N_12304);
xor U13486 (N_13486,N_11681,N_11864);
nor U13487 (N_13487,N_11284,N_11604);
nor U13488 (N_13488,N_11945,N_11889);
or U13489 (N_13489,N_11787,N_11593);
xor U13490 (N_13490,N_11656,N_11622);
xnor U13491 (N_13491,N_12051,N_12469);
nor U13492 (N_13492,N_11711,N_12193);
xnor U13493 (N_13493,N_11788,N_11527);
nor U13494 (N_13494,N_12178,N_11287);
and U13495 (N_13495,N_12440,N_12478);
xnor U13496 (N_13496,N_12130,N_11375);
xor U13497 (N_13497,N_12467,N_11552);
nand U13498 (N_13498,N_12173,N_12304);
and U13499 (N_13499,N_12060,N_12051);
and U13500 (N_13500,N_12104,N_11996);
or U13501 (N_13501,N_12141,N_11799);
and U13502 (N_13502,N_11722,N_11757);
xor U13503 (N_13503,N_11994,N_11387);
nor U13504 (N_13504,N_12438,N_12036);
or U13505 (N_13505,N_11681,N_12442);
nor U13506 (N_13506,N_11386,N_12362);
or U13507 (N_13507,N_12008,N_12110);
and U13508 (N_13508,N_12206,N_11351);
xnor U13509 (N_13509,N_11517,N_12309);
nand U13510 (N_13510,N_12170,N_12369);
nor U13511 (N_13511,N_12465,N_12337);
xnor U13512 (N_13512,N_11886,N_11530);
xor U13513 (N_13513,N_11915,N_12170);
or U13514 (N_13514,N_12078,N_11370);
nand U13515 (N_13515,N_11419,N_12088);
xor U13516 (N_13516,N_11323,N_12202);
nand U13517 (N_13517,N_11983,N_11701);
xor U13518 (N_13518,N_11567,N_11753);
nand U13519 (N_13519,N_12379,N_12417);
nand U13520 (N_13520,N_11935,N_12256);
nor U13521 (N_13521,N_12447,N_11622);
xor U13522 (N_13522,N_12368,N_11593);
xor U13523 (N_13523,N_11512,N_12330);
nand U13524 (N_13524,N_12080,N_12294);
xor U13525 (N_13525,N_12461,N_11635);
nor U13526 (N_13526,N_11602,N_11668);
nor U13527 (N_13527,N_11879,N_11330);
or U13528 (N_13528,N_12467,N_11981);
and U13529 (N_13529,N_11336,N_12471);
or U13530 (N_13530,N_12035,N_12399);
or U13531 (N_13531,N_11649,N_11451);
nand U13532 (N_13532,N_12042,N_11728);
or U13533 (N_13533,N_11324,N_11954);
nor U13534 (N_13534,N_12309,N_11994);
nand U13535 (N_13535,N_11584,N_11502);
nor U13536 (N_13536,N_11725,N_11534);
xnor U13537 (N_13537,N_11486,N_11395);
or U13538 (N_13538,N_12451,N_12078);
or U13539 (N_13539,N_11460,N_11902);
nor U13540 (N_13540,N_12084,N_11871);
nand U13541 (N_13541,N_11455,N_11404);
nand U13542 (N_13542,N_12336,N_11278);
nand U13543 (N_13543,N_12269,N_11406);
nand U13544 (N_13544,N_11759,N_11941);
and U13545 (N_13545,N_11992,N_12197);
nor U13546 (N_13546,N_11759,N_12259);
nand U13547 (N_13547,N_11879,N_11427);
xor U13548 (N_13548,N_11856,N_12491);
or U13549 (N_13549,N_11925,N_12268);
nand U13550 (N_13550,N_11374,N_12416);
or U13551 (N_13551,N_11463,N_11668);
nor U13552 (N_13552,N_11375,N_11466);
and U13553 (N_13553,N_11988,N_11581);
nor U13554 (N_13554,N_11702,N_12465);
xor U13555 (N_13555,N_11304,N_11865);
or U13556 (N_13556,N_12294,N_12379);
nand U13557 (N_13557,N_11338,N_12011);
nor U13558 (N_13558,N_11535,N_12440);
or U13559 (N_13559,N_12443,N_11299);
or U13560 (N_13560,N_12219,N_11676);
and U13561 (N_13561,N_11866,N_11675);
and U13562 (N_13562,N_12497,N_11873);
xor U13563 (N_13563,N_11742,N_12124);
nor U13564 (N_13564,N_12100,N_12002);
nor U13565 (N_13565,N_12058,N_11497);
and U13566 (N_13566,N_11579,N_12217);
or U13567 (N_13567,N_11509,N_11430);
and U13568 (N_13568,N_11604,N_11663);
nand U13569 (N_13569,N_11282,N_12167);
nor U13570 (N_13570,N_11812,N_11713);
nor U13571 (N_13571,N_12436,N_11812);
or U13572 (N_13572,N_12459,N_11593);
xor U13573 (N_13573,N_11296,N_11753);
nor U13574 (N_13574,N_11890,N_11948);
xnor U13575 (N_13575,N_12305,N_11348);
xor U13576 (N_13576,N_11453,N_12043);
nor U13577 (N_13577,N_12088,N_12485);
or U13578 (N_13578,N_12468,N_12424);
and U13579 (N_13579,N_11810,N_12126);
nor U13580 (N_13580,N_11553,N_12479);
or U13581 (N_13581,N_11740,N_11734);
or U13582 (N_13582,N_11602,N_12384);
nor U13583 (N_13583,N_12138,N_11272);
nor U13584 (N_13584,N_12101,N_11670);
and U13585 (N_13585,N_12382,N_12080);
nor U13586 (N_13586,N_12177,N_11968);
nand U13587 (N_13587,N_12003,N_11809);
or U13588 (N_13588,N_11906,N_11940);
or U13589 (N_13589,N_12013,N_11488);
nor U13590 (N_13590,N_12236,N_12459);
nor U13591 (N_13591,N_12084,N_11645);
xor U13592 (N_13592,N_12383,N_12060);
xnor U13593 (N_13593,N_12117,N_11959);
and U13594 (N_13594,N_11615,N_12134);
nand U13595 (N_13595,N_11957,N_11800);
nand U13596 (N_13596,N_12227,N_11805);
nor U13597 (N_13597,N_11596,N_11648);
nand U13598 (N_13598,N_11845,N_11645);
xnor U13599 (N_13599,N_11427,N_11649);
and U13600 (N_13600,N_11870,N_11723);
nor U13601 (N_13601,N_12171,N_11790);
nand U13602 (N_13602,N_12284,N_11511);
nor U13603 (N_13603,N_11954,N_11850);
nor U13604 (N_13604,N_12354,N_11605);
and U13605 (N_13605,N_11856,N_11705);
and U13606 (N_13606,N_11847,N_12178);
and U13607 (N_13607,N_11854,N_12083);
nor U13608 (N_13608,N_11582,N_11458);
and U13609 (N_13609,N_12193,N_12411);
xor U13610 (N_13610,N_11299,N_11414);
xor U13611 (N_13611,N_12109,N_11729);
xor U13612 (N_13612,N_12085,N_11671);
and U13613 (N_13613,N_11725,N_12169);
or U13614 (N_13614,N_12477,N_11890);
and U13615 (N_13615,N_11494,N_11625);
or U13616 (N_13616,N_11861,N_12271);
or U13617 (N_13617,N_11926,N_11381);
nor U13618 (N_13618,N_12238,N_11784);
and U13619 (N_13619,N_11582,N_11423);
or U13620 (N_13620,N_11912,N_11398);
nand U13621 (N_13621,N_11737,N_11774);
nor U13622 (N_13622,N_11306,N_11843);
nor U13623 (N_13623,N_11600,N_11916);
nor U13624 (N_13624,N_12148,N_11367);
or U13625 (N_13625,N_12086,N_11652);
xnor U13626 (N_13626,N_11480,N_12291);
nor U13627 (N_13627,N_11335,N_11741);
xnor U13628 (N_13628,N_11807,N_11500);
xnor U13629 (N_13629,N_11709,N_11937);
nand U13630 (N_13630,N_11870,N_11703);
or U13631 (N_13631,N_12421,N_11945);
xnor U13632 (N_13632,N_11343,N_12035);
xor U13633 (N_13633,N_12242,N_11789);
and U13634 (N_13634,N_11912,N_11487);
and U13635 (N_13635,N_11462,N_12098);
xnor U13636 (N_13636,N_11923,N_12280);
nor U13637 (N_13637,N_12196,N_11557);
and U13638 (N_13638,N_12280,N_11971);
and U13639 (N_13639,N_11683,N_12285);
nor U13640 (N_13640,N_11717,N_11253);
and U13641 (N_13641,N_11836,N_12194);
or U13642 (N_13642,N_11505,N_12021);
nand U13643 (N_13643,N_12232,N_11726);
and U13644 (N_13644,N_11920,N_11463);
and U13645 (N_13645,N_11570,N_12292);
or U13646 (N_13646,N_12461,N_12473);
nand U13647 (N_13647,N_11588,N_12471);
or U13648 (N_13648,N_11877,N_12311);
or U13649 (N_13649,N_11895,N_11296);
nand U13650 (N_13650,N_12374,N_11761);
and U13651 (N_13651,N_11663,N_12402);
nor U13652 (N_13652,N_11882,N_11746);
nor U13653 (N_13653,N_12027,N_11360);
nor U13654 (N_13654,N_11994,N_12007);
and U13655 (N_13655,N_11452,N_11852);
and U13656 (N_13656,N_12447,N_11839);
nand U13657 (N_13657,N_11332,N_12206);
nor U13658 (N_13658,N_12171,N_12128);
and U13659 (N_13659,N_11678,N_11394);
or U13660 (N_13660,N_11518,N_11790);
nand U13661 (N_13661,N_11418,N_12499);
nand U13662 (N_13662,N_12142,N_12448);
nor U13663 (N_13663,N_12430,N_11908);
and U13664 (N_13664,N_11539,N_12126);
xor U13665 (N_13665,N_11641,N_11904);
nand U13666 (N_13666,N_11598,N_11568);
nand U13667 (N_13667,N_11377,N_12459);
xor U13668 (N_13668,N_11318,N_11715);
or U13669 (N_13669,N_11993,N_12216);
nor U13670 (N_13670,N_12105,N_12491);
or U13671 (N_13671,N_12071,N_12315);
nand U13672 (N_13672,N_12254,N_11440);
or U13673 (N_13673,N_11544,N_11956);
nor U13674 (N_13674,N_12484,N_12422);
or U13675 (N_13675,N_12395,N_12310);
or U13676 (N_13676,N_12145,N_12088);
nand U13677 (N_13677,N_11546,N_11359);
nand U13678 (N_13678,N_11519,N_12351);
or U13679 (N_13679,N_12137,N_11541);
or U13680 (N_13680,N_12430,N_12230);
nor U13681 (N_13681,N_11354,N_12200);
or U13682 (N_13682,N_12348,N_12114);
or U13683 (N_13683,N_12432,N_12241);
nand U13684 (N_13684,N_12089,N_11937);
xor U13685 (N_13685,N_11544,N_11524);
nor U13686 (N_13686,N_12493,N_12184);
or U13687 (N_13687,N_11253,N_12152);
nand U13688 (N_13688,N_11365,N_12314);
nor U13689 (N_13689,N_12448,N_12213);
nand U13690 (N_13690,N_11669,N_11470);
and U13691 (N_13691,N_12176,N_11734);
or U13692 (N_13692,N_12337,N_12185);
nor U13693 (N_13693,N_11504,N_12362);
xnor U13694 (N_13694,N_12094,N_12190);
xnor U13695 (N_13695,N_11756,N_11733);
nor U13696 (N_13696,N_12010,N_11682);
nor U13697 (N_13697,N_11361,N_11451);
and U13698 (N_13698,N_12429,N_12107);
or U13699 (N_13699,N_12129,N_11644);
nand U13700 (N_13700,N_12083,N_12388);
xnor U13701 (N_13701,N_12065,N_11837);
xnor U13702 (N_13702,N_11900,N_11788);
or U13703 (N_13703,N_12407,N_11846);
xnor U13704 (N_13704,N_11498,N_12287);
or U13705 (N_13705,N_11383,N_11475);
nor U13706 (N_13706,N_11609,N_12451);
nand U13707 (N_13707,N_12096,N_11572);
xor U13708 (N_13708,N_11785,N_11959);
nand U13709 (N_13709,N_12409,N_11432);
xnor U13710 (N_13710,N_12284,N_12366);
and U13711 (N_13711,N_12377,N_11753);
nand U13712 (N_13712,N_11695,N_11507);
nor U13713 (N_13713,N_11922,N_12296);
and U13714 (N_13714,N_11424,N_11928);
nand U13715 (N_13715,N_11996,N_11729);
or U13716 (N_13716,N_11437,N_12222);
xnor U13717 (N_13717,N_11958,N_11895);
nor U13718 (N_13718,N_12261,N_11275);
nor U13719 (N_13719,N_11358,N_11273);
nand U13720 (N_13720,N_12018,N_11955);
nand U13721 (N_13721,N_12356,N_11730);
and U13722 (N_13722,N_12230,N_12054);
nand U13723 (N_13723,N_11865,N_11452);
and U13724 (N_13724,N_11802,N_12378);
xnor U13725 (N_13725,N_12140,N_11910);
or U13726 (N_13726,N_11694,N_11796);
and U13727 (N_13727,N_12327,N_11318);
or U13728 (N_13728,N_11417,N_11455);
or U13729 (N_13729,N_11914,N_12157);
or U13730 (N_13730,N_12207,N_12329);
and U13731 (N_13731,N_12124,N_11442);
xnor U13732 (N_13732,N_12480,N_11627);
nand U13733 (N_13733,N_12333,N_11857);
xnor U13734 (N_13734,N_12348,N_11878);
nor U13735 (N_13735,N_11437,N_11627);
nand U13736 (N_13736,N_11931,N_11410);
nand U13737 (N_13737,N_12171,N_11799);
or U13738 (N_13738,N_12289,N_12311);
xor U13739 (N_13739,N_11360,N_11420);
and U13740 (N_13740,N_12099,N_11979);
nand U13741 (N_13741,N_12403,N_12282);
nor U13742 (N_13742,N_12229,N_11897);
nand U13743 (N_13743,N_12067,N_11439);
or U13744 (N_13744,N_12186,N_11560);
xor U13745 (N_13745,N_11822,N_11745);
nand U13746 (N_13746,N_12483,N_12399);
xnor U13747 (N_13747,N_12170,N_11456);
and U13748 (N_13748,N_11306,N_11369);
and U13749 (N_13749,N_12336,N_11711);
and U13750 (N_13750,N_13281,N_13577);
xnor U13751 (N_13751,N_13490,N_13479);
or U13752 (N_13752,N_13294,N_12517);
xnor U13753 (N_13753,N_12998,N_13651);
nand U13754 (N_13754,N_12823,N_12813);
and U13755 (N_13755,N_13206,N_13165);
and U13756 (N_13756,N_12801,N_13072);
nand U13757 (N_13757,N_13696,N_13208);
nor U13758 (N_13758,N_13299,N_12982);
nor U13759 (N_13759,N_12554,N_12534);
xor U13760 (N_13760,N_13285,N_12874);
or U13761 (N_13761,N_12533,N_13369);
nand U13762 (N_13762,N_12584,N_12603);
nor U13763 (N_13763,N_13622,N_13424);
nor U13764 (N_13764,N_13460,N_13017);
nor U13765 (N_13765,N_12546,N_13061);
xnor U13766 (N_13766,N_12824,N_12610);
nor U13767 (N_13767,N_12591,N_12588);
xor U13768 (N_13768,N_13446,N_13267);
and U13769 (N_13769,N_13467,N_12582);
or U13770 (N_13770,N_13471,N_12736);
nand U13771 (N_13771,N_13270,N_12864);
or U13772 (N_13772,N_13032,N_12629);
or U13773 (N_13773,N_13404,N_13402);
nor U13774 (N_13774,N_12903,N_13398);
xnor U13775 (N_13775,N_12740,N_12711);
nand U13776 (N_13776,N_13576,N_12835);
xnor U13777 (N_13777,N_13134,N_12741);
nor U13778 (N_13778,N_13192,N_12978);
and U13779 (N_13779,N_12640,N_13125);
xnor U13780 (N_13780,N_13458,N_12726);
nor U13781 (N_13781,N_12605,N_13633);
or U13782 (N_13782,N_13656,N_13305);
and U13783 (N_13783,N_13554,N_12519);
and U13784 (N_13784,N_13002,N_13136);
nand U13785 (N_13785,N_13298,N_13314);
xor U13786 (N_13786,N_12771,N_13496);
nand U13787 (N_13787,N_13198,N_13516);
and U13788 (N_13788,N_13083,N_13033);
xnor U13789 (N_13789,N_12972,N_13105);
xor U13790 (N_13790,N_12722,N_12829);
xnor U13791 (N_13791,N_13413,N_12565);
nor U13792 (N_13792,N_13023,N_13655);
nand U13793 (N_13793,N_13274,N_12785);
and U13794 (N_13794,N_13272,N_13139);
or U13795 (N_13795,N_13171,N_12971);
xor U13796 (N_13796,N_13090,N_13623);
and U13797 (N_13797,N_13532,N_12757);
nor U13798 (N_13798,N_13037,N_13287);
or U13799 (N_13799,N_13191,N_13475);
nor U13800 (N_13800,N_13015,N_13558);
nand U13801 (N_13801,N_13326,N_12849);
and U13802 (N_13802,N_13635,N_12822);
or U13803 (N_13803,N_12875,N_13079);
and U13804 (N_13804,N_13720,N_12936);
nor U13805 (N_13805,N_13617,N_12861);
or U13806 (N_13806,N_12880,N_13324);
xor U13807 (N_13807,N_13268,N_13234);
and U13808 (N_13808,N_12995,N_12963);
nand U13809 (N_13809,N_13440,N_13642);
or U13810 (N_13810,N_13641,N_12983);
and U13811 (N_13811,N_12539,N_12789);
or U13812 (N_13812,N_13086,N_13040);
xnor U13813 (N_13813,N_12745,N_13560);
or U13814 (N_13814,N_12706,N_12516);
nand U13815 (N_13815,N_12887,N_13159);
nand U13816 (N_13816,N_13506,N_13189);
and U13817 (N_13817,N_13379,N_13525);
and U13818 (N_13818,N_13570,N_12670);
xor U13819 (N_13819,N_12797,N_13420);
or U13820 (N_13820,N_12675,N_13618);
nor U13821 (N_13821,N_13556,N_13109);
or U13822 (N_13822,N_13595,N_13010);
or U13823 (N_13823,N_13114,N_12773);
or U13824 (N_13824,N_13135,N_12781);
nor U13825 (N_13825,N_12643,N_13513);
or U13826 (N_13826,N_12889,N_12557);
or U13827 (N_13827,N_13605,N_13749);
nand U13828 (N_13828,N_12809,N_13569);
nor U13829 (N_13829,N_13322,N_13680);
xnor U13830 (N_13830,N_13397,N_13470);
nor U13831 (N_13831,N_12762,N_13162);
nand U13832 (N_13832,N_13190,N_12876);
or U13833 (N_13833,N_13020,N_13223);
and U13834 (N_13834,N_13176,N_12505);
nand U13835 (N_13835,N_13414,N_13627);
xnor U13836 (N_13836,N_13522,N_12597);
or U13837 (N_13837,N_13080,N_13148);
or U13838 (N_13838,N_12676,N_13665);
or U13839 (N_13839,N_13256,N_13473);
nand U13840 (N_13840,N_13687,N_13078);
or U13841 (N_13841,N_13621,N_13207);
xor U13842 (N_13842,N_13710,N_12904);
nor U13843 (N_13843,N_13315,N_12525);
xor U13844 (N_13844,N_13393,N_13663);
xnor U13845 (N_13845,N_12850,N_13110);
nor U13846 (N_13846,N_12622,N_13412);
and U13847 (N_13847,N_13572,N_12716);
xor U13848 (N_13848,N_13368,N_12941);
xor U13849 (N_13849,N_13401,N_13491);
nor U13850 (N_13850,N_13372,N_13505);
nand U13851 (N_13851,N_13484,N_13611);
or U13852 (N_13852,N_13131,N_12820);
xnor U13853 (N_13853,N_13409,N_13047);
and U13854 (N_13854,N_13468,N_13012);
nor U13855 (N_13855,N_13153,N_12614);
nor U13856 (N_13856,N_13297,N_13711);
xnor U13857 (N_13857,N_12947,N_13138);
nand U13858 (N_13858,N_13646,N_13265);
nor U13859 (N_13859,N_13422,N_12916);
and U13860 (N_13860,N_13133,N_13681);
nand U13861 (N_13861,N_12725,N_12713);
nand U13862 (N_13862,N_13673,N_12768);
nor U13863 (N_13863,N_13445,N_12625);
nand U13864 (N_13864,N_12520,N_13250);
or U13865 (N_13865,N_13154,N_13477);
or U13866 (N_13866,N_12949,N_13302);
nand U13867 (N_13867,N_12604,N_13689);
nor U13868 (N_13868,N_12631,N_13310);
nand U13869 (N_13869,N_12727,N_12872);
xnor U13870 (N_13870,N_13524,N_12718);
or U13871 (N_13871,N_13355,N_12923);
or U13872 (N_13872,N_12977,N_12993);
and U13873 (N_13873,N_13518,N_13586);
and U13874 (N_13874,N_12551,N_12833);
or U13875 (N_13875,N_13435,N_13335);
nor U13876 (N_13876,N_12828,N_12693);
or U13877 (N_13877,N_12502,N_12930);
or U13878 (N_13878,N_13249,N_13476);
xnor U13879 (N_13879,N_13193,N_13727);
and U13880 (N_13880,N_13129,N_12894);
and U13881 (N_13881,N_12704,N_13236);
nand U13882 (N_13882,N_13003,N_13046);
nand U13883 (N_13883,N_12843,N_12842);
xor U13884 (N_13884,N_13004,N_13427);
or U13885 (N_13885,N_12994,N_13005);
nor U13886 (N_13886,N_12856,N_13742);
xor U13887 (N_13887,N_13120,N_13459);
nand U13888 (N_13888,N_12883,N_12796);
and U13889 (N_13889,N_13688,N_13116);
nand U13890 (N_13890,N_12900,N_13073);
nand U13891 (N_13891,N_13062,N_13026);
or U13892 (N_13892,N_12668,N_13589);
xnor U13893 (N_13893,N_13247,N_13624);
or U13894 (N_13894,N_12770,N_12553);
or U13895 (N_13895,N_12970,N_12613);
or U13896 (N_13896,N_13312,N_13546);
or U13897 (N_13897,N_13432,N_13735);
nor U13898 (N_13898,N_12538,N_13300);
or U13899 (N_13899,N_13739,N_12737);
and U13900 (N_13900,N_12927,N_12667);
or U13901 (N_13901,N_12576,N_13181);
or U13902 (N_13902,N_13451,N_12961);
and U13903 (N_13903,N_12836,N_12791);
nor U13904 (N_13904,N_12556,N_13466);
nor U13905 (N_13905,N_13151,N_12967);
or U13906 (N_13906,N_12811,N_13018);
xor U13907 (N_13907,N_13500,N_13488);
or U13908 (N_13908,N_12510,N_13241);
nand U13909 (N_13909,N_12608,N_13150);
nand U13910 (N_13910,N_13041,N_12760);
xor U13911 (N_13911,N_12871,N_13504);
nor U13912 (N_13912,N_13564,N_12763);
or U13913 (N_13913,N_12662,N_12599);
and U13914 (N_13914,N_12710,N_12508);
nand U13915 (N_13915,N_13631,N_12687);
or U13916 (N_13916,N_13403,N_13147);
nor U13917 (N_13917,N_13721,N_13231);
xor U13918 (N_13918,N_13140,N_13024);
xnor U13919 (N_13919,N_13678,N_12764);
nor U13920 (N_13920,N_12504,N_12511);
nor U13921 (N_13921,N_12786,N_13647);
xor U13922 (N_13922,N_13196,N_13517);
and U13923 (N_13923,N_12800,N_13666);
and U13924 (N_13924,N_12937,N_12681);
or U13925 (N_13925,N_12761,N_13527);
or U13926 (N_13926,N_12714,N_13694);
or U13927 (N_13927,N_13013,N_13718);
or U13928 (N_13928,N_13685,N_12598);
nor U13929 (N_13929,N_12689,N_13269);
xor U13930 (N_13930,N_12901,N_12717);
and U13931 (N_13931,N_12956,N_12908);
and U13932 (N_13932,N_12924,N_13301);
xnor U13933 (N_13933,N_12543,N_13734);
and U13934 (N_13934,N_12766,N_13657);
xor U13935 (N_13935,N_13229,N_13728);
nor U13936 (N_13936,N_12968,N_13438);
nand U13937 (N_13937,N_13587,N_13474);
nand U13938 (N_13938,N_12688,N_13658);
or U13939 (N_13939,N_13060,N_13156);
and U13940 (N_13940,N_12735,N_12656);
and U13941 (N_13941,N_12780,N_13327);
or U13942 (N_13942,N_13434,N_12902);
or U13943 (N_13943,N_12609,N_13064);
nor U13944 (N_13944,N_13743,N_13308);
xor U13945 (N_13945,N_13709,N_12756);
or U13946 (N_13946,N_12847,N_13723);
or U13947 (N_13947,N_13463,N_12618);
nor U13948 (N_13948,N_13160,N_13701);
nor U13949 (N_13949,N_13000,N_13245);
nand U13950 (N_13950,N_13295,N_12514);
nand U13951 (N_13951,N_13540,N_13482);
nand U13952 (N_13952,N_13058,N_13669);
xor U13953 (N_13953,N_13545,N_12832);
and U13954 (N_13954,N_13132,N_13747);
and U13955 (N_13955,N_13660,N_13199);
xor U13956 (N_13956,N_13653,N_12571);
xnor U13957 (N_13957,N_12996,N_13280);
or U13958 (N_13958,N_12933,N_13009);
nor U13959 (N_13959,N_13008,N_12938);
nand U13960 (N_13960,N_13328,N_13714);
nor U13961 (N_13961,N_13604,N_13194);
nand U13962 (N_13962,N_13130,N_13098);
and U13963 (N_13963,N_13630,N_13523);
or U13964 (N_13964,N_13429,N_12500);
and U13965 (N_13965,N_12803,N_12753);
or U13966 (N_13966,N_13338,N_12729);
nor U13967 (N_13967,N_12863,N_12792);
and U13968 (N_13968,N_13126,N_12953);
xor U13969 (N_13969,N_13279,N_13481);
or U13970 (N_13970,N_13317,N_13386);
and U13971 (N_13971,N_13602,N_13464);
or U13972 (N_13972,N_13498,N_13052);
nand U13973 (N_13973,N_13717,N_13392);
and U13974 (N_13974,N_13497,N_13185);
or U13975 (N_13975,N_13608,N_12945);
and U13976 (N_13976,N_13519,N_13431);
and U13977 (N_13977,N_12660,N_13675);
nor U13978 (N_13978,N_12564,N_13495);
xor U13979 (N_13979,N_12645,N_13145);
nand U13980 (N_13980,N_13515,N_13690);
nand U13981 (N_13981,N_12651,N_13084);
and U13982 (N_13982,N_13699,N_13400);
and U13983 (N_13983,N_13542,N_12795);
xnor U13984 (N_13984,N_13552,N_12547);
xnor U13985 (N_13985,N_13609,N_12585);
or U13986 (N_13986,N_13211,N_13313);
nor U13987 (N_13987,N_13164,N_12862);
or U13988 (N_13988,N_13579,N_13288);
or U13989 (N_13989,N_12881,N_12815);
xnor U13990 (N_13990,N_12913,N_12669);
and U13991 (N_13991,N_13501,N_13691);
nand U13992 (N_13992,N_12733,N_12921);
and U13993 (N_13993,N_12845,N_13296);
xnor U13994 (N_13994,N_12911,N_12653);
xnor U13995 (N_13995,N_13067,N_12981);
nor U13996 (N_13996,N_13447,N_13391);
or U13997 (N_13997,N_13232,N_12805);
nand U13998 (N_13998,N_13365,N_12743);
nor U13999 (N_13999,N_13548,N_12919);
or U14000 (N_14000,N_12991,N_13614);
xor U14001 (N_14001,N_12866,N_13584);
or U14002 (N_14002,N_13538,N_13428);
and U14003 (N_14003,N_13146,N_13492);
xnor U14004 (N_14004,N_13648,N_12744);
nor U14005 (N_14005,N_12952,N_13092);
nand U14006 (N_14006,N_13233,N_13430);
xnor U14007 (N_14007,N_13507,N_13591);
xnor U14008 (N_14008,N_13607,N_12954);
xor U14009 (N_14009,N_13097,N_13662);
xnor U14010 (N_14010,N_13748,N_13354);
and U14011 (N_14011,N_13531,N_13021);
and U14012 (N_14012,N_12635,N_13284);
nand U14013 (N_14013,N_13246,N_13143);
and U14014 (N_14014,N_13104,N_12686);
and U14015 (N_14015,N_12559,N_13186);
nor U14016 (N_14016,N_13347,N_13225);
nand U14017 (N_14017,N_12581,N_12567);
and U14018 (N_14018,N_12708,N_13337);
nand U14019 (N_14019,N_13261,N_13571);
and U14020 (N_14020,N_13228,N_13601);
nand U14021 (N_14021,N_13227,N_13112);
or U14022 (N_14022,N_12917,N_13407);
nor U14023 (N_14023,N_13553,N_13559);
xor U14024 (N_14024,N_12988,N_13535);
nor U14025 (N_14025,N_13119,N_12573);
or U14026 (N_14026,N_12929,N_12989);
or U14027 (N_14027,N_12707,N_13346);
xor U14028 (N_14028,N_13361,N_13426);
xnor U14029 (N_14029,N_13043,N_13273);
and U14030 (N_14030,N_13672,N_13257);
xnor U14031 (N_14031,N_13142,N_13539);
and U14032 (N_14032,N_13082,N_13732);
nor U14033 (N_14033,N_13240,N_12987);
nand U14034 (N_14034,N_13421,N_12626);
and U14035 (N_14035,N_13537,N_13551);
and U14036 (N_14036,N_12526,N_13448);
or U14037 (N_14037,N_13737,N_13209);
and U14038 (N_14038,N_12906,N_13528);
nand U14039 (N_14039,N_13030,N_12672);
and U14040 (N_14040,N_13170,N_13332);
nor U14041 (N_14041,N_13574,N_12657);
nor U14042 (N_14042,N_13321,N_12790);
nand U14043 (N_14043,N_13416,N_13725);
and U14044 (N_14044,N_12531,N_12958);
xor U14045 (N_14045,N_12839,N_12893);
or U14046 (N_14046,N_13529,N_13596);
and U14047 (N_14047,N_12979,N_13059);
or U14048 (N_14048,N_13252,N_12728);
nand U14049 (N_14049,N_13521,N_13550);
or U14050 (N_14050,N_12831,N_13385);
nor U14051 (N_14051,N_13716,N_12617);
and U14052 (N_14052,N_13128,N_13203);
or U14053 (N_14053,N_12999,N_12962);
or U14054 (N_14054,N_12854,N_12819);
nand U14055 (N_14055,N_13638,N_13406);
nand U14056 (N_14056,N_13336,N_13254);
or U14057 (N_14057,N_13307,N_12755);
or U14058 (N_14058,N_13306,N_13330);
or U14059 (N_14059,N_12884,N_12747);
and U14060 (N_14060,N_13544,N_13436);
and U14061 (N_14061,N_13619,N_12623);
nor U14062 (N_14062,N_13668,N_13057);
and U14063 (N_14063,N_13113,N_13102);
nor U14064 (N_14064,N_13025,N_13616);
or U14065 (N_14065,N_13068,N_12868);
and U14066 (N_14066,N_13573,N_13123);
nand U14067 (N_14067,N_13399,N_13697);
and U14068 (N_14068,N_12895,N_12612);
xnor U14069 (N_14069,N_13536,N_13676);
nand U14070 (N_14070,N_12671,N_12548);
and U14071 (N_14071,N_13610,N_12788);
and U14072 (N_14072,N_12851,N_13253);
or U14073 (N_14073,N_13628,N_13715);
or U14074 (N_14074,N_12540,N_12787);
and U14075 (N_14075,N_13634,N_12509);
xor U14076 (N_14076,N_12536,N_13418);
and U14077 (N_14077,N_12709,N_13183);
xnor U14078 (N_14078,N_13100,N_13654);
nand U14079 (N_14079,N_12734,N_13659);
or U14080 (N_14080,N_12992,N_13303);
nand U14081 (N_14081,N_12632,N_12569);
or U14082 (N_14082,N_13698,N_13367);
nand U14083 (N_14083,N_13031,N_13686);
xnor U14084 (N_14084,N_13292,N_12684);
nand U14085 (N_14085,N_12664,N_13417);
nor U14086 (N_14086,N_12928,N_13316);
nand U14087 (N_14087,N_13629,N_13309);
or U14088 (N_14088,N_12939,N_13180);
and U14089 (N_14089,N_12746,N_12891);
or U14090 (N_14090,N_12518,N_13410);
and U14091 (N_14091,N_13039,N_13639);
and U14092 (N_14092,N_12965,N_12821);
nand U14093 (N_14093,N_13244,N_13218);
xor U14094 (N_14094,N_13383,N_12899);
and U14095 (N_14095,N_12860,N_13726);
nor U14096 (N_14096,N_13065,N_13583);
xnor U14097 (N_14097,N_12825,N_12870);
nand U14098 (N_14098,N_12558,N_13472);
and U14099 (N_14099,N_12658,N_13557);
nor U14100 (N_14100,N_12587,N_12951);
and U14101 (N_14101,N_12659,N_13349);
nand U14102 (N_14102,N_12649,N_12973);
nor U14103 (N_14103,N_13599,N_12619);
nand U14104 (N_14104,N_12633,N_13277);
or U14105 (N_14105,N_13351,N_12848);
and U14106 (N_14106,N_13419,N_13323);
nand U14107 (N_14107,N_12985,N_13625);
xor U14108 (N_14108,N_13217,N_12555);
nand U14109 (N_14109,N_12932,N_12877);
nand U14110 (N_14110,N_13543,N_13291);
and U14111 (N_14111,N_13405,N_12777);
and U14112 (N_14112,N_13370,N_13437);
nand U14113 (N_14113,N_13708,N_13028);
and U14114 (N_14114,N_13339,N_13455);
or U14115 (N_14115,N_13415,N_13325);
xnor U14116 (N_14116,N_13375,N_13489);
or U14117 (N_14117,N_13158,N_12654);
nor U14118 (N_14118,N_12544,N_12810);
nand U14119 (N_14119,N_12754,N_12959);
or U14120 (N_14120,N_12697,N_13612);
and U14121 (N_14121,N_13394,N_13585);
or U14122 (N_14122,N_12607,N_13111);
nand U14123 (N_14123,N_13567,N_12804);
and U14124 (N_14124,N_13029,N_12595);
xnor U14125 (N_14125,N_12673,N_13499);
nand U14126 (N_14126,N_13637,N_12909);
and U14127 (N_14127,N_13600,N_13063);
or U14128 (N_14128,N_12507,N_13344);
nor U14129 (N_14129,N_13166,N_13055);
nand U14130 (N_14130,N_12560,N_13106);
xor U14131 (N_14131,N_12580,N_12700);
nand U14132 (N_14132,N_13070,N_12696);
or U14133 (N_14133,N_13318,N_12752);
and U14134 (N_14134,N_13719,N_12568);
nand U14135 (N_14135,N_13243,N_12812);
nand U14136 (N_14136,N_12515,N_13620);
or U14137 (N_14137,N_13271,N_13178);
nand U14138 (N_14138,N_13329,N_13204);
nor U14139 (N_14139,N_12765,N_13568);
or U14140 (N_14140,N_12926,N_13103);
xor U14141 (N_14141,N_13237,N_13074);
and U14142 (N_14142,N_13425,N_13282);
and U14143 (N_14143,N_12637,N_13334);
nand U14144 (N_14144,N_13320,N_13212);
xnor U14145 (N_14145,N_13411,N_12814);
and U14146 (N_14146,N_12885,N_13371);
or U14147 (N_14147,N_12918,N_13377);
or U14148 (N_14148,N_12798,N_13094);
and U14149 (N_14149,N_12898,N_13157);
or U14150 (N_14150,N_13340,N_12550);
nand U14151 (N_14151,N_13179,N_13152);
nand U14152 (N_14152,N_12695,N_13373);
nand U14153 (N_14153,N_13664,N_13091);
nand U14154 (N_14154,N_13478,N_13096);
or U14155 (N_14155,N_13360,N_12719);
and U14156 (N_14156,N_12542,N_12677);
nor U14157 (N_14157,N_13606,N_13107);
or U14158 (N_14158,N_12855,N_12647);
nand U14159 (N_14159,N_13594,N_13045);
nor U14160 (N_14160,N_13457,N_13331);
xor U14161 (N_14161,N_12948,N_12620);
xor U14162 (N_14162,N_13740,N_13396);
and U14163 (N_14163,N_13260,N_12980);
nand U14164 (N_14164,N_13219,N_12665);
and U14165 (N_14165,N_12830,N_13362);
or U14166 (N_14166,N_13382,N_13692);
and U14167 (N_14167,N_13645,N_13289);
nor U14168 (N_14168,N_12524,N_12840);
nand U14169 (N_14169,N_13613,N_12692);
or U14170 (N_14170,N_12865,N_12974);
nor U14171 (N_14171,N_13357,N_13054);
xnor U14172 (N_14172,N_13707,N_13378);
nand U14173 (N_14173,N_13565,N_13235);
xor U14174 (N_14174,N_13118,N_13745);
nand U14175 (N_14175,N_13168,N_13187);
nand U14176 (N_14176,N_12624,N_12639);
nor U14177 (N_14177,N_12846,N_12615);
nor U14178 (N_14178,N_12512,N_13510);
xor U14179 (N_14179,N_12738,N_12589);
xnor U14180 (N_14180,N_12720,N_12644);
xnor U14181 (N_14181,N_13693,N_12691);
xnor U14182 (N_14182,N_12816,N_13069);
nor U14183 (N_14183,N_13049,N_13172);
xnor U14184 (N_14184,N_13441,N_12882);
xnor U14185 (N_14185,N_12794,N_13014);
nor U14186 (N_14186,N_13652,N_13262);
and U14187 (N_14187,N_12818,N_13483);
and U14188 (N_14188,N_12873,N_13333);
nor U14189 (N_14189,N_12907,N_12562);
and U14190 (N_14190,N_13444,N_13242);
xnor U14191 (N_14191,N_12783,N_13580);
nor U14192 (N_14192,N_12826,N_12793);
xor U14193 (N_14193,N_12674,N_13077);
xnor U14194 (N_14194,N_12878,N_13454);
and U14195 (N_14195,N_12506,N_13449);
xnor U14196 (N_14196,N_13149,N_12621);
and U14197 (N_14197,N_13650,N_13514);
or U14198 (N_14198,N_13095,N_12975);
xnor U14199 (N_14199,N_13615,N_13578);
or U14200 (N_14200,N_13075,N_12575);
and U14201 (N_14201,N_13636,N_13342);
and U14202 (N_14202,N_13359,N_12532);
xor U14203 (N_14203,N_13007,N_12636);
nor U14204 (N_14204,N_13487,N_13376);
or U14205 (N_14205,N_13744,N_12966);
xor U14206 (N_14206,N_13290,N_12925);
and U14207 (N_14207,N_12778,N_13216);
nand U14208 (N_14208,N_12986,N_13001);
and U14209 (N_14209,N_12858,N_13705);
nor U14210 (N_14210,N_13713,N_13016);
xnor U14211 (N_14211,N_12552,N_12853);
nor U14212 (N_14212,N_12593,N_12522);
nor U14213 (N_14213,N_13526,N_12606);
xnor U14214 (N_14214,N_12642,N_13184);
and U14215 (N_14215,N_12879,N_12663);
and U14216 (N_14216,N_13038,N_12561);
nand U14217 (N_14217,N_12600,N_12503);
xnor U14218 (N_14218,N_12701,N_13695);
or U14219 (N_14219,N_13640,N_13230);
nand U14220 (N_14220,N_13452,N_13450);
or U14221 (N_14221,N_12890,N_12683);
nand U14222 (N_14222,N_13683,N_12934);
and U14223 (N_14223,N_12579,N_13155);
xnor U14224 (N_14224,N_12774,N_12723);
and U14225 (N_14225,N_13248,N_13733);
and U14226 (N_14226,N_13035,N_13044);
nand U14227 (N_14227,N_12806,N_13278);
nor U14228 (N_14228,N_12944,N_13626);
nand U14229 (N_14229,N_12808,N_12590);
nand U14230 (N_14230,N_12946,N_13239);
nand U14231 (N_14231,N_12844,N_13533);
nand U14232 (N_14232,N_12852,N_13561);
xor U14233 (N_14233,N_12680,N_13343);
nand U14234 (N_14234,N_12931,N_12827);
nand U14235 (N_14235,N_13366,N_13122);
nor U14236 (N_14236,N_13076,N_13433);
nand U14237 (N_14237,N_13210,N_13121);
nor U14238 (N_14238,N_12782,N_13443);
and U14239 (N_14239,N_13549,N_12648);
or U14240 (N_14240,N_13702,N_12712);
nand U14241 (N_14241,N_13163,N_13706);
nand U14242 (N_14242,N_13224,N_13364);
nand U14243 (N_14243,N_13682,N_13036);
nand U14244 (N_14244,N_13387,N_12731);
and U14245 (N_14245,N_13053,N_13541);
nand U14246 (N_14246,N_12838,N_13089);
nor U14247 (N_14247,N_12769,N_13643);
xor U14248 (N_14248,N_13304,N_13311);
and U14249 (N_14249,N_13502,N_13174);
nor U14250 (N_14250,N_13511,N_13006);
and U14251 (N_14251,N_12969,N_13679);
xnor U14252 (N_14252,N_13731,N_12630);
nand U14253 (N_14253,N_12702,N_13081);
or U14254 (N_14254,N_13590,N_12549);
or U14255 (N_14255,N_13712,N_12922);
nand U14256 (N_14256,N_13108,N_13220);
xor U14257 (N_14257,N_13480,N_12976);
nor U14258 (N_14258,N_13746,N_13520);
and U14259 (N_14259,N_13741,N_13205);
nand U14260 (N_14260,N_13341,N_13175);
nor U14261 (N_14261,N_13390,N_12742);
and U14262 (N_14262,N_13222,N_13259);
xor U14263 (N_14263,N_12570,N_12817);
nand U14264 (N_14264,N_12751,N_12748);
and U14265 (N_14265,N_12578,N_13088);
nor U14266 (N_14266,N_13197,N_12732);
and U14267 (N_14267,N_13453,N_13388);
nand U14268 (N_14268,N_12592,N_12586);
nand U14269 (N_14269,N_12940,N_12772);
nor U14270 (N_14270,N_12807,N_12601);
and U14271 (N_14271,N_12694,N_13345);
nand U14272 (N_14272,N_12682,N_13729);
or U14273 (N_14273,N_13465,N_12984);
nand U14274 (N_14274,N_12572,N_13177);
xnor U14275 (N_14275,N_13127,N_12935);
and U14276 (N_14276,N_13182,N_12721);
or U14277 (N_14277,N_13704,N_12679);
nand U14278 (N_14278,N_12920,N_13534);
or U14279 (N_14279,N_12943,N_13019);
xor U14280 (N_14280,N_13071,N_13684);
nand U14281 (N_14281,N_13169,N_13144);
nor U14282 (N_14282,N_12841,N_13442);
xnor U14283 (N_14283,N_13381,N_12739);
xor U14284 (N_14284,N_12652,N_13509);
nor U14285 (N_14285,N_13356,N_12775);
nor U14286 (N_14286,N_13319,N_12779);
nand U14287 (N_14287,N_12759,N_12705);
xor U14288 (N_14288,N_12523,N_13736);
nor U14289 (N_14289,N_12638,N_12802);
nor U14290 (N_14290,N_13581,N_13493);
nand U14291 (N_14291,N_13115,N_13093);
or U14292 (N_14292,N_13603,N_12990);
nor U14293 (N_14293,N_12545,N_13215);
nor U14294 (N_14294,N_13724,N_12834);
and U14295 (N_14295,N_13085,N_12528);
or U14296 (N_14296,N_12646,N_12698);
xor U14297 (N_14297,N_12594,N_13293);
and U14298 (N_14298,N_12892,N_12583);
and U14299 (N_14299,N_13547,N_12857);
and U14300 (N_14300,N_13661,N_13384);
xnor U14301 (N_14301,N_12602,N_12955);
nand U14302 (N_14302,N_13348,N_12513);
and U14303 (N_14303,N_13258,N_12650);
nor U14304 (N_14304,N_12915,N_13508);
nor U14305 (N_14305,N_13195,N_13674);
and U14306 (N_14306,N_13188,N_13530);
nor U14307 (N_14307,N_12501,N_13066);
xnor U14308 (N_14308,N_12699,N_13738);
and U14309 (N_14309,N_12799,N_12897);
and U14310 (N_14310,N_13408,N_13389);
nor U14311 (N_14311,N_12566,N_13512);
nand U14312 (N_14312,N_12837,N_12521);
xor U14313 (N_14313,N_12767,N_13555);
and U14314 (N_14314,N_13563,N_12730);
nand U14315 (N_14315,N_12577,N_13275);
or U14316 (N_14316,N_13700,N_13667);
and U14317 (N_14317,N_13461,N_12957);
nor U14318 (N_14318,N_13439,N_13562);
or U14319 (N_14319,N_13213,N_13101);
and U14320 (N_14320,N_13137,N_13173);
and U14321 (N_14321,N_13374,N_12950);
nor U14322 (N_14322,N_13503,N_12715);
and U14323 (N_14323,N_13592,N_13575);
xnor U14324 (N_14324,N_13263,N_12563);
nor U14325 (N_14325,N_12611,N_13632);
xor U14326 (N_14326,N_12888,N_13048);
or U14327 (N_14327,N_13124,N_12690);
or U14328 (N_14328,N_12960,N_13167);
nand U14329 (N_14329,N_12910,N_13649);
and U14330 (N_14330,N_12678,N_12784);
or U14331 (N_14331,N_13670,N_13251);
nand U14332 (N_14332,N_13276,N_13593);
or U14333 (N_14333,N_12867,N_13597);
xor U14334 (N_14334,N_12537,N_13352);
nand U14335 (N_14335,N_13027,N_13056);
nand U14336 (N_14336,N_13350,N_13486);
and U14337 (N_14337,N_13395,N_13034);
or U14338 (N_14338,N_13566,N_12685);
nor U14339 (N_14339,N_13598,N_13286);
nand U14340 (N_14340,N_13363,N_13099);
or U14341 (N_14341,N_13671,N_13141);
nor U14342 (N_14342,N_12655,N_13582);
and U14343 (N_14343,N_13353,N_13221);
nand U14344 (N_14344,N_12758,N_13042);
xor U14345 (N_14345,N_13485,N_12776);
or U14346 (N_14346,N_12896,N_13494);
nor U14347 (N_14347,N_12964,N_13462);
and U14348 (N_14348,N_12541,N_13456);
or U14349 (N_14349,N_12574,N_13238);
nor U14350 (N_14350,N_13469,N_12905);
and U14351 (N_14351,N_12914,N_13050);
and U14352 (N_14352,N_13051,N_12535);
nor U14353 (N_14353,N_12749,N_13226);
nand U14354 (N_14354,N_12596,N_12641);
xor U14355 (N_14355,N_12869,N_12859);
nand U14356 (N_14356,N_13161,N_12997);
and U14357 (N_14357,N_13358,N_13255);
or U14358 (N_14358,N_13117,N_13283);
nor U14359 (N_14359,N_13730,N_13380);
nor U14360 (N_14360,N_13087,N_12530);
and U14361 (N_14361,N_13644,N_13011);
nor U14362 (N_14362,N_12886,N_12634);
or U14363 (N_14363,N_13200,N_12529);
or U14364 (N_14364,N_13022,N_13588);
and U14365 (N_14365,N_12527,N_13703);
nor U14366 (N_14366,N_12750,N_13266);
nor U14367 (N_14367,N_13214,N_12616);
nor U14368 (N_14368,N_13201,N_12627);
xor U14369 (N_14369,N_12942,N_13677);
nand U14370 (N_14370,N_12912,N_13202);
nand U14371 (N_14371,N_13423,N_13264);
and U14372 (N_14372,N_12628,N_12666);
xnor U14373 (N_14373,N_12661,N_12724);
and U14374 (N_14374,N_13722,N_12703);
nand U14375 (N_14375,N_13429,N_12806);
xnor U14376 (N_14376,N_13100,N_13157);
and U14377 (N_14377,N_12774,N_13414);
xor U14378 (N_14378,N_13381,N_13023);
nor U14379 (N_14379,N_12839,N_13316);
and U14380 (N_14380,N_12589,N_13545);
xor U14381 (N_14381,N_13095,N_13268);
and U14382 (N_14382,N_13376,N_13456);
or U14383 (N_14383,N_12832,N_13703);
xor U14384 (N_14384,N_12553,N_13314);
nand U14385 (N_14385,N_12632,N_13436);
nor U14386 (N_14386,N_12627,N_12529);
nand U14387 (N_14387,N_13212,N_12512);
and U14388 (N_14388,N_12500,N_13248);
xnor U14389 (N_14389,N_12548,N_13665);
and U14390 (N_14390,N_12539,N_12834);
or U14391 (N_14391,N_13077,N_13335);
nor U14392 (N_14392,N_12629,N_13367);
nand U14393 (N_14393,N_12851,N_12609);
and U14394 (N_14394,N_13272,N_13727);
xnor U14395 (N_14395,N_13290,N_12673);
nor U14396 (N_14396,N_12967,N_13605);
nand U14397 (N_14397,N_13190,N_13479);
xnor U14398 (N_14398,N_13509,N_13335);
and U14399 (N_14399,N_13624,N_13291);
and U14400 (N_14400,N_13449,N_12503);
or U14401 (N_14401,N_12978,N_13532);
nor U14402 (N_14402,N_12789,N_12522);
nand U14403 (N_14403,N_13342,N_12919);
nor U14404 (N_14404,N_12782,N_13096);
and U14405 (N_14405,N_13726,N_12556);
xnor U14406 (N_14406,N_13711,N_13744);
or U14407 (N_14407,N_12913,N_13612);
nor U14408 (N_14408,N_13521,N_13361);
xnor U14409 (N_14409,N_13272,N_13290);
nor U14410 (N_14410,N_13136,N_12991);
nand U14411 (N_14411,N_13167,N_13231);
or U14412 (N_14412,N_13617,N_12937);
nor U14413 (N_14413,N_13461,N_13407);
and U14414 (N_14414,N_13213,N_12650);
nor U14415 (N_14415,N_12941,N_12714);
xor U14416 (N_14416,N_13002,N_13550);
nor U14417 (N_14417,N_12829,N_12601);
nand U14418 (N_14418,N_12805,N_12896);
xnor U14419 (N_14419,N_12642,N_13082);
and U14420 (N_14420,N_12916,N_13168);
nand U14421 (N_14421,N_13480,N_13307);
or U14422 (N_14422,N_12880,N_13499);
xor U14423 (N_14423,N_12949,N_13311);
nand U14424 (N_14424,N_12968,N_13584);
nor U14425 (N_14425,N_13003,N_13493);
and U14426 (N_14426,N_13582,N_13180);
or U14427 (N_14427,N_12722,N_13300);
nand U14428 (N_14428,N_13373,N_12538);
xor U14429 (N_14429,N_13004,N_12891);
xor U14430 (N_14430,N_13180,N_12569);
and U14431 (N_14431,N_13597,N_13591);
or U14432 (N_14432,N_13221,N_12949);
or U14433 (N_14433,N_13368,N_12503);
nand U14434 (N_14434,N_12648,N_13369);
nor U14435 (N_14435,N_13645,N_13590);
xor U14436 (N_14436,N_12621,N_13704);
and U14437 (N_14437,N_13429,N_12969);
nor U14438 (N_14438,N_13642,N_12987);
or U14439 (N_14439,N_13149,N_12624);
nand U14440 (N_14440,N_13498,N_13252);
nor U14441 (N_14441,N_12896,N_13415);
nor U14442 (N_14442,N_13488,N_12824);
nor U14443 (N_14443,N_12747,N_13421);
nor U14444 (N_14444,N_13675,N_12798);
xor U14445 (N_14445,N_12935,N_13439);
and U14446 (N_14446,N_12710,N_12533);
or U14447 (N_14447,N_12721,N_12505);
nor U14448 (N_14448,N_12823,N_12926);
nor U14449 (N_14449,N_13158,N_12516);
or U14450 (N_14450,N_13234,N_12777);
and U14451 (N_14451,N_13554,N_13570);
and U14452 (N_14452,N_12664,N_13172);
nor U14453 (N_14453,N_13589,N_13697);
or U14454 (N_14454,N_13400,N_13444);
xnor U14455 (N_14455,N_13127,N_13430);
nor U14456 (N_14456,N_12977,N_12926);
or U14457 (N_14457,N_13309,N_13055);
or U14458 (N_14458,N_12763,N_13353);
or U14459 (N_14459,N_13661,N_13075);
xnor U14460 (N_14460,N_13651,N_13096);
and U14461 (N_14461,N_13056,N_13372);
nor U14462 (N_14462,N_12767,N_12995);
nand U14463 (N_14463,N_13070,N_12802);
nand U14464 (N_14464,N_13317,N_13210);
nand U14465 (N_14465,N_12905,N_12596);
xor U14466 (N_14466,N_13625,N_13308);
nor U14467 (N_14467,N_13320,N_13440);
nor U14468 (N_14468,N_13456,N_12577);
xnor U14469 (N_14469,N_13010,N_13330);
and U14470 (N_14470,N_12856,N_12991);
or U14471 (N_14471,N_13327,N_12822);
and U14472 (N_14472,N_13058,N_12928);
and U14473 (N_14473,N_12550,N_13136);
and U14474 (N_14474,N_13039,N_12590);
and U14475 (N_14475,N_13644,N_12981);
nand U14476 (N_14476,N_12774,N_13647);
xor U14477 (N_14477,N_12821,N_13435);
xor U14478 (N_14478,N_13104,N_13535);
xnor U14479 (N_14479,N_13392,N_12632);
nand U14480 (N_14480,N_13207,N_13083);
or U14481 (N_14481,N_12888,N_13227);
nor U14482 (N_14482,N_12836,N_13636);
or U14483 (N_14483,N_13658,N_13635);
or U14484 (N_14484,N_12865,N_12835);
nand U14485 (N_14485,N_12734,N_13381);
or U14486 (N_14486,N_12811,N_13546);
nor U14487 (N_14487,N_13423,N_13431);
or U14488 (N_14488,N_13438,N_13587);
nor U14489 (N_14489,N_13341,N_12684);
nand U14490 (N_14490,N_13227,N_12811);
or U14491 (N_14491,N_12777,N_12964);
or U14492 (N_14492,N_12745,N_13453);
nand U14493 (N_14493,N_12756,N_13468);
nand U14494 (N_14494,N_13072,N_12554);
nor U14495 (N_14495,N_13669,N_13514);
and U14496 (N_14496,N_13011,N_13215);
nor U14497 (N_14497,N_12884,N_12978);
xnor U14498 (N_14498,N_13480,N_13739);
xor U14499 (N_14499,N_13133,N_12876);
xor U14500 (N_14500,N_13722,N_12669);
xor U14501 (N_14501,N_13643,N_13399);
or U14502 (N_14502,N_13649,N_13312);
nor U14503 (N_14503,N_13748,N_12952);
or U14504 (N_14504,N_12788,N_13411);
xnor U14505 (N_14505,N_13038,N_13261);
nor U14506 (N_14506,N_12917,N_13554);
or U14507 (N_14507,N_13499,N_13331);
xor U14508 (N_14508,N_12614,N_12555);
nand U14509 (N_14509,N_12820,N_12707);
nor U14510 (N_14510,N_13713,N_13282);
nor U14511 (N_14511,N_13323,N_13513);
nand U14512 (N_14512,N_12789,N_13346);
or U14513 (N_14513,N_12561,N_13320);
or U14514 (N_14514,N_12842,N_13249);
nor U14515 (N_14515,N_12775,N_12689);
and U14516 (N_14516,N_12545,N_12606);
or U14517 (N_14517,N_13056,N_12985);
nor U14518 (N_14518,N_12978,N_12676);
nor U14519 (N_14519,N_13249,N_13676);
xnor U14520 (N_14520,N_12570,N_12829);
xnor U14521 (N_14521,N_12757,N_12766);
xor U14522 (N_14522,N_13578,N_12685);
and U14523 (N_14523,N_13560,N_13011);
nor U14524 (N_14524,N_12559,N_12638);
or U14525 (N_14525,N_13540,N_12576);
xor U14526 (N_14526,N_13479,N_13038);
and U14527 (N_14527,N_12846,N_12538);
nor U14528 (N_14528,N_13159,N_13306);
and U14529 (N_14529,N_13220,N_12865);
nor U14530 (N_14530,N_12579,N_13327);
xnor U14531 (N_14531,N_12827,N_13154);
xor U14532 (N_14532,N_13236,N_13087);
or U14533 (N_14533,N_12647,N_13060);
and U14534 (N_14534,N_13206,N_12595);
and U14535 (N_14535,N_13045,N_13397);
nand U14536 (N_14536,N_13688,N_12842);
and U14537 (N_14537,N_13227,N_12786);
nor U14538 (N_14538,N_12996,N_13673);
nor U14539 (N_14539,N_12848,N_13086);
and U14540 (N_14540,N_13663,N_12727);
or U14541 (N_14541,N_13381,N_12747);
and U14542 (N_14542,N_13175,N_13277);
xnor U14543 (N_14543,N_13133,N_13740);
xnor U14544 (N_14544,N_13123,N_13447);
nor U14545 (N_14545,N_13684,N_13191);
and U14546 (N_14546,N_12606,N_13149);
and U14547 (N_14547,N_12977,N_13194);
and U14548 (N_14548,N_13470,N_12829);
or U14549 (N_14549,N_13090,N_13734);
nand U14550 (N_14550,N_12794,N_12766);
xnor U14551 (N_14551,N_12951,N_13542);
and U14552 (N_14552,N_13270,N_12542);
or U14553 (N_14553,N_13302,N_12514);
nor U14554 (N_14554,N_12944,N_13485);
and U14555 (N_14555,N_13617,N_12978);
nand U14556 (N_14556,N_13331,N_13047);
or U14557 (N_14557,N_12525,N_13449);
xor U14558 (N_14558,N_13315,N_12821);
xnor U14559 (N_14559,N_13110,N_12995);
and U14560 (N_14560,N_13319,N_12816);
or U14561 (N_14561,N_13368,N_13090);
xnor U14562 (N_14562,N_12710,N_13334);
xnor U14563 (N_14563,N_13400,N_13053);
or U14564 (N_14564,N_13332,N_13505);
xnor U14565 (N_14565,N_13617,N_13536);
nor U14566 (N_14566,N_13219,N_13724);
nand U14567 (N_14567,N_12626,N_13279);
or U14568 (N_14568,N_13020,N_13571);
or U14569 (N_14569,N_12871,N_13473);
and U14570 (N_14570,N_13571,N_13098);
xnor U14571 (N_14571,N_12531,N_12754);
and U14572 (N_14572,N_12505,N_12631);
and U14573 (N_14573,N_12779,N_12892);
nand U14574 (N_14574,N_13312,N_12904);
nor U14575 (N_14575,N_13513,N_12844);
and U14576 (N_14576,N_13529,N_13038);
nor U14577 (N_14577,N_12772,N_12739);
or U14578 (N_14578,N_13422,N_13127);
xor U14579 (N_14579,N_13070,N_13092);
or U14580 (N_14580,N_13213,N_13279);
xor U14581 (N_14581,N_13251,N_13430);
nand U14582 (N_14582,N_13650,N_13748);
xnor U14583 (N_14583,N_12910,N_13453);
xor U14584 (N_14584,N_12869,N_12870);
nor U14585 (N_14585,N_13134,N_13240);
nor U14586 (N_14586,N_13281,N_13510);
nor U14587 (N_14587,N_12784,N_12521);
xor U14588 (N_14588,N_12995,N_12589);
nand U14589 (N_14589,N_13055,N_13081);
nand U14590 (N_14590,N_12921,N_13400);
xnor U14591 (N_14591,N_12577,N_13362);
and U14592 (N_14592,N_12526,N_12945);
or U14593 (N_14593,N_13573,N_13280);
xnor U14594 (N_14594,N_13189,N_13267);
xor U14595 (N_14595,N_13136,N_13220);
nor U14596 (N_14596,N_13401,N_13217);
nand U14597 (N_14597,N_13454,N_12978);
xnor U14598 (N_14598,N_12547,N_12607);
or U14599 (N_14599,N_13144,N_12987);
nor U14600 (N_14600,N_13065,N_13544);
xnor U14601 (N_14601,N_13277,N_12927);
and U14602 (N_14602,N_13095,N_12722);
and U14603 (N_14603,N_12508,N_12724);
or U14604 (N_14604,N_13193,N_13083);
xor U14605 (N_14605,N_12805,N_13411);
and U14606 (N_14606,N_12615,N_13110);
nor U14607 (N_14607,N_12952,N_13718);
xor U14608 (N_14608,N_13175,N_12563);
xor U14609 (N_14609,N_12834,N_12911);
xor U14610 (N_14610,N_12892,N_13166);
or U14611 (N_14611,N_13014,N_13732);
and U14612 (N_14612,N_12730,N_13150);
nor U14613 (N_14613,N_12858,N_12774);
and U14614 (N_14614,N_13573,N_13463);
nand U14615 (N_14615,N_12722,N_12692);
nand U14616 (N_14616,N_12690,N_13504);
or U14617 (N_14617,N_12719,N_13102);
nor U14618 (N_14618,N_13266,N_13123);
nand U14619 (N_14619,N_13279,N_13215);
and U14620 (N_14620,N_13314,N_12599);
or U14621 (N_14621,N_13138,N_12769);
xnor U14622 (N_14622,N_13089,N_12882);
or U14623 (N_14623,N_13559,N_12610);
nand U14624 (N_14624,N_12690,N_13228);
nor U14625 (N_14625,N_12924,N_13651);
nand U14626 (N_14626,N_13086,N_13703);
or U14627 (N_14627,N_13095,N_12670);
xor U14628 (N_14628,N_12899,N_12987);
or U14629 (N_14629,N_13489,N_12564);
xor U14630 (N_14630,N_13454,N_12518);
and U14631 (N_14631,N_13402,N_12661);
xnor U14632 (N_14632,N_12581,N_12849);
xor U14633 (N_14633,N_13206,N_12619);
or U14634 (N_14634,N_12537,N_12733);
and U14635 (N_14635,N_12715,N_12854);
nand U14636 (N_14636,N_12753,N_12789);
and U14637 (N_14637,N_12667,N_13605);
xor U14638 (N_14638,N_12726,N_12969);
and U14639 (N_14639,N_13497,N_13341);
or U14640 (N_14640,N_13484,N_13011);
or U14641 (N_14641,N_12702,N_13018);
or U14642 (N_14642,N_13234,N_13325);
nor U14643 (N_14643,N_12513,N_12827);
xnor U14644 (N_14644,N_12986,N_12996);
or U14645 (N_14645,N_13302,N_13003);
and U14646 (N_14646,N_13546,N_12970);
nand U14647 (N_14647,N_13339,N_12744);
and U14648 (N_14648,N_12766,N_13381);
and U14649 (N_14649,N_13468,N_12741);
xnor U14650 (N_14650,N_13712,N_13488);
and U14651 (N_14651,N_13301,N_12579);
or U14652 (N_14652,N_13328,N_12621);
xnor U14653 (N_14653,N_12728,N_13052);
or U14654 (N_14654,N_12974,N_12784);
xnor U14655 (N_14655,N_13464,N_13487);
or U14656 (N_14656,N_12846,N_12595);
nor U14657 (N_14657,N_13500,N_13265);
or U14658 (N_14658,N_13747,N_13478);
and U14659 (N_14659,N_13504,N_12530);
or U14660 (N_14660,N_12517,N_12671);
and U14661 (N_14661,N_12773,N_12927);
xor U14662 (N_14662,N_13716,N_13352);
xor U14663 (N_14663,N_12580,N_13288);
nand U14664 (N_14664,N_13586,N_13007);
nand U14665 (N_14665,N_12762,N_13512);
nor U14666 (N_14666,N_13162,N_12729);
or U14667 (N_14667,N_12960,N_13629);
and U14668 (N_14668,N_13449,N_13383);
or U14669 (N_14669,N_12657,N_12807);
and U14670 (N_14670,N_12855,N_13685);
nor U14671 (N_14671,N_13584,N_12755);
or U14672 (N_14672,N_12716,N_12670);
or U14673 (N_14673,N_13471,N_13109);
or U14674 (N_14674,N_12576,N_13088);
nor U14675 (N_14675,N_12866,N_12983);
xnor U14676 (N_14676,N_13029,N_12711);
xnor U14677 (N_14677,N_13270,N_12621);
nand U14678 (N_14678,N_12892,N_13204);
and U14679 (N_14679,N_13367,N_13045);
nor U14680 (N_14680,N_12940,N_13264);
nand U14681 (N_14681,N_12798,N_12525);
xor U14682 (N_14682,N_13725,N_12713);
or U14683 (N_14683,N_12861,N_12922);
xnor U14684 (N_14684,N_13328,N_13201);
and U14685 (N_14685,N_13716,N_13535);
xnor U14686 (N_14686,N_12992,N_13536);
and U14687 (N_14687,N_12938,N_12612);
and U14688 (N_14688,N_12725,N_13410);
xnor U14689 (N_14689,N_12689,N_13102);
xnor U14690 (N_14690,N_13274,N_13240);
nor U14691 (N_14691,N_13275,N_13739);
or U14692 (N_14692,N_13712,N_12752);
and U14693 (N_14693,N_13055,N_13044);
and U14694 (N_14694,N_13135,N_13697);
nand U14695 (N_14695,N_13063,N_13572);
and U14696 (N_14696,N_13443,N_13279);
xor U14697 (N_14697,N_13124,N_13279);
nor U14698 (N_14698,N_12636,N_13114);
xnor U14699 (N_14699,N_13548,N_13398);
or U14700 (N_14700,N_13705,N_13022);
nand U14701 (N_14701,N_12508,N_13267);
nand U14702 (N_14702,N_12717,N_13181);
xnor U14703 (N_14703,N_12679,N_13687);
xnor U14704 (N_14704,N_13390,N_13417);
and U14705 (N_14705,N_13566,N_12728);
and U14706 (N_14706,N_12797,N_13189);
nand U14707 (N_14707,N_13676,N_13534);
xnor U14708 (N_14708,N_12712,N_12940);
and U14709 (N_14709,N_12594,N_12604);
and U14710 (N_14710,N_12627,N_13672);
nand U14711 (N_14711,N_12781,N_13313);
xor U14712 (N_14712,N_12562,N_12791);
and U14713 (N_14713,N_13369,N_13001);
nand U14714 (N_14714,N_13237,N_13346);
nor U14715 (N_14715,N_12763,N_13125);
nand U14716 (N_14716,N_13237,N_12705);
xnor U14717 (N_14717,N_12771,N_13465);
or U14718 (N_14718,N_12721,N_12810);
or U14719 (N_14719,N_12537,N_13600);
xor U14720 (N_14720,N_13018,N_13265);
nor U14721 (N_14721,N_12737,N_13126);
nor U14722 (N_14722,N_13669,N_13151);
or U14723 (N_14723,N_13500,N_13734);
nand U14724 (N_14724,N_13627,N_13424);
and U14725 (N_14725,N_13687,N_13412);
xor U14726 (N_14726,N_13511,N_13348);
or U14727 (N_14727,N_12817,N_13082);
or U14728 (N_14728,N_13109,N_13734);
xor U14729 (N_14729,N_12705,N_13599);
nand U14730 (N_14730,N_12590,N_13002);
or U14731 (N_14731,N_12723,N_13524);
and U14732 (N_14732,N_12931,N_13577);
xor U14733 (N_14733,N_13201,N_12527);
nor U14734 (N_14734,N_12760,N_12548);
nand U14735 (N_14735,N_13458,N_13064);
nand U14736 (N_14736,N_12923,N_13101);
and U14737 (N_14737,N_13005,N_12983);
and U14738 (N_14738,N_13567,N_12702);
nor U14739 (N_14739,N_13009,N_12603);
or U14740 (N_14740,N_13416,N_13357);
xnor U14741 (N_14741,N_12699,N_13309);
xnor U14742 (N_14742,N_12735,N_12601);
and U14743 (N_14743,N_12523,N_13104);
nor U14744 (N_14744,N_13249,N_13131);
nor U14745 (N_14745,N_12855,N_12671);
or U14746 (N_14746,N_13594,N_12670);
or U14747 (N_14747,N_13668,N_12770);
and U14748 (N_14748,N_13148,N_13157);
and U14749 (N_14749,N_13606,N_12533);
nor U14750 (N_14750,N_13669,N_13383);
and U14751 (N_14751,N_12528,N_13434);
nor U14752 (N_14752,N_12868,N_12778);
or U14753 (N_14753,N_13180,N_13462);
and U14754 (N_14754,N_12977,N_13410);
xnor U14755 (N_14755,N_13274,N_13419);
and U14756 (N_14756,N_13562,N_13662);
nor U14757 (N_14757,N_13460,N_13540);
and U14758 (N_14758,N_13592,N_12826);
or U14759 (N_14759,N_13732,N_13617);
nand U14760 (N_14760,N_12670,N_12555);
xor U14761 (N_14761,N_13138,N_13038);
xnor U14762 (N_14762,N_13387,N_12934);
xor U14763 (N_14763,N_12719,N_13736);
or U14764 (N_14764,N_13017,N_12813);
nand U14765 (N_14765,N_13386,N_13646);
nor U14766 (N_14766,N_13440,N_12893);
nor U14767 (N_14767,N_12945,N_12857);
or U14768 (N_14768,N_13387,N_12654);
nand U14769 (N_14769,N_12856,N_12692);
nand U14770 (N_14770,N_12734,N_12686);
and U14771 (N_14771,N_12778,N_13637);
and U14772 (N_14772,N_12640,N_12961);
xnor U14773 (N_14773,N_13685,N_12663);
or U14774 (N_14774,N_12830,N_13554);
or U14775 (N_14775,N_12874,N_12596);
and U14776 (N_14776,N_13103,N_13303);
and U14777 (N_14777,N_13096,N_13436);
nor U14778 (N_14778,N_12744,N_13031);
and U14779 (N_14779,N_13522,N_13455);
or U14780 (N_14780,N_12521,N_12918);
xor U14781 (N_14781,N_13533,N_12912);
nand U14782 (N_14782,N_13173,N_12954);
nand U14783 (N_14783,N_12715,N_13426);
xnor U14784 (N_14784,N_13262,N_12544);
or U14785 (N_14785,N_12668,N_12860);
and U14786 (N_14786,N_13252,N_13748);
xnor U14787 (N_14787,N_12777,N_12956);
and U14788 (N_14788,N_13266,N_13322);
and U14789 (N_14789,N_12907,N_13732);
nor U14790 (N_14790,N_12737,N_12794);
or U14791 (N_14791,N_13107,N_12586);
or U14792 (N_14792,N_12861,N_12698);
or U14793 (N_14793,N_13549,N_12677);
nor U14794 (N_14794,N_13563,N_13244);
and U14795 (N_14795,N_13384,N_13424);
and U14796 (N_14796,N_13236,N_12651);
nand U14797 (N_14797,N_13134,N_12773);
xor U14798 (N_14798,N_12950,N_13032);
nand U14799 (N_14799,N_12609,N_13605);
or U14800 (N_14800,N_12729,N_13010);
nor U14801 (N_14801,N_12597,N_13348);
and U14802 (N_14802,N_12969,N_12505);
and U14803 (N_14803,N_12612,N_12500);
and U14804 (N_14804,N_12507,N_13706);
xor U14805 (N_14805,N_13608,N_13298);
nand U14806 (N_14806,N_13474,N_13092);
xnor U14807 (N_14807,N_13090,N_13076);
nand U14808 (N_14808,N_13643,N_13429);
and U14809 (N_14809,N_13689,N_13074);
or U14810 (N_14810,N_13318,N_13326);
nand U14811 (N_14811,N_12891,N_13332);
nand U14812 (N_14812,N_13724,N_12906);
xor U14813 (N_14813,N_12522,N_12532);
and U14814 (N_14814,N_13435,N_13378);
and U14815 (N_14815,N_13143,N_13254);
and U14816 (N_14816,N_13203,N_12738);
or U14817 (N_14817,N_13445,N_12617);
or U14818 (N_14818,N_13389,N_12768);
xor U14819 (N_14819,N_13100,N_13448);
nand U14820 (N_14820,N_12817,N_13490);
xor U14821 (N_14821,N_13720,N_13143);
xor U14822 (N_14822,N_12764,N_12873);
nor U14823 (N_14823,N_12958,N_12991);
and U14824 (N_14824,N_12819,N_13314);
xnor U14825 (N_14825,N_13551,N_13316);
nand U14826 (N_14826,N_13033,N_13323);
and U14827 (N_14827,N_13359,N_12895);
nand U14828 (N_14828,N_13196,N_13280);
nand U14829 (N_14829,N_12556,N_13060);
nor U14830 (N_14830,N_12994,N_13614);
xor U14831 (N_14831,N_12630,N_12583);
or U14832 (N_14832,N_12767,N_12932);
or U14833 (N_14833,N_13283,N_13734);
or U14834 (N_14834,N_12592,N_13078);
xor U14835 (N_14835,N_13497,N_12950);
nor U14836 (N_14836,N_13465,N_13140);
xor U14837 (N_14837,N_12544,N_12909);
xor U14838 (N_14838,N_13287,N_13436);
xnor U14839 (N_14839,N_12955,N_12783);
nand U14840 (N_14840,N_12622,N_13213);
or U14841 (N_14841,N_13321,N_12698);
xor U14842 (N_14842,N_12980,N_12774);
and U14843 (N_14843,N_13207,N_12514);
nand U14844 (N_14844,N_12842,N_12747);
xnor U14845 (N_14845,N_12577,N_13586);
xnor U14846 (N_14846,N_13235,N_12912);
and U14847 (N_14847,N_13321,N_13523);
or U14848 (N_14848,N_12943,N_13478);
or U14849 (N_14849,N_13247,N_13042);
nor U14850 (N_14850,N_13603,N_12689);
xor U14851 (N_14851,N_13341,N_13176);
nand U14852 (N_14852,N_13356,N_13465);
nand U14853 (N_14853,N_13006,N_13452);
nor U14854 (N_14854,N_13538,N_13530);
xnor U14855 (N_14855,N_13111,N_13397);
nor U14856 (N_14856,N_12833,N_13698);
nor U14857 (N_14857,N_12879,N_12882);
xor U14858 (N_14858,N_12993,N_13500);
nand U14859 (N_14859,N_13440,N_12806);
xnor U14860 (N_14860,N_13358,N_13188);
xnor U14861 (N_14861,N_13001,N_13066);
nor U14862 (N_14862,N_13077,N_13562);
nor U14863 (N_14863,N_13348,N_12598);
or U14864 (N_14864,N_12792,N_12999);
xor U14865 (N_14865,N_13380,N_13367);
or U14866 (N_14866,N_12667,N_12673);
and U14867 (N_14867,N_13011,N_13286);
nor U14868 (N_14868,N_13403,N_13053);
or U14869 (N_14869,N_13520,N_13641);
and U14870 (N_14870,N_13047,N_13239);
or U14871 (N_14871,N_13601,N_13709);
nand U14872 (N_14872,N_13486,N_13186);
and U14873 (N_14873,N_13542,N_12775);
and U14874 (N_14874,N_12988,N_12670);
nor U14875 (N_14875,N_12858,N_13526);
nand U14876 (N_14876,N_13519,N_12584);
and U14877 (N_14877,N_13588,N_13127);
nor U14878 (N_14878,N_13723,N_12841);
or U14879 (N_14879,N_12650,N_13511);
xnor U14880 (N_14880,N_13363,N_13699);
xor U14881 (N_14881,N_12933,N_12530);
nand U14882 (N_14882,N_12918,N_13495);
and U14883 (N_14883,N_12697,N_12899);
or U14884 (N_14884,N_13348,N_12617);
and U14885 (N_14885,N_12941,N_12963);
nand U14886 (N_14886,N_12934,N_13737);
nand U14887 (N_14887,N_12818,N_13625);
or U14888 (N_14888,N_13180,N_13415);
nor U14889 (N_14889,N_12876,N_12945);
and U14890 (N_14890,N_13345,N_13507);
nor U14891 (N_14891,N_13567,N_13565);
nand U14892 (N_14892,N_12600,N_13213);
or U14893 (N_14893,N_13314,N_13672);
nand U14894 (N_14894,N_13106,N_13443);
nor U14895 (N_14895,N_13330,N_13720);
and U14896 (N_14896,N_12886,N_12728);
xor U14897 (N_14897,N_13354,N_12505);
and U14898 (N_14898,N_12671,N_12682);
xor U14899 (N_14899,N_13004,N_12655);
and U14900 (N_14900,N_12509,N_13455);
xor U14901 (N_14901,N_13529,N_12998);
or U14902 (N_14902,N_12689,N_13601);
nand U14903 (N_14903,N_12929,N_12868);
and U14904 (N_14904,N_13613,N_13287);
nand U14905 (N_14905,N_13189,N_13574);
and U14906 (N_14906,N_13633,N_13614);
nand U14907 (N_14907,N_13282,N_13294);
nand U14908 (N_14908,N_13067,N_12973);
or U14909 (N_14909,N_12705,N_13696);
nor U14910 (N_14910,N_12587,N_13591);
nor U14911 (N_14911,N_12933,N_13047);
xnor U14912 (N_14912,N_13168,N_13030);
nand U14913 (N_14913,N_13514,N_13093);
nor U14914 (N_14914,N_13472,N_13227);
xor U14915 (N_14915,N_13156,N_12698);
xnor U14916 (N_14916,N_12835,N_12925);
xnor U14917 (N_14917,N_13543,N_12922);
and U14918 (N_14918,N_13735,N_12897);
xor U14919 (N_14919,N_13626,N_13464);
and U14920 (N_14920,N_13294,N_13210);
xor U14921 (N_14921,N_12936,N_13536);
nor U14922 (N_14922,N_13735,N_12649);
nand U14923 (N_14923,N_13211,N_12689);
nor U14924 (N_14924,N_12646,N_12964);
or U14925 (N_14925,N_12817,N_13416);
xor U14926 (N_14926,N_13455,N_12553);
nor U14927 (N_14927,N_13205,N_13141);
and U14928 (N_14928,N_13209,N_12509);
nor U14929 (N_14929,N_13334,N_13072);
nand U14930 (N_14930,N_12737,N_12913);
xor U14931 (N_14931,N_13605,N_12898);
xor U14932 (N_14932,N_13607,N_12529);
and U14933 (N_14933,N_12833,N_12510);
nand U14934 (N_14934,N_13258,N_13745);
nor U14935 (N_14935,N_13528,N_13524);
nor U14936 (N_14936,N_12969,N_13100);
and U14937 (N_14937,N_13731,N_12800);
nand U14938 (N_14938,N_13502,N_12753);
xor U14939 (N_14939,N_13185,N_13695);
xor U14940 (N_14940,N_12784,N_12537);
nand U14941 (N_14941,N_13019,N_13656);
and U14942 (N_14942,N_13687,N_12904);
nand U14943 (N_14943,N_13304,N_12961);
and U14944 (N_14944,N_12578,N_12947);
nand U14945 (N_14945,N_13409,N_12973);
nand U14946 (N_14946,N_12639,N_13384);
and U14947 (N_14947,N_12983,N_13421);
and U14948 (N_14948,N_13602,N_13470);
or U14949 (N_14949,N_13575,N_12620);
xor U14950 (N_14950,N_12725,N_12779);
or U14951 (N_14951,N_13678,N_13573);
and U14952 (N_14952,N_13378,N_13059);
nor U14953 (N_14953,N_12502,N_13457);
or U14954 (N_14954,N_13080,N_12579);
xor U14955 (N_14955,N_13097,N_13595);
nor U14956 (N_14956,N_13432,N_13014);
and U14957 (N_14957,N_13060,N_12804);
and U14958 (N_14958,N_12973,N_13392);
nand U14959 (N_14959,N_12876,N_13022);
and U14960 (N_14960,N_12891,N_13532);
xnor U14961 (N_14961,N_12643,N_13410);
nor U14962 (N_14962,N_12930,N_13380);
nor U14963 (N_14963,N_13186,N_13278);
xor U14964 (N_14964,N_12526,N_13163);
xor U14965 (N_14965,N_12518,N_13502);
xnor U14966 (N_14966,N_12890,N_12848);
and U14967 (N_14967,N_12552,N_12792);
or U14968 (N_14968,N_13390,N_13010);
nand U14969 (N_14969,N_13137,N_13013);
nor U14970 (N_14970,N_13405,N_13045);
and U14971 (N_14971,N_13633,N_13224);
or U14972 (N_14972,N_13099,N_12625);
xnor U14973 (N_14973,N_13269,N_13121);
xor U14974 (N_14974,N_12824,N_13314);
nand U14975 (N_14975,N_13286,N_13372);
or U14976 (N_14976,N_13482,N_12568);
or U14977 (N_14977,N_13349,N_13216);
nor U14978 (N_14978,N_13261,N_13247);
and U14979 (N_14979,N_12817,N_13578);
nor U14980 (N_14980,N_12996,N_13030);
nor U14981 (N_14981,N_12627,N_13112);
nor U14982 (N_14982,N_13202,N_13325);
nor U14983 (N_14983,N_13000,N_13265);
and U14984 (N_14984,N_13539,N_12580);
nor U14985 (N_14985,N_13300,N_13633);
nand U14986 (N_14986,N_13202,N_13313);
nor U14987 (N_14987,N_13405,N_12858);
and U14988 (N_14988,N_13445,N_13712);
nor U14989 (N_14989,N_12717,N_13341);
xnor U14990 (N_14990,N_12715,N_12898);
or U14991 (N_14991,N_13074,N_12618);
xor U14992 (N_14992,N_12516,N_13645);
or U14993 (N_14993,N_13105,N_12786);
nor U14994 (N_14994,N_12763,N_12847);
nand U14995 (N_14995,N_12883,N_12843);
nor U14996 (N_14996,N_13546,N_13377);
nor U14997 (N_14997,N_13355,N_12813);
nor U14998 (N_14998,N_12741,N_13056);
nand U14999 (N_14999,N_13480,N_13149);
or U15000 (N_15000,N_14648,N_14840);
or U15001 (N_15001,N_14735,N_14704);
xor U15002 (N_15002,N_14792,N_14270);
xor U15003 (N_15003,N_14089,N_14920);
xor U15004 (N_15004,N_13889,N_14467);
or U15005 (N_15005,N_13888,N_13960);
or U15006 (N_15006,N_13971,N_14204);
nand U15007 (N_15007,N_14371,N_14635);
and U15008 (N_15008,N_14520,N_13817);
xnor U15009 (N_15009,N_14340,N_13824);
and U15010 (N_15010,N_13954,N_14529);
xnor U15011 (N_15011,N_14317,N_14572);
or U15012 (N_15012,N_14713,N_13859);
and U15013 (N_15013,N_13987,N_14322);
and U15014 (N_15014,N_14381,N_14212);
xnor U15015 (N_15015,N_13986,N_14856);
nand U15016 (N_15016,N_13810,N_14372);
or U15017 (N_15017,N_14911,N_13899);
xor U15018 (N_15018,N_13957,N_14726);
nand U15019 (N_15019,N_14403,N_14951);
xnor U15020 (N_15020,N_14669,N_14846);
and U15021 (N_15021,N_14473,N_14422);
or U15022 (N_15022,N_14875,N_14079);
xor U15023 (N_15023,N_13902,N_14607);
or U15024 (N_15024,N_14525,N_14755);
or U15025 (N_15025,N_14578,N_14729);
xnor U15026 (N_15026,N_13760,N_14072);
nor U15027 (N_15027,N_14143,N_14182);
and U15028 (N_15028,N_14860,N_14048);
nand U15029 (N_15029,N_14181,N_14560);
or U15030 (N_15030,N_14436,N_14230);
xnor U15031 (N_15031,N_13928,N_14698);
nand U15032 (N_15032,N_14598,N_13794);
nor U15033 (N_15033,N_14519,N_14991);
nand U15034 (N_15034,N_14250,N_13882);
xor U15035 (N_15035,N_14831,N_14099);
nand U15036 (N_15036,N_14214,N_14108);
nor U15037 (N_15037,N_13828,N_14731);
nor U15038 (N_15038,N_14368,N_14500);
xnor U15039 (N_15039,N_14833,N_13929);
nand U15040 (N_15040,N_14565,N_14853);
xnor U15041 (N_15041,N_14925,N_14195);
xnor U15042 (N_15042,N_13913,N_13895);
or U15043 (N_15043,N_14427,N_14061);
and U15044 (N_15044,N_14254,N_14142);
nand U15045 (N_15045,N_14216,N_14398);
nand U15046 (N_15046,N_14998,N_14556);
nand U15047 (N_15047,N_14288,N_13801);
xnor U15048 (N_15048,N_14101,N_13792);
or U15049 (N_15049,N_13967,N_13784);
or U15050 (N_15050,N_14721,N_14830);
nor U15051 (N_15051,N_14834,N_14953);
or U15052 (N_15052,N_14197,N_14802);
nand U15053 (N_15053,N_14878,N_13941);
nor U15054 (N_15054,N_14779,N_14743);
and U15055 (N_15055,N_14417,N_14010);
and U15056 (N_15056,N_14754,N_14468);
nand U15057 (N_15057,N_14313,N_13800);
xnor U15058 (N_15058,N_13822,N_14765);
nor U15059 (N_15059,N_13762,N_14955);
nand U15060 (N_15060,N_14043,N_14431);
nor U15061 (N_15061,N_13809,N_14872);
and U15062 (N_15062,N_14085,N_14518);
nand U15063 (N_15063,N_14155,N_14818);
nor U15064 (N_15064,N_14366,N_14235);
or U15065 (N_15065,N_13980,N_14377);
or U15066 (N_15066,N_14458,N_14133);
and U15067 (N_15067,N_13972,N_14352);
nand U15068 (N_15068,N_13846,N_14938);
xor U15069 (N_15069,N_14348,N_13921);
nor U15070 (N_15070,N_13799,N_14475);
or U15071 (N_15071,N_13862,N_14655);
nor U15072 (N_15072,N_14476,N_14927);
xnor U15073 (N_15073,N_14764,N_13778);
or U15074 (N_15074,N_13780,N_14461);
nand U15075 (N_15075,N_14609,N_14287);
xor U15076 (N_15076,N_14022,N_14205);
nor U15077 (N_15077,N_14612,N_14209);
nand U15078 (N_15078,N_14169,N_13942);
xnor U15079 (N_15079,N_14527,N_13819);
and U15080 (N_15080,N_14027,N_13898);
nor U15081 (N_15081,N_14160,N_14429);
nand U15082 (N_15082,N_14453,N_14187);
xor U15083 (N_15083,N_13861,N_14257);
or U15084 (N_15084,N_14817,N_14739);
nor U15085 (N_15085,N_13992,N_14023);
xor U15086 (N_15086,N_14460,N_14396);
nand U15087 (N_15087,N_14781,N_14662);
nand U15088 (N_15088,N_14981,N_14516);
and U15089 (N_15089,N_14326,N_14865);
xor U15090 (N_15090,N_13901,N_14244);
xnor U15091 (N_15091,N_14379,N_13985);
and U15092 (N_15092,N_14931,N_14213);
nor U15093 (N_15093,N_14630,N_13871);
or U15094 (N_15094,N_14537,N_13943);
xnor U15095 (N_15095,N_14871,N_14986);
nor U15096 (N_15096,N_14354,N_14892);
and U15097 (N_15097,N_14933,N_14447);
nor U15098 (N_15098,N_14245,N_14004);
or U15099 (N_15099,N_13791,N_14869);
nor U15100 (N_15100,N_13878,N_14102);
nor U15101 (N_15101,N_14905,N_14876);
or U15102 (N_15102,N_14693,N_13850);
and U15103 (N_15103,N_14418,N_14080);
xor U15104 (N_15104,N_14059,N_14423);
nand U15105 (N_15105,N_13785,N_14671);
nand U15106 (N_15106,N_14954,N_14980);
nor U15107 (N_15107,N_14452,N_14442);
nand U15108 (N_15108,N_14232,N_13830);
nand U15109 (N_15109,N_14758,N_14446);
and U15110 (N_15110,N_13788,N_14845);
nor U15111 (N_15111,N_14813,N_14026);
or U15112 (N_15112,N_14822,N_14260);
and U15113 (N_15113,N_13781,N_14394);
nor U15114 (N_15114,N_14641,N_13876);
or U15115 (N_15115,N_14801,N_14686);
nor U15116 (N_15116,N_14820,N_14271);
nand U15117 (N_15117,N_14140,N_14046);
or U15118 (N_15118,N_13793,N_14355);
xnor U15119 (N_15119,N_14972,N_14626);
xor U15120 (N_15120,N_13803,N_14137);
or U15121 (N_15121,N_14185,N_14974);
or U15122 (N_15122,N_14649,N_14316);
or U15123 (N_15123,N_14657,N_14740);
xor U15124 (N_15124,N_14367,N_14888);
and U15125 (N_15125,N_14123,N_14310);
or U15126 (N_15126,N_14877,N_14795);
or U15127 (N_15127,N_13961,N_14741);
or U15128 (N_15128,N_14742,N_14425);
xnor U15129 (N_15129,N_14324,N_13877);
xor U15130 (N_15130,N_13969,N_13843);
nand U15131 (N_15131,N_14748,N_14522);
xor U15132 (N_15132,N_14177,N_13886);
nor U15133 (N_15133,N_14485,N_14351);
nand U15134 (N_15134,N_14750,N_13756);
xnor U15135 (N_15135,N_13867,N_14689);
nand U15136 (N_15136,N_14001,N_14575);
and U15137 (N_15137,N_13797,N_14589);
or U15138 (N_15138,N_14218,N_14430);
and U15139 (N_15139,N_14803,N_13770);
nand U15140 (N_15140,N_14203,N_14504);
and U15141 (N_15141,N_14999,N_14175);
xnor U15142 (N_15142,N_14658,N_14725);
or U15143 (N_15143,N_14105,N_14584);
and U15144 (N_15144,N_14733,N_13879);
or U15145 (N_15145,N_14702,N_14646);
or U15146 (N_15146,N_14756,N_14003);
or U15147 (N_15147,N_14014,N_14039);
xor U15148 (N_15148,N_13958,N_14343);
and U15149 (N_15149,N_14676,N_14496);
nor U15150 (N_15150,N_13968,N_14037);
xor U15151 (N_15151,N_14439,N_14791);
nand U15152 (N_15152,N_14361,N_14959);
and U15153 (N_15153,N_14923,N_13844);
nor U15154 (N_15154,N_14388,N_14922);
xnor U15155 (N_15155,N_14344,N_14617);
and U15156 (N_15156,N_14407,N_14499);
nand U15157 (N_15157,N_14402,N_14685);
xnor U15158 (N_15158,N_14070,N_14881);
nor U15159 (N_15159,N_14995,N_14321);
or U15160 (N_15160,N_14688,N_14252);
nor U15161 (N_15161,N_14653,N_14977);
nand U15162 (N_15162,N_14727,N_14996);
and U15163 (N_15163,N_14163,N_14488);
nor U15164 (N_15164,N_14699,N_14031);
or U15165 (N_15165,N_13914,N_14277);
xor U15166 (N_15166,N_14613,N_13955);
xnor U15167 (N_15167,N_14154,N_14349);
and U15168 (N_15168,N_14514,N_14526);
or U15169 (N_15169,N_14406,N_14957);
nand U15170 (N_15170,N_14835,N_14867);
xor U15171 (N_15171,N_14369,N_14749);
xor U15172 (N_15172,N_13779,N_14414);
nor U15173 (N_15173,N_14608,N_14434);
and U15174 (N_15174,N_14814,N_14255);
or U15175 (N_15175,N_14021,N_13912);
nor U15176 (N_15176,N_14563,N_14507);
and U15177 (N_15177,N_14844,N_14283);
nor U15178 (N_15178,N_14062,N_14211);
nand U15179 (N_15179,N_14645,N_14486);
nand U15180 (N_15180,N_14353,N_14852);
and U15181 (N_15181,N_13874,N_13873);
and U15182 (N_15182,N_14292,N_14400);
and U15183 (N_15183,N_13840,N_14152);
and U15184 (N_15184,N_14561,N_14672);
and U15185 (N_15185,N_14628,N_14694);
xnor U15186 (N_15186,N_14437,N_14455);
and U15187 (N_15187,N_13757,N_14828);
nand U15188 (N_15188,N_14586,N_14224);
xor U15189 (N_15189,N_14126,N_14106);
nor U15190 (N_15190,N_14454,N_13996);
nand U15191 (N_15191,N_14640,N_14378);
nand U15192 (N_15192,N_14231,N_14597);
nand U15193 (N_15193,N_13923,N_13755);
or U15194 (N_15194,N_13988,N_14308);
nor U15195 (N_15195,N_14375,N_14604);
nand U15196 (N_15196,N_14930,N_14335);
and U15197 (N_15197,N_14769,N_13906);
xor U15198 (N_15198,N_14839,N_14370);
and U15199 (N_15199,N_14248,N_14842);
and U15200 (N_15200,N_14908,N_14789);
nor U15201 (N_15201,N_14243,N_14363);
nand U15202 (N_15202,N_14189,N_14161);
xor U15203 (N_15203,N_13835,N_14816);
and U15204 (N_15204,N_14706,N_14338);
nor U15205 (N_15205,N_14790,N_13764);
xor U15206 (N_15206,N_14111,N_14052);
xnor U15207 (N_15207,N_13870,N_14280);
and U15208 (N_15208,N_13887,N_14552);
xnor U15209 (N_15209,N_14502,N_14234);
nor U15210 (N_15210,N_14002,N_13920);
and U15211 (N_15211,N_13787,N_13752);
nand U15212 (N_15212,N_14777,N_14896);
or U15213 (N_15213,N_14973,N_14494);
nor U15214 (N_15214,N_14705,N_14602);
nand U15215 (N_15215,N_14510,N_14943);
nor U15216 (N_15216,N_14531,N_14637);
and U15217 (N_15217,N_14557,N_14171);
or U15218 (N_15218,N_14787,N_13880);
nand U15219 (N_15219,N_14382,N_14821);
or U15220 (N_15220,N_13837,N_14415);
nand U15221 (N_15221,N_14498,N_14279);
nor U15222 (N_15222,N_14391,N_14827);
nand U15223 (N_15223,N_13808,N_14376);
or U15224 (N_15224,N_13991,N_14895);
nand U15225 (N_15225,N_14438,N_14360);
or U15226 (N_15226,N_14687,N_14697);
nand U15227 (N_15227,N_14904,N_14483);
nand U15228 (N_15228,N_14334,N_14709);
nor U15229 (N_15229,N_14100,N_14493);
xor U15230 (N_15230,N_14005,N_14906);
xnor U15231 (N_15231,N_14413,N_14544);
xnor U15232 (N_15232,N_14675,N_14681);
and U15233 (N_15233,N_14650,N_14952);
and U15234 (N_15234,N_13807,N_14884);
or U15235 (N_15235,N_13910,N_14985);
xor U15236 (N_15236,N_14112,N_14534);
nor U15237 (N_15237,N_14747,N_14456);
xnor U15238 (N_15238,N_14619,N_14157);
or U15239 (N_15239,N_13798,N_13811);
nor U15240 (N_15240,N_13919,N_13982);
xor U15241 (N_15241,N_14673,N_14759);
nor U15242 (N_15242,N_14859,N_13926);
xor U15243 (N_15243,N_13860,N_14633);
nand U15244 (N_15244,N_13815,N_14139);
and U15245 (N_15245,N_14264,N_14843);
nand U15246 (N_15246,N_14121,N_14517);
or U15247 (N_15247,N_14785,N_14215);
and U15248 (N_15248,N_13813,N_14356);
or U15249 (N_15249,N_13984,N_14129);
nor U15250 (N_15250,N_14549,N_13766);
nand U15251 (N_15251,N_14558,N_14590);
or U15252 (N_15252,N_13818,N_14192);
xor U15253 (N_15253,N_14384,N_13806);
or U15254 (N_15254,N_14007,N_14629);
xor U15255 (N_15255,N_13900,N_14329);
and U15256 (N_15256,N_14325,N_14466);
nand U15257 (N_15257,N_14523,N_14011);
nor U15258 (N_15258,N_14815,N_14994);
or U15259 (N_15259,N_14285,N_14424);
and U15260 (N_15260,N_14236,N_14113);
and U15261 (N_15261,N_13790,N_14762);
or U15262 (N_15262,N_14956,N_14910);
xor U15263 (N_15263,N_14772,N_13977);
or U15264 (N_15264,N_14303,N_14855);
xor U15265 (N_15265,N_14849,N_14937);
nand U15266 (N_15266,N_14753,N_14495);
or U15267 (N_15267,N_14806,N_14201);
nor U15268 (N_15268,N_14272,N_13881);
and U15269 (N_15269,N_14190,N_14393);
and U15270 (N_15270,N_13930,N_14577);
nand U15271 (N_15271,N_14041,N_14678);
or U15272 (N_15272,N_14069,N_13946);
xor U15273 (N_15273,N_14247,N_14847);
nand U15274 (N_15274,N_13863,N_14684);
and U15275 (N_15275,N_14282,N_14767);
and U15276 (N_15276,N_14778,N_13976);
or U15277 (N_15277,N_13868,N_14576);
nand U15278 (N_15278,N_14179,N_14385);
or U15279 (N_15279,N_14807,N_14020);
nor U15280 (N_15280,N_13847,N_14259);
or U15281 (N_15281,N_14744,N_13759);
nand U15282 (N_15282,N_13816,N_14315);
nor U15283 (N_15283,N_13849,N_14297);
xnor U15284 (N_15284,N_13981,N_14532);
nand U15285 (N_15285,N_14104,N_14885);
nand U15286 (N_15286,N_14851,N_13927);
and U15287 (N_15287,N_13885,N_14265);
nor U15288 (N_15288,N_14773,N_13924);
or U15289 (N_15289,N_13965,N_13833);
xor U15290 (N_15290,N_14081,N_14131);
nor U15291 (N_15291,N_13953,N_14470);
or U15292 (N_15292,N_14492,N_13872);
nand U15293 (N_15293,N_14012,N_14331);
nand U15294 (N_15294,N_14408,N_14314);
or U15295 (N_15295,N_14900,N_13777);
nand U15296 (N_15296,N_14284,N_13820);
nor U15297 (N_15297,N_14419,N_14599);
or U15298 (N_15298,N_13856,N_14964);
and U15299 (N_15299,N_14605,N_14667);
nor U15300 (N_15300,N_13962,N_14909);
xnor U15301 (N_15301,N_13936,N_13812);
or U15302 (N_15302,N_14595,N_14226);
xnor U15303 (N_15303,N_13894,N_13995);
xor U15304 (N_15304,N_14950,N_14299);
nand U15305 (N_15305,N_14390,N_13964);
nand U15306 (N_15306,N_14730,N_14266);
and U15307 (N_15307,N_14191,N_14018);
and U15308 (N_15308,N_14768,N_14948);
or U15309 (N_15309,N_14554,N_14714);
nor U15310 (N_15310,N_13896,N_14965);
xnor U15311 (N_15311,N_13892,N_14788);
xnor U15312 (N_15312,N_14032,N_14319);
nor U15313 (N_15313,N_14944,N_13993);
and U15314 (N_15314,N_14125,N_14677);
and U15315 (N_15315,N_14708,N_14239);
nor U15316 (N_15316,N_14665,N_14173);
or U15317 (N_15317,N_14392,N_14634);
xor U15318 (N_15318,N_14374,N_14509);
xnor U15319 (N_15319,N_14083,N_14913);
and U15320 (N_15320,N_14281,N_14639);
nand U15321 (N_15321,N_14887,N_14336);
nand U15322 (N_15322,N_14893,N_14837);
nor U15323 (N_15323,N_14621,N_13768);
and U15324 (N_15324,N_14464,N_14533);
and U15325 (N_15325,N_14984,N_14165);
and U15326 (N_15326,N_14342,N_13829);
xnor U15327 (N_15327,N_14261,N_13997);
and U15328 (N_15328,N_13911,N_14825);
or U15329 (N_15329,N_14075,N_14302);
or U15330 (N_15330,N_14539,N_14903);
and U15331 (N_15331,N_14868,N_13866);
nand U15332 (N_15332,N_14221,N_14016);
or U15333 (N_15333,N_14548,N_13776);
xnor U15334 (N_15334,N_14760,N_14289);
nand U15335 (N_15335,N_14512,N_14134);
nor U15336 (N_15336,N_14968,N_14854);
xor U15337 (N_15337,N_14886,N_14880);
and U15338 (N_15338,N_14794,N_14120);
nor U15339 (N_15339,N_14651,N_14674);
xor U15340 (N_15340,N_14306,N_14652);
nand U15341 (N_15341,N_13821,N_13945);
xor U15342 (N_15342,N_14135,N_14094);
and U15343 (N_15343,N_14841,N_14771);
nor U15344 (N_15344,N_14463,N_13854);
nor U15345 (N_15345,N_14622,N_14793);
nand U15346 (N_15346,N_13783,N_14127);
or U15347 (N_15347,N_14208,N_14963);
and U15348 (N_15348,N_14832,N_14168);
or U15349 (N_15349,N_14044,N_13763);
and U15350 (N_15350,N_13940,N_14065);
nor U15351 (N_15351,N_14627,N_13973);
xor U15352 (N_15352,N_14618,N_14359);
nor U15353 (N_15353,N_14178,N_13802);
nand U15354 (N_15354,N_14656,N_14659);
nor U15355 (N_15355,N_14550,N_14524);
nand U15356 (N_15356,N_14276,N_14130);
or U15357 (N_15357,N_14566,N_14412);
xor U15358 (N_15358,N_14153,N_14623);
nand U15359 (N_15359,N_14696,N_14188);
and U15360 (N_15360,N_14038,N_14426);
nand U15361 (N_15361,N_13998,N_13875);
nor U15362 (N_15362,N_14907,N_13883);
xnor U15363 (N_15363,N_14411,N_14717);
nand U15364 (N_15364,N_14087,N_14217);
nand U15365 (N_15365,N_14535,N_14796);
xnor U15366 (N_15366,N_14914,N_14583);
nor U15367 (N_15367,N_14358,N_14033);
nand U15368 (N_15368,N_14757,N_13834);
and U15369 (N_15369,N_13827,N_14722);
and U15370 (N_15370,N_14588,N_14373);
nor U15371 (N_15371,N_14692,N_14233);
nor U15372 (N_15372,N_13774,N_14863);
nor U15373 (N_15373,N_14812,N_14268);
nor U15374 (N_15374,N_14311,N_13948);
xnor U15375 (N_15375,N_14625,N_14992);
nand U15376 (N_15376,N_14663,N_13934);
nand U15377 (N_15377,N_14547,N_14680);
xor U15378 (N_15378,N_14357,N_14132);
and U15379 (N_15379,N_14158,N_14946);
nor U15380 (N_15380,N_13908,N_14328);
or U15381 (N_15381,N_14976,N_14274);
xor U15382 (N_15382,N_14064,N_14294);
nor U15383 (N_15383,N_13938,N_13857);
and U15384 (N_15384,N_14858,N_13935);
nor U15385 (N_15385,N_14449,N_14958);
xor U15386 (N_15386,N_14076,N_13944);
nand U15387 (N_15387,N_13905,N_14587);
or U15388 (N_15388,N_14114,N_14082);
and U15389 (N_15389,N_14864,N_14724);
nor U15390 (N_15390,N_14862,N_14712);
xor U15391 (N_15391,N_14616,N_13864);
xnor U15392 (N_15392,N_14128,N_14275);
nand U15393 (N_15393,N_14220,N_14448);
and U15394 (N_15394,N_14989,N_14119);
nor U15395 (N_15395,N_13932,N_14136);
or U15396 (N_15396,N_14337,N_13999);
xor U15397 (N_15397,N_13823,N_14200);
nand U15398 (N_15398,N_13937,N_13917);
and U15399 (N_15399,N_14387,N_14763);
nand U15400 (N_15400,N_14715,N_14262);
xor U15401 (N_15401,N_14921,N_14180);
nor U15402 (N_15402,N_14145,N_14732);
nand U15403 (N_15403,N_13796,N_14210);
and U15404 (N_15404,N_14690,N_14484);
nand U15405 (N_15405,N_14810,N_13869);
nor U15406 (N_15406,N_13959,N_14049);
or U15407 (N_15407,N_14611,N_14766);
nor U15408 (N_15408,N_14148,N_14318);
and U15409 (N_15409,N_14567,N_14723);
nand U15410 (N_15410,N_14029,N_14737);
nand U15411 (N_15411,N_14734,N_14186);
xnor U15412 (N_15412,N_14809,N_14350);
and U15413 (N_15413,N_14603,N_14941);
nand U15414 (N_15414,N_14490,N_14477);
or U15415 (N_15415,N_14146,N_14745);
nand U15416 (N_15416,N_14571,N_14122);
or U15417 (N_15417,N_14267,N_14409);
and U15418 (N_15418,N_14278,N_14780);
xor U15419 (N_15419,N_14632,N_14241);
or U15420 (N_15420,N_14568,N_14503);
and U15421 (N_15421,N_13750,N_14078);
and U15422 (N_15422,N_14362,N_14761);
and U15423 (N_15423,N_13907,N_13772);
xnor U15424 (N_15424,N_14090,N_14183);
or U15425 (N_15425,N_14249,N_14471);
nor U15426 (N_15426,N_14253,N_14836);
or U15427 (N_15427,N_14116,N_13839);
nand U15428 (N_15428,N_13831,N_14644);
nand U15429 (N_15429,N_14746,N_14866);
or U15430 (N_15430,N_13939,N_14444);
nand U15431 (N_15431,N_14719,N_14296);
nand U15432 (N_15432,N_14115,N_14481);
or U15433 (N_15433,N_14570,N_14894);
nand U15434 (N_15434,N_14149,N_14228);
or U15435 (N_15435,N_13979,N_13814);
or U15436 (N_15436,N_14162,N_14594);
and U15437 (N_15437,N_14970,N_14932);
and U15438 (N_15438,N_14918,N_14117);
or U15439 (N_15439,N_14600,N_14929);
or U15440 (N_15440,N_13842,N_13775);
nand U15441 (N_15441,N_14988,N_14497);
nand U15442 (N_15442,N_14770,N_14615);
and U15443 (N_15443,N_14960,N_14530);
xor U15444 (N_15444,N_13845,N_14330);
xor U15445 (N_15445,N_13893,N_14462);
or U15446 (N_15446,N_14898,N_14874);
nor U15447 (N_15447,N_14664,N_14819);
and U15448 (N_15448,N_14897,N_14591);
xor U15449 (N_15449,N_13865,N_13903);
xor U15450 (N_15450,N_14207,N_14647);
nor U15451 (N_15451,N_14545,N_14147);
or U15452 (N_15452,N_14093,N_14511);
nor U15453 (N_15453,N_14273,N_14711);
and U15454 (N_15454,N_13978,N_13782);
xnor U15455 (N_15455,N_14596,N_14103);
and U15456 (N_15456,N_14346,N_13994);
and U15457 (N_15457,N_14395,N_14736);
and U15458 (N_15458,N_14540,N_14562);
nand U15459 (N_15459,N_14559,N_14307);
and U15460 (N_15460,N_14312,N_14457);
and U15461 (N_15461,N_14240,N_14636);
nand U15462 (N_15462,N_14459,N_14521);
xor U15463 (N_15463,N_14025,N_14848);
or U15464 (N_15464,N_14095,N_14440);
and U15465 (N_15465,N_13983,N_14474);
xnor U15466 (N_15466,N_14251,N_14800);
nand U15467 (N_15467,N_13832,N_14682);
nor U15468 (N_15468,N_13947,N_14890);
or U15469 (N_15469,N_14784,N_14074);
nor U15470 (N_15470,N_14902,N_14969);
and U15471 (N_15471,N_13950,N_14515);
xnor U15472 (N_15472,N_14942,N_14332);
and U15473 (N_15473,N_14585,N_14501);
nor U15474 (N_15474,N_13974,N_14873);
or U15475 (N_15475,N_13855,N_14364);
nor U15476 (N_15476,N_14738,N_14323);
nand U15477 (N_15477,N_14309,N_14979);
nand U15478 (N_15478,N_14826,N_14024);
nor U15479 (N_15479,N_14624,N_14703);
or U15480 (N_15480,N_13795,N_14056);
nand U15481 (N_15481,N_14786,N_14290);
nand U15482 (N_15482,N_14047,N_13884);
nand U15483 (N_15483,N_14196,N_14246);
xnor U15484 (N_15484,N_14491,N_14679);
and U15485 (N_15485,N_14341,N_13754);
nand U15486 (N_15486,N_14198,N_14776);
xor U15487 (N_15487,N_14850,N_14480);
xor U15488 (N_15488,N_14222,N_14824);
xor U15489 (N_15489,N_14433,N_13765);
nand U15490 (N_15490,N_14917,N_14443);
nand U15491 (N_15491,N_14971,N_14008);
or U15492 (N_15492,N_14574,N_14015);
nor U15493 (N_15493,N_13990,N_14701);
xor U15494 (N_15494,N_14775,N_14720);
xnor U15495 (N_15495,N_14469,N_14138);
and U15496 (N_15496,N_14295,N_13949);
or U15497 (N_15497,N_14432,N_14050);
or U15498 (N_15498,N_14416,N_14949);
and U15499 (N_15499,N_14569,N_14339);
nor U15500 (N_15500,N_14975,N_14141);
nand U15501 (N_15501,N_14728,N_14546);
and U15502 (N_15502,N_14019,N_14066);
and U15503 (N_15503,N_14445,N_14194);
or U15504 (N_15504,N_14164,N_14098);
and U15505 (N_15505,N_14555,N_13956);
nor U15506 (N_15506,N_14034,N_14489);
nor U15507 (N_15507,N_13826,N_14167);
nor U15508 (N_15508,N_14614,N_14654);
nor U15509 (N_15509,N_14983,N_14564);
or U15510 (N_15510,N_14829,N_13825);
or U15511 (N_15511,N_14150,N_14551);
or U15512 (N_15512,N_14399,N_14345);
nand U15513 (N_15513,N_14919,N_14823);
or U15514 (N_15514,N_14219,N_14420);
xor U15515 (N_15515,N_14928,N_14838);
and U15516 (N_15516,N_14237,N_14581);
and U15517 (N_15517,N_13761,N_14472);
or U15518 (N_15518,N_14966,N_14543);
xor U15519 (N_15519,N_14582,N_14263);
and U15520 (N_15520,N_13989,N_14797);
or U15521 (N_15521,N_14683,N_13916);
nor U15522 (N_15522,N_13975,N_14030);
or U15523 (N_15523,N_13841,N_14606);
or U15524 (N_15524,N_14891,N_14320);
xor U15525 (N_15525,N_14118,N_14383);
or U15526 (N_15526,N_13952,N_14088);
or U15527 (N_15527,N_14206,N_13970);
and U15528 (N_15528,N_13767,N_14945);
nand U15529 (N_15529,N_14710,N_14695);
and U15530 (N_15530,N_14799,N_14017);
or U15531 (N_15531,N_14389,N_14199);
or U15532 (N_15532,N_14097,N_13771);
and U15533 (N_15533,N_13966,N_13786);
and U15534 (N_15534,N_14227,N_13751);
xnor U15535 (N_15535,N_14300,N_14916);
or U15536 (N_15536,N_14982,N_14592);
xnor U15537 (N_15537,N_14060,N_14718);
or U15538 (N_15538,N_14553,N_14541);
and U15539 (N_15539,N_14428,N_14170);
nand U15540 (N_15540,N_14305,N_14421);
nor U15541 (N_15541,N_14506,N_14691);
nor U15542 (N_15542,N_14304,N_14298);
xnor U15543 (N_15543,N_14901,N_14404);
and U15544 (N_15544,N_14505,N_14752);
xnor U15545 (N_15545,N_14513,N_14401);
and U15546 (N_15546,N_14610,N_14156);
nor U15547 (N_15547,N_14086,N_14924);
nand U15548 (N_15548,N_14573,N_14202);
xnor U15549 (N_15549,N_13836,N_14940);
nand U15550 (N_15550,N_14631,N_14934);
nand U15551 (N_15551,N_14159,N_14707);
or U15552 (N_15552,N_14380,N_14947);
xor U15553 (N_15553,N_14291,N_14912);
xnor U15554 (N_15554,N_13789,N_13904);
nor U15555 (N_15555,N_14804,N_14405);
nor U15556 (N_15556,N_13804,N_14229);
and U15557 (N_15557,N_14013,N_14058);
xnor U15558 (N_15558,N_14935,N_13891);
nand U15559 (N_15559,N_14528,N_13758);
nand U15560 (N_15560,N_14782,N_14397);
and U15561 (N_15561,N_14110,N_14465);
nor U15562 (N_15562,N_14915,N_13897);
and U15563 (N_15563,N_13753,N_14857);
nor U15564 (N_15564,N_13933,N_14642);
or U15565 (N_15565,N_14700,N_14879);
nand U15566 (N_15566,N_14798,N_13838);
and U15567 (N_15567,N_14035,N_14478);
and U15568 (N_15568,N_14508,N_14092);
xnor U15569 (N_15569,N_14238,N_14883);
nor U15570 (N_15570,N_14077,N_14666);
and U15571 (N_15571,N_14601,N_14071);
nor U15572 (N_15572,N_14939,N_14638);
or U15573 (N_15573,N_14620,N_14978);
and U15574 (N_15574,N_14333,N_14327);
nand U15575 (N_15575,N_14410,N_14242);
and U15576 (N_15576,N_13963,N_13931);
xor U15577 (N_15577,N_14811,N_14670);
nand U15578 (N_15578,N_14990,N_13853);
nand U15579 (N_15579,N_13858,N_14962);
nor U15580 (N_15580,N_13852,N_14774);
nor U15581 (N_15581,N_14347,N_14997);
xor U15582 (N_15582,N_14151,N_14036);
and U15583 (N_15583,N_14000,N_14936);
and U15584 (N_15584,N_14301,N_14643);
xnor U15585 (N_15585,N_14993,N_13890);
xor U15586 (N_15586,N_14124,N_14006);
xor U15587 (N_15587,N_14435,N_14223);
or U15588 (N_15588,N_14256,N_14961);
nand U15589 (N_15589,N_13918,N_14482);
nand U15590 (N_15590,N_14451,N_14450);
and U15591 (N_15591,N_14144,N_14067);
nor U15592 (N_15592,N_14926,N_14293);
xnor U15593 (N_15593,N_14751,N_14967);
xnor U15594 (N_15594,N_14068,N_14783);
nor U15595 (N_15595,N_14109,N_14386);
or U15596 (N_15596,N_14805,N_14889);
and U15597 (N_15597,N_14063,N_13851);
nand U15598 (N_15598,N_14542,N_14172);
xor U15599 (N_15599,N_14861,N_14051);
nor U15600 (N_15600,N_14716,N_14028);
nand U15601 (N_15601,N_13769,N_14269);
nand U15602 (N_15602,N_14174,N_14661);
nor U15603 (N_15603,N_14193,N_14054);
and U15604 (N_15604,N_14176,N_14987);
nand U15605 (N_15605,N_14107,N_14258);
xor U15606 (N_15606,N_14073,N_13915);
nand U15607 (N_15607,N_14042,N_14536);
and U15608 (N_15608,N_14580,N_13773);
or U15609 (N_15609,N_14225,N_14166);
nand U15610 (N_15610,N_14441,N_14084);
nand U15611 (N_15611,N_14184,N_14057);
nor U15612 (N_15612,N_14053,N_13848);
or U15613 (N_15613,N_14055,N_14040);
nand U15614 (N_15614,N_14660,N_13909);
nand U15615 (N_15615,N_14808,N_14538);
nor U15616 (N_15616,N_13922,N_14882);
xor U15617 (N_15617,N_14096,N_13805);
nor U15618 (N_15618,N_14286,N_14487);
xor U15619 (N_15619,N_14668,N_14593);
nand U15620 (N_15620,N_14091,N_14579);
nor U15621 (N_15621,N_14899,N_14045);
and U15622 (N_15622,N_14870,N_14479);
or U15623 (N_15623,N_13951,N_14365);
nor U15624 (N_15624,N_14009,N_13925);
xor U15625 (N_15625,N_14124,N_14400);
or U15626 (N_15626,N_14246,N_14635);
and U15627 (N_15627,N_13848,N_14529);
xor U15628 (N_15628,N_14608,N_14655);
or U15629 (N_15629,N_14423,N_14677);
nand U15630 (N_15630,N_13817,N_14968);
nor U15631 (N_15631,N_14531,N_13847);
or U15632 (N_15632,N_14252,N_13944);
xnor U15633 (N_15633,N_13857,N_14673);
nand U15634 (N_15634,N_14240,N_14553);
nand U15635 (N_15635,N_14055,N_14008);
or U15636 (N_15636,N_14364,N_14248);
xnor U15637 (N_15637,N_14284,N_14495);
and U15638 (N_15638,N_14242,N_14958);
xnor U15639 (N_15639,N_14111,N_14235);
nand U15640 (N_15640,N_14061,N_13927);
xnor U15641 (N_15641,N_14536,N_13864);
nand U15642 (N_15642,N_14133,N_14762);
and U15643 (N_15643,N_14607,N_14845);
or U15644 (N_15644,N_14384,N_14917);
xnor U15645 (N_15645,N_14524,N_14273);
xnor U15646 (N_15646,N_14626,N_14420);
or U15647 (N_15647,N_13948,N_14901);
nor U15648 (N_15648,N_14900,N_14640);
or U15649 (N_15649,N_14428,N_14331);
nor U15650 (N_15650,N_14488,N_14006);
xor U15651 (N_15651,N_14632,N_14371);
or U15652 (N_15652,N_14389,N_14686);
or U15653 (N_15653,N_14903,N_13770);
xor U15654 (N_15654,N_14629,N_14663);
xor U15655 (N_15655,N_14761,N_14658);
nand U15656 (N_15656,N_14523,N_14102);
nor U15657 (N_15657,N_14893,N_14000);
nor U15658 (N_15658,N_13888,N_13869);
xnor U15659 (N_15659,N_14057,N_14221);
and U15660 (N_15660,N_14347,N_14333);
or U15661 (N_15661,N_14841,N_14931);
or U15662 (N_15662,N_13756,N_14463);
or U15663 (N_15663,N_14951,N_14947);
or U15664 (N_15664,N_14727,N_14033);
nor U15665 (N_15665,N_14874,N_14855);
and U15666 (N_15666,N_14716,N_13977);
and U15667 (N_15667,N_13768,N_14750);
xnor U15668 (N_15668,N_14232,N_14205);
or U15669 (N_15669,N_14921,N_13762);
or U15670 (N_15670,N_14119,N_13823);
and U15671 (N_15671,N_13977,N_14894);
and U15672 (N_15672,N_14395,N_13898);
or U15673 (N_15673,N_14241,N_13829);
xnor U15674 (N_15674,N_14629,N_14497);
or U15675 (N_15675,N_14502,N_14005);
xor U15676 (N_15676,N_14052,N_14298);
nand U15677 (N_15677,N_13988,N_13884);
nor U15678 (N_15678,N_14840,N_13834);
and U15679 (N_15679,N_14728,N_14523);
xnor U15680 (N_15680,N_14489,N_14875);
and U15681 (N_15681,N_14095,N_14684);
nor U15682 (N_15682,N_14233,N_14029);
xnor U15683 (N_15683,N_14491,N_14357);
xnor U15684 (N_15684,N_14427,N_14043);
and U15685 (N_15685,N_14940,N_14658);
nor U15686 (N_15686,N_14499,N_14691);
nand U15687 (N_15687,N_14873,N_14158);
or U15688 (N_15688,N_14645,N_14993);
xnor U15689 (N_15689,N_13815,N_13918);
nand U15690 (N_15690,N_14749,N_14686);
and U15691 (N_15691,N_14320,N_14631);
nand U15692 (N_15692,N_13872,N_14808);
nor U15693 (N_15693,N_14535,N_13921);
or U15694 (N_15694,N_13812,N_13848);
or U15695 (N_15695,N_14395,N_14633);
or U15696 (N_15696,N_14436,N_14599);
or U15697 (N_15697,N_14375,N_14629);
and U15698 (N_15698,N_14407,N_13791);
or U15699 (N_15699,N_14789,N_14141);
xor U15700 (N_15700,N_14307,N_14478);
and U15701 (N_15701,N_14304,N_14631);
nor U15702 (N_15702,N_14595,N_14193);
or U15703 (N_15703,N_14671,N_13831);
nor U15704 (N_15704,N_13935,N_14513);
nor U15705 (N_15705,N_14116,N_14180);
or U15706 (N_15706,N_14281,N_14821);
nor U15707 (N_15707,N_14183,N_14638);
or U15708 (N_15708,N_14378,N_14736);
or U15709 (N_15709,N_14533,N_14702);
xor U15710 (N_15710,N_14647,N_14105);
and U15711 (N_15711,N_14015,N_14094);
and U15712 (N_15712,N_13869,N_14106);
nor U15713 (N_15713,N_14655,N_14018);
and U15714 (N_15714,N_14033,N_14155);
or U15715 (N_15715,N_14776,N_14240);
and U15716 (N_15716,N_14720,N_13932);
nor U15717 (N_15717,N_14169,N_14049);
and U15718 (N_15718,N_14895,N_14764);
and U15719 (N_15719,N_14050,N_13891);
nor U15720 (N_15720,N_13840,N_14766);
and U15721 (N_15721,N_14009,N_14036);
nand U15722 (N_15722,N_14478,N_14608);
and U15723 (N_15723,N_14888,N_13840);
xnor U15724 (N_15724,N_13949,N_13915);
and U15725 (N_15725,N_14278,N_14233);
nand U15726 (N_15726,N_14117,N_14022);
nand U15727 (N_15727,N_14521,N_14487);
nor U15728 (N_15728,N_14993,N_14558);
nand U15729 (N_15729,N_14824,N_13862);
nand U15730 (N_15730,N_14160,N_14272);
nor U15731 (N_15731,N_14874,N_14030);
or U15732 (N_15732,N_14316,N_14544);
nand U15733 (N_15733,N_13960,N_14335);
and U15734 (N_15734,N_13882,N_13831);
nor U15735 (N_15735,N_13920,N_14740);
or U15736 (N_15736,N_14459,N_14069);
or U15737 (N_15737,N_14680,N_14395);
nor U15738 (N_15738,N_13875,N_13963);
or U15739 (N_15739,N_13799,N_14801);
xnor U15740 (N_15740,N_14395,N_13969);
or U15741 (N_15741,N_14300,N_14389);
xnor U15742 (N_15742,N_14627,N_14664);
nor U15743 (N_15743,N_14807,N_14554);
or U15744 (N_15744,N_14365,N_13801);
xnor U15745 (N_15745,N_14445,N_14735);
and U15746 (N_15746,N_14825,N_14102);
nand U15747 (N_15747,N_14062,N_14540);
xnor U15748 (N_15748,N_14015,N_14197);
nand U15749 (N_15749,N_14671,N_13801);
nand U15750 (N_15750,N_14106,N_14918);
and U15751 (N_15751,N_14551,N_14599);
nor U15752 (N_15752,N_14556,N_14039);
xor U15753 (N_15753,N_14365,N_13919);
nor U15754 (N_15754,N_13963,N_14081);
nor U15755 (N_15755,N_14236,N_14780);
nand U15756 (N_15756,N_14405,N_14671);
nor U15757 (N_15757,N_14576,N_13925);
nor U15758 (N_15758,N_14529,N_14926);
or U15759 (N_15759,N_14559,N_14441);
nor U15760 (N_15760,N_14258,N_14538);
nand U15761 (N_15761,N_13924,N_14472);
nor U15762 (N_15762,N_14300,N_13839);
and U15763 (N_15763,N_13832,N_14918);
nor U15764 (N_15764,N_13809,N_14709);
or U15765 (N_15765,N_14434,N_13913);
nor U15766 (N_15766,N_14572,N_14933);
nor U15767 (N_15767,N_13874,N_14002);
xor U15768 (N_15768,N_13793,N_14599);
xor U15769 (N_15769,N_13948,N_14812);
nand U15770 (N_15770,N_14631,N_14957);
xor U15771 (N_15771,N_14938,N_14167);
xnor U15772 (N_15772,N_14678,N_14112);
nor U15773 (N_15773,N_14035,N_14340);
and U15774 (N_15774,N_14308,N_14295);
and U15775 (N_15775,N_13914,N_14125);
and U15776 (N_15776,N_14883,N_14653);
xnor U15777 (N_15777,N_14756,N_14906);
xnor U15778 (N_15778,N_14816,N_14659);
or U15779 (N_15779,N_14302,N_13816);
nor U15780 (N_15780,N_14847,N_14722);
and U15781 (N_15781,N_14256,N_14046);
nor U15782 (N_15782,N_13979,N_14464);
xor U15783 (N_15783,N_14992,N_14512);
xnor U15784 (N_15784,N_14371,N_14173);
xnor U15785 (N_15785,N_14875,N_13762);
nand U15786 (N_15786,N_14666,N_14641);
nor U15787 (N_15787,N_14321,N_14458);
nor U15788 (N_15788,N_14509,N_14823);
nor U15789 (N_15789,N_13883,N_13938);
or U15790 (N_15790,N_14316,N_14358);
or U15791 (N_15791,N_14778,N_14241);
nand U15792 (N_15792,N_14741,N_14323);
nand U15793 (N_15793,N_14955,N_14873);
nand U15794 (N_15794,N_14685,N_14158);
and U15795 (N_15795,N_14034,N_14438);
xnor U15796 (N_15796,N_13848,N_13916);
and U15797 (N_15797,N_14697,N_14842);
or U15798 (N_15798,N_13806,N_14253);
xnor U15799 (N_15799,N_14784,N_14545);
and U15800 (N_15800,N_14690,N_13907);
and U15801 (N_15801,N_13802,N_14472);
or U15802 (N_15802,N_14343,N_14183);
or U15803 (N_15803,N_14648,N_14106);
or U15804 (N_15804,N_14292,N_14328);
and U15805 (N_15805,N_14418,N_14893);
or U15806 (N_15806,N_14100,N_14579);
or U15807 (N_15807,N_14612,N_14829);
xor U15808 (N_15808,N_14723,N_14158);
xnor U15809 (N_15809,N_13841,N_14934);
nor U15810 (N_15810,N_14789,N_13947);
and U15811 (N_15811,N_14977,N_13940);
nand U15812 (N_15812,N_14495,N_14903);
xnor U15813 (N_15813,N_14841,N_13817);
nor U15814 (N_15814,N_14426,N_14543);
and U15815 (N_15815,N_13899,N_14412);
nand U15816 (N_15816,N_14889,N_14559);
xnor U15817 (N_15817,N_14779,N_14976);
nor U15818 (N_15818,N_14951,N_14549);
nor U15819 (N_15819,N_13834,N_14158);
nor U15820 (N_15820,N_14980,N_14511);
nand U15821 (N_15821,N_14869,N_14468);
xnor U15822 (N_15822,N_14248,N_14635);
nor U15823 (N_15823,N_14688,N_14487);
nor U15824 (N_15824,N_14553,N_14238);
nand U15825 (N_15825,N_13865,N_13771);
xor U15826 (N_15826,N_13825,N_13998);
nor U15827 (N_15827,N_14403,N_14726);
nand U15828 (N_15828,N_14941,N_14164);
nor U15829 (N_15829,N_14505,N_14376);
nand U15830 (N_15830,N_14400,N_14815);
nand U15831 (N_15831,N_13959,N_14932);
and U15832 (N_15832,N_14347,N_14111);
or U15833 (N_15833,N_14474,N_14228);
nor U15834 (N_15834,N_13825,N_14055);
and U15835 (N_15835,N_14843,N_14826);
and U15836 (N_15836,N_14487,N_14348);
nand U15837 (N_15837,N_14501,N_14846);
nor U15838 (N_15838,N_14119,N_14430);
and U15839 (N_15839,N_13975,N_14413);
or U15840 (N_15840,N_14562,N_13858);
and U15841 (N_15841,N_14906,N_14894);
xor U15842 (N_15842,N_14772,N_14317);
nor U15843 (N_15843,N_14090,N_14207);
or U15844 (N_15844,N_14840,N_13880);
nor U15845 (N_15845,N_13938,N_14560);
nor U15846 (N_15846,N_14243,N_14974);
nand U15847 (N_15847,N_14724,N_13858);
xor U15848 (N_15848,N_14835,N_14351);
nor U15849 (N_15849,N_13991,N_14027);
xor U15850 (N_15850,N_14615,N_13812);
nand U15851 (N_15851,N_14840,N_14002);
xor U15852 (N_15852,N_14384,N_14063);
nand U15853 (N_15853,N_14947,N_14979);
and U15854 (N_15854,N_14421,N_14993);
nor U15855 (N_15855,N_14756,N_13767);
nor U15856 (N_15856,N_14835,N_14000);
or U15857 (N_15857,N_14136,N_14636);
and U15858 (N_15858,N_14383,N_14652);
xor U15859 (N_15859,N_14355,N_14992);
or U15860 (N_15860,N_14476,N_14488);
nand U15861 (N_15861,N_14298,N_14487);
nor U15862 (N_15862,N_14683,N_14694);
or U15863 (N_15863,N_14504,N_14984);
or U15864 (N_15864,N_14936,N_14991);
and U15865 (N_15865,N_14760,N_14703);
nand U15866 (N_15866,N_13756,N_14516);
and U15867 (N_15867,N_14141,N_13883);
and U15868 (N_15868,N_13937,N_14411);
or U15869 (N_15869,N_14717,N_14939);
xnor U15870 (N_15870,N_14999,N_13847);
nand U15871 (N_15871,N_14634,N_14259);
or U15872 (N_15872,N_14967,N_14581);
nor U15873 (N_15873,N_14313,N_13773);
and U15874 (N_15874,N_14295,N_13918);
nor U15875 (N_15875,N_13996,N_14819);
nor U15876 (N_15876,N_14090,N_14557);
nand U15877 (N_15877,N_14529,N_14960);
nor U15878 (N_15878,N_13825,N_14956);
and U15879 (N_15879,N_14120,N_14485);
nor U15880 (N_15880,N_14450,N_14124);
xor U15881 (N_15881,N_14537,N_13812);
xor U15882 (N_15882,N_14011,N_13965);
nor U15883 (N_15883,N_14484,N_14815);
xnor U15884 (N_15884,N_14392,N_14299);
nand U15885 (N_15885,N_14099,N_14594);
xnor U15886 (N_15886,N_14163,N_14627);
nand U15887 (N_15887,N_14619,N_14850);
or U15888 (N_15888,N_14491,N_14836);
nor U15889 (N_15889,N_14442,N_14159);
and U15890 (N_15890,N_14009,N_14506);
or U15891 (N_15891,N_13804,N_13899);
nand U15892 (N_15892,N_14282,N_13979);
nor U15893 (N_15893,N_13793,N_14539);
nand U15894 (N_15894,N_14409,N_14531);
or U15895 (N_15895,N_14125,N_14988);
nand U15896 (N_15896,N_14277,N_14743);
and U15897 (N_15897,N_14421,N_14507);
xnor U15898 (N_15898,N_14172,N_14055);
xor U15899 (N_15899,N_14730,N_13949);
xor U15900 (N_15900,N_14455,N_14118);
or U15901 (N_15901,N_14937,N_14053);
and U15902 (N_15902,N_13868,N_13934);
or U15903 (N_15903,N_14118,N_14426);
or U15904 (N_15904,N_14661,N_14812);
and U15905 (N_15905,N_14887,N_14452);
nor U15906 (N_15906,N_13761,N_13954);
and U15907 (N_15907,N_14629,N_14634);
and U15908 (N_15908,N_14002,N_14671);
xor U15909 (N_15909,N_13812,N_14377);
nand U15910 (N_15910,N_14439,N_14765);
nor U15911 (N_15911,N_14334,N_14917);
or U15912 (N_15912,N_13854,N_13822);
or U15913 (N_15913,N_13892,N_14141);
xor U15914 (N_15914,N_14815,N_14273);
xnor U15915 (N_15915,N_13910,N_13895);
nand U15916 (N_15916,N_14728,N_14958);
nor U15917 (N_15917,N_14308,N_13783);
nand U15918 (N_15918,N_14032,N_14756);
and U15919 (N_15919,N_14351,N_14342);
xnor U15920 (N_15920,N_14265,N_14748);
nor U15921 (N_15921,N_14866,N_14043);
xor U15922 (N_15922,N_14099,N_13838);
nor U15923 (N_15923,N_14686,N_14625);
nand U15924 (N_15924,N_14050,N_14615);
or U15925 (N_15925,N_14932,N_13921);
and U15926 (N_15926,N_13930,N_13861);
and U15927 (N_15927,N_14566,N_14026);
or U15928 (N_15928,N_14971,N_13949);
nor U15929 (N_15929,N_14105,N_14161);
nand U15930 (N_15930,N_13764,N_14965);
xor U15931 (N_15931,N_14869,N_14685);
and U15932 (N_15932,N_14834,N_14536);
nor U15933 (N_15933,N_13849,N_14680);
or U15934 (N_15934,N_14202,N_14744);
and U15935 (N_15935,N_14254,N_14597);
xor U15936 (N_15936,N_14107,N_14483);
or U15937 (N_15937,N_13754,N_14372);
and U15938 (N_15938,N_14505,N_14165);
nand U15939 (N_15939,N_14045,N_14427);
or U15940 (N_15940,N_14979,N_14769);
nor U15941 (N_15941,N_14288,N_14727);
or U15942 (N_15942,N_13813,N_14146);
nor U15943 (N_15943,N_14506,N_14030);
nor U15944 (N_15944,N_14433,N_14183);
nor U15945 (N_15945,N_14612,N_14823);
or U15946 (N_15946,N_14743,N_14438);
and U15947 (N_15947,N_14204,N_14947);
or U15948 (N_15948,N_14872,N_14990);
and U15949 (N_15949,N_14944,N_14020);
and U15950 (N_15950,N_14858,N_14607);
nand U15951 (N_15951,N_14326,N_14084);
or U15952 (N_15952,N_14165,N_14802);
xnor U15953 (N_15953,N_13993,N_14419);
and U15954 (N_15954,N_14447,N_14834);
nand U15955 (N_15955,N_14907,N_13750);
nand U15956 (N_15956,N_14732,N_13802);
nand U15957 (N_15957,N_14919,N_14287);
nor U15958 (N_15958,N_14293,N_13870);
nor U15959 (N_15959,N_14357,N_14891);
and U15960 (N_15960,N_14438,N_14085);
nand U15961 (N_15961,N_14503,N_14780);
nor U15962 (N_15962,N_14577,N_14349);
nor U15963 (N_15963,N_14372,N_13837);
and U15964 (N_15964,N_13960,N_14429);
or U15965 (N_15965,N_14272,N_14099);
nand U15966 (N_15966,N_14037,N_13918);
and U15967 (N_15967,N_14470,N_14300);
nand U15968 (N_15968,N_14887,N_14630);
or U15969 (N_15969,N_14157,N_14133);
and U15970 (N_15970,N_14567,N_14594);
nand U15971 (N_15971,N_14210,N_14402);
nor U15972 (N_15972,N_14313,N_14611);
xor U15973 (N_15973,N_14313,N_13802);
or U15974 (N_15974,N_14712,N_14360);
or U15975 (N_15975,N_14141,N_14901);
and U15976 (N_15976,N_14039,N_14634);
and U15977 (N_15977,N_14773,N_14249);
or U15978 (N_15978,N_14742,N_14745);
and U15979 (N_15979,N_14927,N_14635);
or U15980 (N_15980,N_13775,N_14374);
xnor U15981 (N_15981,N_14776,N_14876);
or U15982 (N_15982,N_14609,N_14043);
xor U15983 (N_15983,N_13967,N_14920);
xnor U15984 (N_15984,N_14026,N_13830);
or U15985 (N_15985,N_14957,N_14918);
nor U15986 (N_15986,N_14816,N_14211);
xnor U15987 (N_15987,N_14678,N_13754);
nand U15988 (N_15988,N_14424,N_14011);
and U15989 (N_15989,N_14448,N_14338);
or U15990 (N_15990,N_14966,N_14564);
xor U15991 (N_15991,N_14843,N_14604);
or U15992 (N_15992,N_14803,N_14334);
xnor U15993 (N_15993,N_14307,N_13989);
nand U15994 (N_15994,N_14278,N_14246);
nand U15995 (N_15995,N_13799,N_14541);
or U15996 (N_15996,N_14092,N_14995);
nor U15997 (N_15997,N_14409,N_14188);
or U15998 (N_15998,N_14684,N_14948);
and U15999 (N_15999,N_14116,N_14345);
or U16000 (N_16000,N_13923,N_14861);
and U16001 (N_16001,N_14653,N_14249);
or U16002 (N_16002,N_13845,N_14230);
and U16003 (N_16003,N_13766,N_14909);
or U16004 (N_16004,N_14820,N_14840);
and U16005 (N_16005,N_14893,N_13751);
nor U16006 (N_16006,N_13839,N_14563);
nor U16007 (N_16007,N_13882,N_13999);
nand U16008 (N_16008,N_13794,N_14459);
and U16009 (N_16009,N_14341,N_13864);
xnor U16010 (N_16010,N_14691,N_14576);
nor U16011 (N_16011,N_14622,N_14182);
nand U16012 (N_16012,N_14508,N_14212);
xnor U16013 (N_16013,N_13999,N_14685);
nand U16014 (N_16014,N_13869,N_14952);
or U16015 (N_16015,N_13877,N_14103);
nand U16016 (N_16016,N_14643,N_14973);
nor U16017 (N_16017,N_14613,N_13770);
and U16018 (N_16018,N_14146,N_14740);
xnor U16019 (N_16019,N_14399,N_13899);
and U16020 (N_16020,N_13871,N_14936);
xor U16021 (N_16021,N_14305,N_13767);
and U16022 (N_16022,N_13941,N_14117);
or U16023 (N_16023,N_14245,N_13785);
nand U16024 (N_16024,N_13773,N_14161);
and U16025 (N_16025,N_14410,N_13760);
nor U16026 (N_16026,N_14846,N_14229);
xnor U16027 (N_16027,N_14167,N_14087);
nand U16028 (N_16028,N_14434,N_14558);
nand U16029 (N_16029,N_14459,N_14871);
xnor U16030 (N_16030,N_14265,N_14217);
and U16031 (N_16031,N_14897,N_14141);
xnor U16032 (N_16032,N_13863,N_14450);
or U16033 (N_16033,N_14303,N_14513);
nor U16034 (N_16034,N_14412,N_14633);
nand U16035 (N_16035,N_14358,N_14659);
nor U16036 (N_16036,N_14801,N_14408);
or U16037 (N_16037,N_14930,N_14861);
and U16038 (N_16038,N_13960,N_14950);
nand U16039 (N_16039,N_14227,N_14813);
xnor U16040 (N_16040,N_14169,N_14138);
and U16041 (N_16041,N_14956,N_14271);
nand U16042 (N_16042,N_14098,N_14249);
or U16043 (N_16043,N_14154,N_14726);
and U16044 (N_16044,N_14423,N_14866);
nor U16045 (N_16045,N_13830,N_14668);
nor U16046 (N_16046,N_14670,N_14116);
and U16047 (N_16047,N_14509,N_13778);
nand U16048 (N_16048,N_14862,N_14904);
xnor U16049 (N_16049,N_13787,N_14347);
nand U16050 (N_16050,N_14982,N_14762);
nand U16051 (N_16051,N_14443,N_14392);
nor U16052 (N_16052,N_13921,N_14236);
or U16053 (N_16053,N_14455,N_14277);
nor U16054 (N_16054,N_14102,N_14977);
nand U16055 (N_16055,N_14872,N_14831);
xnor U16056 (N_16056,N_14451,N_14239);
nor U16057 (N_16057,N_14496,N_14823);
or U16058 (N_16058,N_13977,N_14615);
and U16059 (N_16059,N_14267,N_14884);
nor U16060 (N_16060,N_14668,N_14718);
nor U16061 (N_16061,N_14038,N_13935);
xnor U16062 (N_16062,N_13949,N_14477);
nand U16063 (N_16063,N_14546,N_14131);
xnor U16064 (N_16064,N_14121,N_14725);
nand U16065 (N_16065,N_14333,N_14615);
nor U16066 (N_16066,N_13884,N_14035);
xor U16067 (N_16067,N_14239,N_13804);
nor U16068 (N_16068,N_14997,N_14413);
or U16069 (N_16069,N_14365,N_14064);
nand U16070 (N_16070,N_13775,N_14152);
nand U16071 (N_16071,N_14283,N_14341);
or U16072 (N_16072,N_14781,N_14018);
nor U16073 (N_16073,N_14400,N_14696);
or U16074 (N_16074,N_14533,N_13758);
xnor U16075 (N_16075,N_14562,N_13794);
nor U16076 (N_16076,N_13992,N_14355);
xnor U16077 (N_16077,N_14043,N_14972);
nand U16078 (N_16078,N_14995,N_13859);
nand U16079 (N_16079,N_14946,N_14503);
or U16080 (N_16080,N_14772,N_13984);
nand U16081 (N_16081,N_14088,N_14347);
nand U16082 (N_16082,N_14613,N_14257);
xnor U16083 (N_16083,N_14750,N_14897);
or U16084 (N_16084,N_14614,N_14148);
and U16085 (N_16085,N_14171,N_14919);
and U16086 (N_16086,N_14414,N_13874);
or U16087 (N_16087,N_14952,N_14694);
or U16088 (N_16088,N_14492,N_14686);
and U16089 (N_16089,N_14064,N_14485);
nor U16090 (N_16090,N_14434,N_14034);
nand U16091 (N_16091,N_14516,N_14460);
and U16092 (N_16092,N_14447,N_14558);
or U16093 (N_16093,N_14862,N_14429);
nor U16094 (N_16094,N_14608,N_14115);
or U16095 (N_16095,N_13989,N_14713);
nand U16096 (N_16096,N_14168,N_14303);
and U16097 (N_16097,N_13998,N_14127);
or U16098 (N_16098,N_13881,N_14649);
xnor U16099 (N_16099,N_14166,N_14354);
xor U16100 (N_16100,N_14942,N_14430);
or U16101 (N_16101,N_14440,N_14254);
xnor U16102 (N_16102,N_14896,N_13845);
xnor U16103 (N_16103,N_14256,N_14920);
nor U16104 (N_16104,N_14896,N_14937);
nor U16105 (N_16105,N_14674,N_14546);
nand U16106 (N_16106,N_13775,N_14961);
nor U16107 (N_16107,N_14570,N_14896);
xor U16108 (N_16108,N_14677,N_14097);
or U16109 (N_16109,N_14937,N_14242);
xor U16110 (N_16110,N_14437,N_14074);
and U16111 (N_16111,N_14117,N_14264);
xor U16112 (N_16112,N_14133,N_14255);
nor U16113 (N_16113,N_14353,N_14829);
nor U16114 (N_16114,N_14013,N_14738);
nor U16115 (N_16115,N_14379,N_14895);
or U16116 (N_16116,N_14205,N_14918);
nand U16117 (N_16117,N_14261,N_14319);
nand U16118 (N_16118,N_14735,N_13811);
xor U16119 (N_16119,N_14965,N_13992);
xor U16120 (N_16120,N_14757,N_13983);
and U16121 (N_16121,N_13886,N_14150);
nand U16122 (N_16122,N_14021,N_14358);
nor U16123 (N_16123,N_14428,N_14380);
or U16124 (N_16124,N_14466,N_13816);
nor U16125 (N_16125,N_14968,N_14052);
nor U16126 (N_16126,N_14153,N_14472);
xnor U16127 (N_16127,N_14484,N_14564);
nor U16128 (N_16128,N_14956,N_13995);
nand U16129 (N_16129,N_14708,N_14614);
nand U16130 (N_16130,N_14778,N_14173);
or U16131 (N_16131,N_14943,N_14193);
or U16132 (N_16132,N_14355,N_14677);
nand U16133 (N_16133,N_14491,N_13998);
xor U16134 (N_16134,N_13837,N_14067);
nor U16135 (N_16135,N_13941,N_14827);
or U16136 (N_16136,N_13824,N_14394);
nand U16137 (N_16137,N_13830,N_14382);
and U16138 (N_16138,N_14304,N_14166);
and U16139 (N_16139,N_14640,N_14444);
nor U16140 (N_16140,N_14220,N_14765);
xnor U16141 (N_16141,N_13903,N_14627);
nor U16142 (N_16142,N_14612,N_14142);
nor U16143 (N_16143,N_13776,N_14565);
and U16144 (N_16144,N_14226,N_13969);
or U16145 (N_16145,N_13999,N_14198);
or U16146 (N_16146,N_14195,N_14159);
xor U16147 (N_16147,N_14964,N_14856);
nor U16148 (N_16148,N_14067,N_14534);
xor U16149 (N_16149,N_14326,N_13760);
or U16150 (N_16150,N_14008,N_13759);
and U16151 (N_16151,N_14165,N_14162);
or U16152 (N_16152,N_13810,N_14972);
or U16153 (N_16153,N_14771,N_14625);
or U16154 (N_16154,N_14149,N_14019);
or U16155 (N_16155,N_14654,N_13966);
and U16156 (N_16156,N_14024,N_14861);
nand U16157 (N_16157,N_14104,N_14618);
xor U16158 (N_16158,N_14335,N_14919);
nor U16159 (N_16159,N_14160,N_14825);
and U16160 (N_16160,N_14550,N_14285);
or U16161 (N_16161,N_14178,N_14271);
nor U16162 (N_16162,N_14286,N_13867);
and U16163 (N_16163,N_14963,N_14125);
xnor U16164 (N_16164,N_14227,N_14305);
xnor U16165 (N_16165,N_14333,N_13919);
xnor U16166 (N_16166,N_14033,N_14792);
or U16167 (N_16167,N_14307,N_14368);
nand U16168 (N_16168,N_14831,N_14184);
and U16169 (N_16169,N_14389,N_14007);
or U16170 (N_16170,N_14797,N_14488);
nand U16171 (N_16171,N_13796,N_14367);
and U16172 (N_16172,N_14850,N_14987);
and U16173 (N_16173,N_14266,N_14963);
or U16174 (N_16174,N_14885,N_14556);
and U16175 (N_16175,N_14468,N_14812);
nand U16176 (N_16176,N_14435,N_14643);
and U16177 (N_16177,N_14718,N_14323);
or U16178 (N_16178,N_14414,N_14696);
xor U16179 (N_16179,N_14095,N_14242);
nand U16180 (N_16180,N_14619,N_14492);
nand U16181 (N_16181,N_14113,N_14017);
nand U16182 (N_16182,N_14339,N_14207);
nor U16183 (N_16183,N_14409,N_14171);
nand U16184 (N_16184,N_14732,N_14255);
and U16185 (N_16185,N_13915,N_13885);
and U16186 (N_16186,N_14399,N_13924);
xnor U16187 (N_16187,N_14739,N_14316);
or U16188 (N_16188,N_13799,N_13753);
and U16189 (N_16189,N_14700,N_14306);
and U16190 (N_16190,N_14174,N_14553);
and U16191 (N_16191,N_14409,N_14186);
or U16192 (N_16192,N_14833,N_14534);
nand U16193 (N_16193,N_14248,N_13979);
and U16194 (N_16194,N_14119,N_14441);
and U16195 (N_16195,N_13922,N_14697);
or U16196 (N_16196,N_14460,N_14275);
and U16197 (N_16197,N_14193,N_14023);
nand U16198 (N_16198,N_14869,N_14323);
and U16199 (N_16199,N_14103,N_14083);
xnor U16200 (N_16200,N_13908,N_14729);
xor U16201 (N_16201,N_14856,N_14259);
nor U16202 (N_16202,N_14421,N_14861);
nand U16203 (N_16203,N_14366,N_14362);
and U16204 (N_16204,N_13796,N_14520);
or U16205 (N_16205,N_14982,N_14097);
nor U16206 (N_16206,N_14883,N_14554);
and U16207 (N_16207,N_14778,N_14955);
nand U16208 (N_16208,N_13774,N_14256);
and U16209 (N_16209,N_14220,N_13839);
and U16210 (N_16210,N_14969,N_14976);
or U16211 (N_16211,N_14669,N_13919);
or U16212 (N_16212,N_13893,N_14398);
nor U16213 (N_16213,N_14376,N_14115);
nand U16214 (N_16214,N_14804,N_14337);
or U16215 (N_16215,N_14476,N_13882);
xor U16216 (N_16216,N_14458,N_14092);
nor U16217 (N_16217,N_14073,N_14076);
nand U16218 (N_16218,N_14694,N_14630);
and U16219 (N_16219,N_14276,N_14671);
nand U16220 (N_16220,N_14503,N_14433);
nor U16221 (N_16221,N_14143,N_13981);
or U16222 (N_16222,N_14198,N_14331);
nand U16223 (N_16223,N_14861,N_14067);
nor U16224 (N_16224,N_14766,N_14329);
and U16225 (N_16225,N_13923,N_14289);
nand U16226 (N_16226,N_13755,N_13871);
and U16227 (N_16227,N_14111,N_13936);
nor U16228 (N_16228,N_14940,N_14862);
and U16229 (N_16229,N_14647,N_14394);
nor U16230 (N_16230,N_14409,N_13896);
nor U16231 (N_16231,N_14463,N_14078);
or U16232 (N_16232,N_14465,N_14989);
nand U16233 (N_16233,N_14339,N_14262);
and U16234 (N_16234,N_13962,N_14938);
or U16235 (N_16235,N_14778,N_14593);
xor U16236 (N_16236,N_13975,N_14784);
nor U16237 (N_16237,N_14722,N_14003);
nand U16238 (N_16238,N_13986,N_13899);
or U16239 (N_16239,N_14995,N_14544);
or U16240 (N_16240,N_13892,N_13816);
xor U16241 (N_16241,N_14081,N_13849);
or U16242 (N_16242,N_13987,N_14142);
xor U16243 (N_16243,N_14510,N_14553);
nand U16244 (N_16244,N_14881,N_14787);
and U16245 (N_16245,N_14346,N_14035);
and U16246 (N_16246,N_14016,N_14884);
nand U16247 (N_16247,N_14731,N_14663);
and U16248 (N_16248,N_14715,N_14919);
xnor U16249 (N_16249,N_14633,N_14480);
nand U16250 (N_16250,N_15265,N_16241);
nand U16251 (N_16251,N_15252,N_15411);
nor U16252 (N_16252,N_15450,N_15728);
xor U16253 (N_16253,N_16131,N_15864);
nand U16254 (N_16254,N_15848,N_15125);
nand U16255 (N_16255,N_15374,N_16142);
or U16256 (N_16256,N_15830,N_15973);
and U16257 (N_16257,N_15998,N_15457);
and U16258 (N_16258,N_16206,N_15665);
nand U16259 (N_16259,N_15048,N_15302);
or U16260 (N_16260,N_15805,N_15977);
xnor U16261 (N_16261,N_16176,N_15334);
nor U16262 (N_16262,N_16012,N_15957);
nand U16263 (N_16263,N_16139,N_15837);
or U16264 (N_16264,N_15697,N_15887);
xnor U16265 (N_16265,N_15078,N_16192);
and U16266 (N_16266,N_15505,N_15352);
nor U16267 (N_16267,N_15012,N_15908);
nor U16268 (N_16268,N_15165,N_16108);
nand U16269 (N_16269,N_15490,N_15640);
or U16270 (N_16270,N_15590,N_15239);
xnor U16271 (N_16271,N_15933,N_16039);
nor U16272 (N_16272,N_16185,N_15901);
or U16273 (N_16273,N_15024,N_15788);
and U16274 (N_16274,N_15713,N_15006);
nand U16275 (N_16275,N_15531,N_16095);
nand U16276 (N_16276,N_16088,N_15794);
or U16277 (N_16277,N_15433,N_16002);
nor U16278 (N_16278,N_15199,N_15202);
nor U16279 (N_16279,N_15310,N_16136);
nor U16280 (N_16280,N_15475,N_15154);
and U16281 (N_16281,N_15379,N_15612);
or U16282 (N_16282,N_16147,N_16244);
xnor U16283 (N_16283,N_15312,N_15341);
nor U16284 (N_16284,N_15067,N_15878);
xor U16285 (N_16285,N_15580,N_15288);
or U16286 (N_16286,N_16169,N_15567);
xor U16287 (N_16287,N_15123,N_15255);
nor U16288 (N_16288,N_15421,N_16084);
nand U16289 (N_16289,N_15886,N_15696);
or U16290 (N_16290,N_15645,N_15537);
and U16291 (N_16291,N_15970,N_15711);
or U16292 (N_16292,N_16228,N_15327);
nand U16293 (N_16293,N_15925,N_15553);
or U16294 (N_16294,N_15268,N_15126);
nor U16295 (N_16295,N_15671,N_16209);
nand U16296 (N_16296,N_15384,N_15776);
or U16297 (N_16297,N_15180,N_15008);
and U16298 (N_16298,N_15717,N_16130);
nand U16299 (N_16299,N_15597,N_16051);
and U16300 (N_16300,N_16219,N_15897);
nor U16301 (N_16301,N_15244,N_15927);
nor U16302 (N_16302,N_15122,N_15369);
nor U16303 (N_16303,N_15330,N_15217);
nand U16304 (N_16304,N_16011,N_15349);
or U16305 (N_16305,N_15955,N_15996);
or U16306 (N_16306,N_16031,N_15539);
and U16307 (N_16307,N_15514,N_15907);
xnor U16308 (N_16308,N_15481,N_15285);
or U16309 (N_16309,N_15915,N_15495);
or U16310 (N_16310,N_16210,N_15720);
or U16311 (N_16311,N_15592,N_15113);
nand U16312 (N_16312,N_15695,N_16124);
and U16313 (N_16313,N_15380,N_15183);
or U16314 (N_16314,N_16072,N_16163);
nor U16315 (N_16315,N_15178,N_16216);
or U16316 (N_16316,N_15423,N_16240);
xnor U16317 (N_16317,N_16211,N_15773);
xor U16318 (N_16318,N_15872,N_15503);
nand U16319 (N_16319,N_15545,N_15052);
nor U16320 (N_16320,N_15777,N_16246);
nand U16321 (N_16321,N_15694,N_15354);
and U16322 (N_16322,N_15011,N_15945);
or U16323 (N_16323,N_16069,N_16123);
xnor U16324 (N_16324,N_15118,N_15710);
xnor U16325 (N_16325,N_15809,N_15129);
nand U16326 (N_16326,N_15902,N_15296);
xnor U16327 (N_16327,N_15947,N_15820);
nor U16328 (N_16328,N_15112,N_16135);
nand U16329 (N_16329,N_15443,N_15241);
nand U16330 (N_16330,N_15905,N_15976);
nand U16331 (N_16331,N_15515,N_16125);
nand U16332 (N_16332,N_15845,N_15096);
and U16333 (N_16333,N_15068,N_15863);
xor U16334 (N_16334,N_15922,N_15752);
or U16335 (N_16335,N_15587,N_15541);
nand U16336 (N_16336,N_16243,N_15815);
nor U16337 (N_16337,N_15543,N_15336);
nor U16338 (N_16338,N_15572,N_16188);
xnor U16339 (N_16339,N_15552,N_15859);
xnor U16340 (N_16340,N_15502,N_16153);
nor U16341 (N_16341,N_15045,N_15226);
xor U16342 (N_16342,N_15975,N_16107);
and U16343 (N_16343,N_15677,N_16170);
or U16344 (N_16344,N_15950,N_15037);
nor U16345 (N_16345,N_15600,N_16134);
nor U16346 (N_16346,N_15446,N_15166);
nand U16347 (N_16347,N_15262,N_15232);
xor U16348 (N_16348,N_15281,N_15599);
or U16349 (N_16349,N_15185,N_16221);
nand U16350 (N_16350,N_15127,N_15714);
and U16351 (N_16351,N_16180,N_15066);
nand U16352 (N_16352,N_15023,N_15817);
and U16353 (N_16353,N_15079,N_15134);
or U16354 (N_16354,N_15662,N_16249);
nand U16355 (N_16355,N_15501,N_15753);
xnor U16356 (N_16356,N_16076,N_15210);
and U16357 (N_16357,N_15801,N_15842);
nor U16358 (N_16358,N_15931,N_15570);
nand U16359 (N_16359,N_16214,N_15381);
and U16360 (N_16360,N_16085,N_15478);
and U16361 (N_16361,N_16101,N_15732);
nand U16362 (N_16362,N_16191,N_15028);
or U16363 (N_16363,N_15688,N_15877);
nand U16364 (N_16364,N_16024,N_15781);
xnor U16365 (N_16365,N_16053,N_16202);
xor U16366 (N_16366,N_15988,N_16200);
and U16367 (N_16367,N_15519,N_15004);
and U16368 (N_16368,N_15442,N_16042);
and U16369 (N_16369,N_15147,N_15946);
nand U16370 (N_16370,N_15253,N_15756);
or U16371 (N_16371,N_16046,N_15783);
xor U16372 (N_16372,N_15343,N_15057);
or U16373 (N_16373,N_15787,N_15486);
xor U16374 (N_16374,N_16132,N_15739);
nor U16375 (N_16375,N_15091,N_15974);
and U16376 (N_16376,N_15243,N_15201);
or U16377 (N_16377,N_16043,N_16203);
xor U16378 (N_16378,N_15483,N_16225);
nand U16379 (N_16379,N_16087,N_15420);
nor U16380 (N_16380,N_15063,N_16057);
or U16381 (N_16381,N_15138,N_15642);
nor U16382 (N_16382,N_15621,N_15247);
xor U16383 (N_16383,N_15060,N_15375);
nand U16384 (N_16384,N_15521,N_15811);
xor U16385 (N_16385,N_15992,N_15928);
nand U16386 (N_16386,N_16067,N_16226);
and U16387 (N_16387,N_15387,N_15406);
or U16388 (N_16388,N_15022,N_15629);
xnor U16389 (N_16389,N_15190,N_15814);
and U16390 (N_16390,N_15979,N_16149);
nor U16391 (N_16391,N_15738,N_15342);
or U16392 (N_16392,N_15624,N_16006);
and U16393 (N_16393,N_15293,N_15823);
nand U16394 (N_16394,N_15089,N_16173);
xnor U16395 (N_16395,N_15080,N_15876);
or U16396 (N_16396,N_15598,N_15280);
nand U16397 (N_16397,N_16205,N_15286);
or U16398 (N_16398,N_15359,N_15355);
nand U16399 (N_16399,N_15687,N_15013);
xor U16400 (N_16400,N_15463,N_16034);
nor U16401 (N_16401,N_15526,N_15875);
nor U16402 (N_16402,N_15378,N_15634);
or U16403 (N_16403,N_15167,N_16010);
and U16404 (N_16404,N_15764,N_15750);
nor U16405 (N_16405,N_15292,N_15712);
and U16406 (N_16406,N_16179,N_15661);
or U16407 (N_16407,N_15106,N_15909);
nor U16408 (N_16408,N_15536,N_16190);
and U16409 (N_16409,N_15464,N_15431);
or U16410 (N_16410,N_15276,N_16174);
xnor U16411 (N_16411,N_15718,N_16074);
or U16412 (N_16412,N_15699,N_15520);
nand U16413 (N_16413,N_15110,N_16245);
and U16414 (N_16414,N_15549,N_15758);
and U16415 (N_16415,N_15020,N_16129);
xnor U16416 (N_16416,N_15430,N_16102);
nand U16417 (N_16417,N_15499,N_16030);
nor U16418 (N_16418,N_15492,N_15469);
nand U16419 (N_16419,N_15275,N_15365);
and U16420 (N_16420,N_15193,N_16143);
nor U16421 (N_16421,N_15414,N_16151);
and U16422 (N_16422,N_15324,N_15647);
or U16423 (N_16423,N_15954,N_15216);
or U16424 (N_16424,N_15207,N_15576);
or U16425 (N_16425,N_16196,N_15325);
nand U16426 (N_16426,N_15559,N_16040);
and U16427 (N_16427,N_15831,N_15943);
and U16428 (N_16428,N_15072,N_15615);
or U16429 (N_16429,N_15044,N_15504);
nor U16430 (N_16430,N_15054,N_16213);
and U16431 (N_16431,N_15095,N_15796);
and U16432 (N_16432,N_16155,N_16016);
nand U16433 (N_16433,N_15500,N_16075);
and U16434 (N_16434,N_15938,N_16023);
and U16435 (N_16435,N_15852,N_15754);
xor U16436 (N_16436,N_15186,N_15546);
xor U16437 (N_16437,N_15363,N_15156);
or U16438 (N_16438,N_15610,N_15466);
or U16439 (N_16439,N_16201,N_15672);
xnor U16440 (N_16440,N_15828,N_15120);
nor U16441 (N_16441,N_15358,N_15473);
nor U16442 (N_16442,N_15371,N_15709);
or U16443 (N_16443,N_15248,N_15085);
nand U16444 (N_16444,N_15630,N_15646);
xnor U16445 (N_16445,N_15944,N_15591);
or U16446 (N_16446,N_16027,N_15209);
or U16447 (N_16447,N_15271,N_15757);
or U16448 (N_16448,N_15684,N_15332);
xnor U16449 (N_16449,N_15249,N_15390);
nor U16450 (N_16450,N_15396,N_15398);
nor U16451 (N_16451,N_15264,N_15880);
xor U16452 (N_16452,N_16112,N_15306);
nand U16453 (N_16453,N_15608,N_15935);
and U16454 (N_16454,N_15826,N_15373);
nand U16455 (N_16455,N_16070,N_15159);
and U16456 (N_16456,N_15860,N_16189);
nor U16457 (N_16457,N_15189,N_15569);
xnor U16458 (N_16458,N_15566,N_15222);
nor U16459 (N_16459,N_15219,N_16239);
and U16460 (N_16460,N_15939,N_15214);
and U16461 (N_16461,N_15775,N_15623);
nand U16462 (N_16462,N_15407,N_15769);
nand U16463 (N_16463,N_15124,N_15667);
nor U16464 (N_16464,N_15797,N_15780);
xnor U16465 (N_16465,N_16061,N_15678);
nor U16466 (N_16466,N_15438,N_15512);
and U16467 (N_16467,N_15251,N_15747);
xnor U16468 (N_16468,N_15534,N_16014);
nor U16469 (N_16469,N_15633,N_15338);
nand U16470 (N_16470,N_15192,N_15287);
or U16471 (N_16471,N_15841,N_16117);
or U16472 (N_16472,N_15388,N_15993);
or U16473 (N_16473,N_15040,N_15518);
and U16474 (N_16474,N_15555,N_15857);
nor U16475 (N_16475,N_15238,N_16198);
xor U16476 (N_16476,N_15161,N_15083);
and U16477 (N_16477,N_15191,N_15912);
nor U16478 (N_16478,N_15397,N_15770);
xor U16479 (N_16479,N_15643,N_16148);
xor U16480 (N_16480,N_15997,N_15899);
and U16481 (N_16481,N_16056,N_15227);
nor U16482 (N_16482,N_16032,N_15088);
xnor U16483 (N_16483,N_15451,N_15321);
nor U16484 (N_16484,N_15082,N_16090);
nor U16485 (N_16485,N_15663,N_15454);
xor U16486 (N_16486,N_15485,N_15862);
xor U16487 (N_16487,N_15557,N_15733);
nor U16488 (N_16488,N_15827,N_15272);
and U16489 (N_16489,N_15726,N_15364);
or U16490 (N_16490,N_16082,N_15893);
and U16491 (N_16491,N_15467,N_15003);
nor U16492 (N_16492,N_15700,N_15313);
xor U16493 (N_16493,N_15522,N_15041);
xnor U16494 (N_16494,N_15767,N_15550);
nor U16495 (N_16495,N_15920,N_16197);
or U16496 (N_16496,N_15218,N_15437);
and U16497 (N_16497,N_15344,N_15367);
nor U16498 (N_16498,N_16227,N_15108);
xnor U16499 (N_16499,N_15307,N_16013);
and U16500 (N_16500,N_15188,N_16140);
xnor U16501 (N_16501,N_15985,N_15981);
or U16502 (N_16502,N_15882,N_16000);
nand U16503 (N_16503,N_15668,N_15133);
xnor U16504 (N_16504,N_15991,N_16026);
nor U16505 (N_16505,N_15087,N_15926);
and U16506 (N_16506,N_15162,N_15676);
nor U16507 (N_16507,N_15524,N_15305);
nand U16508 (N_16508,N_16122,N_15683);
nand U16509 (N_16509,N_16005,N_16058);
xor U16510 (N_16510,N_16078,N_16063);
xnor U16511 (N_16511,N_16232,N_15936);
nor U16512 (N_16512,N_16127,N_15212);
nor U16513 (N_16513,N_15273,N_15320);
and U16514 (N_16514,N_16038,N_15840);
nand U16515 (N_16515,N_15058,N_15759);
and U16516 (N_16516,N_15436,N_15101);
and U16517 (N_16517,N_15331,N_15348);
nand U16518 (N_16518,N_15778,N_15056);
xor U16519 (N_16519,N_15737,N_15741);
and U16520 (N_16520,N_15198,N_15429);
nor U16521 (N_16521,N_15871,N_15404);
or U16522 (N_16522,N_15731,N_15018);
or U16523 (N_16523,N_16077,N_15128);
or U16524 (N_16524,N_15213,N_15771);
xnor U16525 (N_16525,N_15477,N_16182);
or U16526 (N_16526,N_15685,N_15861);
or U16527 (N_16527,N_15261,N_15865);
nor U16528 (N_16528,N_15870,N_16086);
nor U16529 (N_16529,N_15808,N_16049);
nand U16530 (N_16530,N_15891,N_15426);
or U16531 (N_16531,N_15489,N_15836);
and U16532 (N_16532,N_16168,N_15328);
nor U16533 (N_16533,N_16094,N_15073);
and U16534 (N_16534,N_15376,N_15804);
nand U16535 (N_16535,N_15391,N_15523);
nor U16536 (N_16536,N_15745,N_15554);
nand U16537 (N_16537,N_15145,N_16138);
or U16538 (N_16538,N_16104,N_16158);
xor U16539 (N_16539,N_15563,N_15641);
nand U16540 (N_16540,N_15205,N_16018);
or U16541 (N_16541,N_16121,N_16033);
nand U16542 (N_16542,N_15829,N_15470);
and U16543 (N_16543,N_15323,N_15626);
nand U16544 (N_16544,N_15196,N_16037);
xor U16545 (N_16545,N_15480,N_15333);
nand U16546 (N_16546,N_15792,N_15723);
nor U16547 (N_16547,N_15279,N_15319);
and U16548 (N_16548,N_15910,N_16161);
or U16549 (N_16549,N_15203,N_15418);
and U16550 (N_16550,N_15229,N_15282);
nand U16551 (N_16551,N_15236,N_15237);
nand U16552 (N_16552,N_15386,N_15652);
xor U16553 (N_16553,N_15000,N_15482);
or U16554 (N_16554,N_15130,N_15158);
or U16555 (N_16555,N_15889,N_16068);
or U16556 (N_16556,N_15560,N_16204);
or U16557 (N_16557,N_15164,N_15881);
nor U16558 (N_16558,N_15806,N_15867);
xnor U16559 (N_16559,N_15176,N_15194);
nor U16560 (N_16560,N_15224,N_15692);
nand U16561 (N_16561,N_15304,N_15742);
nor U16562 (N_16562,N_15493,N_15565);
or U16563 (N_16563,N_16004,N_15989);
or U16564 (N_16564,N_15704,N_16229);
nor U16565 (N_16565,N_15440,N_16022);
xor U16566 (N_16566,N_16089,N_15896);
and U16567 (N_16567,N_15789,N_15220);
nand U16568 (N_16568,N_15150,N_15628);
and U16569 (N_16569,N_15604,N_15370);
xnor U16570 (N_16570,N_15297,N_15744);
and U16571 (N_16571,N_15444,N_16008);
xnor U16572 (N_16572,N_15719,N_16242);
or U16573 (N_16573,N_15674,N_15508);
and U16574 (N_16574,N_15417,N_16156);
and U16575 (N_16575,N_15779,N_15603);
nand U16576 (N_16576,N_16071,N_15289);
xor U16577 (N_16577,N_16103,N_15734);
or U16578 (N_16578,N_15751,N_16021);
or U16579 (N_16579,N_15903,N_16160);
nand U16580 (N_16580,N_16181,N_15152);
nor U16581 (N_16581,N_16047,N_16114);
nor U16582 (N_16582,N_15888,N_15403);
nor U16583 (N_16583,N_15874,N_15529);
or U16584 (N_16584,N_15051,N_15768);
nor U16585 (N_16585,N_15410,N_16166);
and U16586 (N_16586,N_15854,N_15850);
nor U16587 (N_16587,N_16080,N_15448);
xor U16588 (N_16588,N_15602,N_15607);
or U16589 (N_16589,N_15497,N_15791);
or U16590 (N_16590,N_15136,N_15290);
nand U16591 (N_16591,N_15007,N_15472);
xnor U16592 (N_16592,N_15461,N_15743);
nor U16593 (N_16593,N_16111,N_15026);
nor U16594 (N_16594,N_15389,N_15462);
nand U16595 (N_16595,N_15117,N_15551);
or U16596 (N_16596,N_15648,N_16054);
and U16597 (N_16597,N_16144,N_15109);
and U16598 (N_16598,N_15090,N_15356);
nor U16599 (N_16599,N_15727,N_15141);
and U16600 (N_16600,N_15958,N_15547);
and U16601 (N_16601,N_15153,N_15707);
and U16602 (N_16602,N_15225,N_15474);
nor U16603 (N_16603,N_15107,N_15036);
nor U16604 (N_16604,N_16145,N_15027);
or U16605 (N_16605,N_15100,N_15208);
xor U16606 (N_16606,N_15748,N_15131);
and U16607 (N_16607,N_15016,N_15843);
xor U16608 (N_16608,N_15639,N_15966);
or U16609 (N_16609,N_15706,N_15819);
xor U16610 (N_16610,N_15460,N_15813);
nand U16611 (N_16611,N_16195,N_15614);
nand U16612 (N_16612,N_15766,N_15278);
nor U16613 (N_16613,N_15076,N_15969);
xnor U16614 (N_16614,N_16165,N_15844);
nor U16615 (N_16615,N_15835,N_15821);
or U16616 (N_16616,N_15675,N_15182);
nor U16617 (N_16617,N_15335,N_15228);
xnor U16618 (N_16618,N_16230,N_16045);
and U16619 (N_16619,N_15329,N_15119);
or U16620 (N_16620,N_15795,N_15017);
nand U16621 (N_16621,N_15681,N_15419);
or U16622 (N_16622,N_16215,N_15170);
xnor U16623 (N_16623,N_16167,N_15206);
or U16624 (N_16624,N_15772,N_16099);
and U16625 (N_16625,N_15043,N_15479);
or U16626 (N_16626,N_15967,N_15853);
nand U16627 (N_16627,N_16157,N_15031);
and U16628 (N_16628,N_16100,N_15151);
xor U16629 (N_16629,N_15498,N_15673);
nand U16630 (N_16630,N_15858,N_15081);
xnor U16631 (N_16631,N_15097,N_15824);
xor U16632 (N_16632,N_15635,N_15746);
nor U16633 (N_16633,N_15345,N_15509);
nand U16634 (N_16634,N_16113,N_15735);
nor U16635 (N_16635,N_16128,N_16172);
nand U16636 (N_16636,N_15496,N_15653);
xor U16637 (N_16637,N_15010,N_15050);
and U16638 (N_16638,N_15309,N_15964);
or U16639 (N_16639,N_16020,N_15301);
xnor U16640 (N_16640,N_15258,N_16162);
nand U16641 (N_16641,N_15913,N_15868);
nor U16642 (N_16642,N_15434,N_16199);
xnor U16643 (N_16643,N_16003,N_15620);
or U16644 (N_16644,N_15510,N_15855);
or U16645 (N_16645,N_16079,N_16212);
or U16646 (N_16646,N_15468,N_15257);
or U16647 (N_16647,N_16065,N_15507);
nand U16648 (N_16648,N_16098,N_16150);
nand U16649 (N_16649,N_15441,N_15353);
and U16650 (N_16650,N_16133,N_15372);
xnor U16651 (N_16651,N_15730,N_15042);
or U16652 (N_16652,N_16193,N_15394);
nand U16653 (N_16653,N_16092,N_15001);
nor U16654 (N_16654,N_15395,N_15923);
nand U16655 (N_16655,N_16007,N_15246);
and U16656 (N_16656,N_15916,N_15452);
nor U16657 (N_16657,N_15269,N_15061);
xor U16658 (N_16658,N_15021,N_15424);
xnor U16659 (N_16659,N_15245,N_15571);
and U16660 (N_16660,N_15650,N_16141);
nand U16661 (N_16661,N_16119,N_15377);
nand U16662 (N_16662,N_15260,N_15807);
nor U16663 (N_16663,N_15558,N_16050);
and U16664 (N_16664,N_15351,N_15316);
and U16665 (N_16665,N_15049,N_15139);
or U16666 (N_16666,N_15025,N_15574);
and U16667 (N_16667,N_15654,N_15181);
nand U16668 (N_16668,N_15455,N_15339);
nor U16669 (N_16669,N_15074,N_15435);
nor U16670 (N_16670,N_15038,N_15415);
xor U16671 (N_16671,N_15660,N_15693);
or U16672 (N_16672,N_15494,N_15299);
nor U16673 (N_16673,N_15664,N_16178);
xor U16674 (N_16674,N_15885,N_15471);
or U16675 (N_16675,N_15488,N_15721);
nand U16676 (N_16676,N_15235,N_16052);
or U16677 (N_16677,N_16247,N_15884);
xor U16678 (N_16678,N_15919,N_15314);
nand U16679 (N_16679,N_15284,N_15657);
and U16680 (N_16680,N_15691,N_16183);
and U16681 (N_16681,N_15573,N_15725);
nand U16682 (N_16682,N_15283,N_15300);
nor U16683 (N_16683,N_15115,N_16064);
or U16684 (N_16684,N_16146,N_16224);
nand U16685 (N_16685,N_15816,N_15014);
nor U16686 (N_16686,N_15942,N_15658);
nor U16687 (N_16687,N_15790,N_16137);
or U16688 (N_16688,N_15099,N_15822);
and U16689 (N_16689,N_15785,N_15729);
nand U16690 (N_16690,N_15102,N_15894);
and U16691 (N_16691,N_15070,N_15357);
nand U16692 (N_16692,N_15540,N_16096);
xnor U16693 (N_16693,N_15077,N_15636);
and U16694 (N_16694,N_15413,N_15175);
xor U16695 (N_16695,N_15487,N_15892);
xor U16696 (N_16696,N_15978,N_15762);
xor U16697 (N_16697,N_15937,N_15149);
nor U16698 (N_16698,N_15585,N_15157);
nand U16699 (N_16699,N_15086,N_15581);
and U16700 (N_16700,N_15114,N_15039);
and U16701 (N_16701,N_15084,N_15215);
or U16702 (N_16702,N_15266,N_15838);
xnor U16703 (N_16703,N_15263,N_15525);
and U16704 (N_16704,N_15834,N_15135);
xor U16705 (N_16705,N_15303,N_15516);
nor U16706 (N_16706,N_15447,N_15579);
xor U16707 (N_16707,N_15911,N_15484);
and U16708 (N_16708,N_15659,N_15270);
xnor U16709 (N_16709,N_16164,N_16235);
nor U16710 (N_16710,N_15952,N_15530);
or U16711 (N_16711,N_15617,N_15362);
nor U16712 (N_16712,N_15137,N_15613);
nor U16713 (N_16713,N_15986,N_15533);
and U16714 (N_16714,N_15368,N_15968);
xor U16715 (N_16715,N_15317,N_15846);
or U16716 (N_16716,N_16120,N_15995);
and U16717 (N_16717,N_15169,N_15953);
nand U16718 (N_16718,N_15392,N_15983);
nor U16719 (N_16719,N_15098,N_15982);
nand U16720 (N_16720,N_15622,N_15506);
xor U16721 (N_16721,N_16194,N_15578);
and U16722 (N_16722,N_15177,N_16236);
xor U16723 (N_16723,N_15459,N_15595);
nand U16724 (N_16724,N_15517,N_15596);
nor U16725 (N_16725,N_15425,N_15094);
nand U16726 (N_16726,N_15619,N_15715);
or U16727 (N_16727,N_15679,N_15234);
nor U16728 (N_16728,N_16081,N_15940);
xor U16729 (N_16729,N_15046,N_15340);
xnor U16730 (N_16730,N_15231,N_16110);
xor U16731 (N_16731,N_16248,N_15055);
xor U16732 (N_16732,N_15548,N_15948);
xnor U16733 (N_16733,N_15179,N_15941);
xnor U16734 (N_16734,N_15449,N_15618);
or U16735 (N_16735,N_16218,N_15002);
xor U16736 (N_16736,N_15631,N_15168);
and U16737 (N_16737,N_15267,N_15900);
and U16738 (N_16738,N_15337,N_15934);
or U16739 (N_16739,N_15544,N_15793);
nand U16740 (N_16740,N_15143,N_16055);
xor U16741 (N_16741,N_15586,N_15428);
and U16742 (N_16742,N_15812,N_15929);
nor U16743 (N_16743,N_15308,N_15895);
or U16744 (N_16744,N_15071,N_15987);
and U16745 (N_16745,N_15195,N_15705);
nand U16746 (N_16746,N_15786,N_15716);
and U16747 (N_16747,N_16019,N_15918);
and U16748 (N_16748,N_15906,N_15644);
and U16749 (N_16749,N_15187,N_15803);
nor U16750 (N_16750,N_15690,N_15408);
nand U16751 (N_16751,N_16231,N_15616);
or U16752 (N_16752,N_15491,N_16105);
nand U16753 (N_16753,N_15627,N_15670);
xnor U16754 (N_16754,N_15318,N_16009);
and U16755 (N_16755,N_15956,N_15409);
or U16756 (N_16756,N_15075,N_15326);
or U16757 (N_16757,N_15755,N_15535);
or U16758 (N_16758,N_15917,N_15053);
or U16759 (N_16759,N_16035,N_15749);
and U16760 (N_16760,N_16073,N_15065);
xnor U16761 (N_16761,N_16115,N_16106);
nand U16762 (N_16762,N_15637,N_15649);
or U16763 (N_16763,N_15538,N_15259);
xor U16764 (N_16764,N_15172,N_15798);
nor U16765 (N_16765,N_15402,N_15064);
xor U16766 (N_16766,N_15412,N_15009);
nand U16767 (N_16767,N_15360,N_15221);
nand U16768 (N_16768,N_15606,N_15765);
and U16769 (N_16769,N_15810,N_16091);
and U16770 (N_16770,N_15879,N_15401);
and U16771 (N_16771,N_15230,N_15666);
nand U16772 (N_16772,N_16109,N_15103);
nand U16773 (N_16773,N_16184,N_15059);
nand U16774 (N_16774,N_15632,N_15963);
xor U16775 (N_16775,N_15347,N_15104);
nor U16776 (N_16776,N_15625,N_15465);
nand U16777 (N_16777,N_15703,N_15142);
xnor U16778 (N_16778,N_15093,N_15256);
and U16779 (N_16779,N_15211,N_15233);
nor U16780 (N_16780,N_15932,N_15873);
nor U16781 (N_16781,N_15029,N_15869);
xnor U16782 (N_16782,N_15784,N_15924);
and U16783 (N_16783,N_15311,N_15399);
nor U16784 (N_16784,N_15866,N_15062);
and U16785 (N_16785,N_15400,N_16222);
xor U16786 (N_16786,N_15111,N_16059);
and U16787 (N_16787,N_15315,N_15736);
or U16788 (N_16788,N_15047,N_15174);
and U16789 (N_16789,N_15277,N_15930);
or U16790 (N_16790,N_15432,N_15575);
or U16791 (N_16791,N_15949,N_15383);
xnor U16792 (N_16792,N_15476,N_15366);
or U16793 (N_16793,N_16217,N_15382);
or U16794 (N_16794,N_15593,N_15005);
and U16795 (N_16795,N_15972,N_16093);
or U16796 (N_16796,N_15589,N_15416);
xnor U16797 (N_16797,N_15914,N_15116);
nand U16798 (N_16798,N_15984,N_15561);
or U16799 (N_16799,N_15173,N_16234);
nor U16800 (N_16800,N_16237,N_16223);
xnor U16801 (N_16801,N_16066,N_15223);
or U16802 (N_16802,N_15240,N_15564);
nand U16803 (N_16803,N_15030,N_15724);
and U16804 (N_16804,N_15322,N_15999);
and U16805 (N_16805,N_15542,N_15582);
nand U16806 (N_16806,N_15921,N_15962);
xor U16807 (N_16807,N_15689,N_15361);
nor U16808 (N_16808,N_15959,N_16171);
nand U16809 (N_16809,N_15527,N_16028);
or U16810 (N_16810,N_15019,N_15890);
xor U16811 (N_16811,N_15883,N_15638);
and U16812 (N_16812,N_15655,N_15802);
and U16813 (N_16813,N_15708,N_15965);
or U16814 (N_16814,N_15680,N_15656);
nor U16815 (N_16815,N_15761,N_15121);
nor U16816 (N_16816,N_16048,N_15295);
xnor U16817 (N_16817,N_15148,N_15453);
nand U16818 (N_16818,N_16207,N_15197);
nor U16819 (N_16819,N_15160,N_15132);
or U16820 (N_16820,N_15839,N_16060);
or U16821 (N_16821,N_15439,N_15994);
nor U16822 (N_16822,N_16238,N_15960);
nor U16823 (N_16823,N_15763,N_15204);
or U16824 (N_16824,N_15184,N_15799);
nand U16825 (N_16825,N_16036,N_15511);
or U16826 (N_16826,N_16187,N_15961);
and U16827 (N_16827,N_16029,N_16083);
and U16828 (N_16828,N_15528,N_15971);
or U16829 (N_16829,N_15669,N_15033);
xnor U16830 (N_16830,N_15385,N_15594);
nor U16831 (N_16831,N_15562,N_15291);
or U16832 (N_16832,N_15034,N_15980);
nor U16833 (N_16833,N_16062,N_15250);
or U16834 (N_16834,N_15163,N_15583);
nor U16835 (N_16835,N_15847,N_15200);
xnor U16836 (N_16836,N_15532,N_16186);
nor U16837 (N_16837,N_16208,N_15254);
nor U16838 (N_16838,N_15577,N_15740);
nand U16839 (N_16839,N_15092,N_15427);
nand U16840 (N_16840,N_16159,N_15686);
nor U16841 (N_16841,N_16116,N_15898);
nand U16842 (N_16842,N_16118,N_15422);
xor U16843 (N_16843,N_15035,N_15393);
nand U16844 (N_16844,N_15346,N_15760);
and U16845 (N_16845,N_15849,N_15069);
or U16846 (N_16846,N_15032,N_16175);
and U16847 (N_16847,N_15458,N_15105);
nand U16848 (N_16848,N_15856,N_15825);
and U16849 (N_16849,N_15601,N_15682);
nand U16850 (N_16850,N_15298,N_15774);
nand U16851 (N_16851,N_15294,N_15851);
nand U16852 (N_16852,N_16001,N_15722);
or U16853 (N_16853,N_15702,N_15782);
or U16854 (N_16854,N_15146,N_16017);
nand U16855 (N_16855,N_15832,N_15171);
nor U16856 (N_16856,N_15698,N_15990);
nor U16857 (N_16857,N_16097,N_16154);
nor U16858 (N_16858,N_15513,N_15445);
nand U16859 (N_16859,N_15015,N_15588);
xnor U16860 (N_16860,N_15951,N_15605);
and U16861 (N_16861,N_16220,N_16025);
nand U16862 (N_16862,N_15556,N_15568);
nor U16863 (N_16863,N_15833,N_15800);
or U16864 (N_16864,N_15140,N_15405);
and U16865 (N_16865,N_15818,N_16044);
xnor U16866 (N_16866,N_15701,N_15456);
nor U16867 (N_16867,N_15155,N_16233);
or U16868 (N_16868,N_15651,N_15350);
xnor U16869 (N_16869,N_15611,N_15144);
nor U16870 (N_16870,N_15904,N_16177);
xor U16871 (N_16871,N_16015,N_15242);
or U16872 (N_16872,N_16041,N_16152);
nor U16873 (N_16873,N_15609,N_15274);
or U16874 (N_16874,N_16126,N_15584);
xor U16875 (N_16875,N_15560,N_16116);
and U16876 (N_16876,N_15316,N_15817);
and U16877 (N_16877,N_16192,N_15610);
nand U16878 (N_16878,N_15099,N_15399);
or U16879 (N_16879,N_15532,N_15953);
nor U16880 (N_16880,N_15357,N_15161);
nor U16881 (N_16881,N_15975,N_16129);
or U16882 (N_16882,N_15428,N_15052);
and U16883 (N_16883,N_15733,N_15254);
or U16884 (N_16884,N_15216,N_15008);
xor U16885 (N_16885,N_15071,N_15509);
xnor U16886 (N_16886,N_15222,N_15434);
or U16887 (N_16887,N_15360,N_15359);
nand U16888 (N_16888,N_15707,N_16036);
and U16889 (N_16889,N_15329,N_15149);
xnor U16890 (N_16890,N_15373,N_16138);
nor U16891 (N_16891,N_15380,N_15674);
xnor U16892 (N_16892,N_16131,N_15408);
or U16893 (N_16893,N_15915,N_15936);
nand U16894 (N_16894,N_16208,N_16079);
xnor U16895 (N_16895,N_15634,N_16055);
xnor U16896 (N_16896,N_15572,N_15829);
xor U16897 (N_16897,N_15294,N_15857);
or U16898 (N_16898,N_15995,N_15086);
or U16899 (N_16899,N_15213,N_15899);
or U16900 (N_16900,N_15630,N_15339);
or U16901 (N_16901,N_15437,N_15885);
xor U16902 (N_16902,N_16001,N_15813);
or U16903 (N_16903,N_15361,N_15682);
and U16904 (N_16904,N_16164,N_15064);
or U16905 (N_16905,N_15903,N_15038);
xor U16906 (N_16906,N_15800,N_15359);
or U16907 (N_16907,N_15865,N_16159);
nor U16908 (N_16908,N_15633,N_15417);
and U16909 (N_16909,N_15312,N_16156);
and U16910 (N_16910,N_15600,N_15374);
xor U16911 (N_16911,N_15882,N_16068);
xor U16912 (N_16912,N_15373,N_15457);
and U16913 (N_16913,N_16064,N_15927);
nor U16914 (N_16914,N_15152,N_15615);
nor U16915 (N_16915,N_15563,N_15007);
nor U16916 (N_16916,N_15408,N_16161);
or U16917 (N_16917,N_15974,N_15225);
nor U16918 (N_16918,N_15880,N_15269);
nor U16919 (N_16919,N_15907,N_15208);
or U16920 (N_16920,N_15112,N_15411);
xor U16921 (N_16921,N_15044,N_15939);
nand U16922 (N_16922,N_15150,N_15138);
and U16923 (N_16923,N_15262,N_15034);
nor U16924 (N_16924,N_15893,N_15626);
nand U16925 (N_16925,N_15367,N_15397);
nor U16926 (N_16926,N_15269,N_15291);
nor U16927 (N_16927,N_15280,N_16091);
or U16928 (N_16928,N_15530,N_15043);
xnor U16929 (N_16929,N_15143,N_15242);
or U16930 (N_16930,N_15391,N_15076);
and U16931 (N_16931,N_15682,N_15017);
nand U16932 (N_16932,N_15715,N_16206);
nor U16933 (N_16933,N_15273,N_15428);
nor U16934 (N_16934,N_15576,N_15458);
or U16935 (N_16935,N_15571,N_15401);
nand U16936 (N_16936,N_15110,N_15576);
nand U16937 (N_16937,N_15881,N_15536);
or U16938 (N_16938,N_15504,N_15653);
nand U16939 (N_16939,N_16153,N_15911);
nand U16940 (N_16940,N_15515,N_15774);
or U16941 (N_16941,N_16205,N_16085);
nor U16942 (N_16942,N_16057,N_15631);
xnor U16943 (N_16943,N_15451,N_15733);
and U16944 (N_16944,N_15603,N_15543);
nand U16945 (N_16945,N_15155,N_15168);
nand U16946 (N_16946,N_15973,N_15877);
nand U16947 (N_16947,N_16068,N_15101);
nor U16948 (N_16948,N_15013,N_15420);
and U16949 (N_16949,N_15510,N_16125);
nor U16950 (N_16950,N_15579,N_15480);
xnor U16951 (N_16951,N_15955,N_15672);
xnor U16952 (N_16952,N_15856,N_16111);
or U16953 (N_16953,N_15845,N_15144);
nor U16954 (N_16954,N_15030,N_15060);
nor U16955 (N_16955,N_15809,N_16240);
nor U16956 (N_16956,N_15668,N_16015);
or U16957 (N_16957,N_15021,N_15395);
or U16958 (N_16958,N_16181,N_16056);
xor U16959 (N_16959,N_15092,N_15874);
nand U16960 (N_16960,N_15839,N_16144);
nor U16961 (N_16961,N_15265,N_16071);
or U16962 (N_16962,N_15287,N_16188);
and U16963 (N_16963,N_16175,N_15815);
or U16964 (N_16964,N_16229,N_15254);
nor U16965 (N_16965,N_16117,N_15942);
or U16966 (N_16966,N_16229,N_15425);
or U16967 (N_16967,N_15015,N_15536);
xnor U16968 (N_16968,N_15697,N_15330);
xnor U16969 (N_16969,N_15344,N_16159);
and U16970 (N_16970,N_15470,N_15316);
xor U16971 (N_16971,N_16172,N_15715);
nand U16972 (N_16972,N_15682,N_15764);
xnor U16973 (N_16973,N_16046,N_15218);
nand U16974 (N_16974,N_15435,N_15478);
and U16975 (N_16975,N_15499,N_15385);
nand U16976 (N_16976,N_15736,N_15865);
nand U16977 (N_16977,N_15730,N_15171);
nand U16978 (N_16978,N_15921,N_15404);
or U16979 (N_16979,N_15952,N_15552);
and U16980 (N_16980,N_15183,N_16104);
nor U16981 (N_16981,N_16213,N_16246);
nand U16982 (N_16982,N_15508,N_15790);
nand U16983 (N_16983,N_16245,N_15044);
or U16984 (N_16984,N_15398,N_15380);
nor U16985 (N_16985,N_15855,N_15818);
xnor U16986 (N_16986,N_15065,N_15387);
nand U16987 (N_16987,N_15585,N_15333);
nand U16988 (N_16988,N_15765,N_15668);
nor U16989 (N_16989,N_16209,N_15612);
nand U16990 (N_16990,N_15309,N_15815);
nand U16991 (N_16991,N_15744,N_16088);
nand U16992 (N_16992,N_15125,N_15004);
xor U16993 (N_16993,N_15975,N_15653);
xnor U16994 (N_16994,N_16232,N_15889);
xor U16995 (N_16995,N_15274,N_15130);
or U16996 (N_16996,N_16145,N_15930);
or U16997 (N_16997,N_16224,N_15939);
nand U16998 (N_16998,N_16176,N_15732);
xor U16999 (N_16999,N_15815,N_15352);
nor U17000 (N_17000,N_15707,N_16208);
nor U17001 (N_17001,N_15588,N_15353);
xor U17002 (N_17002,N_15930,N_15794);
nand U17003 (N_17003,N_16025,N_15134);
nor U17004 (N_17004,N_15875,N_16004);
nor U17005 (N_17005,N_15942,N_15356);
and U17006 (N_17006,N_15445,N_15544);
nand U17007 (N_17007,N_15133,N_15822);
or U17008 (N_17008,N_15985,N_15964);
nor U17009 (N_17009,N_15483,N_15668);
or U17010 (N_17010,N_15504,N_15472);
nand U17011 (N_17011,N_15825,N_15226);
and U17012 (N_17012,N_15294,N_15719);
xor U17013 (N_17013,N_15152,N_15262);
nor U17014 (N_17014,N_15102,N_16230);
and U17015 (N_17015,N_16121,N_15341);
nand U17016 (N_17016,N_15770,N_15659);
xnor U17017 (N_17017,N_16075,N_15192);
and U17018 (N_17018,N_15593,N_15525);
or U17019 (N_17019,N_15953,N_15099);
and U17020 (N_17020,N_15105,N_15701);
xor U17021 (N_17021,N_15122,N_15346);
or U17022 (N_17022,N_16013,N_15431);
xor U17023 (N_17023,N_15412,N_15012);
and U17024 (N_17024,N_16155,N_15983);
or U17025 (N_17025,N_15972,N_16197);
xnor U17026 (N_17026,N_16078,N_15254);
nor U17027 (N_17027,N_15919,N_16238);
xnor U17028 (N_17028,N_16227,N_15520);
or U17029 (N_17029,N_16137,N_15534);
and U17030 (N_17030,N_15741,N_15642);
nor U17031 (N_17031,N_15506,N_15119);
nor U17032 (N_17032,N_15746,N_15895);
xnor U17033 (N_17033,N_15812,N_16146);
or U17034 (N_17034,N_15481,N_15312);
and U17035 (N_17035,N_15356,N_15112);
xnor U17036 (N_17036,N_15459,N_15932);
xor U17037 (N_17037,N_15108,N_15528);
xnor U17038 (N_17038,N_16033,N_15218);
and U17039 (N_17039,N_16023,N_15820);
and U17040 (N_17040,N_16236,N_15132);
or U17041 (N_17041,N_15270,N_15425);
or U17042 (N_17042,N_15806,N_15710);
or U17043 (N_17043,N_15296,N_15286);
xnor U17044 (N_17044,N_15574,N_15857);
nor U17045 (N_17045,N_15296,N_15148);
nand U17046 (N_17046,N_15437,N_16176);
or U17047 (N_17047,N_15918,N_15201);
nand U17048 (N_17048,N_16230,N_15933);
and U17049 (N_17049,N_15624,N_15126);
nand U17050 (N_17050,N_15674,N_15894);
or U17051 (N_17051,N_15856,N_16114);
or U17052 (N_17052,N_15398,N_16110);
and U17053 (N_17053,N_15611,N_15854);
or U17054 (N_17054,N_15470,N_16013);
and U17055 (N_17055,N_15109,N_15797);
nand U17056 (N_17056,N_15018,N_15700);
or U17057 (N_17057,N_15084,N_15375);
xor U17058 (N_17058,N_16115,N_15730);
nand U17059 (N_17059,N_15329,N_15291);
nor U17060 (N_17060,N_16071,N_15246);
and U17061 (N_17061,N_15259,N_15248);
and U17062 (N_17062,N_16206,N_16222);
nand U17063 (N_17063,N_15190,N_15212);
nor U17064 (N_17064,N_15157,N_16105);
nand U17065 (N_17065,N_16141,N_15805);
nand U17066 (N_17066,N_15519,N_15520);
nand U17067 (N_17067,N_16084,N_15113);
xor U17068 (N_17068,N_15023,N_15781);
and U17069 (N_17069,N_15239,N_15682);
nor U17070 (N_17070,N_15037,N_15737);
xor U17071 (N_17071,N_15456,N_15601);
or U17072 (N_17072,N_16114,N_15199);
and U17073 (N_17073,N_15872,N_15903);
and U17074 (N_17074,N_15142,N_15646);
nor U17075 (N_17075,N_15370,N_15679);
and U17076 (N_17076,N_15211,N_15901);
xor U17077 (N_17077,N_15327,N_15846);
xor U17078 (N_17078,N_15797,N_15331);
nand U17079 (N_17079,N_16134,N_15370);
nor U17080 (N_17080,N_15018,N_15528);
or U17081 (N_17081,N_15824,N_15506);
and U17082 (N_17082,N_15607,N_15713);
nor U17083 (N_17083,N_15212,N_15994);
and U17084 (N_17084,N_15383,N_15366);
or U17085 (N_17085,N_16236,N_15667);
nand U17086 (N_17086,N_15940,N_15376);
xor U17087 (N_17087,N_15096,N_15811);
nand U17088 (N_17088,N_16057,N_16044);
and U17089 (N_17089,N_16100,N_15267);
nand U17090 (N_17090,N_15910,N_15832);
xnor U17091 (N_17091,N_15695,N_15764);
nor U17092 (N_17092,N_15425,N_16143);
xor U17093 (N_17093,N_15551,N_15647);
xor U17094 (N_17094,N_16114,N_16023);
nand U17095 (N_17095,N_15517,N_15074);
and U17096 (N_17096,N_15420,N_15368);
nor U17097 (N_17097,N_15092,N_15547);
and U17098 (N_17098,N_16012,N_15202);
xnor U17099 (N_17099,N_15698,N_16014);
nand U17100 (N_17100,N_15295,N_15350);
nand U17101 (N_17101,N_16020,N_15616);
nor U17102 (N_17102,N_15992,N_15550);
nand U17103 (N_17103,N_15906,N_16198);
xor U17104 (N_17104,N_15275,N_15045);
nor U17105 (N_17105,N_16104,N_15859);
nor U17106 (N_17106,N_15143,N_15472);
nand U17107 (N_17107,N_15251,N_15854);
xnor U17108 (N_17108,N_16099,N_15688);
xor U17109 (N_17109,N_16041,N_15250);
nand U17110 (N_17110,N_15666,N_15346);
nor U17111 (N_17111,N_15970,N_15002);
nand U17112 (N_17112,N_16106,N_15698);
xnor U17113 (N_17113,N_15356,N_15281);
xor U17114 (N_17114,N_15612,N_15406);
nor U17115 (N_17115,N_16213,N_15622);
nand U17116 (N_17116,N_15627,N_15214);
nand U17117 (N_17117,N_15193,N_15223);
xnor U17118 (N_17118,N_16043,N_15226);
nor U17119 (N_17119,N_15070,N_16141);
nor U17120 (N_17120,N_16046,N_15523);
nor U17121 (N_17121,N_15929,N_15078);
and U17122 (N_17122,N_15851,N_15509);
xor U17123 (N_17123,N_15696,N_15537);
and U17124 (N_17124,N_16141,N_15208);
nand U17125 (N_17125,N_15404,N_15727);
and U17126 (N_17126,N_16201,N_15339);
xor U17127 (N_17127,N_15605,N_15757);
nor U17128 (N_17128,N_15538,N_16116);
xnor U17129 (N_17129,N_16172,N_15245);
or U17130 (N_17130,N_16036,N_15125);
or U17131 (N_17131,N_16062,N_15693);
and U17132 (N_17132,N_15944,N_15362);
or U17133 (N_17133,N_15309,N_15344);
nor U17134 (N_17134,N_16134,N_16159);
nand U17135 (N_17135,N_15102,N_16244);
or U17136 (N_17136,N_16057,N_15857);
nor U17137 (N_17137,N_15886,N_15980);
nand U17138 (N_17138,N_15489,N_16048);
nor U17139 (N_17139,N_15789,N_16032);
nor U17140 (N_17140,N_15295,N_15359);
nor U17141 (N_17141,N_15926,N_15350);
or U17142 (N_17142,N_15846,N_15854);
nor U17143 (N_17143,N_15565,N_15715);
or U17144 (N_17144,N_15913,N_15611);
nor U17145 (N_17145,N_15318,N_15636);
or U17146 (N_17146,N_15095,N_16009);
nor U17147 (N_17147,N_15345,N_15286);
or U17148 (N_17148,N_16211,N_15195);
or U17149 (N_17149,N_15281,N_15605);
nor U17150 (N_17150,N_16232,N_15392);
and U17151 (N_17151,N_16207,N_15002);
or U17152 (N_17152,N_15209,N_15848);
nor U17153 (N_17153,N_15370,N_15895);
or U17154 (N_17154,N_15599,N_15898);
xnor U17155 (N_17155,N_15254,N_15276);
or U17156 (N_17156,N_15727,N_16229);
nand U17157 (N_17157,N_16073,N_15393);
xnor U17158 (N_17158,N_15608,N_15345);
nand U17159 (N_17159,N_16040,N_15516);
or U17160 (N_17160,N_15287,N_15992);
nor U17161 (N_17161,N_15774,N_15359);
nand U17162 (N_17162,N_15206,N_16214);
nand U17163 (N_17163,N_15175,N_15223);
nand U17164 (N_17164,N_15621,N_15960);
or U17165 (N_17165,N_15388,N_15670);
nand U17166 (N_17166,N_15828,N_15583);
and U17167 (N_17167,N_15470,N_15396);
nor U17168 (N_17168,N_15965,N_16106);
and U17169 (N_17169,N_15005,N_15961);
or U17170 (N_17170,N_15619,N_16237);
and U17171 (N_17171,N_15284,N_15581);
or U17172 (N_17172,N_15411,N_15912);
or U17173 (N_17173,N_15786,N_15037);
and U17174 (N_17174,N_15872,N_16237);
nand U17175 (N_17175,N_15586,N_15695);
xnor U17176 (N_17176,N_15030,N_16066);
nand U17177 (N_17177,N_15306,N_15509);
xor U17178 (N_17178,N_16130,N_15828);
nand U17179 (N_17179,N_15776,N_15579);
xnor U17180 (N_17180,N_15788,N_15971);
or U17181 (N_17181,N_15841,N_16233);
and U17182 (N_17182,N_15522,N_15450);
and U17183 (N_17183,N_16074,N_16195);
and U17184 (N_17184,N_15988,N_15042);
nor U17185 (N_17185,N_15098,N_15967);
and U17186 (N_17186,N_15435,N_15445);
nor U17187 (N_17187,N_15460,N_15925);
xnor U17188 (N_17188,N_16241,N_16038);
and U17189 (N_17189,N_15700,N_15273);
and U17190 (N_17190,N_15391,N_15667);
or U17191 (N_17191,N_15466,N_16244);
and U17192 (N_17192,N_15514,N_15041);
nor U17193 (N_17193,N_15117,N_16122);
or U17194 (N_17194,N_15023,N_15273);
xnor U17195 (N_17195,N_15083,N_16059);
nor U17196 (N_17196,N_15962,N_15230);
and U17197 (N_17197,N_15115,N_16114);
nand U17198 (N_17198,N_15847,N_16180);
nor U17199 (N_17199,N_15626,N_15570);
nor U17200 (N_17200,N_16125,N_15503);
xnor U17201 (N_17201,N_15222,N_15058);
or U17202 (N_17202,N_15765,N_16059);
and U17203 (N_17203,N_15975,N_15892);
nand U17204 (N_17204,N_15114,N_15696);
nand U17205 (N_17205,N_15475,N_15258);
xor U17206 (N_17206,N_15588,N_15156);
xor U17207 (N_17207,N_15055,N_15746);
or U17208 (N_17208,N_15079,N_16013);
xor U17209 (N_17209,N_15451,N_15214);
or U17210 (N_17210,N_15102,N_16112);
xor U17211 (N_17211,N_16220,N_15526);
nor U17212 (N_17212,N_15866,N_15130);
or U17213 (N_17213,N_15937,N_15370);
and U17214 (N_17214,N_15285,N_15317);
and U17215 (N_17215,N_15277,N_15792);
nand U17216 (N_17216,N_16110,N_15271);
nor U17217 (N_17217,N_15099,N_15041);
xor U17218 (N_17218,N_16103,N_15860);
nand U17219 (N_17219,N_15106,N_16183);
nand U17220 (N_17220,N_15385,N_15258);
and U17221 (N_17221,N_15522,N_16088);
nor U17222 (N_17222,N_15792,N_15766);
or U17223 (N_17223,N_16219,N_16132);
nand U17224 (N_17224,N_15323,N_15326);
or U17225 (N_17225,N_15248,N_15039);
nand U17226 (N_17226,N_15350,N_15999);
nand U17227 (N_17227,N_15129,N_16085);
xor U17228 (N_17228,N_15032,N_16183);
and U17229 (N_17229,N_15347,N_15231);
nor U17230 (N_17230,N_15812,N_15206);
nor U17231 (N_17231,N_15081,N_15928);
xor U17232 (N_17232,N_15308,N_15694);
nand U17233 (N_17233,N_15839,N_15838);
nand U17234 (N_17234,N_15201,N_15823);
nor U17235 (N_17235,N_16179,N_15003);
nand U17236 (N_17236,N_15672,N_16197);
and U17237 (N_17237,N_15141,N_15929);
and U17238 (N_17238,N_16070,N_16100);
nor U17239 (N_17239,N_15067,N_15006);
and U17240 (N_17240,N_15887,N_15213);
or U17241 (N_17241,N_15194,N_15629);
xor U17242 (N_17242,N_15505,N_15696);
nand U17243 (N_17243,N_15721,N_15417);
nor U17244 (N_17244,N_16240,N_15004);
xor U17245 (N_17245,N_15729,N_15728);
nor U17246 (N_17246,N_16241,N_15735);
nor U17247 (N_17247,N_15710,N_15532);
or U17248 (N_17248,N_15764,N_16124);
nand U17249 (N_17249,N_15593,N_15568);
nand U17250 (N_17250,N_15635,N_15319);
xor U17251 (N_17251,N_15029,N_15961);
nand U17252 (N_17252,N_15531,N_15679);
and U17253 (N_17253,N_15234,N_15567);
and U17254 (N_17254,N_16243,N_15660);
and U17255 (N_17255,N_15242,N_15735);
nand U17256 (N_17256,N_15200,N_15999);
nor U17257 (N_17257,N_15099,N_15034);
and U17258 (N_17258,N_15998,N_15079);
and U17259 (N_17259,N_15744,N_15869);
or U17260 (N_17260,N_15452,N_16126);
nor U17261 (N_17261,N_15559,N_15444);
nand U17262 (N_17262,N_15916,N_15925);
nand U17263 (N_17263,N_15693,N_15582);
nor U17264 (N_17264,N_15986,N_16106);
nor U17265 (N_17265,N_15263,N_15951);
or U17266 (N_17266,N_15305,N_15184);
or U17267 (N_17267,N_15298,N_15134);
and U17268 (N_17268,N_16097,N_16095);
nand U17269 (N_17269,N_16198,N_15614);
and U17270 (N_17270,N_15231,N_15409);
nand U17271 (N_17271,N_15568,N_15736);
nor U17272 (N_17272,N_15468,N_16105);
nor U17273 (N_17273,N_15154,N_15963);
nor U17274 (N_17274,N_15586,N_16245);
and U17275 (N_17275,N_15531,N_15201);
or U17276 (N_17276,N_15826,N_15965);
or U17277 (N_17277,N_15157,N_15424);
nand U17278 (N_17278,N_15284,N_15631);
or U17279 (N_17279,N_15312,N_15012);
or U17280 (N_17280,N_15265,N_15225);
or U17281 (N_17281,N_15828,N_15363);
or U17282 (N_17282,N_16102,N_15355);
nand U17283 (N_17283,N_15293,N_15303);
xnor U17284 (N_17284,N_15630,N_15238);
and U17285 (N_17285,N_16173,N_15125);
nor U17286 (N_17286,N_15886,N_15707);
xnor U17287 (N_17287,N_15289,N_15032);
xor U17288 (N_17288,N_15207,N_15615);
xnor U17289 (N_17289,N_16135,N_16178);
and U17290 (N_17290,N_15023,N_15983);
xor U17291 (N_17291,N_15932,N_15434);
nand U17292 (N_17292,N_15523,N_16163);
xor U17293 (N_17293,N_15106,N_15864);
xnor U17294 (N_17294,N_15121,N_15077);
xor U17295 (N_17295,N_16145,N_15013);
xnor U17296 (N_17296,N_15894,N_16004);
and U17297 (N_17297,N_15565,N_15079);
or U17298 (N_17298,N_15030,N_15559);
nor U17299 (N_17299,N_15110,N_15899);
nand U17300 (N_17300,N_15965,N_15772);
and U17301 (N_17301,N_15934,N_15915);
nor U17302 (N_17302,N_15236,N_16173);
and U17303 (N_17303,N_15064,N_15085);
nor U17304 (N_17304,N_15926,N_16121);
and U17305 (N_17305,N_15483,N_15060);
nor U17306 (N_17306,N_15487,N_15369);
nand U17307 (N_17307,N_15267,N_16199);
nand U17308 (N_17308,N_15864,N_15397);
or U17309 (N_17309,N_15743,N_15290);
and U17310 (N_17310,N_15151,N_15028);
or U17311 (N_17311,N_15796,N_16018);
or U17312 (N_17312,N_15493,N_15936);
nand U17313 (N_17313,N_15628,N_15404);
or U17314 (N_17314,N_15727,N_15173);
and U17315 (N_17315,N_15586,N_15597);
or U17316 (N_17316,N_16074,N_15190);
xnor U17317 (N_17317,N_15659,N_15116);
or U17318 (N_17318,N_15655,N_15104);
and U17319 (N_17319,N_15716,N_15328);
or U17320 (N_17320,N_15121,N_16046);
and U17321 (N_17321,N_15591,N_15559);
xnor U17322 (N_17322,N_15550,N_15636);
xor U17323 (N_17323,N_15860,N_15009);
and U17324 (N_17324,N_15629,N_15108);
or U17325 (N_17325,N_15623,N_15038);
or U17326 (N_17326,N_16051,N_15554);
and U17327 (N_17327,N_15442,N_16189);
nor U17328 (N_17328,N_16076,N_15422);
nand U17329 (N_17329,N_15678,N_15739);
and U17330 (N_17330,N_15918,N_15049);
nor U17331 (N_17331,N_15370,N_15050);
nand U17332 (N_17332,N_15281,N_15800);
nor U17333 (N_17333,N_15864,N_15828);
nand U17334 (N_17334,N_15781,N_15062);
xnor U17335 (N_17335,N_16001,N_15888);
nor U17336 (N_17336,N_15585,N_15714);
and U17337 (N_17337,N_15135,N_15040);
nor U17338 (N_17338,N_15612,N_15384);
or U17339 (N_17339,N_16077,N_15389);
or U17340 (N_17340,N_15867,N_15200);
or U17341 (N_17341,N_15146,N_15532);
nor U17342 (N_17342,N_15650,N_15237);
nor U17343 (N_17343,N_15327,N_16110);
nand U17344 (N_17344,N_15948,N_15852);
nand U17345 (N_17345,N_16168,N_15750);
or U17346 (N_17346,N_15447,N_15847);
nor U17347 (N_17347,N_15601,N_15273);
xnor U17348 (N_17348,N_15497,N_15499);
and U17349 (N_17349,N_15914,N_16077);
and U17350 (N_17350,N_15885,N_15307);
or U17351 (N_17351,N_15472,N_15213);
and U17352 (N_17352,N_15781,N_15867);
and U17353 (N_17353,N_15456,N_15873);
xnor U17354 (N_17354,N_15220,N_15443);
or U17355 (N_17355,N_15159,N_16164);
nor U17356 (N_17356,N_16175,N_16202);
and U17357 (N_17357,N_16007,N_15613);
or U17358 (N_17358,N_15017,N_15811);
nor U17359 (N_17359,N_15395,N_15595);
xnor U17360 (N_17360,N_15344,N_15825);
nor U17361 (N_17361,N_15673,N_15476);
nand U17362 (N_17362,N_15223,N_16174);
xor U17363 (N_17363,N_15227,N_15409);
and U17364 (N_17364,N_15292,N_15685);
nor U17365 (N_17365,N_15159,N_16248);
and U17366 (N_17366,N_16032,N_16079);
nand U17367 (N_17367,N_15054,N_16249);
nand U17368 (N_17368,N_15013,N_15159);
and U17369 (N_17369,N_15508,N_15003);
nor U17370 (N_17370,N_15699,N_15597);
nor U17371 (N_17371,N_15192,N_15968);
nand U17372 (N_17372,N_15031,N_15346);
or U17373 (N_17373,N_16160,N_16162);
xor U17374 (N_17374,N_16188,N_15065);
nand U17375 (N_17375,N_15865,N_15914);
and U17376 (N_17376,N_15676,N_15405);
or U17377 (N_17377,N_15186,N_15381);
nand U17378 (N_17378,N_15177,N_15140);
and U17379 (N_17379,N_15372,N_15995);
nand U17380 (N_17380,N_15335,N_15146);
xnor U17381 (N_17381,N_16089,N_15045);
nand U17382 (N_17382,N_15073,N_15525);
or U17383 (N_17383,N_15605,N_15257);
and U17384 (N_17384,N_16072,N_16241);
nand U17385 (N_17385,N_15525,N_15192);
nor U17386 (N_17386,N_15104,N_15802);
nand U17387 (N_17387,N_15838,N_16033);
xnor U17388 (N_17388,N_16071,N_15773);
xnor U17389 (N_17389,N_15755,N_15646);
or U17390 (N_17390,N_15579,N_15607);
and U17391 (N_17391,N_15320,N_15140);
nand U17392 (N_17392,N_15197,N_15257);
nor U17393 (N_17393,N_15662,N_15048);
or U17394 (N_17394,N_15453,N_15813);
or U17395 (N_17395,N_15745,N_15107);
nand U17396 (N_17396,N_15822,N_15750);
nand U17397 (N_17397,N_15088,N_15309);
xor U17398 (N_17398,N_15276,N_16148);
xnor U17399 (N_17399,N_15249,N_15955);
or U17400 (N_17400,N_15154,N_15805);
and U17401 (N_17401,N_15666,N_15660);
and U17402 (N_17402,N_16159,N_16073);
nor U17403 (N_17403,N_15952,N_16003);
or U17404 (N_17404,N_15805,N_15009);
nor U17405 (N_17405,N_16143,N_15848);
xor U17406 (N_17406,N_16211,N_15720);
and U17407 (N_17407,N_15777,N_16162);
xnor U17408 (N_17408,N_15472,N_15059);
and U17409 (N_17409,N_16246,N_15311);
xor U17410 (N_17410,N_15505,N_15521);
nand U17411 (N_17411,N_15726,N_15789);
nor U17412 (N_17412,N_15260,N_15366);
nand U17413 (N_17413,N_16221,N_15907);
and U17414 (N_17414,N_15106,N_15211);
or U17415 (N_17415,N_15256,N_16145);
xnor U17416 (N_17416,N_15368,N_15165);
nor U17417 (N_17417,N_16062,N_15758);
nand U17418 (N_17418,N_16247,N_15896);
and U17419 (N_17419,N_15897,N_16124);
nand U17420 (N_17420,N_15872,N_15415);
or U17421 (N_17421,N_15249,N_15915);
or U17422 (N_17422,N_15644,N_15593);
nor U17423 (N_17423,N_16024,N_15430);
xor U17424 (N_17424,N_15692,N_16017);
or U17425 (N_17425,N_15045,N_15185);
or U17426 (N_17426,N_15291,N_15623);
nor U17427 (N_17427,N_15896,N_15166);
or U17428 (N_17428,N_15327,N_15495);
nor U17429 (N_17429,N_15934,N_16241);
or U17430 (N_17430,N_15179,N_15973);
and U17431 (N_17431,N_15782,N_15913);
and U17432 (N_17432,N_16182,N_15308);
xor U17433 (N_17433,N_15998,N_15394);
nor U17434 (N_17434,N_15634,N_15354);
or U17435 (N_17435,N_15288,N_15658);
nand U17436 (N_17436,N_15566,N_15745);
xor U17437 (N_17437,N_15871,N_15284);
and U17438 (N_17438,N_15510,N_15307);
nor U17439 (N_17439,N_15794,N_15427);
nor U17440 (N_17440,N_15730,N_15704);
or U17441 (N_17441,N_15581,N_15029);
or U17442 (N_17442,N_16239,N_15266);
xor U17443 (N_17443,N_15220,N_15826);
and U17444 (N_17444,N_16012,N_15425);
or U17445 (N_17445,N_15146,N_15657);
and U17446 (N_17446,N_16208,N_15741);
and U17447 (N_17447,N_15325,N_15485);
and U17448 (N_17448,N_15200,N_15759);
and U17449 (N_17449,N_15262,N_16173);
xor U17450 (N_17450,N_15371,N_15247);
nand U17451 (N_17451,N_15191,N_15418);
nor U17452 (N_17452,N_15467,N_15198);
nor U17453 (N_17453,N_15666,N_15424);
nand U17454 (N_17454,N_15026,N_15362);
xnor U17455 (N_17455,N_15136,N_16163);
nand U17456 (N_17456,N_15756,N_15257);
nand U17457 (N_17457,N_15838,N_15765);
xor U17458 (N_17458,N_15036,N_15513);
xor U17459 (N_17459,N_15303,N_15577);
nor U17460 (N_17460,N_15027,N_15903);
or U17461 (N_17461,N_16116,N_16097);
nor U17462 (N_17462,N_16010,N_15622);
xnor U17463 (N_17463,N_15631,N_15533);
and U17464 (N_17464,N_15844,N_16218);
and U17465 (N_17465,N_15469,N_15443);
nand U17466 (N_17466,N_16118,N_15300);
xnor U17467 (N_17467,N_15342,N_15351);
nand U17468 (N_17468,N_15360,N_15689);
and U17469 (N_17469,N_15438,N_15529);
xor U17470 (N_17470,N_16055,N_15990);
nor U17471 (N_17471,N_15347,N_15156);
nand U17472 (N_17472,N_15946,N_15676);
and U17473 (N_17473,N_15096,N_16017);
nand U17474 (N_17474,N_15001,N_15317);
or U17475 (N_17475,N_15696,N_15790);
or U17476 (N_17476,N_15686,N_15637);
xnor U17477 (N_17477,N_15001,N_16062);
xor U17478 (N_17478,N_15108,N_16038);
and U17479 (N_17479,N_15888,N_15466);
nand U17480 (N_17480,N_15498,N_15506);
or U17481 (N_17481,N_15738,N_15607);
and U17482 (N_17482,N_16154,N_15673);
nand U17483 (N_17483,N_16071,N_15752);
nand U17484 (N_17484,N_15430,N_15524);
xor U17485 (N_17485,N_15985,N_15628);
nand U17486 (N_17486,N_15181,N_16238);
xnor U17487 (N_17487,N_15522,N_15820);
nor U17488 (N_17488,N_15353,N_15836);
or U17489 (N_17489,N_15522,N_15381);
nor U17490 (N_17490,N_15557,N_15694);
nor U17491 (N_17491,N_15419,N_15224);
nand U17492 (N_17492,N_15225,N_15343);
and U17493 (N_17493,N_15798,N_16196);
nand U17494 (N_17494,N_15112,N_15191);
xnor U17495 (N_17495,N_15270,N_15876);
nand U17496 (N_17496,N_16229,N_16232);
nand U17497 (N_17497,N_16243,N_15648);
xor U17498 (N_17498,N_15097,N_15616);
xnor U17499 (N_17499,N_15302,N_16218);
nand U17500 (N_17500,N_17459,N_17225);
nor U17501 (N_17501,N_17446,N_16942);
nand U17502 (N_17502,N_16935,N_17261);
nand U17503 (N_17503,N_16770,N_17064);
or U17504 (N_17504,N_17266,N_16609);
and U17505 (N_17505,N_17052,N_16923);
nand U17506 (N_17506,N_17024,N_16685);
or U17507 (N_17507,N_16358,N_17027);
nor U17508 (N_17508,N_16295,N_16768);
and U17509 (N_17509,N_17496,N_16889);
xnor U17510 (N_17510,N_17205,N_17129);
nand U17511 (N_17511,N_16934,N_17499);
and U17512 (N_17512,N_16659,N_17036);
or U17513 (N_17513,N_16418,N_17196);
nand U17514 (N_17514,N_17026,N_16273);
nor U17515 (N_17515,N_16600,N_16477);
and U17516 (N_17516,N_16656,N_17330);
nor U17517 (N_17517,N_16865,N_17344);
xor U17518 (N_17518,N_16349,N_17007);
nor U17519 (N_17519,N_17452,N_16888);
and U17520 (N_17520,N_16338,N_16850);
and U17521 (N_17521,N_17479,N_17341);
xnor U17522 (N_17522,N_16779,N_17000);
nor U17523 (N_17523,N_17003,N_17062);
or U17524 (N_17524,N_16901,N_17059);
xor U17525 (N_17525,N_17079,N_17389);
and U17526 (N_17526,N_16298,N_16705);
xor U17527 (N_17527,N_16830,N_16478);
or U17528 (N_17528,N_16810,N_16846);
or U17529 (N_17529,N_17121,N_16879);
nand U17530 (N_17530,N_17489,N_16907);
xor U17531 (N_17531,N_16854,N_16410);
nand U17532 (N_17532,N_17227,N_17465);
xor U17533 (N_17533,N_17470,N_17339);
nand U17534 (N_17534,N_16252,N_16650);
or U17535 (N_17535,N_17260,N_16636);
nor U17536 (N_17536,N_16796,N_17409);
nor U17537 (N_17537,N_17427,N_16369);
xor U17538 (N_17538,N_16917,N_17136);
and U17539 (N_17539,N_17289,N_16613);
xor U17540 (N_17540,N_17233,N_16627);
xnor U17541 (N_17541,N_16933,N_17222);
and U17542 (N_17542,N_17382,N_16269);
nor U17543 (N_17543,N_17449,N_17399);
xnor U17544 (N_17544,N_17025,N_17301);
xor U17545 (N_17545,N_16937,N_17116);
xor U17546 (N_17546,N_17138,N_16325);
nor U17547 (N_17547,N_16728,N_17429);
and U17548 (N_17548,N_16419,N_17190);
xnor U17549 (N_17549,N_16582,N_17252);
or U17550 (N_17550,N_16357,N_17286);
xor U17551 (N_17551,N_16973,N_17170);
or U17552 (N_17552,N_17104,N_16672);
nand U17553 (N_17553,N_17111,N_17492);
nor U17554 (N_17554,N_16894,N_17397);
nor U17555 (N_17555,N_16734,N_16869);
or U17556 (N_17556,N_17197,N_17012);
nand U17557 (N_17557,N_16741,N_16303);
or U17558 (N_17558,N_16664,N_16317);
xnor U17559 (N_17559,N_17297,N_17189);
xor U17560 (N_17560,N_17472,N_16985);
and U17561 (N_17561,N_16324,N_16355);
and U17562 (N_17562,N_16424,N_16483);
or U17563 (N_17563,N_17114,N_17254);
or U17564 (N_17564,N_16898,N_16794);
and U17565 (N_17565,N_16839,N_16470);
xor U17566 (N_17566,N_16583,N_16361);
and U17567 (N_17567,N_16457,N_16763);
or U17568 (N_17568,N_16944,N_16529);
xnor U17569 (N_17569,N_16399,N_17173);
nand U17570 (N_17570,N_16263,N_16540);
nand U17571 (N_17571,N_16673,N_16864);
and U17572 (N_17572,N_16708,N_16739);
or U17573 (N_17573,N_17274,N_17270);
nand U17574 (N_17574,N_17037,N_16447);
or U17575 (N_17575,N_16517,N_16965);
nand U17576 (N_17576,N_16537,N_16930);
or U17577 (N_17577,N_17065,N_16385);
or U17578 (N_17578,N_16306,N_16595);
nand U17579 (N_17579,N_17185,N_16376);
or U17580 (N_17580,N_16639,N_16799);
nand U17581 (N_17581,N_17383,N_17043);
and U17582 (N_17582,N_17127,N_16863);
nand U17583 (N_17583,N_16653,N_17462);
nand U17584 (N_17584,N_17426,N_16756);
nor U17585 (N_17585,N_17425,N_16534);
xnor U17586 (N_17586,N_16815,N_16738);
and U17587 (N_17587,N_17424,N_16341);
nand U17588 (N_17588,N_16454,N_17223);
nand U17589 (N_17589,N_17366,N_16736);
nor U17590 (N_17590,N_16408,N_16448);
xor U17591 (N_17591,N_17156,N_16755);
or U17592 (N_17592,N_16647,N_16453);
xnor U17593 (N_17593,N_16526,N_17016);
nor U17594 (N_17594,N_16492,N_16841);
or U17595 (N_17595,N_16512,N_17115);
nand U17596 (N_17596,N_16939,N_17308);
nand U17597 (N_17597,N_16749,N_16267);
and U17598 (N_17598,N_16587,N_16891);
xnor U17599 (N_17599,N_16668,N_17258);
nand U17600 (N_17600,N_16747,N_16808);
nor U17601 (N_17601,N_16852,N_16436);
xor U17602 (N_17602,N_16807,N_17186);
nand U17603 (N_17603,N_16695,N_16710);
nand U17604 (N_17604,N_16409,N_17335);
nand U17605 (N_17605,N_17046,N_16919);
or U17606 (N_17606,N_17303,N_16275);
and U17607 (N_17607,N_16764,N_17495);
xor U17608 (N_17608,N_16471,N_16505);
or U17609 (N_17609,N_16569,N_16373);
nand U17610 (N_17610,N_16958,N_16271);
or U17611 (N_17611,N_16828,N_17278);
and U17612 (N_17612,N_16604,N_16746);
nand U17613 (N_17613,N_17483,N_16623);
and U17614 (N_17614,N_16591,N_16918);
xor U17615 (N_17615,N_16825,N_16430);
nor U17616 (N_17616,N_16760,N_16254);
nor U17617 (N_17617,N_16261,N_16397);
and U17618 (N_17618,N_16860,N_16873);
xor U17619 (N_17619,N_16539,N_16284);
and U17620 (N_17620,N_16744,N_17271);
nor U17621 (N_17621,N_16875,N_16380);
nor U17622 (N_17622,N_16510,N_16902);
nand U17623 (N_17623,N_17034,N_17152);
xor U17624 (N_17624,N_16784,N_16922);
nand U17625 (N_17625,N_17091,N_17247);
and U17626 (N_17626,N_17145,N_16844);
nand U17627 (N_17627,N_16559,N_16882);
and U17628 (N_17628,N_16354,N_16750);
or U17629 (N_17629,N_16536,N_16689);
xnor U17630 (N_17630,N_16848,N_17092);
or U17631 (N_17631,N_16753,N_16449);
nand U17632 (N_17632,N_16726,N_16804);
nor U17633 (N_17633,N_16694,N_16851);
nor U17634 (N_17634,N_16472,N_16294);
xor U17635 (N_17635,N_16967,N_17285);
xnor U17636 (N_17636,N_16822,N_17118);
xor U17637 (N_17637,N_16359,N_17105);
xnor U17638 (N_17638,N_17360,N_17432);
xor U17639 (N_17639,N_17228,N_16590);
or U17640 (N_17640,N_17361,N_17178);
xnor U17641 (N_17641,N_17327,N_17216);
nand U17642 (N_17642,N_17172,N_16679);
nand U17643 (N_17643,N_17195,N_16377);
xnor U17644 (N_17644,N_16801,N_17454);
nor U17645 (N_17645,N_17304,N_16811);
nor U17646 (N_17646,N_16482,N_17337);
nand U17647 (N_17647,N_16363,N_17421);
nor U17648 (N_17648,N_16511,N_16723);
nand U17649 (N_17649,N_16840,N_17450);
nand U17650 (N_17650,N_17460,N_17305);
nand U17651 (N_17651,N_16633,N_16730);
nand U17652 (N_17652,N_16250,N_17193);
or U17653 (N_17653,N_17094,N_16733);
and U17654 (N_17654,N_16277,N_16522);
or U17655 (N_17655,N_16999,N_16437);
nand U17656 (N_17656,N_17164,N_17206);
or U17657 (N_17657,N_17182,N_16963);
xnor U17658 (N_17658,N_17191,N_17201);
nor U17659 (N_17659,N_16976,N_16909);
or U17660 (N_17660,N_16713,N_17237);
xnor U17661 (N_17661,N_17469,N_16280);
xor U17662 (N_17662,N_17159,N_16353);
nor U17663 (N_17663,N_16415,N_16315);
nor U17664 (N_17664,N_16964,N_17255);
nor U17665 (N_17665,N_17131,N_17373);
nor U17666 (N_17666,N_17235,N_16698);
or U17667 (N_17667,N_16665,N_16299);
nand U17668 (N_17668,N_16564,N_16304);
nand U17669 (N_17669,N_16578,N_16375);
or U17670 (N_17670,N_17090,N_17180);
or U17671 (N_17671,N_17018,N_16611);
and U17672 (N_17672,N_16836,N_16458);
nand U17673 (N_17673,N_16319,N_16596);
or U17674 (N_17674,N_16971,N_16389);
xor U17675 (N_17675,N_16504,N_17457);
nor U17676 (N_17676,N_17309,N_16684);
or U17677 (N_17677,N_17060,N_17054);
nand U17678 (N_17678,N_16908,N_16778);
xnor U17679 (N_17679,N_16972,N_16987);
or U17680 (N_17680,N_17041,N_16441);
nand U17681 (N_17681,N_16834,N_17396);
xor U17682 (N_17682,N_17244,N_16521);
nor U17683 (N_17683,N_16285,N_16910);
nor U17684 (N_17684,N_16352,N_17374);
nor U17685 (N_17685,N_17434,N_17048);
xnor U17686 (N_17686,N_16843,N_16328);
nand U17687 (N_17687,N_16316,N_16549);
and U17688 (N_17688,N_17153,N_17315);
and U17689 (N_17689,N_16682,N_17443);
and U17690 (N_17690,N_17346,N_17250);
and U17691 (N_17691,N_16988,N_17411);
or U17692 (N_17692,N_17230,N_17110);
nor U17693 (N_17693,N_17467,N_16501);
xnor U17694 (N_17694,N_16631,N_17362);
nor U17695 (N_17695,N_16671,N_17087);
or U17696 (N_17696,N_16646,N_17160);
and U17697 (N_17697,N_17276,N_17493);
nor U17698 (N_17698,N_16374,N_16452);
xor U17699 (N_17699,N_16553,N_17345);
nor U17700 (N_17700,N_17350,N_17137);
nand U17701 (N_17701,N_17453,N_16725);
nor U17702 (N_17702,N_17420,N_17112);
xnor U17703 (N_17703,N_16870,N_16266);
or U17704 (N_17704,N_16669,N_16892);
nand U17705 (N_17705,N_16773,N_16662);
or U17706 (N_17706,N_17298,N_16781);
xnor U17707 (N_17707,N_17010,N_17154);
nand U17708 (N_17708,N_16260,N_17340);
xor U17709 (N_17709,N_17188,N_17219);
xnor U17710 (N_17710,N_17319,N_17168);
or U17711 (N_17711,N_16314,N_16562);
nand U17712 (N_17712,N_17359,N_17093);
or U17713 (N_17713,N_16928,N_17040);
nand U17714 (N_17714,N_16566,N_16524);
nand U17715 (N_17715,N_17192,N_16974);
nand U17716 (N_17716,N_17199,N_16348);
nand U17717 (N_17717,N_16975,N_16509);
xnor U17718 (N_17718,N_16838,N_16890);
nand U17719 (N_17719,N_16495,N_17183);
nor U17720 (N_17720,N_16678,N_17229);
or U17721 (N_17721,N_16500,N_16340);
nand U17722 (N_17722,N_17130,N_16265);
nor U17723 (N_17723,N_16913,N_16996);
or U17724 (N_17724,N_16312,N_17463);
nor U17725 (N_17725,N_17213,N_17476);
and U17726 (N_17726,N_16427,N_16480);
xnor U17727 (N_17727,N_17084,N_16464);
or U17728 (N_17728,N_16620,N_17408);
or U17729 (N_17729,N_16745,N_17405);
or U17730 (N_17730,N_17086,N_17203);
or U17731 (N_17731,N_17273,N_17498);
or U17732 (N_17732,N_16858,N_17353);
nor U17733 (N_17733,N_16608,N_17011);
nand U17734 (N_17734,N_16641,N_17342);
nor U17735 (N_17735,N_16800,N_17272);
xnor U17736 (N_17736,N_16290,N_17068);
nand U17737 (N_17737,N_17140,N_17101);
or U17738 (N_17738,N_16961,N_17014);
xor U17739 (N_17739,N_16962,N_16412);
xor U17740 (N_17740,N_17132,N_16704);
and U17741 (N_17741,N_16816,N_17384);
and U17742 (N_17742,N_17354,N_17021);
or U17743 (N_17743,N_17440,N_17435);
and U17744 (N_17744,N_16551,N_17088);
nand U17745 (N_17745,N_16903,N_16597);
nor U17746 (N_17746,N_16752,N_17263);
nor U17747 (N_17747,N_16817,N_16461);
xnor U17748 (N_17748,N_17045,N_16287);
xor U17749 (N_17749,N_17194,N_17332);
or U17750 (N_17750,N_16833,N_17369);
or U17751 (N_17751,N_17447,N_16398);
or U17752 (N_17752,N_16893,N_17039);
xnor U17753 (N_17753,N_16945,N_16735);
nor U17754 (N_17754,N_16379,N_16829);
nand U17755 (N_17755,N_17422,N_16270);
nand U17756 (N_17756,N_17119,N_16394);
nand U17757 (N_17757,N_16530,N_17394);
and U17758 (N_17758,N_17070,N_16899);
xor U17759 (N_17759,N_17089,N_17458);
or U17760 (N_17760,N_16329,N_16292);
and U17761 (N_17761,N_17055,N_16824);
nor U17762 (N_17762,N_16649,N_16780);
or U17763 (N_17763,N_16494,N_16384);
or U17764 (N_17764,N_16527,N_16383);
and U17765 (N_17765,N_17109,N_16788);
nand U17766 (N_17766,N_16440,N_17076);
nor U17767 (N_17767,N_16616,N_16983);
xnor U17768 (N_17768,N_16518,N_16989);
nor U17769 (N_17769,N_16905,N_17488);
xnor U17770 (N_17770,N_17387,N_17224);
and U17771 (N_17771,N_16949,N_17120);
xnor U17772 (N_17772,N_16856,N_16697);
and U17773 (N_17773,N_17085,N_16463);
xor U17774 (N_17774,N_17403,N_17310);
nand U17775 (N_17775,N_16487,N_16660);
nand U17776 (N_17776,N_16826,N_16484);
xnor U17777 (N_17777,N_16772,N_17307);
xnor U17778 (N_17778,N_16503,N_16282);
nand U17779 (N_17779,N_17311,N_16619);
nor U17780 (N_17780,N_16980,N_16872);
xor U17781 (N_17781,N_17414,N_17200);
xnor U17782 (N_17782,N_16720,N_16567);
or U17783 (N_17783,N_16941,N_17058);
nor U17784 (N_17784,N_16878,N_16481);
and U17785 (N_17785,N_16585,N_17441);
xnor U17786 (N_17786,N_16468,N_17428);
xnor U17787 (N_17787,N_16599,N_16802);
nor U17788 (N_17788,N_16823,N_16652);
or U17789 (N_17789,N_17019,N_16624);
nand U17790 (N_17790,N_16281,N_16871);
xnor U17791 (N_17791,N_16347,N_17126);
and U17792 (N_17792,N_17347,N_16451);
xnor U17793 (N_17793,N_16450,N_17146);
nor U17794 (N_17794,N_17487,N_17442);
nand U17795 (N_17795,N_17069,N_17162);
and U17796 (N_17796,N_16574,N_17143);
nand U17797 (N_17797,N_16791,N_17204);
nor U17798 (N_17798,N_16785,N_16712);
nor U17799 (N_17799,N_17253,N_17128);
or U17800 (N_17800,N_17134,N_16819);
nor U17801 (N_17801,N_17375,N_17209);
and U17802 (N_17802,N_16812,N_16637);
or U17803 (N_17803,N_16895,N_16508);
nand U17804 (N_17804,N_17439,N_16543);
nand U17805 (N_17805,N_16400,N_16683);
or U17806 (N_17806,N_17368,N_16264);
or U17807 (N_17807,N_16663,N_17380);
nor U17808 (N_17808,N_16382,N_16392);
nor U17809 (N_17809,N_16278,N_16262);
or U17810 (N_17810,N_16924,N_16648);
or U17811 (N_17811,N_16491,N_16914);
or U17812 (N_17812,N_16429,N_16425);
or U17813 (N_17813,N_17251,N_17177);
nand U17814 (N_17814,N_17163,N_17035);
and U17815 (N_17815,N_16661,N_17313);
or U17816 (N_17816,N_17407,N_17328);
nor U17817 (N_17817,N_16592,N_17221);
or U17818 (N_17818,N_16628,N_17349);
nand U17819 (N_17819,N_17176,N_16970);
and U17820 (N_17820,N_16777,N_16334);
or U17821 (N_17821,N_16686,N_16442);
nor U17822 (N_17822,N_17316,N_17232);
xor U17823 (N_17823,N_17004,N_17437);
nor U17824 (N_17824,N_16655,N_16900);
and U17825 (N_17825,N_17208,N_17217);
or U17826 (N_17826,N_16925,N_16904);
nor U17827 (N_17827,N_16469,N_17331);
and U17828 (N_17828,N_16283,N_17212);
nor U17829 (N_17829,N_16327,N_16643);
xor U17830 (N_17830,N_16774,N_16541);
or U17831 (N_17831,N_17095,N_16372);
nor U17832 (N_17832,N_17124,N_17283);
or U17833 (N_17833,N_16727,N_16765);
nand U17834 (N_17834,N_16982,N_17484);
xnor U17835 (N_17835,N_16404,N_16326);
or U17836 (N_17836,N_16680,N_16538);
xnor U17837 (N_17837,N_16293,N_16546);
or U17838 (N_17838,N_16343,N_16577);
nor U17839 (N_17839,N_16605,N_16771);
nand U17840 (N_17840,N_16897,N_16434);
or U17841 (N_17841,N_16322,N_17282);
xnor U17842 (N_17842,N_16701,N_16336);
nor U17843 (N_17843,N_16297,N_17220);
nand U17844 (N_17844,N_16929,N_16344);
and U17845 (N_17845,N_17468,N_16896);
and U17846 (N_17846,N_16759,N_16289);
xor U17847 (N_17847,N_16709,N_16992);
and U17848 (N_17848,N_16857,N_17030);
or U17849 (N_17849,N_17378,N_16386);
nor U17850 (N_17850,N_17103,N_16528);
and U17851 (N_17851,N_17256,N_16769);
nand U17852 (N_17852,N_16955,N_17480);
nand U17853 (N_17853,N_16474,N_17169);
or U17854 (N_17854,N_16570,N_16692);
nand U17855 (N_17855,N_16618,N_16940);
or U17856 (N_17856,N_17281,N_17171);
or U17857 (N_17857,N_17401,N_16706);
nand U17858 (N_17858,N_16716,N_16699);
xnor U17859 (N_17859,N_16688,N_17466);
xnor U17860 (N_17860,N_17478,N_16877);
and U17861 (N_17861,N_16795,N_17324);
nor U17862 (N_17862,N_17207,N_16920);
or U17863 (N_17863,N_17343,N_17099);
nor U17864 (N_17864,N_16531,N_16364);
and U17865 (N_17865,N_17245,N_16984);
xnor U17866 (N_17866,N_16423,N_17431);
nand U17867 (N_17867,N_17363,N_17049);
nor U17868 (N_17868,N_16593,N_16335);
or U17869 (N_17869,N_16446,N_16614);
nand U17870 (N_17870,N_17497,N_16651);
nor U17871 (N_17871,N_16790,N_16488);
nor U17872 (N_17872,N_17338,N_17277);
nand U17873 (N_17873,N_16556,N_16431);
and U17874 (N_17874,N_17288,N_16957);
nand U17875 (N_17875,N_16995,N_17317);
nor U17876 (N_17876,N_17264,N_16915);
and U17877 (N_17877,N_17135,N_17370);
and U17878 (N_17878,N_16743,N_17211);
and U17879 (N_17879,N_17202,N_17218);
nand U17880 (N_17880,N_17031,N_17133);
or U17881 (N_17881,N_17367,N_16693);
nand U17882 (N_17882,N_17364,N_16981);
or U17883 (N_17883,N_16979,N_17433);
xnor U17884 (N_17884,N_17071,N_17287);
or U17885 (N_17885,N_17008,N_17234);
or U17886 (N_17886,N_16279,N_16990);
and U17887 (N_17887,N_16853,N_16558);
nand U17888 (N_17888,N_16339,N_17398);
nor U17889 (N_17889,N_17302,N_16560);
and U17890 (N_17890,N_17238,N_16626);
and U17891 (N_17891,N_16571,N_16443);
nor U17892 (N_17892,N_17158,N_17265);
and U17893 (N_17893,N_17392,N_16632);
and U17894 (N_17894,N_17477,N_16584);
or U17895 (N_17895,N_17320,N_17295);
xor U17896 (N_17896,N_17490,N_16438);
or U17897 (N_17897,N_17410,N_16625);
nand U17898 (N_17898,N_16416,N_17322);
and U17899 (N_17899,N_17081,N_16318);
or U17900 (N_17900,N_17107,N_17241);
or U17901 (N_17901,N_16308,N_16792);
nand U17902 (N_17902,N_17292,N_16612);
nor U17903 (N_17903,N_16479,N_16805);
or U17904 (N_17904,N_17009,N_16883);
nand U17905 (N_17905,N_16428,N_17329);
nand U17906 (N_17906,N_16814,N_16542);
or U17907 (N_17907,N_16674,N_16572);
xnor U17908 (N_17908,N_17157,N_17226);
nor U17909 (N_17909,N_16506,N_17314);
and U17910 (N_17910,N_17142,N_16740);
nand U17911 (N_17911,N_16789,N_16555);
or U17912 (N_17912,N_16867,N_16742);
or U17913 (N_17913,N_16952,N_16787);
xnor U17914 (N_17914,N_17017,N_16998);
xnor U17915 (N_17915,N_17358,N_16821);
xnor U17916 (N_17916,N_16960,N_17020);
or U17917 (N_17917,N_16330,N_16420);
nand U17918 (N_17918,N_16737,N_16855);
xor U17919 (N_17919,N_17464,N_16849);
nor U17920 (N_17920,N_16953,N_16251);
and U17921 (N_17921,N_17033,N_16813);
nor U17922 (N_17922,N_17400,N_16381);
nor U17923 (N_17923,N_17321,N_16467);
nor U17924 (N_17924,N_16378,N_16703);
xor U17925 (N_17925,N_16884,N_16622);
nand U17926 (N_17926,N_16337,N_17080);
nand U17927 (N_17927,N_17381,N_16598);
or U17928 (N_17928,N_16466,N_17402);
nand U17929 (N_17929,N_16831,N_16837);
nor U17930 (N_17930,N_16642,N_16321);
or U17931 (N_17931,N_16493,N_17236);
or U17932 (N_17932,N_16601,N_16406);
and U17933 (N_17933,N_17187,N_16258);
xor U17934 (N_17934,N_16758,N_16565);
or U17935 (N_17935,N_17390,N_17356);
xor U17936 (N_17936,N_16422,N_17141);
nand U17937 (N_17937,N_16342,N_17072);
nand U17938 (N_17938,N_17013,N_17150);
xor U17939 (N_17939,N_17106,N_16309);
and U17940 (N_17940,N_16927,N_16388);
nand U17941 (N_17941,N_16700,N_17240);
and U17942 (N_17942,N_16255,N_16654);
xor U17943 (N_17943,N_17057,N_17215);
nand U17944 (N_17944,N_17100,N_17412);
nor U17945 (N_17945,N_17395,N_16702);
nor U17946 (N_17946,N_17481,N_17348);
xnor U17947 (N_17947,N_17293,N_16445);
or U17948 (N_17948,N_16356,N_17248);
nand U17949 (N_17949,N_16581,N_16345);
nand U17950 (N_17950,N_16946,N_16806);
xnor U17951 (N_17951,N_16455,N_16866);
xor U17952 (N_17952,N_16253,N_16496);
xor U17953 (N_17953,N_16489,N_17198);
nor U17954 (N_17954,N_17243,N_16714);
xnor U17955 (N_17955,N_17083,N_16396);
nor U17956 (N_17956,N_16486,N_16615);
xnor U17957 (N_17957,N_16956,N_17098);
nor U17958 (N_17958,N_16847,N_17385);
nand U17959 (N_17959,N_17022,N_17073);
xnor U17960 (N_17960,N_17279,N_16690);
xor U17961 (N_17961,N_17117,N_16576);
nor U17962 (N_17962,N_16405,N_16459);
or U17963 (N_17963,N_16532,N_17249);
nand U17964 (N_17964,N_17056,N_16715);
or U17965 (N_17965,N_17275,N_17376);
nor U17966 (N_17966,N_16786,N_16432);
nor U17967 (N_17967,N_17280,N_16621);
xnor U17968 (N_17968,N_16320,N_17352);
and U17969 (N_17969,N_17474,N_16366);
xor U17970 (N_17970,N_17419,N_16809);
xnor U17971 (N_17971,N_17290,N_17333);
or U17972 (N_17972,N_16594,N_16757);
and U17973 (N_17973,N_16588,N_16391);
or U17974 (N_17974,N_17015,N_16954);
xnor U17975 (N_17975,N_16362,N_16276);
or U17976 (N_17976,N_16640,N_16535);
nand U17977 (N_17977,N_16798,N_16515);
xnor U17978 (N_17978,N_17473,N_17042);
nor U17979 (N_17979,N_16272,N_16658);
or U17980 (N_17980,N_17166,N_17113);
nor U17981 (N_17981,N_16365,N_16368);
and U17982 (N_17982,N_17444,N_17082);
or U17983 (N_17983,N_17365,N_17174);
or U17984 (N_17984,N_16552,N_16676);
xnor U17985 (N_17985,N_16722,N_17455);
nand U17986 (N_17986,N_17318,N_17053);
xor U17987 (N_17987,N_17061,N_17438);
nand U17988 (N_17988,N_17486,N_17482);
nand U17989 (N_17989,N_16301,N_17246);
nand U17990 (N_17990,N_16724,N_17379);
and U17991 (N_17991,N_16473,N_16523);
xor U17992 (N_17992,N_17485,N_16707);
nand U17993 (N_17993,N_16268,N_17144);
and U17994 (N_17994,N_16456,N_16401);
nand U17995 (N_17995,N_16644,N_16256);
or U17996 (N_17996,N_17388,N_17336);
nand U17997 (N_17997,N_17155,N_16943);
nor U17998 (N_17998,N_16402,N_16617);
and U17999 (N_17999,N_16842,N_16311);
nand U18000 (N_18000,N_16497,N_17210);
and U18001 (N_18001,N_17413,N_17097);
or U18002 (N_18002,N_16331,N_17423);
nand U18003 (N_18003,N_17417,N_17139);
or U18004 (N_18004,N_17001,N_16414);
and U18005 (N_18005,N_16775,N_17179);
nand U18006 (N_18006,N_16986,N_16978);
xnor U18007 (N_18007,N_17406,N_16548);
or U18008 (N_18008,N_17002,N_17184);
and U18009 (N_18009,N_16444,N_16721);
xor U18010 (N_18010,N_16610,N_16462);
and U18011 (N_18011,N_16886,N_16332);
xor U18012 (N_18012,N_16520,N_16951);
nand U18013 (N_18013,N_16797,N_16300);
or U18014 (N_18014,N_17494,N_17299);
and U18015 (N_18015,N_17108,N_16666);
nor U18016 (N_18016,N_16731,N_16959);
and U18017 (N_18017,N_17051,N_16513);
and U18018 (N_18018,N_17259,N_16257);
or U18019 (N_18019,N_17386,N_16887);
and U18020 (N_18020,N_17371,N_17451);
and U18021 (N_18021,N_17029,N_16936);
xor U18022 (N_18022,N_17050,N_16426);
or U18023 (N_18023,N_17038,N_17471);
nand U18024 (N_18024,N_16561,N_16994);
and U18025 (N_18025,N_16563,N_16288);
xnor U18026 (N_18026,N_16776,N_16732);
nand U18027 (N_18027,N_17445,N_16645);
nor U18028 (N_18028,N_16387,N_17165);
xor U18029 (N_18029,N_16696,N_16476);
nand U18030 (N_18030,N_16931,N_16947);
xor U18031 (N_18031,N_16490,N_16307);
nand U18032 (N_18032,N_16296,N_16573);
nor U18033 (N_18033,N_17077,N_17006);
and U18034 (N_18034,N_17023,N_17147);
or U18035 (N_18035,N_16291,N_17461);
or U18036 (N_18036,N_17404,N_16435);
nor U18037 (N_18037,N_16390,N_17262);
or U18038 (N_18038,N_16360,N_17323);
nor U18039 (N_18039,N_16845,N_16719);
or U18040 (N_18040,N_17067,N_16783);
and U18041 (N_18041,N_17418,N_17149);
or U18042 (N_18042,N_17284,N_17372);
xor U18043 (N_18043,N_16948,N_16525);
or U18044 (N_18044,N_16393,N_16675);
nand U18045 (N_18045,N_16968,N_16793);
xor U18046 (N_18046,N_16274,N_16677);
and U18047 (N_18047,N_16533,N_16782);
and U18048 (N_18048,N_16302,N_16346);
nand U18049 (N_18049,N_16754,N_16586);
and U18050 (N_18050,N_17312,N_16862);
xnor U18051 (N_18051,N_16761,N_17066);
xor U18052 (N_18052,N_17291,N_16748);
and U18053 (N_18053,N_17325,N_17102);
nand U18054 (N_18054,N_17122,N_17351);
xor U18055 (N_18055,N_16916,N_16544);
or U18056 (N_18056,N_16681,N_16499);
or U18057 (N_18057,N_16603,N_17148);
xor U18058 (N_18058,N_16885,N_16305);
nand U18059 (N_18059,N_16717,N_16507);
nand U18060 (N_18060,N_16323,N_17151);
xor U18061 (N_18061,N_16630,N_16629);
or U18062 (N_18062,N_16803,N_16259);
xnor U18063 (N_18063,N_16460,N_16950);
or U18064 (N_18064,N_16912,N_16286);
or U18065 (N_18065,N_16371,N_16818);
nor U18066 (N_18066,N_16820,N_16465);
nand U18067 (N_18067,N_17357,N_16751);
nand U18068 (N_18068,N_17415,N_16421);
and U18069 (N_18069,N_16859,N_16370);
or U18070 (N_18070,N_17167,N_17239);
and U18071 (N_18071,N_16969,N_17175);
nand U18072 (N_18072,N_17028,N_16514);
and U18073 (N_18073,N_16602,N_17063);
xnor U18074 (N_18074,N_16977,N_17268);
or U18075 (N_18075,N_17074,N_16417);
and U18076 (N_18076,N_16881,N_16606);
nand U18077 (N_18077,N_16485,N_17161);
and U18078 (N_18078,N_17326,N_17475);
xnor U18079 (N_18079,N_17456,N_16413);
nand U18080 (N_18080,N_16827,N_16475);
nor U18081 (N_18081,N_17123,N_16993);
nand U18082 (N_18082,N_17269,N_16687);
xor U18083 (N_18083,N_16550,N_16997);
nor U18084 (N_18084,N_16407,N_16580);
nand U18085 (N_18085,N_17296,N_16350);
nand U18086 (N_18086,N_17306,N_17231);
xor U18087 (N_18087,N_16367,N_16575);
nor U18088 (N_18088,N_16516,N_16861);
or U18089 (N_18089,N_16557,N_16498);
xnor U18090 (N_18090,N_17181,N_16762);
or U18091 (N_18091,N_17044,N_16638);
xor U18092 (N_18092,N_17075,N_16635);
or U18093 (N_18093,N_16868,N_16607);
and U18094 (N_18094,N_16554,N_17257);
and U18095 (N_18095,N_16395,N_16433);
nor U18096 (N_18096,N_16766,N_16921);
or U18097 (N_18097,N_17391,N_17125);
and U18098 (N_18098,N_16718,N_16313);
and U18099 (N_18099,N_16519,N_16876);
and U18100 (N_18100,N_17491,N_17377);
and U18101 (N_18101,N_17294,N_16880);
or U18102 (N_18102,N_17430,N_16667);
nand U18103 (N_18103,N_16991,N_17355);
nand U18104 (N_18104,N_16966,N_17032);
and U18105 (N_18105,N_16832,N_16439);
nand U18106 (N_18106,N_16926,N_16502);
or U18107 (N_18107,N_17436,N_16333);
or U18108 (N_18108,N_16874,N_16589);
or U18109 (N_18109,N_17005,N_16911);
and U18110 (N_18110,N_17448,N_16310);
nor U18111 (N_18111,N_17242,N_16938);
and U18112 (N_18112,N_17078,N_16729);
nor U18113 (N_18113,N_16691,N_16545);
or U18114 (N_18114,N_16767,N_17096);
or U18115 (N_18115,N_17300,N_17334);
xor U18116 (N_18116,N_16932,N_16634);
nand U18117 (N_18117,N_17416,N_17267);
xor U18118 (N_18118,N_16657,N_16351);
xor U18119 (N_18119,N_17393,N_16670);
nor U18120 (N_18120,N_17047,N_16906);
or U18121 (N_18121,N_16547,N_16403);
xnor U18122 (N_18122,N_16711,N_17214);
and U18123 (N_18123,N_16579,N_16835);
nor U18124 (N_18124,N_16568,N_16411);
xnor U18125 (N_18125,N_16268,N_17224);
and U18126 (N_18126,N_17014,N_17178);
and U18127 (N_18127,N_17313,N_16317);
nor U18128 (N_18128,N_17381,N_16768);
nor U18129 (N_18129,N_16327,N_16733);
or U18130 (N_18130,N_17150,N_17426);
nor U18131 (N_18131,N_16993,N_16712);
nor U18132 (N_18132,N_16889,N_16434);
nand U18133 (N_18133,N_16405,N_17155);
and U18134 (N_18134,N_17079,N_16641);
and U18135 (N_18135,N_16455,N_17171);
or U18136 (N_18136,N_16531,N_16701);
nand U18137 (N_18137,N_17022,N_16936);
nor U18138 (N_18138,N_16327,N_17021);
or U18139 (N_18139,N_16741,N_17424);
and U18140 (N_18140,N_17042,N_17370);
or U18141 (N_18141,N_16408,N_16636);
nand U18142 (N_18142,N_17361,N_16954);
nand U18143 (N_18143,N_16444,N_16945);
nor U18144 (N_18144,N_17068,N_17005);
or U18145 (N_18145,N_17239,N_16584);
nor U18146 (N_18146,N_17133,N_17471);
nand U18147 (N_18147,N_16250,N_16397);
and U18148 (N_18148,N_17476,N_16888);
and U18149 (N_18149,N_17010,N_16395);
or U18150 (N_18150,N_16671,N_17297);
and U18151 (N_18151,N_17419,N_17185);
or U18152 (N_18152,N_17154,N_16960);
and U18153 (N_18153,N_16399,N_17456);
or U18154 (N_18154,N_16600,N_16418);
and U18155 (N_18155,N_16904,N_16274);
or U18156 (N_18156,N_16486,N_17349);
nor U18157 (N_18157,N_16711,N_17412);
nand U18158 (N_18158,N_16637,N_16734);
nor U18159 (N_18159,N_16768,N_17230);
and U18160 (N_18160,N_16843,N_16805);
nor U18161 (N_18161,N_17327,N_17450);
and U18162 (N_18162,N_16637,N_17158);
or U18163 (N_18163,N_16463,N_17494);
xor U18164 (N_18164,N_17121,N_16787);
nor U18165 (N_18165,N_17217,N_17297);
xor U18166 (N_18166,N_16412,N_16585);
and U18167 (N_18167,N_17083,N_16430);
nand U18168 (N_18168,N_16837,N_17149);
nand U18169 (N_18169,N_17368,N_16904);
and U18170 (N_18170,N_16436,N_16950);
nor U18171 (N_18171,N_16798,N_17096);
and U18172 (N_18172,N_17259,N_16782);
or U18173 (N_18173,N_16796,N_16894);
nor U18174 (N_18174,N_16634,N_17126);
and U18175 (N_18175,N_16798,N_17219);
nor U18176 (N_18176,N_16660,N_16723);
or U18177 (N_18177,N_17382,N_17275);
xnor U18178 (N_18178,N_17036,N_16346);
nor U18179 (N_18179,N_17281,N_17099);
or U18180 (N_18180,N_16810,N_17034);
or U18181 (N_18181,N_16976,N_17150);
nor U18182 (N_18182,N_17489,N_17385);
or U18183 (N_18183,N_17421,N_16725);
xnor U18184 (N_18184,N_16366,N_16386);
and U18185 (N_18185,N_16999,N_16294);
and U18186 (N_18186,N_16448,N_17268);
or U18187 (N_18187,N_16922,N_17251);
and U18188 (N_18188,N_16929,N_16730);
nand U18189 (N_18189,N_16393,N_16284);
xnor U18190 (N_18190,N_16618,N_17060);
nand U18191 (N_18191,N_17006,N_16756);
nor U18192 (N_18192,N_16704,N_16817);
and U18193 (N_18193,N_17224,N_16280);
nand U18194 (N_18194,N_17422,N_17061);
nor U18195 (N_18195,N_16479,N_16624);
nand U18196 (N_18196,N_17441,N_17297);
or U18197 (N_18197,N_17193,N_17306);
nor U18198 (N_18198,N_17092,N_16577);
and U18199 (N_18199,N_16423,N_16440);
and U18200 (N_18200,N_16758,N_17031);
xnor U18201 (N_18201,N_16996,N_16487);
and U18202 (N_18202,N_17057,N_16656);
nand U18203 (N_18203,N_16592,N_17140);
xor U18204 (N_18204,N_16339,N_16740);
nand U18205 (N_18205,N_16717,N_16297);
nand U18206 (N_18206,N_17051,N_16797);
nand U18207 (N_18207,N_16292,N_17386);
xnor U18208 (N_18208,N_17491,N_17080);
nand U18209 (N_18209,N_17028,N_17329);
or U18210 (N_18210,N_16624,N_16883);
nand U18211 (N_18211,N_16359,N_16713);
nor U18212 (N_18212,N_16513,N_17269);
nand U18213 (N_18213,N_17195,N_17050);
nor U18214 (N_18214,N_16932,N_16758);
nand U18215 (N_18215,N_16756,N_16905);
nand U18216 (N_18216,N_16905,N_16664);
and U18217 (N_18217,N_16823,N_16662);
nor U18218 (N_18218,N_16777,N_17361);
nor U18219 (N_18219,N_17063,N_17051);
or U18220 (N_18220,N_17387,N_16982);
nand U18221 (N_18221,N_16450,N_16265);
xor U18222 (N_18222,N_16609,N_17476);
or U18223 (N_18223,N_16688,N_16816);
xnor U18224 (N_18224,N_17351,N_16279);
or U18225 (N_18225,N_17314,N_16956);
nor U18226 (N_18226,N_16737,N_16589);
and U18227 (N_18227,N_17045,N_16496);
nand U18228 (N_18228,N_17156,N_17249);
xor U18229 (N_18229,N_17145,N_16702);
nand U18230 (N_18230,N_17103,N_16373);
xor U18231 (N_18231,N_16591,N_16416);
and U18232 (N_18232,N_17008,N_17196);
and U18233 (N_18233,N_16736,N_16754);
nand U18234 (N_18234,N_17032,N_16800);
nand U18235 (N_18235,N_16691,N_16776);
xor U18236 (N_18236,N_17399,N_17345);
nor U18237 (N_18237,N_16544,N_17007);
and U18238 (N_18238,N_16462,N_17267);
xnor U18239 (N_18239,N_16818,N_16380);
and U18240 (N_18240,N_16682,N_17433);
xnor U18241 (N_18241,N_16348,N_16326);
nand U18242 (N_18242,N_17289,N_16814);
xnor U18243 (N_18243,N_16530,N_16755);
nor U18244 (N_18244,N_16373,N_17035);
nand U18245 (N_18245,N_17221,N_16641);
and U18246 (N_18246,N_16918,N_16442);
xnor U18247 (N_18247,N_16392,N_17277);
or U18248 (N_18248,N_16597,N_16498);
or U18249 (N_18249,N_17280,N_17346);
or U18250 (N_18250,N_17066,N_17449);
and U18251 (N_18251,N_16390,N_17240);
and U18252 (N_18252,N_16783,N_16758);
or U18253 (N_18253,N_17229,N_16537);
or U18254 (N_18254,N_16410,N_17013);
and U18255 (N_18255,N_17011,N_16641);
xor U18256 (N_18256,N_17373,N_17261);
nor U18257 (N_18257,N_16608,N_16745);
xnor U18258 (N_18258,N_16327,N_17341);
or U18259 (N_18259,N_16636,N_16731);
xor U18260 (N_18260,N_16428,N_16313);
nand U18261 (N_18261,N_16407,N_16828);
nand U18262 (N_18262,N_16511,N_17414);
and U18263 (N_18263,N_17039,N_17414);
nand U18264 (N_18264,N_16519,N_16515);
and U18265 (N_18265,N_16250,N_16962);
nand U18266 (N_18266,N_16763,N_16557);
and U18267 (N_18267,N_16950,N_16690);
nand U18268 (N_18268,N_16750,N_16890);
nand U18269 (N_18269,N_16806,N_16831);
or U18270 (N_18270,N_16929,N_16382);
nand U18271 (N_18271,N_16468,N_16803);
and U18272 (N_18272,N_16683,N_16792);
or U18273 (N_18273,N_17020,N_16424);
xnor U18274 (N_18274,N_16573,N_16815);
or U18275 (N_18275,N_17185,N_17467);
nand U18276 (N_18276,N_16314,N_16817);
and U18277 (N_18277,N_16399,N_17300);
nand U18278 (N_18278,N_17076,N_16345);
nor U18279 (N_18279,N_17299,N_16733);
nand U18280 (N_18280,N_16266,N_17186);
and U18281 (N_18281,N_17424,N_17167);
xnor U18282 (N_18282,N_16358,N_16690);
or U18283 (N_18283,N_17076,N_16802);
nand U18284 (N_18284,N_16338,N_17179);
xnor U18285 (N_18285,N_16978,N_16803);
nand U18286 (N_18286,N_16396,N_16642);
or U18287 (N_18287,N_16625,N_16312);
and U18288 (N_18288,N_16361,N_17125);
and U18289 (N_18289,N_16540,N_16361);
and U18290 (N_18290,N_16396,N_17213);
nor U18291 (N_18291,N_16751,N_16945);
xnor U18292 (N_18292,N_16276,N_16522);
and U18293 (N_18293,N_17442,N_17399);
xor U18294 (N_18294,N_16977,N_16793);
nor U18295 (N_18295,N_16318,N_17197);
or U18296 (N_18296,N_16949,N_17254);
or U18297 (N_18297,N_17470,N_16430);
xnor U18298 (N_18298,N_16374,N_17006);
nand U18299 (N_18299,N_17451,N_17152);
and U18300 (N_18300,N_16792,N_16914);
nand U18301 (N_18301,N_16700,N_16777);
nor U18302 (N_18302,N_16707,N_16925);
xor U18303 (N_18303,N_17256,N_16401);
and U18304 (N_18304,N_16672,N_16401);
nor U18305 (N_18305,N_16978,N_16671);
nand U18306 (N_18306,N_16792,N_16662);
xnor U18307 (N_18307,N_17089,N_16485);
or U18308 (N_18308,N_16951,N_17353);
nand U18309 (N_18309,N_16816,N_16373);
or U18310 (N_18310,N_17091,N_17270);
nand U18311 (N_18311,N_16484,N_16864);
nor U18312 (N_18312,N_16264,N_16351);
or U18313 (N_18313,N_17357,N_16987);
and U18314 (N_18314,N_16871,N_16700);
nor U18315 (N_18315,N_17190,N_16314);
xnor U18316 (N_18316,N_17319,N_17203);
nand U18317 (N_18317,N_16481,N_16897);
xnor U18318 (N_18318,N_16650,N_17180);
nor U18319 (N_18319,N_16604,N_16481);
or U18320 (N_18320,N_17086,N_16648);
nor U18321 (N_18321,N_16371,N_17169);
xor U18322 (N_18322,N_17272,N_16903);
or U18323 (N_18323,N_17363,N_17169);
or U18324 (N_18324,N_16312,N_17217);
xor U18325 (N_18325,N_16914,N_17419);
or U18326 (N_18326,N_17219,N_16513);
nor U18327 (N_18327,N_17420,N_17321);
xor U18328 (N_18328,N_16538,N_16745);
xnor U18329 (N_18329,N_16919,N_17324);
xnor U18330 (N_18330,N_17091,N_17424);
nand U18331 (N_18331,N_17091,N_16880);
and U18332 (N_18332,N_16601,N_16271);
nand U18333 (N_18333,N_17141,N_16358);
nand U18334 (N_18334,N_16281,N_17453);
or U18335 (N_18335,N_17313,N_16644);
nand U18336 (N_18336,N_16538,N_17163);
nand U18337 (N_18337,N_17431,N_16415);
nand U18338 (N_18338,N_16507,N_17283);
nor U18339 (N_18339,N_17342,N_17059);
and U18340 (N_18340,N_16469,N_16710);
nor U18341 (N_18341,N_17252,N_17378);
and U18342 (N_18342,N_16911,N_16499);
and U18343 (N_18343,N_16292,N_16429);
xor U18344 (N_18344,N_16774,N_17003);
nand U18345 (N_18345,N_16710,N_16761);
xnor U18346 (N_18346,N_16487,N_17028);
or U18347 (N_18347,N_16514,N_16511);
xor U18348 (N_18348,N_16681,N_17325);
nand U18349 (N_18349,N_16500,N_16635);
nor U18350 (N_18350,N_17439,N_16639);
xor U18351 (N_18351,N_16365,N_17436);
or U18352 (N_18352,N_16503,N_17487);
xor U18353 (N_18353,N_17447,N_16791);
nor U18354 (N_18354,N_17427,N_17221);
nor U18355 (N_18355,N_17030,N_17179);
nor U18356 (N_18356,N_17317,N_16531);
nand U18357 (N_18357,N_16407,N_16803);
nor U18358 (N_18358,N_17469,N_16944);
or U18359 (N_18359,N_16597,N_16661);
nor U18360 (N_18360,N_16997,N_17049);
xor U18361 (N_18361,N_16361,N_16739);
xnor U18362 (N_18362,N_17146,N_16506);
xnor U18363 (N_18363,N_17214,N_17472);
xor U18364 (N_18364,N_16365,N_17070);
xnor U18365 (N_18365,N_16411,N_16540);
xnor U18366 (N_18366,N_16751,N_16720);
xor U18367 (N_18367,N_16662,N_16388);
nor U18368 (N_18368,N_16877,N_16970);
and U18369 (N_18369,N_16253,N_17166);
or U18370 (N_18370,N_17366,N_16819);
or U18371 (N_18371,N_17393,N_16256);
xor U18372 (N_18372,N_16620,N_16501);
xnor U18373 (N_18373,N_16993,N_17466);
xnor U18374 (N_18374,N_16874,N_17305);
nand U18375 (N_18375,N_17031,N_16879);
and U18376 (N_18376,N_16441,N_16398);
and U18377 (N_18377,N_17181,N_16506);
nand U18378 (N_18378,N_17260,N_17284);
or U18379 (N_18379,N_16739,N_17284);
nand U18380 (N_18380,N_16521,N_16891);
xor U18381 (N_18381,N_16386,N_17267);
and U18382 (N_18382,N_16425,N_16948);
nor U18383 (N_18383,N_16559,N_17076);
or U18384 (N_18384,N_16508,N_16281);
and U18385 (N_18385,N_16675,N_17200);
nand U18386 (N_18386,N_17021,N_17437);
nand U18387 (N_18387,N_17234,N_16272);
or U18388 (N_18388,N_16989,N_16556);
xor U18389 (N_18389,N_17193,N_16420);
or U18390 (N_18390,N_16836,N_17045);
nor U18391 (N_18391,N_16619,N_17147);
nand U18392 (N_18392,N_16764,N_16682);
or U18393 (N_18393,N_16801,N_16298);
nor U18394 (N_18394,N_16934,N_17026);
xor U18395 (N_18395,N_16375,N_16521);
nand U18396 (N_18396,N_17251,N_17472);
nor U18397 (N_18397,N_16368,N_16963);
or U18398 (N_18398,N_16950,N_16869);
nand U18399 (N_18399,N_16898,N_17424);
nor U18400 (N_18400,N_16254,N_16506);
and U18401 (N_18401,N_17117,N_16970);
nor U18402 (N_18402,N_17417,N_17389);
or U18403 (N_18403,N_17089,N_16500);
and U18404 (N_18404,N_16563,N_17209);
and U18405 (N_18405,N_16346,N_16541);
nor U18406 (N_18406,N_16724,N_16566);
and U18407 (N_18407,N_16889,N_17403);
or U18408 (N_18408,N_16946,N_16885);
nor U18409 (N_18409,N_16608,N_17262);
nor U18410 (N_18410,N_16468,N_16258);
or U18411 (N_18411,N_16487,N_17182);
nor U18412 (N_18412,N_17319,N_17240);
nand U18413 (N_18413,N_16827,N_16817);
nand U18414 (N_18414,N_16320,N_16271);
or U18415 (N_18415,N_16396,N_17383);
and U18416 (N_18416,N_16778,N_16476);
nand U18417 (N_18417,N_16460,N_17222);
or U18418 (N_18418,N_17445,N_16876);
and U18419 (N_18419,N_17305,N_16252);
or U18420 (N_18420,N_17315,N_17407);
nand U18421 (N_18421,N_16649,N_16254);
nand U18422 (N_18422,N_17047,N_16933);
nor U18423 (N_18423,N_17362,N_16612);
or U18424 (N_18424,N_16380,N_16577);
or U18425 (N_18425,N_16368,N_16977);
and U18426 (N_18426,N_16550,N_17072);
nor U18427 (N_18427,N_16563,N_16749);
xnor U18428 (N_18428,N_16423,N_17055);
and U18429 (N_18429,N_16548,N_16815);
or U18430 (N_18430,N_16743,N_17127);
nand U18431 (N_18431,N_16423,N_17494);
nor U18432 (N_18432,N_17073,N_16633);
or U18433 (N_18433,N_17127,N_17013);
xnor U18434 (N_18434,N_17402,N_16788);
nor U18435 (N_18435,N_16879,N_17385);
and U18436 (N_18436,N_16272,N_16330);
xnor U18437 (N_18437,N_16603,N_16377);
and U18438 (N_18438,N_16470,N_16880);
xor U18439 (N_18439,N_16727,N_16885);
xor U18440 (N_18440,N_17176,N_16620);
and U18441 (N_18441,N_16887,N_16583);
xnor U18442 (N_18442,N_16577,N_17011);
nor U18443 (N_18443,N_16921,N_16375);
nand U18444 (N_18444,N_16402,N_17163);
nor U18445 (N_18445,N_16678,N_16790);
and U18446 (N_18446,N_16339,N_16948);
nor U18447 (N_18447,N_16400,N_17469);
and U18448 (N_18448,N_16295,N_17253);
or U18449 (N_18449,N_16942,N_16451);
nor U18450 (N_18450,N_17256,N_16957);
nor U18451 (N_18451,N_17490,N_17076);
and U18452 (N_18452,N_16542,N_17090);
and U18453 (N_18453,N_16342,N_17479);
and U18454 (N_18454,N_17270,N_16569);
xor U18455 (N_18455,N_16973,N_16546);
xnor U18456 (N_18456,N_16285,N_17306);
or U18457 (N_18457,N_17320,N_16584);
and U18458 (N_18458,N_16713,N_16973);
nand U18459 (N_18459,N_16253,N_16656);
and U18460 (N_18460,N_17038,N_17007);
nand U18461 (N_18461,N_17356,N_16396);
nand U18462 (N_18462,N_16556,N_16625);
nand U18463 (N_18463,N_17064,N_17139);
nand U18464 (N_18464,N_17489,N_17458);
or U18465 (N_18465,N_16704,N_17405);
and U18466 (N_18466,N_16921,N_17004);
xor U18467 (N_18467,N_17202,N_16548);
or U18468 (N_18468,N_16387,N_16575);
nand U18469 (N_18469,N_17399,N_17191);
xor U18470 (N_18470,N_16408,N_17087);
xnor U18471 (N_18471,N_16957,N_17141);
and U18472 (N_18472,N_16984,N_16947);
xor U18473 (N_18473,N_17419,N_16492);
or U18474 (N_18474,N_16491,N_17392);
nand U18475 (N_18475,N_17010,N_17087);
and U18476 (N_18476,N_17255,N_17109);
and U18477 (N_18477,N_17395,N_16587);
and U18478 (N_18478,N_17284,N_16293);
and U18479 (N_18479,N_17079,N_17286);
xor U18480 (N_18480,N_17391,N_16635);
nand U18481 (N_18481,N_17409,N_17434);
nor U18482 (N_18482,N_16868,N_16789);
xnor U18483 (N_18483,N_16379,N_16792);
xor U18484 (N_18484,N_17188,N_16317);
and U18485 (N_18485,N_16787,N_17471);
xor U18486 (N_18486,N_17182,N_16627);
or U18487 (N_18487,N_16561,N_16291);
or U18488 (N_18488,N_16367,N_16395);
nor U18489 (N_18489,N_16392,N_17345);
nand U18490 (N_18490,N_17486,N_16750);
or U18491 (N_18491,N_16567,N_16899);
or U18492 (N_18492,N_17268,N_16653);
nor U18493 (N_18493,N_17010,N_16750);
nor U18494 (N_18494,N_16296,N_17389);
nor U18495 (N_18495,N_17081,N_16992);
nand U18496 (N_18496,N_16353,N_17242);
xor U18497 (N_18497,N_17280,N_17138);
nor U18498 (N_18498,N_17178,N_17078);
nor U18499 (N_18499,N_16886,N_16253);
and U18500 (N_18500,N_17152,N_17032);
nand U18501 (N_18501,N_16984,N_16371);
or U18502 (N_18502,N_16823,N_17180);
nor U18503 (N_18503,N_16879,N_17398);
nor U18504 (N_18504,N_16667,N_17492);
and U18505 (N_18505,N_16687,N_17271);
nor U18506 (N_18506,N_16780,N_16666);
nor U18507 (N_18507,N_17331,N_16521);
nor U18508 (N_18508,N_17296,N_16344);
or U18509 (N_18509,N_17205,N_16553);
nand U18510 (N_18510,N_16412,N_16939);
and U18511 (N_18511,N_17039,N_17417);
nor U18512 (N_18512,N_16403,N_16271);
xor U18513 (N_18513,N_17366,N_17332);
or U18514 (N_18514,N_17239,N_17093);
and U18515 (N_18515,N_16464,N_17154);
and U18516 (N_18516,N_16262,N_16564);
nor U18517 (N_18517,N_16985,N_16758);
nor U18518 (N_18518,N_17476,N_16473);
and U18519 (N_18519,N_17007,N_17197);
nand U18520 (N_18520,N_17141,N_16579);
and U18521 (N_18521,N_16341,N_17183);
nand U18522 (N_18522,N_17104,N_17208);
nand U18523 (N_18523,N_16570,N_17100);
or U18524 (N_18524,N_17377,N_16635);
or U18525 (N_18525,N_16493,N_17123);
nand U18526 (N_18526,N_16983,N_16459);
nor U18527 (N_18527,N_16785,N_17115);
or U18528 (N_18528,N_16280,N_17214);
nand U18529 (N_18529,N_16987,N_17254);
or U18530 (N_18530,N_17136,N_16601);
xor U18531 (N_18531,N_16568,N_16954);
and U18532 (N_18532,N_16999,N_17401);
xnor U18533 (N_18533,N_16850,N_17174);
or U18534 (N_18534,N_16624,N_17104);
nor U18535 (N_18535,N_17271,N_16473);
xor U18536 (N_18536,N_16315,N_16477);
and U18537 (N_18537,N_16903,N_16464);
nand U18538 (N_18538,N_17376,N_16575);
or U18539 (N_18539,N_16411,N_16384);
nor U18540 (N_18540,N_16343,N_16295);
or U18541 (N_18541,N_17338,N_17114);
or U18542 (N_18542,N_16925,N_16874);
nand U18543 (N_18543,N_17351,N_16347);
and U18544 (N_18544,N_17253,N_17300);
nor U18545 (N_18545,N_17356,N_16940);
nand U18546 (N_18546,N_16342,N_16931);
and U18547 (N_18547,N_17358,N_16777);
nand U18548 (N_18548,N_17219,N_16703);
and U18549 (N_18549,N_16604,N_17075);
and U18550 (N_18550,N_16745,N_17106);
nand U18551 (N_18551,N_16819,N_16619);
xor U18552 (N_18552,N_17447,N_16365);
xor U18553 (N_18553,N_17100,N_16540);
or U18554 (N_18554,N_17228,N_16353);
xor U18555 (N_18555,N_17040,N_16839);
or U18556 (N_18556,N_16553,N_16778);
nand U18557 (N_18557,N_16890,N_16279);
or U18558 (N_18558,N_16254,N_17380);
or U18559 (N_18559,N_17482,N_17131);
nor U18560 (N_18560,N_16276,N_16932);
xnor U18561 (N_18561,N_16984,N_17257);
xor U18562 (N_18562,N_16812,N_17378);
or U18563 (N_18563,N_16902,N_17312);
xor U18564 (N_18564,N_16662,N_17419);
and U18565 (N_18565,N_17254,N_16286);
or U18566 (N_18566,N_17495,N_16791);
nor U18567 (N_18567,N_16971,N_17194);
xor U18568 (N_18568,N_16839,N_16671);
nand U18569 (N_18569,N_16983,N_16525);
and U18570 (N_18570,N_16425,N_16606);
or U18571 (N_18571,N_17349,N_16388);
or U18572 (N_18572,N_16576,N_16844);
and U18573 (N_18573,N_17354,N_16607);
xnor U18574 (N_18574,N_16343,N_16809);
or U18575 (N_18575,N_16861,N_16482);
nand U18576 (N_18576,N_17442,N_17130);
or U18577 (N_18577,N_17091,N_17144);
and U18578 (N_18578,N_16987,N_17290);
nor U18579 (N_18579,N_17073,N_17226);
or U18580 (N_18580,N_17133,N_17306);
xnor U18581 (N_18581,N_17010,N_16724);
or U18582 (N_18582,N_16672,N_16977);
xor U18583 (N_18583,N_16337,N_17433);
and U18584 (N_18584,N_16763,N_17446);
xor U18585 (N_18585,N_16881,N_16267);
xnor U18586 (N_18586,N_17380,N_16882);
nor U18587 (N_18587,N_16452,N_16527);
xnor U18588 (N_18588,N_17031,N_16995);
nor U18589 (N_18589,N_16992,N_17187);
nor U18590 (N_18590,N_16441,N_17367);
and U18591 (N_18591,N_17000,N_16589);
nand U18592 (N_18592,N_17446,N_16305);
xor U18593 (N_18593,N_16772,N_17089);
xnor U18594 (N_18594,N_17492,N_17499);
and U18595 (N_18595,N_16652,N_16858);
xor U18596 (N_18596,N_17392,N_17357);
or U18597 (N_18597,N_17403,N_16811);
and U18598 (N_18598,N_16849,N_16688);
nand U18599 (N_18599,N_16754,N_16365);
nor U18600 (N_18600,N_16979,N_16759);
or U18601 (N_18601,N_17216,N_16751);
xnor U18602 (N_18602,N_17447,N_16749);
xor U18603 (N_18603,N_17483,N_16866);
and U18604 (N_18604,N_17071,N_17238);
nor U18605 (N_18605,N_16521,N_17472);
xor U18606 (N_18606,N_17025,N_16570);
xnor U18607 (N_18607,N_17441,N_17402);
or U18608 (N_18608,N_17056,N_17226);
and U18609 (N_18609,N_16776,N_17245);
nand U18610 (N_18610,N_16458,N_17463);
nand U18611 (N_18611,N_16469,N_16938);
nand U18612 (N_18612,N_16915,N_16444);
nand U18613 (N_18613,N_16570,N_17431);
nor U18614 (N_18614,N_16443,N_16987);
nor U18615 (N_18615,N_16489,N_17190);
or U18616 (N_18616,N_16465,N_16788);
or U18617 (N_18617,N_16398,N_16834);
xnor U18618 (N_18618,N_16479,N_17272);
and U18619 (N_18619,N_16643,N_17413);
nor U18620 (N_18620,N_16929,N_17259);
nor U18621 (N_18621,N_17019,N_17104);
nand U18622 (N_18622,N_16276,N_16589);
xnor U18623 (N_18623,N_16837,N_17115);
xnor U18624 (N_18624,N_16438,N_16651);
or U18625 (N_18625,N_17210,N_16468);
and U18626 (N_18626,N_17352,N_17043);
nor U18627 (N_18627,N_16738,N_17434);
xor U18628 (N_18628,N_17426,N_16260);
nand U18629 (N_18629,N_17441,N_16661);
and U18630 (N_18630,N_16551,N_16484);
or U18631 (N_18631,N_16638,N_16884);
and U18632 (N_18632,N_16357,N_16812);
nor U18633 (N_18633,N_17304,N_17121);
nor U18634 (N_18634,N_17493,N_16464);
nand U18635 (N_18635,N_16700,N_17461);
nor U18636 (N_18636,N_17382,N_16858);
xnor U18637 (N_18637,N_16511,N_17260);
or U18638 (N_18638,N_16627,N_16793);
nor U18639 (N_18639,N_17108,N_16851);
xor U18640 (N_18640,N_16945,N_16380);
and U18641 (N_18641,N_17261,N_17499);
nor U18642 (N_18642,N_17274,N_16939);
xnor U18643 (N_18643,N_17459,N_17008);
and U18644 (N_18644,N_17347,N_17249);
or U18645 (N_18645,N_17392,N_16786);
xnor U18646 (N_18646,N_16772,N_16663);
and U18647 (N_18647,N_17205,N_16741);
or U18648 (N_18648,N_17015,N_16313);
or U18649 (N_18649,N_17316,N_16277);
nand U18650 (N_18650,N_17302,N_16976);
nor U18651 (N_18651,N_17104,N_17492);
and U18652 (N_18652,N_17177,N_16647);
or U18653 (N_18653,N_16438,N_16816);
nor U18654 (N_18654,N_17461,N_17045);
and U18655 (N_18655,N_17124,N_16720);
nor U18656 (N_18656,N_17473,N_16657);
and U18657 (N_18657,N_17366,N_16988);
and U18658 (N_18658,N_16862,N_17102);
xor U18659 (N_18659,N_16935,N_16610);
or U18660 (N_18660,N_17087,N_16561);
xnor U18661 (N_18661,N_16918,N_16305);
nand U18662 (N_18662,N_17291,N_16505);
or U18663 (N_18663,N_17283,N_17007);
and U18664 (N_18664,N_16942,N_17149);
and U18665 (N_18665,N_16757,N_16915);
and U18666 (N_18666,N_16958,N_17432);
nor U18667 (N_18667,N_16337,N_16654);
and U18668 (N_18668,N_16339,N_16567);
or U18669 (N_18669,N_17286,N_16458);
xnor U18670 (N_18670,N_17486,N_16937);
nand U18671 (N_18671,N_17180,N_16911);
nand U18672 (N_18672,N_16273,N_16530);
or U18673 (N_18673,N_17462,N_16822);
or U18674 (N_18674,N_17324,N_16521);
xor U18675 (N_18675,N_17420,N_16887);
nand U18676 (N_18676,N_17487,N_16890);
xor U18677 (N_18677,N_17300,N_17484);
nor U18678 (N_18678,N_16736,N_16499);
nand U18679 (N_18679,N_16414,N_17441);
nor U18680 (N_18680,N_16817,N_16434);
nand U18681 (N_18681,N_17226,N_17233);
nand U18682 (N_18682,N_17231,N_16356);
xnor U18683 (N_18683,N_17383,N_16585);
nand U18684 (N_18684,N_16557,N_17189);
xor U18685 (N_18685,N_16351,N_17285);
nand U18686 (N_18686,N_17242,N_16263);
or U18687 (N_18687,N_16404,N_17399);
nand U18688 (N_18688,N_17003,N_16878);
nor U18689 (N_18689,N_16878,N_17457);
and U18690 (N_18690,N_17352,N_16649);
nor U18691 (N_18691,N_16616,N_17202);
xor U18692 (N_18692,N_16566,N_17146);
and U18693 (N_18693,N_17306,N_16815);
nand U18694 (N_18694,N_17290,N_17073);
nor U18695 (N_18695,N_16422,N_16513);
or U18696 (N_18696,N_16776,N_17116);
nand U18697 (N_18697,N_17337,N_16953);
nor U18698 (N_18698,N_17117,N_17322);
nand U18699 (N_18699,N_17460,N_16947);
and U18700 (N_18700,N_16679,N_17362);
nand U18701 (N_18701,N_16695,N_17242);
and U18702 (N_18702,N_16359,N_16858);
nand U18703 (N_18703,N_17088,N_17293);
or U18704 (N_18704,N_16649,N_17244);
or U18705 (N_18705,N_16840,N_17415);
xnor U18706 (N_18706,N_17082,N_16655);
nand U18707 (N_18707,N_17460,N_16673);
and U18708 (N_18708,N_16990,N_16710);
and U18709 (N_18709,N_17230,N_16747);
xnor U18710 (N_18710,N_17201,N_16799);
xnor U18711 (N_18711,N_17365,N_16532);
and U18712 (N_18712,N_16895,N_16525);
or U18713 (N_18713,N_17213,N_16651);
and U18714 (N_18714,N_17474,N_16816);
nand U18715 (N_18715,N_16553,N_16870);
or U18716 (N_18716,N_16428,N_16295);
nand U18717 (N_18717,N_16782,N_16829);
xor U18718 (N_18718,N_16495,N_16992);
nand U18719 (N_18719,N_17111,N_16506);
xnor U18720 (N_18720,N_16289,N_17076);
or U18721 (N_18721,N_16823,N_16755);
or U18722 (N_18722,N_16625,N_17011);
nor U18723 (N_18723,N_16676,N_17329);
xor U18724 (N_18724,N_16568,N_17420);
xnor U18725 (N_18725,N_17368,N_16586);
nor U18726 (N_18726,N_16823,N_17338);
or U18727 (N_18727,N_16428,N_16954);
nand U18728 (N_18728,N_17275,N_16714);
nor U18729 (N_18729,N_16730,N_16524);
nor U18730 (N_18730,N_16444,N_16640);
xnor U18731 (N_18731,N_16537,N_16996);
nand U18732 (N_18732,N_16692,N_16803);
or U18733 (N_18733,N_16436,N_17204);
nor U18734 (N_18734,N_16858,N_16857);
nand U18735 (N_18735,N_16520,N_16811);
nand U18736 (N_18736,N_17287,N_17212);
and U18737 (N_18737,N_16392,N_17378);
nand U18738 (N_18738,N_17215,N_17435);
xnor U18739 (N_18739,N_17349,N_17040);
nand U18740 (N_18740,N_17048,N_16391);
xor U18741 (N_18741,N_16909,N_16493);
or U18742 (N_18742,N_16942,N_17084);
nand U18743 (N_18743,N_17019,N_16902);
xnor U18744 (N_18744,N_16293,N_16615);
nor U18745 (N_18745,N_17153,N_17253);
or U18746 (N_18746,N_16562,N_16370);
and U18747 (N_18747,N_17054,N_17118);
nand U18748 (N_18748,N_16559,N_17418);
and U18749 (N_18749,N_17467,N_16640);
nand U18750 (N_18750,N_18098,N_17623);
nor U18751 (N_18751,N_18429,N_18146);
nand U18752 (N_18752,N_17651,N_17565);
nand U18753 (N_18753,N_18400,N_18413);
or U18754 (N_18754,N_18699,N_17551);
or U18755 (N_18755,N_17774,N_17770);
nor U18756 (N_18756,N_17611,N_17967);
nand U18757 (N_18757,N_18077,N_17691);
nand U18758 (N_18758,N_18023,N_17573);
nor U18759 (N_18759,N_18067,N_17723);
xor U18760 (N_18760,N_17510,N_18397);
xnor U18761 (N_18761,N_17643,N_18608);
xor U18762 (N_18762,N_18483,N_17619);
xor U18763 (N_18763,N_17513,N_17872);
and U18764 (N_18764,N_18063,N_18702);
or U18765 (N_18765,N_17583,N_17804);
and U18766 (N_18766,N_17563,N_17602);
xnor U18767 (N_18767,N_17989,N_18124);
nor U18768 (N_18768,N_18671,N_18561);
nand U18769 (N_18769,N_17598,N_17720);
nand U18770 (N_18770,N_17843,N_18485);
xnor U18771 (N_18771,N_18481,N_17839);
and U18772 (N_18772,N_17557,N_17854);
or U18773 (N_18773,N_17820,N_17696);
nor U18774 (N_18774,N_18548,N_17825);
and U18775 (N_18775,N_17517,N_18352);
nand U18776 (N_18776,N_18669,N_17836);
nand U18777 (N_18777,N_18004,N_18234);
xor U18778 (N_18778,N_18290,N_18208);
nand U18779 (N_18779,N_17706,N_17961);
xor U18780 (N_18780,N_18594,N_18450);
nand U18781 (N_18781,N_17960,N_18261);
xnor U18782 (N_18782,N_18334,N_17558);
or U18783 (N_18783,N_17639,N_17986);
nand U18784 (N_18784,N_18595,N_17586);
nand U18785 (N_18785,N_18630,N_17549);
and U18786 (N_18786,N_17742,N_18042);
nor U18787 (N_18787,N_18617,N_18428);
or U18788 (N_18788,N_18218,N_18366);
nand U18789 (N_18789,N_18125,N_18027);
and U18790 (N_18790,N_18011,N_17682);
nor U18791 (N_18791,N_18094,N_18133);
nand U18792 (N_18792,N_18165,N_18618);
nor U18793 (N_18793,N_18256,N_18323);
and U18794 (N_18794,N_18742,N_17846);
xnor U18795 (N_18795,N_18328,N_18647);
xor U18796 (N_18796,N_17615,N_18663);
nor U18797 (N_18797,N_18335,N_17750);
and U18798 (N_18798,N_18733,N_18705);
nand U18799 (N_18799,N_18221,N_18112);
xor U18800 (N_18800,N_18641,N_17731);
and U18801 (N_18801,N_18628,N_17959);
or U18802 (N_18802,N_18097,N_18638);
xnor U18803 (N_18803,N_17727,N_18721);
nand U18804 (N_18804,N_18205,N_18744);
xor U18805 (N_18805,N_18532,N_18372);
nand U18806 (N_18806,N_18521,N_17625);
and U18807 (N_18807,N_18048,N_18391);
and U18808 (N_18808,N_17660,N_18609);
or U18809 (N_18809,N_17859,N_18664);
nor U18810 (N_18810,N_18237,N_18028);
or U18811 (N_18811,N_18231,N_18403);
nand U18812 (N_18812,N_18039,N_18259);
nand U18813 (N_18813,N_18229,N_18667);
or U18814 (N_18814,N_18476,N_17789);
nand U18815 (N_18815,N_18108,N_18126);
nor U18816 (N_18816,N_18121,N_18272);
xor U18817 (N_18817,N_17648,N_17894);
nand U18818 (N_18818,N_17624,N_17605);
nand U18819 (N_18819,N_18387,N_18085);
nor U18820 (N_18820,N_18519,N_18310);
nand U18821 (N_18821,N_18631,N_18072);
or U18822 (N_18822,N_18245,N_17932);
and U18823 (N_18823,N_17988,N_17866);
xnor U18824 (N_18824,N_18244,N_18465);
and U18825 (N_18825,N_18657,N_18251);
and U18826 (N_18826,N_17955,N_17555);
and U18827 (N_18827,N_17926,N_18696);
or U18828 (N_18828,N_17924,N_18566);
nand U18829 (N_18829,N_18402,N_17943);
nand U18830 (N_18830,N_18529,N_18083);
nand U18831 (N_18831,N_17858,N_18713);
nor U18832 (N_18832,N_18613,N_17613);
xor U18833 (N_18833,N_18639,N_17977);
xor U18834 (N_18834,N_18567,N_18061);
or U18835 (N_18835,N_17994,N_18740);
nor U18836 (N_18836,N_18140,N_18430);
xor U18837 (N_18837,N_18507,N_17952);
and U18838 (N_18838,N_17920,N_18535);
nand U18839 (N_18839,N_18314,N_17728);
or U18840 (N_18840,N_17515,N_17975);
xnor U18841 (N_18841,N_17949,N_18190);
and U18842 (N_18842,N_17936,N_17860);
nand U18843 (N_18843,N_18526,N_17685);
or U18844 (N_18844,N_18687,N_18636);
or U18845 (N_18845,N_18344,N_18203);
xor U18846 (N_18846,N_18252,N_17528);
nor U18847 (N_18847,N_18374,N_18348);
nand U18848 (N_18848,N_18555,N_17701);
nor U18849 (N_18849,N_18053,N_18729);
nand U18850 (N_18850,N_17791,N_18032);
nand U18851 (N_18851,N_17522,N_17751);
and U18852 (N_18852,N_17543,N_17892);
nand U18853 (N_18853,N_18349,N_17637);
xnor U18854 (N_18854,N_18068,N_18401);
or U18855 (N_18855,N_17883,N_17628);
or U18856 (N_18856,N_17678,N_17566);
or U18857 (N_18857,N_18116,N_17950);
and U18858 (N_18858,N_17579,N_18444);
nor U18859 (N_18859,N_18632,N_17969);
nor U18860 (N_18860,N_18188,N_18212);
nor U18861 (N_18861,N_18484,N_18474);
or U18862 (N_18862,N_18267,N_18722);
nor U18863 (N_18863,N_18606,N_18065);
nor U18864 (N_18864,N_17787,N_17601);
nand U18865 (N_18865,N_17607,N_18357);
nor U18866 (N_18866,N_18496,N_17785);
nor U18867 (N_18867,N_17689,N_17876);
nand U18868 (N_18868,N_17603,N_18487);
nand U18869 (N_18869,N_17600,N_18747);
nand U18870 (N_18870,N_18029,N_18327);
nor U18871 (N_18871,N_18652,N_17903);
nand U18872 (N_18872,N_18573,N_18451);
nand U18873 (N_18873,N_18017,N_18191);
or U18874 (N_18874,N_18223,N_18354);
and U18875 (N_18875,N_18533,N_18179);
or U18876 (N_18876,N_18051,N_17738);
nor U18877 (N_18877,N_18367,N_17963);
and U18878 (N_18878,N_18497,N_18250);
and U18879 (N_18879,N_18684,N_17564);
nand U18880 (N_18880,N_18719,N_17881);
and U18881 (N_18881,N_17874,N_18625);
and U18882 (N_18882,N_17996,N_17606);
or U18883 (N_18883,N_18688,N_18297);
nor U18884 (N_18884,N_18572,N_17928);
or U18885 (N_18885,N_18422,N_17627);
nor U18886 (N_18886,N_17992,N_18610);
or U18887 (N_18887,N_18731,N_18010);
xor U18888 (N_18888,N_17962,N_17794);
nor U18889 (N_18889,N_18135,N_18270);
nor U18890 (N_18890,N_17533,N_17783);
nand U18891 (N_18891,N_17906,N_18622);
nand U18892 (N_18892,N_18534,N_18393);
nor U18893 (N_18893,N_18074,N_17542);
xor U18894 (N_18894,N_17652,N_18087);
and U18895 (N_18895,N_18166,N_18281);
nor U18896 (N_18896,N_17550,N_17500);
nor U18897 (N_18897,N_17818,N_17585);
nor U18898 (N_18898,N_17524,N_18291);
or U18899 (N_18899,N_17879,N_18308);
xor U18900 (N_18900,N_17835,N_18509);
or U18901 (N_18901,N_18536,N_18425);
and U18902 (N_18902,N_17801,N_17939);
nand U18903 (N_18903,N_17878,N_17805);
nor U18904 (N_18904,N_17740,N_17869);
nor U18905 (N_18905,N_17594,N_18350);
or U18906 (N_18906,N_17703,N_18215);
nor U18907 (N_18907,N_18173,N_17978);
nand U18908 (N_18908,N_18346,N_17645);
xor U18909 (N_18909,N_18274,N_17833);
nor U18910 (N_18910,N_18342,N_18439);
or U18911 (N_18911,N_18480,N_18524);
nand U18912 (N_18912,N_17762,N_18064);
and U18913 (N_18913,N_18523,N_17856);
nor U18914 (N_18914,N_18390,N_18193);
and U18915 (N_18915,N_17875,N_18624);
nand U18916 (N_18916,N_18187,N_17741);
nor U18917 (N_18917,N_18662,N_18182);
and U18918 (N_18918,N_17807,N_18093);
xnor U18919 (N_18919,N_17838,N_18356);
nor U18920 (N_18920,N_17655,N_18046);
and U18921 (N_18921,N_17616,N_17958);
and U18922 (N_18922,N_18681,N_18394);
xnor U18923 (N_18923,N_17849,N_18668);
xor U18924 (N_18924,N_18445,N_17845);
nor U18925 (N_18925,N_17813,N_18576);
and U18926 (N_18926,N_17571,N_18512);
or U18927 (N_18927,N_17744,N_18253);
and U18928 (N_18928,N_17912,N_18745);
nand U18929 (N_18929,N_18463,N_18537);
nor U18930 (N_18930,N_18665,N_18047);
and U18931 (N_18931,N_18726,N_18605);
or U18932 (N_18932,N_18707,N_18260);
nand U18933 (N_18933,N_18544,N_18607);
or U18934 (N_18934,N_17529,N_18635);
and U18935 (N_18935,N_18727,N_18404);
xnor U18936 (N_18936,N_17743,N_18706);
and U18937 (N_18937,N_18007,N_17540);
xnor U18938 (N_18938,N_18238,N_17898);
or U18939 (N_18939,N_17589,N_18492);
nor U18940 (N_18940,N_18220,N_17886);
or U18941 (N_18941,N_17861,N_17811);
and U18942 (N_18942,N_17831,N_18648);
nand U18943 (N_18943,N_17755,N_18192);
nor U18944 (N_18944,N_18282,N_18358);
nand U18945 (N_18945,N_17942,N_18184);
nand U18946 (N_18946,N_17568,N_17654);
nand U18947 (N_18947,N_17999,N_18739);
and U18948 (N_18948,N_17908,N_18575);
nand U18949 (N_18949,N_18510,N_18482);
and U18950 (N_18950,N_18325,N_18286);
and U18951 (N_18951,N_17930,N_18157);
nand U18952 (N_18952,N_18351,N_17972);
and U18953 (N_18953,N_17521,N_18306);
and U18954 (N_18954,N_17681,N_17917);
xor U18955 (N_18955,N_17739,N_18710);
and U18956 (N_18956,N_18141,N_17803);
or U18957 (N_18957,N_18037,N_18131);
and U18958 (N_18958,N_18224,N_17931);
nor U18959 (N_18959,N_17509,N_17629);
or U18960 (N_18960,N_17748,N_17553);
or U18961 (N_18961,N_17633,N_17590);
and U18962 (N_18962,N_18611,N_18194);
nor U18963 (N_18963,N_17690,N_17640);
and U18964 (N_18964,N_17984,N_18672);
nand U18965 (N_18965,N_17631,N_18383);
nand U18966 (N_18966,N_17851,N_18202);
and U18967 (N_18967,N_18491,N_18170);
nor U18968 (N_18968,N_17526,N_17954);
nand U18969 (N_18969,N_17848,N_18649);
xnor U18970 (N_18970,N_18525,N_18033);
xnor U18971 (N_18971,N_18115,N_17788);
nor U18972 (N_18972,N_18619,N_17729);
and U18973 (N_18973,N_18433,N_18441);
nor U18974 (N_18974,N_17890,N_18155);
xnor U18975 (N_18975,N_17576,N_17502);
and U18976 (N_18976,N_17925,N_18339);
nor U18977 (N_18977,N_17552,N_18315);
xor U18978 (N_18978,N_18447,N_18436);
xnor U18979 (N_18979,N_17895,N_17888);
and U18980 (N_18980,N_18373,N_18734);
xnor U18981 (N_18981,N_18409,N_18694);
or U18982 (N_18982,N_18353,N_18650);
or U18983 (N_18983,N_17541,N_18030);
and U18984 (N_18984,N_18278,N_18217);
nand U18985 (N_18985,N_17772,N_17980);
nand U18986 (N_18986,N_18380,N_18511);
nor U18987 (N_18987,N_18152,N_17665);
nor U18988 (N_18988,N_18324,N_18162);
nand U18989 (N_18989,N_18147,N_17519);
and U18990 (N_18990,N_18082,N_17864);
and U18991 (N_18991,N_18232,N_18642);
nor U18992 (N_18992,N_17819,N_18545);
or U18993 (N_18993,N_18045,N_17990);
nor U18994 (N_18994,N_18311,N_18295);
or U18995 (N_18995,N_17938,N_18498);
nand U18996 (N_18996,N_17844,N_17777);
nand U18997 (N_18997,N_18596,N_18364);
nand U18998 (N_18998,N_17656,N_17709);
nand U18999 (N_18999,N_18110,N_17592);
nor U19000 (N_19000,N_18009,N_18612);
or U19001 (N_19001,N_18299,N_17561);
xor U19002 (N_19002,N_18411,N_17698);
nand U19003 (N_19003,N_18118,N_17934);
xor U19004 (N_19004,N_18503,N_17756);
nand U19005 (N_19005,N_17667,N_18076);
xor U19006 (N_19006,N_17810,N_17945);
or U19007 (N_19007,N_18593,N_18105);
xor U19008 (N_19008,N_18159,N_18096);
xnor U19009 (N_19009,N_18103,N_18542);
or U19010 (N_19010,N_18435,N_18120);
nand U19011 (N_19011,N_18541,N_17534);
nand U19012 (N_19012,N_18580,N_18214);
nor U19013 (N_19013,N_18177,N_18031);
nand U19014 (N_19014,N_17686,N_17661);
nor U19015 (N_19015,N_17713,N_17596);
nand U19016 (N_19016,N_18459,N_18002);
nor U19017 (N_19017,N_17578,N_18216);
nand U19018 (N_19018,N_18102,N_17862);
nand U19019 (N_19019,N_18725,N_17976);
or U19020 (N_19020,N_17900,N_18528);
and U19021 (N_19021,N_17918,N_17567);
or U19022 (N_19022,N_18160,N_18717);
nand U19023 (N_19023,N_18081,N_18375);
nor U19024 (N_19024,N_17973,N_18467);
and U19025 (N_19025,N_18691,N_18407);
nand U19026 (N_19026,N_18736,N_18377);
or U19027 (N_19027,N_18686,N_18458);
or U19028 (N_19028,N_18122,N_18005);
and U19029 (N_19029,N_17781,N_18369);
nand U19030 (N_19030,N_18200,N_17636);
or U19031 (N_19031,N_17580,N_17951);
nor U19032 (N_19032,N_18737,N_18185);
or U19033 (N_19033,N_18543,N_18326);
nor U19034 (N_19034,N_17718,N_18262);
and U19035 (N_19035,N_17916,N_18629);
and U19036 (N_19036,N_17786,N_17733);
nand U19037 (N_19037,N_17653,N_18106);
and U19038 (N_19038,N_18499,N_17614);
and U19039 (N_19039,N_18239,N_18038);
and U19040 (N_19040,N_18360,N_17798);
or U19041 (N_19041,N_17897,N_17808);
nand U19042 (N_19042,N_18025,N_18438);
nand U19043 (N_19043,N_18302,N_18461);
or U19044 (N_19044,N_17675,N_18181);
and U19045 (N_19045,N_17736,N_17901);
nand U19046 (N_19046,N_17621,N_18175);
xnor U19047 (N_19047,N_18701,N_17516);
nand U19048 (N_19048,N_18129,N_17767);
nand U19049 (N_19049,N_18058,N_17507);
and U19050 (N_19050,N_18195,N_17981);
and U19051 (N_19051,N_17546,N_17520);
nand U19052 (N_19052,N_18018,N_17688);
nor U19053 (N_19053,N_17705,N_17674);
or U19054 (N_19054,N_18225,N_18582);
or U19055 (N_19055,N_17599,N_18587);
nor U19056 (N_19056,N_17768,N_18440);
nand U19057 (N_19057,N_17581,N_18294);
xor U19058 (N_19058,N_18560,N_17577);
and U19059 (N_19059,N_18044,N_18520);
nor U19060 (N_19060,N_17670,N_18059);
xor U19061 (N_19061,N_17760,N_18257);
or U19062 (N_19062,N_18597,N_18183);
xnor U19063 (N_19063,N_18514,N_18254);
nor U19064 (N_19064,N_18341,N_18099);
nor U19065 (N_19065,N_17997,N_17821);
or U19066 (N_19066,N_18716,N_17799);
xnor U19067 (N_19067,N_17909,N_18207);
and U19068 (N_19068,N_17946,N_18264);
nor U19069 (N_19069,N_18266,N_18735);
nor U19070 (N_19070,N_17717,N_18634);
nand U19071 (N_19071,N_17608,N_17868);
or U19072 (N_19072,N_17933,N_17921);
nor U19073 (N_19073,N_18211,N_18198);
xnor U19074 (N_19074,N_18586,N_17915);
nand U19075 (N_19075,N_17889,N_18204);
xnor U19076 (N_19076,N_17865,N_18199);
nor U19077 (N_19077,N_18084,N_17692);
and U19078 (N_19078,N_17714,N_17712);
nand U19079 (N_19079,N_18055,N_17971);
or U19080 (N_19080,N_17504,N_18718);
nand U19081 (N_19081,N_18453,N_18653);
xor U19082 (N_19082,N_17684,N_17560);
nand U19083 (N_19083,N_18709,N_18599);
or U19084 (N_19084,N_18104,N_17779);
xor U19085 (N_19085,N_18590,N_17642);
nor U19086 (N_19086,N_18079,N_18362);
nor U19087 (N_19087,N_18284,N_18693);
xor U19088 (N_19088,N_17823,N_18329);
and U19089 (N_19089,N_18405,N_18034);
or U19090 (N_19090,N_18139,N_18434);
nor U19091 (N_19091,N_18448,N_18673);
nor U19092 (N_19092,N_18690,N_18574);
or U19093 (N_19093,N_17834,N_18470);
and U19094 (N_19094,N_17970,N_17732);
or U19095 (N_19095,N_17896,N_17940);
nor U19096 (N_19096,N_17947,N_18583);
nand U19097 (N_19097,N_17545,N_18263);
or U19098 (N_19098,N_18488,N_18248);
nor U19099 (N_19099,N_18398,N_17735);
or U19100 (N_19100,N_17699,N_18178);
nor U19101 (N_19101,N_18305,N_18723);
nand U19102 (N_19102,N_17852,N_17979);
nand U19103 (N_19103,N_17855,N_17531);
or U19104 (N_19104,N_17508,N_17626);
or U19105 (N_19105,N_18557,N_18677);
xnor U19106 (N_19106,N_18001,N_18410);
nor U19107 (N_19107,N_17658,N_17944);
and U19108 (N_19108,N_18304,N_17663);
xor U19109 (N_19109,N_18502,N_18714);
or U19110 (N_19110,N_18592,N_18080);
and U19111 (N_19111,N_17523,N_17679);
xor U19112 (N_19112,N_18708,N_17983);
and U19113 (N_19113,N_17870,N_17814);
xnor U19114 (N_19114,N_18119,N_17597);
nor U19115 (N_19115,N_17704,N_18227);
nor U19116 (N_19116,N_17582,N_18388);
and U19117 (N_19117,N_18516,N_18703);
nor U19118 (N_19118,N_17761,N_18288);
xor U19119 (N_19119,N_18347,N_18236);
xor U19120 (N_19120,N_17863,N_17724);
or U19121 (N_19121,N_18381,N_17715);
nor U19122 (N_19122,N_17782,N_18389);
and U19123 (N_19123,N_18728,N_18564);
nand U19124 (N_19124,N_18589,N_18666);
nor U19125 (N_19125,N_18466,N_18505);
and U19126 (N_19126,N_17792,N_18550);
xnor U19127 (N_19127,N_18167,N_17800);
nor U19128 (N_19128,N_18562,N_18395);
nand U19129 (N_19129,N_17711,N_18442);
xnor U19130 (N_19130,N_18475,N_18500);
xnor U19131 (N_19131,N_18382,N_18384);
xnor U19132 (N_19132,N_18554,N_17802);
nor U19133 (N_19133,N_17604,N_18456);
or U19134 (N_19134,N_18412,N_18164);
nor U19135 (N_19135,N_18359,N_18621);
or U19136 (N_19136,N_18602,N_18303);
nor U19137 (N_19137,N_17773,N_17877);
or U19138 (N_19138,N_17671,N_18469);
xnor U19139 (N_19139,N_17588,N_18421);
or U19140 (N_19140,N_18700,N_18276);
xor U19141 (N_19141,N_18538,N_18697);
and U19142 (N_19142,N_18035,N_17857);
nand U19143 (N_19143,N_18163,N_18222);
xnor U19144 (N_19144,N_17525,N_17919);
xnor U19145 (N_19145,N_18585,N_18645);
xor U19146 (N_19146,N_18540,N_17530);
nand U19147 (N_19147,N_18015,N_18614);
nand U19148 (N_19148,N_18454,N_18678);
nand U19149 (N_19149,N_17650,N_18089);
nand U19150 (N_19150,N_17548,N_17638);
or U19151 (N_19151,N_17885,N_18138);
nand U19152 (N_19152,N_17880,N_18660);
and U19153 (N_19153,N_17511,N_18109);
xor U19154 (N_19154,N_17764,N_18633);
nand U19155 (N_19155,N_18340,N_18128);
and U19156 (N_19156,N_18396,N_17935);
and U19157 (N_19157,N_17827,N_18692);
nor U19158 (N_19158,N_18741,N_17669);
nor U19159 (N_19159,N_18591,N_18016);
or U19160 (N_19160,N_18013,N_18659);
and U19161 (N_19161,N_18069,N_18517);
or U19162 (N_19162,N_17815,N_18240);
or U19163 (N_19163,N_18003,N_18655);
nand U19164 (N_19164,N_18026,N_17584);
or U19165 (N_19165,N_17673,N_17687);
xor U19166 (N_19166,N_17754,N_17937);
nand U19167 (N_19167,N_18019,N_17829);
or U19168 (N_19168,N_17795,N_17995);
nand U19169 (N_19169,N_18732,N_17752);
and U19170 (N_19170,N_18501,N_18268);
nand U19171 (N_19171,N_18022,N_18000);
or U19172 (N_19172,N_18432,N_18551);
nand U19173 (N_19173,N_17612,N_17775);
nor U19174 (N_19174,N_18014,N_18313);
nor U19175 (N_19175,N_18418,N_18515);
nor U19176 (N_19176,N_18494,N_18273);
or U19177 (N_19177,N_18457,N_18423);
or U19178 (N_19178,N_18249,N_18312);
nor U19179 (N_19179,N_17780,N_17641);
and U19180 (N_19180,N_18209,N_17753);
and U19181 (N_19181,N_18241,N_18616);
nor U19182 (N_19182,N_18640,N_18424);
xor U19183 (N_19183,N_18309,N_18603);
and U19184 (N_19184,N_18683,N_17902);
nor U19185 (N_19185,N_18743,N_17593);
nor U19186 (N_19186,N_17758,N_18615);
and U19187 (N_19187,N_17929,N_18330);
nor U19188 (N_19188,N_18552,N_18134);
nand U19189 (N_19189,N_18553,N_18531);
nor U19190 (N_19190,N_18588,N_18539);
xor U19191 (N_19191,N_17506,N_18661);
and U19192 (N_19192,N_18365,N_18489);
or U19193 (N_19193,N_17884,N_17887);
nand U19194 (N_19194,N_18078,N_18041);
nor U19195 (N_19195,N_18558,N_18154);
xnor U19196 (N_19196,N_17956,N_17662);
and U19197 (N_19197,N_17595,N_17797);
and U19198 (N_19198,N_18427,N_17556);
nor U19199 (N_19199,N_17559,N_17694);
or U19200 (N_19200,N_17617,N_17657);
xnor U19201 (N_19201,N_17708,N_18008);
or U19202 (N_19202,N_18604,N_18345);
and U19203 (N_19203,N_17609,N_18623);
xnor U19204 (N_19204,N_18452,N_17527);
or U19205 (N_19205,N_18095,N_18449);
xnor U19206 (N_19206,N_18565,N_18527);
nand U19207 (N_19207,N_18292,N_17745);
nor U19208 (N_19208,N_18255,N_17635);
nor U19209 (N_19209,N_18235,N_18689);
nor U19210 (N_19210,N_18654,N_17644);
nor U19211 (N_19211,N_18477,N_18738);
nand U19212 (N_19212,N_17518,N_17749);
xnor U19213 (N_19213,N_18176,N_18143);
nor U19214 (N_19214,N_18598,N_18130);
xor U19215 (N_19215,N_18651,N_18101);
and U19216 (N_19216,N_18336,N_18100);
nand U19217 (N_19217,N_18420,N_17659);
nor U19218 (N_19218,N_17649,N_17850);
xor U19219 (N_19219,N_18571,N_18376);
nand U19220 (N_19220,N_18724,N_17676);
or U19221 (N_19221,N_18414,N_18050);
nand U19222 (N_19222,N_17948,N_18150);
xnor U19223 (N_19223,N_17867,N_18233);
nand U19224 (N_19224,N_17793,N_17702);
and U19225 (N_19225,N_18443,N_17769);
and U19226 (N_19226,N_18518,N_18021);
or U19227 (N_19227,N_18283,N_18333);
xor U19228 (N_19228,N_17725,N_18298);
and U19229 (N_19229,N_17991,N_18137);
nand U19230 (N_19230,N_18601,N_18680);
or U19231 (N_19231,N_18479,N_18361);
and U19232 (N_19232,N_18417,N_17680);
nor U19233 (N_19233,N_18493,N_17710);
or U19234 (N_19234,N_17871,N_18040);
or U19235 (N_19235,N_18711,N_17683);
nor U19236 (N_19236,N_18054,N_17746);
or U19237 (N_19237,N_17817,N_17847);
xor U19238 (N_19238,N_18293,N_18426);
and U19239 (N_19239,N_18584,N_17677);
nor U19240 (N_19240,N_18371,N_18674);
xor U19241 (N_19241,N_17911,N_17893);
nand U19242 (N_19242,N_17904,N_17505);
and U19243 (N_19243,N_18337,N_17905);
nand U19244 (N_19244,N_17809,N_17666);
and U19245 (N_19245,N_18549,N_18071);
nor U19246 (N_19246,N_17974,N_17634);
nand U19247 (N_19247,N_18730,N_18219);
xnor U19248 (N_19248,N_18392,N_18577);
or U19249 (N_19249,N_17841,N_17927);
and U19250 (N_19250,N_18012,N_17832);
xor U19251 (N_19251,N_18464,N_18145);
and U19252 (N_19252,N_18111,N_18563);
nand U19253 (N_19253,N_18406,N_17514);
nor U19254 (N_19254,N_18246,N_18189);
or U19255 (N_19255,N_18092,N_17899);
nand U19256 (N_19256,N_18066,N_17716);
nand U19257 (N_19257,N_18036,N_17574);
and U19258 (N_19258,N_18287,N_17622);
nor U19259 (N_19259,N_17757,N_18114);
and U19260 (N_19260,N_17840,N_18153);
nor U19261 (N_19261,N_18148,N_18473);
nand U19262 (N_19262,N_18468,N_18471);
nand U19263 (N_19263,N_17982,N_18695);
nor U19264 (N_19264,N_18578,N_18280);
nor U19265 (N_19265,N_17693,N_18156);
xor U19266 (N_19266,N_17512,N_18024);
and U19267 (N_19267,N_18620,N_17730);
or U19268 (N_19268,N_18363,N_18446);
and U19269 (N_19269,N_18158,N_17790);
nor U19270 (N_19270,N_18196,N_18151);
nor U19271 (N_19271,N_18289,N_17964);
nand U19272 (N_19272,N_17882,N_18242);
nor U19273 (N_19273,N_17503,N_17778);
or U19274 (N_19274,N_17993,N_18269);
and U19275 (N_19275,N_17721,N_18478);
nor U19276 (N_19276,N_17828,N_17538);
and U19277 (N_19277,N_17587,N_18161);
or U19278 (N_19278,N_18715,N_18378);
xnor U19279 (N_19279,N_17646,N_18644);
xnor U19280 (N_19280,N_18559,N_17968);
and U19281 (N_19281,N_18416,N_17697);
nor U19282 (N_19282,N_18057,N_18331);
nor U19283 (N_19283,N_18643,N_17668);
and U19284 (N_19284,N_17591,N_18495);
or U19285 (N_19285,N_17647,N_18508);
and U19286 (N_19286,N_18437,N_17569);
nand U19287 (N_19287,N_18399,N_18144);
xnor U19288 (N_19288,N_18052,N_18285);
or U19289 (N_19289,N_18316,N_17998);
nor U19290 (N_19290,N_17562,N_18142);
xor U19291 (N_19291,N_17759,N_18568);
and U19292 (N_19292,N_17822,N_18332);
or U19293 (N_19293,N_18149,N_17910);
nor U19294 (N_19294,N_18462,N_18321);
xnor U19295 (N_19295,N_17784,N_17953);
or U19296 (N_19296,N_18676,N_17610);
nor U19297 (N_19297,N_17501,N_17575);
or U19298 (N_19298,N_18169,N_17873);
nand U19299 (N_19299,N_18228,N_18279);
nand U19300 (N_19300,N_17726,N_18455);
xnor U19301 (N_19301,N_18460,N_17913);
nor U19302 (N_19302,N_17842,N_17957);
nand U19303 (N_19303,N_17816,N_17776);
nor U19304 (N_19304,N_17554,N_17734);
and U19305 (N_19305,N_18419,N_18117);
xor U19306 (N_19306,N_18547,N_18338);
or U19307 (N_19307,N_18258,N_18712);
xnor U19308 (N_19308,N_18277,N_18123);
or U19309 (N_19309,N_18658,N_18086);
nor U19310 (N_19310,N_18171,N_17923);
nor U19311 (N_19311,N_18174,N_18343);
nand U19312 (N_19312,N_18749,N_17771);
xor U19313 (N_19313,N_17664,N_18060);
or U19314 (N_19314,N_18213,N_17695);
or U19315 (N_19315,N_18062,N_17766);
xnor U19316 (N_19316,N_18197,N_18682);
nand U19317 (N_19317,N_18070,N_17532);
and U19318 (N_19318,N_18296,N_17722);
nand U19319 (N_19319,N_18319,N_18132);
nand U19320 (N_19320,N_17618,N_17853);
or U19321 (N_19321,N_17796,N_17535);
xnor U19322 (N_19322,N_18243,N_18720);
nand U19323 (N_19323,N_17763,N_18090);
and U19324 (N_19324,N_18556,N_18322);
xnor U19325 (N_19325,N_18020,N_18355);
nor U19326 (N_19326,N_18210,N_17907);
or U19327 (N_19327,N_18186,N_18522);
xor U19328 (N_19328,N_18247,N_18271);
nor U19329 (N_19329,N_18746,N_18107);
nand U19330 (N_19330,N_17632,N_17672);
nor U19331 (N_19331,N_18472,N_18656);
xor U19332 (N_19332,N_18091,N_17700);
and U19333 (N_19333,N_17826,N_17914);
nor U19334 (N_19334,N_18265,N_18675);
or U19335 (N_19335,N_17544,N_17922);
or U19336 (N_19336,N_18570,N_18379);
or U19337 (N_19337,N_18088,N_18704);
nor U19338 (N_19338,N_17965,N_18581);
nor U19339 (N_19339,N_18386,N_18113);
and U19340 (N_19340,N_18486,N_17985);
nor U19341 (N_19341,N_18748,N_17837);
or U19342 (N_19342,N_18230,N_18127);
nor U19343 (N_19343,N_18579,N_18275);
and U19344 (N_19344,N_17537,N_17966);
or U19345 (N_19345,N_18415,N_18073);
xnor U19346 (N_19346,N_18006,N_18698);
nor U19347 (N_19347,N_17536,N_17539);
nor U19348 (N_19348,N_18506,N_18301);
nor U19349 (N_19349,N_17824,N_18385);
nor U19350 (N_19350,N_17737,N_17630);
or U19351 (N_19351,N_18513,N_17620);
nor U19352 (N_19352,N_18546,N_18408);
and U19353 (N_19353,N_18627,N_18172);
nand U19354 (N_19354,N_17765,N_18600);
xnor U19355 (N_19355,N_18504,N_18056);
or U19356 (N_19356,N_17570,N_17987);
xnor U19357 (N_19357,N_18646,N_18043);
nand U19358 (N_19358,N_18307,N_17747);
or U19359 (N_19359,N_18049,N_17707);
nand U19360 (N_19360,N_18431,N_18670);
nand U19361 (N_19361,N_17830,N_18490);
nor U19362 (N_19362,N_18637,N_18168);
and U19363 (N_19363,N_18300,N_18075);
and U19364 (N_19364,N_18136,N_18180);
nor U19365 (N_19365,N_18370,N_18368);
nor U19366 (N_19366,N_17719,N_17547);
xor U19367 (N_19367,N_17806,N_17891);
xor U19368 (N_19368,N_18679,N_18206);
and U19369 (N_19369,N_18530,N_18320);
or U19370 (N_19370,N_18626,N_17572);
or U19371 (N_19371,N_17812,N_18317);
xnor U19372 (N_19372,N_18318,N_18226);
xor U19373 (N_19373,N_18569,N_18685);
or U19374 (N_19374,N_17941,N_18201);
nor U19375 (N_19375,N_17788,N_18735);
and U19376 (N_19376,N_18343,N_18607);
nor U19377 (N_19377,N_17681,N_18402);
or U19378 (N_19378,N_18315,N_18024);
and U19379 (N_19379,N_17556,N_17707);
nand U19380 (N_19380,N_18169,N_17518);
nor U19381 (N_19381,N_18415,N_18598);
xnor U19382 (N_19382,N_18311,N_17685);
xor U19383 (N_19383,N_17816,N_17606);
and U19384 (N_19384,N_17814,N_17849);
nand U19385 (N_19385,N_18646,N_18747);
and U19386 (N_19386,N_18119,N_18197);
nor U19387 (N_19387,N_17578,N_18017);
nor U19388 (N_19388,N_18009,N_18269);
nand U19389 (N_19389,N_17643,N_17522);
xor U19390 (N_19390,N_17867,N_17635);
or U19391 (N_19391,N_18182,N_18033);
and U19392 (N_19392,N_17624,N_17943);
nand U19393 (N_19393,N_18685,N_18698);
or U19394 (N_19394,N_18233,N_18344);
and U19395 (N_19395,N_18559,N_18136);
and U19396 (N_19396,N_17823,N_18063);
nand U19397 (N_19397,N_18438,N_18046);
xnor U19398 (N_19398,N_17801,N_17871);
nor U19399 (N_19399,N_17950,N_17957);
xnor U19400 (N_19400,N_17733,N_17916);
nor U19401 (N_19401,N_17787,N_18704);
or U19402 (N_19402,N_18426,N_18667);
nand U19403 (N_19403,N_18453,N_18428);
or U19404 (N_19404,N_17835,N_18456);
or U19405 (N_19405,N_17859,N_18632);
xor U19406 (N_19406,N_18510,N_18655);
or U19407 (N_19407,N_17745,N_18464);
and U19408 (N_19408,N_18027,N_17701);
or U19409 (N_19409,N_18356,N_18363);
and U19410 (N_19410,N_17618,N_17873);
nand U19411 (N_19411,N_17945,N_18474);
nor U19412 (N_19412,N_17899,N_17635);
or U19413 (N_19413,N_18077,N_18703);
nand U19414 (N_19414,N_18441,N_17963);
or U19415 (N_19415,N_18560,N_17787);
or U19416 (N_19416,N_17596,N_17882);
nand U19417 (N_19417,N_18493,N_18473);
or U19418 (N_19418,N_18487,N_18036);
nand U19419 (N_19419,N_18080,N_18278);
and U19420 (N_19420,N_17536,N_18593);
nand U19421 (N_19421,N_17564,N_18350);
and U19422 (N_19422,N_17546,N_18652);
xor U19423 (N_19423,N_18425,N_18564);
nor U19424 (N_19424,N_18643,N_18185);
nand U19425 (N_19425,N_18716,N_18721);
and U19426 (N_19426,N_18491,N_17732);
nor U19427 (N_19427,N_18279,N_17655);
nor U19428 (N_19428,N_17655,N_18166);
nand U19429 (N_19429,N_17881,N_18540);
nor U19430 (N_19430,N_18218,N_18568);
and U19431 (N_19431,N_18346,N_17827);
nand U19432 (N_19432,N_17583,N_17999);
or U19433 (N_19433,N_18647,N_17716);
nand U19434 (N_19434,N_18506,N_17967);
nand U19435 (N_19435,N_17733,N_18342);
nand U19436 (N_19436,N_18710,N_18393);
xnor U19437 (N_19437,N_18337,N_17923);
and U19438 (N_19438,N_18377,N_18677);
or U19439 (N_19439,N_18324,N_17604);
and U19440 (N_19440,N_18688,N_18430);
or U19441 (N_19441,N_17907,N_18401);
or U19442 (N_19442,N_17969,N_17581);
xor U19443 (N_19443,N_17866,N_17859);
xor U19444 (N_19444,N_18123,N_18540);
or U19445 (N_19445,N_17884,N_18020);
nor U19446 (N_19446,N_18240,N_17839);
nand U19447 (N_19447,N_17920,N_17841);
nand U19448 (N_19448,N_18332,N_18176);
nor U19449 (N_19449,N_18014,N_18486);
nand U19450 (N_19450,N_17777,N_18236);
nor U19451 (N_19451,N_17687,N_17603);
and U19452 (N_19452,N_17912,N_18111);
xnor U19453 (N_19453,N_18210,N_18217);
nor U19454 (N_19454,N_18005,N_17767);
nand U19455 (N_19455,N_18506,N_17811);
nand U19456 (N_19456,N_18739,N_18650);
nor U19457 (N_19457,N_17924,N_18504);
nor U19458 (N_19458,N_17796,N_17949);
xnor U19459 (N_19459,N_17812,N_17759);
and U19460 (N_19460,N_17742,N_17781);
xnor U19461 (N_19461,N_18000,N_18144);
nor U19462 (N_19462,N_18495,N_18697);
or U19463 (N_19463,N_18596,N_17576);
nor U19464 (N_19464,N_18565,N_18172);
nand U19465 (N_19465,N_18069,N_17886);
xnor U19466 (N_19466,N_18399,N_18413);
and U19467 (N_19467,N_17502,N_18109);
or U19468 (N_19468,N_17504,N_18116);
xnor U19469 (N_19469,N_17514,N_18619);
nand U19470 (N_19470,N_17705,N_17966);
or U19471 (N_19471,N_18149,N_18324);
xor U19472 (N_19472,N_18663,N_18334);
or U19473 (N_19473,N_18694,N_17896);
nor U19474 (N_19474,N_18709,N_17561);
xor U19475 (N_19475,N_18042,N_17642);
xnor U19476 (N_19476,N_17515,N_18466);
nand U19477 (N_19477,N_18082,N_17602);
nand U19478 (N_19478,N_18031,N_17749);
nor U19479 (N_19479,N_17697,N_18305);
nand U19480 (N_19480,N_18692,N_17707);
or U19481 (N_19481,N_17834,N_18701);
nor U19482 (N_19482,N_17534,N_17648);
nand U19483 (N_19483,N_18048,N_17613);
or U19484 (N_19484,N_18247,N_18624);
or U19485 (N_19485,N_18510,N_17643);
or U19486 (N_19486,N_18236,N_17575);
and U19487 (N_19487,N_18209,N_17662);
xnor U19488 (N_19488,N_18586,N_17746);
or U19489 (N_19489,N_17760,N_17979);
or U19490 (N_19490,N_18181,N_18745);
or U19491 (N_19491,N_18385,N_17678);
xor U19492 (N_19492,N_17537,N_18019);
nand U19493 (N_19493,N_18607,N_18007);
nand U19494 (N_19494,N_18607,N_18553);
or U19495 (N_19495,N_17610,N_18202);
xnor U19496 (N_19496,N_17991,N_18278);
or U19497 (N_19497,N_17730,N_18659);
or U19498 (N_19498,N_17588,N_17601);
nand U19499 (N_19499,N_17654,N_17770);
nand U19500 (N_19500,N_18614,N_18678);
nand U19501 (N_19501,N_17738,N_18038);
xor U19502 (N_19502,N_18680,N_18312);
nand U19503 (N_19503,N_18183,N_17583);
or U19504 (N_19504,N_17797,N_18592);
nand U19505 (N_19505,N_18413,N_17511);
and U19506 (N_19506,N_18401,N_18317);
nor U19507 (N_19507,N_17814,N_18325);
and U19508 (N_19508,N_17721,N_18183);
xnor U19509 (N_19509,N_18656,N_17923);
or U19510 (N_19510,N_18631,N_18130);
nand U19511 (N_19511,N_17890,N_18472);
nand U19512 (N_19512,N_18348,N_18533);
nand U19513 (N_19513,N_18086,N_17988);
nand U19514 (N_19514,N_18329,N_17708);
or U19515 (N_19515,N_18425,N_18545);
or U19516 (N_19516,N_18142,N_17790);
and U19517 (N_19517,N_18379,N_17732);
xnor U19518 (N_19518,N_18228,N_17785);
nand U19519 (N_19519,N_17631,N_18386);
or U19520 (N_19520,N_17896,N_18570);
nand U19521 (N_19521,N_18215,N_18212);
nor U19522 (N_19522,N_18272,N_18616);
or U19523 (N_19523,N_18092,N_18405);
xnor U19524 (N_19524,N_18593,N_18540);
xor U19525 (N_19525,N_18035,N_18454);
or U19526 (N_19526,N_17663,N_17884);
or U19527 (N_19527,N_17987,N_17894);
nor U19528 (N_19528,N_18484,N_17944);
or U19529 (N_19529,N_18126,N_17879);
or U19530 (N_19530,N_18209,N_18165);
nand U19531 (N_19531,N_17609,N_17768);
or U19532 (N_19532,N_18453,N_18730);
nand U19533 (N_19533,N_17985,N_18359);
nor U19534 (N_19534,N_18104,N_17909);
nor U19535 (N_19535,N_18564,N_17516);
and U19536 (N_19536,N_17900,N_17606);
nand U19537 (N_19537,N_17792,N_17743);
or U19538 (N_19538,N_18196,N_18313);
nand U19539 (N_19539,N_18209,N_18299);
or U19540 (N_19540,N_17893,N_17703);
xnor U19541 (N_19541,N_17912,N_18194);
or U19542 (N_19542,N_18616,N_17837);
nand U19543 (N_19543,N_17821,N_17710);
and U19544 (N_19544,N_18197,N_18088);
xor U19545 (N_19545,N_17838,N_17619);
xor U19546 (N_19546,N_18039,N_18162);
xor U19547 (N_19547,N_18685,N_17612);
nor U19548 (N_19548,N_18323,N_18290);
nor U19549 (N_19549,N_17753,N_18174);
or U19550 (N_19550,N_17863,N_18504);
nand U19551 (N_19551,N_17518,N_18737);
nand U19552 (N_19552,N_18036,N_18168);
and U19553 (N_19553,N_17859,N_18399);
nand U19554 (N_19554,N_18592,N_18417);
xor U19555 (N_19555,N_18278,N_17736);
nor U19556 (N_19556,N_17884,N_17698);
nor U19557 (N_19557,N_17756,N_18716);
and U19558 (N_19558,N_18349,N_17638);
and U19559 (N_19559,N_18204,N_17590);
nand U19560 (N_19560,N_18228,N_18330);
nand U19561 (N_19561,N_17741,N_18159);
nor U19562 (N_19562,N_18554,N_17673);
and U19563 (N_19563,N_17746,N_17734);
nand U19564 (N_19564,N_17647,N_18273);
nor U19565 (N_19565,N_17793,N_18330);
and U19566 (N_19566,N_18661,N_17923);
nor U19567 (N_19567,N_17747,N_18192);
or U19568 (N_19568,N_17682,N_17866);
nand U19569 (N_19569,N_18364,N_18490);
and U19570 (N_19570,N_18567,N_18498);
nand U19571 (N_19571,N_18516,N_17511);
and U19572 (N_19572,N_18333,N_17662);
and U19573 (N_19573,N_18322,N_17597);
nor U19574 (N_19574,N_17760,N_18100);
nand U19575 (N_19575,N_18340,N_18101);
nor U19576 (N_19576,N_18059,N_17609);
and U19577 (N_19577,N_18613,N_18550);
or U19578 (N_19578,N_17912,N_18043);
or U19579 (N_19579,N_18108,N_18499);
and U19580 (N_19580,N_18156,N_18344);
or U19581 (N_19581,N_17677,N_18399);
xnor U19582 (N_19582,N_18372,N_17838);
xor U19583 (N_19583,N_18409,N_18705);
xor U19584 (N_19584,N_18257,N_17914);
and U19585 (N_19585,N_17950,N_18493);
nor U19586 (N_19586,N_18295,N_17550);
and U19587 (N_19587,N_17515,N_18700);
xor U19588 (N_19588,N_17509,N_17603);
nor U19589 (N_19589,N_17804,N_18052);
nor U19590 (N_19590,N_18303,N_17649);
nor U19591 (N_19591,N_18210,N_17967);
nand U19592 (N_19592,N_18197,N_17567);
nor U19593 (N_19593,N_18327,N_17977);
nor U19594 (N_19594,N_18530,N_18588);
nor U19595 (N_19595,N_17567,N_18299);
nor U19596 (N_19596,N_18622,N_18207);
nor U19597 (N_19597,N_17666,N_18120);
xnor U19598 (N_19598,N_17644,N_18075);
or U19599 (N_19599,N_18318,N_17754);
nand U19600 (N_19600,N_17564,N_18256);
nand U19601 (N_19601,N_18203,N_17754);
xnor U19602 (N_19602,N_18682,N_18049);
and U19603 (N_19603,N_17799,N_17994);
nand U19604 (N_19604,N_17985,N_17600);
and U19605 (N_19605,N_17921,N_18118);
and U19606 (N_19606,N_18658,N_18379);
nand U19607 (N_19607,N_18208,N_17505);
or U19608 (N_19608,N_17946,N_18267);
and U19609 (N_19609,N_18021,N_17543);
and U19610 (N_19610,N_18494,N_18492);
nand U19611 (N_19611,N_18541,N_17899);
and U19612 (N_19612,N_17520,N_17612);
or U19613 (N_19613,N_17648,N_18544);
xor U19614 (N_19614,N_18521,N_17634);
and U19615 (N_19615,N_17947,N_18358);
or U19616 (N_19616,N_17569,N_17900);
and U19617 (N_19617,N_17644,N_18538);
nor U19618 (N_19618,N_18455,N_17516);
and U19619 (N_19619,N_18300,N_18256);
or U19620 (N_19620,N_18335,N_18633);
xnor U19621 (N_19621,N_18004,N_17733);
and U19622 (N_19622,N_17999,N_18685);
xor U19623 (N_19623,N_17964,N_18638);
and U19624 (N_19624,N_18521,N_18366);
and U19625 (N_19625,N_18426,N_18065);
or U19626 (N_19626,N_18602,N_18650);
nor U19627 (N_19627,N_18553,N_18038);
nand U19628 (N_19628,N_17903,N_18498);
and U19629 (N_19629,N_17960,N_18697);
or U19630 (N_19630,N_18611,N_18635);
nand U19631 (N_19631,N_18182,N_18334);
xor U19632 (N_19632,N_17833,N_17727);
and U19633 (N_19633,N_18627,N_18114);
nand U19634 (N_19634,N_18384,N_18343);
nor U19635 (N_19635,N_17654,N_17760);
nor U19636 (N_19636,N_18677,N_17653);
nor U19637 (N_19637,N_18189,N_18057);
xnor U19638 (N_19638,N_18284,N_17983);
xor U19639 (N_19639,N_17859,N_18146);
and U19640 (N_19640,N_17529,N_17823);
or U19641 (N_19641,N_17530,N_18455);
nand U19642 (N_19642,N_18584,N_17841);
nor U19643 (N_19643,N_17738,N_18416);
and U19644 (N_19644,N_18151,N_18706);
or U19645 (N_19645,N_17672,N_17788);
or U19646 (N_19646,N_18745,N_17599);
or U19647 (N_19647,N_18625,N_17534);
nor U19648 (N_19648,N_17532,N_18035);
or U19649 (N_19649,N_17563,N_18018);
or U19650 (N_19650,N_17772,N_17902);
or U19651 (N_19651,N_17674,N_18305);
xnor U19652 (N_19652,N_18500,N_18505);
and U19653 (N_19653,N_18339,N_18649);
and U19654 (N_19654,N_18057,N_17917);
or U19655 (N_19655,N_18595,N_18098);
or U19656 (N_19656,N_18026,N_17775);
nor U19657 (N_19657,N_18272,N_18508);
nand U19658 (N_19658,N_17646,N_17958);
or U19659 (N_19659,N_18531,N_18340);
nor U19660 (N_19660,N_17942,N_17793);
and U19661 (N_19661,N_18233,N_17718);
or U19662 (N_19662,N_18383,N_18537);
and U19663 (N_19663,N_18282,N_17556);
or U19664 (N_19664,N_17871,N_18157);
nand U19665 (N_19665,N_17550,N_18546);
nand U19666 (N_19666,N_18440,N_17515);
nand U19667 (N_19667,N_18288,N_17733);
xnor U19668 (N_19668,N_18532,N_18514);
nor U19669 (N_19669,N_18250,N_18358);
nor U19670 (N_19670,N_18639,N_18693);
or U19671 (N_19671,N_18058,N_18605);
or U19672 (N_19672,N_17565,N_17834);
xor U19673 (N_19673,N_18154,N_17770);
nor U19674 (N_19674,N_18677,N_18132);
nand U19675 (N_19675,N_18553,N_18645);
xnor U19676 (N_19676,N_18566,N_18099);
nand U19677 (N_19677,N_17529,N_17685);
or U19678 (N_19678,N_17848,N_18660);
and U19679 (N_19679,N_18145,N_17779);
xor U19680 (N_19680,N_18132,N_18639);
or U19681 (N_19681,N_18270,N_17553);
xor U19682 (N_19682,N_18361,N_17704);
or U19683 (N_19683,N_17538,N_18654);
nand U19684 (N_19684,N_17824,N_18046);
nor U19685 (N_19685,N_18253,N_18356);
nand U19686 (N_19686,N_18452,N_18370);
or U19687 (N_19687,N_18102,N_17641);
nand U19688 (N_19688,N_17941,N_17981);
and U19689 (N_19689,N_17791,N_17501);
nor U19690 (N_19690,N_18430,N_18739);
and U19691 (N_19691,N_18040,N_17537);
nor U19692 (N_19692,N_18376,N_18403);
nor U19693 (N_19693,N_18495,N_17539);
and U19694 (N_19694,N_18240,N_18096);
nor U19695 (N_19695,N_18173,N_17995);
nor U19696 (N_19696,N_18601,N_18308);
and U19697 (N_19697,N_18010,N_18591);
and U19698 (N_19698,N_18485,N_18434);
xnor U19699 (N_19699,N_17952,N_18377);
or U19700 (N_19700,N_18109,N_17718);
or U19701 (N_19701,N_17553,N_17951);
xor U19702 (N_19702,N_18422,N_18546);
and U19703 (N_19703,N_17751,N_18265);
xnor U19704 (N_19704,N_17710,N_18312);
nor U19705 (N_19705,N_17659,N_18047);
xor U19706 (N_19706,N_17957,N_18111);
nor U19707 (N_19707,N_18553,N_18021);
or U19708 (N_19708,N_18094,N_18499);
nor U19709 (N_19709,N_17923,N_18444);
or U19710 (N_19710,N_17867,N_17768);
nand U19711 (N_19711,N_17974,N_18070);
xor U19712 (N_19712,N_17931,N_18542);
nand U19713 (N_19713,N_17654,N_18464);
or U19714 (N_19714,N_17893,N_18098);
or U19715 (N_19715,N_18185,N_18240);
nand U19716 (N_19716,N_17794,N_17597);
nor U19717 (N_19717,N_18013,N_18244);
or U19718 (N_19718,N_17893,N_18148);
nand U19719 (N_19719,N_18227,N_17758);
and U19720 (N_19720,N_18688,N_18082);
xnor U19721 (N_19721,N_18466,N_18383);
nor U19722 (N_19722,N_18346,N_18298);
nor U19723 (N_19723,N_18092,N_18349);
and U19724 (N_19724,N_17546,N_18598);
nor U19725 (N_19725,N_17730,N_17912);
nand U19726 (N_19726,N_17519,N_18117);
and U19727 (N_19727,N_17703,N_17602);
and U19728 (N_19728,N_17614,N_17944);
nand U19729 (N_19729,N_18217,N_17648);
and U19730 (N_19730,N_18604,N_17659);
xor U19731 (N_19731,N_18319,N_17862);
nor U19732 (N_19732,N_17815,N_18521);
xor U19733 (N_19733,N_18662,N_18579);
xor U19734 (N_19734,N_18052,N_17730);
nand U19735 (N_19735,N_17844,N_17770);
nor U19736 (N_19736,N_18239,N_18330);
nor U19737 (N_19737,N_18139,N_18339);
xor U19738 (N_19738,N_18327,N_17592);
nand U19739 (N_19739,N_18071,N_18641);
and U19740 (N_19740,N_18204,N_17967);
nor U19741 (N_19741,N_18731,N_18432);
and U19742 (N_19742,N_17721,N_17881);
nor U19743 (N_19743,N_18275,N_17906);
or U19744 (N_19744,N_18098,N_17962);
and U19745 (N_19745,N_18227,N_17629);
nor U19746 (N_19746,N_18399,N_18388);
xor U19747 (N_19747,N_18225,N_17963);
or U19748 (N_19748,N_18244,N_17599);
or U19749 (N_19749,N_18627,N_17529);
nand U19750 (N_19750,N_18426,N_17502);
and U19751 (N_19751,N_18657,N_17525);
nor U19752 (N_19752,N_18105,N_18178);
nor U19753 (N_19753,N_17645,N_18364);
and U19754 (N_19754,N_17950,N_18484);
xor U19755 (N_19755,N_18023,N_18269);
xnor U19756 (N_19756,N_18319,N_18255);
and U19757 (N_19757,N_17734,N_18344);
nand U19758 (N_19758,N_18653,N_17879);
and U19759 (N_19759,N_18393,N_17609);
nor U19760 (N_19760,N_18460,N_18126);
nand U19761 (N_19761,N_18044,N_17501);
nor U19762 (N_19762,N_18402,N_17544);
and U19763 (N_19763,N_18113,N_17859);
xnor U19764 (N_19764,N_18201,N_17750);
nor U19765 (N_19765,N_18623,N_18233);
and U19766 (N_19766,N_17876,N_18569);
xor U19767 (N_19767,N_18068,N_17792);
nor U19768 (N_19768,N_17878,N_17882);
nor U19769 (N_19769,N_18050,N_18471);
and U19770 (N_19770,N_18692,N_18166);
or U19771 (N_19771,N_18478,N_18507);
and U19772 (N_19772,N_18171,N_17941);
or U19773 (N_19773,N_18504,N_18135);
xnor U19774 (N_19774,N_18202,N_18516);
and U19775 (N_19775,N_18610,N_18389);
xor U19776 (N_19776,N_17520,N_18085);
nor U19777 (N_19777,N_18186,N_18060);
nor U19778 (N_19778,N_18720,N_18048);
xnor U19779 (N_19779,N_17668,N_17879);
or U19780 (N_19780,N_18546,N_17586);
nand U19781 (N_19781,N_18706,N_18645);
nand U19782 (N_19782,N_17622,N_17767);
and U19783 (N_19783,N_18514,N_18140);
nor U19784 (N_19784,N_17658,N_18265);
nand U19785 (N_19785,N_18182,N_17911);
or U19786 (N_19786,N_18617,N_17869);
nor U19787 (N_19787,N_17721,N_17923);
xnor U19788 (N_19788,N_17857,N_18506);
nor U19789 (N_19789,N_17669,N_18014);
nor U19790 (N_19790,N_17995,N_18518);
nor U19791 (N_19791,N_17775,N_18482);
xnor U19792 (N_19792,N_17921,N_18116);
nand U19793 (N_19793,N_17721,N_18162);
and U19794 (N_19794,N_18400,N_17962);
nand U19795 (N_19795,N_18638,N_17775);
xor U19796 (N_19796,N_17560,N_18212);
and U19797 (N_19797,N_18491,N_17977);
and U19798 (N_19798,N_17905,N_18536);
nand U19799 (N_19799,N_18663,N_18235);
nand U19800 (N_19800,N_17626,N_17617);
nand U19801 (N_19801,N_17926,N_17771);
nand U19802 (N_19802,N_18395,N_17918);
or U19803 (N_19803,N_17558,N_18066);
and U19804 (N_19804,N_17952,N_18393);
or U19805 (N_19805,N_17914,N_17830);
or U19806 (N_19806,N_18666,N_18553);
nand U19807 (N_19807,N_17792,N_18088);
xor U19808 (N_19808,N_17592,N_17922);
xnor U19809 (N_19809,N_17679,N_18566);
xor U19810 (N_19810,N_18448,N_18737);
and U19811 (N_19811,N_18252,N_17808);
xnor U19812 (N_19812,N_18684,N_18733);
xor U19813 (N_19813,N_17725,N_18622);
nand U19814 (N_19814,N_18726,N_18465);
and U19815 (N_19815,N_17525,N_18614);
xor U19816 (N_19816,N_18232,N_18667);
nand U19817 (N_19817,N_18374,N_18684);
and U19818 (N_19818,N_18598,N_17948);
nor U19819 (N_19819,N_17920,N_17664);
nor U19820 (N_19820,N_18363,N_18545);
and U19821 (N_19821,N_17868,N_17659);
and U19822 (N_19822,N_17665,N_17618);
nand U19823 (N_19823,N_18066,N_18048);
xnor U19824 (N_19824,N_17504,N_17516);
nor U19825 (N_19825,N_18284,N_18429);
xnor U19826 (N_19826,N_18372,N_17835);
xnor U19827 (N_19827,N_18206,N_18139);
and U19828 (N_19828,N_18049,N_18260);
or U19829 (N_19829,N_17564,N_17500);
xnor U19830 (N_19830,N_18556,N_17832);
and U19831 (N_19831,N_17562,N_18333);
nor U19832 (N_19832,N_18463,N_18152);
nor U19833 (N_19833,N_17969,N_17576);
xnor U19834 (N_19834,N_18568,N_18662);
or U19835 (N_19835,N_17615,N_18468);
and U19836 (N_19836,N_18257,N_17628);
xnor U19837 (N_19837,N_17823,N_17974);
or U19838 (N_19838,N_17960,N_17773);
nand U19839 (N_19839,N_18321,N_18511);
xor U19840 (N_19840,N_18078,N_17894);
xor U19841 (N_19841,N_17897,N_18416);
nor U19842 (N_19842,N_18169,N_18149);
and U19843 (N_19843,N_18552,N_17767);
and U19844 (N_19844,N_18110,N_17997);
and U19845 (N_19845,N_18524,N_17691);
xnor U19846 (N_19846,N_18402,N_18092);
nand U19847 (N_19847,N_17696,N_17553);
and U19848 (N_19848,N_17998,N_17599);
or U19849 (N_19849,N_18488,N_17766);
and U19850 (N_19850,N_18252,N_18190);
or U19851 (N_19851,N_18074,N_17777);
nand U19852 (N_19852,N_17898,N_17799);
or U19853 (N_19853,N_17712,N_18171);
nor U19854 (N_19854,N_17755,N_17668);
and U19855 (N_19855,N_17593,N_18003);
nand U19856 (N_19856,N_17646,N_18034);
or U19857 (N_19857,N_17620,N_18278);
and U19858 (N_19858,N_18524,N_18601);
nand U19859 (N_19859,N_18399,N_18593);
xor U19860 (N_19860,N_18067,N_17604);
xnor U19861 (N_19861,N_18340,N_18569);
nor U19862 (N_19862,N_18212,N_17936);
nand U19863 (N_19863,N_17753,N_18437);
and U19864 (N_19864,N_18297,N_18434);
xnor U19865 (N_19865,N_17857,N_18403);
nor U19866 (N_19866,N_18387,N_18207);
and U19867 (N_19867,N_18439,N_18256);
xnor U19868 (N_19868,N_18104,N_18298);
xor U19869 (N_19869,N_17897,N_18047);
and U19870 (N_19870,N_17662,N_17784);
and U19871 (N_19871,N_18637,N_18415);
or U19872 (N_19872,N_17811,N_17941);
and U19873 (N_19873,N_18061,N_18631);
nor U19874 (N_19874,N_18228,N_18018);
xnor U19875 (N_19875,N_18166,N_18054);
nor U19876 (N_19876,N_18563,N_17551);
or U19877 (N_19877,N_18195,N_18660);
nand U19878 (N_19878,N_17577,N_18354);
nor U19879 (N_19879,N_18497,N_18288);
or U19880 (N_19880,N_18482,N_18544);
nor U19881 (N_19881,N_17614,N_17804);
or U19882 (N_19882,N_18555,N_18619);
and U19883 (N_19883,N_17560,N_18306);
or U19884 (N_19884,N_18172,N_18163);
xnor U19885 (N_19885,N_18589,N_17704);
nand U19886 (N_19886,N_18514,N_17652);
and U19887 (N_19887,N_17537,N_17829);
and U19888 (N_19888,N_18146,N_17693);
nand U19889 (N_19889,N_18591,N_18462);
nand U19890 (N_19890,N_18585,N_18186);
nor U19891 (N_19891,N_18723,N_18484);
xnor U19892 (N_19892,N_17793,N_17610);
and U19893 (N_19893,N_18445,N_17682);
nor U19894 (N_19894,N_17738,N_18662);
nor U19895 (N_19895,N_17594,N_17670);
or U19896 (N_19896,N_18535,N_17611);
xor U19897 (N_19897,N_17656,N_18011);
or U19898 (N_19898,N_18607,N_17774);
nor U19899 (N_19899,N_17779,N_17906);
xnor U19900 (N_19900,N_17670,N_17997);
xor U19901 (N_19901,N_18314,N_17805);
xor U19902 (N_19902,N_18267,N_18725);
nand U19903 (N_19903,N_18455,N_17987);
nand U19904 (N_19904,N_17666,N_18063);
nor U19905 (N_19905,N_18241,N_18139);
xor U19906 (N_19906,N_17733,N_18436);
xor U19907 (N_19907,N_18561,N_18577);
nand U19908 (N_19908,N_18042,N_17576);
or U19909 (N_19909,N_17774,N_18164);
and U19910 (N_19910,N_17858,N_18565);
nand U19911 (N_19911,N_18714,N_17966);
nand U19912 (N_19912,N_18252,N_18468);
and U19913 (N_19913,N_18304,N_18440);
xor U19914 (N_19914,N_17828,N_17798);
nor U19915 (N_19915,N_18097,N_18528);
xnor U19916 (N_19916,N_18268,N_18669);
and U19917 (N_19917,N_18118,N_17617);
or U19918 (N_19918,N_17833,N_18540);
xor U19919 (N_19919,N_18026,N_17548);
xnor U19920 (N_19920,N_18490,N_17610);
xnor U19921 (N_19921,N_18009,N_18036);
and U19922 (N_19922,N_18406,N_17546);
nor U19923 (N_19923,N_17508,N_18643);
nor U19924 (N_19924,N_18494,N_18056);
and U19925 (N_19925,N_17545,N_18646);
nand U19926 (N_19926,N_18348,N_18636);
nor U19927 (N_19927,N_17995,N_17863);
or U19928 (N_19928,N_17817,N_18589);
and U19929 (N_19929,N_17512,N_18386);
nor U19930 (N_19930,N_18343,N_17697);
nor U19931 (N_19931,N_17626,N_17721);
xor U19932 (N_19932,N_18541,N_17989);
or U19933 (N_19933,N_18133,N_18195);
nand U19934 (N_19934,N_18319,N_18054);
xnor U19935 (N_19935,N_18707,N_18247);
and U19936 (N_19936,N_18452,N_18518);
nand U19937 (N_19937,N_17787,N_18150);
xor U19938 (N_19938,N_17504,N_18600);
nor U19939 (N_19939,N_17831,N_18556);
and U19940 (N_19940,N_17796,N_18309);
xnor U19941 (N_19941,N_18548,N_18472);
xnor U19942 (N_19942,N_18662,N_17527);
nand U19943 (N_19943,N_17872,N_18465);
and U19944 (N_19944,N_18242,N_18081);
nor U19945 (N_19945,N_18210,N_18051);
xnor U19946 (N_19946,N_18182,N_18040);
xnor U19947 (N_19947,N_18469,N_18512);
xnor U19948 (N_19948,N_17932,N_17899);
nor U19949 (N_19949,N_18481,N_17570);
nor U19950 (N_19950,N_18588,N_17543);
or U19951 (N_19951,N_18211,N_18228);
nand U19952 (N_19952,N_18184,N_18348);
xnor U19953 (N_19953,N_17851,N_18546);
nor U19954 (N_19954,N_17823,N_18617);
and U19955 (N_19955,N_17512,N_18728);
nand U19956 (N_19956,N_18405,N_18586);
xor U19957 (N_19957,N_18135,N_18227);
and U19958 (N_19958,N_18298,N_17822);
nor U19959 (N_19959,N_17881,N_17684);
xnor U19960 (N_19960,N_17997,N_18729);
nor U19961 (N_19961,N_17973,N_18406);
nor U19962 (N_19962,N_18087,N_18706);
xnor U19963 (N_19963,N_17950,N_18440);
nand U19964 (N_19964,N_17933,N_17555);
nor U19965 (N_19965,N_18075,N_18382);
and U19966 (N_19966,N_17530,N_17625);
and U19967 (N_19967,N_18155,N_17703);
xor U19968 (N_19968,N_18616,N_18519);
or U19969 (N_19969,N_18340,N_17792);
or U19970 (N_19970,N_18366,N_18577);
and U19971 (N_19971,N_18739,N_18449);
or U19972 (N_19972,N_18259,N_18099);
nand U19973 (N_19973,N_18140,N_18498);
and U19974 (N_19974,N_17698,N_17746);
nand U19975 (N_19975,N_17787,N_18495);
xnor U19976 (N_19976,N_18641,N_17850);
or U19977 (N_19977,N_18495,N_17752);
nand U19978 (N_19978,N_17599,N_18514);
xnor U19979 (N_19979,N_17903,N_18181);
or U19980 (N_19980,N_18463,N_18558);
nor U19981 (N_19981,N_18491,N_17504);
and U19982 (N_19982,N_18166,N_18667);
or U19983 (N_19983,N_18493,N_17696);
or U19984 (N_19984,N_18156,N_17720);
nor U19985 (N_19985,N_18331,N_18595);
xor U19986 (N_19986,N_17947,N_18700);
and U19987 (N_19987,N_18091,N_18074);
nand U19988 (N_19988,N_18635,N_18487);
and U19989 (N_19989,N_18416,N_18602);
nand U19990 (N_19990,N_17522,N_17864);
and U19991 (N_19991,N_17582,N_18489);
or U19992 (N_19992,N_18314,N_18449);
or U19993 (N_19993,N_18064,N_18686);
or U19994 (N_19994,N_18115,N_17987);
xnor U19995 (N_19995,N_18698,N_17958);
xor U19996 (N_19996,N_18222,N_17830);
nor U19997 (N_19997,N_18626,N_18315);
or U19998 (N_19998,N_17983,N_17741);
or U19999 (N_19999,N_17842,N_18342);
or U20000 (N_20000,N_19827,N_19854);
or U20001 (N_20001,N_19253,N_19336);
or U20002 (N_20002,N_19770,N_18796);
nand U20003 (N_20003,N_18845,N_19126);
nor U20004 (N_20004,N_19276,N_19756);
or U20005 (N_20005,N_19286,N_19605);
nand U20006 (N_20006,N_19759,N_19178);
and U20007 (N_20007,N_19179,N_19504);
nor U20008 (N_20008,N_19769,N_19739);
nand U20009 (N_20009,N_19071,N_19172);
and U20010 (N_20010,N_19238,N_18899);
nor U20011 (N_20011,N_19628,N_19439);
nor U20012 (N_20012,N_19932,N_18959);
xor U20013 (N_20013,N_19965,N_19988);
nand U20014 (N_20014,N_19799,N_19395);
or U20015 (N_20015,N_18925,N_19197);
nor U20016 (N_20016,N_19270,N_19714);
nor U20017 (N_20017,N_18986,N_19948);
or U20018 (N_20018,N_19680,N_19506);
nor U20019 (N_20019,N_19423,N_19529);
or U20020 (N_20020,N_19848,N_19855);
or U20021 (N_20021,N_18963,N_19791);
nand U20022 (N_20022,N_19852,N_19562);
nand U20023 (N_20023,N_19694,N_19331);
nand U20024 (N_20024,N_19184,N_19260);
nand U20025 (N_20025,N_19840,N_19925);
and U20026 (N_20026,N_19732,N_19100);
and U20027 (N_20027,N_19899,N_19651);
or U20028 (N_20028,N_18926,N_19895);
or U20029 (N_20029,N_19746,N_19048);
or U20030 (N_20030,N_18768,N_19715);
and U20031 (N_20031,N_19356,N_18888);
nand U20032 (N_20032,N_19523,N_18822);
or U20033 (N_20033,N_19365,N_18785);
or U20034 (N_20034,N_18983,N_19877);
and U20035 (N_20035,N_19914,N_19296);
nand U20036 (N_20036,N_18827,N_19979);
nand U20037 (N_20037,N_18901,N_19836);
nor U20038 (N_20038,N_19552,N_19265);
nand U20039 (N_20039,N_19986,N_18981);
xnor U20040 (N_20040,N_19316,N_19291);
xor U20041 (N_20041,N_19751,N_19239);
or U20042 (N_20042,N_18994,N_19707);
nor U20043 (N_20043,N_18880,N_19340);
nor U20044 (N_20044,N_19224,N_19460);
and U20045 (N_20045,N_19020,N_19893);
nor U20046 (N_20046,N_19273,N_19226);
nor U20047 (N_20047,N_19377,N_19962);
or U20048 (N_20048,N_19322,N_19402);
and U20049 (N_20049,N_19109,N_19674);
nand U20050 (N_20050,N_19061,N_19691);
nor U20051 (N_20051,N_19210,N_19474);
xnor U20052 (N_20052,N_19931,N_19897);
xor U20053 (N_20053,N_19404,N_19361);
nand U20054 (N_20054,N_19718,N_19440);
xnor U20055 (N_20055,N_19611,N_18951);
nand U20056 (N_20056,N_19119,N_19295);
xnor U20057 (N_20057,N_19704,N_19645);
or U20058 (N_20058,N_18988,N_18887);
or U20059 (N_20059,N_19234,N_19810);
nand U20060 (N_20060,N_19868,N_19505);
or U20061 (N_20061,N_19266,N_19441);
or U20062 (N_20062,N_19698,N_19211);
xnor U20063 (N_20063,N_19060,N_19851);
nand U20064 (N_20064,N_19695,N_19304);
nor U20065 (N_20065,N_19157,N_19194);
and U20066 (N_20066,N_19815,N_19251);
nor U20067 (N_20067,N_18977,N_19442);
nor U20068 (N_20068,N_19149,N_19864);
nor U20069 (N_20069,N_18933,N_18914);
nand U20070 (N_20070,N_19901,N_19632);
or U20071 (N_20071,N_18857,N_19867);
nor U20072 (N_20072,N_19880,N_19987);
and U20073 (N_20073,N_19189,N_19761);
nor U20074 (N_20074,N_19067,N_19950);
xor U20075 (N_20075,N_19713,N_18777);
nand U20076 (N_20076,N_19858,N_19937);
and U20077 (N_20077,N_19958,N_19831);
nand U20078 (N_20078,N_19603,N_19724);
nor U20079 (N_20079,N_19596,N_19127);
xnor U20080 (N_20080,N_19911,N_18776);
nor U20081 (N_20081,N_19064,N_18818);
or U20082 (N_20082,N_19777,N_19982);
nor U20083 (N_20083,N_18786,N_19412);
or U20084 (N_20084,N_19920,N_18831);
nor U20085 (N_20085,N_19472,N_18832);
and U20086 (N_20086,N_19641,N_18945);
nor U20087 (N_20087,N_19470,N_19346);
nor U20088 (N_20088,N_19731,N_19708);
or U20089 (N_20089,N_19215,N_19405);
and U20090 (N_20090,N_19323,N_18927);
or U20091 (N_20091,N_19923,N_19083);
nand U20092 (N_20092,N_19057,N_18921);
and U20093 (N_20093,N_18908,N_19183);
or U20094 (N_20094,N_18979,N_19294);
or U20095 (N_20095,N_19092,N_19499);
nand U20096 (N_20096,N_19495,N_19003);
xor U20097 (N_20097,N_18969,N_19491);
nand U20098 (N_20098,N_19550,N_19303);
nor U20099 (N_20099,N_18974,N_19916);
xnor U20100 (N_20100,N_19776,N_18895);
and U20101 (N_20101,N_19146,N_19298);
nor U20102 (N_20102,N_19383,N_19849);
xnor U20103 (N_20103,N_18987,N_19409);
and U20104 (N_20104,N_19185,N_18837);
and U20105 (N_20105,N_19534,N_19585);
xnor U20106 (N_20106,N_19110,N_19314);
and U20107 (N_20107,N_19106,N_19587);
nor U20108 (N_20108,N_19391,N_19445);
nand U20109 (N_20109,N_19835,N_19271);
or U20110 (N_20110,N_19640,N_19220);
or U20111 (N_20111,N_19861,N_19337);
or U20112 (N_20112,N_19588,N_19050);
nand U20113 (N_20113,N_19249,N_19168);
nor U20114 (N_20114,N_19737,N_19629);
xnor U20115 (N_20115,N_19686,N_19281);
nor U20116 (N_20116,N_19334,N_19417);
or U20117 (N_20117,N_19828,N_19150);
and U20118 (N_20118,N_19556,N_18976);
xnor U20119 (N_20119,N_19338,N_19765);
or U20120 (N_20120,N_19516,N_19188);
or U20121 (N_20121,N_19860,N_19447);
nand U20122 (N_20122,N_19977,N_19614);
nor U20123 (N_20123,N_19859,N_19206);
and U20124 (N_20124,N_18817,N_19221);
or U20125 (N_20125,N_19646,N_19572);
nand U20126 (N_20126,N_18999,N_19151);
or U20127 (N_20127,N_19597,N_18767);
or U20128 (N_20128,N_19915,N_18897);
or U20129 (N_20129,N_19566,N_19021);
nand U20130 (N_20130,N_19584,N_19205);
xnor U20131 (N_20131,N_19526,N_18828);
xor U20132 (N_20132,N_19382,N_18788);
xnor U20133 (N_20133,N_19532,N_18771);
and U20134 (N_20134,N_19175,N_19466);
nand U20135 (N_20135,N_19326,N_19002);
and U20136 (N_20136,N_18756,N_19033);
nand U20137 (N_20137,N_19519,N_19075);
and U20138 (N_20138,N_18755,N_19991);
xor U20139 (N_20139,N_19501,N_19481);
nand U20140 (N_20140,N_18902,N_19803);
nand U20141 (N_20141,N_19652,N_19077);
nor U20142 (N_20142,N_19560,N_18973);
nand U20143 (N_20143,N_19623,N_19236);
or U20144 (N_20144,N_18968,N_19416);
and U20145 (N_20145,N_19606,N_19421);
and U20146 (N_20146,N_18795,N_18890);
or U20147 (N_20147,N_19872,N_19881);
and U20148 (N_20148,N_19009,N_19284);
nand U20149 (N_20149,N_18836,N_19288);
nand U20150 (N_20150,N_19181,N_19689);
or U20151 (N_20151,N_19531,N_19613);
nor U20152 (N_20152,N_19419,N_19863);
or U20153 (N_20153,N_19414,N_19829);
nor U20154 (N_20154,N_19214,N_19318);
xor U20155 (N_20155,N_18884,N_19463);
nor U20156 (N_20156,N_18790,N_19424);
or U20157 (N_20157,N_19263,N_19115);
xor U20158 (N_20158,N_19943,N_19927);
xor U20159 (N_20159,N_19237,N_19794);
nand U20160 (N_20160,N_19299,N_19166);
or U20161 (N_20161,N_19575,N_19679);
nor U20162 (N_20162,N_18970,N_19600);
or U20163 (N_20163,N_19653,N_19685);
nand U20164 (N_20164,N_19367,N_19553);
or U20165 (N_20165,N_19489,N_18954);
or U20166 (N_20166,N_19257,N_19569);
xor U20167 (N_20167,N_19242,N_19443);
xor U20168 (N_20168,N_19480,N_18995);
or U20169 (N_20169,N_19591,N_19675);
nand U20170 (N_20170,N_19204,N_19593);
and U20171 (N_20171,N_19980,N_18784);
or U20172 (N_20172,N_18962,N_19567);
nor U20173 (N_20173,N_19586,N_18851);
nor U20174 (N_20174,N_19687,N_19734);
xor U20175 (N_20175,N_19193,N_19933);
nor U20176 (N_20176,N_18932,N_19153);
and U20177 (N_20177,N_19152,N_19132);
nor U20178 (N_20178,N_19701,N_19929);
nor U20179 (N_20179,N_19969,N_19186);
or U20180 (N_20180,N_19143,N_19045);
or U20181 (N_20181,N_18842,N_19040);
or U20182 (N_20182,N_19388,N_19426);
xor U20183 (N_20183,N_19354,N_18750);
and U20184 (N_20184,N_19428,N_19612);
xnor U20185 (N_20185,N_19887,N_19017);
nand U20186 (N_20186,N_19174,N_19906);
nor U20187 (N_20187,N_19312,N_19216);
and U20188 (N_20188,N_18975,N_19102);
or U20189 (N_20189,N_18775,N_19578);
nand U20190 (N_20190,N_19306,N_19098);
and U20191 (N_20191,N_19961,N_19865);
and U20192 (N_20192,N_19144,N_19742);
nor U20193 (N_20193,N_18953,N_19942);
or U20194 (N_20194,N_18939,N_19026);
nand U20195 (N_20195,N_18798,N_19511);
nand U20196 (N_20196,N_18824,N_19247);
nor U20197 (N_20197,N_19627,N_19219);
xnor U20198 (N_20198,N_19535,N_18773);
nor U20199 (N_20199,N_19207,N_18863);
xnor U20200 (N_20200,N_19250,N_19664);
nand U20201 (N_20201,N_19070,N_19305);
or U20202 (N_20202,N_19408,N_18924);
nand U20203 (N_20203,N_18905,N_18805);
nor U20204 (N_20204,N_19332,N_19778);
or U20205 (N_20205,N_19444,N_18811);
xnor U20206 (N_20206,N_19010,N_19771);
nand U20207 (N_20207,N_19107,N_19710);
nor U20208 (N_20208,N_18993,N_19817);
nand U20209 (N_20209,N_19894,N_19293);
nor U20210 (N_20210,N_19994,N_19477);
xnor U20211 (N_20211,N_19544,N_19957);
or U20212 (N_20212,N_18812,N_19838);
nor U20213 (N_20213,N_19468,N_19648);
xor U20214 (N_20214,N_19022,N_18825);
nand U20215 (N_20215,N_19093,N_19384);
and U20216 (N_20216,N_19317,N_19904);
or U20217 (N_20217,N_19359,N_19345);
or U20218 (N_20218,N_19747,N_18772);
nand U20219 (N_20219,N_18866,N_19728);
nor U20220 (N_20220,N_18966,N_19310);
xor U20221 (N_20221,N_19936,N_19081);
or U20222 (N_20222,N_18759,N_19705);
and U20223 (N_20223,N_19407,N_19085);
xnor U20224 (N_20224,N_19065,N_19967);
xor U20225 (N_20225,N_19403,N_19913);
nand U20226 (N_20226,N_19088,N_18808);
nor U20227 (N_20227,N_19103,N_19608);
nor U20228 (N_20228,N_19741,N_19386);
nor U20229 (N_20229,N_19420,N_19034);
nor U20230 (N_20230,N_19371,N_19479);
nand U20231 (N_20231,N_19580,N_19520);
and U20232 (N_20232,N_18849,N_18942);
and U20233 (N_20233,N_19981,N_19287);
xnor U20234 (N_20234,N_19430,N_19454);
xor U20235 (N_20235,N_19720,N_19393);
xor U20236 (N_20236,N_19753,N_19094);
xnor U20237 (N_20237,N_19773,N_19389);
or U20238 (N_20238,N_18766,N_19124);
or U20239 (N_20239,N_19108,N_19133);
or U20240 (N_20240,N_19521,N_19467);
and U20241 (N_20241,N_19258,N_18829);
nand U20242 (N_20242,N_18950,N_19160);
nor U20243 (N_20243,N_18938,N_19368);
nor U20244 (N_20244,N_18807,N_18778);
nor U20245 (N_20245,N_19830,N_19955);
xor U20246 (N_20246,N_18990,N_19683);
nand U20247 (N_20247,N_19947,N_19524);
nor U20248 (N_20248,N_19438,N_19418);
nor U20249 (N_20249,N_19330,N_19768);
and U20250 (N_20250,N_19825,N_19311);
or U20251 (N_20251,N_19329,N_19999);
or U20252 (N_20252,N_18934,N_19946);
or U20253 (N_20253,N_19624,N_19926);
xnor U20254 (N_20254,N_18952,N_19381);
nand U20255 (N_20255,N_19984,N_19978);
nand U20256 (N_20256,N_19824,N_19039);
or U20257 (N_20257,N_19537,N_18958);
nor U20258 (N_20258,N_18877,N_19804);
xnor U20259 (N_20259,N_18997,N_19826);
or U20260 (N_20260,N_19661,N_19644);
or U20261 (N_20261,N_19610,N_19668);
xnor U20262 (N_20262,N_19167,N_19677);
and U20263 (N_20263,N_19658,N_19573);
xnor U20264 (N_20264,N_19351,N_18848);
nor U20265 (N_20265,N_19973,N_19726);
nor U20266 (N_20266,N_19432,N_18978);
and U20267 (N_20267,N_19058,N_19764);
and U20268 (N_20268,N_19814,N_19199);
or U20269 (N_20269,N_18846,N_18781);
nor U20270 (N_20270,N_19464,N_19788);
nor U20271 (N_20271,N_19775,N_18865);
nand U20272 (N_20272,N_19729,N_19767);
xor U20273 (N_20273,N_19372,N_18876);
or U20274 (N_20274,N_19577,N_19822);
and U20275 (N_20275,N_19650,N_19079);
xor U20276 (N_20276,N_19795,N_19169);
xor U20277 (N_20277,N_19750,N_19869);
or U20278 (N_20278,N_19390,N_19013);
nand U20279 (N_20279,N_19676,N_18918);
xor U20280 (N_20280,N_18874,N_19452);
or U20281 (N_20281,N_18910,N_19053);
xnor U20282 (N_20282,N_19012,N_19530);
xor U20283 (N_20283,N_19069,N_19555);
nand U20284 (N_20284,N_19666,N_19745);
and U20285 (N_20285,N_18816,N_19131);
xor U20286 (N_20286,N_19551,N_19785);
and U20287 (N_20287,N_19949,N_19527);
nor U20288 (N_20288,N_18774,N_19008);
xnor U20289 (N_20289,N_18912,N_19394);
nand U20290 (N_20290,N_18944,N_19170);
nand U20291 (N_20291,N_18847,N_19128);
nand U20292 (N_20292,N_19319,N_19811);
xnor U20293 (N_20293,N_19787,N_19086);
nand U20294 (N_20294,N_19684,N_19528);
and U20295 (N_20295,N_18861,N_19410);
and U20296 (N_20296,N_19248,N_19222);
nor U20297 (N_20297,N_19582,N_19862);
nor U20298 (N_20298,N_18937,N_19755);
nand U20299 (N_20299,N_19252,N_19669);
or U20300 (N_20300,N_19997,N_18792);
nand U20301 (N_20301,N_18900,N_18753);
xnor U20302 (N_20302,N_19900,N_19841);
and U20303 (N_20303,N_19839,N_18971);
or U20304 (N_20304,N_19374,N_19866);
or U20305 (N_20305,N_19935,N_19941);
nor U20306 (N_20306,N_19522,N_19801);
nor U20307 (N_20307,N_18803,N_19954);
or U20308 (N_20308,N_18765,N_19781);
or U20309 (N_20309,N_18989,N_19235);
nor U20310 (N_20310,N_19177,N_19590);
nand U20311 (N_20311,N_19592,N_19154);
nor U20312 (N_20312,N_19320,N_19607);
or U20313 (N_20313,N_19721,N_18935);
and U20314 (N_20314,N_19233,N_19043);
and U20315 (N_20315,N_18814,N_19482);
xnor U20316 (N_20316,N_19264,N_19812);
nand U20317 (N_20317,N_18907,N_19047);
or U20318 (N_20318,N_18813,N_19921);
or U20319 (N_20319,N_18823,N_19618);
xor U20320 (N_20320,N_19502,N_19800);
nand U20321 (N_20321,N_19995,N_19007);
or U20322 (N_20322,N_18919,N_18799);
nand U20323 (N_20323,N_19654,N_18955);
nand U20324 (N_20324,N_18929,N_19892);
nor U20325 (N_20325,N_19000,N_19285);
nor U20326 (N_20326,N_19437,N_19883);
and U20327 (N_20327,N_18948,N_19376);
nand U20328 (N_20328,N_19503,N_19457);
nor U20329 (N_20329,N_19633,N_19123);
xnor U20330 (N_20330,N_19321,N_18841);
nor U20331 (N_20331,N_19244,N_19031);
xor U20332 (N_20332,N_19696,N_19819);
and U20333 (N_20333,N_19362,N_19028);
nand U20334 (N_20334,N_19125,N_19492);
nand U20335 (N_20335,N_18913,N_19515);
or U20336 (N_20336,N_19375,N_19080);
nor U20337 (N_20337,N_19735,N_19016);
and U20338 (N_20338,N_19952,N_18992);
xnor U20339 (N_20339,N_19114,N_19972);
and U20340 (N_20340,N_19908,N_19693);
nand U20341 (N_20341,N_19917,N_19379);
nor U20342 (N_20342,N_19754,N_19171);
nor U20343 (N_20343,N_19400,N_19096);
nand U20344 (N_20344,N_19275,N_19163);
xor U20345 (N_20345,N_19643,N_19968);
and U20346 (N_20346,N_19557,N_19889);
or U20347 (N_20347,N_19162,N_19784);
nand U20348 (N_20348,N_19996,N_19462);
xor U20349 (N_20349,N_18843,N_19870);
and U20350 (N_20350,N_19542,N_19843);
nand U20351 (N_20351,N_19717,N_19399);
xor U20352 (N_20352,N_18872,N_18820);
xnor U20353 (N_20353,N_18909,N_19625);
xnor U20354 (N_20354,N_18893,N_18940);
nand U20355 (N_20355,N_18898,N_19173);
xnor U20356 (N_20356,N_19548,N_18838);
nor U20357 (N_20357,N_19875,N_19790);
and U20358 (N_20358,N_19660,N_19837);
nand U20359 (N_20359,N_18835,N_18762);
nand U20360 (N_20360,N_19719,N_19657);
xor U20361 (N_20361,N_19422,N_18802);
nand U20362 (N_20362,N_19019,N_19190);
nand U20363 (N_20363,N_19682,N_18862);
xnor U20364 (N_20364,N_19155,N_19201);
or U20365 (N_20365,N_19960,N_18985);
and U20366 (N_20366,N_19156,N_19042);
nor U20367 (N_20367,N_19533,N_19525);
and U20368 (N_20368,N_19993,N_19267);
or U20369 (N_20369,N_19315,N_19366);
and U20370 (N_20370,N_18791,N_19052);
nor U20371 (N_20371,N_18794,N_19129);
xnor U20372 (N_20372,N_19082,N_19148);
or U20373 (N_20373,N_19290,N_18764);
or U20374 (N_20374,N_19891,N_18991);
xnor U20375 (N_20375,N_19667,N_18961);
or U20376 (N_20376,N_19062,N_19363);
nand U20377 (N_20377,N_19262,N_19763);
xor U20378 (N_20378,N_19446,N_18998);
and U20379 (N_20379,N_19974,N_19313);
nor U20380 (N_20380,N_19066,N_19111);
nand U20381 (N_20381,N_19576,N_19637);
and U20382 (N_20382,N_19571,N_18923);
or U20383 (N_20383,N_18752,N_18965);
xor U20384 (N_20384,N_18982,N_19411);
nand U20385 (N_20385,N_19035,N_19909);
or U20386 (N_20386,N_19325,N_19833);
nor U20387 (N_20387,N_18867,N_19918);
and U20388 (N_20388,N_19796,N_19113);
nor U20389 (N_20389,N_19766,N_19493);
nor U20390 (N_20390,N_19546,N_19230);
nand U20391 (N_20391,N_19938,N_19581);
xnor U20392 (N_20392,N_19789,N_19044);
xnor U20393 (N_20393,N_19678,N_19561);
nor U20394 (N_20394,N_19985,N_19135);
nand U20395 (N_20395,N_19165,N_19090);
nand U20396 (N_20396,N_18770,N_19087);
nor U20397 (N_20397,N_18763,N_19269);
nand U20398 (N_20398,N_19736,N_19760);
nand U20399 (N_20399,N_19436,N_19626);
nand U20400 (N_20400,N_19634,N_19089);
and U20401 (N_20401,N_19360,N_18839);
or U20402 (N_20402,N_19015,N_19018);
xor U20403 (N_20403,N_18896,N_19198);
or U20404 (N_20404,N_19348,N_19964);
or U20405 (N_20405,N_19622,N_19397);
nand U20406 (N_20406,N_18875,N_19091);
nor U20407 (N_20407,N_19324,N_19902);
nor U20408 (N_20408,N_19335,N_19509);
xnor U20409 (N_20409,N_18957,N_19353);
or U20410 (N_20410,N_19037,N_19656);
or U20411 (N_20411,N_19583,N_19655);
nand U20412 (N_20412,N_19642,N_19117);
nor U20413 (N_20413,N_19011,N_19748);
or U20414 (N_20414,N_19398,N_19782);
nand U20415 (N_20415,N_19343,N_19023);
and U20416 (N_20416,N_19792,N_19970);
and U20417 (N_20417,N_19699,N_19456);
nor U20418 (N_20418,N_19873,N_19212);
nor U20419 (N_20419,N_19097,N_19568);
nor U20420 (N_20420,N_19118,N_19380);
nor U20421 (N_20421,N_19112,N_19073);
nand U20422 (N_20422,N_19615,N_19068);
nor U20423 (N_20423,N_19821,N_18996);
and U20424 (N_20424,N_18972,N_18928);
nor U20425 (N_20425,N_19500,N_19029);
nor U20426 (N_20426,N_19496,N_19099);
nor U20427 (N_20427,N_19453,N_19488);
and U20428 (N_20428,N_19638,N_19448);
xnor U20429 (N_20429,N_19730,N_18870);
or U20430 (N_20430,N_19145,N_19558);
nor U20431 (N_20431,N_19944,N_19574);
xor U20432 (N_20432,N_19038,N_18967);
nand U20433 (N_20433,N_19844,N_19342);
or U20434 (N_20434,N_18949,N_18854);
nand U20435 (N_20435,N_18787,N_18984);
and U20436 (N_20436,N_18853,N_19497);
xor U20437 (N_20437,N_19347,N_19966);
nand U20438 (N_20438,N_19278,N_19518);
xor U20439 (N_20439,N_19939,N_19141);
nor U20440 (N_20440,N_19805,N_19469);
and U20441 (N_20441,N_18809,N_18757);
nand U20442 (N_20442,N_19876,N_19934);
xnor U20443 (N_20443,N_18964,N_19054);
and U20444 (N_20444,N_19475,N_19601);
nand U20445 (N_20445,N_19898,N_19589);
nand U20446 (N_20446,N_19649,N_19120);
and U20447 (N_20447,N_18761,N_19543);
nand U20448 (N_20448,N_18754,N_19779);
or U20449 (N_20449,N_19998,N_19554);
nor U20450 (N_20450,N_19241,N_18922);
xnor U20451 (N_20451,N_19218,N_19191);
and U20452 (N_20452,N_19619,N_19200);
xnor U20453 (N_20453,N_19147,N_19232);
or U20454 (N_20454,N_18886,N_19886);
nand U20455 (N_20455,N_19006,N_19850);
or U20456 (N_20456,N_19030,N_19989);
xnor U20457 (N_20457,N_18806,N_18830);
nor U20458 (N_20458,N_19341,N_19681);
nand U20459 (N_20459,N_19159,N_19300);
and U20460 (N_20460,N_19243,N_19369);
nor U20461 (N_20461,N_19919,N_19549);
and U20462 (N_20462,N_19227,N_18826);
nor U20463 (N_20463,N_19429,N_19225);
nor U20464 (N_20464,N_19401,N_19256);
or U20465 (N_20465,N_19621,N_19486);
xnor U20466 (N_20466,N_19142,N_19032);
or U20467 (N_20467,N_18850,N_19808);
nor U20468 (N_20468,N_19922,N_19333);
nand U20469 (N_20469,N_19277,N_19302);
xor U20470 (N_20470,N_18780,N_19924);
nand U20471 (N_20471,N_18917,N_19871);
nor U20472 (N_20472,N_19772,N_19283);
xor U20473 (N_20473,N_19358,N_18980);
and U20474 (N_20474,N_18894,N_19565);
nor U20475 (N_20475,N_19539,N_19879);
and U20476 (N_20476,N_18797,N_19425);
nor U20477 (N_20477,N_18859,N_19339);
or U20478 (N_20478,N_19209,N_19823);
nor U20479 (N_20479,N_19672,N_19261);
and U20480 (N_20480,N_19059,N_19195);
xor U20481 (N_20481,N_18915,N_18834);
xnor U20482 (N_20482,N_19255,N_19274);
xnor U20483 (N_20483,N_19807,N_19845);
xnor U20484 (N_20484,N_19415,N_19140);
and U20485 (N_20485,N_19308,N_19594);
nand U20486 (N_20486,N_19912,N_19223);
and U20487 (N_20487,N_19538,N_19727);
nand U20488 (N_20488,N_19636,N_18904);
and U20489 (N_20489,N_19884,N_19078);
and U20490 (N_20490,N_19272,N_19164);
and U20491 (N_20491,N_19352,N_18936);
and U20492 (N_20492,N_18760,N_18871);
xor U20493 (N_20493,N_18883,N_19749);
and U20494 (N_20494,N_19254,N_18920);
or U20495 (N_20495,N_19579,N_18800);
and U20496 (N_20496,N_19945,N_19890);
or U20497 (N_20497,N_19540,N_19617);
and U20498 (N_20498,N_19297,N_19630);
nor U20499 (N_20499,N_18844,N_19396);
nand U20500 (N_20500,N_19910,N_18956);
nand U20501 (N_20501,N_19136,N_19063);
nand U20502 (N_20502,N_19856,N_19104);
and U20503 (N_20503,N_19604,N_19975);
nor U20504 (N_20504,N_19176,N_19663);
and U20505 (N_20505,N_19536,N_19599);
nand U20506 (N_20506,N_19072,N_19427);
nand U20507 (N_20507,N_18941,N_19158);
nor U20508 (N_20508,N_19953,N_19231);
nor U20509 (N_20509,N_19182,N_19056);
or U20510 (N_20510,N_19857,N_19971);
xor U20511 (N_20511,N_19616,N_19956);
xor U20512 (N_20512,N_18815,N_19963);
nand U20513 (N_20513,N_19213,N_18931);
xor U20514 (N_20514,N_18911,N_19690);
and U20515 (N_20515,N_19545,N_19494);
and U20516 (N_20516,N_19279,N_19027);
nand U20517 (N_20517,N_19834,N_19004);
nand U20518 (N_20518,N_19122,N_19292);
or U20519 (N_20519,N_19138,N_19510);
or U20520 (N_20520,N_19798,N_19740);
xnor U20521 (N_20521,N_19797,N_19282);
nand U20522 (N_20522,N_19307,N_19435);
and U20523 (N_20523,N_19711,N_19116);
and U20524 (N_20524,N_19309,N_19507);
or U20525 (N_20525,N_19378,N_19541);
or U20526 (N_20526,N_19490,N_18804);
or U20527 (N_20527,N_19344,N_19121);
or U20528 (N_20528,N_19670,N_19387);
and U20529 (N_20529,N_19413,N_19882);
nor U20530 (N_20530,N_19025,N_19802);
xor U20531 (N_20531,N_19990,N_19793);
nor U20532 (N_20532,N_19928,N_19458);
or U20533 (N_20533,N_19385,N_19631);
nand U20534 (N_20534,N_19780,N_19449);
nor U20535 (N_20535,N_18855,N_19846);
xnor U20536 (N_20536,N_19559,N_19716);
xor U20537 (N_20537,N_19180,N_19598);
nor U20538 (N_20538,N_19595,N_19700);
or U20539 (N_20539,N_19547,N_19671);
and U20540 (N_20540,N_19992,N_18793);
xor U20541 (N_20541,N_19280,N_19289);
or U20542 (N_20542,N_19885,N_19357);
nor U20543 (N_20543,N_19101,N_19473);
and U20544 (N_20544,N_18769,N_19455);
nand U20545 (N_20545,N_18916,N_19809);
or U20546 (N_20546,N_19514,N_19659);
xor U20547 (N_20547,N_19433,N_19476);
and U20548 (N_20548,N_19635,N_19878);
nor U20549 (N_20549,N_18946,N_19228);
or U20550 (N_20550,N_19259,N_18819);
or U20551 (N_20551,N_18960,N_18930);
or U20552 (N_20552,N_18821,N_19051);
nand U20553 (N_20553,N_19327,N_19005);
and U20554 (N_20554,N_19874,N_19905);
and U20555 (N_20555,N_18783,N_19095);
nor U20556 (N_20556,N_19041,N_19105);
or U20557 (N_20557,N_18860,N_19431);
nand U20558 (N_20558,N_19465,N_19301);
and U20559 (N_20559,N_19888,N_19161);
nor U20560 (N_20560,N_19762,N_19245);
and U20561 (N_20561,N_19722,N_19709);
and U20562 (N_20562,N_19229,N_19697);
nand U20563 (N_20563,N_18869,N_18782);
nor U20564 (N_20564,N_18903,N_18906);
or U20565 (N_20565,N_19940,N_18810);
xnor U20566 (N_20566,N_19951,N_19471);
xnor U20567 (N_20567,N_19847,N_19842);
or U20568 (N_20568,N_19485,N_19498);
xnor U20569 (N_20569,N_18878,N_18789);
xnor U20570 (N_20570,N_18801,N_19774);
or U20571 (N_20571,N_19036,N_19703);
nor U20572 (N_20572,N_19046,N_19513);
or U20573 (N_20573,N_19983,N_19001);
nand U20574 (N_20574,N_19786,N_18881);
and U20575 (N_20575,N_18779,N_18879);
and U20576 (N_20576,N_19487,N_18868);
nor U20577 (N_20577,N_18858,N_19373);
nand U20578 (N_20578,N_19187,N_19459);
xor U20579 (N_20579,N_19758,N_19461);
nand U20580 (N_20580,N_19478,N_19662);
nand U20581 (N_20581,N_18864,N_19451);
or U20582 (N_20582,N_19406,N_19349);
or U20583 (N_20583,N_18882,N_18852);
xnor U20584 (N_20584,N_19609,N_19930);
or U20585 (N_20585,N_19907,N_19483);
xnor U20586 (N_20586,N_19328,N_18885);
or U20587 (N_20587,N_19139,N_19896);
xor U20588 (N_20588,N_19024,N_19049);
nand U20589 (N_20589,N_19564,N_18856);
or U20590 (N_20590,N_19570,N_18840);
and U20591 (N_20591,N_19202,N_19074);
nor U20592 (N_20592,N_19602,N_19084);
nand U20593 (N_20593,N_19673,N_19692);
and U20594 (N_20594,N_19508,N_19647);
xnor U20595 (N_20595,N_19688,N_19355);
xnor U20596 (N_20596,N_19806,N_19203);
or U20597 (N_20597,N_19130,N_19706);
nor U20598 (N_20598,N_18758,N_19738);
nor U20599 (N_20599,N_19192,N_19959);
nand U20600 (N_20600,N_19240,N_19744);
or U20601 (N_20601,N_18873,N_19853);
and U20602 (N_20602,N_19620,N_19903);
nand U20603 (N_20603,N_19364,N_19450);
or U20604 (N_20604,N_19733,N_18751);
and U20605 (N_20605,N_19217,N_19702);
nor U20606 (N_20606,N_18947,N_19392);
nand U20607 (N_20607,N_19832,N_19350);
or U20608 (N_20608,N_19783,N_19134);
or U20609 (N_20609,N_19055,N_19757);
and U20610 (N_20610,N_18891,N_18943);
nor U20611 (N_20611,N_19752,N_19813);
xor U20612 (N_20612,N_19820,N_19563);
nand U20613 (N_20613,N_19818,N_19723);
or U20614 (N_20614,N_19246,N_19484);
xnor U20615 (N_20615,N_19712,N_19512);
or U20616 (N_20616,N_19268,N_19816);
or U20617 (N_20617,N_19370,N_19076);
or U20618 (N_20618,N_19665,N_19743);
nand U20619 (N_20619,N_19517,N_19014);
nand U20620 (N_20620,N_19208,N_19976);
nand U20621 (N_20621,N_19725,N_19434);
and U20622 (N_20622,N_19196,N_19137);
xor U20623 (N_20623,N_18889,N_19639);
xnor U20624 (N_20624,N_18892,N_18833);
or U20625 (N_20625,N_19664,N_19966);
or U20626 (N_20626,N_19886,N_19480);
and U20627 (N_20627,N_19812,N_19572);
nor U20628 (N_20628,N_19222,N_19179);
nand U20629 (N_20629,N_18850,N_19249);
and U20630 (N_20630,N_19384,N_19860);
xor U20631 (N_20631,N_19148,N_19842);
nand U20632 (N_20632,N_19231,N_18756);
or U20633 (N_20633,N_19273,N_19810);
nor U20634 (N_20634,N_18878,N_19018);
xor U20635 (N_20635,N_19954,N_19574);
and U20636 (N_20636,N_19849,N_19546);
and U20637 (N_20637,N_19021,N_19862);
or U20638 (N_20638,N_18998,N_19167);
nor U20639 (N_20639,N_19783,N_19778);
nand U20640 (N_20640,N_19779,N_19255);
xnor U20641 (N_20641,N_19936,N_19370);
and U20642 (N_20642,N_18797,N_18977);
nor U20643 (N_20643,N_19014,N_19091);
xor U20644 (N_20644,N_19134,N_19650);
xor U20645 (N_20645,N_19155,N_19934);
nand U20646 (N_20646,N_19556,N_19986);
nor U20647 (N_20647,N_19026,N_18834);
or U20648 (N_20648,N_19871,N_19522);
or U20649 (N_20649,N_18994,N_19540);
nor U20650 (N_20650,N_19285,N_19052);
nand U20651 (N_20651,N_19042,N_19304);
xor U20652 (N_20652,N_19636,N_19550);
xor U20653 (N_20653,N_19559,N_18761);
or U20654 (N_20654,N_19359,N_19136);
or U20655 (N_20655,N_19309,N_19999);
nand U20656 (N_20656,N_19221,N_19169);
or U20657 (N_20657,N_19519,N_19029);
or U20658 (N_20658,N_19018,N_19171);
xnor U20659 (N_20659,N_19646,N_19719);
or U20660 (N_20660,N_19644,N_19786);
nand U20661 (N_20661,N_18835,N_19862);
or U20662 (N_20662,N_19198,N_19692);
or U20663 (N_20663,N_18756,N_19294);
or U20664 (N_20664,N_19488,N_19662);
nor U20665 (N_20665,N_18882,N_19294);
and U20666 (N_20666,N_19972,N_18755);
xor U20667 (N_20667,N_19953,N_18797);
and U20668 (N_20668,N_19360,N_19561);
or U20669 (N_20669,N_19454,N_18983);
nor U20670 (N_20670,N_19488,N_19812);
nor U20671 (N_20671,N_18965,N_19989);
nand U20672 (N_20672,N_19436,N_19258);
xor U20673 (N_20673,N_19577,N_19640);
nand U20674 (N_20674,N_19044,N_19309);
nor U20675 (N_20675,N_19529,N_19672);
or U20676 (N_20676,N_19562,N_18925);
or U20677 (N_20677,N_19673,N_19956);
nor U20678 (N_20678,N_19898,N_19466);
or U20679 (N_20679,N_18763,N_19537);
nand U20680 (N_20680,N_19638,N_19514);
and U20681 (N_20681,N_19583,N_19054);
and U20682 (N_20682,N_19812,N_19070);
nor U20683 (N_20683,N_19726,N_18915);
or U20684 (N_20684,N_18753,N_19698);
or U20685 (N_20685,N_18805,N_19798);
nand U20686 (N_20686,N_19788,N_19254);
nand U20687 (N_20687,N_19756,N_18780);
or U20688 (N_20688,N_19500,N_19940);
and U20689 (N_20689,N_19591,N_19334);
nor U20690 (N_20690,N_19143,N_19411);
or U20691 (N_20691,N_18784,N_18810);
or U20692 (N_20692,N_18885,N_19546);
xor U20693 (N_20693,N_19366,N_18834);
or U20694 (N_20694,N_19579,N_19213);
xor U20695 (N_20695,N_19678,N_19484);
xor U20696 (N_20696,N_19517,N_19663);
nor U20697 (N_20697,N_19899,N_19471);
nor U20698 (N_20698,N_19688,N_19463);
or U20699 (N_20699,N_19999,N_18937);
or U20700 (N_20700,N_19262,N_19961);
nor U20701 (N_20701,N_19684,N_19112);
xnor U20702 (N_20702,N_19561,N_19881);
nor U20703 (N_20703,N_19888,N_19890);
nand U20704 (N_20704,N_19009,N_19583);
xor U20705 (N_20705,N_19019,N_19024);
and U20706 (N_20706,N_19815,N_19135);
or U20707 (N_20707,N_18875,N_19724);
nand U20708 (N_20708,N_19372,N_19482);
or U20709 (N_20709,N_19172,N_19464);
nand U20710 (N_20710,N_18819,N_19784);
xor U20711 (N_20711,N_18757,N_18898);
or U20712 (N_20712,N_19609,N_19440);
or U20713 (N_20713,N_19169,N_19302);
nor U20714 (N_20714,N_19785,N_19693);
or U20715 (N_20715,N_19769,N_19802);
nand U20716 (N_20716,N_19910,N_19510);
or U20717 (N_20717,N_18996,N_18826);
and U20718 (N_20718,N_19097,N_19215);
nor U20719 (N_20719,N_18886,N_19903);
or U20720 (N_20720,N_19335,N_18794);
nor U20721 (N_20721,N_19283,N_19497);
or U20722 (N_20722,N_19909,N_18773);
xnor U20723 (N_20723,N_19868,N_19576);
nand U20724 (N_20724,N_19686,N_18902);
and U20725 (N_20725,N_19403,N_19683);
xor U20726 (N_20726,N_19999,N_19269);
and U20727 (N_20727,N_19885,N_19019);
nor U20728 (N_20728,N_19617,N_19187);
and U20729 (N_20729,N_18998,N_19288);
nor U20730 (N_20730,N_18818,N_19775);
xor U20731 (N_20731,N_19010,N_19945);
nand U20732 (N_20732,N_19981,N_18974);
and U20733 (N_20733,N_19332,N_19750);
and U20734 (N_20734,N_19867,N_19679);
and U20735 (N_20735,N_19655,N_19206);
nand U20736 (N_20736,N_18861,N_19558);
or U20737 (N_20737,N_19103,N_19303);
and U20738 (N_20738,N_18969,N_18891);
or U20739 (N_20739,N_19358,N_19230);
or U20740 (N_20740,N_18756,N_19483);
or U20741 (N_20741,N_19341,N_19394);
xnor U20742 (N_20742,N_19184,N_19517);
and U20743 (N_20743,N_19258,N_19748);
or U20744 (N_20744,N_19920,N_19452);
xnor U20745 (N_20745,N_19785,N_19601);
or U20746 (N_20746,N_19922,N_19322);
and U20747 (N_20747,N_19461,N_19201);
xnor U20748 (N_20748,N_19118,N_19454);
nor U20749 (N_20749,N_19979,N_19552);
nand U20750 (N_20750,N_19070,N_19017);
nor U20751 (N_20751,N_18764,N_19633);
nand U20752 (N_20752,N_19976,N_19059);
nor U20753 (N_20753,N_18906,N_19159);
nand U20754 (N_20754,N_19261,N_19689);
nand U20755 (N_20755,N_19476,N_19942);
or U20756 (N_20756,N_18873,N_19751);
and U20757 (N_20757,N_19223,N_18874);
xor U20758 (N_20758,N_19474,N_19142);
and U20759 (N_20759,N_19174,N_19414);
xnor U20760 (N_20760,N_19067,N_19817);
and U20761 (N_20761,N_19880,N_18828);
xor U20762 (N_20762,N_18887,N_19764);
nor U20763 (N_20763,N_19612,N_19100);
or U20764 (N_20764,N_18992,N_19363);
nand U20765 (N_20765,N_19603,N_19390);
or U20766 (N_20766,N_19793,N_18804);
and U20767 (N_20767,N_19277,N_18949);
or U20768 (N_20768,N_18952,N_19362);
and U20769 (N_20769,N_19205,N_19625);
nor U20770 (N_20770,N_19946,N_19124);
or U20771 (N_20771,N_19833,N_19533);
xnor U20772 (N_20772,N_19056,N_19457);
and U20773 (N_20773,N_19557,N_19318);
nor U20774 (N_20774,N_19547,N_19388);
xor U20775 (N_20775,N_19175,N_19568);
nand U20776 (N_20776,N_19208,N_19482);
xor U20777 (N_20777,N_19233,N_19321);
nor U20778 (N_20778,N_19234,N_19324);
xor U20779 (N_20779,N_19327,N_19925);
nand U20780 (N_20780,N_18898,N_19610);
and U20781 (N_20781,N_18934,N_19733);
nor U20782 (N_20782,N_19729,N_18882);
nor U20783 (N_20783,N_19098,N_19115);
nor U20784 (N_20784,N_19213,N_19262);
and U20785 (N_20785,N_19395,N_19968);
nor U20786 (N_20786,N_19628,N_19747);
nor U20787 (N_20787,N_19356,N_19593);
xnor U20788 (N_20788,N_19072,N_19062);
nand U20789 (N_20789,N_18971,N_19121);
nand U20790 (N_20790,N_19207,N_19326);
xnor U20791 (N_20791,N_18901,N_18792);
nand U20792 (N_20792,N_19399,N_19561);
xnor U20793 (N_20793,N_18752,N_19635);
xnor U20794 (N_20794,N_19379,N_19843);
nand U20795 (N_20795,N_19484,N_19347);
or U20796 (N_20796,N_19390,N_18923);
and U20797 (N_20797,N_18995,N_19261);
nor U20798 (N_20798,N_19072,N_19484);
nor U20799 (N_20799,N_19314,N_19623);
xor U20800 (N_20800,N_19189,N_18808);
or U20801 (N_20801,N_19609,N_18759);
xnor U20802 (N_20802,N_18897,N_18832);
or U20803 (N_20803,N_19117,N_19111);
or U20804 (N_20804,N_19563,N_18776);
nor U20805 (N_20805,N_19919,N_19682);
or U20806 (N_20806,N_19620,N_19533);
xnor U20807 (N_20807,N_19059,N_19961);
xnor U20808 (N_20808,N_19134,N_19202);
xnor U20809 (N_20809,N_19946,N_19293);
nand U20810 (N_20810,N_19960,N_19634);
nor U20811 (N_20811,N_19854,N_19365);
and U20812 (N_20812,N_19622,N_19403);
nor U20813 (N_20813,N_19991,N_19971);
xnor U20814 (N_20814,N_19246,N_19314);
xor U20815 (N_20815,N_19802,N_19497);
and U20816 (N_20816,N_19665,N_19267);
xnor U20817 (N_20817,N_19702,N_19771);
nor U20818 (N_20818,N_18935,N_19247);
nor U20819 (N_20819,N_19356,N_19341);
nand U20820 (N_20820,N_18951,N_18881);
nand U20821 (N_20821,N_19456,N_19436);
nor U20822 (N_20822,N_19448,N_19975);
and U20823 (N_20823,N_19516,N_19170);
nand U20824 (N_20824,N_18950,N_18844);
xor U20825 (N_20825,N_19737,N_19990);
or U20826 (N_20826,N_19695,N_19030);
nor U20827 (N_20827,N_19302,N_19988);
or U20828 (N_20828,N_19664,N_19783);
nor U20829 (N_20829,N_18967,N_18754);
nand U20830 (N_20830,N_19490,N_19661);
nor U20831 (N_20831,N_18901,N_19282);
nor U20832 (N_20832,N_19977,N_19646);
nor U20833 (N_20833,N_19915,N_19125);
and U20834 (N_20834,N_19862,N_19583);
nand U20835 (N_20835,N_19607,N_19147);
and U20836 (N_20836,N_19597,N_19086);
or U20837 (N_20837,N_19470,N_19145);
xor U20838 (N_20838,N_18786,N_19772);
xor U20839 (N_20839,N_19893,N_18907);
or U20840 (N_20840,N_19779,N_19552);
or U20841 (N_20841,N_19887,N_19710);
or U20842 (N_20842,N_19921,N_19672);
and U20843 (N_20843,N_18894,N_19202);
or U20844 (N_20844,N_19291,N_19505);
and U20845 (N_20845,N_18995,N_18859);
nand U20846 (N_20846,N_18840,N_19124);
or U20847 (N_20847,N_19753,N_19719);
xor U20848 (N_20848,N_19039,N_19330);
nand U20849 (N_20849,N_18873,N_19603);
and U20850 (N_20850,N_19029,N_19719);
nand U20851 (N_20851,N_19709,N_19401);
nor U20852 (N_20852,N_19668,N_18789);
nand U20853 (N_20853,N_19573,N_19271);
or U20854 (N_20854,N_19712,N_19304);
and U20855 (N_20855,N_19024,N_19452);
or U20856 (N_20856,N_19450,N_19182);
xor U20857 (N_20857,N_19274,N_19786);
and U20858 (N_20858,N_19648,N_18985);
nand U20859 (N_20859,N_19633,N_19535);
xnor U20860 (N_20860,N_19743,N_19233);
xnor U20861 (N_20861,N_19342,N_18907);
nor U20862 (N_20862,N_18976,N_18790);
nand U20863 (N_20863,N_19901,N_19370);
xnor U20864 (N_20864,N_19306,N_18754);
or U20865 (N_20865,N_19334,N_19498);
xor U20866 (N_20866,N_19570,N_18978);
or U20867 (N_20867,N_19814,N_18762);
nand U20868 (N_20868,N_18956,N_19088);
nand U20869 (N_20869,N_19075,N_18784);
and U20870 (N_20870,N_18842,N_19490);
nand U20871 (N_20871,N_19417,N_19644);
and U20872 (N_20872,N_18825,N_18911);
nor U20873 (N_20873,N_19655,N_19979);
nor U20874 (N_20874,N_18951,N_19283);
nor U20875 (N_20875,N_19619,N_19855);
xor U20876 (N_20876,N_19079,N_19923);
nor U20877 (N_20877,N_19987,N_19777);
nor U20878 (N_20878,N_19528,N_19546);
xnor U20879 (N_20879,N_19035,N_19207);
xnor U20880 (N_20880,N_19361,N_18804);
xnor U20881 (N_20881,N_19719,N_19071);
nand U20882 (N_20882,N_19646,N_19937);
nand U20883 (N_20883,N_19566,N_19315);
nor U20884 (N_20884,N_19394,N_19427);
xor U20885 (N_20885,N_19391,N_19209);
xnor U20886 (N_20886,N_19364,N_18856);
nor U20887 (N_20887,N_19642,N_19735);
nor U20888 (N_20888,N_19173,N_19010);
or U20889 (N_20889,N_19968,N_19831);
and U20890 (N_20890,N_19282,N_19969);
and U20891 (N_20891,N_19986,N_19774);
nand U20892 (N_20892,N_19697,N_18843);
and U20893 (N_20893,N_19548,N_19461);
nor U20894 (N_20894,N_19118,N_18911);
xor U20895 (N_20895,N_19061,N_19454);
or U20896 (N_20896,N_19655,N_18767);
xor U20897 (N_20897,N_19730,N_19099);
nand U20898 (N_20898,N_18995,N_19439);
nor U20899 (N_20899,N_19900,N_19611);
xor U20900 (N_20900,N_18872,N_19333);
xor U20901 (N_20901,N_19833,N_19724);
nand U20902 (N_20902,N_19317,N_19149);
and U20903 (N_20903,N_19119,N_19265);
nand U20904 (N_20904,N_19986,N_19600);
nand U20905 (N_20905,N_19232,N_19242);
or U20906 (N_20906,N_19142,N_19615);
or U20907 (N_20907,N_19140,N_19221);
xnor U20908 (N_20908,N_19471,N_19514);
xnor U20909 (N_20909,N_19845,N_19371);
nand U20910 (N_20910,N_18839,N_18882);
nor U20911 (N_20911,N_18948,N_19940);
nor U20912 (N_20912,N_19400,N_19320);
nand U20913 (N_20913,N_18826,N_19869);
or U20914 (N_20914,N_19005,N_18990);
or U20915 (N_20915,N_18828,N_19606);
or U20916 (N_20916,N_19160,N_19122);
xor U20917 (N_20917,N_19969,N_19586);
xor U20918 (N_20918,N_19599,N_19907);
nand U20919 (N_20919,N_19271,N_18819);
or U20920 (N_20920,N_19928,N_19664);
and U20921 (N_20921,N_18776,N_19412);
nand U20922 (N_20922,N_19124,N_19364);
nand U20923 (N_20923,N_19936,N_19800);
or U20924 (N_20924,N_19503,N_19869);
nor U20925 (N_20925,N_19539,N_19324);
and U20926 (N_20926,N_19630,N_18925);
and U20927 (N_20927,N_19803,N_18879);
and U20928 (N_20928,N_19523,N_19140);
nor U20929 (N_20929,N_18909,N_19400);
xor U20930 (N_20930,N_19371,N_19874);
nor U20931 (N_20931,N_19370,N_19415);
and U20932 (N_20932,N_19757,N_19772);
and U20933 (N_20933,N_19258,N_19136);
xnor U20934 (N_20934,N_19372,N_19129);
xnor U20935 (N_20935,N_19352,N_18932);
or U20936 (N_20936,N_19564,N_19540);
nor U20937 (N_20937,N_19546,N_19898);
xnor U20938 (N_20938,N_19705,N_18853);
and U20939 (N_20939,N_18920,N_19449);
and U20940 (N_20940,N_19244,N_19883);
and U20941 (N_20941,N_19063,N_19749);
or U20942 (N_20942,N_19588,N_19266);
xnor U20943 (N_20943,N_19435,N_18768);
xnor U20944 (N_20944,N_19640,N_19527);
nor U20945 (N_20945,N_19207,N_18998);
or U20946 (N_20946,N_19938,N_19224);
nor U20947 (N_20947,N_19510,N_19552);
nor U20948 (N_20948,N_19501,N_18792);
nand U20949 (N_20949,N_19230,N_19026);
and U20950 (N_20950,N_19814,N_19083);
or U20951 (N_20951,N_19031,N_19896);
nand U20952 (N_20952,N_19370,N_19273);
or U20953 (N_20953,N_18833,N_18751);
xnor U20954 (N_20954,N_19987,N_19021);
or U20955 (N_20955,N_19910,N_19788);
and U20956 (N_20956,N_19940,N_19583);
nand U20957 (N_20957,N_18882,N_19212);
or U20958 (N_20958,N_19264,N_19857);
or U20959 (N_20959,N_18916,N_19248);
or U20960 (N_20960,N_19672,N_19247);
xnor U20961 (N_20961,N_18890,N_18886);
nand U20962 (N_20962,N_19933,N_18759);
and U20963 (N_20963,N_18845,N_19630);
xor U20964 (N_20964,N_19016,N_19433);
and U20965 (N_20965,N_19852,N_19345);
and U20966 (N_20966,N_19396,N_19593);
nand U20967 (N_20967,N_19322,N_19499);
xor U20968 (N_20968,N_18933,N_19840);
nand U20969 (N_20969,N_18879,N_19188);
nor U20970 (N_20970,N_18928,N_18858);
nor U20971 (N_20971,N_19977,N_19150);
nand U20972 (N_20972,N_18866,N_19127);
nor U20973 (N_20973,N_19619,N_19832);
nand U20974 (N_20974,N_19242,N_19571);
xnor U20975 (N_20975,N_19682,N_18778);
or U20976 (N_20976,N_19289,N_19129);
or U20977 (N_20977,N_19968,N_19126);
and U20978 (N_20978,N_19445,N_19349);
and U20979 (N_20979,N_18904,N_19699);
xnor U20980 (N_20980,N_19773,N_19999);
xor U20981 (N_20981,N_18899,N_18975);
nor U20982 (N_20982,N_19335,N_19146);
nor U20983 (N_20983,N_19639,N_19721);
and U20984 (N_20984,N_19094,N_19779);
nor U20985 (N_20985,N_19594,N_19532);
and U20986 (N_20986,N_19052,N_19975);
or U20987 (N_20987,N_19850,N_18922);
or U20988 (N_20988,N_18997,N_19970);
xnor U20989 (N_20989,N_18928,N_19498);
or U20990 (N_20990,N_19963,N_19867);
nand U20991 (N_20991,N_19268,N_19485);
and U20992 (N_20992,N_19649,N_19965);
xor U20993 (N_20993,N_19789,N_19199);
xnor U20994 (N_20994,N_18956,N_19422);
nor U20995 (N_20995,N_19212,N_19963);
nor U20996 (N_20996,N_19988,N_19283);
xnor U20997 (N_20997,N_19887,N_18853);
or U20998 (N_20998,N_19646,N_19636);
nand U20999 (N_20999,N_19978,N_19612);
nor U21000 (N_21000,N_19757,N_19615);
nand U21001 (N_21001,N_19270,N_19713);
or U21002 (N_21002,N_19699,N_18916);
nor U21003 (N_21003,N_19611,N_19395);
nor U21004 (N_21004,N_19216,N_19812);
nor U21005 (N_21005,N_19588,N_19003);
or U21006 (N_21006,N_19839,N_19829);
and U21007 (N_21007,N_18865,N_19722);
and U21008 (N_21008,N_18799,N_19623);
and U21009 (N_21009,N_19899,N_19747);
nor U21010 (N_21010,N_19651,N_19867);
nor U21011 (N_21011,N_19144,N_19005);
nor U21012 (N_21012,N_18782,N_19003);
xnor U21013 (N_21013,N_18810,N_18940);
xnor U21014 (N_21014,N_18931,N_19986);
or U21015 (N_21015,N_19036,N_19363);
or U21016 (N_21016,N_19124,N_19452);
nand U21017 (N_21017,N_19842,N_19977);
nor U21018 (N_21018,N_18977,N_19193);
nand U21019 (N_21019,N_18771,N_19464);
or U21020 (N_21020,N_19664,N_18885);
or U21021 (N_21021,N_19070,N_19096);
or U21022 (N_21022,N_19315,N_19915);
and U21023 (N_21023,N_19256,N_19480);
xor U21024 (N_21024,N_19975,N_18998);
or U21025 (N_21025,N_19138,N_19318);
and U21026 (N_21026,N_19441,N_19893);
nor U21027 (N_21027,N_19790,N_19837);
and U21028 (N_21028,N_19268,N_19142);
nand U21029 (N_21029,N_19567,N_19342);
xor U21030 (N_21030,N_19141,N_19311);
nand U21031 (N_21031,N_19858,N_19779);
nor U21032 (N_21032,N_19701,N_19647);
and U21033 (N_21033,N_19791,N_19529);
or U21034 (N_21034,N_19731,N_19933);
or U21035 (N_21035,N_19370,N_19534);
and U21036 (N_21036,N_19347,N_19314);
nor U21037 (N_21037,N_19238,N_19917);
nor U21038 (N_21038,N_19433,N_18865);
nand U21039 (N_21039,N_19591,N_19975);
or U21040 (N_21040,N_19309,N_19559);
and U21041 (N_21041,N_19330,N_19451);
nand U21042 (N_21042,N_19777,N_19463);
xnor U21043 (N_21043,N_19932,N_19576);
nor U21044 (N_21044,N_19252,N_19962);
nand U21045 (N_21045,N_19634,N_19449);
nand U21046 (N_21046,N_19550,N_19181);
and U21047 (N_21047,N_19203,N_19617);
xor U21048 (N_21048,N_18945,N_19408);
and U21049 (N_21049,N_19726,N_19169);
and U21050 (N_21050,N_19888,N_19410);
and U21051 (N_21051,N_19226,N_18787);
xnor U21052 (N_21052,N_18930,N_19868);
nand U21053 (N_21053,N_18793,N_18860);
nor U21054 (N_21054,N_19052,N_19946);
and U21055 (N_21055,N_19981,N_19627);
and U21056 (N_21056,N_19620,N_18767);
nand U21057 (N_21057,N_18849,N_19645);
nand U21058 (N_21058,N_18810,N_19723);
nor U21059 (N_21059,N_19016,N_19128);
and U21060 (N_21060,N_19993,N_19560);
and U21061 (N_21061,N_19282,N_19621);
and U21062 (N_21062,N_19131,N_19143);
nand U21063 (N_21063,N_18754,N_19871);
nor U21064 (N_21064,N_19772,N_19318);
or U21065 (N_21065,N_19317,N_19727);
nor U21066 (N_21066,N_19229,N_18815);
or U21067 (N_21067,N_19094,N_19185);
nand U21068 (N_21068,N_19174,N_19245);
nor U21069 (N_21069,N_19423,N_19358);
or U21070 (N_21070,N_19668,N_19399);
or U21071 (N_21071,N_19153,N_19975);
nor U21072 (N_21072,N_19511,N_19822);
nand U21073 (N_21073,N_19119,N_19689);
nor U21074 (N_21074,N_19243,N_19656);
or U21075 (N_21075,N_19711,N_19500);
xor U21076 (N_21076,N_18778,N_19628);
nor U21077 (N_21077,N_18958,N_19296);
and U21078 (N_21078,N_18899,N_19418);
xnor U21079 (N_21079,N_19326,N_18857);
and U21080 (N_21080,N_18853,N_19785);
xnor U21081 (N_21081,N_19095,N_18982);
xor U21082 (N_21082,N_19692,N_19154);
nand U21083 (N_21083,N_19105,N_19451);
or U21084 (N_21084,N_19087,N_19980);
nand U21085 (N_21085,N_19743,N_19654);
nor U21086 (N_21086,N_18893,N_19477);
or U21087 (N_21087,N_19139,N_19761);
nor U21088 (N_21088,N_19539,N_18778);
nor U21089 (N_21089,N_19512,N_19516);
or U21090 (N_21090,N_18960,N_19058);
nand U21091 (N_21091,N_19303,N_18992);
nor U21092 (N_21092,N_19009,N_19884);
or U21093 (N_21093,N_19152,N_19870);
nand U21094 (N_21094,N_19395,N_18999);
or U21095 (N_21095,N_19920,N_18857);
nand U21096 (N_21096,N_18995,N_19788);
nor U21097 (N_21097,N_18767,N_19458);
nor U21098 (N_21098,N_19220,N_19703);
and U21099 (N_21099,N_19303,N_19194);
and U21100 (N_21100,N_18829,N_18940);
nor U21101 (N_21101,N_19542,N_19487);
and U21102 (N_21102,N_18806,N_19018);
nand U21103 (N_21103,N_19620,N_18938);
nand U21104 (N_21104,N_19259,N_18779);
xnor U21105 (N_21105,N_19486,N_19915);
and U21106 (N_21106,N_19188,N_19951);
and U21107 (N_21107,N_19142,N_18902);
nand U21108 (N_21108,N_19001,N_19348);
xor U21109 (N_21109,N_19276,N_19449);
or U21110 (N_21110,N_19205,N_19612);
nand U21111 (N_21111,N_19106,N_19619);
nand U21112 (N_21112,N_19425,N_19798);
nand U21113 (N_21113,N_19282,N_19267);
nand U21114 (N_21114,N_19132,N_19860);
and U21115 (N_21115,N_18795,N_19053);
or U21116 (N_21116,N_19286,N_19671);
nand U21117 (N_21117,N_19561,N_18957);
nor U21118 (N_21118,N_19283,N_18808);
xnor U21119 (N_21119,N_19520,N_18796);
and U21120 (N_21120,N_19216,N_19928);
and U21121 (N_21121,N_19080,N_18898);
nand U21122 (N_21122,N_18862,N_19888);
and U21123 (N_21123,N_18797,N_18950);
or U21124 (N_21124,N_19425,N_19464);
xnor U21125 (N_21125,N_19173,N_18960);
xnor U21126 (N_21126,N_19490,N_19973);
or U21127 (N_21127,N_19249,N_19391);
nor U21128 (N_21128,N_19096,N_19272);
and U21129 (N_21129,N_19829,N_18975);
nor U21130 (N_21130,N_19307,N_18763);
nor U21131 (N_21131,N_19165,N_19057);
xor U21132 (N_21132,N_19288,N_19451);
and U21133 (N_21133,N_18851,N_18790);
xor U21134 (N_21134,N_19483,N_19979);
or U21135 (N_21135,N_19919,N_19629);
nand U21136 (N_21136,N_18835,N_19636);
or U21137 (N_21137,N_19875,N_19930);
nor U21138 (N_21138,N_19326,N_18971);
nor U21139 (N_21139,N_19156,N_19477);
nor U21140 (N_21140,N_19471,N_19759);
nand U21141 (N_21141,N_19303,N_19081);
nand U21142 (N_21142,N_19250,N_19985);
nor U21143 (N_21143,N_19829,N_19441);
or U21144 (N_21144,N_19241,N_19722);
xor U21145 (N_21145,N_19618,N_19869);
nor U21146 (N_21146,N_18948,N_19248);
nor U21147 (N_21147,N_19489,N_19715);
or U21148 (N_21148,N_18753,N_19390);
nor U21149 (N_21149,N_19455,N_19145);
nor U21150 (N_21150,N_19071,N_19728);
xnor U21151 (N_21151,N_19961,N_19895);
nand U21152 (N_21152,N_19634,N_19236);
nor U21153 (N_21153,N_18864,N_19158);
and U21154 (N_21154,N_19434,N_19036);
or U21155 (N_21155,N_19135,N_19324);
nand U21156 (N_21156,N_19325,N_19915);
xor U21157 (N_21157,N_19055,N_19587);
nand U21158 (N_21158,N_19649,N_19563);
xnor U21159 (N_21159,N_18833,N_19932);
nor U21160 (N_21160,N_19731,N_19090);
nor U21161 (N_21161,N_19555,N_19613);
xor U21162 (N_21162,N_19870,N_19362);
xor U21163 (N_21163,N_19919,N_18860);
xnor U21164 (N_21164,N_19531,N_19283);
or U21165 (N_21165,N_19144,N_19113);
or U21166 (N_21166,N_19297,N_19511);
nand U21167 (N_21167,N_19540,N_19147);
and U21168 (N_21168,N_18983,N_19344);
and U21169 (N_21169,N_19172,N_18912);
and U21170 (N_21170,N_19119,N_19414);
or U21171 (N_21171,N_19569,N_18891);
nand U21172 (N_21172,N_19945,N_19663);
or U21173 (N_21173,N_19409,N_18826);
nor U21174 (N_21174,N_19850,N_18859);
nor U21175 (N_21175,N_19235,N_19326);
nor U21176 (N_21176,N_19439,N_19009);
and U21177 (N_21177,N_19128,N_19605);
nand U21178 (N_21178,N_19095,N_19675);
or U21179 (N_21179,N_18958,N_19875);
nand U21180 (N_21180,N_19233,N_19522);
xor U21181 (N_21181,N_18765,N_19825);
or U21182 (N_21182,N_19653,N_19328);
and U21183 (N_21183,N_19605,N_19452);
or U21184 (N_21184,N_19017,N_19625);
xor U21185 (N_21185,N_18982,N_19133);
nand U21186 (N_21186,N_18887,N_18942);
xnor U21187 (N_21187,N_18774,N_18913);
nor U21188 (N_21188,N_19850,N_19324);
or U21189 (N_21189,N_18922,N_19070);
nand U21190 (N_21190,N_18882,N_18953);
or U21191 (N_21191,N_18958,N_19206);
xnor U21192 (N_21192,N_19005,N_19396);
and U21193 (N_21193,N_19954,N_18923);
nor U21194 (N_21194,N_19544,N_19534);
nor U21195 (N_21195,N_19422,N_19109);
xor U21196 (N_21196,N_19801,N_19428);
nor U21197 (N_21197,N_19089,N_19175);
nand U21198 (N_21198,N_19621,N_19093);
and U21199 (N_21199,N_19519,N_19044);
xor U21200 (N_21200,N_19085,N_19275);
xnor U21201 (N_21201,N_19801,N_19655);
nor U21202 (N_21202,N_19461,N_19533);
nor U21203 (N_21203,N_18966,N_19144);
nand U21204 (N_21204,N_18987,N_18998);
xnor U21205 (N_21205,N_19348,N_19280);
nand U21206 (N_21206,N_18971,N_19534);
and U21207 (N_21207,N_19848,N_19360);
and U21208 (N_21208,N_19861,N_19664);
and U21209 (N_21209,N_18809,N_19183);
xor U21210 (N_21210,N_19020,N_19170);
or U21211 (N_21211,N_18837,N_19106);
and U21212 (N_21212,N_19721,N_19321);
xnor U21213 (N_21213,N_19405,N_19058);
or U21214 (N_21214,N_19353,N_18786);
or U21215 (N_21215,N_19714,N_19314);
nor U21216 (N_21216,N_18998,N_19408);
xnor U21217 (N_21217,N_19107,N_19105);
nand U21218 (N_21218,N_19160,N_19207);
nand U21219 (N_21219,N_19907,N_19031);
nand U21220 (N_21220,N_19799,N_19427);
nor U21221 (N_21221,N_19752,N_19458);
nor U21222 (N_21222,N_18929,N_19664);
or U21223 (N_21223,N_19911,N_19446);
nor U21224 (N_21224,N_19833,N_18811);
or U21225 (N_21225,N_18792,N_19328);
xor U21226 (N_21226,N_19747,N_19801);
nor U21227 (N_21227,N_19369,N_19357);
xor U21228 (N_21228,N_19931,N_19153);
nor U21229 (N_21229,N_19196,N_19739);
nand U21230 (N_21230,N_19295,N_19286);
and U21231 (N_21231,N_18832,N_19340);
or U21232 (N_21232,N_19693,N_19492);
xnor U21233 (N_21233,N_19905,N_19386);
and U21234 (N_21234,N_18786,N_19533);
xor U21235 (N_21235,N_19255,N_18905);
and U21236 (N_21236,N_19726,N_19417);
nor U21237 (N_21237,N_19496,N_19810);
nand U21238 (N_21238,N_19751,N_19482);
nor U21239 (N_21239,N_19028,N_19882);
and U21240 (N_21240,N_18979,N_19750);
xor U21241 (N_21241,N_19503,N_19105);
xnor U21242 (N_21242,N_18878,N_19122);
nand U21243 (N_21243,N_19803,N_19236);
or U21244 (N_21244,N_19497,N_19549);
and U21245 (N_21245,N_18801,N_19910);
or U21246 (N_21246,N_19146,N_19454);
nand U21247 (N_21247,N_19931,N_19919);
or U21248 (N_21248,N_19077,N_18776);
xnor U21249 (N_21249,N_18960,N_19129);
xnor U21250 (N_21250,N_20262,N_20427);
nand U21251 (N_21251,N_20714,N_20197);
nor U21252 (N_21252,N_20784,N_20046);
nand U21253 (N_21253,N_21106,N_20214);
and U21254 (N_21254,N_20162,N_20238);
or U21255 (N_21255,N_20710,N_20827);
and U21256 (N_21256,N_21127,N_21019);
and U21257 (N_21257,N_20057,N_20289);
and U21258 (N_21258,N_20861,N_20912);
or U21259 (N_21259,N_20587,N_20292);
and U21260 (N_21260,N_20791,N_21072);
nor U21261 (N_21261,N_20750,N_20481);
and U21262 (N_21262,N_21008,N_20561);
or U21263 (N_21263,N_20053,N_20319);
nand U21264 (N_21264,N_20568,N_20439);
and U21265 (N_21265,N_21213,N_20550);
and U21266 (N_21266,N_21104,N_20217);
or U21267 (N_21267,N_20735,N_20064);
nand U21268 (N_21268,N_20233,N_20258);
nand U21269 (N_21269,N_20456,N_20573);
nand U21270 (N_21270,N_20286,N_20694);
nor U21271 (N_21271,N_20876,N_20728);
xor U21272 (N_21272,N_20212,N_20186);
or U21273 (N_21273,N_20285,N_21047);
nor U21274 (N_21274,N_20535,N_21099);
or U21275 (N_21275,N_20756,N_20613);
nor U21276 (N_21276,N_20173,N_21087);
and U21277 (N_21277,N_20668,N_20744);
nor U21278 (N_21278,N_20158,N_21188);
or U21279 (N_21279,N_20007,N_20591);
xor U21280 (N_21280,N_20371,N_20108);
or U21281 (N_21281,N_20468,N_20880);
or U21282 (N_21282,N_20828,N_20630);
nor U21283 (N_21283,N_20265,N_20216);
xor U21284 (N_21284,N_20628,N_20224);
nor U21285 (N_21285,N_20365,N_21064);
and U21286 (N_21286,N_20625,N_20070);
or U21287 (N_21287,N_20316,N_20247);
and U21288 (N_21288,N_20367,N_20690);
xnor U21289 (N_21289,N_21229,N_20418);
or U21290 (N_21290,N_20801,N_20860);
nor U21291 (N_21291,N_20649,N_20723);
nand U21292 (N_21292,N_20597,N_20871);
nand U21293 (N_21293,N_20362,N_20603);
nand U21294 (N_21294,N_20766,N_20101);
or U21295 (N_21295,N_21235,N_20038);
or U21296 (N_21296,N_20395,N_21172);
or U21297 (N_21297,N_20875,N_20726);
nor U21298 (N_21298,N_20127,N_21012);
nand U21299 (N_21299,N_20229,N_20522);
xnor U21300 (N_21300,N_21114,N_20093);
nand U21301 (N_21301,N_20052,N_21002);
nand U21302 (N_21302,N_20202,N_20375);
xnor U21303 (N_21303,N_20817,N_21025);
xnor U21304 (N_21304,N_20465,N_20678);
nor U21305 (N_21305,N_20517,N_20097);
xor U21306 (N_21306,N_20109,N_20176);
and U21307 (N_21307,N_20933,N_21043);
nor U21308 (N_21308,N_20204,N_20949);
nand U21309 (N_21309,N_20156,N_20639);
or U21310 (N_21310,N_20823,N_20960);
nand U21311 (N_21311,N_21111,N_20161);
nor U21312 (N_21312,N_21065,N_20620);
nand U21313 (N_21313,N_21187,N_20048);
and U21314 (N_21314,N_20011,N_20488);
nand U21315 (N_21315,N_21095,N_20434);
nor U21316 (N_21316,N_21158,N_20842);
xor U21317 (N_21317,N_20157,N_20938);
or U21318 (N_21318,N_21112,N_20808);
nand U21319 (N_21319,N_20719,N_20453);
xor U21320 (N_21320,N_20058,N_20026);
nand U21321 (N_21321,N_20687,N_20255);
and U21322 (N_21322,N_21196,N_20899);
nand U21323 (N_21323,N_20961,N_20650);
xnor U21324 (N_21324,N_21199,N_20996);
nand U21325 (N_21325,N_20235,N_20787);
and U21326 (N_21326,N_20742,N_20672);
nand U21327 (N_21327,N_20629,N_20356);
and U21328 (N_21328,N_21056,N_20745);
xnor U21329 (N_21329,N_21139,N_20777);
nand U21330 (N_21330,N_20187,N_20922);
or U21331 (N_21331,N_20018,N_20049);
nand U21332 (N_21332,N_20703,N_20680);
and U21333 (N_21333,N_20581,N_21046);
xor U21334 (N_21334,N_20815,N_20270);
or U21335 (N_21335,N_20479,N_21226);
nor U21336 (N_21336,N_21244,N_20409);
nand U21337 (N_21337,N_20394,N_20849);
xor U21338 (N_21338,N_20106,N_21118);
nand U21339 (N_21339,N_20884,N_21146);
nand U21340 (N_21340,N_20490,N_20373);
nor U21341 (N_21341,N_20866,N_20067);
or U21342 (N_21342,N_20227,N_20753);
xor U21343 (N_21343,N_20492,N_20724);
nor U21344 (N_21344,N_20775,N_20600);
nand U21345 (N_21345,N_20306,N_20565);
and U21346 (N_21346,N_20413,N_20612);
or U21347 (N_21347,N_20772,N_20245);
nor U21348 (N_21348,N_20722,N_20334);
xor U21349 (N_21349,N_20196,N_20201);
nor U21350 (N_21350,N_20976,N_21137);
and U21351 (N_21351,N_20877,N_20607);
or U21352 (N_21352,N_20206,N_20814);
and U21353 (N_21353,N_20741,N_20405);
xor U21354 (N_21354,N_20647,N_21058);
xor U21355 (N_21355,N_20389,N_20303);
nor U21356 (N_21356,N_20354,N_20429);
xnor U21357 (N_21357,N_20177,N_20061);
nor U21358 (N_21358,N_20448,N_20623);
and U21359 (N_21359,N_21030,N_20034);
and U21360 (N_21360,N_20361,N_21132);
xor U21361 (N_21361,N_20560,N_20077);
xnor U21362 (N_21362,N_20614,N_20952);
xor U21363 (N_21363,N_21084,N_20717);
nor U21364 (N_21364,N_20886,N_20805);
nand U21365 (N_21365,N_20256,N_21067);
and U21366 (N_21366,N_20919,N_20858);
nor U21367 (N_21367,N_21153,N_20326);
xnor U21368 (N_21368,N_20888,N_20896);
xor U21369 (N_21369,N_21221,N_21133);
or U21370 (N_21370,N_20622,N_20348);
and U21371 (N_21371,N_20205,N_20435);
xor U21372 (N_21372,N_20243,N_21219);
and U21373 (N_21373,N_21097,N_20540);
or U21374 (N_21374,N_20733,N_21026);
and U21375 (N_21375,N_20826,N_20529);
nor U21376 (N_21376,N_20758,N_20044);
nor U21377 (N_21377,N_20763,N_20019);
nor U21378 (N_21378,N_20720,N_20004);
nand U21379 (N_21379,N_21128,N_20194);
or U21380 (N_21380,N_20115,N_20679);
and U21381 (N_21381,N_20638,N_20845);
or U21382 (N_21382,N_20892,N_20583);
and U21383 (N_21383,N_20898,N_20426);
and U21384 (N_21384,N_21242,N_20313);
and U21385 (N_21385,N_20921,N_20795);
nand U21386 (N_21386,N_20520,N_20513);
xnor U21387 (N_21387,N_21131,N_20928);
nor U21388 (N_21388,N_21232,N_20139);
or U21389 (N_21389,N_20515,N_21005);
xor U21390 (N_21390,N_20037,N_21107);
or U21391 (N_21391,N_20979,N_21037);
nor U21392 (N_21392,N_20589,N_20980);
or U21393 (N_21393,N_20116,N_20611);
nand U21394 (N_21394,N_20022,N_20219);
or U21395 (N_21395,N_21203,N_20015);
and U21396 (N_21396,N_20489,N_20605);
nand U21397 (N_21397,N_21222,N_21238);
or U21398 (N_21398,N_20799,N_20510);
nand U21399 (N_21399,N_20103,N_21171);
and U21400 (N_21400,N_20916,N_20183);
and U21401 (N_21401,N_21062,N_20908);
or U21402 (N_21402,N_20910,N_20014);
nand U21403 (N_21403,N_21050,N_20800);
xor U21404 (N_21404,N_20001,N_20006);
and U21405 (N_21405,N_20191,N_20331);
xor U21406 (N_21406,N_20080,N_21006);
or U21407 (N_21407,N_20350,N_20830);
xor U21408 (N_21408,N_20125,N_20478);
or U21409 (N_21409,N_20447,N_20463);
nand U21410 (N_21410,N_20946,N_20947);
or U21411 (N_21411,N_21053,N_20953);
xor U21412 (N_21412,N_20360,N_20152);
xnor U21413 (N_21413,N_20914,N_20287);
or U21414 (N_21414,N_20382,N_20170);
or U21415 (N_21415,N_21068,N_20838);
or U21416 (N_21416,N_20280,N_20084);
or U21417 (N_21417,N_20344,N_21079);
or U21418 (N_21418,N_20905,N_20786);
or U21419 (N_21419,N_20768,N_20856);
and U21420 (N_21420,N_21191,N_20959);
nand U21421 (N_21421,N_20254,N_20543);
xnor U21422 (N_21422,N_21020,N_21011);
and U21423 (N_21423,N_20918,N_20577);
or U21424 (N_21424,N_21181,N_21208);
and U21425 (N_21425,N_20132,N_20738);
nor U21426 (N_21426,N_20220,N_21023);
and U21427 (N_21427,N_21215,N_20472);
or U21428 (N_21428,N_20062,N_20269);
nand U21429 (N_21429,N_20123,N_20047);
and U21430 (N_21430,N_21078,N_20904);
nand U21431 (N_21431,N_20552,N_20785);
or U21432 (N_21432,N_20562,N_20819);
and U21433 (N_21433,N_20137,N_21141);
xnor U21434 (N_21434,N_20120,N_20844);
xnor U21435 (N_21435,N_20988,N_20083);
nand U21436 (N_21436,N_20652,N_20634);
or U21437 (N_21437,N_20477,N_21123);
and U21438 (N_21438,N_20221,N_20782);
and U21439 (N_21439,N_20347,N_20748);
nor U21440 (N_21440,N_21063,N_20767);
nor U21441 (N_21441,N_21200,N_20383);
xor U21442 (N_21442,N_20151,N_20537);
nor U21443 (N_21443,N_20755,N_20230);
or U21444 (N_21444,N_20190,N_20119);
nor U21445 (N_21445,N_21246,N_20110);
and U21446 (N_21446,N_20602,N_20760);
xnor U21447 (N_21447,N_20803,N_21041);
and U21448 (N_21448,N_20297,N_20182);
nor U21449 (N_21449,N_20259,N_20915);
xor U21450 (N_21450,N_20284,N_21166);
and U21451 (N_21451,N_21113,N_20764);
and U21452 (N_21452,N_20480,N_21057);
xnor U21453 (N_21453,N_20731,N_20962);
and U21454 (N_21454,N_20374,N_20497);
or U21455 (N_21455,N_20700,N_20539);
nor U21456 (N_21456,N_20820,N_20833);
nor U21457 (N_21457,N_20525,N_21098);
nor U21458 (N_21458,N_20536,N_20295);
xnor U21459 (N_21459,N_20706,N_21180);
nor U21460 (N_21460,N_20094,N_21243);
or U21461 (N_21461,N_20407,N_21125);
or U21462 (N_21462,N_20086,N_20797);
or U21463 (N_21463,N_20812,N_20872);
and U21464 (N_21464,N_20163,N_20288);
nor U21465 (N_21465,N_20926,N_21070);
or U21466 (N_21466,N_20692,N_20563);
nor U21467 (N_21467,N_20707,N_20586);
xnor U21468 (N_21468,N_20521,N_20958);
or U21469 (N_21469,N_21239,N_20232);
or U21470 (N_21470,N_20166,N_20894);
nand U21471 (N_21471,N_20020,N_20364);
nand U21472 (N_21472,N_21224,N_21186);
xor U21473 (N_21473,N_21152,N_20032);
or U21474 (N_21474,N_20028,N_20400);
or U21475 (N_21475,N_20148,N_20403);
xor U21476 (N_21476,N_21103,N_20693);
xnor U21477 (N_21477,N_21124,N_20927);
and U21478 (N_21478,N_20301,N_20829);
xnor U21479 (N_21479,N_20740,N_21044);
xor U21480 (N_21480,N_20831,N_20111);
nor U21481 (N_21481,N_20516,N_20462);
nor U21482 (N_21482,N_20601,N_21147);
and U21483 (N_21483,N_20683,N_20903);
or U21484 (N_21484,N_20322,N_20832);
xor U21485 (N_21485,N_20566,N_20174);
or U21486 (N_21486,N_20199,N_20008);
nand U21487 (N_21487,N_20632,N_21110);
nand U21488 (N_21488,N_21143,N_20276);
and U21489 (N_21489,N_20974,N_21201);
nor U21490 (N_21490,N_20822,N_20495);
nor U21491 (N_21491,N_20160,N_20913);
nand U21492 (N_21492,N_20428,N_20935);
nand U21493 (N_21493,N_20957,N_20633);
nand U21494 (N_21494,N_20443,N_20130);
nand U21495 (N_21495,N_20185,N_20095);
xnor U21496 (N_21496,N_20423,N_20684);
nor U21497 (N_21497,N_20983,N_20171);
and U21498 (N_21498,N_20941,N_20792);
and U21499 (N_21499,N_20518,N_20266);
and U21500 (N_21500,N_20937,N_20340);
xor U21501 (N_21501,N_20482,N_20604);
nand U21502 (N_21502,N_20511,N_21119);
and U21503 (N_21503,N_21059,N_20016);
nand U21504 (N_21504,N_20392,N_20328);
xnor U21505 (N_21505,N_20847,N_20757);
nand U21506 (N_21506,N_20655,N_20925);
xnor U21507 (N_21507,N_20461,N_20549);
and U21508 (N_21508,N_20762,N_20711);
or U21509 (N_21509,N_20725,N_20734);
xnor U21510 (N_21510,N_21082,N_20942);
or U21511 (N_21511,N_20385,N_20716);
nand U21512 (N_21512,N_20027,N_21129);
or U21513 (N_21513,N_21135,N_20642);
and U21514 (N_21514,N_20404,N_21231);
or U21515 (N_21515,N_20260,N_21134);
and U21516 (N_21516,N_20451,N_20977);
nor U21517 (N_21517,N_20090,N_20105);
nand U21518 (N_21518,N_20487,N_21149);
nor U21519 (N_21519,N_20596,N_20907);
or U21520 (N_21520,N_21175,N_20682);
nand U21521 (N_21521,N_20494,N_20558);
or U21522 (N_21522,N_21066,N_20923);
or U21523 (N_21523,N_21193,N_20689);
xor U21524 (N_21524,N_21090,N_20211);
or U21525 (N_21525,N_20144,N_20437);
xor U21526 (N_21526,N_20442,N_20834);
or U21527 (N_21527,N_20155,N_20865);
nor U21528 (N_21528,N_20851,N_20593);
nor U21529 (N_21529,N_20023,N_20180);
xnor U21530 (N_21530,N_21016,N_20342);
xnor U21531 (N_21531,N_20388,N_20878);
xor U21532 (N_21532,N_20121,N_20685);
nor U21533 (N_21533,N_20450,N_20721);
or U21534 (N_21534,N_20474,N_20029);
xor U21535 (N_21535,N_20298,N_20751);
and U21536 (N_21536,N_21197,N_20496);
nor U21537 (N_21537,N_20493,N_21048);
xnor U21538 (N_21538,N_20664,N_20159);
or U21539 (N_21539,N_20718,N_20533);
nor U21540 (N_21540,N_20778,N_20055);
xnor U21541 (N_21541,N_21086,N_21045);
or U21542 (N_21542,N_20794,N_20261);
xor U21543 (N_21543,N_20686,N_20984);
nand U21544 (N_21544,N_20631,N_20291);
nor U21545 (N_21545,N_20075,N_20353);
nor U21546 (N_21546,N_20126,N_20370);
and U21547 (N_21547,N_20882,N_20397);
nand U21548 (N_21548,N_21077,N_20452);
or U21549 (N_21549,N_20372,N_21209);
and U21550 (N_21550,N_21102,N_20730);
nor U21551 (N_21551,N_20645,N_20141);
nand U21552 (N_21552,N_20341,N_20239);
nand U21553 (N_21553,N_20338,N_20060);
and U21554 (N_21554,N_21055,N_20867);
and U21555 (N_21555,N_21126,N_20272);
and U21556 (N_21556,N_20868,N_20594);
or U21557 (N_21557,N_21145,N_21073);
or U21558 (N_21558,N_20242,N_20635);
and U21559 (N_21559,N_21021,N_20131);
nor U21560 (N_21560,N_21051,N_20906);
nor U21561 (N_21561,N_20499,N_20747);
or U21562 (N_21562,N_20050,N_20327);
xor U21563 (N_21563,N_21100,N_21009);
nand U21564 (N_21564,N_20500,N_20853);
or U21565 (N_21565,N_20809,N_20530);
nand U21566 (N_21566,N_20615,N_21085);
or U21567 (N_21567,N_20088,N_21092);
nor U21568 (N_21568,N_20556,N_21202);
nand U21569 (N_21569,N_20749,N_20253);
nor U21570 (N_21570,N_20323,N_20967);
xnor U21571 (N_21571,N_20042,N_20930);
nor U21572 (N_21572,N_20352,N_20897);
xnor U21573 (N_21573,N_20396,N_21151);
nand U21574 (N_21574,N_20311,N_20512);
nand U21575 (N_21575,N_20358,N_21237);
xor U21576 (N_21576,N_20349,N_21015);
and U21577 (N_21577,N_20788,N_21109);
nor U21578 (N_21578,N_20172,N_20329);
or U21579 (N_21579,N_20267,N_20699);
and U21580 (N_21580,N_20430,N_20807);
xnor U21581 (N_21581,N_20134,N_21184);
nand U21582 (N_21582,N_20676,N_20653);
and U21583 (N_21583,N_20818,N_20454);
or U21584 (N_21584,N_21083,N_20932);
nor U21585 (N_21585,N_20595,N_20293);
nand U21586 (N_21586,N_20641,N_20440);
or U21587 (N_21587,N_21168,N_20455);
nor U21588 (N_21588,N_20471,N_20688);
xor U21589 (N_21589,N_21182,N_20142);
and U21590 (N_21590,N_20290,N_20165);
xnor U21591 (N_21591,N_20574,N_21211);
and U21592 (N_21592,N_20950,N_20965);
nor U21593 (N_21593,N_20781,N_20491);
nand U21594 (N_21594,N_20609,N_21121);
and U21595 (N_21595,N_21052,N_20945);
or U21596 (N_21596,N_20459,N_20357);
or U21597 (N_21597,N_20841,N_21003);
nor U21598 (N_21598,N_20436,N_20863);
nor U21599 (N_21599,N_20542,N_20376);
nand U21600 (N_21600,N_21013,N_21154);
or U21601 (N_21601,N_21160,N_20143);
nand U21602 (N_21602,N_20296,N_20765);
xor U21603 (N_21603,N_20909,N_20585);
and U21604 (N_21604,N_21198,N_21130);
nor U21605 (N_21605,N_20599,N_20986);
nor U21606 (N_21606,N_20104,N_20264);
xor U21607 (N_21607,N_20729,N_20770);
nor U21608 (N_21608,N_20534,N_20963);
or U21609 (N_21609,N_20790,N_20508);
nor U21610 (N_21610,N_20059,N_20954);
nor U21611 (N_21611,N_20982,N_20231);
or U21612 (N_21612,N_20846,N_20502);
xnor U21613 (N_21613,N_20637,N_21225);
nand U21614 (N_21614,N_20030,N_20704);
xnor U21615 (N_21615,N_20147,N_20773);
and U21616 (N_21616,N_20627,N_20040);
and U21617 (N_21617,N_20793,N_20900);
and U21618 (N_21618,N_20228,N_20249);
nand U21619 (N_21619,N_20616,N_20314);
nor U21620 (N_21620,N_20324,N_20154);
nor U21621 (N_21621,N_20325,N_20643);
and U21622 (N_21622,N_20852,N_21069);
xnor U21623 (N_21623,N_20387,N_20063);
nor U21624 (N_21624,N_20505,N_20210);
nor U21625 (N_21625,N_21206,N_21105);
xor U21626 (N_21626,N_20662,N_20691);
nand U21627 (N_21627,N_21101,N_20895);
and U21628 (N_21628,N_21207,N_21178);
xnor U21629 (N_21629,N_20582,N_20263);
xnor U21630 (N_21630,N_21228,N_21165);
nand U21631 (N_21631,N_20332,N_20971);
or U21632 (N_21632,N_21122,N_20570);
nor U21633 (N_21633,N_21108,N_20506);
or U21634 (N_21634,N_21024,N_20567);
nand U21635 (N_21635,N_21223,N_20660);
xor U21636 (N_21636,N_20003,N_21000);
nand U21637 (N_21637,N_20771,N_21039);
nand U21638 (N_21638,N_20975,N_20779);
nor U21639 (N_21639,N_20114,N_20990);
xnor U21640 (N_21640,N_20416,N_21230);
xnor U21641 (N_21641,N_20117,N_20420);
nand U21642 (N_21642,N_20002,N_20449);
nor U21643 (N_21643,N_20519,N_21138);
nand U21644 (N_21644,N_20369,N_20695);
xnor U21645 (N_21645,N_21049,N_20780);
or U21646 (N_21646,N_21216,N_20079);
xor U21647 (N_21647,N_20864,N_20355);
xor U21648 (N_21648,N_21032,N_20207);
or U21649 (N_21649,N_20215,N_20544);
nor U21650 (N_21650,N_20802,N_20939);
or U21651 (N_21651,N_20661,N_20065);
nand U21652 (N_21652,N_20066,N_20712);
xor U21653 (N_21653,N_20398,N_20315);
or U21654 (N_21654,N_20318,N_21014);
nor U21655 (N_21655,N_21150,N_20610);
and U21656 (N_21656,N_20564,N_20309);
and U21657 (N_21657,N_21117,N_21081);
and U21658 (N_21658,N_20783,N_20124);
and U21659 (N_21659,N_21233,N_21115);
and U21660 (N_21660,N_20769,N_20806);
and U21661 (N_21661,N_20981,N_20244);
nor U21662 (N_21662,N_20943,N_20091);
or U21663 (N_21663,N_20545,N_20366);
nor U21664 (N_21664,N_20789,N_20483);
or U21665 (N_21665,N_20598,N_20969);
and U21666 (N_21666,N_20346,N_20917);
xor U21667 (N_21667,N_21093,N_20054);
xor U21668 (N_21668,N_20624,N_20636);
nor U21669 (N_21669,N_20879,N_20862);
nand U21670 (N_21670,N_20514,N_20705);
nor U21671 (N_21671,N_21035,N_20994);
or U21672 (N_21672,N_20133,N_20071);
and U21673 (N_21673,N_21240,N_20317);
and U21674 (N_21674,N_20074,N_20445);
nor U21675 (N_21675,N_20150,N_21116);
xnor U21676 (N_21676,N_21094,N_20709);
nand U21677 (N_21677,N_20485,N_20476);
nor U21678 (N_21678,N_20648,N_20417);
and U21679 (N_21679,N_20363,N_21169);
or U21680 (N_21680,N_20275,N_21157);
xnor U21681 (N_21681,N_20881,N_20218);
and U21682 (N_21682,N_20701,N_20464);
or U21683 (N_21683,N_21148,N_20246);
nand U21684 (N_21684,N_20532,N_20393);
xnor U21685 (N_21685,N_21004,N_20282);
nor U21686 (N_21686,N_20466,N_21010);
nand U21687 (N_21687,N_20608,N_20368);
xor U21688 (N_21688,N_20248,N_20901);
or U21689 (N_21689,N_21185,N_20069);
nor U21690 (N_21690,N_20667,N_20811);
nand U21691 (N_21691,N_20874,N_21120);
nor U21692 (N_21692,N_20840,N_20796);
and U21693 (N_21693,N_20848,N_20873);
nor U21694 (N_21694,N_20359,N_20209);
nor U21695 (N_21695,N_20056,N_20200);
xnor U21696 (N_21696,N_20675,N_20893);
and U21697 (N_21697,N_20527,N_20618);
or U21698 (N_21698,N_21162,N_20619);
and U21699 (N_21699,N_21174,N_20526);
nor U21700 (N_21700,N_20569,N_21210);
and U21701 (N_21701,N_20300,N_20081);
nor U21702 (N_21702,N_20135,N_20198);
and U21703 (N_21703,N_20970,N_20934);
xnor U21704 (N_21704,N_20005,N_21142);
nor U21705 (N_21705,N_21227,N_20145);
nand U21706 (N_21706,N_20089,N_20911);
xor U21707 (N_21707,N_20681,N_20551);
or U21708 (N_21708,N_20955,N_20531);
xnor U21709 (N_21709,N_20113,N_20665);
xnor U21710 (N_21710,N_20136,N_20237);
nor U21711 (N_21711,N_20181,N_20924);
nand U21712 (N_21712,N_20669,N_20737);
nand U21713 (N_21713,N_20484,N_20754);
nor U21714 (N_21714,N_20013,N_20989);
nor U21715 (N_21715,N_20978,N_20441);
xnor U21716 (N_21716,N_20887,N_20250);
nor U21717 (N_21717,N_20039,N_20336);
nor U21718 (N_21718,N_20225,N_20128);
or U21719 (N_21719,N_20837,N_20855);
xor U21720 (N_21720,N_20998,N_20257);
and U21721 (N_21721,N_20333,N_20951);
and U21722 (N_21722,N_20509,N_20548);
or U21723 (N_21723,N_20412,N_20241);
nand U21724 (N_21724,N_20184,N_20761);
xnor U21725 (N_21725,N_20944,N_21029);
or U21726 (N_21726,N_20072,N_21183);
and U21727 (N_21727,N_20107,N_20178);
nor U21728 (N_21728,N_20415,N_20964);
xnor U21729 (N_21729,N_20281,N_20175);
xor U21730 (N_21730,N_20816,N_20621);
nand U21731 (N_21731,N_20438,N_20379);
nand U21732 (N_21732,N_20213,N_20697);
or U21733 (N_21733,N_21033,N_20671);
and U21734 (N_21734,N_20674,N_21071);
nand U21735 (N_21735,N_20966,N_21195);
xor U21736 (N_21736,N_20592,N_21212);
or U21737 (N_21737,N_20017,N_21089);
nor U21738 (N_21738,N_20885,N_20335);
nand U21739 (N_21739,N_21249,N_21245);
or U21740 (N_21740,N_20626,N_20188);
nor U21741 (N_21741,N_20920,N_20223);
and U21742 (N_21742,N_20985,N_20743);
nor U21743 (N_21743,N_21054,N_21234);
nand U21744 (N_21744,N_20657,N_20195);
xor U21745 (N_21745,N_20859,N_20553);
nor U21746 (N_21746,N_20078,N_20138);
xor U21747 (N_21747,N_20226,N_21159);
or U21748 (N_21748,N_20644,N_20992);
nand U21749 (N_21749,N_20843,N_20098);
and U21750 (N_21750,N_20000,N_20702);
or U21751 (N_21751,N_20713,N_20384);
and U21752 (N_21752,N_20351,N_20475);
or U21753 (N_21753,N_20045,N_20422);
or U21754 (N_21754,N_20677,N_20473);
and U21755 (N_21755,N_20559,N_20425);
or U21756 (N_21756,N_20798,N_20824);
and U21757 (N_21757,N_20854,N_21022);
nor U21758 (N_21758,N_21034,N_21144);
nand U21759 (N_21759,N_20240,N_20554);
nor U21760 (N_21760,N_20759,N_20321);
nand U21761 (N_21761,N_20192,N_21163);
xor U21762 (N_21762,N_20189,N_20839);
and U21763 (N_21763,N_20659,N_21189);
nor U21764 (N_21764,N_20575,N_20997);
or U21765 (N_21765,N_21236,N_21038);
nand U21766 (N_21766,N_20024,N_20337);
xnor U21767 (N_21767,N_20857,N_21218);
xnor U21768 (N_21768,N_21164,N_20129);
nor U21769 (N_21769,N_20654,N_20294);
xnor U21770 (N_21770,N_20410,N_20033);
nand U21771 (N_21771,N_20305,N_20414);
xnor U21772 (N_21772,N_20009,N_20572);
xnor U21773 (N_21773,N_20401,N_20169);
xnor U21774 (N_21774,N_20715,N_20696);
and U21775 (N_21775,N_20835,N_21247);
nor U21776 (N_21776,N_20076,N_20087);
and U21777 (N_21777,N_20390,N_20578);
xnor U21778 (N_21778,N_20419,N_20666);
and U21779 (N_21779,N_20617,N_20339);
nor U21780 (N_21780,N_20698,N_20739);
nand U21781 (N_21781,N_20956,N_20646);
xnor U21782 (N_21782,N_20774,N_20467);
xor U21783 (N_21783,N_20557,N_20252);
nand U21784 (N_21784,N_20547,N_20082);
or U21785 (N_21785,N_20085,N_21220);
xor U21786 (N_21786,N_20528,N_20523);
nor U21787 (N_21787,N_20579,N_21192);
nand U21788 (N_21788,N_20279,N_20460);
xnor U21789 (N_21789,N_21248,N_21028);
nand U21790 (N_21790,N_20444,N_20498);
xor U21791 (N_21791,N_20068,N_21205);
and U21792 (N_21792,N_20973,N_20380);
nor U21793 (N_21793,N_20102,N_20968);
nor U21794 (N_21794,N_20931,N_20164);
or U21795 (N_21795,N_20277,N_20651);
xor U21796 (N_21796,N_20821,N_20889);
nand U21797 (N_21797,N_21018,N_20524);
or U21798 (N_21798,N_20810,N_21001);
nand U21799 (N_21799,N_21091,N_20036);
and U21800 (N_21800,N_21161,N_21088);
nand U21801 (N_21801,N_20051,N_21036);
xnor U21802 (N_21802,N_20268,N_20936);
nor U21803 (N_21803,N_20283,N_20271);
nand U21804 (N_21804,N_20776,N_20140);
and U21805 (N_21805,N_20940,N_20399);
xor U21806 (N_21806,N_20883,N_20555);
and U21807 (N_21807,N_20274,N_20096);
nor U21808 (N_21808,N_20501,N_21074);
nor U21809 (N_21809,N_20580,N_20411);
and U21810 (N_21810,N_20991,N_20836);
and U21811 (N_21811,N_20606,N_20993);
nand U21812 (N_21812,N_20458,N_21214);
nor U21813 (N_21813,N_20948,N_20663);
and U21814 (N_21814,N_21177,N_20588);
xnor U21815 (N_21815,N_21040,N_20343);
and U21816 (N_21816,N_21173,N_21156);
xnor U21817 (N_21817,N_20732,N_20402);
xnor U21818 (N_21818,N_20869,N_20307);
and U21819 (N_21819,N_20010,N_20179);
and U21820 (N_21820,N_20122,N_20149);
nor U21821 (N_21821,N_20999,N_20073);
and U21822 (N_21822,N_20146,N_21170);
nor U21823 (N_21823,N_20486,N_21241);
and U21824 (N_21824,N_20406,N_21204);
or U21825 (N_21825,N_20391,N_20386);
or U21826 (N_21826,N_20656,N_20433);
nor U21827 (N_21827,N_20092,N_20446);
nor U21828 (N_21828,N_20278,N_21076);
nor U21829 (N_21829,N_20584,N_20538);
nand U21830 (N_21830,N_20850,N_21096);
nand U21831 (N_21831,N_21167,N_21027);
or U21832 (N_21832,N_20987,N_21176);
or U21833 (N_21833,N_20752,N_21080);
nor U21834 (N_21834,N_20995,N_20902);
nand U21835 (N_21835,N_20470,N_20118);
or U21836 (N_21836,N_20432,N_20302);
nor U21837 (N_21837,N_21136,N_20308);
or U21838 (N_21838,N_20100,N_20021);
or U21839 (N_21839,N_20312,N_20236);
nand U21840 (N_21840,N_20043,N_20112);
nor U21841 (N_21841,N_20431,N_20424);
nor U21842 (N_21842,N_20099,N_20035);
nor U21843 (N_21843,N_20571,N_20727);
nand U21844 (N_21844,N_20736,N_21217);
nand U21845 (N_21845,N_20469,N_20273);
and U21846 (N_21846,N_20503,N_20804);
and U21847 (N_21847,N_21007,N_20299);
nor U21848 (N_21848,N_21140,N_21031);
and U21849 (N_21849,N_20234,N_20222);
nand U21850 (N_21850,N_20345,N_20590);
and U21851 (N_21851,N_20972,N_20310);
or U21852 (N_21852,N_20658,N_20193);
and U21853 (N_21853,N_20320,N_20670);
xnor U21854 (N_21854,N_21061,N_21190);
nand U21855 (N_21855,N_20304,N_20421);
nand U21856 (N_21856,N_21179,N_20167);
nor U21857 (N_21857,N_20813,N_20168);
nor U21858 (N_21858,N_20890,N_20330);
nor U21859 (N_21859,N_20041,N_20457);
or U21860 (N_21860,N_20825,N_20507);
or U21861 (N_21861,N_20012,N_20546);
or U21862 (N_21862,N_21075,N_20541);
nor U21863 (N_21863,N_20378,N_21060);
or U21864 (N_21864,N_20251,N_20891);
nand U21865 (N_21865,N_20870,N_20708);
nand U21866 (N_21866,N_20153,N_20576);
xnor U21867 (N_21867,N_20381,N_20673);
nand U21868 (N_21868,N_21017,N_20208);
xnor U21869 (N_21869,N_20640,N_20025);
and U21870 (N_21870,N_21155,N_20929);
or U21871 (N_21871,N_20408,N_20031);
nand U21872 (N_21872,N_21042,N_20504);
nand U21873 (N_21873,N_20377,N_20746);
xor U21874 (N_21874,N_21194,N_20203);
nand U21875 (N_21875,N_20363,N_20793);
xor U21876 (N_21876,N_20044,N_20844);
or U21877 (N_21877,N_20842,N_20662);
and U21878 (N_21878,N_20956,N_21238);
xnor U21879 (N_21879,N_20683,N_20548);
xor U21880 (N_21880,N_21170,N_20455);
and U21881 (N_21881,N_20245,N_20105);
and U21882 (N_21882,N_20634,N_20866);
nand U21883 (N_21883,N_20889,N_20817);
or U21884 (N_21884,N_20876,N_21062);
nor U21885 (N_21885,N_20015,N_20146);
or U21886 (N_21886,N_20417,N_20197);
nor U21887 (N_21887,N_21187,N_20267);
nand U21888 (N_21888,N_20838,N_20139);
nand U21889 (N_21889,N_20991,N_20970);
or U21890 (N_21890,N_21185,N_20338);
and U21891 (N_21891,N_20871,N_20035);
and U21892 (N_21892,N_20310,N_20394);
or U21893 (N_21893,N_21094,N_21070);
nand U21894 (N_21894,N_20178,N_20732);
nand U21895 (N_21895,N_20828,N_20605);
and U21896 (N_21896,N_20787,N_20935);
and U21897 (N_21897,N_20445,N_20455);
or U21898 (N_21898,N_21174,N_20211);
and U21899 (N_21899,N_21044,N_21232);
and U21900 (N_21900,N_20178,N_20003);
xnor U21901 (N_21901,N_20926,N_20744);
xnor U21902 (N_21902,N_20410,N_20242);
nor U21903 (N_21903,N_20787,N_20900);
xor U21904 (N_21904,N_20409,N_20398);
nor U21905 (N_21905,N_21236,N_20465);
nand U21906 (N_21906,N_21163,N_21133);
nor U21907 (N_21907,N_20187,N_20996);
and U21908 (N_21908,N_20163,N_20796);
and U21909 (N_21909,N_20875,N_20149);
or U21910 (N_21910,N_20202,N_20444);
nand U21911 (N_21911,N_20668,N_21094);
xnor U21912 (N_21912,N_20871,N_20160);
and U21913 (N_21913,N_20558,N_20851);
and U21914 (N_21914,N_20395,N_20196);
nor U21915 (N_21915,N_20973,N_20972);
and U21916 (N_21916,N_20333,N_21229);
nor U21917 (N_21917,N_20598,N_20700);
nand U21918 (N_21918,N_20882,N_20713);
xnor U21919 (N_21919,N_20742,N_20454);
nand U21920 (N_21920,N_20981,N_20436);
xor U21921 (N_21921,N_20787,N_20533);
and U21922 (N_21922,N_20518,N_20311);
nand U21923 (N_21923,N_20809,N_20090);
or U21924 (N_21924,N_20639,N_20293);
nand U21925 (N_21925,N_20226,N_20950);
xnor U21926 (N_21926,N_20580,N_20152);
nand U21927 (N_21927,N_21156,N_21088);
xnor U21928 (N_21928,N_20600,N_21013);
nand U21929 (N_21929,N_20421,N_21243);
and U21930 (N_21930,N_21059,N_21090);
nor U21931 (N_21931,N_20407,N_20214);
nand U21932 (N_21932,N_20928,N_21136);
nand U21933 (N_21933,N_20229,N_20610);
nor U21934 (N_21934,N_20812,N_20777);
or U21935 (N_21935,N_20466,N_20898);
nor U21936 (N_21936,N_21107,N_20685);
and U21937 (N_21937,N_20879,N_20905);
nand U21938 (N_21938,N_21157,N_20537);
xnor U21939 (N_21939,N_20693,N_21166);
nand U21940 (N_21940,N_20181,N_21004);
and U21941 (N_21941,N_20244,N_20628);
nor U21942 (N_21942,N_20430,N_20279);
xor U21943 (N_21943,N_20301,N_20350);
xnor U21944 (N_21944,N_20288,N_21041);
and U21945 (N_21945,N_20975,N_20380);
nor U21946 (N_21946,N_20837,N_20345);
nor U21947 (N_21947,N_21227,N_20001);
or U21948 (N_21948,N_20704,N_20286);
nor U21949 (N_21949,N_20480,N_20839);
xnor U21950 (N_21950,N_21004,N_20095);
nand U21951 (N_21951,N_20894,N_20537);
nand U21952 (N_21952,N_20122,N_21082);
xnor U21953 (N_21953,N_20815,N_20874);
nand U21954 (N_21954,N_20800,N_20484);
nand U21955 (N_21955,N_20305,N_20001);
and U21956 (N_21956,N_21203,N_20667);
nor U21957 (N_21957,N_20547,N_21065);
and U21958 (N_21958,N_20256,N_20694);
and U21959 (N_21959,N_20073,N_21140);
and U21960 (N_21960,N_20824,N_20738);
nand U21961 (N_21961,N_21242,N_20689);
xnor U21962 (N_21962,N_20313,N_20201);
xnor U21963 (N_21963,N_20324,N_20185);
or U21964 (N_21964,N_20685,N_20859);
nor U21965 (N_21965,N_20409,N_20248);
nor U21966 (N_21966,N_20714,N_20712);
or U21967 (N_21967,N_20966,N_20217);
nor U21968 (N_21968,N_21129,N_20174);
nor U21969 (N_21969,N_20756,N_20790);
nor U21970 (N_21970,N_20593,N_20655);
and U21971 (N_21971,N_20247,N_20824);
xnor U21972 (N_21972,N_20346,N_20454);
or U21973 (N_21973,N_21004,N_20447);
nor U21974 (N_21974,N_20055,N_20144);
or U21975 (N_21975,N_20465,N_20810);
xnor U21976 (N_21976,N_20164,N_20439);
nor U21977 (N_21977,N_20113,N_21106);
xor U21978 (N_21978,N_20167,N_20920);
nand U21979 (N_21979,N_20772,N_21151);
or U21980 (N_21980,N_21150,N_20412);
or U21981 (N_21981,N_20968,N_20789);
and U21982 (N_21982,N_20199,N_21000);
nor U21983 (N_21983,N_20381,N_21179);
nor U21984 (N_21984,N_21041,N_21216);
nand U21985 (N_21985,N_20781,N_21157);
or U21986 (N_21986,N_20074,N_21016);
xor U21987 (N_21987,N_21186,N_21159);
xor U21988 (N_21988,N_20504,N_20496);
and U21989 (N_21989,N_20142,N_20069);
or U21990 (N_21990,N_21008,N_20748);
nand U21991 (N_21991,N_20817,N_20877);
xor U21992 (N_21992,N_20093,N_21163);
nor U21993 (N_21993,N_20815,N_21063);
nor U21994 (N_21994,N_20964,N_20288);
xor U21995 (N_21995,N_21169,N_20359);
or U21996 (N_21996,N_21204,N_20062);
and U21997 (N_21997,N_21019,N_21033);
and U21998 (N_21998,N_21066,N_20474);
xnor U21999 (N_21999,N_20678,N_20262);
xnor U22000 (N_22000,N_20238,N_20105);
nand U22001 (N_22001,N_20813,N_20601);
nand U22002 (N_22002,N_21237,N_20641);
or U22003 (N_22003,N_20211,N_20081);
or U22004 (N_22004,N_20687,N_20980);
xnor U22005 (N_22005,N_21020,N_20265);
xnor U22006 (N_22006,N_20766,N_20510);
and U22007 (N_22007,N_21119,N_20042);
nor U22008 (N_22008,N_21184,N_20297);
xor U22009 (N_22009,N_20484,N_21179);
or U22010 (N_22010,N_20199,N_21206);
nand U22011 (N_22011,N_21180,N_20410);
nand U22012 (N_22012,N_20428,N_20911);
xnor U22013 (N_22013,N_20399,N_20479);
nand U22014 (N_22014,N_21146,N_20334);
nand U22015 (N_22015,N_21246,N_20442);
and U22016 (N_22016,N_20451,N_21158);
nand U22017 (N_22017,N_20290,N_20837);
or U22018 (N_22018,N_21101,N_20950);
nor U22019 (N_22019,N_21158,N_20025);
nand U22020 (N_22020,N_21127,N_21157);
xnor U22021 (N_22021,N_20275,N_20045);
nand U22022 (N_22022,N_20526,N_20836);
nor U22023 (N_22023,N_21178,N_20909);
or U22024 (N_22024,N_20040,N_20823);
xnor U22025 (N_22025,N_20351,N_20197);
xnor U22026 (N_22026,N_20682,N_21048);
and U22027 (N_22027,N_20110,N_20283);
nand U22028 (N_22028,N_20172,N_20344);
nand U22029 (N_22029,N_20754,N_20337);
nand U22030 (N_22030,N_20365,N_20092);
nand U22031 (N_22031,N_20836,N_20605);
nand U22032 (N_22032,N_20767,N_20531);
and U22033 (N_22033,N_20275,N_20088);
or U22034 (N_22034,N_20382,N_20679);
nor U22035 (N_22035,N_21168,N_20705);
and U22036 (N_22036,N_20007,N_21021);
and U22037 (N_22037,N_20458,N_20377);
xor U22038 (N_22038,N_20538,N_21004);
and U22039 (N_22039,N_21248,N_20469);
and U22040 (N_22040,N_20669,N_20176);
and U22041 (N_22041,N_20039,N_20306);
nand U22042 (N_22042,N_20051,N_20274);
and U22043 (N_22043,N_20916,N_21023);
and U22044 (N_22044,N_20181,N_21232);
xnor U22045 (N_22045,N_20235,N_20604);
and U22046 (N_22046,N_20145,N_20805);
and U22047 (N_22047,N_21234,N_21110);
or U22048 (N_22048,N_20372,N_20306);
nor U22049 (N_22049,N_21126,N_20804);
nand U22050 (N_22050,N_20513,N_21151);
xor U22051 (N_22051,N_20615,N_21022);
or U22052 (N_22052,N_20122,N_20912);
or U22053 (N_22053,N_20127,N_20386);
nor U22054 (N_22054,N_20837,N_20638);
xor U22055 (N_22055,N_20971,N_20620);
xor U22056 (N_22056,N_20136,N_20202);
and U22057 (N_22057,N_20614,N_20805);
nor U22058 (N_22058,N_20505,N_20075);
nor U22059 (N_22059,N_20440,N_21193);
xnor U22060 (N_22060,N_21176,N_21084);
and U22061 (N_22061,N_20598,N_20314);
nor U22062 (N_22062,N_21103,N_20668);
or U22063 (N_22063,N_20974,N_20291);
and U22064 (N_22064,N_20805,N_20607);
xor U22065 (N_22065,N_20706,N_21221);
and U22066 (N_22066,N_20265,N_20346);
xnor U22067 (N_22067,N_21195,N_21056);
or U22068 (N_22068,N_20456,N_20940);
nor U22069 (N_22069,N_20043,N_20770);
or U22070 (N_22070,N_20910,N_20020);
nor U22071 (N_22071,N_20477,N_20908);
or U22072 (N_22072,N_20296,N_20090);
or U22073 (N_22073,N_20906,N_20087);
and U22074 (N_22074,N_20648,N_20267);
xnor U22075 (N_22075,N_20525,N_20508);
or U22076 (N_22076,N_20722,N_21030);
and U22077 (N_22077,N_20710,N_20306);
nand U22078 (N_22078,N_21045,N_20354);
and U22079 (N_22079,N_20519,N_20623);
xnor U22080 (N_22080,N_20098,N_20530);
nor U22081 (N_22081,N_20989,N_20074);
nor U22082 (N_22082,N_20367,N_20390);
or U22083 (N_22083,N_20868,N_20808);
or U22084 (N_22084,N_20079,N_21214);
xnor U22085 (N_22085,N_20857,N_20678);
nand U22086 (N_22086,N_20257,N_21104);
and U22087 (N_22087,N_20470,N_20849);
nor U22088 (N_22088,N_20481,N_20001);
nand U22089 (N_22089,N_20039,N_20232);
nand U22090 (N_22090,N_20552,N_20385);
xnor U22091 (N_22091,N_20548,N_21172);
xor U22092 (N_22092,N_20055,N_20701);
nand U22093 (N_22093,N_21186,N_20604);
or U22094 (N_22094,N_20513,N_20463);
or U22095 (N_22095,N_20037,N_20431);
and U22096 (N_22096,N_21160,N_20456);
nor U22097 (N_22097,N_20040,N_20266);
nand U22098 (N_22098,N_20566,N_20323);
or U22099 (N_22099,N_20215,N_20198);
and U22100 (N_22100,N_20839,N_20625);
nand U22101 (N_22101,N_20938,N_20067);
xor U22102 (N_22102,N_21139,N_20902);
nor U22103 (N_22103,N_20151,N_20962);
nor U22104 (N_22104,N_20202,N_21169);
or U22105 (N_22105,N_21142,N_20649);
nand U22106 (N_22106,N_21227,N_20489);
or U22107 (N_22107,N_20648,N_21004);
and U22108 (N_22108,N_20135,N_20484);
and U22109 (N_22109,N_20074,N_20513);
nor U22110 (N_22110,N_20798,N_21139);
xor U22111 (N_22111,N_20114,N_20942);
nor U22112 (N_22112,N_21026,N_21024);
and U22113 (N_22113,N_21158,N_20522);
and U22114 (N_22114,N_21060,N_21053);
xor U22115 (N_22115,N_21198,N_20813);
nor U22116 (N_22116,N_20687,N_21149);
nor U22117 (N_22117,N_20798,N_20895);
xor U22118 (N_22118,N_20455,N_20284);
nand U22119 (N_22119,N_20553,N_21088);
and U22120 (N_22120,N_20589,N_20225);
nand U22121 (N_22121,N_20116,N_21244);
nor U22122 (N_22122,N_20091,N_21119);
and U22123 (N_22123,N_21086,N_21123);
nand U22124 (N_22124,N_21103,N_20729);
xor U22125 (N_22125,N_20414,N_20611);
nor U22126 (N_22126,N_20811,N_20403);
or U22127 (N_22127,N_20194,N_20732);
and U22128 (N_22128,N_20779,N_20744);
nor U22129 (N_22129,N_20685,N_20458);
or U22130 (N_22130,N_20485,N_20921);
or U22131 (N_22131,N_20868,N_20405);
xor U22132 (N_22132,N_20631,N_20111);
xnor U22133 (N_22133,N_20214,N_20409);
or U22134 (N_22134,N_20199,N_20237);
or U22135 (N_22135,N_20957,N_20716);
and U22136 (N_22136,N_20853,N_20333);
and U22137 (N_22137,N_20210,N_20113);
xnor U22138 (N_22138,N_20955,N_20114);
nor U22139 (N_22139,N_20988,N_20970);
xor U22140 (N_22140,N_20255,N_20044);
or U22141 (N_22141,N_21045,N_20576);
and U22142 (N_22142,N_20641,N_20786);
nand U22143 (N_22143,N_20381,N_20997);
xor U22144 (N_22144,N_20317,N_20372);
or U22145 (N_22145,N_20020,N_20750);
or U22146 (N_22146,N_20233,N_21034);
or U22147 (N_22147,N_20074,N_20006);
nand U22148 (N_22148,N_20556,N_20235);
xnor U22149 (N_22149,N_20540,N_20693);
nand U22150 (N_22150,N_20309,N_20413);
nor U22151 (N_22151,N_20282,N_20941);
nand U22152 (N_22152,N_20667,N_20621);
nor U22153 (N_22153,N_20932,N_20568);
xnor U22154 (N_22154,N_20584,N_20742);
and U22155 (N_22155,N_20196,N_20002);
nand U22156 (N_22156,N_20142,N_20586);
nand U22157 (N_22157,N_20845,N_20129);
nand U22158 (N_22158,N_21123,N_20933);
or U22159 (N_22159,N_21004,N_20764);
xor U22160 (N_22160,N_20936,N_20198);
xnor U22161 (N_22161,N_20988,N_20474);
and U22162 (N_22162,N_20132,N_20767);
or U22163 (N_22163,N_21088,N_20582);
nand U22164 (N_22164,N_20943,N_20107);
nand U22165 (N_22165,N_20715,N_21160);
nor U22166 (N_22166,N_20159,N_20817);
nand U22167 (N_22167,N_21229,N_20519);
nor U22168 (N_22168,N_20512,N_20353);
or U22169 (N_22169,N_20643,N_21212);
xnor U22170 (N_22170,N_20698,N_20892);
and U22171 (N_22171,N_21030,N_21029);
nand U22172 (N_22172,N_21114,N_20805);
or U22173 (N_22173,N_20493,N_20261);
or U22174 (N_22174,N_20918,N_20302);
or U22175 (N_22175,N_20257,N_20589);
xor U22176 (N_22176,N_21087,N_20059);
nand U22177 (N_22177,N_20738,N_20508);
nand U22178 (N_22178,N_20502,N_20458);
xor U22179 (N_22179,N_21106,N_20426);
or U22180 (N_22180,N_21005,N_20714);
nor U22181 (N_22181,N_20574,N_20837);
xor U22182 (N_22182,N_21038,N_20759);
nand U22183 (N_22183,N_20390,N_21139);
nor U22184 (N_22184,N_20878,N_21054);
nand U22185 (N_22185,N_21035,N_20929);
xor U22186 (N_22186,N_21029,N_20576);
xor U22187 (N_22187,N_21084,N_20287);
or U22188 (N_22188,N_20261,N_20244);
nand U22189 (N_22189,N_20206,N_21197);
and U22190 (N_22190,N_20403,N_21139);
nand U22191 (N_22191,N_20160,N_21190);
and U22192 (N_22192,N_20344,N_21085);
xnor U22193 (N_22193,N_21021,N_21048);
nor U22194 (N_22194,N_21189,N_20760);
xor U22195 (N_22195,N_21101,N_20559);
xor U22196 (N_22196,N_21003,N_20832);
and U22197 (N_22197,N_20884,N_20232);
nor U22198 (N_22198,N_20786,N_20561);
or U22199 (N_22199,N_20790,N_20210);
and U22200 (N_22200,N_20439,N_20365);
nor U22201 (N_22201,N_20729,N_20473);
and U22202 (N_22202,N_20268,N_20959);
xnor U22203 (N_22203,N_20290,N_20015);
nand U22204 (N_22204,N_20920,N_20634);
nor U22205 (N_22205,N_20347,N_20014);
or U22206 (N_22206,N_20034,N_20687);
nand U22207 (N_22207,N_20413,N_20696);
nand U22208 (N_22208,N_20419,N_20614);
nand U22209 (N_22209,N_20661,N_20847);
and U22210 (N_22210,N_21067,N_20443);
or U22211 (N_22211,N_20695,N_20511);
xor U22212 (N_22212,N_20793,N_20734);
nor U22213 (N_22213,N_20549,N_21177);
nor U22214 (N_22214,N_21125,N_20894);
nand U22215 (N_22215,N_20530,N_20511);
nor U22216 (N_22216,N_20914,N_20536);
and U22217 (N_22217,N_20940,N_20539);
xor U22218 (N_22218,N_20122,N_20058);
or U22219 (N_22219,N_20301,N_20216);
and U22220 (N_22220,N_20037,N_20621);
nand U22221 (N_22221,N_21239,N_20801);
xnor U22222 (N_22222,N_21047,N_21204);
and U22223 (N_22223,N_20966,N_20400);
nand U22224 (N_22224,N_21002,N_20006);
xnor U22225 (N_22225,N_20342,N_20986);
or U22226 (N_22226,N_21024,N_20141);
nor U22227 (N_22227,N_20523,N_20152);
xor U22228 (N_22228,N_20229,N_20491);
and U22229 (N_22229,N_20741,N_20553);
nor U22230 (N_22230,N_20605,N_20280);
and U22231 (N_22231,N_20724,N_20937);
xnor U22232 (N_22232,N_20343,N_21079);
xor U22233 (N_22233,N_20995,N_20406);
and U22234 (N_22234,N_21042,N_20863);
and U22235 (N_22235,N_20448,N_20409);
nor U22236 (N_22236,N_20945,N_20048);
or U22237 (N_22237,N_20909,N_20051);
or U22238 (N_22238,N_20224,N_21052);
nor U22239 (N_22239,N_20299,N_21195);
nor U22240 (N_22240,N_21097,N_20348);
xor U22241 (N_22241,N_20134,N_20853);
or U22242 (N_22242,N_20164,N_20791);
nor U22243 (N_22243,N_21111,N_20997);
nor U22244 (N_22244,N_20137,N_20813);
or U22245 (N_22245,N_21167,N_20583);
xnor U22246 (N_22246,N_20604,N_20992);
nor U22247 (N_22247,N_20920,N_20886);
nor U22248 (N_22248,N_20659,N_21060);
xor U22249 (N_22249,N_20375,N_21219);
or U22250 (N_22250,N_20485,N_20763);
xor U22251 (N_22251,N_20229,N_20706);
nand U22252 (N_22252,N_20918,N_21036);
or U22253 (N_22253,N_20011,N_20932);
nor U22254 (N_22254,N_20762,N_20428);
and U22255 (N_22255,N_20512,N_20896);
and U22256 (N_22256,N_21061,N_20156);
nand U22257 (N_22257,N_20949,N_21137);
or U22258 (N_22258,N_20448,N_20201);
xnor U22259 (N_22259,N_21033,N_21128);
xnor U22260 (N_22260,N_20789,N_20919);
nor U22261 (N_22261,N_20776,N_20695);
xnor U22262 (N_22262,N_20592,N_20771);
and U22263 (N_22263,N_21204,N_20040);
or U22264 (N_22264,N_20447,N_20608);
and U22265 (N_22265,N_20475,N_20908);
nand U22266 (N_22266,N_20339,N_21001);
or U22267 (N_22267,N_20954,N_20831);
xor U22268 (N_22268,N_20733,N_20481);
nand U22269 (N_22269,N_20380,N_21135);
and U22270 (N_22270,N_21024,N_21009);
xor U22271 (N_22271,N_20298,N_20659);
or U22272 (N_22272,N_20360,N_21085);
nand U22273 (N_22273,N_20641,N_21030);
xnor U22274 (N_22274,N_21032,N_20278);
xnor U22275 (N_22275,N_20667,N_20647);
xnor U22276 (N_22276,N_20817,N_20967);
nor U22277 (N_22277,N_20417,N_20026);
xnor U22278 (N_22278,N_20973,N_20883);
xnor U22279 (N_22279,N_20077,N_20463);
xnor U22280 (N_22280,N_20546,N_20115);
or U22281 (N_22281,N_20676,N_20787);
and U22282 (N_22282,N_20045,N_20979);
or U22283 (N_22283,N_20293,N_20222);
nand U22284 (N_22284,N_21038,N_20225);
or U22285 (N_22285,N_21209,N_20222);
or U22286 (N_22286,N_21215,N_21238);
xor U22287 (N_22287,N_20141,N_20824);
xor U22288 (N_22288,N_20269,N_21222);
xor U22289 (N_22289,N_20098,N_20048);
nand U22290 (N_22290,N_20540,N_20032);
or U22291 (N_22291,N_20875,N_20331);
nand U22292 (N_22292,N_20636,N_20215);
and U22293 (N_22293,N_20235,N_20234);
or U22294 (N_22294,N_20263,N_20272);
or U22295 (N_22295,N_20232,N_20817);
nor U22296 (N_22296,N_20303,N_20213);
and U22297 (N_22297,N_20971,N_20713);
and U22298 (N_22298,N_20855,N_20838);
and U22299 (N_22299,N_20472,N_20780);
nand U22300 (N_22300,N_21097,N_21089);
xnor U22301 (N_22301,N_20970,N_20558);
or U22302 (N_22302,N_20316,N_20848);
and U22303 (N_22303,N_20200,N_21115);
nor U22304 (N_22304,N_20360,N_20408);
xor U22305 (N_22305,N_20830,N_21190);
or U22306 (N_22306,N_20448,N_20847);
nor U22307 (N_22307,N_20494,N_20803);
nor U22308 (N_22308,N_20434,N_20792);
xor U22309 (N_22309,N_20084,N_20799);
nor U22310 (N_22310,N_21073,N_20574);
xor U22311 (N_22311,N_21243,N_20763);
nor U22312 (N_22312,N_20406,N_20342);
nor U22313 (N_22313,N_20888,N_20033);
and U22314 (N_22314,N_20449,N_20882);
and U22315 (N_22315,N_20624,N_20078);
nand U22316 (N_22316,N_20354,N_20934);
nor U22317 (N_22317,N_20148,N_21220);
and U22318 (N_22318,N_20893,N_20404);
and U22319 (N_22319,N_21133,N_20865);
nand U22320 (N_22320,N_21213,N_20011);
or U22321 (N_22321,N_20911,N_20106);
xor U22322 (N_22322,N_21129,N_21152);
nor U22323 (N_22323,N_20710,N_20205);
nor U22324 (N_22324,N_20488,N_20516);
and U22325 (N_22325,N_20368,N_20627);
and U22326 (N_22326,N_20445,N_20869);
nand U22327 (N_22327,N_20789,N_20849);
nand U22328 (N_22328,N_21053,N_20976);
nor U22329 (N_22329,N_20001,N_20713);
xnor U22330 (N_22330,N_20493,N_20786);
nand U22331 (N_22331,N_20153,N_20527);
or U22332 (N_22332,N_20671,N_20273);
or U22333 (N_22333,N_21138,N_20525);
nor U22334 (N_22334,N_20826,N_20905);
and U22335 (N_22335,N_20234,N_21219);
or U22336 (N_22336,N_20440,N_20072);
xnor U22337 (N_22337,N_21086,N_21203);
or U22338 (N_22338,N_21170,N_20466);
nand U22339 (N_22339,N_21049,N_20512);
xnor U22340 (N_22340,N_21148,N_20161);
xor U22341 (N_22341,N_21122,N_20606);
nand U22342 (N_22342,N_20144,N_20448);
and U22343 (N_22343,N_20297,N_20071);
and U22344 (N_22344,N_20135,N_21184);
nand U22345 (N_22345,N_20689,N_20032);
or U22346 (N_22346,N_20901,N_20681);
or U22347 (N_22347,N_20675,N_20451);
xor U22348 (N_22348,N_20759,N_21099);
and U22349 (N_22349,N_20528,N_21003);
xnor U22350 (N_22350,N_20464,N_21188);
nand U22351 (N_22351,N_21188,N_20580);
or U22352 (N_22352,N_20839,N_20785);
and U22353 (N_22353,N_21030,N_20805);
and U22354 (N_22354,N_20328,N_21032);
and U22355 (N_22355,N_21162,N_20550);
and U22356 (N_22356,N_20910,N_21165);
xnor U22357 (N_22357,N_20573,N_20755);
nand U22358 (N_22358,N_20925,N_20036);
nand U22359 (N_22359,N_20828,N_20072);
xor U22360 (N_22360,N_20007,N_21169);
xnor U22361 (N_22361,N_20693,N_20279);
and U22362 (N_22362,N_20134,N_20320);
or U22363 (N_22363,N_20668,N_20537);
xnor U22364 (N_22364,N_20897,N_21045);
nor U22365 (N_22365,N_21214,N_20696);
xnor U22366 (N_22366,N_21042,N_20804);
and U22367 (N_22367,N_20149,N_20831);
nand U22368 (N_22368,N_20020,N_20077);
or U22369 (N_22369,N_21180,N_20036);
nor U22370 (N_22370,N_20661,N_21028);
xor U22371 (N_22371,N_20395,N_20954);
xnor U22372 (N_22372,N_20158,N_21132);
nor U22373 (N_22373,N_21134,N_20887);
nor U22374 (N_22374,N_21065,N_20516);
nor U22375 (N_22375,N_20958,N_20925);
or U22376 (N_22376,N_20521,N_20433);
and U22377 (N_22377,N_20244,N_20520);
xnor U22378 (N_22378,N_21175,N_20418);
and U22379 (N_22379,N_21047,N_20539);
and U22380 (N_22380,N_20613,N_20725);
or U22381 (N_22381,N_20405,N_21222);
nor U22382 (N_22382,N_20625,N_20302);
xnor U22383 (N_22383,N_20255,N_20458);
nand U22384 (N_22384,N_20884,N_21119);
nor U22385 (N_22385,N_20854,N_20608);
nand U22386 (N_22386,N_21111,N_21165);
and U22387 (N_22387,N_20777,N_20749);
xor U22388 (N_22388,N_21131,N_20659);
xnor U22389 (N_22389,N_21058,N_20698);
xor U22390 (N_22390,N_20505,N_20038);
nand U22391 (N_22391,N_20907,N_20452);
nand U22392 (N_22392,N_20649,N_20844);
or U22393 (N_22393,N_20745,N_20124);
and U22394 (N_22394,N_20390,N_20631);
nand U22395 (N_22395,N_20119,N_20522);
xnor U22396 (N_22396,N_20173,N_21234);
nand U22397 (N_22397,N_20095,N_20866);
xor U22398 (N_22398,N_20896,N_21249);
or U22399 (N_22399,N_21110,N_20392);
nor U22400 (N_22400,N_20412,N_20249);
nand U22401 (N_22401,N_20510,N_20309);
nand U22402 (N_22402,N_20481,N_20755);
nand U22403 (N_22403,N_20062,N_20383);
or U22404 (N_22404,N_20242,N_20978);
nand U22405 (N_22405,N_21012,N_21000);
nor U22406 (N_22406,N_20265,N_20184);
nand U22407 (N_22407,N_20332,N_20616);
nand U22408 (N_22408,N_20922,N_20366);
and U22409 (N_22409,N_20136,N_20906);
and U22410 (N_22410,N_20896,N_20824);
or U22411 (N_22411,N_21147,N_20987);
nor U22412 (N_22412,N_20508,N_20558);
xnor U22413 (N_22413,N_21000,N_20087);
nand U22414 (N_22414,N_20852,N_21231);
xnor U22415 (N_22415,N_20540,N_20164);
or U22416 (N_22416,N_20028,N_21159);
or U22417 (N_22417,N_20304,N_20570);
or U22418 (N_22418,N_20410,N_21162);
and U22419 (N_22419,N_20671,N_20647);
and U22420 (N_22420,N_21027,N_21043);
xor U22421 (N_22421,N_21004,N_20796);
xor U22422 (N_22422,N_21206,N_20739);
xnor U22423 (N_22423,N_20708,N_20635);
and U22424 (N_22424,N_20715,N_20336);
xnor U22425 (N_22425,N_20211,N_20726);
xnor U22426 (N_22426,N_21021,N_20108);
nor U22427 (N_22427,N_20414,N_20902);
nand U22428 (N_22428,N_21143,N_21126);
nor U22429 (N_22429,N_20072,N_20375);
and U22430 (N_22430,N_21120,N_20495);
xnor U22431 (N_22431,N_20833,N_20787);
nor U22432 (N_22432,N_20683,N_20447);
nand U22433 (N_22433,N_20119,N_20056);
or U22434 (N_22434,N_21087,N_20464);
or U22435 (N_22435,N_20104,N_20572);
nor U22436 (N_22436,N_21247,N_20261);
and U22437 (N_22437,N_20685,N_21207);
nand U22438 (N_22438,N_20456,N_20270);
nand U22439 (N_22439,N_21038,N_20435);
nand U22440 (N_22440,N_20088,N_20585);
nor U22441 (N_22441,N_21180,N_20746);
or U22442 (N_22442,N_20455,N_20130);
nand U22443 (N_22443,N_20689,N_20562);
nand U22444 (N_22444,N_20703,N_20095);
nand U22445 (N_22445,N_20505,N_20269);
nand U22446 (N_22446,N_20545,N_20141);
nor U22447 (N_22447,N_20545,N_20154);
or U22448 (N_22448,N_20113,N_20832);
and U22449 (N_22449,N_20157,N_20732);
nor U22450 (N_22450,N_20963,N_20996);
and U22451 (N_22451,N_20548,N_21121);
or U22452 (N_22452,N_20001,N_20278);
and U22453 (N_22453,N_20095,N_20362);
or U22454 (N_22454,N_20719,N_21114);
xor U22455 (N_22455,N_20663,N_20593);
nor U22456 (N_22456,N_20343,N_20360);
nor U22457 (N_22457,N_20370,N_20204);
xnor U22458 (N_22458,N_20256,N_20242);
nand U22459 (N_22459,N_20674,N_20097);
or U22460 (N_22460,N_20341,N_20417);
nand U22461 (N_22461,N_20083,N_21214);
xnor U22462 (N_22462,N_20432,N_20013);
xnor U22463 (N_22463,N_20422,N_20800);
xnor U22464 (N_22464,N_21007,N_20145);
nand U22465 (N_22465,N_21234,N_20787);
nor U22466 (N_22466,N_20550,N_20013);
nor U22467 (N_22467,N_20621,N_21239);
or U22468 (N_22468,N_20278,N_20969);
nor U22469 (N_22469,N_20748,N_20230);
and U22470 (N_22470,N_20502,N_20622);
xnor U22471 (N_22471,N_20124,N_20699);
nand U22472 (N_22472,N_20466,N_21109);
xor U22473 (N_22473,N_20914,N_20463);
xnor U22474 (N_22474,N_20018,N_21094);
or U22475 (N_22475,N_20475,N_21080);
nand U22476 (N_22476,N_20528,N_20074);
or U22477 (N_22477,N_20681,N_20179);
or U22478 (N_22478,N_20249,N_20966);
or U22479 (N_22479,N_20895,N_20824);
and U22480 (N_22480,N_21055,N_20648);
nand U22481 (N_22481,N_20678,N_20023);
or U22482 (N_22482,N_20604,N_20593);
nor U22483 (N_22483,N_20982,N_20377);
xnor U22484 (N_22484,N_20757,N_21009);
or U22485 (N_22485,N_20528,N_20115);
nand U22486 (N_22486,N_20069,N_20030);
nand U22487 (N_22487,N_21221,N_20849);
nor U22488 (N_22488,N_20293,N_20689);
nand U22489 (N_22489,N_20189,N_21216);
nand U22490 (N_22490,N_20459,N_20435);
nor U22491 (N_22491,N_20097,N_20322);
nand U22492 (N_22492,N_20757,N_20732);
xor U22493 (N_22493,N_20750,N_20743);
and U22494 (N_22494,N_20499,N_20075);
nand U22495 (N_22495,N_20018,N_20244);
xor U22496 (N_22496,N_20606,N_20411);
nor U22497 (N_22497,N_20476,N_20057);
and U22498 (N_22498,N_20520,N_20248);
nand U22499 (N_22499,N_20927,N_20973);
nand U22500 (N_22500,N_22045,N_22070);
nor U22501 (N_22501,N_22318,N_22341);
and U22502 (N_22502,N_21941,N_21712);
or U22503 (N_22503,N_22424,N_22368);
and U22504 (N_22504,N_21441,N_21393);
nor U22505 (N_22505,N_22384,N_21311);
or U22506 (N_22506,N_22118,N_21748);
and U22507 (N_22507,N_21260,N_22097);
nand U22508 (N_22508,N_21648,N_21438);
and U22509 (N_22509,N_21733,N_22495);
or U22510 (N_22510,N_22272,N_21873);
and U22511 (N_22511,N_22480,N_22254);
nor U22512 (N_22512,N_22081,N_21286);
nand U22513 (N_22513,N_21863,N_21284);
or U22514 (N_22514,N_21854,N_21650);
nor U22515 (N_22515,N_21993,N_21930);
and U22516 (N_22516,N_21497,N_21932);
or U22517 (N_22517,N_22294,N_22449);
or U22518 (N_22518,N_21995,N_21295);
and U22519 (N_22519,N_22265,N_22134);
nand U22520 (N_22520,N_22052,N_22270);
nand U22521 (N_22521,N_22478,N_21399);
nand U22522 (N_22522,N_22428,N_21395);
and U22523 (N_22523,N_21695,N_21546);
xor U22524 (N_22524,N_21798,N_21988);
or U22525 (N_22525,N_22435,N_22320);
and U22526 (N_22526,N_22119,N_21455);
xnor U22527 (N_22527,N_21836,N_22337);
nor U22528 (N_22528,N_22485,N_21338);
nor U22529 (N_22529,N_22240,N_22359);
and U22530 (N_22530,N_21453,N_22315);
xor U22531 (N_22531,N_21264,N_22444);
nor U22532 (N_22532,N_21968,N_22126);
nand U22533 (N_22533,N_21850,N_21586);
nand U22534 (N_22534,N_22417,N_21825);
nand U22535 (N_22535,N_22021,N_22044);
nand U22536 (N_22536,N_22441,N_21525);
or U22537 (N_22537,N_22105,N_22224);
nor U22538 (N_22538,N_21406,N_22128);
nand U22539 (N_22539,N_21711,N_21339);
and U22540 (N_22540,N_21686,N_21560);
or U22541 (N_22541,N_21547,N_22187);
and U22542 (N_22542,N_21327,N_21769);
and U22543 (N_22543,N_22088,N_21565);
and U22544 (N_22544,N_21449,N_22192);
nor U22545 (N_22545,N_22396,N_21529);
nor U22546 (N_22546,N_21583,N_22403);
or U22547 (N_22547,N_21346,N_21394);
nor U22548 (N_22548,N_22133,N_21559);
and U22549 (N_22549,N_22189,N_22141);
nand U22550 (N_22550,N_21544,N_21580);
or U22551 (N_22551,N_22271,N_22380);
nor U22552 (N_22552,N_21978,N_21548);
and U22553 (N_22553,N_21690,N_22106);
nor U22554 (N_22554,N_22082,N_21920);
or U22555 (N_22555,N_21813,N_21640);
or U22556 (N_22556,N_21635,N_21591);
xnor U22557 (N_22557,N_21288,N_21549);
or U22558 (N_22558,N_21313,N_22237);
and U22559 (N_22559,N_21522,N_22350);
and U22560 (N_22560,N_22139,N_21613);
or U22561 (N_22561,N_22220,N_22232);
nand U22562 (N_22562,N_21957,N_21922);
xor U22563 (N_22563,N_21402,N_21875);
nor U22564 (N_22564,N_21259,N_22029);
nor U22565 (N_22565,N_21360,N_22094);
or U22566 (N_22566,N_22353,N_21716);
nand U22567 (N_22567,N_21723,N_21964);
or U22568 (N_22568,N_21936,N_22217);
nand U22569 (N_22569,N_21507,N_21514);
nand U22570 (N_22570,N_22140,N_22412);
nor U22571 (N_22571,N_22074,N_21958);
nor U22572 (N_22572,N_22297,N_21664);
xor U22573 (N_22573,N_22223,N_22303);
nand U22574 (N_22574,N_22479,N_21676);
or U22575 (N_22575,N_22323,N_22429);
xor U22576 (N_22576,N_21281,N_22159);
nand U22577 (N_22577,N_22282,N_22103);
nor U22578 (N_22578,N_21483,N_22151);
nor U22579 (N_22579,N_22028,N_21280);
or U22580 (N_22580,N_22110,N_22226);
xnor U22581 (N_22581,N_21779,N_21600);
xnor U22582 (N_22582,N_22124,N_22132);
or U22583 (N_22583,N_21786,N_21643);
or U22584 (N_22584,N_21762,N_21715);
nand U22585 (N_22585,N_21476,N_22243);
or U22586 (N_22586,N_21421,N_22002);
nor U22587 (N_22587,N_22431,N_21979);
nor U22588 (N_22588,N_22342,N_21835);
nor U22589 (N_22589,N_21261,N_21887);
nand U22590 (N_22590,N_21921,N_21322);
and U22591 (N_22591,N_21305,N_21361);
nor U22592 (N_22592,N_21963,N_21777);
nor U22593 (N_22593,N_21608,N_21253);
xnor U22594 (N_22594,N_21692,N_22459);
or U22595 (N_22595,N_22286,N_21975);
nand U22596 (N_22596,N_21597,N_21627);
xnor U22597 (N_22597,N_22125,N_21364);
nor U22598 (N_22598,N_21859,N_22392);
nand U22599 (N_22599,N_21300,N_22123);
and U22600 (N_22600,N_21869,N_21423);
nor U22601 (N_22601,N_21925,N_21734);
or U22602 (N_22602,N_21701,N_22014);
xor U22603 (N_22603,N_21403,N_21894);
and U22604 (N_22604,N_22379,N_21742);
and U22605 (N_22605,N_21458,N_21343);
and U22606 (N_22606,N_21636,N_22405);
nand U22607 (N_22607,N_22075,N_21381);
and U22608 (N_22608,N_22031,N_21900);
nand U22609 (N_22609,N_21362,N_22180);
or U22610 (N_22610,N_22206,N_22114);
nand U22611 (N_22611,N_22036,N_22229);
nor U22612 (N_22612,N_21951,N_21982);
and U22613 (N_22613,N_22461,N_21299);
nand U22614 (N_22614,N_21658,N_22190);
or U22615 (N_22615,N_22212,N_21707);
and U22616 (N_22616,N_22312,N_21397);
or U22617 (N_22617,N_22207,N_21290);
or U22618 (N_22618,N_21782,N_21326);
nor U22619 (N_22619,N_21749,N_21689);
or U22620 (N_22620,N_21384,N_22016);
or U22621 (N_22621,N_22457,N_22344);
and U22622 (N_22622,N_22161,N_21639);
and U22623 (N_22623,N_21916,N_21902);
and U22624 (N_22624,N_21289,N_21509);
and U22625 (N_22625,N_21751,N_22409);
or U22626 (N_22626,N_21845,N_22283);
nor U22627 (N_22627,N_21541,N_21294);
nand U22628 (N_22628,N_22108,N_21358);
nor U22629 (N_22629,N_22005,N_21839);
xor U22630 (N_22630,N_21917,N_21759);
nor U22631 (N_22631,N_21886,N_22292);
and U22632 (N_22632,N_21575,N_21466);
xor U22633 (N_22633,N_21410,N_21841);
or U22634 (N_22634,N_21444,N_22084);
xor U22635 (N_22635,N_21878,N_22136);
and U22636 (N_22636,N_22456,N_21770);
nand U22637 (N_22637,N_22474,N_22242);
and U22638 (N_22638,N_21536,N_22117);
xor U22639 (N_22639,N_21756,N_21699);
or U22640 (N_22640,N_21852,N_21436);
nor U22641 (N_22641,N_21537,N_21414);
and U22642 (N_22642,N_21459,N_21931);
nand U22643 (N_22643,N_21587,N_22410);
nor U22644 (N_22644,N_22169,N_22493);
and U22645 (N_22645,N_22146,N_21771);
xor U22646 (N_22646,N_22238,N_22176);
xor U22647 (N_22647,N_21735,N_21484);
nand U22648 (N_22648,N_22372,N_21687);
nor U22649 (N_22649,N_21793,N_22404);
or U22650 (N_22650,N_22481,N_22277);
and U22651 (N_22651,N_21903,N_21523);
nand U22652 (N_22652,N_21604,N_21721);
xor U22653 (N_22653,N_21528,N_21746);
and U22654 (N_22654,N_21325,N_21334);
nand U22655 (N_22655,N_22090,N_21611);
nor U22656 (N_22656,N_21959,N_21685);
nand U22657 (N_22657,N_21888,N_21494);
or U22658 (N_22658,N_21316,N_22038);
and U22659 (N_22659,N_21336,N_21697);
or U22660 (N_22660,N_21367,N_21871);
nand U22661 (N_22661,N_22400,N_21610);
xor U22662 (N_22662,N_21969,N_22087);
or U22663 (N_22663,N_21987,N_22445);
or U22664 (N_22664,N_22200,N_21574);
nor U22665 (N_22665,N_21630,N_22421);
xnor U22666 (N_22666,N_21601,N_22371);
xor U22667 (N_22667,N_22390,N_21981);
or U22668 (N_22668,N_22023,N_22017);
xor U22669 (N_22669,N_21838,N_22316);
and U22670 (N_22670,N_21991,N_21614);
or U22671 (N_22671,N_21372,N_21652);
nand U22672 (N_22672,N_22058,N_22361);
or U22673 (N_22673,N_21628,N_21709);
or U22674 (N_22674,N_21961,N_21719);
or U22675 (N_22675,N_21732,N_21785);
nand U22676 (N_22676,N_22049,N_21463);
xnor U22677 (N_22677,N_22116,N_21933);
nor U22678 (N_22678,N_21815,N_21858);
nand U22679 (N_22679,N_21764,N_21829);
and U22680 (N_22680,N_21542,N_22386);
and U22681 (N_22681,N_21772,N_22195);
xor U22682 (N_22682,N_22280,N_22309);
nand U22683 (N_22683,N_22263,N_22347);
nand U22684 (N_22684,N_22009,N_21532);
nor U22685 (N_22685,N_21504,N_21910);
xnor U22686 (N_22686,N_22436,N_21892);
nor U22687 (N_22687,N_22250,N_21940);
nor U22688 (N_22688,N_21739,N_22067);
and U22689 (N_22689,N_21434,N_21267);
and U22690 (N_22690,N_21582,N_22137);
nor U22691 (N_22691,N_22443,N_22402);
and U22692 (N_22692,N_21743,N_21807);
xor U22693 (N_22693,N_21477,N_22113);
nor U22694 (N_22694,N_21866,N_22248);
nor U22695 (N_22695,N_22162,N_21857);
xor U22696 (N_22696,N_21952,N_22198);
or U22697 (N_22697,N_21501,N_22092);
xor U22698 (N_22698,N_21823,N_21446);
and U22699 (N_22699,N_21589,N_22202);
xnor U22700 (N_22700,N_22334,N_21622);
and U22701 (N_22701,N_22324,N_22033);
nor U22702 (N_22702,N_21853,N_22246);
and U22703 (N_22703,N_22304,N_22155);
or U22704 (N_22704,N_22120,N_22471);
and U22705 (N_22705,N_21479,N_21268);
or U22706 (N_22706,N_22335,N_22231);
xnor U22707 (N_22707,N_22488,N_21669);
and U22708 (N_22708,N_21837,N_22227);
or U22709 (N_22709,N_21344,N_22184);
nor U22710 (N_22710,N_22260,N_22193);
and U22711 (N_22711,N_21661,N_22111);
xor U22712 (N_22712,N_21561,N_21847);
nor U22713 (N_22713,N_22487,N_21820);
nand U22714 (N_22714,N_21708,N_22467);
xnor U22715 (N_22715,N_22152,N_21439);
and U22716 (N_22716,N_22022,N_21623);
and U22717 (N_22717,N_21277,N_22325);
xor U22718 (N_22718,N_21505,N_21893);
xnor U22719 (N_22719,N_21896,N_21263);
nor U22720 (N_22720,N_21330,N_21655);
or U22721 (N_22721,N_21255,N_21320);
and U22722 (N_22722,N_21555,N_21578);
nor U22723 (N_22723,N_21520,N_22095);
and U22724 (N_22724,N_22285,N_21365);
and U22725 (N_22725,N_22245,N_22486);
xor U22726 (N_22726,N_21703,N_21727);
nor U22727 (N_22727,N_22030,N_22298);
nor U22728 (N_22728,N_21947,N_21949);
nand U22729 (N_22729,N_22149,N_21323);
nor U22730 (N_22730,N_22210,N_21867);
xor U22731 (N_22731,N_21341,N_22196);
or U22732 (N_22732,N_21673,N_22369);
nand U22733 (N_22733,N_21375,N_21803);
nand U22734 (N_22734,N_22153,N_21832);
xor U22735 (N_22735,N_22476,N_21674);
or U22736 (N_22736,N_21496,N_21706);
nand U22737 (N_22737,N_21447,N_22004);
and U22738 (N_22738,N_21659,N_21513);
nor U22739 (N_22739,N_21366,N_22469);
nand U22740 (N_22740,N_21297,N_21763);
and U22741 (N_22741,N_21812,N_22276);
or U22742 (N_22742,N_22219,N_21452);
xor U22743 (N_22743,N_22043,N_21448);
xnor U22744 (N_22744,N_22145,N_21480);
or U22745 (N_22745,N_21368,N_21524);
nand U22746 (N_22746,N_21595,N_22354);
nor U22747 (N_22747,N_21870,N_21306);
or U22748 (N_22748,N_21303,N_22351);
xor U22749 (N_22749,N_21332,N_22258);
xnor U22750 (N_22750,N_21543,N_22266);
and U22751 (N_22751,N_21570,N_22062);
and U22752 (N_22752,N_22050,N_21353);
xnor U22753 (N_22753,N_22267,N_21607);
nor U22754 (N_22754,N_21262,N_21943);
and U22755 (N_22755,N_22378,N_22374);
xnor U22756 (N_22756,N_22496,N_22305);
or U22757 (N_22757,N_22201,N_22208);
nand U22758 (N_22758,N_21540,N_21319);
or U22759 (N_22759,N_22348,N_21956);
nor U22760 (N_22760,N_22452,N_22173);
xnor U22761 (N_22761,N_21654,N_21495);
nor U22762 (N_22762,N_22046,N_22364);
and U22763 (N_22763,N_22458,N_21817);
or U22764 (N_22764,N_21577,N_21412);
nand U22765 (N_22765,N_21626,N_21398);
and U22766 (N_22766,N_21539,N_22089);
nor U22767 (N_22767,N_22253,N_22446);
and U22768 (N_22768,N_22131,N_21774);
xnor U22769 (N_22769,N_21405,N_21273);
xor U22770 (N_22770,N_22321,N_21791);
nor U22771 (N_22771,N_21533,N_21806);
nor U22772 (N_22772,N_21800,N_21666);
or U22773 (N_22773,N_21848,N_22453);
nor U22774 (N_22774,N_21919,N_21876);
xnor U22775 (N_22775,N_21389,N_21445);
or U22776 (N_22776,N_21554,N_22419);
and U22777 (N_22777,N_21909,N_22440);
xnor U22778 (N_22778,N_22274,N_22408);
or U22779 (N_22779,N_21581,N_21265);
or U22780 (N_22780,N_22389,N_21474);
and U22781 (N_22781,N_22104,N_21811);
xnor U22782 (N_22782,N_22163,N_22057);
nor U22783 (N_22783,N_21747,N_22204);
and U22784 (N_22784,N_22415,N_22313);
or U22785 (N_22785,N_21293,N_22096);
and U22786 (N_22786,N_22352,N_21517);
nor U22787 (N_22787,N_21973,N_22255);
nand U22788 (N_22788,N_21795,N_22437);
xor U22789 (N_22789,N_22291,N_21741);
xnor U22790 (N_22790,N_22194,N_21730);
or U22791 (N_22791,N_21391,N_21783);
nor U22792 (N_22792,N_22182,N_22156);
xnor U22793 (N_22793,N_21967,N_21307);
xor U22794 (N_22794,N_21482,N_21766);
nor U22795 (N_22795,N_22426,N_21461);
and U22796 (N_22796,N_21616,N_21884);
nor U22797 (N_22797,N_22393,N_22477);
and U22798 (N_22798,N_22284,N_22042);
or U22799 (N_22799,N_22470,N_21799);
and U22800 (N_22800,N_21849,N_21714);
or U22801 (N_22801,N_22071,N_21621);
or U22802 (N_22802,N_22383,N_22222);
or U22803 (N_22803,N_21998,N_22239);
xor U22804 (N_22804,N_22262,N_22019);
nand U22805 (N_22805,N_22215,N_21258);
and U22806 (N_22806,N_22244,N_21726);
nor U22807 (N_22807,N_21442,N_21424);
and U22808 (N_22808,N_22358,N_21374);
or U22809 (N_22809,N_21725,N_21752);
nor U22810 (N_22810,N_21939,N_21370);
or U22811 (N_22811,N_21913,N_21645);
or U22812 (N_22812,N_21906,N_21328);
and U22813 (N_22813,N_21252,N_22295);
nor U22814 (N_22814,N_22015,N_22185);
or U22815 (N_22815,N_22264,N_21926);
xnor U22816 (N_22816,N_21457,N_21702);
or U22817 (N_22817,N_22366,N_21790);
and U22818 (N_22818,N_21912,N_22491);
nand U22819 (N_22819,N_21373,N_22073);
nor U22820 (N_22820,N_21638,N_21983);
nor U22821 (N_22821,N_21724,N_22241);
nand U22822 (N_22822,N_22279,N_21821);
nor U22823 (N_22823,N_21805,N_21422);
and U22824 (N_22824,N_21704,N_21437);
nand U22825 (N_22825,N_22330,N_22012);
and U22826 (N_22826,N_21301,N_21728);
xor U22827 (N_22827,N_21312,N_22010);
nor U22828 (N_22828,N_22439,N_22460);
xnor U22829 (N_22829,N_21787,N_21450);
nor U22830 (N_22830,N_21696,N_21451);
or U22831 (N_22831,N_21443,N_21460);
nor U22832 (N_22832,N_22115,N_21378);
or U22833 (N_22833,N_22080,N_21927);
or U22834 (N_22834,N_22235,N_21566);
or U22835 (N_22835,N_21499,N_21419);
and U22836 (N_22836,N_21433,N_21994);
xor U22837 (N_22837,N_21371,N_21409);
nor U22838 (N_22838,N_21590,N_22466);
or U22839 (N_22839,N_21997,N_22102);
nor U22840 (N_22840,N_22069,N_21773);
nand U22841 (N_22841,N_22332,N_22099);
or U22842 (N_22842,N_21500,N_22259);
and U22843 (N_22843,N_22112,N_22221);
nor U22844 (N_22844,N_21416,N_22154);
or U22845 (N_22845,N_22177,N_21429);
xnor U22846 (N_22846,N_22451,N_22473);
nand U22847 (N_22847,N_22026,N_22061);
and U22848 (N_22848,N_21526,N_21901);
and U22849 (N_22849,N_21472,N_22107);
nor U22850 (N_22850,N_21340,N_21681);
nor U22851 (N_22851,N_22209,N_21620);
or U22852 (N_22852,N_21283,N_22308);
and U22853 (N_22853,N_22310,N_22158);
or U22854 (N_22854,N_22365,N_21573);
nand U22855 (N_22855,N_22191,N_21737);
nor U22856 (N_22856,N_21950,N_21647);
nor U22857 (N_22857,N_22287,N_22455);
nor U22858 (N_22858,N_21274,N_21948);
nor U22859 (N_22859,N_21602,N_21700);
nand U22860 (N_22860,N_21382,N_21473);
nor U22861 (N_22861,N_22000,N_21625);
nand U22862 (N_22862,N_22385,N_22339);
and U22863 (N_22863,N_21953,N_21984);
nand U22864 (N_22864,N_21468,N_21464);
xor U22865 (N_22865,N_21637,N_22413);
nand U22866 (N_22866,N_22376,N_22065);
nand U22867 (N_22867,N_21462,N_22381);
nor U22868 (N_22868,N_21347,N_21584);
or U22869 (N_22869,N_21606,N_21485);
or U22870 (N_22870,N_21470,N_21745);
nor U22871 (N_22871,N_21804,N_22032);
nand U22872 (N_22872,N_21929,N_21872);
nand U22873 (N_22873,N_21996,N_21331);
and U22874 (N_22874,N_21415,N_22037);
or U22875 (N_22875,N_22234,N_21915);
nand U22876 (N_22876,N_21492,N_21302);
nand U22877 (N_22877,N_21683,N_21515);
and U22878 (N_22878,N_21914,N_22373);
nand U22879 (N_22879,N_21531,N_22482);
nor U22880 (N_22880,N_21562,N_21844);
and U22881 (N_22881,N_21989,N_21568);
nand U22882 (N_22882,N_21558,N_21599);
nor U22883 (N_22883,N_22174,N_22211);
xnor U22884 (N_22884,N_22175,N_22363);
and U22885 (N_22885,N_21855,N_22394);
xnor U22886 (N_22886,N_21380,N_21563);
nand U22887 (N_22887,N_21891,N_22498);
or U22888 (N_22888,N_22382,N_22472);
or U22889 (N_22889,N_21899,N_21808);
xor U22890 (N_22890,N_21435,N_22377);
nand U22891 (N_22891,N_22434,N_21842);
or U22892 (N_22892,N_21298,N_21335);
and U22893 (N_22893,N_21918,N_22047);
and U22894 (N_22894,N_22317,N_21407);
xnor U22895 (N_22895,N_22322,N_22468);
and U22896 (N_22896,N_22293,N_21516);
and U22897 (N_22897,N_21881,N_22367);
nor U22898 (N_22898,N_22340,N_21877);
nand U22899 (N_22899,N_21907,N_21675);
nand U22900 (N_22900,N_22003,N_21498);
xnor U22901 (N_22901,N_22236,N_22171);
nor U22902 (N_22902,N_22035,N_22414);
xor U22903 (N_22903,N_22462,N_22079);
or U22904 (N_22904,N_21355,N_22034);
or U22905 (N_22905,N_21310,N_21833);
or U22906 (N_22906,N_21481,N_21491);
and U22907 (N_22907,N_21809,N_21617);
nand U22908 (N_22908,N_21792,N_21720);
or U22909 (N_22909,N_21960,N_22233);
nor U22910 (N_22910,N_22039,N_21651);
or U22911 (N_22911,N_22343,N_22018);
and U22912 (N_22912,N_22051,N_21883);
nand U22913 (N_22913,N_21816,N_21388);
nand U22914 (N_22914,N_21275,N_21646);
or U22915 (N_22915,N_22432,N_21618);
and U22916 (N_22916,N_21801,N_22165);
or U22917 (N_22917,N_21634,N_21392);
nor U22918 (N_22918,N_22290,N_21889);
nand U22919 (N_22919,N_21831,N_22225);
nor U22920 (N_22920,N_21810,N_21944);
and U22921 (N_22921,N_22307,N_22370);
nor U22922 (N_22922,N_21612,N_21418);
xor U22923 (N_22923,N_22027,N_21430);
or U22924 (N_22924,N_21569,N_21677);
nor U22925 (N_22925,N_21999,N_22091);
and U22926 (N_22926,N_22060,N_21758);
xnor U22927 (N_22927,N_21588,N_22170);
nor U22928 (N_22928,N_21846,N_21649);
xnor U22929 (N_22929,N_21521,N_22213);
and U22930 (N_22930,N_21860,N_22416);
or U22931 (N_22931,N_21974,N_22406);
or U22932 (N_22932,N_22338,N_21408);
xnor U22933 (N_22933,N_21934,N_21354);
or U22934 (N_22934,N_22100,N_21924);
xnor U22935 (N_22935,N_22064,N_21928);
and U22936 (N_22936,N_21668,N_21309);
nand U22937 (N_22937,N_21624,N_21986);
xor U22938 (N_22938,N_22076,N_21778);
nor U22939 (N_22939,N_22122,N_21768);
or U22940 (N_22940,N_21722,N_22362);
nor U22941 (N_22941,N_22391,N_21456);
xnor U22942 (N_22942,N_22450,N_21256);
nor U22943 (N_22943,N_22066,N_21337);
nand U22944 (N_22944,N_22007,N_21885);
and U22945 (N_22945,N_22078,N_21400);
nand U22946 (N_22946,N_21880,N_22261);
xnor U22947 (N_22947,N_21557,N_22401);
or U22948 (N_22948,N_21576,N_21656);
xnor U22949 (N_22949,N_21665,N_21369);
xor U22950 (N_22950,N_21680,N_22001);
nand U22951 (N_22951,N_21551,N_21552);
or U22952 (N_22952,N_22388,N_21490);
or U22953 (N_22953,N_21396,N_21254);
or U22954 (N_22954,N_22300,N_22166);
nand U22955 (N_22955,N_21465,N_21644);
nand U22956 (N_22956,N_22179,N_21897);
nand U22957 (N_22957,N_21657,N_22072);
nand U22958 (N_22958,N_21511,N_21619);
xnor U22959 (N_22959,N_22167,N_22257);
xor U22960 (N_22960,N_21879,N_21342);
nand U22961 (N_22961,N_21304,N_21754);
nand U22962 (N_22962,N_21535,N_22138);
and U22963 (N_22963,N_22164,N_22181);
and U22964 (N_22964,N_22494,N_21753);
xor U22965 (N_22965,N_21527,N_22306);
or U22966 (N_22966,N_21486,N_21824);
xnor U22967 (N_22967,N_21670,N_21980);
nor U22968 (N_22968,N_21386,N_22127);
and U22969 (N_22969,N_21428,N_21882);
or U22970 (N_22970,N_22346,N_21615);
nor U22971 (N_22971,N_21672,N_21904);
and U22972 (N_22972,N_22142,N_22329);
nor U22973 (N_22973,N_21976,N_22463);
and U22974 (N_22974,N_21351,N_22454);
nor U22975 (N_22975,N_22020,N_22288);
nor U22976 (N_22976,N_21868,N_21510);
or U22977 (N_22977,N_21321,N_22144);
nand U22978 (N_22978,N_21861,N_22356);
nand U22979 (N_22979,N_21788,N_22448);
xor U22980 (N_22980,N_22251,N_22186);
and U22981 (N_22981,N_21518,N_22150);
xor U22982 (N_22982,N_22407,N_21270);
nor U22983 (N_22983,N_21761,N_21251);
or U22984 (N_22984,N_21572,N_21781);
nor U22985 (N_22985,N_22314,N_21740);
nor U22986 (N_22986,N_21970,N_21592);
nor U22987 (N_22987,N_21945,N_22275);
nand U22988 (N_22988,N_21818,N_22319);
nor U22989 (N_22989,N_21411,N_21478);
and U22990 (N_22990,N_21757,N_21315);
nor U22991 (N_22991,N_21667,N_21285);
and U22992 (N_22992,N_21318,N_21840);
nor U22993 (N_22993,N_21417,N_22497);
nand U22994 (N_22994,N_21596,N_22301);
nor U22995 (N_22995,N_21905,N_22214);
or U22996 (N_22996,N_21794,N_21363);
and U22997 (N_22997,N_21663,N_22077);
xnor U22998 (N_22998,N_21605,N_21985);
xnor U22999 (N_22999,N_22218,N_22135);
and U23000 (N_23000,N_21865,N_21556);
nor U23001 (N_23001,N_21938,N_22281);
nor U23002 (N_23002,N_22345,N_21349);
nor U23003 (N_23003,N_21705,N_22147);
and U23004 (N_23004,N_21890,N_22053);
xnor U23005 (N_23005,N_21296,N_21856);
or U23006 (N_23006,N_22484,N_21431);
and U23007 (N_23007,N_22422,N_22395);
nand U23008 (N_23008,N_21377,N_21534);
nand U23009 (N_23009,N_21350,N_21508);
xnor U23010 (N_23010,N_21851,N_22423);
or U23011 (N_23011,N_21862,N_21632);
nand U23012 (N_23012,N_21911,N_21356);
nand U23013 (N_23013,N_22121,N_22430);
xor U23014 (N_23014,N_22326,N_22357);
nand U23015 (N_23015,N_22296,N_21731);
and U23016 (N_23016,N_22269,N_22398);
xor U23017 (N_23017,N_22013,N_21834);
xnor U23018 (N_23018,N_21413,N_21895);
and U23019 (N_23019,N_21693,N_22205);
and U23020 (N_23020,N_21502,N_21710);
nor U23021 (N_23021,N_21401,N_22216);
xor U23022 (N_23022,N_21698,N_22328);
and U23023 (N_23023,N_21765,N_22054);
and U23024 (N_23024,N_21454,N_21308);
xor U23025 (N_23025,N_22499,N_21662);
xnor U23026 (N_23026,N_21519,N_21291);
and U23027 (N_23027,N_21935,N_22333);
nand U23028 (N_23028,N_22157,N_21488);
or U23029 (N_23029,N_22256,N_21642);
nor U23030 (N_23030,N_21688,N_22268);
nor U23031 (N_23031,N_21718,N_21329);
xor U23032 (N_23032,N_21977,N_22464);
nor U23033 (N_23033,N_22387,N_22433);
and U23034 (N_23034,N_21545,N_21828);
xnor U23035 (N_23035,N_22492,N_21660);
xnor U23036 (N_23036,N_21784,N_22129);
xor U23037 (N_23037,N_22349,N_21830);
nor U23038 (N_23038,N_21767,N_21603);
nand U23039 (N_23039,N_21276,N_21553);
nor U23040 (N_23040,N_21598,N_21631);
xnor U23041 (N_23041,N_22311,N_22041);
nand U23042 (N_23042,N_22199,N_21333);
xor U23043 (N_23043,N_21822,N_21420);
xnor U23044 (N_23044,N_22168,N_22278);
nor U23045 (N_23045,N_21387,N_22148);
or U23046 (N_23046,N_22101,N_21990);
nor U23047 (N_23047,N_21682,N_22475);
nor U23048 (N_23048,N_21279,N_22109);
nand U23049 (N_23049,N_22442,N_21946);
nor U23050 (N_23050,N_22063,N_21564);
nor U23051 (N_23051,N_21567,N_22068);
or U23052 (N_23052,N_21593,N_21629);
or U23053 (N_23053,N_21609,N_21489);
nor U23054 (N_23054,N_21348,N_21359);
nor U23055 (N_23055,N_21250,N_22427);
xnor U23056 (N_23056,N_21426,N_21898);
and U23057 (N_23057,N_21755,N_21471);
nand U23058 (N_23058,N_21512,N_21390);
nor U23059 (N_23059,N_22086,N_22399);
xnor U23060 (N_23060,N_21376,N_21671);
xnor U23061 (N_23061,N_22130,N_21972);
nor U23062 (N_23062,N_22420,N_21684);
nand U23063 (N_23063,N_21775,N_22024);
and U23064 (N_23064,N_21314,N_21923);
nand U23065 (N_23065,N_21345,N_22447);
nor U23066 (N_23066,N_22438,N_21467);
and U23067 (N_23067,N_22289,N_21404);
and U23068 (N_23068,N_22008,N_21955);
nand U23069 (N_23069,N_21469,N_21962);
nand U23070 (N_23070,N_22011,N_21780);
and U23071 (N_23071,N_22336,N_21550);
or U23072 (N_23072,N_22083,N_21379);
nor U23073 (N_23073,N_21257,N_21736);
nor U23074 (N_23074,N_21908,N_21760);
nor U23075 (N_23075,N_21475,N_22040);
or U23076 (N_23076,N_21653,N_21352);
and U23077 (N_23077,N_22252,N_21954);
xnor U23078 (N_23078,N_22397,N_21694);
nand U23079 (N_23079,N_22230,N_21750);
or U23080 (N_23080,N_21503,N_22197);
and U23081 (N_23081,N_22483,N_21942);
nand U23082 (N_23082,N_21287,N_21937);
nor U23083 (N_23083,N_22411,N_22172);
nand U23084 (N_23084,N_22056,N_22249);
nor U23085 (N_23085,N_21282,N_21425);
or U23086 (N_23086,N_21357,N_21324);
xor U23087 (N_23087,N_22355,N_21432);
xor U23088 (N_23088,N_22055,N_21965);
xnor U23089 (N_23089,N_22228,N_21802);
and U23090 (N_23090,N_22048,N_21966);
or U23091 (N_23091,N_21594,N_21738);
and U23092 (N_23092,N_22299,N_21530);
or U23093 (N_23093,N_21317,N_21679);
xnor U23094 (N_23094,N_21292,N_21691);
xor U23095 (N_23095,N_22006,N_22425);
nand U23096 (N_23096,N_22059,N_21789);
xnor U23097 (N_23097,N_21383,N_21971);
or U23098 (N_23098,N_21797,N_21571);
and U23099 (N_23099,N_21864,N_21678);
and U23100 (N_23100,N_22331,N_21843);
or U23101 (N_23101,N_21427,N_22273);
xor U23102 (N_23102,N_21992,N_22160);
nand U23103 (N_23103,N_21271,N_21278);
nand U23104 (N_23104,N_21269,N_22098);
nand U23105 (N_23105,N_21641,N_22302);
xor U23106 (N_23106,N_21487,N_22093);
nor U23107 (N_23107,N_22490,N_21827);
or U23108 (N_23108,N_21440,N_21744);
nand U23109 (N_23109,N_21585,N_21729);
and U23110 (N_23110,N_21538,N_22143);
or U23111 (N_23111,N_21874,N_22188);
nand U23112 (N_23112,N_22489,N_21776);
xnor U23113 (N_23113,N_21796,N_21493);
and U23114 (N_23114,N_21826,N_21814);
nand U23115 (N_23115,N_22375,N_22178);
xor U23116 (N_23116,N_21272,N_22085);
nor U23117 (N_23117,N_22247,N_21579);
or U23118 (N_23118,N_21266,N_22025);
and U23119 (N_23119,N_22465,N_22203);
or U23120 (N_23120,N_22418,N_22327);
nand U23121 (N_23121,N_21506,N_21717);
and U23122 (N_23122,N_21819,N_21633);
or U23123 (N_23123,N_22183,N_22360);
and U23124 (N_23124,N_21385,N_21713);
xor U23125 (N_23125,N_21538,N_21478);
nor U23126 (N_23126,N_22115,N_21737);
nor U23127 (N_23127,N_21554,N_22263);
nor U23128 (N_23128,N_21763,N_21474);
xor U23129 (N_23129,N_21421,N_21840);
nand U23130 (N_23130,N_22405,N_21277);
or U23131 (N_23131,N_22067,N_21987);
xor U23132 (N_23132,N_22117,N_21868);
or U23133 (N_23133,N_22456,N_22358);
nor U23134 (N_23134,N_21977,N_21783);
and U23135 (N_23135,N_21384,N_22416);
xor U23136 (N_23136,N_21428,N_22236);
or U23137 (N_23137,N_22393,N_21687);
nand U23138 (N_23138,N_21408,N_21741);
nand U23139 (N_23139,N_21356,N_22476);
and U23140 (N_23140,N_22330,N_22383);
and U23141 (N_23141,N_22474,N_21540);
nor U23142 (N_23142,N_22225,N_21432);
or U23143 (N_23143,N_22098,N_22452);
or U23144 (N_23144,N_22344,N_21452);
xor U23145 (N_23145,N_22026,N_22009);
and U23146 (N_23146,N_21944,N_21400);
nor U23147 (N_23147,N_22028,N_21494);
and U23148 (N_23148,N_21680,N_21525);
or U23149 (N_23149,N_22162,N_22145);
nor U23150 (N_23150,N_21878,N_21728);
nand U23151 (N_23151,N_22053,N_22195);
and U23152 (N_23152,N_22256,N_22252);
xor U23153 (N_23153,N_22056,N_22000);
xnor U23154 (N_23154,N_21421,N_22333);
and U23155 (N_23155,N_22457,N_21321);
nand U23156 (N_23156,N_22031,N_21651);
nor U23157 (N_23157,N_22387,N_22144);
or U23158 (N_23158,N_21459,N_21992);
or U23159 (N_23159,N_22445,N_21952);
or U23160 (N_23160,N_22256,N_21434);
nor U23161 (N_23161,N_22119,N_21450);
and U23162 (N_23162,N_22248,N_21891);
nand U23163 (N_23163,N_21779,N_21499);
xor U23164 (N_23164,N_21469,N_21853);
and U23165 (N_23165,N_22051,N_22410);
nor U23166 (N_23166,N_22077,N_21862);
nand U23167 (N_23167,N_21566,N_22085);
nand U23168 (N_23168,N_21899,N_22138);
xnor U23169 (N_23169,N_21491,N_22392);
nand U23170 (N_23170,N_21552,N_21299);
or U23171 (N_23171,N_22422,N_21412);
and U23172 (N_23172,N_21506,N_21781);
and U23173 (N_23173,N_22053,N_21724);
or U23174 (N_23174,N_21405,N_21637);
nand U23175 (N_23175,N_21945,N_21793);
nor U23176 (N_23176,N_22304,N_21809);
and U23177 (N_23177,N_22188,N_22392);
xnor U23178 (N_23178,N_21620,N_22429);
and U23179 (N_23179,N_21886,N_22358);
nor U23180 (N_23180,N_22212,N_21766);
nor U23181 (N_23181,N_22169,N_22442);
and U23182 (N_23182,N_22427,N_22408);
nand U23183 (N_23183,N_21757,N_21440);
nor U23184 (N_23184,N_22300,N_22431);
xor U23185 (N_23185,N_21901,N_21531);
or U23186 (N_23186,N_22292,N_21310);
nand U23187 (N_23187,N_21818,N_21623);
or U23188 (N_23188,N_21396,N_21713);
nor U23189 (N_23189,N_22180,N_21581);
xor U23190 (N_23190,N_21488,N_21361);
nand U23191 (N_23191,N_22074,N_22471);
nor U23192 (N_23192,N_21846,N_22479);
nand U23193 (N_23193,N_21371,N_21657);
xnor U23194 (N_23194,N_22277,N_21964);
nand U23195 (N_23195,N_21355,N_21324);
xnor U23196 (N_23196,N_21898,N_22367);
and U23197 (N_23197,N_21487,N_22061);
or U23198 (N_23198,N_22098,N_22432);
or U23199 (N_23199,N_21510,N_22010);
or U23200 (N_23200,N_21942,N_21570);
nand U23201 (N_23201,N_22398,N_21875);
nand U23202 (N_23202,N_22014,N_21991);
xor U23203 (N_23203,N_21639,N_21602);
and U23204 (N_23204,N_21874,N_22186);
and U23205 (N_23205,N_21908,N_22307);
or U23206 (N_23206,N_22034,N_22334);
xor U23207 (N_23207,N_21456,N_21320);
nand U23208 (N_23208,N_21680,N_21768);
nand U23209 (N_23209,N_21749,N_22098);
nand U23210 (N_23210,N_21519,N_21875);
xnor U23211 (N_23211,N_22327,N_21574);
nor U23212 (N_23212,N_22414,N_22242);
nand U23213 (N_23213,N_21496,N_22410);
and U23214 (N_23214,N_22370,N_22460);
nand U23215 (N_23215,N_22109,N_22396);
nor U23216 (N_23216,N_22407,N_22200);
or U23217 (N_23217,N_21450,N_21590);
and U23218 (N_23218,N_21705,N_21559);
nand U23219 (N_23219,N_22285,N_22349);
nand U23220 (N_23220,N_22099,N_21699);
and U23221 (N_23221,N_22065,N_22294);
nor U23222 (N_23222,N_21964,N_21511);
nor U23223 (N_23223,N_21784,N_22162);
nor U23224 (N_23224,N_21335,N_21844);
nand U23225 (N_23225,N_21671,N_22392);
nor U23226 (N_23226,N_21299,N_21599);
or U23227 (N_23227,N_21997,N_21646);
nor U23228 (N_23228,N_21292,N_22389);
xor U23229 (N_23229,N_22350,N_22146);
xnor U23230 (N_23230,N_21502,N_22431);
and U23231 (N_23231,N_22030,N_22103);
and U23232 (N_23232,N_21673,N_22287);
nor U23233 (N_23233,N_21566,N_21560);
xnor U23234 (N_23234,N_22255,N_21343);
nor U23235 (N_23235,N_21586,N_21727);
and U23236 (N_23236,N_22312,N_21663);
nand U23237 (N_23237,N_22206,N_21344);
nand U23238 (N_23238,N_21761,N_22309);
nor U23239 (N_23239,N_22200,N_21728);
nor U23240 (N_23240,N_21949,N_21917);
nand U23241 (N_23241,N_21280,N_22079);
xnor U23242 (N_23242,N_22268,N_22455);
xor U23243 (N_23243,N_21580,N_22227);
xor U23244 (N_23244,N_21348,N_22395);
or U23245 (N_23245,N_22402,N_22331);
or U23246 (N_23246,N_21444,N_22440);
nor U23247 (N_23247,N_21261,N_21980);
or U23248 (N_23248,N_21905,N_22357);
and U23249 (N_23249,N_22306,N_22098);
and U23250 (N_23250,N_21264,N_22066);
and U23251 (N_23251,N_21463,N_21275);
nor U23252 (N_23252,N_21524,N_21897);
xnor U23253 (N_23253,N_21978,N_21671);
nor U23254 (N_23254,N_21743,N_21495);
nand U23255 (N_23255,N_21946,N_22012);
nor U23256 (N_23256,N_21626,N_22463);
nor U23257 (N_23257,N_21487,N_21683);
and U23258 (N_23258,N_22324,N_22484);
or U23259 (N_23259,N_21371,N_22380);
or U23260 (N_23260,N_21526,N_21774);
nand U23261 (N_23261,N_22204,N_21345);
nand U23262 (N_23262,N_21320,N_22071);
nand U23263 (N_23263,N_21372,N_22296);
nand U23264 (N_23264,N_22062,N_21404);
xor U23265 (N_23265,N_21702,N_21646);
and U23266 (N_23266,N_21463,N_21655);
nor U23267 (N_23267,N_21743,N_21645);
and U23268 (N_23268,N_21257,N_22254);
xor U23269 (N_23269,N_21693,N_21317);
nor U23270 (N_23270,N_21587,N_21473);
nand U23271 (N_23271,N_21742,N_21775);
nand U23272 (N_23272,N_21484,N_22117);
nor U23273 (N_23273,N_21918,N_21262);
nor U23274 (N_23274,N_21573,N_21996);
xnor U23275 (N_23275,N_21416,N_21567);
xor U23276 (N_23276,N_21350,N_21381);
and U23277 (N_23277,N_21922,N_21833);
xor U23278 (N_23278,N_21910,N_22498);
and U23279 (N_23279,N_22013,N_22333);
or U23280 (N_23280,N_21481,N_21708);
nand U23281 (N_23281,N_22101,N_21578);
xnor U23282 (N_23282,N_21993,N_21860);
and U23283 (N_23283,N_21656,N_22402);
and U23284 (N_23284,N_21739,N_21308);
xnor U23285 (N_23285,N_22203,N_22353);
and U23286 (N_23286,N_22013,N_21515);
xor U23287 (N_23287,N_21257,N_21457);
nor U23288 (N_23288,N_22177,N_21647);
and U23289 (N_23289,N_22295,N_21928);
xor U23290 (N_23290,N_21477,N_21389);
nor U23291 (N_23291,N_21722,N_22108);
and U23292 (N_23292,N_22354,N_22486);
and U23293 (N_23293,N_21817,N_22088);
xor U23294 (N_23294,N_22495,N_22061);
nor U23295 (N_23295,N_22222,N_22353);
nand U23296 (N_23296,N_21544,N_22426);
or U23297 (N_23297,N_21796,N_22057);
nor U23298 (N_23298,N_21666,N_22302);
xnor U23299 (N_23299,N_21278,N_22407);
and U23300 (N_23300,N_22182,N_22235);
xor U23301 (N_23301,N_21778,N_21652);
nand U23302 (N_23302,N_22471,N_22164);
nand U23303 (N_23303,N_22398,N_21612);
nor U23304 (N_23304,N_22398,N_21623);
nand U23305 (N_23305,N_21624,N_21901);
or U23306 (N_23306,N_21706,N_22247);
xnor U23307 (N_23307,N_21728,N_21271);
and U23308 (N_23308,N_21439,N_21320);
or U23309 (N_23309,N_22114,N_21954);
or U23310 (N_23310,N_21855,N_21673);
nor U23311 (N_23311,N_22343,N_21527);
nor U23312 (N_23312,N_21799,N_21557);
nand U23313 (N_23313,N_21943,N_21667);
nor U23314 (N_23314,N_21869,N_21672);
and U23315 (N_23315,N_21519,N_22434);
and U23316 (N_23316,N_22374,N_21738);
nand U23317 (N_23317,N_22255,N_21651);
xor U23318 (N_23318,N_21588,N_21999);
xor U23319 (N_23319,N_22311,N_21639);
xnor U23320 (N_23320,N_21783,N_22201);
and U23321 (N_23321,N_21673,N_21987);
and U23322 (N_23322,N_21954,N_21462);
nor U23323 (N_23323,N_21893,N_21381);
or U23324 (N_23324,N_21723,N_21916);
nand U23325 (N_23325,N_21361,N_21255);
or U23326 (N_23326,N_21284,N_21435);
xor U23327 (N_23327,N_21649,N_22107);
and U23328 (N_23328,N_22484,N_22113);
and U23329 (N_23329,N_22422,N_21592);
or U23330 (N_23330,N_21829,N_21406);
and U23331 (N_23331,N_22321,N_21400);
and U23332 (N_23332,N_22227,N_22461);
and U23333 (N_23333,N_21521,N_21251);
nor U23334 (N_23334,N_22180,N_21947);
and U23335 (N_23335,N_22301,N_21933);
or U23336 (N_23336,N_21820,N_22114);
and U23337 (N_23337,N_21365,N_21912);
xnor U23338 (N_23338,N_21684,N_21386);
and U23339 (N_23339,N_22209,N_21868);
or U23340 (N_23340,N_21361,N_21451);
nand U23341 (N_23341,N_21914,N_22204);
nor U23342 (N_23342,N_22474,N_22409);
nor U23343 (N_23343,N_21432,N_22019);
xnor U23344 (N_23344,N_22062,N_22072);
xnor U23345 (N_23345,N_21640,N_22298);
or U23346 (N_23346,N_21831,N_21538);
xnor U23347 (N_23347,N_21694,N_22385);
or U23348 (N_23348,N_21559,N_22482);
and U23349 (N_23349,N_22144,N_21838);
xor U23350 (N_23350,N_22065,N_22159);
nand U23351 (N_23351,N_21588,N_21712);
nor U23352 (N_23352,N_21499,N_21647);
and U23353 (N_23353,N_21999,N_22094);
nand U23354 (N_23354,N_22458,N_22214);
or U23355 (N_23355,N_22428,N_21649);
nor U23356 (N_23356,N_21919,N_22045);
and U23357 (N_23357,N_22110,N_21663);
nand U23358 (N_23358,N_22400,N_22003);
nand U23359 (N_23359,N_22402,N_22398);
xor U23360 (N_23360,N_21690,N_21770);
and U23361 (N_23361,N_22324,N_21918);
and U23362 (N_23362,N_22116,N_22106);
and U23363 (N_23363,N_21810,N_21430);
xor U23364 (N_23364,N_21834,N_21816);
nand U23365 (N_23365,N_21364,N_22281);
and U23366 (N_23366,N_21756,N_21451);
xor U23367 (N_23367,N_21349,N_21782);
nand U23368 (N_23368,N_22028,N_22320);
nor U23369 (N_23369,N_21682,N_21265);
xor U23370 (N_23370,N_21919,N_22374);
and U23371 (N_23371,N_22220,N_22174);
and U23372 (N_23372,N_21955,N_21875);
nand U23373 (N_23373,N_22132,N_21343);
and U23374 (N_23374,N_22496,N_22348);
and U23375 (N_23375,N_21303,N_21267);
and U23376 (N_23376,N_21706,N_21433);
nand U23377 (N_23377,N_21648,N_21998);
nand U23378 (N_23378,N_22032,N_21473);
nand U23379 (N_23379,N_22182,N_22365);
and U23380 (N_23380,N_21961,N_22076);
nand U23381 (N_23381,N_21443,N_21389);
nand U23382 (N_23382,N_21624,N_21641);
xnor U23383 (N_23383,N_21284,N_22359);
xnor U23384 (N_23384,N_21535,N_21481);
xnor U23385 (N_23385,N_22355,N_21545);
xnor U23386 (N_23386,N_21260,N_22302);
nand U23387 (N_23387,N_22282,N_21996);
and U23388 (N_23388,N_22138,N_21735);
and U23389 (N_23389,N_21944,N_22361);
nor U23390 (N_23390,N_21890,N_21268);
nand U23391 (N_23391,N_22287,N_22444);
or U23392 (N_23392,N_22059,N_22413);
or U23393 (N_23393,N_21253,N_21682);
nor U23394 (N_23394,N_21998,N_22231);
nand U23395 (N_23395,N_21270,N_22075);
nor U23396 (N_23396,N_22478,N_21350);
nand U23397 (N_23397,N_21466,N_22023);
nor U23398 (N_23398,N_22240,N_22272);
and U23399 (N_23399,N_21444,N_21270);
nand U23400 (N_23400,N_21989,N_21407);
nor U23401 (N_23401,N_22495,N_21634);
xnor U23402 (N_23402,N_21454,N_21951);
and U23403 (N_23403,N_22020,N_22390);
nand U23404 (N_23404,N_21347,N_21545);
xor U23405 (N_23405,N_21859,N_21932);
nor U23406 (N_23406,N_21514,N_22138);
xor U23407 (N_23407,N_22321,N_22148);
xor U23408 (N_23408,N_22018,N_21612);
xnor U23409 (N_23409,N_21933,N_22209);
nor U23410 (N_23410,N_22018,N_22374);
or U23411 (N_23411,N_21619,N_22024);
xor U23412 (N_23412,N_22223,N_21728);
xor U23413 (N_23413,N_21563,N_21373);
or U23414 (N_23414,N_21970,N_22354);
nor U23415 (N_23415,N_21273,N_22457);
nor U23416 (N_23416,N_22269,N_21530);
and U23417 (N_23417,N_22376,N_21629);
nand U23418 (N_23418,N_21656,N_21666);
nand U23419 (N_23419,N_22241,N_21621);
xor U23420 (N_23420,N_21487,N_21578);
nor U23421 (N_23421,N_21527,N_21656);
xnor U23422 (N_23422,N_21548,N_21971);
or U23423 (N_23423,N_21286,N_21588);
and U23424 (N_23424,N_21825,N_21523);
nor U23425 (N_23425,N_22158,N_22363);
nand U23426 (N_23426,N_21699,N_21335);
nor U23427 (N_23427,N_21306,N_22314);
or U23428 (N_23428,N_21589,N_22239);
nor U23429 (N_23429,N_21430,N_21279);
nand U23430 (N_23430,N_21540,N_22280);
xnor U23431 (N_23431,N_21815,N_22210);
and U23432 (N_23432,N_21317,N_21311);
nand U23433 (N_23433,N_22307,N_22368);
xnor U23434 (N_23434,N_22040,N_21500);
and U23435 (N_23435,N_22160,N_22368);
nand U23436 (N_23436,N_22440,N_21473);
nor U23437 (N_23437,N_21910,N_21839);
nand U23438 (N_23438,N_21997,N_22183);
nor U23439 (N_23439,N_21861,N_21709);
nand U23440 (N_23440,N_22381,N_22132);
or U23441 (N_23441,N_21477,N_21525);
or U23442 (N_23442,N_21950,N_22195);
or U23443 (N_23443,N_21291,N_21691);
nor U23444 (N_23444,N_21334,N_21327);
and U23445 (N_23445,N_21832,N_21640);
xor U23446 (N_23446,N_21540,N_22449);
nor U23447 (N_23447,N_22254,N_21885);
nor U23448 (N_23448,N_21559,N_22113);
nand U23449 (N_23449,N_21679,N_21346);
nor U23450 (N_23450,N_21299,N_22112);
xor U23451 (N_23451,N_22017,N_21977);
xnor U23452 (N_23452,N_22206,N_21399);
xnor U23453 (N_23453,N_22495,N_22016);
nor U23454 (N_23454,N_21516,N_21377);
nor U23455 (N_23455,N_22162,N_22043);
or U23456 (N_23456,N_21696,N_22378);
nand U23457 (N_23457,N_22418,N_21859);
and U23458 (N_23458,N_22034,N_22173);
or U23459 (N_23459,N_22111,N_21864);
nand U23460 (N_23460,N_21795,N_21976);
or U23461 (N_23461,N_22376,N_22164);
or U23462 (N_23462,N_21270,N_22162);
or U23463 (N_23463,N_21923,N_21388);
or U23464 (N_23464,N_21706,N_22029);
and U23465 (N_23465,N_21816,N_21773);
and U23466 (N_23466,N_21654,N_22288);
and U23467 (N_23467,N_22117,N_22010);
or U23468 (N_23468,N_21360,N_21579);
xnor U23469 (N_23469,N_21463,N_22310);
or U23470 (N_23470,N_21775,N_21698);
xnor U23471 (N_23471,N_22056,N_21298);
nand U23472 (N_23472,N_22142,N_21816);
and U23473 (N_23473,N_21637,N_21603);
or U23474 (N_23474,N_21502,N_21377);
and U23475 (N_23475,N_21848,N_21332);
nand U23476 (N_23476,N_22193,N_22231);
or U23477 (N_23477,N_21741,N_22325);
nand U23478 (N_23478,N_21357,N_21767);
and U23479 (N_23479,N_22119,N_22452);
or U23480 (N_23480,N_22092,N_21255);
and U23481 (N_23481,N_22390,N_22458);
nor U23482 (N_23482,N_21567,N_21423);
nor U23483 (N_23483,N_21450,N_21596);
nor U23484 (N_23484,N_21632,N_22033);
nor U23485 (N_23485,N_21517,N_22367);
and U23486 (N_23486,N_21822,N_21282);
and U23487 (N_23487,N_21711,N_21755);
nand U23488 (N_23488,N_22312,N_22499);
and U23489 (N_23489,N_21363,N_21267);
or U23490 (N_23490,N_22497,N_22046);
or U23491 (N_23491,N_22082,N_22337);
and U23492 (N_23492,N_21689,N_22095);
and U23493 (N_23493,N_21912,N_21858);
xnor U23494 (N_23494,N_21800,N_21680);
nand U23495 (N_23495,N_21826,N_22161);
and U23496 (N_23496,N_21774,N_22431);
nor U23497 (N_23497,N_21929,N_22379);
or U23498 (N_23498,N_21631,N_21713);
or U23499 (N_23499,N_22346,N_21811);
or U23500 (N_23500,N_21690,N_22089);
nor U23501 (N_23501,N_22277,N_21457);
xor U23502 (N_23502,N_22063,N_21612);
nor U23503 (N_23503,N_21919,N_21525);
xnor U23504 (N_23504,N_21547,N_21553);
and U23505 (N_23505,N_21469,N_22440);
and U23506 (N_23506,N_22281,N_21583);
and U23507 (N_23507,N_21866,N_22396);
nand U23508 (N_23508,N_22428,N_22261);
nand U23509 (N_23509,N_22293,N_22439);
nor U23510 (N_23510,N_22097,N_22117);
or U23511 (N_23511,N_21981,N_22423);
or U23512 (N_23512,N_22120,N_21367);
xor U23513 (N_23513,N_22293,N_22305);
or U23514 (N_23514,N_21648,N_22216);
or U23515 (N_23515,N_22188,N_21354);
xnor U23516 (N_23516,N_22210,N_21595);
and U23517 (N_23517,N_21610,N_21661);
and U23518 (N_23518,N_21656,N_21967);
xnor U23519 (N_23519,N_22450,N_22157);
or U23520 (N_23520,N_22439,N_21959);
nor U23521 (N_23521,N_21280,N_22404);
and U23522 (N_23522,N_21776,N_22289);
nor U23523 (N_23523,N_21312,N_22186);
xnor U23524 (N_23524,N_21945,N_21641);
nor U23525 (N_23525,N_22477,N_22003);
and U23526 (N_23526,N_22324,N_21501);
or U23527 (N_23527,N_22052,N_21659);
or U23528 (N_23528,N_21271,N_22450);
and U23529 (N_23529,N_21271,N_21570);
or U23530 (N_23530,N_21711,N_22418);
xnor U23531 (N_23531,N_22220,N_22469);
nand U23532 (N_23532,N_22156,N_22259);
nand U23533 (N_23533,N_21497,N_22304);
nor U23534 (N_23534,N_21532,N_22368);
xor U23535 (N_23535,N_22410,N_21782);
or U23536 (N_23536,N_22104,N_21615);
nand U23537 (N_23537,N_21941,N_21536);
nand U23538 (N_23538,N_21443,N_22051);
xnor U23539 (N_23539,N_21488,N_21820);
nand U23540 (N_23540,N_22402,N_21524);
nor U23541 (N_23541,N_22243,N_22199);
xnor U23542 (N_23542,N_21682,N_21495);
nor U23543 (N_23543,N_22460,N_21679);
or U23544 (N_23544,N_22134,N_22473);
nor U23545 (N_23545,N_22275,N_21935);
nor U23546 (N_23546,N_22066,N_21810);
nor U23547 (N_23547,N_21784,N_22253);
and U23548 (N_23548,N_21727,N_21370);
nand U23549 (N_23549,N_22419,N_22470);
or U23550 (N_23550,N_21515,N_22030);
xor U23551 (N_23551,N_21270,N_21581);
nor U23552 (N_23552,N_21669,N_22011);
and U23553 (N_23553,N_21730,N_21304);
or U23554 (N_23554,N_21410,N_21290);
xnor U23555 (N_23555,N_21406,N_21392);
nand U23556 (N_23556,N_22415,N_21483);
or U23557 (N_23557,N_22185,N_22206);
nand U23558 (N_23558,N_21861,N_21789);
xor U23559 (N_23559,N_21907,N_21815);
xor U23560 (N_23560,N_21803,N_22117);
xor U23561 (N_23561,N_21447,N_21502);
and U23562 (N_23562,N_22161,N_21637);
or U23563 (N_23563,N_21779,N_21503);
or U23564 (N_23564,N_22225,N_22453);
nor U23565 (N_23565,N_21656,N_21842);
nand U23566 (N_23566,N_22227,N_21843);
nor U23567 (N_23567,N_21758,N_22470);
nand U23568 (N_23568,N_21538,N_22335);
nand U23569 (N_23569,N_21284,N_21680);
nand U23570 (N_23570,N_22388,N_22331);
and U23571 (N_23571,N_21915,N_22406);
xor U23572 (N_23572,N_21875,N_22203);
nand U23573 (N_23573,N_22112,N_21900);
and U23574 (N_23574,N_22327,N_21276);
xnor U23575 (N_23575,N_21407,N_21552);
xnor U23576 (N_23576,N_21275,N_21336);
nand U23577 (N_23577,N_21854,N_21721);
xor U23578 (N_23578,N_21582,N_22371);
or U23579 (N_23579,N_21864,N_21407);
nand U23580 (N_23580,N_22000,N_22404);
or U23581 (N_23581,N_21322,N_21654);
or U23582 (N_23582,N_21257,N_21853);
or U23583 (N_23583,N_21976,N_21353);
and U23584 (N_23584,N_22286,N_22499);
nand U23585 (N_23585,N_21450,N_21544);
and U23586 (N_23586,N_21962,N_22130);
or U23587 (N_23587,N_21586,N_21744);
and U23588 (N_23588,N_21521,N_21735);
or U23589 (N_23589,N_21439,N_22006);
or U23590 (N_23590,N_22312,N_22373);
xor U23591 (N_23591,N_21270,N_22030);
or U23592 (N_23592,N_21921,N_22161);
nand U23593 (N_23593,N_22236,N_22476);
and U23594 (N_23594,N_22035,N_22478);
or U23595 (N_23595,N_22097,N_21559);
and U23596 (N_23596,N_22192,N_22210);
or U23597 (N_23597,N_21828,N_22083);
nand U23598 (N_23598,N_21960,N_21934);
xnor U23599 (N_23599,N_21897,N_22190);
nand U23600 (N_23600,N_21636,N_21866);
xnor U23601 (N_23601,N_22339,N_22335);
nor U23602 (N_23602,N_21675,N_21731);
nand U23603 (N_23603,N_21833,N_21454);
nand U23604 (N_23604,N_21311,N_21686);
and U23605 (N_23605,N_21986,N_22326);
xnor U23606 (N_23606,N_22106,N_22034);
or U23607 (N_23607,N_22455,N_22153);
or U23608 (N_23608,N_22283,N_21879);
nand U23609 (N_23609,N_22171,N_22029);
or U23610 (N_23610,N_21281,N_21853);
nand U23611 (N_23611,N_22112,N_21971);
or U23612 (N_23612,N_21753,N_21664);
or U23613 (N_23613,N_22159,N_22022);
and U23614 (N_23614,N_21396,N_21852);
xor U23615 (N_23615,N_21744,N_21329);
nor U23616 (N_23616,N_21785,N_21720);
and U23617 (N_23617,N_21719,N_22127);
or U23618 (N_23618,N_21808,N_22145);
nand U23619 (N_23619,N_22465,N_22491);
or U23620 (N_23620,N_21820,N_21822);
xor U23621 (N_23621,N_22241,N_21600);
nor U23622 (N_23622,N_21627,N_21599);
nor U23623 (N_23623,N_21688,N_21405);
nand U23624 (N_23624,N_22056,N_21710);
and U23625 (N_23625,N_21830,N_21758);
nor U23626 (N_23626,N_21931,N_22028);
and U23627 (N_23627,N_22350,N_21570);
or U23628 (N_23628,N_21694,N_21834);
xnor U23629 (N_23629,N_21372,N_21899);
or U23630 (N_23630,N_22033,N_22243);
nor U23631 (N_23631,N_21843,N_22298);
nand U23632 (N_23632,N_21636,N_21587);
xor U23633 (N_23633,N_21724,N_22468);
nor U23634 (N_23634,N_21793,N_21580);
nor U23635 (N_23635,N_22401,N_21551);
nor U23636 (N_23636,N_21500,N_22039);
or U23637 (N_23637,N_21383,N_21934);
and U23638 (N_23638,N_21890,N_21593);
xnor U23639 (N_23639,N_21539,N_21262);
nor U23640 (N_23640,N_22269,N_22325);
or U23641 (N_23641,N_22359,N_22307);
xnor U23642 (N_23642,N_21884,N_22407);
nor U23643 (N_23643,N_21461,N_21369);
xnor U23644 (N_23644,N_21300,N_21713);
nand U23645 (N_23645,N_21393,N_22377);
nor U23646 (N_23646,N_21745,N_21406);
nor U23647 (N_23647,N_21678,N_21845);
and U23648 (N_23648,N_21593,N_21278);
xor U23649 (N_23649,N_21549,N_22460);
xnor U23650 (N_23650,N_21444,N_21859);
and U23651 (N_23651,N_21393,N_21887);
nor U23652 (N_23652,N_21284,N_21758);
xnor U23653 (N_23653,N_21299,N_22200);
and U23654 (N_23654,N_22236,N_21258);
or U23655 (N_23655,N_21954,N_21359);
nor U23656 (N_23656,N_21725,N_21996);
or U23657 (N_23657,N_21586,N_21614);
nor U23658 (N_23658,N_21794,N_21474);
xor U23659 (N_23659,N_21833,N_22188);
nand U23660 (N_23660,N_22042,N_21472);
or U23661 (N_23661,N_21314,N_21368);
and U23662 (N_23662,N_21641,N_21767);
nand U23663 (N_23663,N_21932,N_22211);
nand U23664 (N_23664,N_22010,N_21759);
nor U23665 (N_23665,N_22079,N_21380);
or U23666 (N_23666,N_21306,N_22332);
xor U23667 (N_23667,N_21861,N_21731);
and U23668 (N_23668,N_22303,N_21623);
xor U23669 (N_23669,N_22473,N_22267);
or U23670 (N_23670,N_22494,N_21435);
or U23671 (N_23671,N_21502,N_21627);
or U23672 (N_23672,N_22444,N_21961);
and U23673 (N_23673,N_21522,N_22071);
and U23674 (N_23674,N_21422,N_22011);
and U23675 (N_23675,N_22482,N_21528);
or U23676 (N_23676,N_21862,N_21490);
xnor U23677 (N_23677,N_22182,N_21505);
nand U23678 (N_23678,N_21895,N_22214);
nand U23679 (N_23679,N_22224,N_22491);
nor U23680 (N_23680,N_21636,N_21811);
xor U23681 (N_23681,N_21748,N_22176);
or U23682 (N_23682,N_21955,N_22369);
xnor U23683 (N_23683,N_22240,N_21414);
or U23684 (N_23684,N_21331,N_21734);
nor U23685 (N_23685,N_21378,N_21597);
xnor U23686 (N_23686,N_21583,N_22101);
xor U23687 (N_23687,N_21509,N_21584);
xor U23688 (N_23688,N_22372,N_21359);
or U23689 (N_23689,N_22481,N_22344);
or U23690 (N_23690,N_21736,N_22354);
and U23691 (N_23691,N_21647,N_22277);
xnor U23692 (N_23692,N_22280,N_21436);
or U23693 (N_23693,N_21527,N_21476);
and U23694 (N_23694,N_22139,N_21528);
nand U23695 (N_23695,N_22216,N_22333);
nor U23696 (N_23696,N_21967,N_22282);
nor U23697 (N_23697,N_21654,N_22460);
nor U23698 (N_23698,N_22254,N_22402);
xnor U23699 (N_23699,N_21894,N_21765);
and U23700 (N_23700,N_22360,N_21358);
nand U23701 (N_23701,N_22421,N_21699);
and U23702 (N_23702,N_22217,N_21279);
xor U23703 (N_23703,N_21722,N_21662);
nor U23704 (N_23704,N_22311,N_22252);
and U23705 (N_23705,N_22259,N_21563);
xor U23706 (N_23706,N_21584,N_21778);
and U23707 (N_23707,N_22067,N_22286);
nand U23708 (N_23708,N_21763,N_21485);
nor U23709 (N_23709,N_21657,N_21499);
nand U23710 (N_23710,N_21611,N_21772);
xnor U23711 (N_23711,N_22115,N_22489);
xnor U23712 (N_23712,N_22240,N_22464);
nor U23713 (N_23713,N_21889,N_22086);
xor U23714 (N_23714,N_21751,N_21555);
and U23715 (N_23715,N_21884,N_21453);
nor U23716 (N_23716,N_22210,N_22081);
xor U23717 (N_23717,N_21283,N_22421);
xor U23718 (N_23718,N_21297,N_22358);
or U23719 (N_23719,N_22387,N_21371);
xnor U23720 (N_23720,N_21611,N_22339);
and U23721 (N_23721,N_22062,N_22411);
and U23722 (N_23722,N_21356,N_22053);
and U23723 (N_23723,N_22483,N_21366);
xor U23724 (N_23724,N_22034,N_21942);
xnor U23725 (N_23725,N_21544,N_21346);
xor U23726 (N_23726,N_22372,N_22069);
nand U23727 (N_23727,N_22434,N_21783);
xnor U23728 (N_23728,N_22236,N_21254);
xor U23729 (N_23729,N_22332,N_22294);
and U23730 (N_23730,N_21394,N_21905);
or U23731 (N_23731,N_21578,N_21307);
xnor U23732 (N_23732,N_21463,N_21653);
or U23733 (N_23733,N_21925,N_21756);
xor U23734 (N_23734,N_21963,N_21255);
nand U23735 (N_23735,N_21748,N_21887);
nor U23736 (N_23736,N_22085,N_21488);
or U23737 (N_23737,N_22161,N_22088);
xnor U23738 (N_23738,N_22258,N_22418);
nor U23739 (N_23739,N_21794,N_21623);
and U23740 (N_23740,N_21673,N_21907);
xnor U23741 (N_23741,N_21603,N_22222);
or U23742 (N_23742,N_21255,N_21900);
nand U23743 (N_23743,N_22471,N_21490);
nor U23744 (N_23744,N_21894,N_22435);
nor U23745 (N_23745,N_21978,N_22148);
xnor U23746 (N_23746,N_22252,N_21826);
nor U23747 (N_23747,N_22476,N_22304);
and U23748 (N_23748,N_21250,N_21620);
nand U23749 (N_23749,N_21557,N_21838);
xor U23750 (N_23750,N_22513,N_23426);
nand U23751 (N_23751,N_22507,N_23141);
xnor U23752 (N_23752,N_22964,N_23335);
or U23753 (N_23753,N_23558,N_23056);
nor U23754 (N_23754,N_23130,N_23533);
and U23755 (N_23755,N_22841,N_23009);
xor U23756 (N_23756,N_22697,N_22858);
and U23757 (N_23757,N_22685,N_22860);
and U23758 (N_23758,N_22832,N_23715);
nor U23759 (N_23759,N_23718,N_23495);
nand U23760 (N_23760,N_22517,N_22777);
nand U23761 (N_23761,N_23396,N_22966);
and U23762 (N_23762,N_22885,N_23494);
nand U23763 (N_23763,N_22505,N_23236);
or U23764 (N_23764,N_22625,N_23380);
and U23765 (N_23765,N_23344,N_23617);
nand U23766 (N_23766,N_22552,N_22710);
and U23767 (N_23767,N_23207,N_23687);
nand U23768 (N_23768,N_22615,N_22642);
nor U23769 (N_23769,N_23389,N_22742);
or U23770 (N_23770,N_23322,N_23387);
and U23771 (N_23771,N_22597,N_23278);
xor U23772 (N_23772,N_22867,N_23382);
or U23773 (N_23773,N_22870,N_23279);
xnor U23774 (N_23774,N_22871,N_22994);
xnor U23775 (N_23775,N_23457,N_23662);
xnor U23776 (N_23776,N_23571,N_23485);
nand U23777 (N_23777,N_23593,N_22959);
or U23778 (N_23778,N_22820,N_22603);
xnor U23779 (N_23779,N_23291,N_23492);
or U23780 (N_23780,N_23104,N_23047);
or U23781 (N_23781,N_23476,N_22881);
or U23782 (N_23782,N_22690,N_22947);
nand U23783 (N_23783,N_23181,N_23117);
and U23784 (N_23784,N_22772,N_22812);
nand U23785 (N_23785,N_22981,N_23039);
nor U23786 (N_23786,N_23602,N_22923);
xor U23787 (N_23787,N_22712,N_23468);
nand U23788 (N_23788,N_22795,N_23345);
nand U23789 (N_23789,N_22617,N_22894);
and U23790 (N_23790,N_22606,N_22982);
nand U23791 (N_23791,N_22588,N_23459);
nor U23792 (N_23792,N_22636,N_23452);
xnor U23793 (N_23793,N_23626,N_22883);
or U23794 (N_23794,N_23230,N_22511);
or U23795 (N_23795,N_22839,N_22586);
nor U23796 (N_23796,N_23266,N_23700);
and U23797 (N_23797,N_23247,N_23337);
and U23798 (N_23798,N_22691,N_22957);
or U23799 (N_23799,N_23615,N_22596);
nand U23800 (N_23800,N_22949,N_23084);
nor U23801 (N_23801,N_22549,N_23397);
xnor U23802 (N_23802,N_23562,N_22918);
nor U23803 (N_23803,N_22991,N_22605);
nor U23804 (N_23804,N_23362,N_23560);
or U23805 (N_23805,N_23164,N_22925);
xor U23806 (N_23806,N_23467,N_23106);
nor U23807 (N_23807,N_23512,N_22921);
nand U23808 (N_23808,N_23025,N_22791);
nand U23809 (N_23809,N_22533,N_23388);
and U23810 (N_23810,N_23111,N_23381);
nor U23811 (N_23811,N_23371,N_22581);
and U23812 (N_23812,N_22590,N_23689);
nand U23813 (N_23813,N_23237,N_22518);
and U23814 (N_23814,N_23270,N_23641);
and U23815 (N_23815,N_23638,N_23108);
nor U23816 (N_23816,N_23282,N_23366);
xnor U23817 (N_23817,N_22847,N_23475);
xnor U23818 (N_23818,N_22848,N_23050);
and U23819 (N_23819,N_22919,N_23660);
nand U23820 (N_23820,N_22593,N_23343);
nand U23821 (N_23821,N_23434,N_22626);
and U23822 (N_23822,N_22656,N_23409);
nand U23823 (N_23823,N_22506,N_22988);
xor U23824 (N_23824,N_22724,N_23550);
nand U23825 (N_23825,N_23098,N_22530);
nor U23826 (N_23826,N_23131,N_23392);
or U23827 (N_23827,N_22736,N_23599);
nand U23828 (N_23828,N_23256,N_22749);
nor U23829 (N_23829,N_23515,N_22818);
and U23830 (N_23830,N_23324,N_23124);
nand U23831 (N_23831,N_23724,N_23151);
nand U23832 (N_23832,N_22531,N_22732);
nand U23833 (N_23833,N_22864,N_22936);
nand U23834 (N_23834,N_22700,N_23316);
xor U23835 (N_23835,N_23243,N_22560);
nand U23836 (N_23836,N_23506,N_23307);
nand U23837 (N_23837,N_23020,N_23676);
xor U23838 (N_23838,N_22608,N_22575);
nor U23839 (N_23839,N_23450,N_22905);
or U23840 (N_23840,N_22973,N_23711);
or U23841 (N_23841,N_23206,N_23358);
xor U23842 (N_23842,N_22933,N_23139);
and U23843 (N_23843,N_23632,N_22859);
and U23844 (N_23844,N_22904,N_23294);
nor U23845 (N_23845,N_22790,N_22670);
or U23846 (N_23846,N_23422,N_22601);
xnor U23847 (N_23847,N_23437,N_23037);
nor U23848 (N_23848,N_23348,N_22713);
or U23849 (N_23849,N_23157,N_23746);
or U23850 (N_23850,N_23581,N_22579);
xnor U23851 (N_23851,N_22971,N_23144);
xnor U23852 (N_23852,N_22932,N_22683);
nand U23853 (N_23853,N_22693,N_23691);
and U23854 (N_23854,N_23138,N_23481);
and U23855 (N_23855,N_23351,N_23150);
and U23856 (N_23856,N_23140,N_22726);
xor U23857 (N_23857,N_23717,N_23738);
xnor U23858 (N_23858,N_23684,N_22613);
and U23859 (N_23859,N_23579,N_22715);
or U23860 (N_23860,N_23167,N_23233);
nand U23861 (N_23861,N_22663,N_23285);
nor U23862 (N_23862,N_22644,N_23624);
and U23863 (N_23863,N_22938,N_22676);
nor U23864 (N_23864,N_23707,N_23603);
xor U23865 (N_23865,N_23162,N_23209);
nand U23866 (N_23866,N_23100,N_22872);
and U23867 (N_23867,N_23716,N_23538);
and U23868 (N_23868,N_23545,N_23591);
and U23869 (N_23869,N_22532,N_23143);
nor U23870 (N_23870,N_22708,N_22861);
xor U23871 (N_23871,N_23188,N_23187);
xor U23872 (N_23872,N_23401,N_23504);
or U23873 (N_23873,N_23186,N_23745);
and U23874 (N_23874,N_23260,N_23673);
and U23875 (N_23875,N_23491,N_23511);
nor U23876 (N_23876,N_22942,N_23318);
and U23877 (N_23877,N_22559,N_23336);
nand U23878 (N_23878,N_22621,N_23465);
and U23879 (N_23879,N_23722,N_23415);
nor U23880 (N_23880,N_23184,N_23532);
xor U23881 (N_23881,N_23274,N_23079);
and U23882 (N_23882,N_22900,N_23120);
nand U23883 (N_23883,N_22696,N_23369);
nor U23884 (N_23884,N_23419,N_23589);
nor U23885 (N_23885,N_23478,N_23175);
nand U23886 (N_23886,N_23298,N_22884);
or U23887 (N_23887,N_23379,N_22849);
or U23888 (N_23888,N_22875,N_22598);
xnor U23889 (N_23889,N_23542,N_22521);
xnor U23890 (N_23890,N_23099,N_23672);
xnor U23891 (N_23891,N_22512,N_23611);
nand U23892 (N_23892,N_23577,N_22672);
and U23893 (N_23893,N_22874,N_23502);
nor U23894 (N_23894,N_22682,N_22716);
xor U23895 (N_23895,N_22928,N_23172);
nor U23896 (N_23896,N_23251,N_22567);
xnor U23897 (N_23897,N_23086,N_23010);
nand U23898 (N_23898,N_22709,N_22563);
nand U23899 (N_23899,N_22535,N_22536);
and U23900 (N_23900,N_22844,N_23384);
and U23901 (N_23901,N_23173,N_23059);
xnor U23902 (N_23902,N_23651,N_23212);
or U23903 (N_23903,N_22523,N_22969);
or U23904 (N_23904,N_23202,N_22831);
xor U23905 (N_23905,N_22999,N_23352);
nand U23906 (N_23906,N_23564,N_23101);
xor U23907 (N_23907,N_23516,N_23650);
nor U23908 (N_23908,N_23364,N_23326);
and U23909 (N_23909,N_22826,N_23161);
nand U23910 (N_23910,N_23623,N_23547);
and U23911 (N_23911,N_23613,N_22734);
xor U23912 (N_23912,N_23122,N_23634);
xor U23913 (N_23913,N_23429,N_23176);
nand U23914 (N_23914,N_23040,N_23472);
nor U23915 (N_23915,N_22631,N_22610);
or U23916 (N_23916,N_22781,N_22722);
or U23917 (N_23917,N_23166,N_23540);
xnor U23918 (N_23918,N_22935,N_22771);
xor U23919 (N_23919,N_22720,N_23372);
nand U23920 (N_23920,N_23749,N_23303);
and U23921 (N_23921,N_23527,N_22876);
nand U23922 (N_23922,N_22972,N_23290);
nor U23923 (N_23923,N_23304,N_23147);
nand U23924 (N_23924,N_23563,N_23462);
nand U23925 (N_23925,N_22748,N_23425);
nor U23926 (N_23926,N_22646,N_23310);
nor U23927 (N_23927,N_23735,N_22851);
nor U23928 (N_23928,N_23311,N_22721);
and U23929 (N_23929,N_22930,N_22660);
xor U23930 (N_23930,N_22502,N_22850);
and U23931 (N_23931,N_23529,N_23199);
or U23932 (N_23932,N_23618,N_23639);
nor U23933 (N_23933,N_23067,N_22886);
xor U23934 (N_23934,N_22892,N_23596);
nor U23935 (N_23935,N_23661,N_23035);
xor U23936 (N_23936,N_23435,N_22604);
xor U23937 (N_23937,N_22951,N_23081);
and U23938 (N_23938,N_22703,N_23391);
nand U23939 (N_23939,N_23240,N_23667);
xor U23940 (N_23940,N_23097,N_23178);
xnor U23941 (N_23941,N_23567,N_22714);
nand U23942 (N_23942,N_23442,N_23604);
or U23943 (N_23943,N_22809,N_22554);
nor U23944 (N_23944,N_23216,N_23286);
or U23945 (N_23945,N_23353,N_23407);
and U23946 (N_23946,N_22687,N_22706);
nor U23947 (N_23947,N_23329,N_23284);
nor U23948 (N_23948,N_22882,N_23701);
xor U23949 (N_23949,N_23091,N_23729);
nand U23950 (N_23950,N_22728,N_22576);
and U23951 (N_23951,N_22992,N_22985);
nor U23952 (N_23952,N_23622,N_23685);
nor U23953 (N_23953,N_22577,N_22757);
xor U23954 (N_23954,N_22829,N_22842);
or U23955 (N_23955,N_23696,N_22784);
nor U23956 (N_23956,N_23671,N_23552);
nand U23957 (N_23957,N_23438,N_23049);
nand U23958 (N_23958,N_23554,N_22569);
nor U23959 (N_23959,N_23447,N_23509);
xnor U23960 (N_23960,N_22673,N_23683);
nand U23961 (N_23961,N_23261,N_23417);
or U23962 (N_23962,N_22624,N_23073);
or U23963 (N_23963,N_23300,N_23289);
nand U23964 (N_23964,N_23231,N_22853);
and U23965 (N_23965,N_23356,N_23228);
xor U23966 (N_23966,N_23249,N_22797);
nor U23967 (N_23967,N_22580,N_23340);
nand U23968 (N_23968,N_22671,N_23680);
nand U23969 (N_23969,N_23454,N_23395);
and U23970 (N_23970,N_23017,N_23062);
and U23971 (N_23971,N_23486,N_23620);
or U23972 (N_23972,N_22802,N_22774);
and U23973 (N_23973,N_23193,N_22856);
nand U23974 (N_23974,N_22783,N_23332);
or U23975 (N_23975,N_22561,N_23133);
or U23976 (N_23976,N_23460,N_23730);
xnor U23977 (N_23977,N_23649,N_23349);
and U23978 (N_23978,N_22640,N_23728);
and U23979 (N_23979,N_23219,N_23619);
or U23980 (N_23980,N_23721,N_23016);
and U23981 (N_23981,N_23499,N_22753);
xnor U23982 (N_23982,N_22557,N_23148);
nand U23983 (N_23983,N_23125,N_22595);
nand U23984 (N_23984,N_23276,N_23713);
nor U23985 (N_23985,N_23555,N_22801);
or U23986 (N_23986,N_23664,N_23484);
xnor U23987 (N_23987,N_22768,N_22987);
or U23988 (N_23988,N_22934,N_23399);
xor U23989 (N_23989,N_23094,N_22838);
xor U23990 (N_23990,N_23076,N_22759);
nor U23991 (N_23991,N_22611,N_23706);
and U23992 (N_23992,N_23678,N_23112);
or U23993 (N_23993,N_23085,N_22995);
nor U23994 (N_23994,N_22955,N_23192);
nand U23995 (N_23995,N_22914,N_22537);
nand U23996 (N_23996,N_23648,N_22741);
nor U23997 (N_23997,N_23627,N_22819);
xor U23998 (N_23998,N_23183,N_23292);
nor U23999 (N_23999,N_22633,N_23393);
nor U24000 (N_24000,N_22718,N_23584);
or U24001 (N_24001,N_22863,N_23220);
and U24002 (N_24002,N_23065,N_23269);
and U24003 (N_24003,N_23005,N_23046);
and U24004 (N_24004,N_23403,N_23235);
xnor U24005 (N_24005,N_22527,N_23258);
nand U24006 (N_24006,N_23018,N_22571);
nor U24007 (N_24007,N_23090,N_23553);
xnor U24008 (N_24008,N_23296,N_22762);
and U24009 (N_24009,N_23674,N_23208);
xor U24010 (N_24010,N_23297,N_23275);
or U24011 (N_24011,N_23314,N_23606);
or U24012 (N_24012,N_23496,N_23742);
nand U24013 (N_24013,N_22983,N_23410);
or U24014 (N_24014,N_23609,N_22931);
nand U24015 (N_24015,N_22740,N_23497);
or U24016 (N_24016,N_23692,N_23185);
xnor U24017 (N_24017,N_23347,N_23110);
xor U24018 (N_24018,N_22952,N_22570);
xnor U24019 (N_24019,N_23182,N_22692);
nand U24020 (N_24020,N_23211,N_23030);
and U24021 (N_24021,N_23402,N_22619);
nand U24022 (N_24022,N_22767,N_23573);
and U24023 (N_24023,N_23083,N_23338);
xor U24024 (N_24024,N_22998,N_23656);
xor U24025 (N_24025,N_22578,N_23537);
xnor U24026 (N_24026,N_22778,N_23000);
or U24027 (N_24027,N_23312,N_22846);
nor U24028 (N_24028,N_23154,N_23413);
nand U24029 (N_24029,N_22655,N_22543);
nor U24030 (N_24030,N_22622,N_23521);
or U24031 (N_24031,N_23528,N_23375);
nand U24032 (N_24032,N_23668,N_23077);
xor U24033 (N_24033,N_23234,N_23224);
xor U24034 (N_24034,N_23473,N_22540);
nor U24035 (N_24035,N_23149,N_23498);
nand U24036 (N_24036,N_22912,N_23666);
xor U24037 (N_24037,N_23013,N_23203);
xnor U24038 (N_24038,N_22669,N_23041);
nor U24039 (N_24039,N_23232,N_23739);
or U24040 (N_24040,N_23424,N_22776);
nor U24041 (N_24041,N_23360,N_22747);
nand U24042 (N_24042,N_22953,N_23002);
or U24043 (N_24043,N_22893,N_23214);
nand U24044 (N_24044,N_23445,N_23483);
nand U24045 (N_24045,N_23440,N_23163);
or U24046 (N_24046,N_22843,N_22654);
xnor U24047 (N_24047,N_22970,N_22589);
or U24048 (N_24048,N_22524,N_23608);
nor U24049 (N_24049,N_23339,N_22873);
nand U24050 (N_24050,N_23204,N_23663);
xnor U24051 (N_24051,N_23588,N_23404);
nor U24052 (N_24052,N_22616,N_23658);
or U24053 (N_24053,N_22810,N_23451);
and U24054 (N_24054,N_23293,N_23510);
or U24055 (N_24055,N_23694,N_22701);
nand U24056 (N_24056,N_23458,N_23734);
and U24057 (N_24057,N_23569,N_22585);
or U24058 (N_24058,N_23268,N_22739);
nand U24059 (N_24059,N_23042,N_23536);
nor U24060 (N_24060,N_23686,N_22545);
or U24061 (N_24061,N_23054,N_23518);
nand U24062 (N_24062,N_22827,N_22804);
and U24063 (N_24063,N_23582,N_22792);
nand U24064 (N_24064,N_23408,N_23262);
and U24065 (N_24065,N_22584,N_23514);
nand U24066 (N_24066,N_22763,N_23309);
nor U24067 (N_24067,N_22564,N_22594);
or U24068 (N_24068,N_22745,N_23023);
xnor U24069 (N_24069,N_22565,N_23610);
nor U24070 (N_24070,N_22824,N_23334);
and U24071 (N_24071,N_23190,N_22727);
xor U24072 (N_24072,N_22775,N_23743);
and U24073 (N_24073,N_23531,N_23586);
nand U24074 (N_24074,N_23263,N_23313);
nand U24075 (N_24075,N_23549,N_22600);
or U24076 (N_24076,N_23652,N_23535);
and U24077 (N_24077,N_22854,N_22539);
xnor U24078 (N_24078,N_22694,N_23646);
nand U24079 (N_24079,N_22704,N_22520);
or U24080 (N_24080,N_22558,N_23180);
xor U24081 (N_24081,N_22946,N_23045);
or U24082 (N_24082,N_23027,N_22572);
or U24083 (N_24083,N_22711,N_22816);
or U24084 (N_24084,N_23200,N_23082);
and U24085 (N_24085,N_22773,N_22990);
and U24086 (N_24086,N_23398,N_22815);
and U24087 (N_24087,N_22754,N_23058);
nor U24088 (N_24088,N_23597,N_23169);
nor U24089 (N_24089,N_23625,N_22553);
or U24090 (N_24090,N_23014,N_23281);
nand U24091 (N_24091,N_22555,N_23080);
nor U24092 (N_24092,N_22977,N_23636);
xnor U24093 (N_24093,N_22735,N_22865);
nand U24094 (N_24094,N_23443,N_22504);
nor U24095 (N_24095,N_23559,N_23733);
xnor U24096 (N_24096,N_22653,N_23576);
or U24097 (N_24097,N_23317,N_23523);
nand U24098 (N_24098,N_23241,N_23225);
or U24099 (N_24099,N_23116,N_23069);
nand U24100 (N_24100,N_23341,N_23378);
or U24101 (N_24101,N_22766,N_22659);
or U24102 (N_24102,N_22650,N_23001);
nor U24103 (N_24103,N_23119,N_22939);
nand U24104 (N_24104,N_22917,N_23034);
or U24105 (N_24105,N_23598,N_22927);
and U24106 (N_24106,N_22976,N_22677);
and U24107 (N_24107,N_22943,N_22612);
or U24108 (N_24108,N_23115,N_23146);
nor U24109 (N_24109,N_22896,N_23160);
or U24110 (N_24110,N_22744,N_22916);
or U24111 (N_24111,N_23325,N_23534);
nand U24112 (N_24112,N_23189,N_22780);
and U24113 (N_24113,N_23118,N_22719);
nor U24114 (N_24114,N_23061,N_22627);
and U24115 (N_24115,N_22993,N_22828);
nand U24116 (N_24116,N_23070,N_23423);
nand U24117 (N_24117,N_23105,N_22913);
and U24118 (N_24118,N_23704,N_23021);
or U24119 (N_24119,N_22707,N_23719);
and U24120 (N_24120,N_22830,N_22582);
nor U24121 (N_24121,N_23517,N_23354);
and U24122 (N_24122,N_22974,N_23078);
xor U24123 (N_24123,N_23328,N_23698);
xor U24124 (N_24124,N_22538,N_23205);
nand U24125 (N_24125,N_23109,N_23436);
nand U24126 (N_24126,N_23267,N_23583);
nor U24127 (N_24127,N_23412,N_23288);
and U24128 (N_24128,N_23655,N_22920);
xnor U24129 (N_24129,N_23548,N_22911);
nand U24130 (N_24130,N_23355,N_23508);
or U24131 (N_24131,N_23507,N_23007);
nor U24132 (N_24132,N_23640,N_23556);
nor U24133 (N_24133,N_23682,N_22688);
nor U24134 (N_24134,N_22591,N_23321);
nand U24135 (N_24135,N_23740,N_23570);
xnor U24136 (N_24136,N_23330,N_23469);
and U24137 (N_24137,N_23038,N_22628);
xnor U24138 (N_24138,N_23633,N_22629);
nand U24139 (N_24139,N_22817,N_23229);
and U24140 (N_24140,N_23320,N_23725);
or U24141 (N_24141,N_22509,N_22632);
and U24142 (N_24142,N_23129,N_22678);
xnor U24143 (N_24143,N_23487,N_23127);
nor U24144 (N_24144,N_23474,N_22665);
xnor U24145 (N_24145,N_23227,N_22525);
nor U24146 (N_24146,N_22899,N_23075);
xnor U24147 (N_24147,N_23088,N_23132);
and U24148 (N_24148,N_22834,N_22765);
or U24149 (N_24149,N_22643,N_23390);
and U24150 (N_24150,N_23222,N_23418);
nor U24151 (N_24151,N_23595,N_23406);
nand U24152 (N_24152,N_23259,N_22960);
xnor U24153 (N_24153,N_23530,N_23741);
nand U24154 (N_24154,N_22746,N_23136);
nor U24155 (N_24155,N_22779,N_23463);
nor U24156 (N_24156,N_23365,N_22794);
nand U24157 (N_24157,N_23302,N_23333);
nor U24158 (N_24158,N_22587,N_22750);
and U24159 (N_24159,N_23367,N_23702);
nor U24160 (N_24160,N_22755,N_23068);
nand U24161 (N_24161,N_22737,N_23196);
xor U24162 (N_24162,N_23137,N_23607);
xor U24163 (N_24163,N_23519,N_23373);
or U24164 (N_24164,N_23159,N_23170);
and U24165 (N_24165,N_22980,N_23690);
xor U24166 (N_24166,N_23004,N_23357);
and U24167 (N_24167,N_23433,N_22649);
xor U24168 (N_24168,N_22910,N_23128);
xor U24169 (N_24169,N_22806,N_22796);
or U24170 (N_24170,N_22890,N_23561);
nand U24171 (N_24171,N_23179,N_23019);
nor U24172 (N_24172,N_23654,N_22534);
nand U24173 (N_24173,N_23114,N_22551);
nand U24174 (N_24174,N_23411,N_23031);
or U24175 (N_24175,N_23102,N_22907);
nand U24176 (N_24176,N_23226,N_22510);
or U24177 (N_24177,N_23405,N_23165);
nand U24178 (N_24178,N_22837,N_22680);
nand U24179 (N_24179,N_23223,N_23156);
or U24180 (N_24180,N_23659,N_22730);
nand U24181 (N_24181,N_22514,N_22997);
nor U24182 (N_24182,N_22902,N_23201);
or U24183 (N_24183,N_22702,N_22909);
xor U24184 (N_24184,N_23374,N_23265);
or U24185 (N_24185,N_23350,N_22800);
or U24186 (N_24186,N_22785,N_23605);
xor U24187 (N_24187,N_22877,N_23568);
and U24188 (N_24188,N_23526,N_23544);
and U24189 (N_24189,N_23574,N_23253);
nor U24190 (N_24190,N_23414,N_23500);
or U24191 (N_24191,N_23726,N_23063);
xnor U24192 (N_24192,N_23255,N_23113);
and U24193 (N_24193,N_23747,N_23520);
xor U24194 (N_24194,N_22752,N_22618);
nand U24195 (N_24195,N_23250,N_22634);
and U24196 (N_24196,N_23103,N_22743);
xor U24197 (N_24197,N_23244,N_23637);
xor U24198 (N_24198,N_23455,N_23283);
nand U24199 (N_24199,N_22963,N_23096);
nand U24200 (N_24200,N_23446,N_23669);
or U24201 (N_24201,N_23400,N_22835);
or U24202 (N_24202,N_23697,N_23217);
nor U24203 (N_24203,N_22852,N_23029);
nand U24204 (N_24204,N_23688,N_23557);
or U24205 (N_24205,N_22808,N_23456);
and U24206 (N_24206,N_23427,N_23489);
xnor U24207 (N_24207,N_23479,N_23008);
nand U24208 (N_24208,N_22751,N_23430);
and U24209 (N_24209,N_23587,N_23197);
xnor U24210 (N_24210,N_22623,N_23003);
xor U24211 (N_24211,N_23714,N_22840);
nor U24212 (N_24212,N_22764,N_23048);
nand U24213 (N_24213,N_22607,N_23064);
nand U24214 (N_24214,N_22500,N_22508);
xnor U24215 (N_24215,N_22901,N_23287);
nor U24216 (N_24216,N_22630,N_23657);
nor U24217 (N_24217,N_22542,N_22529);
or U24218 (N_24218,N_22889,N_22967);
or U24219 (N_24219,N_23195,N_22651);
and U24220 (N_24220,N_22956,N_23394);
nor U24221 (N_24221,N_22729,N_22805);
or U24222 (N_24222,N_22705,N_23383);
nor U24223 (N_24223,N_22641,N_23616);
nor U24224 (N_24224,N_22662,N_22550);
nor U24225 (N_24225,N_23466,N_23732);
xnor U24226 (N_24226,N_23239,N_23600);
and U24227 (N_24227,N_23028,N_23171);
xor U24228 (N_24228,N_23093,N_23645);
xor U24229 (N_24229,N_23693,N_23305);
nand U24230 (N_24230,N_23575,N_22965);
nand U24231 (N_24231,N_23679,N_23614);
nor U24232 (N_24232,N_23012,N_22674);
nor U24233 (N_24233,N_23503,N_23107);
nor U24234 (N_24234,N_22862,N_22855);
and U24235 (N_24235,N_23731,N_22679);
xnor U24236 (N_24236,N_23126,N_23152);
nor U24237 (N_24237,N_23543,N_23051);
and U24238 (N_24238,N_23428,N_22813);
nand U24239 (N_24239,N_23033,N_23449);
and U24240 (N_24240,N_23134,N_22526);
nand U24241 (N_24241,N_23319,N_23416);
and U24242 (N_24242,N_23464,N_22887);
xor U24243 (N_24243,N_22667,N_23477);
xnor U24244 (N_24244,N_23022,N_23024);
or U24245 (N_24245,N_22895,N_23720);
nor U24246 (N_24246,N_22503,N_23621);
and U24247 (N_24247,N_22979,N_22937);
nor U24248 (N_24248,N_22638,N_22733);
and U24249 (N_24249,N_23541,N_23566);
nor U24250 (N_24250,N_23708,N_23376);
nand U24251 (N_24251,N_23439,N_22731);
xnor U24252 (N_24252,N_22948,N_22769);
or U24253 (N_24253,N_22756,N_22546);
or U24254 (N_24254,N_22789,N_22599);
xnor U24255 (N_24255,N_23032,N_23145);
nand U24256 (N_24256,N_22866,N_22723);
xor U24257 (N_24257,N_23342,N_23444);
and U24258 (N_24258,N_23026,N_23248);
or U24259 (N_24259,N_23301,N_22799);
and U24260 (N_24260,N_22975,N_23448);
nor U24261 (N_24261,N_23072,N_22880);
and U24262 (N_24262,N_23174,N_23629);
or U24263 (N_24263,N_22941,N_22945);
nor U24264 (N_24264,N_22978,N_22548);
or U24265 (N_24265,N_23331,N_23238);
nor U24266 (N_24266,N_23327,N_23386);
nand U24267 (N_24267,N_23277,N_23699);
and U24268 (N_24268,N_23089,N_23363);
and U24269 (N_24269,N_22647,N_22652);
nor U24270 (N_24270,N_23385,N_23431);
nor U24271 (N_24271,N_23675,N_22968);
or U24272 (N_24272,N_22782,N_23295);
or U24273 (N_24273,N_23006,N_22556);
and U24274 (N_24274,N_22544,N_23215);
and U24275 (N_24275,N_23525,N_22573);
and U24276 (N_24276,N_22833,N_22823);
xnor U24277 (N_24277,N_23737,N_23264);
nand U24278 (N_24278,N_22926,N_23585);
nor U24279 (N_24279,N_22950,N_22522);
xor U24280 (N_24280,N_23191,N_23480);
nor U24281 (N_24281,N_23346,N_22639);
or U24282 (N_24282,N_22924,N_23420);
or U24283 (N_24283,N_22803,N_23123);
nor U24284 (N_24284,N_23361,N_23194);
nand U24285 (N_24285,N_23221,N_22658);
or U24286 (N_24286,N_23580,N_23524);
nand U24287 (N_24287,N_23368,N_23710);
nand U24288 (N_24288,N_23308,N_23488);
nand U24289 (N_24289,N_23074,N_22684);
xor U24290 (N_24290,N_23242,N_22620);
nor U24291 (N_24291,N_22695,N_23723);
or U24292 (N_24292,N_22788,N_23644);
or U24293 (N_24293,N_23471,N_23280);
nor U24294 (N_24294,N_23601,N_23736);
nand U24295 (N_24295,N_23647,N_23218);
or U24296 (N_24296,N_22519,N_23168);
or U24297 (N_24297,N_22614,N_23095);
or U24298 (N_24298,N_23015,N_23630);
nand U24299 (N_24299,N_23501,N_22547);
nor U24300 (N_24300,N_22592,N_23551);
nand U24301 (N_24301,N_23703,N_22566);
xnor U24302 (N_24302,N_23271,N_23210);
or U24303 (N_24303,N_22760,N_22637);
and U24304 (N_24304,N_23470,N_23299);
xnor U24305 (N_24305,N_23441,N_23546);
nor U24306 (N_24306,N_22501,N_22915);
nand U24307 (N_24307,N_23153,N_22668);
and U24308 (N_24308,N_23135,N_23744);
and U24309 (N_24309,N_22940,N_22574);
nand U24310 (N_24310,N_22825,N_22836);
nor U24311 (N_24311,N_22609,N_22528);
xor U24312 (N_24312,N_23315,N_22891);
nand U24313 (N_24313,N_23142,N_22689);
xnor U24314 (N_24314,N_23246,N_22868);
nand U24315 (N_24315,N_23323,N_23493);
xnor U24316 (N_24316,N_23590,N_23522);
nor U24317 (N_24317,N_22814,N_23011);
and U24318 (N_24318,N_23198,N_22906);
or U24319 (N_24319,N_22958,N_23252);
nand U24320 (N_24320,N_23060,N_22686);
xnor U24321 (N_24321,N_22699,N_23213);
and U24322 (N_24322,N_23421,N_23681);
nor U24323 (N_24323,N_22761,N_22793);
nand U24324 (N_24324,N_22787,N_23612);
or U24325 (N_24325,N_23705,N_22583);
xor U24326 (N_24326,N_23539,N_23155);
and U24327 (N_24327,N_22666,N_22954);
nand U24328 (N_24328,N_22897,N_23709);
nor U24329 (N_24329,N_23306,N_23071);
xnor U24330 (N_24330,N_23635,N_22515);
or U24331 (N_24331,N_23695,N_23490);
and U24332 (N_24332,N_23043,N_23482);
and U24333 (N_24333,N_22986,N_22798);
xnor U24334 (N_24334,N_23432,N_23245);
nor U24335 (N_24335,N_23036,N_23377);
nand U24336 (N_24336,N_22562,N_22984);
and U24337 (N_24337,N_23177,N_22989);
nand U24338 (N_24338,N_23513,N_23254);
nor U24339 (N_24339,N_22648,N_22962);
xor U24340 (N_24340,N_23453,N_22888);
or U24341 (N_24341,N_23158,N_23712);
nor U24342 (N_24342,N_22898,N_22961);
nor U24343 (N_24343,N_23272,N_23727);
nand U24344 (N_24344,N_23044,N_22681);
nor U24345 (N_24345,N_23592,N_22758);
xnor U24346 (N_24346,N_23665,N_23087);
and U24347 (N_24347,N_22903,N_22878);
nor U24348 (N_24348,N_23370,N_22786);
xor U24349 (N_24349,N_23653,N_23053);
xnor U24350 (N_24350,N_22944,N_22811);
nand U24351 (N_24351,N_23066,N_23643);
xnor U24352 (N_24352,N_23565,N_22717);
nor U24353 (N_24353,N_23055,N_22807);
nor U24354 (N_24354,N_22922,N_22869);
xor U24355 (N_24355,N_23748,N_23257);
or U24356 (N_24356,N_23670,N_22738);
or U24357 (N_24357,N_22698,N_22516);
nor U24358 (N_24358,N_23052,N_22675);
and U24359 (N_24359,N_23642,N_23359);
xnor U24360 (N_24360,N_23677,N_23092);
nor U24361 (N_24361,N_22770,N_23505);
nor U24362 (N_24362,N_23628,N_22568);
nand U24363 (N_24363,N_22635,N_22645);
xnor U24364 (N_24364,N_23273,N_23572);
and U24365 (N_24365,N_22664,N_22845);
or U24366 (N_24366,N_22821,N_22602);
nor U24367 (N_24367,N_22879,N_22929);
nor U24368 (N_24368,N_23057,N_22996);
or U24369 (N_24369,N_22725,N_23461);
nor U24370 (N_24370,N_23594,N_22908);
nand U24371 (N_24371,N_23631,N_22661);
xnor U24372 (N_24372,N_22541,N_23578);
nand U24373 (N_24373,N_23121,N_22857);
or U24374 (N_24374,N_22822,N_22657);
and U24375 (N_24375,N_22737,N_22802);
nand U24376 (N_24376,N_23531,N_23328);
nand U24377 (N_24377,N_22921,N_23624);
or U24378 (N_24378,N_22996,N_22650);
nor U24379 (N_24379,N_22670,N_23113);
xnor U24380 (N_24380,N_23111,N_23116);
nor U24381 (N_24381,N_22888,N_22742);
or U24382 (N_24382,N_22529,N_23294);
nor U24383 (N_24383,N_23392,N_22996);
xnor U24384 (N_24384,N_22704,N_22697);
xnor U24385 (N_24385,N_22661,N_23249);
and U24386 (N_24386,N_22615,N_22516);
xnor U24387 (N_24387,N_22606,N_23731);
xnor U24388 (N_24388,N_23251,N_23497);
nand U24389 (N_24389,N_23537,N_22504);
and U24390 (N_24390,N_22694,N_22881);
or U24391 (N_24391,N_23115,N_23472);
nor U24392 (N_24392,N_22829,N_22976);
or U24393 (N_24393,N_22958,N_22653);
and U24394 (N_24394,N_23707,N_23299);
nand U24395 (N_24395,N_22946,N_22822);
xnor U24396 (N_24396,N_23259,N_23188);
nor U24397 (N_24397,N_23265,N_22525);
nand U24398 (N_24398,N_22511,N_23144);
nand U24399 (N_24399,N_22847,N_22708);
and U24400 (N_24400,N_22881,N_22561);
nand U24401 (N_24401,N_23208,N_22644);
nand U24402 (N_24402,N_23146,N_23544);
xor U24403 (N_24403,N_22673,N_23545);
and U24404 (N_24404,N_22679,N_23299);
or U24405 (N_24405,N_22519,N_23434);
nor U24406 (N_24406,N_22948,N_23737);
nor U24407 (N_24407,N_22659,N_22543);
and U24408 (N_24408,N_22750,N_22718);
or U24409 (N_24409,N_23024,N_23455);
nand U24410 (N_24410,N_23622,N_22902);
and U24411 (N_24411,N_23191,N_23040);
xor U24412 (N_24412,N_23293,N_22663);
xor U24413 (N_24413,N_23517,N_23613);
or U24414 (N_24414,N_23559,N_23209);
xor U24415 (N_24415,N_23537,N_23360);
nand U24416 (N_24416,N_22923,N_22629);
and U24417 (N_24417,N_23642,N_23453);
xor U24418 (N_24418,N_23491,N_23400);
or U24419 (N_24419,N_23396,N_23473);
nand U24420 (N_24420,N_22687,N_22537);
xnor U24421 (N_24421,N_22937,N_23420);
and U24422 (N_24422,N_23288,N_23311);
xor U24423 (N_24423,N_23006,N_23117);
nor U24424 (N_24424,N_22831,N_22989);
and U24425 (N_24425,N_23463,N_22656);
xor U24426 (N_24426,N_23561,N_23283);
xor U24427 (N_24427,N_23281,N_23570);
nand U24428 (N_24428,N_22829,N_22696);
nand U24429 (N_24429,N_23127,N_22913);
or U24430 (N_24430,N_23673,N_23209);
xnor U24431 (N_24431,N_22757,N_22691);
or U24432 (N_24432,N_23651,N_23159);
nand U24433 (N_24433,N_23306,N_23302);
xor U24434 (N_24434,N_22901,N_23129);
nand U24435 (N_24435,N_22649,N_23180);
or U24436 (N_24436,N_23160,N_22503);
nand U24437 (N_24437,N_23303,N_23148);
or U24438 (N_24438,N_23117,N_22978);
and U24439 (N_24439,N_22594,N_23222);
nand U24440 (N_24440,N_23068,N_23736);
or U24441 (N_24441,N_23572,N_22986);
and U24442 (N_24442,N_23427,N_23412);
nand U24443 (N_24443,N_23191,N_23036);
or U24444 (N_24444,N_23028,N_22732);
or U24445 (N_24445,N_22921,N_23152);
or U24446 (N_24446,N_22755,N_23741);
xnor U24447 (N_24447,N_22725,N_23596);
nand U24448 (N_24448,N_23443,N_22815);
nand U24449 (N_24449,N_23498,N_22910);
xnor U24450 (N_24450,N_23239,N_22858);
or U24451 (N_24451,N_23172,N_22631);
nor U24452 (N_24452,N_23228,N_22910);
or U24453 (N_24453,N_23298,N_22788);
nor U24454 (N_24454,N_22630,N_22641);
or U24455 (N_24455,N_22650,N_22625);
nor U24456 (N_24456,N_22574,N_22606);
nand U24457 (N_24457,N_22914,N_22812);
and U24458 (N_24458,N_22747,N_23072);
or U24459 (N_24459,N_23611,N_22574);
or U24460 (N_24460,N_23084,N_23327);
or U24461 (N_24461,N_23180,N_22989);
and U24462 (N_24462,N_23450,N_23367);
nand U24463 (N_24463,N_22886,N_23232);
or U24464 (N_24464,N_23400,N_23622);
xor U24465 (N_24465,N_22808,N_23547);
and U24466 (N_24466,N_23404,N_23102);
nor U24467 (N_24467,N_22917,N_22812);
xor U24468 (N_24468,N_23218,N_23645);
or U24469 (N_24469,N_23342,N_22624);
nor U24470 (N_24470,N_23447,N_23526);
nand U24471 (N_24471,N_23133,N_23701);
nand U24472 (N_24472,N_22800,N_23341);
and U24473 (N_24473,N_23642,N_23631);
and U24474 (N_24474,N_23031,N_23214);
and U24475 (N_24475,N_23214,N_23737);
or U24476 (N_24476,N_23027,N_23268);
nor U24477 (N_24477,N_23529,N_22518);
nand U24478 (N_24478,N_22822,N_23275);
or U24479 (N_24479,N_23254,N_23718);
or U24480 (N_24480,N_22878,N_23601);
nand U24481 (N_24481,N_22785,N_23540);
and U24482 (N_24482,N_23251,N_23312);
or U24483 (N_24483,N_22764,N_23702);
and U24484 (N_24484,N_22818,N_23018);
or U24485 (N_24485,N_23336,N_22871);
or U24486 (N_24486,N_22712,N_22855);
nor U24487 (N_24487,N_23443,N_23482);
nand U24488 (N_24488,N_23050,N_22553);
or U24489 (N_24489,N_23157,N_22688);
xor U24490 (N_24490,N_22830,N_22736);
or U24491 (N_24491,N_23219,N_22545);
and U24492 (N_24492,N_23438,N_22529);
xnor U24493 (N_24493,N_22656,N_22586);
or U24494 (N_24494,N_23446,N_22932);
or U24495 (N_24495,N_22539,N_23101);
xnor U24496 (N_24496,N_22960,N_22565);
nor U24497 (N_24497,N_22955,N_23107);
or U24498 (N_24498,N_23251,N_23169);
nand U24499 (N_24499,N_23594,N_23068);
or U24500 (N_24500,N_23502,N_23030);
or U24501 (N_24501,N_22979,N_23384);
or U24502 (N_24502,N_23457,N_22598);
nand U24503 (N_24503,N_22971,N_22998);
xnor U24504 (N_24504,N_23240,N_22698);
nor U24505 (N_24505,N_22706,N_22531);
nand U24506 (N_24506,N_22580,N_23029);
nor U24507 (N_24507,N_22750,N_23182);
or U24508 (N_24508,N_22759,N_23077);
xor U24509 (N_24509,N_22500,N_22619);
and U24510 (N_24510,N_23474,N_22844);
nor U24511 (N_24511,N_23412,N_23342);
and U24512 (N_24512,N_22877,N_23287);
nand U24513 (N_24513,N_22754,N_23060);
or U24514 (N_24514,N_22955,N_22601);
xor U24515 (N_24515,N_23636,N_23719);
and U24516 (N_24516,N_23581,N_22979);
or U24517 (N_24517,N_23429,N_22514);
xnor U24518 (N_24518,N_23725,N_23173);
and U24519 (N_24519,N_22697,N_22933);
and U24520 (N_24520,N_23458,N_22615);
nand U24521 (N_24521,N_23154,N_23096);
and U24522 (N_24522,N_22984,N_23002);
xor U24523 (N_24523,N_23078,N_22623);
nand U24524 (N_24524,N_22841,N_23477);
xnor U24525 (N_24525,N_23495,N_23537);
or U24526 (N_24526,N_22644,N_23608);
nand U24527 (N_24527,N_22833,N_23058);
and U24528 (N_24528,N_23175,N_22589);
xor U24529 (N_24529,N_22500,N_22970);
or U24530 (N_24530,N_22773,N_23730);
nand U24531 (N_24531,N_22905,N_23502);
and U24532 (N_24532,N_23307,N_23078);
nand U24533 (N_24533,N_22800,N_22695);
nor U24534 (N_24534,N_23366,N_22617);
or U24535 (N_24535,N_23720,N_23350);
nand U24536 (N_24536,N_23582,N_22948);
and U24537 (N_24537,N_23304,N_22822);
nor U24538 (N_24538,N_23625,N_23172);
xor U24539 (N_24539,N_23567,N_22785);
nor U24540 (N_24540,N_22982,N_23402);
nand U24541 (N_24541,N_23566,N_22909);
nand U24542 (N_24542,N_22872,N_22565);
nand U24543 (N_24543,N_23666,N_23454);
nor U24544 (N_24544,N_22531,N_23537);
nor U24545 (N_24545,N_23016,N_22780);
and U24546 (N_24546,N_22656,N_22565);
or U24547 (N_24547,N_23089,N_22918);
xnor U24548 (N_24548,N_23218,N_23270);
and U24549 (N_24549,N_23399,N_23233);
or U24550 (N_24550,N_23598,N_23626);
or U24551 (N_24551,N_23141,N_22994);
nand U24552 (N_24552,N_23434,N_22921);
nand U24553 (N_24553,N_23139,N_22878);
xnor U24554 (N_24554,N_23625,N_22850);
or U24555 (N_24555,N_23068,N_23634);
xor U24556 (N_24556,N_23041,N_23423);
nand U24557 (N_24557,N_23683,N_22668);
or U24558 (N_24558,N_23535,N_22956);
nand U24559 (N_24559,N_23367,N_23073);
and U24560 (N_24560,N_23256,N_23568);
and U24561 (N_24561,N_23469,N_23030);
or U24562 (N_24562,N_22501,N_23047);
or U24563 (N_24563,N_23049,N_23429);
and U24564 (N_24564,N_22885,N_23304);
nand U24565 (N_24565,N_23455,N_23329);
xnor U24566 (N_24566,N_22657,N_22766);
and U24567 (N_24567,N_23228,N_23016);
and U24568 (N_24568,N_23349,N_23335);
nand U24569 (N_24569,N_22781,N_23270);
or U24570 (N_24570,N_23508,N_23627);
xor U24571 (N_24571,N_23040,N_23697);
nand U24572 (N_24572,N_23608,N_23066);
or U24573 (N_24573,N_23178,N_23590);
nand U24574 (N_24574,N_22652,N_23113);
nor U24575 (N_24575,N_23395,N_23116);
nand U24576 (N_24576,N_23679,N_23473);
xnor U24577 (N_24577,N_23263,N_23275);
xnor U24578 (N_24578,N_22631,N_23133);
or U24579 (N_24579,N_23326,N_23504);
nor U24580 (N_24580,N_22593,N_23071);
nor U24581 (N_24581,N_23657,N_22919);
xor U24582 (N_24582,N_23695,N_23405);
xnor U24583 (N_24583,N_22664,N_22714);
xnor U24584 (N_24584,N_23414,N_23675);
nand U24585 (N_24585,N_23182,N_23084);
and U24586 (N_24586,N_23330,N_23008);
and U24587 (N_24587,N_23364,N_23029);
or U24588 (N_24588,N_23601,N_22724);
nor U24589 (N_24589,N_22668,N_22607);
nor U24590 (N_24590,N_23350,N_23613);
xnor U24591 (N_24591,N_22655,N_22798);
nor U24592 (N_24592,N_22834,N_23426);
or U24593 (N_24593,N_22538,N_22693);
or U24594 (N_24594,N_23410,N_23491);
nor U24595 (N_24595,N_23377,N_22584);
nor U24596 (N_24596,N_22804,N_23193);
xor U24597 (N_24597,N_23555,N_22530);
nand U24598 (N_24598,N_23119,N_22512);
and U24599 (N_24599,N_22968,N_23358);
nor U24600 (N_24600,N_22756,N_23446);
xor U24601 (N_24601,N_23441,N_22892);
nand U24602 (N_24602,N_23450,N_22932);
or U24603 (N_24603,N_22931,N_23702);
and U24604 (N_24604,N_22837,N_23126);
or U24605 (N_24605,N_23678,N_22602);
or U24606 (N_24606,N_23168,N_22850);
and U24607 (N_24607,N_23356,N_22839);
or U24608 (N_24608,N_23244,N_23087);
and U24609 (N_24609,N_22836,N_23147);
xnor U24610 (N_24610,N_22703,N_23101);
or U24611 (N_24611,N_23434,N_23522);
xnor U24612 (N_24612,N_23095,N_22605);
and U24613 (N_24613,N_23739,N_23749);
nor U24614 (N_24614,N_22719,N_23513);
or U24615 (N_24615,N_23590,N_23194);
nor U24616 (N_24616,N_23646,N_23171);
and U24617 (N_24617,N_23623,N_23416);
and U24618 (N_24618,N_22839,N_22773);
nor U24619 (N_24619,N_23644,N_22864);
and U24620 (N_24620,N_22648,N_22848);
nor U24621 (N_24621,N_22820,N_23721);
nand U24622 (N_24622,N_22535,N_23470);
or U24623 (N_24623,N_23640,N_22641);
nor U24624 (N_24624,N_22587,N_22557);
nand U24625 (N_24625,N_23600,N_23675);
or U24626 (N_24626,N_23671,N_23242);
nor U24627 (N_24627,N_23291,N_22746);
xor U24628 (N_24628,N_22957,N_23718);
xor U24629 (N_24629,N_23292,N_22815);
and U24630 (N_24630,N_23729,N_22947);
nor U24631 (N_24631,N_23744,N_22654);
and U24632 (N_24632,N_23160,N_23051);
xnor U24633 (N_24633,N_23025,N_22602);
nor U24634 (N_24634,N_23644,N_22868);
xnor U24635 (N_24635,N_22577,N_23152);
or U24636 (N_24636,N_23320,N_22963);
nor U24637 (N_24637,N_23419,N_23285);
xor U24638 (N_24638,N_23063,N_23432);
xnor U24639 (N_24639,N_22531,N_22925);
nor U24640 (N_24640,N_22860,N_23545);
or U24641 (N_24641,N_22720,N_23554);
or U24642 (N_24642,N_23572,N_22588);
xnor U24643 (N_24643,N_23088,N_23238);
and U24644 (N_24644,N_22557,N_22619);
nand U24645 (N_24645,N_23616,N_23078);
xnor U24646 (N_24646,N_23451,N_23239);
nand U24647 (N_24647,N_23470,N_23365);
xnor U24648 (N_24648,N_22991,N_22563);
nand U24649 (N_24649,N_23442,N_23383);
xnor U24650 (N_24650,N_23204,N_22981);
and U24651 (N_24651,N_23176,N_23617);
or U24652 (N_24652,N_23316,N_23063);
and U24653 (N_24653,N_23437,N_22892);
nand U24654 (N_24654,N_22560,N_22543);
nor U24655 (N_24655,N_23368,N_22861);
nand U24656 (N_24656,N_23729,N_22789);
nor U24657 (N_24657,N_22877,N_23235);
nor U24658 (N_24658,N_23288,N_22990);
nand U24659 (N_24659,N_23337,N_23537);
and U24660 (N_24660,N_23349,N_23425);
xnor U24661 (N_24661,N_22735,N_22861);
nor U24662 (N_24662,N_23377,N_23723);
and U24663 (N_24663,N_23585,N_22751);
nand U24664 (N_24664,N_23453,N_23349);
nor U24665 (N_24665,N_23531,N_22561);
nor U24666 (N_24666,N_23660,N_23378);
nor U24667 (N_24667,N_23150,N_22776);
or U24668 (N_24668,N_22885,N_23057);
nor U24669 (N_24669,N_23193,N_23499);
xor U24670 (N_24670,N_22582,N_23342);
nor U24671 (N_24671,N_23462,N_22675);
or U24672 (N_24672,N_23091,N_23691);
or U24673 (N_24673,N_23567,N_22695);
nor U24674 (N_24674,N_23355,N_23373);
nand U24675 (N_24675,N_22774,N_22528);
nor U24676 (N_24676,N_23216,N_22861);
nor U24677 (N_24677,N_22865,N_23445);
and U24678 (N_24678,N_23435,N_22992);
xnor U24679 (N_24679,N_22686,N_23596);
xor U24680 (N_24680,N_23415,N_23688);
nand U24681 (N_24681,N_22867,N_23558);
xor U24682 (N_24682,N_23347,N_22717);
nand U24683 (N_24683,N_23082,N_22887);
and U24684 (N_24684,N_23479,N_22788);
nor U24685 (N_24685,N_22954,N_22979);
or U24686 (N_24686,N_22834,N_22819);
and U24687 (N_24687,N_23326,N_22954);
or U24688 (N_24688,N_23178,N_22926);
nand U24689 (N_24689,N_23196,N_23118);
nor U24690 (N_24690,N_23605,N_22925);
nor U24691 (N_24691,N_22567,N_22989);
and U24692 (N_24692,N_23452,N_23466);
or U24693 (N_24693,N_23602,N_22695);
or U24694 (N_24694,N_23046,N_23345);
nand U24695 (N_24695,N_23568,N_23238);
nand U24696 (N_24696,N_23131,N_23448);
and U24697 (N_24697,N_23050,N_23094);
nor U24698 (N_24698,N_23331,N_23631);
xnor U24699 (N_24699,N_22728,N_23392);
nor U24700 (N_24700,N_23490,N_23261);
nand U24701 (N_24701,N_22799,N_22795);
or U24702 (N_24702,N_22534,N_23194);
xnor U24703 (N_24703,N_23723,N_23159);
nor U24704 (N_24704,N_22975,N_23609);
and U24705 (N_24705,N_22574,N_23507);
nor U24706 (N_24706,N_23145,N_23390);
nor U24707 (N_24707,N_23491,N_23747);
or U24708 (N_24708,N_23442,N_22745);
nand U24709 (N_24709,N_22600,N_22756);
nor U24710 (N_24710,N_23291,N_23402);
xnor U24711 (N_24711,N_23417,N_22730);
and U24712 (N_24712,N_22701,N_23334);
and U24713 (N_24713,N_22628,N_22692);
and U24714 (N_24714,N_23400,N_23152);
or U24715 (N_24715,N_22983,N_22612);
and U24716 (N_24716,N_23465,N_23551);
nand U24717 (N_24717,N_22547,N_23480);
or U24718 (N_24718,N_22909,N_22723);
and U24719 (N_24719,N_22995,N_23547);
xnor U24720 (N_24720,N_23304,N_22681);
or U24721 (N_24721,N_22868,N_23163);
and U24722 (N_24722,N_23182,N_22924);
nand U24723 (N_24723,N_22672,N_22802);
xnor U24724 (N_24724,N_23176,N_22905);
or U24725 (N_24725,N_23228,N_23583);
or U24726 (N_24726,N_22533,N_22745);
xnor U24727 (N_24727,N_23043,N_22845);
and U24728 (N_24728,N_22713,N_23580);
nand U24729 (N_24729,N_22915,N_23676);
xor U24730 (N_24730,N_22681,N_22521);
nand U24731 (N_24731,N_23590,N_23686);
and U24732 (N_24732,N_23385,N_23616);
and U24733 (N_24733,N_23510,N_23118);
nor U24734 (N_24734,N_23634,N_22897);
or U24735 (N_24735,N_23252,N_23686);
nor U24736 (N_24736,N_22591,N_23718);
or U24737 (N_24737,N_23119,N_23363);
xor U24738 (N_24738,N_23450,N_22931);
and U24739 (N_24739,N_22899,N_23390);
or U24740 (N_24740,N_22541,N_22851);
nand U24741 (N_24741,N_22629,N_22978);
nor U24742 (N_24742,N_23407,N_23621);
xor U24743 (N_24743,N_23268,N_22551);
and U24744 (N_24744,N_23311,N_22759);
or U24745 (N_24745,N_23226,N_23119);
xor U24746 (N_24746,N_22906,N_23698);
xor U24747 (N_24747,N_22611,N_23684);
or U24748 (N_24748,N_23536,N_22755);
nand U24749 (N_24749,N_22890,N_22520);
xor U24750 (N_24750,N_23101,N_22540);
nand U24751 (N_24751,N_22973,N_22987);
nand U24752 (N_24752,N_23604,N_23051);
nand U24753 (N_24753,N_22500,N_23538);
or U24754 (N_24754,N_23441,N_22884);
or U24755 (N_24755,N_23515,N_23356);
and U24756 (N_24756,N_23391,N_23597);
or U24757 (N_24757,N_23442,N_23070);
or U24758 (N_24758,N_23660,N_23352);
nand U24759 (N_24759,N_23084,N_22588);
nand U24760 (N_24760,N_23428,N_22607);
nand U24761 (N_24761,N_22821,N_23160);
nand U24762 (N_24762,N_23687,N_23654);
xnor U24763 (N_24763,N_23552,N_23117);
xnor U24764 (N_24764,N_22623,N_23722);
xnor U24765 (N_24765,N_23705,N_23478);
nand U24766 (N_24766,N_22516,N_22811);
xor U24767 (N_24767,N_23586,N_23417);
nand U24768 (N_24768,N_23741,N_23075);
nand U24769 (N_24769,N_22713,N_23623);
and U24770 (N_24770,N_23551,N_22959);
or U24771 (N_24771,N_22674,N_22561);
xor U24772 (N_24772,N_22709,N_23005);
and U24773 (N_24773,N_23106,N_22571);
nor U24774 (N_24774,N_23129,N_22751);
nor U24775 (N_24775,N_23340,N_23133);
or U24776 (N_24776,N_22574,N_22521);
and U24777 (N_24777,N_23071,N_22896);
or U24778 (N_24778,N_22626,N_22642);
nand U24779 (N_24779,N_23047,N_23177);
nor U24780 (N_24780,N_23205,N_22568);
xor U24781 (N_24781,N_23281,N_22948);
nand U24782 (N_24782,N_22674,N_22874);
or U24783 (N_24783,N_22981,N_22944);
and U24784 (N_24784,N_23365,N_23630);
or U24785 (N_24785,N_22778,N_22585);
nand U24786 (N_24786,N_22603,N_23317);
nand U24787 (N_24787,N_22764,N_23279);
nand U24788 (N_24788,N_22592,N_22542);
xnor U24789 (N_24789,N_23247,N_23162);
nand U24790 (N_24790,N_22692,N_22635);
nor U24791 (N_24791,N_23207,N_22755);
nand U24792 (N_24792,N_23215,N_23137);
nand U24793 (N_24793,N_23424,N_23315);
nor U24794 (N_24794,N_23409,N_22663);
or U24795 (N_24795,N_23117,N_23565);
or U24796 (N_24796,N_23736,N_23478);
nor U24797 (N_24797,N_22607,N_23357);
nand U24798 (N_24798,N_22570,N_23533);
and U24799 (N_24799,N_22607,N_22724);
nand U24800 (N_24800,N_22915,N_23321);
nor U24801 (N_24801,N_23236,N_23230);
xor U24802 (N_24802,N_23549,N_22797);
or U24803 (N_24803,N_23410,N_22775);
xor U24804 (N_24804,N_23667,N_23156);
and U24805 (N_24805,N_23210,N_22858);
and U24806 (N_24806,N_23340,N_23098);
nand U24807 (N_24807,N_22757,N_23277);
xor U24808 (N_24808,N_23299,N_23077);
or U24809 (N_24809,N_22774,N_23031);
xnor U24810 (N_24810,N_23584,N_23286);
xor U24811 (N_24811,N_23007,N_23665);
xor U24812 (N_24812,N_22524,N_22969);
nand U24813 (N_24813,N_23452,N_23105);
and U24814 (N_24814,N_22790,N_23377);
nand U24815 (N_24815,N_22756,N_22849);
and U24816 (N_24816,N_23188,N_22521);
and U24817 (N_24817,N_23330,N_23183);
xor U24818 (N_24818,N_22829,N_23547);
and U24819 (N_24819,N_23623,N_23053);
nor U24820 (N_24820,N_23046,N_23678);
and U24821 (N_24821,N_23310,N_23696);
and U24822 (N_24822,N_22690,N_22741);
or U24823 (N_24823,N_23673,N_23319);
nand U24824 (N_24824,N_23451,N_23034);
nor U24825 (N_24825,N_23616,N_22748);
and U24826 (N_24826,N_22631,N_23099);
nand U24827 (N_24827,N_23118,N_23464);
and U24828 (N_24828,N_23566,N_22885);
nor U24829 (N_24829,N_23353,N_22915);
nand U24830 (N_24830,N_23113,N_23134);
nor U24831 (N_24831,N_23141,N_22640);
nor U24832 (N_24832,N_22651,N_23735);
or U24833 (N_24833,N_22515,N_23552);
and U24834 (N_24834,N_22736,N_22856);
xor U24835 (N_24835,N_23691,N_22553);
or U24836 (N_24836,N_23528,N_22996);
or U24837 (N_24837,N_23366,N_23144);
xnor U24838 (N_24838,N_23673,N_22837);
and U24839 (N_24839,N_22934,N_23250);
and U24840 (N_24840,N_22793,N_22701);
nor U24841 (N_24841,N_23060,N_22615);
nor U24842 (N_24842,N_22803,N_23287);
or U24843 (N_24843,N_23233,N_23311);
nand U24844 (N_24844,N_23091,N_23110);
xnor U24845 (N_24845,N_22553,N_23634);
xnor U24846 (N_24846,N_23420,N_22540);
xnor U24847 (N_24847,N_22960,N_23507);
xnor U24848 (N_24848,N_23727,N_23690);
nor U24849 (N_24849,N_23298,N_23357);
xnor U24850 (N_24850,N_23505,N_22788);
nor U24851 (N_24851,N_23405,N_23201);
nor U24852 (N_24852,N_23307,N_23649);
nand U24853 (N_24853,N_22507,N_23550);
nand U24854 (N_24854,N_22982,N_23166);
and U24855 (N_24855,N_23491,N_22756);
xnor U24856 (N_24856,N_23476,N_23009);
or U24857 (N_24857,N_22641,N_23620);
or U24858 (N_24858,N_23366,N_23369);
nand U24859 (N_24859,N_23210,N_22503);
xnor U24860 (N_24860,N_22556,N_23410);
and U24861 (N_24861,N_23553,N_23069);
nand U24862 (N_24862,N_23561,N_22744);
xor U24863 (N_24863,N_22658,N_22789);
nand U24864 (N_24864,N_23139,N_23690);
nor U24865 (N_24865,N_22861,N_23134);
nor U24866 (N_24866,N_23275,N_23639);
and U24867 (N_24867,N_23187,N_22977);
or U24868 (N_24868,N_23422,N_22965);
or U24869 (N_24869,N_22816,N_23291);
and U24870 (N_24870,N_23000,N_22981);
nor U24871 (N_24871,N_22548,N_22584);
nand U24872 (N_24872,N_22585,N_23061);
and U24873 (N_24873,N_23486,N_23146);
and U24874 (N_24874,N_22563,N_22587);
or U24875 (N_24875,N_23576,N_23633);
and U24876 (N_24876,N_23166,N_23381);
and U24877 (N_24877,N_22837,N_23318);
or U24878 (N_24878,N_23121,N_23472);
and U24879 (N_24879,N_23715,N_23192);
or U24880 (N_24880,N_22843,N_23581);
nor U24881 (N_24881,N_23039,N_23220);
nor U24882 (N_24882,N_23280,N_22979);
nand U24883 (N_24883,N_22901,N_23103);
nand U24884 (N_24884,N_23306,N_22708);
nor U24885 (N_24885,N_22728,N_23125);
or U24886 (N_24886,N_23643,N_22706);
nand U24887 (N_24887,N_23308,N_22768);
xor U24888 (N_24888,N_23608,N_22729);
nor U24889 (N_24889,N_23612,N_22601);
nor U24890 (N_24890,N_22672,N_22695);
or U24891 (N_24891,N_23290,N_22542);
nor U24892 (N_24892,N_22510,N_23634);
or U24893 (N_24893,N_22827,N_23331);
or U24894 (N_24894,N_22793,N_23169);
nand U24895 (N_24895,N_23161,N_23649);
nor U24896 (N_24896,N_22927,N_23211);
or U24897 (N_24897,N_23396,N_22818);
xnor U24898 (N_24898,N_23368,N_23430);
and U24899 (N_24899,N_22647,N_22698);
nand U24900 (N_24900,N_22683,N_23301);
and U24901 (N_24901,N_22613,N_22927);
nor U24902 (N_24902,N_22518,N_23703);
or U24903 (N_24903,N_22733,N_22754);
xor U24904 (N_24904,N_23247,N_23735);
or U24905 (N_24905,N_22513,N_23130);
and U24906 (N_24906,N_23476,N_23613);
nand U24907 (N_24907,N_23739,N_23208);
nand U24908 (N_24908,N_22916,N_23232);
or U24909 (N_24909,N_23687,N_22802);
nor U24910 (N_24910,N_22800,N_23410);
nand U24911 (N_24911,N_23217,N_23047);
nand U24912 (N_24912,N_22849,N_23384);
or U24913 (N_24913,N_22814,N_23172);
xor U24914 (N_24914,N_23043,N_23306);
nor U24915 (N_24915,N_23167,N_23231);
xnor U24916 (N_24916,N_23567,N_23477);
and U24917 (N_24917,N_22731,N_23244);
and U24918 (N_24918,N_23320,N_23302);
and U24919 (N_24919,N_22833,N_23352);
xnor U24920 (N_24920,N_23379,N_22933);
nor U24921 (N_24921,N_23197,N_23661);
xor U24922 (N_24922,N_22661,N_22948);
or U24923 (N_24923,N_23043,N_22639);
or U24924 (N_24924,N_22529,N_22916);
xnor U24925 (N_24925,N_22537,N_22614);
xor U24926 (N_24926,N_23487,N_23427);
or U24927 (N_24927,N_22985,N_22526);
xnor U24928 (N_24928,N_23744,N_22722);
nor U24929 (N_24929,N_23312,N_23055);
nor U24930 (N_24930,N_23544,N_23399);
xor U24931 (N_24931,N_22560,N_23336);
or U24932 (N_24932,N_22739,N_23331);
xor U24933 (N_24933,N_23673,N_23566);
and U24934 (N_24934,N_22783,N_22594);
nor U24935 (N_24935,N_23515,N_23068);
and U24936 (N_24936,N_23186,N_22873);
nor U24937 (N_24937,N_22844,N_23345);
and U24938 (N_24938,N_23720,N_23020);
nor U24939 (N_24939,N_23606,N_22854);
xnor U24940 (N_24940,N_22573,N_22550);
nand U24941 (N_24941,N_23315,N_22702);
or U24942 (N_24942,N_23091,N_22732);
xor U24943 (N_24943,N_23308,N_22655);
nor U24944 (N_24944,N_22928,N_23045);
nor U24945 (N_24945,N_22970,N_22653);
nand U24946 (N_24946,N_23175,N_23558);
xor U24947 (N_24947,N_22848,N_22758);
and U24948 (N_24948,N_23616,N_23166);
nand U24949 (N_24949,N_23452,N_23545);
nand U24950 (N_24950,N_23513,N_23402);
or U24951 (N_24951,N_22729,N_22568);
nor U24952 (N_24952,N_22838,N_23725);
nor U24953 (N_24953,N_23509,N_23555);
nand U24954 (N_24954,N_22823,N_22622);
and U24955 (N_24955,N_22895,N_23034);
xor U24956 (N_24956,N_23367,N_23049);
and U24957 (N_24957,N_22983,N_22794);
xor U24958 (N_24958,N_23748,N_23535);
xor U24959 (N_24959,N_23097,N_23622);
and U24960 (N_24960,N_22645,N_22553);
and U24961 (N_24961,N_22622,N_22924);
nor U24962 (N_24962,N_23430,N_23583);
and U24963 (N_24963,N_22769,N_22543);
nor U24964 (N_24964,N_22789,N_23511);
xnor U24965 (N_24965,N_23144,N_23367);
xor U24966 (N_24966,N_23304,N_22920);
and U24967 (N_24967,N_23447,N_23737);
xor U24968 (N_24968,N_23207,N_22665);
xnor U24969 (N_24969,N_23510,N_22932);
nand U24970 (N_24970,N_23219,N_22727);
or U24971 (N_24971,N_23573,N_22582);
xnor U24972 (N_24972,N_22512,N_23143);
nor U24973 (N_24973,N_23082,N_23219);
xor U24974 (N_24974,N_22563,N_23459);
nor U24975 (N_24975,N_22723,N_23395);
nor U24976 (N_24976,N_23469,N_22661);
nor U24977 (N_24977,N_23225,N_23586);
or U24978 (N_24978,N_23161,N_23002);
or U24979 (N_24979,N_22520,N_22620);
or U24980 (N_24980,N_22773,N_22845);
xor U24981 (N_24981,N_23045,N_23401);
or U24982 (N_24982,N_22929,N_22847);
or U24983 (N_24983,N_23264,N_23100);
and U24984 (N_24984,N_23059,N_22619);
and U24985 (N_24985,N_23676,N_22852);
or U24986 (N_24986,N_23062,N_23695);
xor U24987 (N_24987,N_23118,N_23643);
or U24988 (N_24988,N_22527,N_23131);
or U24989 (N_24989,N_23312,N_22560);
nand U24990 (N_24990,N_23613,N_23399);
or U24991 (N_24991,N_22587,N_23184);
xnor U24992 (N_24992,N_23173,N_22787);
or U24993 (N_24993,N_23370,N_23506);
nor U24994 (N_24994,N_23054,N_23529);
nand U24995 (N_24995,N_22863,N_23193);
xnor U24996 (N_24996,N_23250,N_23710);
xnor U24997 (N_24997,N_23225,N_22884);
nand U24998 (N_24998,N_22777,N_22954);
and U24999 (N_24999,N_22536,N_22773);
nand UO_0 (O_0,N_24722,N_24021);
and UO_1 (O_1,N_24554,N_24429);
nand UO_2 (O_2,N_24744,N_23921);
nor UO_3 (O_3,N_23915,N_24896);
xor UO_4 (O_4,N_24037,N_24934);
xor UO_5 (O_5,N_24854,N_24797);
or UO_6 (O_6,N_24424,N_23975);
nand UO_7 (O_7,N_24386,N_24763);
or UO_8 (O_8,N_24053,N_24309);
or UO_9 (O_9,N_24777,N_24518);
and UO_10 (O_10,N_24732,N_24778);
and UO_11 (O_11,N_24809,N_24653);
or UO_12 (O_12,N_24752,N_23978);
nor UO_13 (O_13,N_24709,N_24378);
nor UO_14 (O_14,N_24706,N_24750);
or UO_15 (O_15,N_24235,N_24676);
and UO_16 (O_16,N_24137,N_24519);
or UO_17 (O_17,N_24263,N_24132);
and UO_18 (O_18,N_24177,N_24087);
nor UO_19 (O_19,N_23785,N_24899);
nand UO_20 (O_20,N_24320,N_24463);
and UO_21 (O_21,N_24115,N_24711);
or UO_22 (O_22,N_24344,N_24028);
nor UO_23 (O_23,N_23814,N_24611);
nor UO_24 (O_24,N_24216,N_24520);
or UO_25 (O_25,N_24567,N_24033);
or UO_26 (O_26,N_24716,N_23988);
nand UO_27 (O_27,N_24580,N_24764);
and UO_28 (O_28,N_24472,N_24772);
nor UO_29 (O_29,N_24039,N_24907);
nand UO_30 (O_30,N_24470,N_23926);
nor UO_31 (O_31,N_24064,N_24274);
nand UO_32 (O_32,N_24984,N_24484);
and UO_33 (O_33,N_23910,N_24953);
nor UO_34 (O_34,N_23872,N_23912);
and UO_35 (O_35,N_24566,N_24747);
xnor UO_36 (O_36,N_23962,N_24074);
nor UO_37 (O_37,N_23781,N_24831);
and UO_38 (O_38,N_24393,N_24371);
xor UO_39 (O_39,N_24635,N_24718);
nor UO_40 (O_40,N_24364,N_23955);
nand UO_41 (O_41,N_24333,N_24766);
and UO_42 (O_42,N_23974,N_24169);
and UO_43 (O_43,N_24358,N_23956);
nand UO_44 (O_44,N_24650,N_24858);
or UO_45 (O_45,N_24079,N_24691);
or UO_46 (O_46,N_24803,N_24278);
or UO_47 (O_47,N_24806,N_24419);
or UO_48 (O_48,N_24559,N_23854);
nand UO_49 (O_49,N_24590,N_24546);
or UO_50 (O_50,N_23901,N_24671);
xor UO_51 (O_51,N_23755,N_23971);
or UO_52 (O_52,N_24724,N_24659);
xor UO_53 (O_53,N_24893,N_23940);
nand UO_54 (O_54,N_23900,N_24909);
xnor UO_55 (O_55,N_24459,N_24946);
nor UO_56 (O_56,N_23809,N_24765);
nand UO_57 (O_57,N_24636,N_24193);
xnor UO_58 (O_58,N_24355,N_23994);
xnor UO_59 (O_59,N_23906,N_23796);
nor UO_60 (O_60,N_24295,N_23864);
or UO_61 (O_61,N_24703,N_23946);
or UO_62 (O_62,N_24890,N_23892);
nor UO_63 (O_63,N_24160,N_23977);
or UO_64 (O_64,N_23983,N_24867);
xor UO_65 (O_65,N_24165,N_24754);
and UO_66 (O_66,N_24989,N_24599);
or UO_67 (O_67,N_24618,N_24849);
nor UO_68 (O_68,N_24434,N_24349);
nor UO_69 (O_69,N_23758,N_24439);
or UO_70 (O_70,N_23986,N_24385);
nand UO_71 (O_71,N_24258,N_23828);
nand UO_72 (O_72,N_24904,N_24242);
xnor UO_73 (O_73,N_24810,N_24297);
nor UO_74 (O_74,N_24886,N_24897);
and UO_75 (O_75,N_24197,N_24228);
and UO_76 (O_76,N_24960,N_23839);
nor UO_77 (O_77,N_24964,N_24581);
nand UO_78 (O_78,N_24374,N_24432);
xor UO_79 (O_79,N_24129,N_23862);
xor UO_80 (O_80,N_24102,N_24044);
nand UO_81 (O_81,N_24638,N_24577);
nor UO_82 (O_82,N_24503,N_24479);
nand UO_83 (O_83,N_24512,N_23858);
or UO_84 (O_84,N_24663,N_24642);
nand UO_85 (O_85,N_24623,N_23855);
xnor UO_86 (O_86,N_24875,N_24549);
or UO_87 (O_87,N_24668,N_24633);
nor UO_88 (O_88,N_24521,N_24413);
xor UO_89 (O_89,N_24713,N_24931);
and UO_90 (O_90,N_24701,N_23762);
or UO_91 (O_91,N_24901,N_24001);
nor UO_92 (O_92,N_24843,N_24330);
or UO_93 (O_93,N_24200,N_24202);
nand UO_94 (O_94,N_23919,N_23846);
nand UO_95 (O_95,N_24687,N_24558);
or UO_96 (O_96,N_23773,N_24194);
nor UO_97 (O_97,N_24510,N_24442);
and UO_98 (O_98,N_24234,N_24773);
xnor UO_99 (O_99,N_24625,N_24878);
xnor UO_100 (O_100,N_24277,N_24133);
nand UO_101 (O_101,N_24070,N_24226);
nand UO_102 (O_102,N_24485,N_23776);
nand UO_103 (O_103,N_24534,N_24059);
xor UO_104 (O_104,N_24798,N_23754);
and UO_105 (O_105,N_24103,N_24130);
xor UO_106 (O_106,N_24446,N_24308);
or UO_107 (O_107,N_24082,N_23866);
xor UO_108 (O_108,N_24532,N_24557);
xnor UO_109 (O_109,N_24621,N_24086);
or UO_110 (O_110,N_24090,N_24092);
or UO_111 (O_111,N_24865,N_24312);
nor UO_112 (O_112,N_24517,N_24016);
or UO_113 (O_113,N_24981,N_23979);
nor UO_114 (O_114,N_23907,N_24829);
nand UO_115 (O_115,N_24579,N_24927);
or UO_116 (O_116,N_24820,N_23806);
or UO_117 (O_117,N_23938,N_24551);
or UO_118 (O_118,N_24648,N_23765);
and UO_119 (O_119,N_24298,N_24816);
nor UO_120 (O_120,N_24008,N_24376);
nand UO_121 (O_121,N_24093,N_23861);
or UO_122 (O_122,N_24830,N_24832);
xor UO_123 (O_123,N_24607,N_24664);
or UO_124 (O_124,N_24814,N_23869);
xnor UO_125 (O_125,N_24950,N_23816);
or UO_126 (O_126,N_24218,N_24533);
and UO_127 (O_127,N_24708,N_24695);
xnor UO_128 (O_128,N_24221,N_23997);
nand UO_129 (O_129,N_23894,N_24328);
nor UO_130 (O_130,N_23859,N_24608);
and UO_131 (O_131,N_23774,N_24911);
and UO_132 (O_132,N_24537,N_23952);
or UO_133 (O_133,N_24208,N_24509);
nand UO_134 (O_134,N_24321,N_24247);
nor UO_135 (O_135,N_23980,N_24801);
xor UO_136 (O_136,N_24455,N_24780);
xor UO_137 (O_137,N_24665,N_24003);
and UO_138 (O_138,N_24781,N_24451);
nand UO_139 (O_139,N_24857,N_24322);
or UO_140 (O_140,N_24464,N_24051);
xor UO_141 (O_141,N_24405,N_24027);
xor UO_142 (O_142,N_24220,N_24351);
nand UO_143 (O_143,N_24756,N_24932);
and UO_144 (O_144,N_24883,N_24284);
and UO_145 (O_145,N_24576,N_24493);
and UO_146 (O_146,N_24341,N_24057);
and UO_147 (O_147,N_24977,N_24768);
and UO_148 (O_148,N_24501,N_24997);
nand UO_149 (O_149,N_24229,N_24631);
or UO_150 (O_150,N_24880,N_24850);
nand UO_151 (O_151,N_24739,N_24162);
or UO_152 (O_152,N_23860,N_24141);
nand UO_153 (O_153,N_24416,N_23820);
nor UO_154 (O_154,N_24678,N_23752);
and UO_155 (O_155,N_24660,N_24224);
nand UO_156 (O_156,N_24054,N_23884);
xnor UO_157 (O_157,N_24006,N_24753);
xor UO_158 (O_158,N_24868,N_24187);
xnor UO_159 (O_159,N_24751,N_24004);
nor UO_160 (O_160,N_24529,N_24646);
and UO_161 (O_161,N_24406,N_24882);
or UO_162 (O_162,N_24073,N_24467);
nand UO_163 (O_163,N_24415,N_24861);
and UO_164 (O_164,N_23803,N_23769);
and UO_165 (O_165,N_24589,N_23779);
and UO_166 (O_166,N_24626,N_23879);
nor UO_167 (O_167,N_24921,N_24720);
nor UO_168 (O_168,N_24178,N_24367);
or UO_169 (O_169,N_24474,N_24758);
nand UO_170 (O_170,N_24817,N_23768);
nand UO_171 (O_171,N_24370,N_24049);
xor UO_172 (O_172,N_23964,N_23924);
nand UO_173 (O_173,N_24494,N_24507);
or UO_174 (O_174,N_24404,N_24855);
xor UO_175 (O_175,N_24261,N_24099);
nand UO_176 (O_176,N_24276,N_24571);
and UO_177 (O_177,N_24531,N_24641);
or UO_178 (O_178,N_24561,N_24615);
and UO_179 (O_179,N_24124,N_24114);
xor UO_180 (O_180,N_24998,N_24612);
or UO_181 (O_181,N_24856,N_24238);
xnor UO_182 (O_182,N_24267,N_24199);
nor UO_183 (O_183,N_24800,N_24588);
nor UO_184 (O_184,N_24598,N_23972);
nand UO_185 (O_185,N_23914,N_24433);
nand UO_186 (O_186,N_24179,N_24030);
nand UO_187 (O_187,N_24941,N_24223);
nor UO_188 (O_188,N_24435,N_24346);
or UO_189 (O_189,N_24991,N_23794);
xnor UO_190 (O_190,N_23909,N_24444);
nand UO_191 (O_191,N_24840,N_24259);
nor UO_192 (O_192,N_24755,N_23985);
or UO_193 (O_193,N_24245,N_24913);
and UO_194 (O_194,N_24210,N_23984);
nand UO_195 (O_195,N_24154,N_24682);
and UO_196 (O_196,N_24654,N_24696);
nor UO_197 (O_197,N_23941,N_24275);
nand UO_198 (O_198,N_24879,N_23958);
xor UO_199 (O_199,N_24083,N_24852);
and UO_200 (O_200,N_24380,N_24975);
xor UO_201 (O_201,N_24523,N_24990);
xnor UO_202 (O_202,N_24388,N_24905);
nand UO_203 (O_203,N_24914,N_24134);
or UO_204 (O_204,N_23760,N_24399);
nand UO_205 (O_205,N_24918,N_24481);
and UO_206 (O_206,N_24478,N_24895);
or UO_207 (O_207,N_24982,N_24301);
or UO_208 (O_208,N_23871,N_23947);
and UO_209 (O_209,N_24637,N_24847);
xor UO_210 (O_210,N_24915,N_24101);
and UO_211 (O_211,N_24155,N_24294);
nor UO_212 (O_212,N_24604,N_23804);
nand UO_213 (O_213,N_23832,N_24354);
and UO_214 (O_214,N_24552,N_23782);
nor UO_215 (O_215,N_24573,N_24859);
or UO_216 (O_216,N_23996,N_24900);
nor UO_217 (O_217,N_24230,N_24425);
nor UO_218 (O_218,N_24995,N_23793);
and UO_219 (O_219,N_24569,N_23904);
nor UO_220 (O_220,N_24910,N_24372);
and UO_221 (O_221,N_23825,N_24318);
and UO_222 (O_222,N_24822,N_24452);
and UO_223 (O_223,N_24397,N_24017);
and UO_224 (O_224,N_24384,N_24793);
and UO_225 (O_225,N_24782,N_24236);
and UO_226 (O_226,N_23953,N_24863);
nor UO_227 (O_227,N_24215,N_23949);
nand UO_228 (O_228,N_24749,N_24575);
or UO_229 (O_229,N_24689,N_24787);
nor UO_230 (O_230,N_24462,N_24401);
xor UO_231 (O_231,N_23911,N_24465);
nand UO_232 (O_232,N_24656,N_24675);
nor UO_233 (O_233,N_23930,N_24839);
nor UO_234 (O_234,N_24348,N_24808);
and UO_235 (O_235,N_24311,N_24304);
or UO_236 (O_236,N_23927,N_23998);
or UO_237 (O_237,N_24336,N_23827);
xor UO_238 (O_238,N_23948,N_24319);
xnor UO_239 (O_239,N_24201,N_24527);
nor UO_240 (O_240,N_24343,N_24545);
nand UO_241 (O_241,N_24805,N_24723);
xor UO_242 (O_242,N_24771,N_24988);
nor UO_243 (O_243,N_24672,N_24145);
or UO_244 (O_244,N_23759,N_23791);
or UO_245 (O_245,N_24585,N_24273);
xor UO_246 (O_246,N_23943,N_24978);
and UO_247 (O_247,N_23870,N_24395);
and UO_248 (O_248,N_24151,N_24593);
nand UO_249 (O_249,N_24996,N_24338);
nor UO_250 (O_250,N_24126,N_24624);
nand UO_251 (O_251,N_24707,N_24955);
and UO_252 (O_252,N_24884,N_24106);
xnor UO_253 (O_253,N_24644,N_23857);
nor UO_254 (O_254,N_24680,N_24310);
or UO_255 (O_255,N_23918,N_24342);
nand UO_256 (O_256,N_24345,N_24390);
or UO_257 (O_257,N_23811,N_24186);
nor UO_258 (O_258,N_24933,N_24524);
or UO_259 (O_259,N_24379,N_24835);
and UO_260 (O_260,N_24649,N_24191);
or UO_261 (O_261,N_24556,N_23792);
nand UO_262 (O_262,N_24231,N_24119);
xnor UO_263 (O_263,N_24281,N_24564);
nor UO_264 (O_264,N_24712,N_24587);
and UO_265 (O_265,N_23995,N_24323);
xor UO_266 (O_266,N_24741,N_24757);
and UO_267 (O_267,N_23824,N_24502);
and UO_268 (O_268,N_24418,N_24340);
nor UO_269 (O_269,N_23812,N_24919);
or UO_270 (O_270,N_24299,N_24457);
and UO_271 (O_271,N_24357,N_24036);
xnor UO_272 (O_272,N_24436,N_24568);
and UO_273 (O_273,N_24136,N_23881);
and UO_274 (O_274,N_24917,N_24110);
nand UO_275 (O_275,N_24702,N_23981);
nand UO_276 (O_276,N_24725,N_24775);
xnor UO_277 (O_277,N_24227,N_23838);
and UO_278 (O_278,N_24735,N_23784);
nand UO_279 (O_279,N_24440,N_23976);
or UO_280 (O_280,N_24733,N_24591);
or UO_281 (O_281,N_24111,N_24080);
nand UO_282 (O_282,N_23935,N_23891);
or UO_283 (O_283,N_24833,N_23987);
or UO_284 (O_284,N_24640,N_24968);
and UO_285 (O_285,N_24572,N_24091);
xor UO_286 (O_286,N_24407,N_24067);
nor UO_287 (O_287,N_24109,N_24293);
xor UO_288 (O_288,N_24123,N_24838);
and UO_289 (O_289,N_24205,N_24113);
nor UO_290 (O_290,N_24889,N_24072);
xor UO_291 (O_291,N_24251,N_23992);
and UO_292 (O_292,N_24595,N_24783);
or UO_293 (O_293,N_23888,N_24441);
or UO_294 (O_294,N_24959,N_24736);
xor UO_295 (O_295,N_24266,N_24704);
xnor UO_296 (O_296,N_24062,N_23982);
nand UO_297 (O_297,N_24738,N_24032);
or UO_298 (O_298,N_24306,N_24525);
nand UO_299 (O_299,N_24870,N_24873);
xor UO_300 (O_300,N_24973,N_24948);
or UO_301 (O_301,N_23886,N_24375);
or UO_302 (O_302,N_24402,N_24892);
and UO_303 (O_303,N_23767,N_24505);
and UO_304 (O_304,N_24862,N_24597);
or UO_305 (O_305,N_24290,N_24690);
xnor UO_306 (O_306,N_24325,N_23932);
nand UO_307 (O_307,N_23991,N_24335);
and UO_308 (O_308,N_23837,N_23963);
nor UO_309 (O_309,N_23868,N_24254);
and UO_310 (O_310,N_23753,N_24596);
or UO_311 (O_311,N_24476,N_23756);
xnor UO_312 (O_312,N_24853,N_24986);
or UO_313 (O_313,N_24734,N_23856);
nor UO_314 (O_314,N_24740,N_23801);
and UO_315 (O_315,N_24065,N_24842);
or UO_316 (O_316,N_24547,N_24877);
or UO_317 (O_317,N_24458,N_24951);
nor UO_318 (O_318,N_24746,N_24104);
xnor UO_319 (O_319,N_24243,N_24548);
xor UO_320 (O_320,N_24282,N_24289);
xnor UO_321 (O_321,N_24207,N_24204);
xnor UO_322 (O_322,N_24887,N_24606);
nor UO_323 (O_323,N_24430,N_24769);
nor UO_324 (O_324,N_24128,N_24622);
nor UO_325 (O_325,N_23954,N_24737);
nor UO_326 (O_326,N_24369,N_24412);
nand UO_327 (O_327,N_24147,N_24674);
xnor UO_328 (O_328,N_24480,N_24477);
xor UO_329 (O_329,N_24392,N_24448);
and UO_330 (O_330,N_24098,N_24655);
nor UO_331 (O_331,N_24287,N_24985);
nand UO_332 (O_332,N_24292,N_24730);
nor UO_333 (O_333,N_24670,N_24270);
xor UO_334 (O_334,N_24694,N_24860);
or UO_335 (O_335,N_24965,N_23783);
nand UO_336 (O_336,N_24601,N_24940);
and UO_337 (O_337,N_24048,N_24632);
nand UO_338 (O_338,N_24876,N_24423);
and UO_339 (O_339,N_23848,N_24639);
nand UO_340 (O_340,N_24813,N_24761);
nor UO_341 (O_341,N_24156,N_24329);
or UO_342 (O_342,N_24167,N_24466);
nor UO_343 (O_343,N_23797,N_24025);
xor UO_344 (O_344,N_24012,N_24987);
nor UO_345 (O_345,N_24609,N_24992);
and UO_346 (O_346,N_23908,N_24410);
and UO_347 (O_347,N_24963,N_24958);
nor UO_348 (O_348,N_24779,N_24408);
or UO_349 (O_349,N_24945,N_23903);
nor UO_350 (O_350,N_24339,N_24184);
xnor UO_351 (O_351,N_24232,N_24020);
and UO_352 (O_352,N_24190,N_24071);
nor UO_353 (O_353,N_24239,N_24490);
nor UO_354 (O_354,N_23931,N_24976);
xnor UO_355 (O_355,N_24891,N_24872);
nand UO_356 (O_356,N_24094,N_24947);
nand UO_357 (O_357,N_24908,N_24928);
xnor UO_358 (O_358,N_24180,N_23818);
and UO_359 (O_359,N_23934,N_24821);
xnor UO_360 (O_360,N_24967,N_24888);
xnor UO_361 (O_361,N_24420,N_24834);
nor UO_362 (O_362,N_24952,N_24500);
xor UO_363 (O_363,N_23834,N_24089);
or UO_364 (O_364,N_24195,N_24373);
xor UO_365 (O_365,N_23965,N_24540);
nand UO_366 (O_366,N_24634,N_24192);
and UO_367 (O_367,N_24240,N_24954);
and UO_368 (O_368,N_23898,N_24010);
nand UO_369 (O_369,N_24745,N_24693);
nor UO_370 (O_370,N_23882,N_24361);
and UO_371 (O_371,N_24799,N_23899);
and UO_372 (O_372,N_24031,N_24443);
or UO_373 (O_373,N_24492,N_24881);
nand UO_374 (O_374,N_24498,N_24078);
and UO_375 (O_375,N_24149,N_24922);
nor UO_376 (O_376,N_24482,N_23750);
nand UO_377 (O_377,N_24776,N_24923);
or UO_378 (O_378,N_24600,N_24213);
or UO_379 (O_379,N_24303,N_23802);
or UO_380 (O_380,N_23808,N_24288);
nand UO_381 (O_381,N_24314,N_23905);
nand UO_382 (O_382,N_24047,N_24851);
nand UO_383 (O_383,N_23770,N_24906);
nor UO_384 (O_384,N_24255,N_23990);
nor UO_385 (O_385,N_24324,N_24539);
and UO_386 (O_386,N_24185,N_24514);
and UO_387 (O_387,N_23786,N_24553);
or UO_388 (O_388,N_23817,N_24356);
xor UO_389 (O_389,N_23969,N_23922);
xnor UO_390 (O_390,N_24454,N_24422);
nand UO_391 (O_391,N_24748,N_24785);
nand UO_392 (O_392,N_23875,N_24513);
or UO_393 (O_393,N_23772,N_23863);
or UO_394 (O_394,N_24957,N_24560);
nor UO_395 (O_395,N_24456,N_23841);
nor UO_396 (O_396,N_24045,N_24864);
or UO_397 (O_397,N_24052,N_24060);
nand UO_398 (O_398,N_24826,N_23878);
xnor UO_399 (O_399,N_24935,N_24774);
nand UO_400 (O_400,N_24291,N_24999);
and UO_401 (O_401,N_23936,N_23873);
and UO_402 (O_402,N_24866,N_24506);
nand UO_403 (O_403,N_24302,N_24943);
nand UO_404 (O_404,N_24331,N_23851);
and UO_405 (O_405,N_24211,N_24076);
nor UO_406 (O_406,N_24836,N_24206);
nor UO_407 (O_407,N_24815,N_24511);
and UO_408 (O_408,N_24497,N_24026);
xor UO_409 (O_409,N_23885,N_24337);
xor UO_410 (O_410,N_24305,N_24926);
or UO_411 (O_411,N_24770,N_24453);
and UO_412 (O_412,N_24979,N_24972);
nor UO_413 (O_413,N_24100,N_24096);
nand UO_414 (O_414,N_24280,N_24619);
nor UO_415 (O_415,N_24152,N_24142);
xor UO_416 (O_416,N_24353,N_24669);
or UO_417 (O_417,N_24144,N_23815);
nor UO_418 (O_418,N_23895,N_24143);
and UO_419 (O_419,N_24938,N_24869);
or UO_420 (O_420,N_24125,N_24264);
xor UO_421 (O_421,N_24651,N_24726);
and UO_422 (O_422,N_24686,N_23766);
nand UO_423 (O_423,N_23880,N_24828);
nand UO_424 (O_424,N_24819,N_24056);
and UO_425 (O_425,N_24790,N_24645);
or UO_426 (O_426,N_24643,N_24673);
or UO_427 (O_427,N_24473,N_24956);
and UO_428 (O_428,N_24874,N_23993);
and UO_429 (O_429,N_24647,N_24666);
nor UO_430 (O_430,N_24538,N_24760);
xor UO_431 (O_431,N_24391,N_24792);
xor UO_432 (O_432,N_23944,N_24685);
and UO_433 (O_433,N_23836,N_24426);
and UO_434 (O_434,N_24555,N_24942);
nand UO_435 (O_435,N_23973,N_24212);
and UO_436 (O_436,N_23923,N_24252);
or UO_437 (O_437,N_24069,N_23897);
nand UO_438 (O_438,N_24743,N_24962);
xor UO_439 (O_439,N_24974,N_24018);
nand UO_440 (O_440,N_24661,N_23877);
nor UO_441 (O_441,N_24225,N_24802);
xnor UO_442 (O_442,N_24562,N_24944);
nand UO_443 (O_443,N_23819,N_24489);
or UO_444 (O_444,N_24846,N_24475);
nand UO_445 (O_445,N_24447,N_24616);
nand UO_446 (O_446,N_24930,N_23831);
nor UO_447 (O_447,N_24161,N_23761);
nor UO_448 (O_448,N_24000,N_24714);
and UO_449 (O_449,N_24542,N_24677);
xor UO_450 (O_450,N_24628,N_23777);
xor UO_451 (O_451,N_24409,N_24387);
nand UO_452 (O_452,N_23787,N_23798);
and UO_453 (O_453,N_23968,N_24159);
and UO_454 (O_454,N_24789,N_23842);
and UO_455 (O_455,N_24495,N_24710);
nand UO_456 (O_456,N_24368,N_24683);
xnor UO_457 (O_457,N_24382,N_24170);
xor UO_458 (O_458,N_24788,N_23883);
or UO_459 (O_459,N_24574,N_24719);
xnor UO_460 (O_460,N_24181,N_24657);
or UO_461 (O_461,N_24414,N_24767);
nor UO_462 (O_462,N_23966,N_24034);
nor UO_463 (O_463,N_24286,N_24445);
nor UO_464 (O_464,N_24460,N_24920);
or UO_465 (O_465,N_23896,N_23807);
nor UO_466 (O_466,N_24818,N_24085);
and UO_467 (O_467,N_24403,N_24692);
or UO_468 (O_468,N_24347,N_24841);
or UO_469 (O_469,N_24313,N_24417);
nor UO_470 (O_470,N_24279,N_24784);
and UO_471 (O_471,N_24198,N_24487);
nor UO_472 (O_472,N_24584,N_23950);
nand UO_473 (O_473,N_24035,N_24256);
nand UO_474 (O_474,N_24250,N_24317);
or UO_475 (O_475,N_24150,N_24118);
and UO_476 (O_476,N_23876,N_24271);
and UO_477 (O_477,N_24171,N_24400);
xor UO_478 (O_478,N_24437,N_24807);
nor UO_479 (O_479,N_24728,N_23961);
or UO_480 (O_480,N_24486,N_24427);
and UO_481 (O_481,N_24189,N_23942);
nor UO_482 (O_482,N_23960,N_24582);
nand UO_483 (O_483,N_24411,N_24158);
nor UO_484 (O_484,N_24488,N_24535);
nor UO_485 (O_485,N_24088,N_23999);
nand UO_486 (O_486,N_23799,N_24352);
or UO_487 (O_487,N_23821,N_23833);
xnor UO_488 (O_488,N_24837,N_24570);
nand UO_489 (O_489,N_24164,N_24176);
nor UO_490 (O_490,N_24217,N_24617);
or UO_491 (O_491,N_24362,N_24848);
nand UO_492 (O_492,N_24009,N_24762);
nor UO_493 (O_493,N_24937,N_24925);
and UO_494 (O_494,N_24122,N_24804);
nor UO_495 (O_495,N_24667,N_23822);
xnor UO_496 (O_496,N_24050,N_23835);
nand UO_497 (O_497,N_24269,N_24586);
and UO_498 (O_498,N_24383,N_24327);
and UO_499 (O_499,N_24658,N_24980);
and UO_500 (O_500,N_23951,N_24994);
nand UO_501 (O_501,N_24602,N_24222);
nor UO_502 (O_502,N_24268,N_24684);
nand UO_503 (O_503,N_24679,N_24366);
nor UO_504 (O_504,N_23790,N_24244);
or UO_505 (O_505,N_23778,N_24061);
nor UO_506 (O_506,N_24583,N_24796);
nand UO_507 (O_507,N_24097,N_24717);
and UO_508 (O_508,N_23928,N_24024);
nor UO_509 (O_509,N_23775,N_24491);
or UO_510 (O_510,N_24172,N_24698);
nand UO_511 (O_511,N_24175,N_24438);
nand UO_512 (O_512,N_24262,N_23826);
nand UO_513 (O_513,N_24285,N_23780);
nor UO_514 (O_514,N_24248,N_24214);
and UO_515 (O_515,N_23989,N_24272);
xor UO_516 (O_516,N_23925,N_23795);
nor UO_517 (O_517,N_24283,N_24759);
xnor UO_518 (O_518,N_24068,N_24139);
xnor UO_519 (O_519,N_23865,N_24105);
nand UO_520 (O_520,N_23893,N_24138);
or UO_521 (O_521,N_24522,N_24700);
or UO_522 (O_522,N_24449,N_24731);
nand UO_523 (O_523,N_24233,N_24063);
nand UO_524 (O_524,N_23939,N_24360);
and UO_525 (O_525,N_24182,N_23957);
nand UO_526 (O_526,N_24013,N_24007);
nand UO_527 (O_527,N_24483,N_23867);
nand UO_528 (O_528,N_23902,N_24949);
or UO_529 (O_529,N_24163,N_24108);
nand UO_530 (O_530,N_24075,N_24871);
or UO_531 (O_531,N_24398,N_24127);
and UO_532 (O_532,N_24112,N_24153);
and UO_533 (O_533,N_24116,N_23844);
nand UO_534 (O_534,N_24971,N_24146);
or UO_535 (O_535,N_24929,N_24699);
nor UO_536 (O_536,N_24970,N_24365);
nand UO_537 (O_537,N_24040,N_23887);
nand UO_538 (O_538,N_24058,N_23889);
or UO_539 (O_539,N_24468,N_24203);
nor UO_540 (O_540,N_24526,N_24043);
or UO_541 (O_541,N_23874,N_24334);
and UO_542 (O_542,N_24496,N_23751);
nand UO_543 (O_543,N_24396,N_24681);
nor UO_544 (O_544,N_24823,N_24469);
nand UO_545 (O_545,N_24095,N_23853);
or UO_546 (O_546,N_24844,N_24508);
nand UO_547 (O_547,N_23945,N_24620);
nor UO_548 (O_548,N_24924,N_24652);
nor UO_549 (O_549,N_24107,N_24183);
nor UO_550 (O_550,N_24249,N_24038);
xnor UO_551 (O_551,N_24055,N_23913);
and UO_552 (O_552,N_23967,N_24359);
nor UO_553 (O_553,N_24550,N_23959);
or UO_554 (O_554,N_24903,N_24196);
nor UO_555 (O_555,N_24041,N_24898);
and UO_556 (O_556,N_23920,N_24168);
nand UO_557 (O_557,N_24721,N_24363);
nor UO_558 (O_558,N_24536,N_24389);
nand UO_559 (O_559,N_24983,N_24326);
and UO_560 (O_560,N_24042,N_24246);
xor UO_561 (O_561,N_24121,N_23852);
and UO_562 (O_562,N_24845,N_24461);
and UO_563 (O_563,N_24729,N_23810);
and UO_564 (O_564,N_24742,N_24265);
nand UO_565 (O_565,N_24381,N_24791);
nor UO_566 (O_566,N_24241,N_24015);
nand UO_567 (O_567,N_24135,N_24544);
or UO_568 (O_568,N_24630,N_24812);
or UO_569 (O_569,N_24961,N_24257);
or UO_570 (O_570,N_24578,N_24936);
nor UO_571 (O_571,N_24117,N_24029);
and UO_572 (O_572,N_24157,N_24629);
nand UO_573 (O_573,N_24614,N_24120);
nor UO_574 (O_574,N_23970,N_24894);
xor UO_575 (O_575,N_24428,N_24697);
or UO_576 (O_576,N_24969,N_24046);
and UO_577 (O_577,N_24014,N_24662);
or UO_578 (O_578,N_23847,N_23823);
xor UO_579 (O_579,N_24603,N_24563);
xnor UO_580 (O_580,N_24022,N_24912);
and UO_581 (O_581,N_23764,N_24530);
or UO_582 (O_582,N_24613,N_24077);
nand UO_583 (O_583,N_24795,N_23845);
xnor UO_584 (O_584,N_24727,N_23813);
nor UO_585 (O_585,N_24188,N_24605);
xnor UO_586 (O_586,N_24431,N_24966);
and UO_587 (O_587,N_23929,N_24173);
nand UO_588 (O_588,N_24705,N_24237);
nor UO_589 (O_589,N_24594,N_24824);
nor UO_590 (O_590,N_24066,N_23800);
xor UO_591 (O_591,N_24516,N_23830);
nand UO_592 (O_592,N_24084,N_23843);
xnor UO_593 (O_593,N_24316,N_23771);
or UO_594 (O_594,N_24939,N_24504);
nor UO_595 (O_595,N_24332,N_24902);
nor UO_596 (O_596,N_23850,N_24627);
or UO_597 (O_597,N_24131,N_24993);
nand UO_598 (O_598,N_23840,N_24350);
nand UO_599 (O_599,N_24174,N_24825);
xnor UO_600 (O_600,N_24565,N_24002);
or UO_601 (O_601,N_23890,N_24515);
nand UO_602 (O_602,N_24811,N_24315);
and UO_603 (O_603,N_24541,N_24916);
or UO_604 (O_604,N_24081,N_24786);
and UO_605 (O_605,N_24827,N_24140);
and UO_606 (O_606,N_24019,N_24885);
nand UO_607 (O_607,N_24592,N_24688);
or UO_608 (O_608,N_24005,N_23917);
nor UO_609 (O_609,N_23849,N_23763);
xor UO_610 (O_610,N_24499,N_23937);
nor UO_611 (O_611,N_24377,N_24528);
nand UO_612 (O_612,N_24794,N_24219);
and UO_613 (O_613,N_24610,N_24209);
xnor UO_614 (O_614,N_24023,N_24148);
nor UO_615 (O_615,N_23933,N_24300);
or UO_616 (O_616,N_24421,N_24260);
nand UO_617 (O_617,N_24394,N_24296);
nand UO_618 (O_618,N_23788,N_23916);
nand UO_619 (O_619,N_23757,N_24011);
xor UO_620 (O_620,N_23805,N_24450);
xnor UO_621 (O_621,N_24307,N_24166);
nand UO_622 (O_622,N_24253,N_23789);
nor UO_623 (O_623,N_24471,N_24543);
nor UO_624 (O_624,N_24715,N_23829);
and UO_625 (O_625,N_24587,N_24127);
or UO_626 (O_626,N_24587,N_24364);
and UO_627 (O_627,N_24554,N_24906);
xnor UO_628 (O_628,N_24619,N_24628);
xor UO_629 (O_629,N_24791,N_24769);
nor UO_630 (O_630,N_24875,N_23765);
and UO_631 (O_631,N_24808,N_24999);
and UO_632 (O_632,N_24422,N_24802);
xnor UO_633 (O_633,N_23960,N_24498);
and UO_634 (O_634,N_24636,N_24409);
xnor UO_635 (O_635,N_24758,N_23803);
nor UO_636 (O_636,N_24918,N_24488);
and UO_637 (O_637,N_24641,N_24675);
and UO_638 (O_638,N_24143,N_23824);
and UO_639 (O_639,N_24520,N_23915);
xnor UO_640 (O_640,N_24698,N_24254);
xnor UO_641 (O_641,N_23976,N_23775);
or UO_642 (O_642,N_23804,N_24815);
or UO_643 (O_643,N_24518,N_24220);
and UO_644 (O_644,N_24776,N_23859);
xor UO_645 (O_645,N_24067,N_24885);
nand UO_646 (O_646,N_24208,N_24411);
xor UO_647 (O_647,N_24694,N_23890);
or UO_648 (O_648,N_23845,N_23860);
xnor UO_649 (O_649,N_24750,N_24030);
nor UO_650 (O_650,N_24068,N_24533);
xnor UO_651 (O_651,N_23902,N_23917);
and UO_652 (O_652,N_24962,N_24364);
nor UO_653 (O_653,N_24312,N_24793);
nor UO_654 (O_654,N_24011,N_23789);
nand UO_655 (O_655,N_23999,N_24761);
and UO_656 (O_656,N_24743,N_24690);
or UO_657 (O_657,N_24580,N_23916);
and UO_658 (O_658,N_23984,N_24313);
nand UO_659 (O_659,N_23822,N_24179);
and UO_660 (O_660,N_24304,N_24687);
or UO_661 (O_661,N_24537,N_24434);
or UO_662 (O_662,N_24913,N_24520);
nor UO_663 (O_663,N_24892,N_24182);
and UO_664 (O_664,N_24056,N_24429);
nand UO_665 (O_665,N_24882,N_23878);
nor UO_666 (O_666,N_24540,N_24821);
and UO_667 (O_667,N_24170,N_23871);
nor UO_668 (O_668,N_23914,N_24659);
and UO_669 (O_669,N_24899,N_24314);
nand UO_670 (O_670,N_24752,N_24201);
nor UO_671 (O_671,N_24031,N_24268);
nor UO_672 (O_672,N_24147,N_23938);
nor UO_673 (O_673,N_24212,N_23902);
and UO_674 (O_674,N_24906,N_24203);
xnor UO_675 (O_675,N_24939,N_24075);
xnor UO_676 (O_676,N_24261,N_23919);
or UO_677 (O_677,N_24159,N_24810);
nor UO_678 (O_678,N_23998,N_24630);
or UO_679 (O_679,N_24926,N_23779);
xnor UO_680 (O_680,N_23954,N_24663);
nor UO_681 (O_681,N_23778,N_24530);
and UO_682 (O_682,N_24569,N_24696);
nor UO_683 (O_683,N_24304,N_23974);
nand UO_684 (O_684,N_24039,N_24914);
and UO_685 (O_685,N_23937,N_24821);
or UO_686 (O_686,N_24724,N_24149);
or UO_687 (O_687,N_23970,N_24087);
or UO_688 (O_688,N_24732,N_24753);
and UO_689 (O_689,N_24728,N_24341);
and UO_690 (O_690,N_24319,N_24641);
xor UO_691 (O_691,N_24913,N_24648);
or UO_692 (O_692,N_23946,N_24440);
or UO_693 (O_693,N_24899,N_24356);
nor UO_694 (O_694,N_24159,N_23831);
and UO_695 (O_695,N_24466,N_24937);
nand UO_696 (O_696,N_24984,N_24554);
xnor UO_697 (O_697,N_24721,N_24167);
nor UO_698 (O_698,N_24570,N_24892);
and UO_699 (O_699,N_24128,N_23829);
nand UO_700 (O_700,N_23945,N_24088);
or UO_701 (O_701,N_23866,N_24863);
and UO_702 (O_702,N_24964,N_24240);
and UO_703 (O_703,N_24352,N_23797);
and UO_704 (O_704,N_24742,N_24881);
nand UO_705 (O_705,N_24838,N_24326);
or UO_706 (O_706,N_24774,N_24745);
nor UO_707 (O_707,N_24662,N_24191);
nor UO_708 (O_708,N_24926,N_23969);
and UO_709 (O_709,N_24905,N_24646);
or UO_710 (O_710,N_24985,N_24089);
and UO_711 (O_711,N_24919,N_24557);
nand UO_712 (O_712,N_24542,N_23859);
nor UO_713 (O_713,N_24976,N_24458);
or UO_714 (O_714,N_24404,N_24379);
nand UO_715 (O_715,N_24342,N_24053);
xor UO_716 (O_716,N_23791,N_24000);
and UO_717 (O_717,N_24194,N_24820);
or UO_718 (O_718,N_23936,N_24453);
xnor UO_719 (O_719,N_24662,N_24551);
nand UO_720 (O_720,N_24502,N_23894);
nand UO_721 (O_721,N_23777,N_24839);
xnor UO_722 (O_722,N_24124,N_23960);
nor UO_723 (O_723,N_23779,N_24655);
xnor UO_724 (O_724,N_24105,N_24298);
or UO_725 (O_725,N_24589,N_24825);
nand UO_726 (O_726,N_23817,N_24416);
or UO_727 (O_727,N_23812,N_24904);
nand UO_728 (O_728,N_23948,N_24757);
nor UO_729 (O_729,N_24235,N_24047);
and UO_730 (O_730,N_24048,N_24151);
or UO_731 (O_731,N_24789,N_23768);
xor UO_732 (O_732,N_24234,N_23964);
and UO_733 (O_733,N_23887,N_24253);
and UO_734 (O_734,N_24729,N_24188);
nor UO_735 (O_735,N_23833,N_24486);
nor UO_736 (O_736,N_23974,N_24203);
xor UO_737 (O_737,N_24362,N_24569);
nor UO_738 (O_738,N_24881,N_23870);
nor UO_739 (O_739,N_24943,N_24810);
xnor UO_740 (O_740,N_24972,N_23777);
and UO_741 (O_741,N_24176,N_24689);
or UO_742 (O_742,N_24284,N_23952);
xor UO_743 (O_743,N_23818,N_24395);
or UO_744 (O_744,N_23776,N_23867);
and UO_745 (O_745,N_24299,N_24855);
or UO_746 (O_746,N_24639,N_24012);
or UO_747 (O_747,N_24191,N_24495);
and UO_748 (O_748,N_24000,N_23899);
xnor UO_749 (O_749,N_24780,N_24958);
or UO_750 (O_750,N_24697,N_24199);
nor UO_751 (O_751,N_24046,N_24482);
and UO_752 (O_752,N_23896,N_24723);
xor UO_753 (O_753,N_24481,N_24888);
nor UO_754 (O_754,N_24788,N_23797);
nand UO_755 (O_755,N_24200,N_24508);
nor UO_756 (O_756,N_24637,N_24083);
or UO_757 (O_757,N_24720,N_24911);
and UO_758 (O_758,N_24332,N_24863);
and UO_759 (O_759,N_24109,N_24677);
and UO_760 (O_760,N_23946,N_24077);
xor UO_761 (O_761,N_24386,N_24174);
nand UO_762 (O_762,N_24271,N_24029);
and UO_763 (O_763,N_24293,N_24027);
nor UO_764 (O_764,N_24180,N_24522);
and UO_765 (O_765,N_24484,N_23994);
and UO_766 (O_766,N_24400,N_24920);
nand UO_767 (O_767,N_24885,N_24823);
xor UO_768 (O_768,N_24265,N_24481);
xnor UO_769 (O_769,N_24207,N_24824);
xnor UO_770 (O_770,N_23845,N_24541);
nor UO_771 (O_771,N_24986,N_24482);
or UO_772 (O_772,N_24997,N_24000);
and UO_773 (O_773,N_24307,N_24122);
nor UO_774 (O_774,N_24408,N_23801);
xnor UO_775 (O_775,N_24364,N_24503);
or UO_776 (O_776,N_24857,N_24821);
xor UO_777 (O_777,N_24524,N_23830);
or UO_778 (O_778,N_24424,N_24758);
nand UO_779 (O_779,N_24696,N_24662);
or UO_780 (O_780,N_24617,N_23856);
and UO_781 (O_781,N_23978,N_24029);
and UO_782 (O_782,N_23769,N_24206);
and UO_783 (O_783,N_24129,N_24160);
nand UO_784 (O_784,N_24956,N_24194);
xnor UO_785 (O_785,N_24082,N_24169);
xnor UO_786 (O_786,N_24021,N_23970);
xnor UO_787 (O_787,N_24274,N_24628);
and UO_788 (O_788,N_24777,N_23784);
nor UO_789 (O_789,N_24572,N_23957);
nor UO_790 (O_790,N_24193,N_24686);
nor UO_791 (O_791,N_24566,N_24863);
xnor UO_792 (O_792,N_24382,N_23921);
nand UO_793 (O_793,N_24637,N_24979);
and UO_794 (O_794,N_24227,N_24603);
nand UO_795 (O_795,N_24391,N_24180);
and UO_796 (O_796,N_24274,N_24042);
nor UO_797 (O_797,N_24343,N_24690);
nand UO_798 (O_798,N_24714,N_24224);
nand UO_799 (O_799,N_24136,N_24810);
nand UO_800 (O_800,N_24286,N_23839);
xor UO_801 (O_801,N_23843,N_23877);
xnor UO_802 (O_802,N_24804,N_24406);
xor UO_803 (O_803,N_24510,N_24895);
nor UO_804 (O_804,N_24938,N_24137);
nor UO_805 (O_805,N_24194,N_24969);
xnor UO_806 (O_806,N_23833,N_24716);
or UO_807 (O_807,N_24118,N_24642);
or UO_808 (O_808,N_24192,N_24594);
nand UO_809 (O_809,N_24483,N_24924);
nand UO_810 (O_810,N_24821,N_24758);
and UO_811 (O_811,N_24308,N_23996);
or UO_812 (O_812,N_24269,N_24609);
nor UO_813 (O_813,N_24302,N_24140);
nor UO_814 (O_814,N_23862,N_24556);
nor UO_815 (O_815,N_24782,N_24337);
nor UO_816 (O_816,N_24020,N_24915);
xor UO_817 (O_817,N_24046,N_23847);
and UO_818 (O_818,N_24830,N_24596);
and UO_819 (O_819,N_24127,N_23874);
nor UO_820 (O_820,N_23841,N_24747);
or UO_821 (O_821,N_24142,N_24293);
and UO_822 (O_822,N_24931,N_24617);
xor UO_823 (O_823,N_24908,N_24494);
or UO_824 (O_824,N_24839,N_24908);
nor UO_825 (O_825,N_23823,N_24584);
and UO_826 (O_826,N_24164,N_24505);
nor UO_827 (O_827,N_24865,N_24356);
or UO_828 (O_828,N_24641,N_24630);
or UO_829 (O_829,N_24016,N_24786);
and UO_830 (O_830,N_24400,N_24391);
nor UO_831 (O_831,N_24016,N_24736);
nand UO_832 (O_832,N_24146,N_24539);
and UO_833 (O_833,N_23823,N_23770);
or UO_834 (O_834,N_24490,N_24492);
or UO_835 (O_835,N_24216,N_24965);
nor UO_836 (O_836,N_24795,N_24884);
nand UO_837 (O_837,N_24439,N_23798);
and UO_838 (O_838,N_24461,N_24665);
xnor UO_839 (O_839,N_24029,N_24487);
or UO_840 (O_840,N_24240,N_23806);
xnor UO_841 (O_841,N_24070,N_24021);
or UO_842 (O_842,N_24992,N_24897);
xnor UO_843 (O_843,N_24692,N_24826);
xor UO_844 (O_844,N_24962,N_23764);
nor UO_845 (O_845,N_24039,N_24193);
or UO_846 (O_846,N_23793,N_23810);
or UO_847 (O_847,N_24440,N_24902);
and UO_848 (O_848,N_23958,N_24148);
and UO_849 (O_849,N_24387,N_24561);
nor UO_850 (O_850,N_24213,N_24811);
nand UO_851 (O_851,N_24570,N_24902);
nor UO_852 (O_852,N_24888,N_23898);
nand UO_853 (O_853,N_24492,N_24454);
and UO_854 (O_854,N_24039,N_23948);
nand UO_855 (O_855,N_24176,N_23815);
and UO_856 (O_856,N_24829,N_24580);
or UO_857 (O_857,N_24880,N_24616);
xnor UO_858 (O_858,N_24619,N_24350);
xor UO_859 (O_859,N_24017,N_24118);
or UO_860 (O_860,N_24590,N_24583);
nand UO_861 (O_861,N_24436,N_23904);
nand UO_862 (O_862,N_24808,N_24927);
xor UO_863 (O_863,N_24685,N_23969);
nand UO_864 (O_864,N_24297,N_24705);
nand UO_865 (O_865,N_24773,N_24955);
nand UO_866 (O_866,N_24937,N_24762);
xor UO_867 (O_867,N_24197,N_24132);
or UO_868 (O_868,N_23765,N_24247);
and UO_869 (O_869,N_24147,N_24727);
and UO_870 (O_870,N_23999,N_24897);
nor UO_871 (O_871,N_23977,N_24920);
and UO_872 (O_872,N_24022,N_24466);
nor UO_873 (O_873,N_24501,N_24744);
nand UO_874 (O_874,N_23905,N_24528);
xnor UO_875 (O_875,N_24420,N_23839);
nor UO_876 (O_876,N_23812,N_24912);
nor UO_877 (O_877,N_24178,N_23846);
nor UO_878 (O_878,N_24655,N_23958);
or UO_879 (O_879,N_24600,N_24318);
or UO_880 (O_880,N_24318,N_24782);
xor UO_881 (O_881,N_24799,N_23984);
or UO_882 (O_882,N_24577,N_24311);
or UO_883 (O_883,N_23974,N_24215);
and UO_884 (O_884,N_24221,N_24865);
or UO_885 (O_885,N_23853,N_24493);
or UO_886 (O_886,N_24866,N_24819);
xor UO_887 (O_887,N_24031,N_24762);
nor UO_888 (O_888,N_24781,N_24947);
and UO_889 (O_889,N_24772,N_24830);
and UO_890 (O_890,N_23777,N_23913);
nor UO_891 (O_891,N_24003,N_23840);
and UO_892 (O_892,N_24044,N_24987);
and UO_893 (O_893,N_24529,N_24946);
nand UO_894 (O_894,N_24275,N_24994);
xor UO_895 (O_895,N_24087,N_23777);
nor UO_896 (O_896,N_23785,N_24259);
and UO_897 (O_897,N_24066,N_24962);
nor UO_898 (O_898,N_23982,N_23993);
and UO_899 (O_899,N_23943,N_24622);
or UO_900 (O_900,N_24364,N_24090);
or UO_901 (O_901,N_24706,N_24748);
nor UO_902 (O_902,N_24186,N_24051);
xnor UO_903 (O_903,N_24795,N_24985);
xor UO_904 (O_904,N_24353,N_24792);
and UO_905 (O_905,N_24697,N_24279);
nor UO_906 (O_906,N_24365,N_24072);
nor UO_907 (O_907,N_24655,N_24814);
and UO_908 (O_908,N_24385,N_24228);
and UO_909 (O_909,N_24282,N_24516);
xor UO_910 (O_910,N_23816,N_24373);
xor UO_911 (O_911,N_24639,N_24662);
xnor UO_912 (O_912,N_24211,N_24351);
or UO_913 (O_913,N_24957,N_24859);
and UO_914 (O_914,N_24837,N_24306);
xnor UO_915 (O_915,N_24113,N_24226);
nand UO_916 (O_916,N_24554,N_24830);
or UO_917 (O_917,N_24910,N_23898);
nor UO_918 (O_918,N_24003,N_24449);
nor UO_919 (O_919,N_24807,N_24928);
xnor UO_920 (O_920,N_24059,N_24855);
and UO_921 (O_921,N_24469,N_24968);
nand UO_922 (O_922,N_23808,N_24468);
xnor UO_923 (O_923,N_23899,N_24374);
and UO_924 (O_924,N_24732,N_24536);
nor UO_925 (O_925,N_24946,N_24807);
nor UO_926 (O_926,N_24357,N_24620);
nor UO_927 (O_927,N_23883,N_23786);
and UO_928 (O_928,N_24213,N_24791);
or UO_929 (O_929,N_24625,N_23969);
nor UO_930 (O_930,N_24804,N_24067);
xor UO_931 (O_931,N_24678,N_24716);
nor UO_932 (O_932,N_24111,N_24082);
xor UO_933 (O_933,N_24372,N_24698);
or UO_934 (O_934,N_24756,N_23969);
or UO_935 (O_935,N_24937,N_24437);
nand UO_936 (O_936,N_24458,N_24521);
xor UO_937 (O_937,N_24477,N_24522);
and UO_938 (O_938,N_24156,N_24833);
xnor UO_939 (O_939,N_24295,N_23798);
or UO_940 (O_940,N_24943,N_24759);
and UO_941 (O_941,N_24612,N_24288);
xor UO_942 (O_942,N_23886,N_24028);
and UO_943 (O_943,N_24917,N_24844);
nand UO_944 (O_944,N_24099,N_24341);
xnor UO_945 (O_945,N_24112,N_24465);
nand UO_946 (O_946,N_24222,N_24142);
xnor UO_947 (O_947,N_24131,N_24459);
and UO_948 (O_948,N_24990,N_23752);
and UO_949 (O_949,N_24902,N_24601);
or UO_950 (O_950,N_24554,N_24926);
or UO_951 (O_951,N_24038,N_24791);
nand UO_952 (O_952,N_23955,N_24182);
nand UO_953 (O_953,N_23764,N_24051);
xnor UO_954 (O_954,N_24544,N_24034);
nor UO_955 (O_955,N_24430,N_24389);
nand UO_956 (O_956,N_24385,N_23768);
nor UO_957 (O_957,N_24078,N_24991);
nor UO_958 (O_958,N_24164,N_24918);
or UO_959 (O_959,N_24310,N_24925);
nor UO_960 (O_960,N_24811,N_24776);
nor UO_961 (O_961,N_24513,N_24936);
and UO_962 (O_962,N_23800,N_23811);
or UO_963 (O_963,N_24791,N_24183);
nand UO_964 (O_964,N_23986,N_24873);
or UO_965 (O_965,N_24829,N_24212);
xnor UO_966 (O_966,N_24370,N_24829);
xnor UO_967 (O_967,N_24819,N_24892);
xor UO_968 (O_968,N_24876,N_24024);
nand UO_969 (O_969,N_23763,N_24719);
nand UO_970 (O_970,N_24065,N_24589);
xor UO_971 (O_971,N_23921,N_23867);
or UO_972 (O_972,N_23948,N_24802);
nand UO_973 (O_973,N_23969,N_23883);
xor UO_974 (O_974,N_24068,N_23960);
nor UO_975 (O_975,N_24911,N_24688);
and UO_976 (O_976,N_24673,N_24116);
xnor UO_977 (O_977,N_24447,N_23952);
nand UO_978 (O_978,N_23876,N_24932);
and UO_979 (O_979,N_24036,N_24779);
and UO_980 (O_980,N_24847,N_24194);
and UO_981 (O_981,N_24945,N_24087);
nand UO_982 (O_982,N_24142,N_24143);
and UO_983 (O_983,N_24294,N_24224);
nor UO_984 (O_984,N_24075,N_24511);
or UO_985 (O_985,N_23791,N_24516);
nand UO_986 (O_986,N_24996,N_24692);
and UO_987 (O_987,N_24598,N_24367);
and UO_988 (O_988,N_24401,N_23751);
xor UO_989 (O_989,N_24315,N_24148);
nand UO_990 (O_990,N_24786,N_23898);
xor UO_991 (O_991,N_24955,N_23808);
and UO_992 (O_992,N_24448,N_24880);
or UO_993 (O_993,N_24002,N_24966);
nand UO_994 (O_994,N_24041,N_24845);
nand UO_995 (O_995,N_24873,N_24372);
xor UO_996 (O_996,N_24227,N_23869);
nor UO_997 (O_997,N_23834,N_24423);
or UO_998 (O_998,N_24733,N_24353);
xor UO_999 (O_999,N_24852,N_24255);
or UO_1000 (O_1000,N_24399,N_24040);
and UO_1001 (O_1001,N_24451,N_24073);
and UO_1002 (O_1002,N_24583,N_23909);
or UO_1003 (O_1003,N_24932,N_24296);
xor UO_1004 (O_1004,N_24704,N_24297);
nor UO_1005 (O_1005,N_24726,N_24535);
or UO_1006 (O_1006,N_24132,N_24313);
or UO_1007 (O_1007,N_24958,N_24619);
or UO_1008 (O_1008,N_24195,N_24201);
nand UO_1009 (O_1009,N_23987,N_24222);
and UO_1010 (O_1010,N_23809,N_24851);
or UO_1011 (O_1011,N_24013,N_23831);
xnor UO_1012 (O_1012,N_24051,N_24342);
nor UO_1013 (O_1013,N_24366,N_24383);
nor UO_1014 (O_1014,N_24458,N_24120);
and UO_1015 (O_1015,N_24510,N_24155);
nand UO_1016 (O_1016,N_24634,N_24995);
nand UO_1017 (O_1017,N_24724,N_24368);
or UO_1018 (O_1018,N_24295,N_23868);
xnor UO_1019 (O_1019,N_24056,N_24196);
or UO_1020 (O_1020,N_24589,N_23912);
and UO_1021 (O_1021,N_24940,N_24780);
nand UO_1022 (O_1022,N_24812,N_24470);
and UO_1023 (O_1023,N_24097,N_24419);
nor UO_1024 (O_1024,N_23850,N_24760);
nor UO_1025 (O_1025,N_23830,N_24839);
or UO_1026 (O_1026,N_24911,N_24124);
and UO_1027 (O_1027,N_24355,N_24446);
nor UO_1028 (O_1028,N_24650,N_24198);
xnor UO_1029 (O_1029,N_24051,N_24547);
nand UO_1030 (O_1030,N_23996,N_24237);
or UO_1031 (O_1031,N_24802,N_23760);
or UO_1032 (O_1032,N_24959,N_24611);
nand UO_1033 (O_1033,N_23780,N_24664);
nor UO_1034 (O_1034,N_24739,N_24000);
xor UO_1035 (O_1035,N_24729,N_24497);
or UO_1036 (O_1036,N_23947,N_24187);
nor UO_1037 (O_1037,N_24713,N_24666);
xnor UO_1038 (O_1038,N_24512,N_24312);
or UO_1039 (O_1039,N_24500,N_23959);
nand UO_1040 (O_1040,N_24672,N_24742);
nor UO_1041 (O_1041,N_23945,N_24221);
xor UO_1042 (O_1042,N_24275,N_24481);
or UO_1043 (O_1043,N_24884,N_24070);
nor UO_1044 (O_1044,N_24486,N_24695);
and UO_1045 (O_1045,N_24953,N_23756);
or UO_1046 (O_1046,N_24225,N_24636);
or UO_1047 (O_1047,N_24497,N_24658);
xor UO_1048 (O_1048,N_24126,N_24914);
nand UO_1049 (O_1049,N_24227,N_24978);
and UO_1050 (O_1050,N_23857,N_24370);
nor UO_1051 (O_1051,N_24449,N_24520);
nand UO_1052 (O_1052,N_24493,N_24754);
and UO_1053 (O_1053,N_24172,N_24898);
nor UO_1054 (O_1054,N_24015,N_24984);
and UO_1055 (O_1055,N_23831,N_24374);
nor UO_1056 (O_1056,N_24215,N_24932);
nand UO_1057 (O_1057,N_24914,N_24116);
nand UO_1058 (O_1058,N_24941,N_24118);
nor UO_1059 (O_1059,N_24954,N_24779);
and UO_1060 (O_1060,N_24461,N_24516);
and UO_1061 (O_1061,N_24477,N_24706);
or UO_1062 (O_1062,N_23838,N_24999);
nand UO_1063 (O_1063,N_24103,N_24160);
or UO_1064 (O_1064,N_24919,N_23767);
nand UO_1065 (O_1065,N_24978,N_24433);
nand UO_1066 (O_1066,N_24030,N_24541);
or UO_1067 (O_1067,N_24045,N_23905);
and UO_1068 (O_1068,N_24844,N_24289);
nor UO_1069 (O_1069,N_24776,N_23751);
and UO_1070 (O_1070,N_24789,N_24947);
xnor UO_1071 (O_1071,N_23772,N_24632);
or UO_1072 (O_1072,N_23860,N_23877);
xor UO_1073 (O_1073,N_24906,N_24196);
xnor UO_1074 (O_1074,N_23830,N_24163);
nor UO_1075 (O_1075,N_24878,N_23992);
nor UO_1076 (O_1076,N_24807,N_24664);
and UO_1077 (O_1077,N_24983,N_24827);
nor UO_1078 (O_1078,N_24242,N_24248);
or UO_1079 (O_1079,N_24773,N_23887);
and UO_1080 (O_1080,N_24395,N_24275);
and UO_1081 (O_1081,N_24345,N_24014);
nor UO_1082 (O_1082,N_24366,N_24670);
and UO_1083 (O_1083,N_23900,N_24613);
xnor UO_1084 (O_1084,N_24587,N_24822);
nor UO_1085 (O_1085,N_24043,N_24009);
and UO_1086 (O_1086,N_24748,N_24686);
nand UO_1087 (O_1087,N_24207,N_23776);
and UO_1088 (O_1088,N_24122,N_24692);
or UO_1089 (O_1089,N_24364,N_24333);
or UO_1090 (O_1090,N_24365,N_24946);
and UO_1091 (O_1091,N_24107,N_24836);
and UO_1092 (O_1092,N_23919,N_24063);
xnor UO_1093 (O_1093,N_24253,N_24281);
nor UO_1094 (O_1094,N_24738,N_24742);
and UO_1095 (O_1095,N_23844,N_23937);
and UO_1096 (O_1096,N_24833,N_23917);
nor UO_1097 (O_1097,N_23986,N_24151);
nand UO_1098 (O_1098,N_24315,N_24384);
and UO_1099 (O_1099,N_24869,N_23866);
nand UO_1100 (O_1100,N_24472,N_24572);
xnor UO_1101 (O_1101,N_24709,N_24552);
nor UO_1102 (O_1102,N_24520,N_23768);
and UO_1103 (O_1103,N_24340,N_24873);
xor UO_1104 (O_1104,N_24295,N_24835);
xor UO_1105 (O_1105,N_24123,N_24754);
nor UO_1106 (O_1106,N_24145,N_23882);
and UO_1107 (O_1107,N_24765,N_24193);
xor UO_1108 (O_1108,N_23825,N_24797);
or UO_1109 (O_1109,N_24722,N_23901);
nand UO_1110 (O_1110,N_23939,N_23970);
nor UO_1111 (O_1111,N_24149,N_24751);
or UO_1112 (O_1112,N_24246,N_23938);
and UO_1113 (O_1113,N_24371,N_24293);
nand UO_1114 (O_1114,N_24125,N_24345);
nand UO_1115 (O_1115,N_23982,N_24355);
xor UO_1116 (O_1116,N_24223,N_24046);
nor UO_1117 (O_1117,N_24255,N_23953);
nand UO_1118 (O_1118,N_24550,N_24588);
nor UO_1119 (O_1119,N_23959,N_24361);
or UO_1120 (O_1120,N_23805,N_24777);
xor UO_1121 (O_1121,N_24448,N_24607);
or UO_1122 (O_1122,N_24831,N_24779);
nand UO_1123 (O_1123,N_24116,N_24763);
or UO_1124 (O_1124,N_23914,N_24235);
and UO_1125 (O_1125,N_23794,N_24127);
and UO_1126 (O_1126,N_23998,N_24005);
nand UO_1127 (O_1127,N_23972,N_24624);
nor UO_1128 (O_1128,N_23886,N_23837);
nand UO_1129 (O_1129,N_24561,N_24327);
xnor UO_1130 (O_1130,N_23924,N_24351);
and UO_1131 (O_1131,N_23990,N_24018);
nand UO_1132 (O_1132,N_24157,N_24790);
nor UO_1133 (O_1133,N_24591,N_24281);
and UO_1134 (O_1134,N_24071,N_24156);
and UO_1135 (O_1135,N_24274,N_23809);
xnor UO_1136 (O_1136,N_24290,N_24870);
nand UO_1137 (O_1137,N_23979,N_24683);
nor UO_1138 (O_1138,N_24452,N_23755);
and UO_1139 (O_1139,N_24587,N_24803);
and UO_1140 (O_1140,N_24129,N_24628);
or UO_1141 (O_1141,N_23963,N_24019);
xor UO_1142 (O_1142,N_24643,N_24612);
nand UO_1143 (O_1143,N_24503,N_24425);
and UO_1144 (O_1144,N_24493,N_24227);
and UO_1145 (O_1145,N_24286,N_24910);
xor UO_1146 (O_1146,N_24678,N_24477);
nand UO_1147 (O_1147,N_23992,N_23959);
or UO_1148 (O_1148,N_23808,N_24836);
xnor UO_1149 (O_1149,N_24346,N_24041);
xor UO_1150 (O_1150,N_24598,N_24020);
nor UO_1151 (O_1151,N_24547,N_23794);
nor UO_1152 (O_1152,N_24749,N_24810);
or UO_1153 (O_1153,N_24987,N_23863);
or UO_1154 (O_1154,N_23860,N_24663);
or UO_1155 (O_1155,N_24390,N_24323);
nor UO_1156 (O_1156,N_23777,N_23833);
or UO_1157 (O_1157,N_24291,N_24961);
nor UO_1158 (O_1158,N_24095,N_24826);
nand UO_1159 (O_1159,N_24952,N_24591);
xnor UO_1160 (O_1160,N_24198,N_23757);
xnor UO_1161 (O_1161,N_24607,N_23786);
nand UO_1162 (O_1162,N_24210,N_24348);
or UO_1163 (O_1163,N_24521,N_24311);
nor UO_1164 (O_1164,N_24600,N_24826);
or UO_1165 (O_1165,N_23848,N_24384);
and UO_1166 (O_1166,N_24821,N_24865);
and UO_1167 (O_1167,N_24496,N_24214);
nand UO_1168 (O_1168,N_24034,N_24087);
and UO_1169 (O_1169,N_23962,N_23926);
nor UO_1170 (O_1170,N_24335,N_23918);
nand UO_1171 (O_1171,N_24178,N_23855);
nor UO_1172 (O_1172,N_24497,N_24555);
nand UO_1173 (O_1173,N_24636,N_24955);
or UO_1174 (O_1174,N_23969,N_23916);
and UO_1175 (O_1175,N_24557,N_24464);
nor UO_1176 (O_1176,N_24905,N_24543);
nor UO_1177 (O_1177,N_24391,N_24438);
and UO_1178 (O_1178,N_24874,N_24776);
nor UO_1179 (O_1179,N_23864,N_24927);
or UO_1180 (O_1180,N_24375,N_24039);
or UO_1181 (O_1181,N_24988,N_24993);
or UO_1182 (O_1182,N_24799,N_24297);
xor UO_1183 (O_1183,N_24096,N_24441);
or UO_1184 (O_1184,N_24511,N_24695);
and UO_1185 (O_1185,N_24250,N_23873);
and UO_1186 (O_1186,N_24467,N_24770);
or UO_1187 (O_1187,N_24028,N_24084);
xor UO_1188 (O_1188,N_23959,N_24321);
or UO_1189 (O_1189,N_24294,N_24511);
nor UO_1190 (O_1190,N_24239,N_24767);
xor UO_1191 (O_1191,N_24399,N_23992);
or UO_1192 (O_1192,N_24794,N_24701);
nor UO_1193 (O_1193,N_24226,N_24904);
xnor UO_1194 (O_1194,N_24515,N_23986);
nor UO_1195 (O_1195,N_24599,N_24385);
xor UO_1196 (O_1196,N_24496,N_24974);
xnor UO_1197 (O_1197,N_23949,N_24116);
nor UO_1198 (O_1198,N_24451,N_23969);
and UO_1199 (O_1199,N_23759,N_24381);
and UO_1200 (O_1200,N_23970,N_24192);
or UO_1201 (O_1201,N_24185,N_24959);
or UO_1202 (O_1202,N_24166,N_24422);
and UO_1203 (O_1203,N_24161,N_23990);
and UO_1204 (O_1204,N_23822,N_23909);
or UO_1205 (O_1205,N_24325,N_24703);
nand UO_1206 (O_1206,N_23975,N_24567);
or UO_1207 (O_1207,N_24589,N_24440);
or UO_1208 (O_1208,N_24860,N_23947);
and UO_1209 (O_1209,N_24893,N_23771);
or UO_1210 (O_1210,N_24909,N_24297);
and UO_1211 (O_1211,N_24651,N_23863);
xnor UO_1212 (O_1212,N_24233,N_24060);
xor UO_1213 (O_1213,N_24375,N_23906);
nor UO_1214 (O_1214,N_24097,N_24637);
xnor UO_1215 (O_1215,N_24848,N_24940);
and UO_1216 (O_1216,N_24546,N_23788);
nor UO_1217 (O_1217,N_24160,N_24560);
nand UO_1218 (O_1218,N_24076,N_23829);
xor UO_1219 (O_1219,N_24306,N_24720);
nor UO_1220 (O_1220,N_24179,N_24191);
nor UO_1221 (O_1221,N_24160,N_24193);
nand UO_1222 (O_1222,N_24253,N_23794);
or UO_1223 (O_1223,N_24029,N_24582);
and UO_1224 (O_1224,N_23874,N_24411);
nand UO_1225 (O_1225,N_24198,N_24312);
xor UO_1226 (O_1226,N_23840,N_23827);
xnor UO_1227 (O_1227,N_23859,N_23910);
nor UO_1228 (O_1228,N_23814,N_23810);
or UO_1229 (O_1229,N_24371,N_24819);
and UO_1230 (O_1230,N_24487,N_23874);
and UO_1231 (O_1231,N_24509,N_23921);
or UO_1232 (O_1232,N_23750,N_23954);
nor UO_1233 (O_1233,N_24536,N_24038);
nor UO_1234 (O_1234,N_24989,N_24049);
nand UO_1235 (O_1235,N_24826,N_24574);
xor UO_1236 (O_1236,N_24010,N_24412);
or UO_1237 (O_1237,N_23826,N_24141);
nor UO_1238 (O_1238,N_24173,N_24493);
or UO_1239 (O_1239,N_24217,N_24102);
and UO_1240 (O_1240,N_24362,N_23992);
xor UO_1241 (O_1241,N_24437,N_23853);
and UO_1242 (O_1242,N_24712,N_24268);
and UO_1243 (O_1243,N_24725,N_24501);
or UO_1244 (O_1244,N_24929,N_24550);
or UO_1245 (O_1245,N_24313,N_24563);
and UO_1246 (O_1246,N_24701,N_24907);
nor UO_1247 (O_1247,N_24465,N_24165);
xnor UO_1248 (O_1248,N_24057,N_24097);
and UO_1249 (O_1249,N_23966,N_24544);
xnor UO_1250 (O_1250,N_24247,N_24732);
and UO_1251 (O_1251,N_24501,N_24433);
and UO_1252 (O_1252,N_24387,N_24369);
and UO_1253 (O_1253,N_24667,N_24951);
xor UO_1254 (O_1254,N_24146,N_24953);
nor UO_1255 (O_1255,N_23923,N_24664);
nor UO_1256 (O_1256,N_24193,N_24795);
nand UO_1257 (O_1257,N_24331,N_24575);
xor UO_1258 (O_1258,N_24690,N_24331);
and UO_1259 (O_1259,N_23906,N_23873);
nand UO_1260 (O_1260,N_24311,N_24623);
nand UO_1261 (O_1261,N_24295,N_24467);
xnor UO_1262 (O_1262,N_24039,N_24061);
nand UO_1263 (O_1263,N_24882,N_24901);
nand UO_1264 (O_1264,N_24196,N_24596);
xor UO_1265 (O_1265,N_24132,N_24128);
nand UO_1266 (O_1266,N_24047,N_24188);
xnor UO_1267 (O_1267,N_24963,N_24642);
and UO_1268 (O_1268,N_23956,N_23964);
nand UO_1269 (O_1269,N_24815,N_24181);
nand UO_1270 (O_1270,N_24242,N_24023);
or UO_1271 (O_1271,N_24375,N_24810);
or UO_1272 (O_1272,N_24956,N_24878);
nor UO_1273 (O_1273,N_23877,N_24242);
nor UO_1274 (O_1274,N_24246,N_24531);
and UO_1275 (O_1275,N_24166,N_23873);
or UO_1276 (O_1276,N_24552,N_24691);
nand UO_1277 (O_1277,N_23940,N_24314);
or UO_1278 (O_1278,N_24111,N_24993);
or UO_1279 (O_1279,N_23912,N_24164);
nand UO_1280 (O_1280,N_23994,N_23978);
nor UO_1281 (O_1281,N_24823,N_24149);
and UO_1282 (O_1282,N_24369,N_23938);
nand UO_1283 (O_1283,N_24321,N_23871);
nor UO_1284 (O_1284,N_24906,N_23958);
or UO_1285 (O_1285,N_23950,N_24446);
xnor UO_1286 (O_1286,N_24338,N_24375);
and UO_1287 (O_1287,N_24354,N_23943);
or UO_1288 (O_1288,N_24208,N_23854);
xor UO_1289 (O_1289,N_24459,N_24000);
nor UO_1290 (O_1290,N_24984,N_24516);
xnor UO_1291 (O_1291,N_24262,N_23846);
or UO_1292 (O_1292,N_24536,N_23808);
and UO_1293 (O_1293,N_23933,N_24959);
xnor UO_1294 (O_1294,N_24599,N_23815);
nor UO_1295 (O_1295,N_24861,N_24044);
nor UO_1296 (O_1296,N_23977,N_23836);
or UO_1297 (O_1297,N_24605,N_24443);
xor UO_1298 (O_1298,N_23891,N_24438);
or UO_1299 (O_1299,N_24971,N_23954);
nor UO_1300 (O_1300,N_24147,N_24627);
and UO_1301 (O_1301,N_24760,N_24366);
nor UO_1302 (O_1302,N_23862,N_24433);
nand UO_1303 (O_1303,N_24251,N_23950);
nand UO_1304 (O_1304,N_24803,N_23858);
or UO_1305 (O_1305,N_24072,N_24328);
xor UO_1306 (O_1306,N_23891,N_24257);
or UO_1307 (O_1307,N_24404,N_24659);
and UO_1308 (O_1308,N_24634,N_24786);
xnor UO_1309 (O_1309,N_24213,N_24140);
xnor UO_1310 (O_1310,N_24383,N_24320);
xor UO_1311 (O_1311,N_23930,N_24766);
nor UO_1312 (O_1312,N_23830,N_24953);
xnor UO_1313 (O_1313,N_24250,N_24426);
and UO_1314 (O_1314,N_24441,N_24046);
nor UO_1315 (O_1315,N_24529,N_24449);
and UO_1316 (O_1316,N_24309,N_24220);
xor UO_1317 (O_1317,N_24648,N_24557);
and UO_1318 (O_1318,N_24084,N_24371);
or UO_1319 (O_1319,N_24200,N_24947);
or UO_1320 (O_1320,N_24963,N_23888);
or UO_1321 (O_1321,N_23936,N_24576);
and UO_1322 (O_1322,N_24135,N_24082);
nor UO_1323 (O_1323,N_24985,N_24792);
nand UO_1324 (O_1324,N_24935,N_24170);
nor UO_1325 (O_1325,N_24114,N_24545);
or UO_1326 (O_1326,N_24096,N_24228);
nor UO_1327 (O_1327,N_24163,N_24190);
nor UO_1328 (O_1328,N_24586,N_24490);
nand UO_1329 (O_1329,N_24018,N_24654);
nand UO_1330 (O_1330,N_24067,N_24900);
nand UO_1331 (O_1331,N_24403,N_24280);
nor UO_1332 (O_1332,N_24004,N_24081);
xnor UO_1333 (O_1333,N_24726,N_23903);
nor UO_1334 (O_1334,N_24172,N_24435);
or UO_1335 (O_1335,N_24789,N_24243);
nand UO_1336 (O_1336,N_24767,N_24646);
xor UO_1337 (O_1337,N_24593,N_24134);
nand UO_1338 (O_1338,N_24526,N_24875);
nor UO_1339 (O_1339,N_24239,N_23802);
nand UO_1340 (O_1340,N_24890,N_24782);
xor UO_1341 (O_1341,N_24612,N_24465);
or UO_1342 (O_1342,N_24181,N_24873);
nand UO_1343 (O_1343,N_24524,N_24758);
xor UO_1344 (O_1344,N_24566,N_23780);
nor UO_1345 (O_1345,N_23910,N_24709);
and UO_1346 (O_1346,N_23943,N_24080);
nor UO_1347 (O_1347,N_24148,N_24953);
nor UO_1348 (O_1348,N_24946,N_24228);
xnor UO_1349 (O_1349,N_24146,N_24362);
xor UO_1350 (O_1350,N_24149,N_24404);
or UO_1351 (O_1351,N_24557,N_24437);
and UO_1352 (O_1352,N_24579,N_23886);
nor UO_1353 (O_1353,N_24711,N_24139);
nor UO_1354 (O_1354,N_24529,N_23941);
nand UO_1355 (O_1355,N_24320,N_24475);
and UO_1356 (O_1356,N_24244,N_24437);
nand UO_1357 (O_1357,N_24356,N_24812);
xnor UO_1358 (O_1358,N_24479,N_24586);
or UO_1359 (O_1359,N_23900,N_24061);
and UO_1360 (O_1360,N_24597,N_24348);
nand UO_1361 (O_1361,N_24475,N_24871);
and UO_1362 (O_1362,N_24102,N_24529);
nor UO_1363 (O_1363,N_24565,N_24381);
nand UO_1364 (O_1364,N_24501,N_24049);
nand UO_1365 (O_1365,N_24769,N_23935);
nand UO_1366 (O_1366,N_24548,N_24442);
xnor UO_1367 (O_1367,N_23752,N_24108);
xnor UO_1368 (O_1368,N_24706,N_24808);
nand UO_1369 (O_1369,N_24352,N_24439);
xor UO_1370 (O_1370,N_24994,N_24311);
nand UO_1371 (O_1371,N_24994,N_24071);
nor UO_1372 (O_1372,N_23915,N_24728);
or UO_1373 (O_1373,N_23775,N_24486);
nor UO_1374 (O_1374,N_23766,N_24487);
and UO_1375 (O_1375,N_23827,N_24962);
xnor UO_1376 (O_1376,N_24269,N_24076);
xor UO_1377 (O_1377,N_24707,N_24754);
xnor UO_1378 (O_1378,N_23900,N_24294);
xnor UO_1379 (O_1379,N_24690,N_24634);
xor UO_1380 (O_1380,N_24131,N_24820);
nand UO_1381 (O_1381,N_24947,N_24170);
and UO_1382 (O_1382,N_24278,N_23812);
nand UO_1383 (O_1383,N_24904,N_24377);
nor UO_1384 (O_1384,N_24756,N_24231);
or UO_1385 (O_1385,N_24345,N_24256);
or UO_1386 (O_1386,N_24705,N_24665);
xor UO_1387 (O_1387,N_24581,N_23842);
xnor UO_1388 (O_1388,N_23797,N_24155);
nor UO_1389 (O_1389,N_24732,N_24830);
or UO_1390 (O_1390,N_24808,N_24058);
or UO_1391 (O_1391,N_24815,N_24973);
and UO_1392 (O_1392,N_24847,N_24515);
nor UO_1393 (O_1393,N_24288,N_24929);
or UO_1394 (O_1394,N_23866,N_24100);
and UO_1395 (O_1395,N_24753,N_24985);
or UO_1396 (O_1396,N_24341,N_24918);
and UO_1397 (O_1397,N_24742,N_24468);
and UO_1398 (O_1398,N_24063,N_24010);
nor UO_1399 (O_1399,N_24146,N_24239);
or UO_1400 (O_1400,N_23859,N_24950);
or UO_1401 (O_1401,N_24914,N_24502);
xor UO_1402 (O_1402,N_24005,N_24835);
nor UO_1403 (O_1403,N_24582,N_23778);
nor UO_1404 (O_1404,N_24675,N_23829);
nor UO_1405 (O_1405,N_24335,N_23961);
nand UO_1406 (O_1406,N_24853,N_24807);
nor UO_1407 (O_1407,N_24300,N_23917);
xnor UO_1408 (O_1408,N_24910,N_24062);
nand UO_1409 (O_1409,N_24906,N_24606);
xor UO_1410 (O_1410,N_24421,N_23912);
and UO_1411 (O_1411,N_24323,N_24896);
xor UO_1412 (O_1412,N_24376,N_24586);
nor UO_1413 (O_1413,N_24010,N_24918);
xor UO_1414 (O_1414,N_23888,N_24330);
or UO_1415 (O_1415,N_24786,N_23934);
nor UO_1416 (O_1416,N_24735,N_24209);
and UO_1417 (O_1417,N_24999,N_24126);
and UO_1418 (O_1418,N_24653,N_24035);
nor UO_1419 (O_1419,N_24435,N_24654);
nand UO_1420 (O_1420,N_24425,N_24473);
or UO_1421 (O_1421,N_24652,N_24751);
xnor UO_1422 (O_1422,N_24112,N_23978);
nand UO_1423 (O_1423,N_24256,N_24545);
or UO_1424 (O_1424,N_24492,N_24065);
and UO_1425 (O_1425,N_24758,N_24847);
and UO_1426 (O_1426,N_24676,N_24734);
nor UO_1427 (O_1427,N_24195,N_24146);
or UO_1428 (O_1428,N_24976,N_24150);
xor UO_1429 (O_1429,N_24710,N_24866);
xnor UO_1430 (O_1430,N_24720,N_24581);
or UO_1431 (O_1431,N_24467,N_24409);
nor UO_1432 (O_1432,N_24904,N_24096);
nor UO_1433 (O_1433,N_24697,N_24291);
and UO_1434 (O_1434,N_24242,N_24331);
nand UO_1435 (O_1435,N_24463,N_24220);
or UO_1436 (O_1436,N_23769,N_24228);
and UO_1437 (O_1437,N_23769,N_24279);
and UO_1438 (O_1438,N_24316,N_24955);
or UO_1439 (O_1439,N_23966,N_24539);
or UO_1440 (O_1440,N_23914,N_24539);
nor UO_1441 (O_1441,N_23773,N_24124);
xnor UO_1442 (O_1442,N_24213,N_24555);
xnor UO_1443 (O_1443,N_23882,N_23757);
nor UO_1444 (O_1444,N_23878,N_24277);
and UO_1445 (O_1445,N_24722,N_24755);
and UO_1446 (O_1446,N_23939,N_24956);
nand UO_1447 (O_1447,N_24389,N_24327);
and UO_1448 (O_1448,N_24332,N_24602);
xor UO_1449 (O_1449,N_23859,N_23895);
and UO_1450 (O_1450,N_24942,N_24367);
xor UO_1451 (O_1451,N_24820,N_24816);
and UO_1452 (O_1452,N_24557,N_24158);
and UO_1453 (O_1453,N_24988,N_23858);
nor UO_1454 (O_1454,N_24554,N_24837);
nor UO_1455 (O_1455,N_23867,N_23888);
xor UO_1456 (O_1456,N_24858,N_24389);
xor UO_1457 (O_1457,N_24614,N_24058);
nand UO_1458 (O_1458,N_24648,N_23916);
nand UO_1459 (O_1459,N_24663,N_24792);
or UO_1460 (O_1460,N_23840,N_24557);
or UO_1461 (O_1461,N_24554,N_24726);
xor UO_1462 (O_1462,N_24814,N_24782);
and UO_1463 (O_1463,N_24051,N_24910);
nor UO_1464 (O_1464,N_24133,N_24475);
nand UO_1465 (O_1465,N_23931,N_24511);
xor UO_1466 (O_1466,N_24619,N_24825);
or UO_1467 (O_1467,N_24893,N_24884);
xnor UO_1468 (O_1468,N_24617,N_24150);
or UO_1469 (O_1469,N_23878,N_24713);
or UO_1470 (O_1470,N_23767,N_24912);
xor UO_1471 (O_1471,N_23978,N_24148);
xnor UO_1472 (O_1472,N_24382,N_24189);
xnor UO_1473 (O_1473,N_24926,N_23806);
xor UO_1474 (O_1474,N_24781,N_24631);
and UO_1475 (O_1475,N_23757,N_24503);
or UO_1476 (O_1476,N_23823,N_23979);
and UO_1477 (O_1477,N_23921,N_24708);
xor UO_1478 (O_1478,N_24815,N_23783);
and UO_1479 (O_1479,N_24665,N_24558);
and UO_1480 (O_1480,N_24759,N_24576);
nand UO_1481 (O_1481,N_23977,N_23751);
nor UO_1482 (O_1482,N_23834,N_24892);
and UO_1483 (O_1483,N_24192,N_24368);
or UO_1484 (O_1484,N_24807,N_24102);
nor UO_1485 (O_1485,N_24407,N_23878);
or UO_1486 (O_1486,N_24435,N_24258);
xnor UO_1487 (O_1487,N_23867,N_24698);
or UO_1488 (O_1488,N_24452,N_23986);
nand UO_1489 (O_1489,N_24417,N_24967);
nor UO_1490 (O_1490,N_24988,N_24198);
and UO_1491 (O_1491,N_24781,N_24323);
nand UO_1492 (O_1492,N_24127,N_24547);
nor UO_1493 (O_1493,N_24695,N_24340);
and UO_1494 (O_1494,N_24008,N_24494);
nor UO_1495 (O_1495,N_24641,N_23878);
nor UO_1496 (O_1496,N_23814,N_23972);
and UO_1497 (O_1497,N_24975,N_24052);
nor UO_1498 (O_1498,N_24823,N_24540);
xor UO_1499 (O_1499,N_24645,N_23920);
nor UO_1500 (O_1500,N_23914,N_24553);
nor UO_1501 (O_1501,N_23981,N_24908);
xor UO_1502 (O_1502,N_23975,N_24576);
and UO_1503 (O_1503,N_24927,N_24804);
xor UO_1504 (O_1504,N_23816,N_24088);
nor UO_1505 (O_1505,N_24465,N_23774);
nor UO_1506 (O_1506,N_24534,N_24714);
or UO_1507 (O_1507,N_24238,N_24366);
xor UO_1508 (O_1508,N_24580,N_24190);
and UO_1509 (O_1509,N_24090,N_24470);
or UO_1510 (O_1510,N_24818,N_24604);
nand UO_1511 (O_1511,N_23765,N_24264);
xor UO_1512 (O_1512,N_23921,N_24347);
or UO_1513 (O_1513,N_24017,N_24470);
or UO_1514 (O_1514,N_24443,N_23930);
and UO_1515 (O_1515,N_24742,N_24880);
or UO_1516 (O_1516,N_24531,N_24177);
and UO_1517 (O_1517,N_24960,N_24756);
and UO_1518 (O_1518,N_23780,N_24584);
and UO_1519 (O_1519,N_23939,N_24983);
nor UO_1520 (O_1520,N_23905,N_24004);
or UO_1521 (O_1521,N_24564,N_24274);
nor UO_1522 (O_1522,N_23847,N_24419);
or UO_1523 (O_1523,N_24692,N_24635);
xnor UO_1524 (O_1524,N_23869,N_24761);
nand UO_1525 (O_1525,N_24467,N_24625);
nor UO_1526 (O_1526,N_24126,N_23806);
nand UO_1527 (O_1527,N_24936,N_24524);
and UO_1528 (O_1528,N_24488,N_24213);
nand UO_1529 (O_1529,N_24601,N_24900);
and UO_1530 (O_1530,N_24480,N_24328);
or UO_1531 (O_1531,N_23904,N_24547);
or UO_1532 (O_1532,N_24546,N_24312);
xnor UO_1533 (O_1533,N_24648,N_23917);
nor UO_1534 (O_1534,N_24480,N_23875);
and UO_1535 (O_1535,N_23841,N_24537);
xor UO_1536 (O_1536,N_23806,N_24222);
or UO_1537 (O_1537,N_24143,N_24439);
xnor UO_1538 (O_1538,N_24152,N_23955);
and UO_1539 (O_1539,N_24689,N_24990);
nor UO_1540 (O_1540,N_24684,N_24087);
or UO_1541 (O_1541,N_24944,N_24672);
nand UO_1542 (O_1542,N_24734,N_24570);
nor UO_1543 (O_1543,N_24213,N_23999);
xor UO_1544 (O_1544,N_24433,N_24397);
or UO_1545 (O_1545,N_24460,N_24052);
xor UO_1546 (O_1546,N_24767,N_24083);
xnor UO_1547 (O_1547,N_24671,N_24698);
nand UO_1548 (O_1548,N_24887,N_24711);
xor UO_1549 (O_1549,N_24106,N_24763);
or UO_1550 (O_1550,N_23763,N_24301);
or UO_1551 (O_1551,N_24949,N_24186);
or UO_1552 (O_1552,N_23838,N_24252);
xor UO_1553 (O_1553,N_24859,N_24256);
nand UO_1554 (O_1554,N_24370,N_24649);
or UO_1555 (O_1555,N_24638,N_24409);
xor UO_1556 (O_1556,N_24279,N_24224);
and UO_1557 (O_1557,N_24488,N_24627);
nand UO_1558 (O_1558,N_24783,N_24424);
and UO_1559 (O_1559,N_24744,N_24795);
and UO_1560 (O_1560,N_24145,N_23987);
and UO_1561 (O_1561,N_24349,N_24629);
nor UO_1562 (O_1562,N_24464,N_24646);
and UO_1563 (O_1563,N_24170,N_24679);
nor UO_1564 (O_1564,N_23927,N_24356);
nor UO_1565 (O_1565,N_24053,N_24034);
and UO_1566 (O_1566,N_24647,N_24522);
nor UO_1567 (O_1567,N_24793,N_24279);
nand UO_1568 (O_1568,N_24655,N_24276);
nand UO_1569 (O_1569,N_24555,N_24144);
nor UO_1570 (O_1570,N_24170,N_24523);
or UO_1571 (O_1571,N_24602,N_24105);
nor UO_1572 (O_1572,N_24435,N_24279);
or UO_1573 (O_1573,N_24684,N_24119);
and UO_1574 (O_1574,N_23773,N_24801);
or UO_1575 (O_1575,N_24206,N_24318);
or UO_1576 (O_1576,N_24557,N_24122);
nand UO_1577 (O_1577,N_24646,N_24664);
or UO_1578 (O_1578,N_24417,N_24622);
xnor UO_1579 (O_1579,N_24473,N_24204);
and UO_1580 (O_1580,N_23772,N_24592);
nand UO_1581 (O_1581,N_24278,N_24387);
and UO_1582 (O_1582,N_24659,N_24416);
and UO_1583 (O_1583,N_24192,N_24948);
nor UO_1584 (O_1584,N_24635,N_24793);
xor UO_1585 (O_1585,N_24826,N_24963);
nand UO_1586 (O_1586,N_24996,N_24008);
or UO_1587 (O_1587,N_24007,N_24550);
nor UO_1588 (O_1588,N_24405,N_23780);
and UO_1589 (O_1589,N_24143,N_24026);
and UO_1590 (O_1590,N_24417,N_23898);
xnor UO_1591 (O_1591,N_23895,N_24608);
or UO_1592 (O_1592,N_24548,N_24531);
nor UO_1593 (O_1593,N_23772,N_24444);
nor UO_1594 (O_1594,N_24184,N_24694);
nand UO_1595 (O_1595,N_24829,N_24868);
or UO_1596 (O_1596,N_24260,N_24562);
nand UO_1597 (O_1597,N_24161,N_24287);
nor UO_1598 (O_1598,N_24340,N_23794);
and UO_1599 (O_1599,N_24631,N_24911);
nor UO_1600 (O_1600,N_24098,N_24027);
nor UO_1601 (O_1601,N_23774,N_23822);
nor UO_1602 (O_1602,N_24812,N_24926);
nand UO_1603 (O_1603,N_24492,N_24745);
xnor UO_1604 (O_1604,N_23962,N_23927);
nor UO_1605 (O_1605,N_24736,N_24607);
and UO_1606 (O_1606,N_24838,N_24724);
nor UO_1607 (O_1607,N_24687,N_24144);
and UO_1608 (O_1608,N_24934,N_24325);
nor UO_1609 (O_1609,N_23767,N_24016);
nor UO_1610 (O_1610,N_24396,N_24912);
and UO_1611 (O_1611,N_24621,N_23758);
nand UO_1612 (O_1612,N_23815,N_24654);
nor UO_1613 (O_1613,N_24837,N_23792);
and UO_1614 (O_1614,N_24919,N_24487);
xnor UO_1615 (O_1615,N_24392,N_24962);
xnor UO_1616 (O_1616,N_24387,N_24329);
or UO_1617 (O_1617,N_23838,N_24718);
or UO_1618 (O_1618,N_24964,N_24589);
nor UO_1619 (O_1619,N_24942,N_24238);
and UO_1620 (O_1620,N_24008,N_24200);
and UO_1621 (O_1621,N_24619,N_24644);
nand UO_1622 (O_1622,N_24594,N_23859);
or UO_1623 (O_1623,N_24818,N_23790);
or UO_1624 (O_1624,N_24530,N_24629);
and UO_1625 (O_1625,N_24285,N_24573);
or UO_1626 (O_1626,N_24559,N_24696);
nor UO_1627 (O_1627,N_24529,N_23828);
nor UO_1628 (O_1628,N_24276,N_24322);
or UO_1629 (O_1629,N_24596,N_24198);
and UO_1630 (O_1630,N_24546,N_24834);
or UO_1631 (O_1631,N_23909,N_24627);
or UO_1632 (O_1632,N_23790,N_24420);
or UO_1633 (O_1633,N_24116,N_24787);
xor UO_1634 (O_1634,N_24946,N_24940);
and UO_1635 (O_1635,N_24967,N_24672);
xor UO_1636 (O_1636,N_24015,N_24961);
nor UO_1637 (O_1637,N_23875,N_23866);
and UO_1638 (O_1638,N_23842,N_24377);
or UO_1639 (O_1639,N_24769,N_24264);
xnor UO_1640 (O_1640,N_23927,N_23806);
nor UO_1641 (O_1641,N_24598,N_23893);
nand UO_1642 (O_1642,N_24569,N_24504);
and UO_1643 (O_1643,N_24169,N_24246);
or UO_1644 (O_1644,N_24063,N_23850);
and UO_1645 (O_1645,N_23837,N_24460);
and UO_1646 (O_1646,N_24077,N_24051);
xnor UO_1647 (O_1647,N_24159,N_24336);
nor UO_1648 (O_1648,N_23985,N_24151);
nor UO_1649 (O_1649,N_23773,N_24610);
xnor UO_1650 (O_1650,N_24093,N_24741);
xor UO_1651 (O_1651,N_24272,N_24987);
xnor UO_1652 (O_1652,N_24912,N_24672);
nor UO_1653 (O_1653,N_24419,N_23893);
and UO_1654 (O_1654,N_24976,N_23941);
nand UO_1655 (O_1655,N_24312,N_23851);
nor UO_1656 (O_1656,N_24350,N_23869);
xnor UO_1657 (O_1657,N_24064,N_24137);
nor UO_1658 (O_1658,N_24723,N_24694);
or UO_1659 (O_1659,N_24633,N_24297);
nand UO_1660 (O_1660,N_24891,N_23965);
and UO_1661 (O_1661,N_24986,N_24051);
nand UO_1662 (O_1662,N_24649,N_24494);
and UO_1663 (O_1663,N_24798,N_24944);
nand UO_1664 (O_1664,N_23822,N_24727);
and UO_1665 (O_1665,N_24759,N_24679);
nor UO_1666 (O_1666,N_23755,N_24136);
nand UO_1667 (O_1667,N_24636,N_24459);
nand UO_1668 (O_1668,N_23985,N_23754);
nor UO_1669 (O_1669,N_24772,N_24177);
and UO_1670 (O_1670,N_24275,N_24555);
nor UO_1671 (O_1671,N_23942,N_24282);
xor UO_1672 (O_1672,N_24342,N_24973);
nor UO_1673 (O_1673,N_24251,N_24940);
nand UO_1674 (O_1674,N_24022,N_24519);
nand UO_1675 (O_1675,N_23939,N_24823);
and UO_1676 (O_1676,N_24516,N_23916);
nor UO_1677 (O_1677,N_24807,N_24356);
and UO_1678 (O_1678,N_24455,N_24146);
xor UO_1679 (O_1679,N_24083,N_24130);
xor UO_1680 (O_1680,N_24750,N_24503);
nand UO_1681 (O_1681,N_24273,N_24649);
and UO_1682 (O_1682,N_24427,N_24941);
and UO_1683 (O_1683,N_24121,N_24482);
and UO_1684 (O_1684,N_24877,N_24745);
nand UO_1685 (O_1685,N_24715,N_24968);
nor UO_1686 (O_1686,N_24402,N_24668);
xor UO_1687 (O_1687,N_24320,N_24959);
and UO_1688 (O_1688,N_24782,N_23787);
nand UO_1689 (O_1689,N_24092,N_24448);
nor UO_1690 (O_1690,N_24183,N_23809);
or UO_1691 (O_1691,N_23767,N_24382);
nor UO_1692 (O_1692,N_24924,N_24446);
nand UO_1693 (O_1693,N_24591,N_24864);
nand UO_1694 (O_1694,N_24033,N_24627);
nand UO_1695 (O_1695,N_23975,N_24464);
nand UO_1696 (O_1696,N_24600,N_24177);
xor UO_1697 (O_1697,N_24999,N_23899);
xnor UO_1698 (O_1698,N_24777,N_24574);
nand UO_1699 (O_1699,N_24124,N_24311);
or UO_1700 (O_1700,N_23891,N_24726);
and UO_1701 (O_1701,N_24112,N_24050);
nand UO_1702 (O_1702,N_24658,N_23977);
or UO_1703 (O_1703,N_24008,N_24416);
nor UO_1704 (O_1704,N_24602,N_24683);
nor UO_1705 (O_1705,N_24426,N_24203);
nor UO_1706 (O_1706,N_24118,N_24979);
nand UO_1707 (O_1707,N_23952,N_24157);
nand UO_1708 (O_1708,N_24197,N_24970);
nor UO_1709 (O_1709,N_24435,N_24143);
and UO_1710 (O_1710,N_23794,N_23936);
or UO_1711 (O_1711,N_24720,N_24915);
and UO_1712 (O_1712,N_24939,N_23956);
xor UO_1713 (O_1713,N_23978,N_24633);
or UO_1714 (O_1714,N_24470,N_23855);
or UO_1715 (O_1715,N_24308,N_24481);
nor UO_1716 (O_1716,N_24078,N_24344);
nor UO_1717 (O_1717,N_24337,N_24284);
or UO_1718 (O_1718,N_24280,N_24811);
nor UO_1719 (O_1719,N_24892,N_24203);
nand UO_1720 (O_1720,N_24923,N_24019);
and UO_1721 (O_1721,N_23886,N_24356);
xor UO_1722 (O_1722,N_24620,N_24192);
or UO_1723 (O_1723,N_24911,N_23799);
and UO_1724 (O_1724,N_23754,N_24619);
xor UO_1725 (O_1725,N_23794,N_24661);
xnor UO_1726 (O_1726,N_23987,N_24240);
nor UO_1727 (O_1727,N_24778,N_24768);
nor UO_1728 (O_1728,N_24597,N_23879);
or UO_1729 (O_1729,N_24249,N_24422);
xor UO_1730 (O_1730,N_24996,N_24544);
or UO_1731 (O_1731,N_24001,N_24515);
and UO_1732 (O_1732,N_24747,N_24814);
nor UO_1733 (O_1733,N_24944,N_24265);
nor UO_1734 (O_1734,N_24303,N_23837);
and UO_1735 (O_1735,N_24444,N_24529);
and UO_1736 (O_1736,N_24239,N_24472);
or UO_1737 (O_1737,N_24281,N_24128);
and UO_1738 (O_1738,N_24389,N_24183);
nand UO_1739 (O_1739,N_24402,N_24443);
and UO_1740 (O_1740,N_23750,N_24074);
xnor UO_1741 (O_1741,N_24377,N_24330);
nor UO_1742 (O_1742,N_24909,N_23784);
xor UO_1743 (O_1743,N_24995,N_23855);
or UO_1744 (O_1744,N_23835,N_24133);
xnor UO_1745 (O_1745,N_24680,N_24758);
or UO_1746 (O_1746,N_24610,N_24314);
and UO_1747 (O_1747,N_23989,N_24972);
xnor UO_1748 (O_1748,N_24314,N_23789);
nand UO_1749 (O_1749,N_24050,N_24584);
or UO_1750 (O_1750,N_23751,N_24842);
nor UO_1751 (O_1751,N_24178,N_23827);
nand UO_1752 (O_1752,N_24369,N_24506);
xor UO_1753 (O_1753,N_24630,N_24393);
and UO_1754 (O_1754,N_24568,N_24176);
nand UO_1755 (O_1755,N_24555,N_24896);
xor UO_1756 (O_1756,N_24680,N_24588);
nor UO_1757 (O_1757,N_23918,N_23864);
xor UO_1758 (O_1758,N_24086,N_24686);
nand UO_1759 (O_1759,N_24903,N_24545);
and UO_1760 (O_1760,N_24141,N_24904);
and UO_1761 (O_1761,N_24426,N_23775);
nand UO_1762 (O_1762,N_24464,N_24731);
or UO_1763 (O_1763,N_24102,N_23916);
or UO_1764 (O_1764,N_24450,N_24624);
and UO_1765 (O_1765,N_24267,N_23889);
or UO_1766 (O_1766,N_24810,N_24236);
or UO_1767 (O_1767,N_24324,N_24136);
nand UO_1768 (O_1768,N_24197,N_24500);
nand UO_1769 (O_1769,N_24342,N_24205);
nand UO_1770 (O_1770,N_23829,N_24533);
nor UO_1771 (O_1771,N_23984,N_24640);
or UO_1772 (O_1772,N_24992,N_24555);
and UO_1773 (O_1773,N_24808,N_24500);
nor UO_1774 (O_1774,N_24747,N_24578);
and UO_1775 (O_1775,N_24665,N_24878);
nor UO_1776 (O_1776,N_23841,N_24696);
and UO_1777 (O_1777,N_23872,N_23758);
and UO_1778 (O_1778,N_24442,N_24264);
nor UO_1779 (O_1779,N_24059,N_24694);
nand UO_1780 (O_1780,N_24276,N_24008);
nor UO_1781 (O_1781,N_24846,N_23861);
xor UO_1782 (O_1782,N_24599,N_24285);
xor UO_1783 (O_1783,N_24771,N_24328);
nor UO_1784 (O_1784,N_24272,N_24334);
nor UO_1785 (O_1785,N_24397,N_24253);
and UO_1786 (O_1786,N_23956,N_24958);
nand UO_1787 (O_1787,N_24804,N_24941);
and UO_1788 (O_1788,N_24092,N_24083);
nor UO_1789 (O_1789,N_23967,N_24005);
and UO_1790 (O_1790,N_24820,N_24439);
nand UO_1791 (O_1791,N_24259,N_24290);
or UO_1792 (O_1792,N_24790,N_24365);
nand UO_1793 (O_1793,N_23881,N_24733);
and UO_1794 (O_1794,N_24336,N_24663);
and UO_1795 (O_1795,N_24237,N_23831);
nand UO_1796 (O_1796,N_24794,N_23861);
nand UO_1797 (O_1797,N_24592,N_24508);
nor UO_1798 (O_1798,N_24854,N_23909);
nor UO_1799 (O_1799,N_24596,N_24379);
xor UO_1800 (O_1800,N_24705,N_24084);
and UO_1801 (O_1801,N_24129,N_24694);
nor UO_1802 (O_1802,N_23884,N_23868);
or UO_1803 (O_1803,N_24980,N_24836);
and UO_1804 (O_1804,N_24666,N_23874);
or UO_1805 (O_1805,N_23905,N_24588);
xnor UO_1806 (O_1806,N_24398,N_24182);
nand UO_1807 (O_1807,N_24052,N_24564);
nand UO_1808 (O_1808,N_24806,N_24597);
nand UO_1809 (O_1809,N_23876,N_24545);
xnor UO_1810 (O_1810,N_24524,N_24484);
nor UO_1811 (O_1811,N_24349,N_24900);
nor UO_1812 (O_1812,N_24603,N_24877);
nor UO_1813 (O_1813,N_24164,N_24776);
nor UO_1814 (O_1814,N_24066,N_23832);
or UO_1815 (O_1815,N_24451,N_24496);
xor UO_1816 (O_1816,N_24152,N_23758);
xnor UO_1817 (O_1817,N_23953,N_24274);
nand UO_1818 (O_1818,N_24484,N_24784);
nor UO_1819 (O_1819,N_24642,N_24426);
or UO_1820 (O_1820,N_24017,N_24316);
nand UO_1821 (O_1821,N_24881,N_23858);
xor UO_1822 (O_1822,N_24352,N_23963);
nor UO_1823 (O_1823,N_24766,N_24699);
nor UO_1824 (O_1824,N_24899,N_24020);
and UO_1825 (O_1825,N_24859,N_23994);
and UO_1826 (O_1826,N_24252,N_24113);
xnor UO_1827 (O_1827,N_24440,N_23778);
nor UO_1828 (O_1828,N_24932,N_24050);
or UO_1829 (O_1829,N_23841,N_24993);
nand UO_1830 (O_1830,N_24929,N_24709);
xnor UO_1831 (O_1831,N_24684,N_24301);
nand UO_1832 (O_1832,N_24744,N_24041);
nor UO_1833 (O_1833,N_24467,N_23941);
nand UO_1834 (O_1834,N_24905,N_24582);
or UO_1835 (O_1835,N_24903,N_24221);
nor UO_1836 (O_1836,N_24737,N_23924);
nor UO_1837 (O_1837,N_23903,N_24986);
nand UO_1838 (O_1838,N_24697,N_24618);
xnor UO_1839 (O_1839,N_24122,N_24600);
xor UO_1840 (O_1840,N_24150,N_23759);
or UO_1841 (O_1841,N_24907,N_24232);
or UO_1842 (O_1842,N_24689,N_24421);
or UO_1843 (O_1843,N_24252,N_24432);
nand UO_1844 (O_1844,N_24351,N_24352);
xnor UO_1845 (O_1845,N_24354,N_24319);
xor UO_1846 (O_1846,N_24408,N_23889);
and UO_1847 (O_1847,N_23995,N_24481);
nor UO_1848 (O_1848,N_24332,N_24894);
nand UO_1849 (O_1849,N_24057,N_24516);
nand UO_1850 (O_1850,N_23911,N_24050);
nand UO_1851 (O_1851,N_23778,N_24270);
nor UO_1852 (O_1852,N_24892,N_24527);
nor UO_1853 (O_1853,N_23856,N_24334);
nor UO_1854 (O_1854,N_24646,N_24407);
nor UO_1855 (O_1855,N_24453,N_24785);
nor UO_1856 (O_1856,N_23869,N_24219);
or UO_1857 (O_1857,N_24108,N_23966);
or UO_1858 (O_1858,N_24082,N_24949);
or UO_1859 (O_1859,N_24731,N_23851);
nand UO_1860 (O_1860,N_24188,N_23859);
and UO_1861 (O_1861,N_24112,N_24779);
xnor UO_1862 (O_1862,N_24191,N_24471);
nor UO_1863 (O_1863,N_24026,N_23824);
xor UO_1864 (O_1864,N_24625,N_24775);
nand UO_1865 (O_1865,N_23984,N_24882);
nand UO_1866 (O_1866,N_24764,N_24491);
and UO_1867 (O_1867,N_23840,N_24152);
nor UO_1868 (O_1868,N_24443,N_24459);
or UO_1869 (O_1869,N_24821,N_24866);
xnor UO_1870 (O_1870,N_24027,N_24612);
nor UO_1871 (O_1871,N_24540,N_24955);
nand UO_1872 (O_1872,N_23803,N_23866);
and UO_1873 (O_1873,N_24740,N_24102);
and UO_1874 (O_1874,N_24204,N_24496);
and UO_1875 (O_1875,N_24979,N_24332);
nand UO_1876 (O_1876,N_24027,N_24351);
nand UO_1877 (O_1877,N_23832,N_24909);
xnor UO_1878 (O_1878,N_24497,N_23985);
xor UO_1879 (O_1879,N_24345,N_23809);
xnor UO_1880 (O_1880,N_24708,N_24842);
and UO_1881 (O_1881,N_23863,N_24474);
or UO_1882 (O_1882,N_24443,N_24869);
and UO_1883 (O_1883,N_24530,N_23795);
xnor UO_1884 (O_1884,N_24946,N_24685);
or UO_1885 (O_1885,N_24917,N_24848);
nand UO_1886 (O_1886,N_23838,N_24753);
xnor UO_1887 (O_1887,N_23862,N_24194);
nand UO_1888 (O_1888,N_23806,N_24937);
nor UO_1889 (O_1889,N_23983,N_23816);
xor UO_1890 (O_1890,N_24190,N_24821);
xor UO_1891 (O_1891,N_24239,N_24837);
xnor UO_1892 (O_1892,N_24462,N_23812);
xnor UO_1893 (O_1893,N_24887,N_24677);
nor UO_1894 (O_1894,N_24597,N_24564);
and UO_1895 (O_1895,N_24123,N_23815);
or UO_1896 (O_1896,N_24767,N_24564);
and UO_1897 (O_1897,N_24717,N_24988);
or UO_1898 (O_1898,N_23884,N_24584);
nor UO_1899 (O_1899,N_24700,N_24450);
nand UO_1900 (O_1900,N_24283,N_24514);
xor UO_1901 (O_1901,N_24913,N_24739);
and UO_1902 (O_1902,N_24993,N_24016);
xor UO_1903 (O_1903,N_23879,N_24834);
or UO_1904 (O_1904,N_24020,N_24632);
or UO_1905 (O_1905,N_24645,N_24759);
nand UO_1906 (O_1906,N_24512,N_24330);
nand UO_1907 (O_1907,N_23878,N_24939);
nand UO_1908 (O_1908,N_24770,N_23838);
xor UO_1909 (O_1909,N_24178,N_24157);
nor UO_1910 (O_1910,N_24176,N_23980);
or UO_1911 (O_1911,N_23869,N_23925);
xor UO_1912 (O_1912,N_24366,N_23909);
xnor UO_1913 (O_1913,N_23956,N_23857);
and UO_1914 (O_1914,N_24002,N_24413);
or UO_1915 (O_1915,N_23930,N_23918);
and UO_1916 (O_1916,N_24402,N_24153);
and UO_1917 (O_1917,N_24533,N_24038);
nand UO_1918 (O_1918,N_24652,N_24733);
nand UO_1919 (O_1919,N_23870,N_24287);
xnor UO_1920 (O_1920,N_24392,N_23784);
and UO_1921 (O_1921,N_24836,N_24615);
or UO_1922 (O_1922,N_24199,N_23968);
and UO_1923 (O_1923,N_24377,N_24893);
or UO_1924 (O_1924,N_24079,N_23935);
nand UO_1925 (O_1925,N_24418,N_24092);
nand UO_1926 (O_1926,N_24499,N_24097);
nor UO_1927 (O_1927,N_24563,N_24000);
nand UO_1928 (O_1928,N_24167,N_24692);
and UO_1929 (O_1929,N_24644,N_24112);
xnor UO_1930 (O_1930,N_24970,N_24352);
or UO_1931 (O_1931,N_24271,N_24333);
nor UO_1932 (O_1932,N_24746,N_24658);
nor UO_1933 (O_1933,N_24422,N_23760);
xnor UO_1934 (O_1934,N_24099,N_24692);
nand UO_1935 (O_1935,N_24973,N_24924);
nor UO_1936 (O_1936,N_23758,N_24540);
nand UO_1937 (O_1937,N_24159,N_23982);
or UO_1938 (O_1938,N_24378,N_23926);
nand UO_1939 (O_1939,N_24036,N_24654);
and UO_1940 (O_1940,N_23763,N_23883);
and UO_1941 (O_1941,N_24039,N_24617);
nand UO_1942 (O_1942,N_24326,N_24383);
and UO_1943 (O_1943,N_24601,N_24377);
nor UO_1944 (O_1944,N_24991,N_24948);
nor UO_1945 (O_1945,N_24486,N_24280);
nor UO_1946 (O_1946,N_24915,N_24743);
nand UO_1947 (O_1947,N_24691,N_24591);
nor UO_1948 (O_1948,N_24488,N_24189);
nor UO_1949 (O_1949,N_24415,N_24950);
and UO_1950 (O_1950,N_23769,N_24583);
xor UO_1951 (O_1951,N_24053,N_24279);
nor UO_1952 (O_1952,N_24439,N_24667);
and UO_1953 (O_1953,N_24906,N_23882);
nand UO_1954 (O_1954,N_24555,N_24227);
nor UO_1955 (O_1955,N_24763,N_24253);
and UO_1956 (O_1956,N_24623,N_24641);
nor UO_1957 (O_1957,N_24773,N_24271);
nand UO_1958 (O_1958,N_24682,N_24090);
nand UO_1959 (O_1959,N_24096,N_24319);
nor UO_1960 (O_1960,N_23915,N_23780);
nand UO_1961 (O_1961,N_24870,N_24798);
and UO_1962 (O_1962,N_24739,N_23855);
nor UO_1963 (O_1963,N_24429,N_24556);
nand UO_1964 (O_1964,N_24660,N_24986);
or UO_1965 (O_1965,N_24816,N_24363);
and UO_1966 (O_1966,N_24124,N_23761);
and UO_1967 (O_1967,N_23982,N_24160);
and UO_1968 (O_1968,N_24682,N_24127);
or UO_1969 (O_1969,N_24826,N_24616);
nand UO_1970 (O_1970,N_24484,N_24468);
or UO_1971 (O_1971,N_24784,N_24152);
and UO_1972 (O_1972,N_24382,N_24856);
and UO_1973 (O_1973,N_23970,N_23786);
nor UO_1974 (O_1974,N_23988,N_24347);
or UO_1975 (O_1975,N_24481,N_24394);
and UO_1976 (O_1976,N_24862,N_24234);
xor UO_1977 (O_1977,N_24574,N_23892);
nor UO_1978 (O_1978,N_23776,N_24109);
nand UO_1979 (O_1979,N_24373,N_23875);
nand UO_1980 (O_1980,N_24979,N_23817);
and UO_1981 (O_1981,N_24186,N_24965);
or UO_1982 (O_1982,N_24034,N_23943);
and UO_1983 (O_1983,N_24428,N_23951);
xnor UO_1984 (O_1984,N_24458,N_24840);
nor UO_1985 (O_1985,N_24825,N_24244);
nor UO_1986 (O_1986,N_24965,N_24983);
nand UO_1987 (O_1987,N_24535,N_24348);
or UO_1988 (O_1988,N_24561,N_24761);
xor UO_1989 (O_1989,N_23924,N_24581);
xnor UO_1990 (O_1990,N_24812,N_24539);
or UO_1991 (O_1991,N_23794,N_24352);
nor UO_1992 (O_1992,N_23812,N_24871);
nor UO_1993 (O_1993,N_24850,N_23938);
or UO_1994 (O_1994,N_24576,N_24612);
xnor UO_1995 (O_1995,N_23957,N_24060);
nand UO_1996 (O_1996,N_24096,N_23930);
nor UO_1997 (O_1997,N_24336,N_24525);
nor UO_1998 (O_1998,N_24342,N_24865);
xnor UO_1999 (O_1999,N_24201,N_23923);
and UO_2000 (O_2000,N_24270,N_24086);
or UO_2001 (O_2001,N_23958,N_24431);
xnor UO_2002 (O_2002,N_24224,N_24151);
xor UO_2003 (O_2003,N_24222,N_24049);
nor UO_2004 (O_2004,N_24838,N_24298);
or UO_2005 (O_2005,N_24910,N_24763);
and UO_2006 (O_2006,N_23856,N_23800);
xor UO_2007 (O_2007,N_24596,N_24584);
xnor UO_2008 (O_2008,N_24288,N_24864);
nand UO_2009 (O_2009,N_24922,N_23769);
or UO_2010 (O_2010,N_24879,N_24412);
xor UO_2011 (O_2011,N_24566,N_24853);
nor UO_2012 (O_2012,N_24483,N_24602);
or UO_2013 (O_2013,N_23999,N_23918);
nand UO_2014 (O_2014,N_24335,N_23843);
xnor UO_2015 (O_2015,N_24607,N_23762);
nor UO_2016 (O_2016,N_24271,N_23930);
nor UO_2017 (O_2017,N_23865,N_24367);
and UO_2018 (O_2018,N_23917,N_24819);
and UO_2019 (O_2019,N_23865,N_24819);
and UO_2020 (O_2020,N_24312,N_24738);
xnor UO_2021 (O_2021,N_24690,N_24472);
xnor UO_2022 (O_2022,N_24252,N_24111);
xor UO_2023 (O_2023,N_24537,N_24476);
and UO_2024 (O_2024,N_24213,N_24329);
nor UO_2025 (O_2025,N_23861,N_24901);
xnor UO_2026 (O_2026,N_24725,N_24924);
and UO_2027 (O_2027,N_24604,N_24785);
xor UO_2028 (O_2028,N_24139,N_23951);
xnor UO_2029 (O_2029,N_24016,N_23964);
or UO_2030 (O_2030,N_24869,N_24091);
nand UO_2031 (O_2031,N_24084,N_23861);
nand UO_2032 (O_2032,N_24657,N_24587);
nand UO_2033 (O_2033,N_24340,N_24189);
nor UO_2034 (O_2034,N_24908,N_24627);
xor UO_2035 (O_2035,N_24074,N_24314);
or UO_2036 (O_2036,N_24312,N_24411);
or UO_2037 (O_2037,N_24367,N_24634);
and UO_2038 (O_2038,N_24749,N_24304);
and UO_2039 (O_2039,N_23924,N_24847);
nor UO_2040 (O_2040,N_23892,N_24794);
nand UO_2041 (O_2041,N_24301,N_23757);
nand UO_2042 (O_2042,N_24998,N_24025);
nor UO_2043 (O_2043,N_24598,N_24545);
nor UO_2044 (O_2044,N_24443,N_23809);
or UO_2045 (O_2045,N_23918,N_23798);
and UO_2046 (O_2046,N_24067,N_24105);
xor UO_2047 (O_2047,N_24512,N_23944);
nor UO_2048 (O_2048,N_24606,N_24688);
or UO_2049 (O_2049,N_24330,N_23871);
xnor UO_2050 (O_2050,N_24403,N_23802);
or UO_2051 (O_2051,N_24841,N_24631);
nor UO_2052 (O_2052,N_23994,N_24940);
nor UO_2053 (O_2053,N_24254,N_23943);
or UO_2054 (O_2054,N_23990,N_24619);
xnor UO_2055 (O_2055,N_24148,N_24639);
xnor UO_2056 (O_2056,N_24563,N_24728);
and UO_2057 (O_2057,N_24535,N_24328);
and UO_2058 (O_2058,N_24404,N_24704);
xor UO_2059 (O_2059,N_24806,N_23900);
xnor UO_2060 (O_2060,N_24653,N_24951);
and UO_2061 (O_2061,N_24849,N_24365);
nand UO_2062 (O_2062,N_24602,N_24203);
xnor UO_2063 (O_2063,N_24576,N_23844);
or UO_2064 (O_2064,N_24917,N_23766);
and UO_2065 (O_2065,N_24545,N_24029);
or UO_2066 (O_2066,N_24362,N_24222);
nand UO_2067 (O_2067,N_23923,N_23762);
or UO_2068 (O_2068,N_24428,N_24094);
nor UO_2069 (O_2069,N_23942,N_23851);
xnor UO_2070 (O_2070,N_24611,N_23965);
nand UO_2071 (O_2071,N_24368,N_24710);
and UO_2072 (O_2072,N_24265,N_23923);
or UO_2073 (O_2073,N_23866,N_24793);
nand UO_2074 (O_2074,N_24137,N_23881);
nor UO_2075 (O_2075,N_24435,N_24566);
nor UO_2076 (O_2076,N_23870,N_23761);
and UO_2077 (O_2077,N_24577,N_24857);
nand UO_2078 (O_2078,N_24090,N_24314);
and UO_2079 (O_2079,N_24934,N_24629);
xor UO_2080 (O_2080,N_23976,N_24503);
or UO_2081 (O_2081,N_24928,N_24792);
nand UO_2082 (O_2082,N_24836,N_23935);
nand UO_2083 (O_2083,N_23889,N_23879);
nor UO_2084 (O_2084,N_24109,N_24936);
nand UO_2085 (O_2085,N_23961,N_24793);
nand UO_2086 (O_2086,N_24158,N_24272);
and UO_2087 (O_2087,N_23988,N_24188);
and UO_2088 (O_2088,N_24840,N_24558);
and UO_2089 (O_2089,N_24339,N_23791);
xor UO_2090 (O_2090,N_24254,N_24359);
nand UO_2091 (O_2091,N_24254,N_24978);
or UO_2092 (O_2092,N_24934,N_23981);
xor UO_2093 (O_2093,N_24743,N_23987);
and UO_2094 (O_2094,N_24200,N_23999);
xnor UO_2095 (O_2095,N_24179,N_24824);
or UO_2096 (O_2096,N_24930,N_24565);
and UO_2097 (O_2097,N_24972,N_24448);
and UO_2098 (O_2098,N_23914,N_24501);
xor UO_2099 (O_2099,N_23853,N_24735);
nand UO_2100 (O_2100,N_24822,N_23812);
nor UO_2101 (O_2101,N_24914,N_24096);
and UO_2102 (O_2102,N_24473,N_24658);
nor UO_2103 (O_2103,N_24652,N_24033);
nor UO_2104 (O_2104,N_23782,N_24148);
or UO_2105 (O_2105,N_24770,N_24078);
xor UO_2106 (O_2106,N_23965,N_24708);
or UO_2107 (O_2107,N_23919,N_24217);
nand UO_2108 (O_2108,N_23844,N_23777);
nand UO_2109 (O_2109,N_24797,N_24740);
and UO_2110 (O_2110,N_24110,N_24916);
xor UO_2111 (O_2111,N_24352,N_24886);
and UO_2112 (O_2112,N_24086,N_24667);
or UO_2113 (O_2113,N_24770,N_24906);
xnor UO_2114 (O_2114,N_24000,N_24401);
xnor UO_2115 (O_2115,N_24088,N_24572);
xor UO_2116 (O_2116,N_24860,N_24864);
or UO_2117 (O_2117,N_24960,N_24384);
xnor UO_2118 (O_2118,N_23938,N_23805);
and UO_2119 (O_2119,N_24190,N_24926);
nand UO_2120 (O_2120,N_24839,N_24059);
nand UO_2121 (O_2121,N_24604,N_24117);
and UO_2122 (O_2122,N_23887,N_24044);
nor UO_2123 (O_2123,N_24594,N_24783);
nor UO_2124 (O_2124,N_24215,N_24410);
or UO_2125 (O_2125,N_23776,N_24380);
or UO_2126 (O_2126,N_24809,N_24912);
nor UO_2127 (O_2127,N_24459,N_23898);
nor UO_2128 (O_2128,N_24685,N_23774);
or UO_2129 (O_2129,N_24052,N_24572);
or UO_2130 (O_2130,N_24202,N_24748);
nand UO_2131 (O_2131,N_24290,N_24839);
xor UO_2132 (O_2132,N_23787,N_23879);
xor UO_2133 (O_2133,N_24153,N_24852);
nor UO_2134 (O_2134,N_24875,N_24289);
or UO_2135 (O_2135,N_24765,N_23911);
nand UO_2136 (O_2136,N_24679,N_23988);
or UO_2137 (O_2137,N_23936,N_24288);
nand UO_2138 (O_2138,N_24193,N_23932);
and UO_2139 (O_2139,N_23884,N_24419);
xnor UO_2140 (O_2140,N_24814,N_24964);
nand UO_2141 (O_2141,N_23881,N_24332);
and UO_2142 (O_2142,N_24840,N_24742);
and UO_2143 (O_2143,N_24388,N_24221);
xnor UO_2144 (O_2144,N_24946,N_24410);
nand UO_2145 (O_2145,N_24127,N_24561);
xnor UO_2146 (O_2146,N_24112,N_23887);
or UO_2147 (O_2147,N_24837,N_24329);
nand UO_2148 (O_2148,N_24527,N_23799);
or UO_2149 (O_2149,N_23874,N_24810);
nand UO_2150 (O_2150,N_24270,N_24847);
and UO_2151 (O_2151,N_23951,N_24119);
or UO_2152 (O_2152,N_23908,N_24313);
nor UO_2153 (O_2153,N_24067,N_24150);
and UO_2154 (O_2154,N_24768,N_24195);
nand UO_2155 (O_2155,N_23766,N_24932);
and UO_2156 (O_2156,N_24705,N_23846);
xnor UO_2157 (O_2157,N_23932,N_24492);
xnor UO_2158 (O_2158,N_24096,N_24122);
or UO_2159 (O_2159,N_24339,N_23799);
nor UO_2160 (O_2160,N_23840,N_24103);
nand UO_2161 (O_2161,N_24695,N_24809);
xor UO_2162 (O_2162,N_23942,N_24613);
xor UO_2163 (O_2163,N_24222,N_24653);
nand UO_2164 (O_2164,N_24214,N_24023);
and UO_2165 (O_2165,N_23932,N_24034);
xnor UO_2166 (O_2166,N_24143,N_24144);
nand UO_2167 (O_2167,N_24771,N_24319);
xor UO_2168 (O_2168,N_24213,N_24591);
nor UO_2169 (O_2169,N_24867,N_24493);
or UO_2170 (O_2170,N_24369,N_24719);
xnor UO_2171 (O_2171,N_23896,N_24174);
nand UO_2172 (O_2172,N_24931,N_24916);
nand UO_2173 (O_2173,N_24694,N_23888);
and UO_2174 (O_2174,N_24146,N_24854);
nand UO_2175 (O_2175,N_24866,N_24458);
nor UO_2176 (O_2176,N_23752,N_24405);
or UO_2177 (O_2177,N_23884,N_24863);
nand UO_2178 (O_2178,N_24849,N_24256);
or UO_2179 (O_2179,N_24975,N_23925);
nor UO_2180 (O_2180,N_24021,N_24160);
nor UO_2181 (O_2181,N_23887,N_24805);
and UO_2182 (O_2182,N_24771,N_24357);
xor UO_2183 (O_2183,N_24488,N_24685);
or UO_2184 (O_2184,N_24394,N_24316);
or UO_2185 (O_2185,N_24857,N_24838);
nand UO_2186 (O_2186,N_23812,N_23912);
xor UO_2187 (O_2187,N_23817,N_24863);
nand UO_2188 (O_2188,N_23977,N_24845);
and UO_2189 (O_2189,N_24625,N_24461);
or UO_2190 (O_2190,N_24354,N_24317);
and UO_2191 (O_2191,N_24837,N_23827);
nand UO_2192 (O_2192,N_24682,N_23927);
xnor UO_2193 (O_2193,N_24766,N_24066);
or UO_2194 (O_2194,N_24788,N_23956);
and UO_2195 (O_2195,N_23854,N_24168);
xor UO_2196 (O_2196,N_24878,N_24763);
xnor UO_2197 (O_2197,N_24028,N_24603);
nand UO_2198 (O_2198,N_23984,N_23787);
and UO_2199 (O_2199,N_24323,N_23830);
and UO_2200 (O_2200,N_24079,N_24374);
xnor UO_2201 (O_2201,N_23914,N_24149);
and UO_2202 (O_2202,N_23905,N_24723);
and UO_2203 (O_2203,N_24871,N_24625);
nand UO_2204 (O_2204,N_24234,N_24127);
xnor UO_2205 (O_2205,N_24325,N_24111);
or UO_2206 (O_2206,N_24322,N_24402);
xor UO_2207 (O_2207,N_24437,N_24273);
nand UO_2208 (O_2208,N_24169,N_24399);
or UO_2209 (O_2209,N_23924,N_24347);
or UO_2210 (O_2210,N_23907,N_23976);
nand UO_2211 (O_2211,N_24396,N_24291);
or UO_2212 (O_2212,N_23934,N_24133);
or UO_2213 (O_2213,N_24407,N_24583);
and UO_2214 (O_2214,N_24090,N_24249);
nand UO_2215 (O_2215,N_23867,N_24038);
nor UO_2216 (O_2216,N_24233,N_24138);
nand UO_2217 (O_2217,N_24150,N_23795);
and UO_2218 (O_2218,N_23814,N_23853);
xor UO_2219 (O_2219,N_24525,N_24865);
or UO_2220 (O_2220,N_23752,N_23833);
nor UO_2221 (O_2221,N_24712,N_24071);
and UO_2222 (O_2222,N_24017,N_24688);
and UO_2223 (O_2223,N_24209,N_24058);
nand UO_2224 (O_2224,N_24255,N_23844);
nor UO_2225 (O_2225,N_24892,N_24855);
or UO_2226 (O_2226,N_24335,N_24447);
or UO_2227 (O_2227,N_23902,N_24543);
or UO_2228 (O_2228,N_23878,N_23967);
xor UO_2229 (O_2229,N_24800,N_24216);
nand UO_2230 (O_2230,N_24235,N_24565);
nand UO_2231 (O_2231,N_24122,N_23854);
nand UO_2232 (O_2232,N_24472,N_24190);
and UO_2233 (O_2233,N_23877,N_24131);
nand UO_2234 (O_2234,N_24909,N_23928);
nand UO_2235 (O_2235,N_24934,N_24947);
xnor UO_2236 (O_2236,N_24583,N_24832);
or UO_2237 (O_2237,N_23957,N_23770);
or UO_2238 (O_2238,N_24501,N_24710);
and UO_2239 (O_2239,N_24092,N_24023);
xor UO_2240 (O_2240,N_24713,N_24249);
xor UO_2241 (O_2241,N_24453,N_24964);
xnor UO_2242 (O_2242,N_23882,N_24513);
and UO_2243 (O_2243,N_24751,N_24504);
xnor UO_2244 (O_2244,N_24701,N_24003);
or UO_2245 (O_2245,N_23972,N_24021);
xnor UO_2246 (O_2246,N_24427,N_24806);
and UO_2247 (O_2247,N_24955,N_23840);
nor UO_2248 (O_2248,N_24067,N_24899);
nor UO_2249 (O_2249,N_23905,N_24914);
xnor UO_2250 (O_2250,N_24302,N_24276);
nor UO_2251 (O_2251,N_24601,N_23951);
nand UO_2252 (O_2252,N_24815,N_24489);
and UO_2253 (O_2253,N_23941,N_23751);
and UO_2254 (O_2254,N_23753,N_23763);
nor UO_2255 (O_2255,N_24435,N_24318);
and UO_2256 (O_2256,N_24841,N_24866);
nor UO_2257 (O_2257,N_24835,N_24774);
nand UO_2258 (O_2258,N_24164,N_24083);
and UO_2259 (O_2259,N_23967,N_24442);
xor UO_2260 (O_2260,N_24001,N_24205);
nand UO_2261 (O_2261,N_24834,N_24240);
or UO_2262 (O_2262,N_24501,N_23910);
and UO_2263 (O_2263,N_24436,N_24654);
nand UO_2264 (O_2264,N_23785,N_24405);
or UO_2265 (O_2265,N_24080,N_23774);
nand UO_2266 (O_2266,N_24726,N_24478);
or UO_2267 (O_2267,N_24905,N_24594);
or UO_2268 (O_2268,N_24877,N_23987);
or UO_2269 (O_2269,N_24900,N_24189);
nor UO_2270 (O_2270,N_24292,N_24295);
or UO_2271 (O_2271,N_24419,N_24176);
or UO_2272 (O_2272,N_24878,N_24622);
nand UO_2273 (O_2273,N_24591,N_24935);
nand UO_2274 (O_2274,N_23940,N_24004);
nand UO_2275 (O_2275,N_24658,N_24284);
and UO_2276 (O_2276,N_23853,N_24849);
nor UO_2277 (O_2277,N_24213,N_24630);
xor UO_2278 (O_2278,N_24856,N_24096);
nor UO_2279 (O_2279,N_24488,N_23836);
nand UO_2280 (O_2280,N_24464,N_24990);
nand UO_2281 (O_2281,N_24317,N_23952);
nor UO_2282 (O_2282,N_23849,N_24043);
or UO_2283 (O_2283,N_24055,N_24571);
xor UO_2284 (O_2284,N_24897,N_24627);
xor UO_2285 (O_2285,N_24973,N_23981);
and UO_2286 (O_2286,N_24266,N_24792);
or UO_2287 (O_2287,N_23875,N_24950);
xnor UO_2288 (O_2288,N_24332,N_24956);
or UO_2289 (O_2289,N_23999,N_24075);
or UO_2290 (O_2290,N_24673,N_23805);
nand UO_2291 (O_2291,N_23808,N_24948);
nor UO_2292 (O_2292,N_24625,N_24620);
and UO_2293 (O_2293,N_24332,N_24682);
and UO_2294 (O_2294,N_24550,N_24146);
xor UO_2295 (O_2295,N_23899,N_24583);
or UO_2296 (O_2296,N_24091,N_24134);
xnor UO_2297 (O_2297,N_24320,N_24548);
or UO_2298 (O_2298,N_24293,N_24412);
nor UO_2299 (O_2299,N_24126,N_23823);
nand UO_2300 (O_2300,N_24013,N_24512);
and UO_2301 (O_2301,N_24766,N_24134);
nor UO_2302 (O_2302,N_24332,N_24262);
and UO_2303 (O_2303,N_24267,N_24780);
xor UO_2304 (O_2304,N_24493,N_24298);
or UO_2305 (O_2305,N_24567,N_23996);
and UO_2306 (O_2306,N_24759,N_23973);
nor UO_2307 (O_2307,N_24214,N_24002);
nand UO_2308 (O_2308,N_24325,N_24258);
xor UO_2309 (O_2309,N_23874,N_24968);
xnor UO_2310 (O_2310,N_24018,N_24528);
xor UO_2311 (O_2311,N_24408,N_24527);
xor UO_2312 (O_2312,N_23908,N_24648);
nand UO_2313 (O_2313,N_24399,N_24739);
and UO_2314 (O_2314,N_24433,N_24975);
and UO_2315 (O_2315,N_23760,N_24692);
xnor UO_2316 (O_2316,N_24642,N_23822);
xor UO_2317 (O_2317,N_24439,N_24361);
and UO_2318 (O_2318,N_24848,N_24040);
nor UO_2319 (O_2319,N_24024,N_24918);
nor UO_2320 (O_2320,N_23992,N_24545);
and UO_2321 (O_2321,N_23853,N_24341);
nand UO_2322 (O_2322,N_23961,N_24163);
nor UO_2323 (O_2323,N_24730,N_24950);
nand UO_2324 (O_2324,N_24318,N_24999);
or UO_2325 (O_2325,N_24416,N_24770);
xor UO_2326 (O_2326,N_24047,N_24706);
or UO_2327 (O_2327,N_24491,N_24033);
nand UO_2328 (O_2328,N_24528,N_23848);
and UO_2329 (O_2329,N_24511,N_24990);
nor UO_2330 (O_2330,N_24184,N_24690);
nand UO_2331 (O_2331,N_24798,N_24572);
xnor UO_2332 (O_2332,N_23869,N_24077);
and UO_2333 (O_2333,N_24282,N_24021);
and UO_2334 (O_2334,N_24230,N_24919);
or UO_2335 (O_2335,N_24350,N_23923);
or UO_2336 (O_2336,N_24213,N_24515);
or UO_2337 (O_2337,N_24774,N_23909);
and UO_2338 (O_2338,N_24973,N_24611);
or UO_2339 (O_2339,N_24040,N_24870);
or UO_2340 (O_2340,N_24104,N_24894);
and UO_2341 (O_2341,N_24130,N_23836);
nand UO_2342 (O_2342,N_24575,N_24811);
xor UO_2343 (O_2343,N_23879,N_24858);
xnor UO_2344 (O_2344,N_24669,N_24578);
or UO_2345 (O_2345,N_24920,N_24137);
xor UO_2346 (O_2346,N_24417,N_23761);
xor UO_2347 (O_2347,N_24486,N_24378);
nand UO_2348 (O_2348,N_24058,N_24659);
nor UO_2349 (O_2349,N_24575,N_23948);
xnor UO_2350 (O_2350,N_24616,N_23859);
or UO_2351 (O_2351,N_23873,N_24965);
and UO_2352 (O_2352,N_24029,N_24330);
or UO_2353 (O_2353,N_23882,N_24870);
nand UO_2354 (O_2354,N_23956,N_24903);
xor UO_2355 (O_2355,N_24223,N_24636);
nor UO_2356 (O_2356,N_24698,N_24794);
xor UO_2357 (O_2357,N_24886,N_24465);
nor UO_2358 (O_2358,N_23936,N_24176);
xor UO_2359 (O_2359,N_23948,N_24638);
xnor UO_2360 (O_2360,N_24566,N_23806);
nand UO_2361 (O_2361,N_24830,N_24398);
nand UO_2362 (O_2362,N_24512,N_23873);
nand UO_2363 (O_2363,N_23922,N_24113);
nor UO_2364 (O_2364,N_24872,N_23914);
or UO_2365 (O_2365,N_24611,N_24972);
and UO_2366 (O_2366,N_24113,N_24513);
nand UO_2367 (O_2367,N_24547,N_24724);
xnor UO_2368 (O_2368,N_23871,N_24037);
or UO_2369 (O_2369,N_24747,N_24082);
xnor UO_2370 (O_2370,N_23860,N_24193);
nand UO_2371 (O_2371,N_24933,N_24279);
and UO_2372 (O_2372,N_23820,N_24108);
nand UO_2373 (O_2373,N_23879,N_24302);
and UO_2374 (O_2374,N_23756,N_24070);
or UO_2375 (O_2375,N_23784,N_24819);
nor UO_2376 (O_2376,N_23795,N_23898);
nand UO_2377 (O_2377,N_24614,N_24186);
xor UO_2378 (O_2378,N_23795,N_24239);
nor UO_2379 (O_2379,N_23946,N_24652);
or UO_2380 (O_2380,N_24664,N_24608);
nor UO_2381 (O_2381,N_24977,N_24175);
and UO_2382 (O_2382,N_24022,N_24498);
nand UO_2383 (O_2383,N_24457,N_24118);
or UO_2384 (O_2384,N_24379,N_24331);
nand UO_2385 (O_2385,N_24228,N_24893);
or UO_2386 (O_2386,N_24188,N_24750);
nor UO_2387 (O_2387,N_24435,N_24414);
nand UO_2388 (O_2388,N_24916,N_24671);
nand UO_2389 (O_2389,N_24051,N_24642);
or UO_2390 (O_2390,N_24902,N_24553);
nor UO_2391 (O_2391,N_24642,N_24049);
xor UO_2392 (O_2392,N_23850,N_24939);
nor UO_2393 (O_2393,N_24238,N_23932);
xor UO_2394 (O_2394,N_24081,N_24244);
nand UO_2395 (O_2395,N_23881,N_23782);
and UO_2396 (O_2396,N_24924,N_24544);
xor UO_2397 (O_2397,N_24612,N_24080);
nand UO_2398 (O_2398,N_23840,N_24030);
xor UO_2399 (O_2399,N_24536,N_24808);
nor UO_2400 (O_2400,N_24836,N_23900);
xnor UO_2401 (O_2401,N_24280,N_24620);
nand UO_2402 (O_2402,N_24611,N_24579);
nand UO_2403 (O_2403,N_24826,N_24202);
xnor UO_2404 (O_2404,N_24785,N_23757);
xnor UO_2405 (O_2405,N_24052,N_24295);
or UO_2406 (O_2406,N_23845,N_24219);
and UO_2407 (O_2407,N_24767,N_24459);
nor UO_2408 (O_2408,N_24558,N_23882);
and UO_2409 (O_2409,N_23872,N_24803);
and UO_2410 (O_2410,N_24774,N_23897);
nor UO_2411 (O_2411,N_24077,N_24079);
nand UO_2412 (O_2412,N_24445,N_23905);
or UO_2413 (O_2413,N_24708,N_23755);
nor UO_2414 (O_2414,N_24085,N_24169);
nor UO_2415 (O_2415,N_24291,N_24765);
nand UO_2416 (O_2416,N_23753,N_24441);
and UO_2417 (O_2417,N_24194,N_23992);
or UO_2418 (O_2418,N_23806,N_24037);
nor UO_2419 (O_2419,N_24094,N_23805);
or UO_2420 (O_2420,N_24886,N_23914);
nand UO_2421 (O_2421,N_24942,N_24525);
xnor UO_2422 (O_2422,N_24015,N_24585);
nor UO_2423 (O_2423,N_24048,N_24010);
or UO_2424 (O_2424,N_24319,N_24302);
and UO_2425 (O_2425,N_24215,N_23893);
or UO_2426 (O_2426,N_24167,N_23862);
xor UO_2427 (O_2427,N_23817,N_23996);
xor UO_2428 (O_2428,N_24135,N_23825);
xor UO_2429 (O_2429,N_24621,N_23975);
and UO_2430 (O_2430,N_24608,N_24579);
and UO_2431 (O_2431,N_23876,N_23976);
nand UO_2432 (O_2432,N_24162,N_24279);
nor UO_2433 (O_2433,N_24993,N_24750);
nand UO_2434 (O_2434,N_24662,N_24093);
nor UO_2435 (O_2435,N_24456,N_23779);
and UO_2436 (O_2436,N_24239,N_24087);
xor UO_2437 (O_2437,N_24083,N_24249);
nor UO_2438 (O_2438,N_23817,N_24109);
xnor UO_2439 (O_2439,N_24825,N_23910);
nor UO_2440 (O_2440,N_24125,N_24676);
nand UO_2441 (O_2441,N_24265,N_23972);
nor UO_2442 (O_2442,N_24670,N_24749);
nor UO_2443 (O_2443,N_24842,N_24752);
and UO_2444 (O_2444,N_24692,N_24805);
and UO_2445 (O_2445,N_24859,N_24545);
nand UO_2446 (O_2446,N_24646,N_24622);
nand UO_2447 (O_2447,N_24483,N_23814);
xnor UO_2448 (O_2448,N_24722,N_24177);
and UO_2449 (O_2449,N_24864,N_24758);
or UO_2450 (O_2450,N_23902,N_24089);
nand UO_2451 (O_2451,N_23956,N_23848);
and UO_2452 (O_2452,N_24408,N_24656);
or UO_2453 (O_2453,N_24730,N_23793);
or UO_2454 (O_2454,N_23937,N_24407);
and UO_2455 (O_2455,N_24269,N_24843);
xor UO_2456 (O_2456,N_24223,N_24092);
nand UO_2457 (O_2457,N_24218,N_24761);
xnor UO_2458 (O_2458,N_24262,N_24373);
nand UO_2459 (O_2459,N_24514,N_23970);
nand UO_2460 (O_2460,N_24655,N_24203);
xnor UO_2461 (O_2461,N_24702,N_23834);
nor UO_2462 (O_2462,N_24730,N_24569);
nor UO_2463 (O_2463,N_24164,N_24156);
nand UO_2464 (O_2464,N_24908,N_24051);
nor UO_2465 (O_2465,N_23967,N_23938);
nor UO_2466 (O_2466,N_23760,N_24889);
nor UO_2467 (O_2467,N_23919,N_23789);
nand UO_2468 (O_2468,N_24037,N_24051);
or UO_2469 (O_2469,N_24170,N_23977);
and UO_2470 (O_2470,N_24279,N_24211);
and UO_2471 (O_2471,N_24835,N_24048);
and UO_2472 (O_2472,N_23813,N_24765);
or UO_2473 (O_2473,N_24189,N_23810);
xnor UO_2474 (O_2474,N_24095,N_24655);
xnor UO_2475 (O_2475,N_24331,N_24656);
and UO_2476 (O_2476,N_24456,N_24767);
xor UO_2477 (O_2477,N_23896,N_24013);
or UO_2478 (O_2478,N_24060,N_24218);
nor UO_2479 (O_2479,N_24712,N_24093);
xor UO_2480 (O_2480,N_24820,N_24367);
and UO_2481 (O_2481,N_23811,N_24706);
and UO_2482 (O_2482,N_23986,N_24872);
xor UO_2483 (O_2483,N_24681,N_24179);
and UO_2484 (O_2484,N_24204,N_24086);
nand UO_2485 (O_2485,N_24187,N_24213);
xor UO_2486 (O_2486,N_23785,N_24757);
nor UO_2487 (O_2487,N_24034,N_24579);
and UO_2488 (O_2488,N_24187,N_24548);
nand UO_2489 (O_2489,N_24711,N_24678);
nor UO_2490 (O_2490,N_24477,N_24529);
nor UO_2491 (O_2491,N_24109,N_24204);
nand UO_2492 (O_2492,N_24701,N_24310);
or UO_2493 (O_2493,N_23985,N_24378);
or UO_2494 (O_2494,N_24203,N_24894);
and UO_2495 (O_2495,N_24892,N_24513);
or UO_2496 (O_2496,N_24053,N_24540);
nor UO_2497 (O_2497,N_23832,N_24536);
nor UO_2498 (O_2498,N_23790,N_24819);
xnor UO_2499 (O_2499,N_24539,N_23807);
or UO_2500 (O_2500,N_24628,N_24608);
nand UO_2501 (O_2501,N_23756,N_24819);
xor UO_2502 (O_2502,N_24784,N_24606);
nor UO_2503 (O_2503,N_23825,N_24759);
and UO_2504 (O_2504,N_24070,N_24775);
and UO_2505 (O_2505,N_24019,N_23876);
or UO_2506 (O_2506,N_24473,N_24264);
and UO_2507 (O_2507,N_24612,N_24258);
and UO_2508 (O_2508,N_24308,N_24171);
nor UO_2509 (O_2509,N_24886,N_24871);
nand UO_2510 (O_2510,N_24198,N_23858);
or UO_2511 (O_2511,N_24055,N_24400);
xor UO_2512 (O_2512,N_24427,N_24008);
or UO_2513 (O_2513,N_23760,N_24931);
or UO_2514 (O_2514,N_24384,N_24895);
or UO_2515 (O_2515,N_24236,N_24012);
xor UO_2516 (O_2516,N_24702,N_24671);
nor UO_2517 (O_2517,N_24787,N_24515);
xor UO_2518 (O_2518,N_23858,N_24386);
and UO_2519 (O_2519,N_23916,N_24354);
and UO_2520 (O_2520,N_24856,N_24407);
xor UO_2521 (O_2521,N_24199,N_23846);
or UO_2522 (O_2522,N_24871,N_24033);
or UO_2523 (O_2523,N_24830,N_24402);
and UO_2524 (O_2524,N_24663,N_24468);
or UO_2525 (O_2525,N_24484,N_24861);
nand UO_2526 (O_2526,N_24127,N_23930);
or UO_2527 (O_2527,N_24613,N_24631);
or UO_2528 (O_2528,N_24989,N_24597);
and UO_2529 (O_2529,N_24207,N_24303);
xor UO_2530 (O_2530,N_24624,N_24320);
nor UO_2531 (O_2531,N_23919,N_24651);
and UO_2532 (O_2532,N_24298,N_24712);
or UO_2533 (O_2533,N_24588,N_24502);
xnor UO_2534 (O_2534,N_24167,N_24584);
and UO_2535 (O_2535,N_24281,N_24790);
nor UO_2536 (O_2536,N_23762,N_24388);
and UO_2537 (O_2537,N_24858,N_24962);
xor UO_2538 (O_2538,N_24273,N_24704);
nand UO_2539 (O_2539,N_24418,N_24242);
nor UO_2540 (O_2540,N_24244,N_24363);
nand UO_2541 (O_2541,N_24430,N_23844);
nand UO_2542 (O_2542,N_24930,N_24230);
xor UO_2543 (O_2543,N_24593,N_23836);
nand UO_2544 (O_2544,N_24060,N_24360);
or UO_2545 (O_2545,N_24334,N_24028);
or UO_2546 (O_2546,N_23959,N_24223);
xnor UO_2547 (O_2547,N_24446,N_24356);
nand UO_2548 (O_2548,N_24762,N_24825);
xor UO_2549 (O_2549,N_23877,N_24203);
nand UO_2550 (O_2550,N_23789,N_23821);
nor UO_2551 (O_2551,N_24163,N_23904);
nand UO_2552 (O_2552,N_24196,N_23914);
xnor UO_2553 (O_2553,N_24691,N_23882);
and UO_2554 (O_2554,N_24469,N_24458);
nand UO_2555 (O_2555,N_23794,N_24630);
xnor UO_2556 (O_2556,N_24080,N_24749);
and UO_2557 (O_2557,N_24215,N_23889);
or UO_2558 (O_2558,N_24066,N_24549);
nor UO_2559 (O_2559,N_23990,N_24022);
nor UO_2560 (O_2560,N_24515,N_24512);
xnor UO_2561 (O_2561,N_24511,N_24938);
or UO_2562 (O_2562,N_24509,N_24138);
nand UO_2563 (O_2563,N_23862,N_24905);
xor UO_2564 (O_2564,N_23958,N_23756);
or UO_2565 (O_2565,N_24307,N_24736);
or UO_2566 (O_2566,N_24688,N_24801);
nor UO_2567 (O_2567,N_24782,N_23750);
xor UO_2568 (O_2568,N_24499,N_24310);
nand UO_2569 (O_2569,N_24939,N_24832);
or UO_2570 (O_2570,N_23777,N_24023);
nand UO_2571 (O_2571,N_24506,N_24129);
and UO_2572 (O_2572,N_24452,N_24149);
nand UO_2573 (O_2573,N_24409,N_23866);
or UO_2574 (O_2574,N_24153,N_24550);
nand UO_2575 (O_2575,N_24395,N_24501);
or UO_2576 (O_2576,N_24198,N_24984);
xor UO_2577 (O_2577,N_24335,N_24407);
nor UO_2578 (O_2578,N_24962,N_24801);
nor UO_2579 (O_2579,N_24268,N_23861);
xor UO_2580 (O_2580,N_24826,N_24358);
nor UO_2581 (O_2581,N_23940,N_24710);
xnor UO_2582 (O_2582,N_24460,N_24264);
nor UO_2583 (O_2583,N_23972,N_24895);
and UO_2584 (O_2584,N_24721,N_23911);
nand UO_2585 (O_2585,N_24409,N_24740);
nor UO_2586 (O_2586,N_23888,N_24364);
nand UO_2587 (O_2587,N_24693,N_24453);
xnor UO_2588 (O_2588,N_24844,N_24099);
xnor UO_2589 (O_2589,N_24198,N_24139);
xor UO_2590 (O_2590,N_24010,N_24237);
or UO_2591 (O_2591,N_23917,N_24960);
nor UO_2592 (O_2592,N_24430,N_24226);
nor UO_2593 (O_2593,N_24311,N_24714);
or UO_2594 (O_2594,N_24451,N_24605);
and UO_2595 (O_2595,N_24575,N_24488);
xnor UO_2596 (O_2596,N_24413,N_24928);
nor UO_2597 (O_2597,N_24919,N_24247);
and UO_2598 (O_2598,N_24591,N_24928);
or UO_2599 (O_2599,N_24634,N_24438);
xor UO_2600 (O_2600,N_24821,N_24969);
xnor UO_2601 (O_2601,N_23955,N_24948);
nand UO_2602 (O_2602,N_24596,N_24923);
and UO_2603 (O_2603,N_24597,N_24119);
and UO_2604 (O_2604,N_24688,N_24534);
nand UO_2605 (O_2605,N_24592,N_24327);
nor UO_2606 (O_2606,N_24328,N_24457);
xnor UO_2607 (O_2607,N_24120,N_24379);
xor UO_2608 (O_2608,N_24415,N_24729);
nor UO_2609 (O_2609,N_24045,N_24468);
nand UO_2610 (O_2610,N_24578,N_24819);
xor UO_2611 (O_2611,N_24977,N_24626);
nand UO_2612 (O_2612,N_24097,N_24149);
or UO_2613 (O_2613,N_24586,N_23804);
and UO_2614 (O_2614,N_23902,N_24561);
nand UO_2615 (O_2615,N_23818,N_24695);
and UO_2616 (O_2616,N_24834,N_23776);
xnor UO_2617 (O_2617,N_24576,N_23807);
or UO_2618 (O_2618,N_24815,N_23825);
xnor UO_2619 (O_2619,N_23983,N_24118);
and UO_2620 (O_2620,N_24883,N_24259);
and UO_2621 (O_2621,N_24032,N_24005);
nand UO_2622 (O_2622,N_24801,N_24376);
nand UO_2623 (O_2623,N_24787,N_24312);
and UO_2624 (O_2624,N_24938,N_24831);
nor UO_2625 (O_2625,N_24285,N_24173);
or UO_2626 (O_2626,N_24091,N_24015);
or UO_2627 (O_2627,N_24965,N_23774);
or UO_2628 (O_2628,N_24842,N_24357);
nand UO_2629 (O_2629,N_24568,N_23938);
nand UO_2630 (O_2630,N_23951,N_24161);
xor UO_2631 (O_2631,N_24300,N_24448);
and UO_2632 (O_2632,N_24578,N_24032);
and UO_2633 (O_2633,N_24091,N_24529);
xnor UO_2634 (O_2634,N_24580,N_23807);
or UO_2635 (O_2635,N_23991,N_24692);
nor UO_2636 (O_2636,N_24692,N_24778);
nor UO_2637 (O_2637,N_24599,N_24827);
nor UO_2638 (O_2638,N_23985,N_24877);
nor UO_2639 (O_2639,N_24684,N_24542);
xnor UO_2640 (O_2640,N_24649,N_24055);
xnor UO_2641 (O_2641,N_24047,N_23934);
and UO_2642 (O_2642,N_24890,N_24179);
nor UO_2643 (O_2643,N_24128,N_24901);
nor UO_2644 (O_2644,N_24451,N_24228);
nand UO_2645 (O_2645,N_23974,N_24720);
xor UO_2646 (O_2646,N_23846,N_24293);
nor UO_2647 (O_2647,N_24221,N_24408);
or UO_2648 (O_2648,N_24664,N_24556);
xnor UO_2649 (O_2649,N_24564,N_24159);
xnor UO_2650 (O_2650,N_23864,N_24169);
nor UO_2651 (O_2651,N_23922,N_23905);
xor UO_2652 (O_2652,N_24711,N_24564);
and UO_2653 (O_2653,N_24022,N_24081);
xnor UO_2654 (O_2654,N_24716,N_24318);
nand UO_2655 (O_2655,N_23755,N_24898);
xor UO_2656 (O_2656,N_24465,N_24172);
nand UO_2657 (O_2657,N_24576,N_23855);
and UO_2658 (O_2658,N_24833,N_24773);
and UO_2659 (O_2659,N_24646,N_24693);
nand UO_2660 (O_2660,N_24117,N_24503);
nor UO_2661 (O_2661,N_24335,N_24355);
xor UO_2662 (O_2662,N_23923,N_24128);
or UO_2663 (O_2663,N_24028,N_24916);
nor UO_2664 (O_2664,N_24913,N_24308);
nand UO_2665 (O_2665,N_24454,N_24421);
nor UO_2666 (O_2666,N_24755,N_24953);
nand UO_2667 (O_2667,N_24425,N_24967);
or UO_2668 (O_2668,N_23933,N_24980);
nor UO_2669 (O_2669,N_23960,N_23927);
xnor UO_2670 (O_2670,N_24235,N_24366);
nand UO_2671 (O_2671,N_24708,N_23790);
nand UO_2672 (O_2672,N_24908,N_24866);
and UO_2673 (O_2673,N_24420,N_24310);
nor UO_2674 (O_2674,N_24299,N_24688);
or UO_2675 (O_2675,N_24714,N_24538);
xnor UO_2676 (O_2676,N_24794,N_24526);
nor UO_2677 (O_2677,N_24547,N_24896);
xnor UO_2678 (O_2678,N_24634,N_24676);
nor UO_2679 (O_2679,N_23998,N_24898);
xnor UO_2680 (O_2680,N_24833,N_24149);
xnor UO_2681 (O_2681,N_23981,N_23909);
or UO_2682 (O_2682,N_24532,N_24172);
nand UO_2683 (O_2683,N_24995,N_24980);
nand UO_2684 (O_2684,N_24173,N_24406);
xor UO_2685 (O_2685,N_24636,N_24682);
nand UO_2686 (O_2686,N_24874,N_24834);
nand UO_2687 (O_2687,N_24101,N_24053);
nand UO_2688 (O_2688,N_23850,N_24600);
nand UO_2689 (O_2689,N_24704,N_24202);
nand UO_2690 (O_2690,N_24946,N_24763);
nor UO_2691 (O_2691,N_24746,N_23943);
xnor UO_2692 (O_2692,N_24137,N_24927);
nand UO_2693 (O_2693,N_24255,N_24938);
and UO_2694 (O_2694,N_24915,N_24853);
nand UO_2695 (O_2695,N_24978,N_24935);
xnor UO_2696 (O_2696,N_24046,N_24217);
and UO_2697 (O_2697,N_24248,N_23857);
nor UO_2698 (O_2698,N_24190,N_24346);
or UO_2699 (O_2699,N_24750,N_24117);
or UO_2700 (O_2700,N_24300,N_23851);
nand UO_2701 (O_2701,N_24904,N_24776);
xor UO_2702 (O_2702,N_24001,N_24212);
nor UO_2703 (O_2703,N_23778,N_24702);
and UO_2704 (O_2704,N_24374,N_24401);
and UO_2705 (O_2705,N_24933,N_24073);
nor UO_2706 (O_2706,N_24444,N_24320);
or UO_2707 (O_2707,N_24822,N_23825);
nand UO_2708 (O_2708,N_23956,N_24458);
or UO_2709 (O_2709,N_24644,N_24506);
nor UO_2710 (O_2710,N_24704,N_24635);
xnor UO_2711 (O_2711,N_24479,N_24549);
nand UO_2712 (O_2712,N_24609,N_24802);
and UO_2713 (O_2713,N_24359,N_24702);
or UO_2714 (O_2714,N_23956,N_23957);
nand UO_2715 (O_2715,N_24285,N_24300);
or UO_2716 (O_2716,N_24371,N_24723);
and UO_2717 (O_2717,N_24418,N_24670);
or UO_2718 (O_2718,N_23962,N_23981);
nand UO_2719 (O_2719,N_24706,N_24342);
or UO_2720 (O_2720,N_24746,N_24031);
and UO_2721 (O_2721,N_24136,N_24042);
or UO_2722 (O_2722,N_24877,N_24288);
or UO_2723 (O_2723,N_24571,N_24732);
or UO_2724 (O_2724,N_23863,N_23823);
xor UO_2725 (O_2725,N_24425,N_24750);
or UO_2726 (O_2726,N_23874,N_24912);
nand UO_2727 (O_2727,N_24669,N_24826);
or UO_2728 (O_2728,N_24282,N_24737);
xor UO_2729 (O_2729,N_24905,N_24080);
and UO_2730 (O_2730,N_24308,N_24825);
nor UO_2731 (O_2731,N_24020,N_23987);
nor UO_2732 (O_2732,N_24496,N_24228);
xnor UO_2733 (O_2733,N_24926,N_24214);
nor UO_2734 (O_2734,N_24773,N_24195);
nand UO_2735 (O_2735,N_24470,N_24006);
nor UO_2736 (O_2736,N_24551,N_24621);
or UO_2737 (O_2737,N_23900,N_24224);
xnor UO_2738 (O_2738,N_24368,N_24984);
nand UO_2739 (O_2739,N_23908,N_24692);
xnor UO_2740 (O_2740,N_24610,N_24971);
nand UO_2741 (O_2741,N_24266,N_24980);
nor UO_2742 (O_2742,N_24339,N_24694);
nor UO_2743 (O_2743,N_24426,N_24716);
xnor UO_2744 (O_2744,N_24176,N_24442);
nand UO_2745 (O_2745,N_24975,N_24095);
xnor UO_2746 (O_2746,N_23827,N_23798);
nor UO_2747 (O_2747,N_24880,N_24948);
and UO_2748 (O_2748,N_24528,N_24318);
nor UO_2749 (O_2749,N_24783,N_24068);
nand UO_2750 (O_2750,N_24514,N_24006);
xor UO_2751 (O_2751,N_24743,N_24163);
nor UO_2752 (O_2752,N_23884,N_24218);
nand UO_2753 (O_2753,N_24993,N_24469);
or UO_2754 (O_2754,N_24221,N_24075);
and UO_2755 (O_2755,N_24867,N_24054);
nand UO_2756 (O_2756,N_24816,N_24027);
and UO_2757 (O_2757,N_24403,N_24346);
and UO_2758 (O_2758,N_24713,N_24999);
xor UO_2759 (O_2759,N_24447,N_24220);
nor UO_2760 (O_2760,N_23783,N_24635);
nor UO_2761 (O_2761,N_24797,N_23788);
and UO_2762 (O_2762,N_24516,N_24208);
or UO_2763 (O_2763,N_23995,N_24909);
xnor UO_2764 (O_2764,N_23944,N_24090);
nand UO_2765 (O_2765,N_23908,N_24349);
and UO_2766 (O_2766,N_24238,N_23824);
nand UO_2767 (O_2767,N_23966,N_23972);
xnor UO_2768 (O_2768,N_23854,N_24390);
and UO_2769 (O_2769,N_24005,N_24942);
nand UO_2770 (O_2770,N_23907,N_24405);
nand UO_2771 (O_2771,N_24796,N_24954);
and UO_2772 (O_2772,N_24665,N_24975);
or UO_2773 (O_2773,N_24682,N_24578);
or UO_2774 (O_2774,N_24132,N_24006);
and UO_2775 (O_2775,N_24881,N_24200);
nand UO_2776 (O_2776,N_24328,N_23769);
or UO_2777 (O_2777,N_24437,N_24673);
or UO_2778 (O_2778,N_24357,N_24449);
xnor UO_2779 (O_2779,N_24604,N_24653);
and UO_2780 (O_2780,N_24313,N_24288);
or UO_2781 (O_2781,N_24582,N_24816);
or UO_2782 (O_2782,N_24629,N_23979);
or UO_2783 (O_2783,N_24867,N_24383);
nor UO_2784 (O_2784,N_24390,N_24298);
and UO_2785 (O_2785,N_24908,N_24692);
or UO_2786 (O_2786,N_24490,N_23823);
nand UO_2787 (O_2787,N_24919,N_24781);
xnor UO_2788 (O_2788,N_24939,N_24925);
xnor UO_2789 (O_2789,N_24000,N_24923);
or UO_2790 (O_2790,N_24959,N_24033);
and UO_2791 (O_2791,N_23864,N_24930);
nand UO_2792 (O_2792,N_24984,N_24353);
nand UO_2793 (O_2793,N_23837,N_24572);
xor UO_2794 (O_2794,N_24265,N_24559);
xnor UO_2795 (O_2795,N_23838,N_23857);
nand UO_2796 (O_2796,N_24576,N_23944);
nor UO_2797 (O_2797,N_24178,N_24505);
and UO_2798 (O_2798,N_24842,N_24308);
or UO_2799 (O_2799,N_24879,N_23940);
xnor UO_2800 (O_2800,N_23880,N_24453);
nand UO_2801 (O_2801,N_24714,N_24918);
nor UO_2802 (O_2802,N_24174,N_24861);
nand UO_2803 (O_2803,N_24032,N_24256);
xnor UO_2804 (O_2804,N_23848,N_24875);
xor UO_2805 (O_2805,N_23919,N_24012);
nand UO_2806 (O_2806,N_24688,N_24130);
and UO_2807 (O_2807,N_24717,N_24910);
nor UO_2808 (O_2808,N_24080,N_24025);
xnor UO_2809 (O_2809,N_24417,N_24482);
xor UO_2810 (O_2810,N_24037,N_23809);
xnor UO_2811 (O_2811,N_24450,N_24198);
or UO_2812 (O_2812,N_24822,N_24544);
nand UO_2813 (O_2813,N_24361,N_24482);
nor UO_2814 (O_2814,N_24803,N_24343);
nand UO_2815 (O_2815,N_24753,N_24557);
nand UO_2816 (O_2816,N_24556,N_23765);
and UO_2817 (O_2817,N_24067,N_24051);
xor UO_2818 (O_2818,N_24146,N_24756);
or UO_2819 (O_2819,N_24312,N_23938);
nand UO_2820 (O_2820,N_24852,N_24649);
nor UO_2821 (O_2821,N_23879,N_24501);
nand UO_2822 (O_2822,N_24933,N_24274);
or UO_2823 (O_2823,N_23849,N_24069);
and UO_2824 (O_2824,N_24341,N_23945);
and UO_2825 (O_2825,N_23825,N_24328);
or UO_2826 (O_2826,N_24066,N_24671);
or UO_2827 (O_2827,N_24863,N_24998);
xor UO_2828 (O_2828,N_24429,N_23911);
and UO_2829 (O_2829,N_23885,N_24753);
xor UO_2830 (O_2830,N_23983,N_24886);
and UO_2831 (O_2831,N_24592,N_23966);
or UO_2832 (O_2832,N_24772,N_24376);
or UO_2833 (O_2833,N_24478,N_24044);
nand UO_2834 (O_2834,N_23781,N_24550);
xnor UO_2835 (O_2835,N_24093,N_24309);
or UO_2836 (O_2836,N_23871,N_24314);
or UO_2837 (O_2837,N_24424,N_23991);
nor UO_2838 (O_2838,N_24209,N_23955);
or UO_2839 (O_2839,N_24974,N_24506);
nor UO_2840 (O_2840,N_24095,N_24972);
nor UO_2841 (O_2841,N_24809,N_24891);
xnor UO_2842 (O_2842,N_24324,N_23879);
xor UO_2843 (O_2843,N_24514,N_24864);
nor UO_2844 (O_2844,N_24212,N_24825);
or UO_2845 (O_2845,N_24583,N_23796);
or UO_2846 (O_2846,N_24737,N_24528);
nand UO_2847 (O_2847,N_24847,N_24148);
and UO_2848 (O_2848,N_24858,N_24454);
nand UO_2849 (O_2849,N_24253,N_24058);
xor UO_2850 (O_2850,N_24868,N_24734);
nor UO_2851 (O_2851,N_24754,N_23928);
xnor UO_2852 (O_2852,N_24225,N_24434);
and UO_2853 (O_2853,N_24558,N_24905);
nand UO_2854 (O_2854,N_24425,N_24819);
and UO_2855 (O_2855,N_23765,N_24753);
or UO_2856 (O_2856,N_24749,N_24822);
and UO_2857 (O_2857,N_24508,N_23880);
or UO_2858 (O_2858,N_24496,N_24459);
nand UO_2859 (O_2859,N_24120,N_24690);
nand UO_2860 (O_2860,N_24693,N_23772);
nor UO_2861 (O_2861,N_24191,N_24643);
nor UO_2862 (O_2862,N_24388,N_24978);
or UO_2863 (O_2863,N_24258,N_23830);
xor UO_2864 (O_2864,N_23902,N_24786);
or UO_2865 (O_2865,N_24413,N_24480);
xor UO_2866 (O_2866,N_24702,N_24302);
xor UO_2867 (O_2867,N_24698,N_24279);
nand UO_2868 (O_2868,N_23883,N_24507);
xnor UO_2869 (O_2869,N_24168,N_24935);
xor UO_2870 (O_2870,N_24540,N_24525);
and UO_2871 (O_2871,N_24000,N_24259);
and UO_2872 (O_2872,N_24394,N_24323);
xnor UO_2873 (O_2873,N_23904,N_23839);
nand UO_2874 (O_2874,N_24102,N_24303);
xor UO_2875 (O_2875,N_24692,N_24046);
xor UO_2876 (O_2876,N_24627,N_24510);
nand UO_2877 (O_2877,N_24251,N_23899);
or UO_2878 (O_2878,N_24751,N_24494);
and UO_2879 (O_2879,N_24571,N_24139);
xnor UO_2880 (O_2880,N_24231,N_24792);
nor UO_2881 (O_2881,N_24907,N_23760);
and UO_2882 (O_2882,N_24218,N_24586);
xnor UO_2883 (O_2883,N_23952,N_24554);
and UO_2884 (O_2884,N_24664,N_24577);
or UO_2885 (O_2885,N_24468,N_23799);
or UO_2886 (O_2886,N_23929,N_24188);
nand UO_2887 (O_2887,N_24138,N_24474);
nand UO_2888 (O_2888,N_24982,N_24563);
nor UO_2889 (O_2889,N_23863,N_24637);
nand UO_2890 (O_2890,N_24628,N_24830);
nand UO_2891 (O_2891,N_24649,N_23809);
or UO_2892 (O_2892,N_24815,N_24505);
or UO_2893 (O_2893,N_24228,N_24665);
xnor UO_2894 (O_2894,N_24773,N_24644);
nor UO_2895 (O_2895,N_24120,N_24479);
xor UO_2896 (O_2896,N_24569,N_24104);
or UO_2897 (O_2897,N_24027,N_24968);
xor UO_2898 (O_2898,N_24591,N_24451);
and UO_2899 (O_2899,N_24222,N_24165);
or UO_2900 (O_2900,N_24371,N_24450);
nand UO_2901 (O_2901,N_24349,N_24135);
nor UO_2902 (O_2902,N_24945,N_23794);
or UO_2903 (O_2903,N_24347,N_24885);
nor UO_2904 (O_2904,N_24993,N_24412);
or UO_2905 (O_2905,N_24467,N_23921);
nor UO_2906 (O_2906,N_24423,N_23778);
and UO_2907 (O_2907,N_24345,N_24339);
nor UO_2908 (O_2908,N_24894,N_24716);
nor UO_2909 (O_2909,N_24291,N_23868);
xnor UO_2910 (O_2910,N_24315,N_24797);
xor UO_2911 (O_2911,N_24840,N_23858);
xnor UO_2912 (O_2912,N_24618,N_24762);
xnor UO_2913 (O_2913,N_24620,N_24186);
nor UO_2914 (O_2914,N_23810,N_24202);
nor UO_2915 (O_2915,N_24975,N_24255);
nand UO_2916 (O_2916,N_24610,N_23809);
nor UO_2917 (O_2917,N_24396,N_23963);
or UO_2918 (O_2918,N_24052,N_24285);
or UO_2919 (O_2919,N_23940,N_23816);
or UO_2920 (O_2920,N_24802,N_24830);
nand UO_2921 (O_2921,N_24400,N_24780);
xor UO_2922 (O_2922,N_24958,N_24613);
nand UO_2923 (O_2923,N_24367,N_24856);
nor UO_2924 (O_2924,N_23989,N_24799);
or UO_2925 (O_2925,N_24555,N_24828);
or UO_2926 (O_2926,N_24588,N_24918);
and UO_2927 (O_2927,N_24058,N_24959);
nand UO_2928 (O_2928,N_24291,N_24381);
nand UO_2929 (O_2929,N_23754,N_23978);
xnor UO_2930 (O_2930,N_24332,N_24508);
nand UO_2931 (O_2931,N_24886,N_24032);
nand UO_2932 (O_2932,N_24492,N_24508);
and UO_2933 (O_2933,N_24851,N_24876);
nor UO_2934 (O_2934,N_24350,N_23844);
nor UO_2935 (O_2935,N_24043,N_24122);
and UO_2936 (O_2936,N_24386,N_24185);
or UO_2937 (O_2937,N_23840,N_24243);
or UO_2938 (O_2938,N_24310,N_24119);
nand UO_2939 (O_2939,N_24962,N_24516);
xor UO_2940 (O_2940,N_24791,N_24497);
nand UO_2941 (O_2941,N_24501,N_23783);
or UO_2942 (O_2942,N_23771,N_24672);
and UO_2943 (O_2943,N_23986,N_24644);
nor UO_2944 (O_2944,N_23901,N_24769);
or UO_2945 (O_2945,N_24442,N_24786);
and UO_2946 (O_2946,N_24141,N_24659);
nor UO_2947 (O_2947,N_24196,N_24217);
and UO_2948 (O_2948,N_24791,N_24628);
or UO_2949 (O_2949,N_24656,N_24267);
nor UO_2950 (O_2950,N_24928,N_24520);
nor UO_2951 (O_2951,N_24934,N_24433);
nand UO_2952 (O_2952,N_23762,N_24179);
and UO_2953 (O_2953,N_24440,N_24025);
nand UO_2954 (O_2954,N_24769,N_24581);
nand UO_2955 (O_2955,N_24846,N_24057);
xor UO_2956 (O_2956,N_24492,N_24872);
and UO_2957 (O_2957,N_23942,N_23974);
nand UO_2958 (O_2958,N_24761,N_24008);
xnor UO_2959 (O_2959,N_23772,N_24178);
xnor UO_2960 (O_2960,N_24931,N_24548);
nor UO_2961 (O_2961,N_24548,N_24769);
xor UO_2962 (O_2962,N_24825,N_24627);
and UO_2963 (O_2963,N_24098,N_24011);
nor UO_2964 (O_2964,N_24275,N_24620);
nor UO_2965 (O_2965,N_24545,N_23785);
or UO_2966 (O_2966,N_24393,N_24303);
nor UO_2967 (O_2967,N_23829,N_24690);
and UO_2968 (O_2968,N_24288,N_24316);
nor UO_2969 (O_2969,N_24905,N_24432);
nor UO_2970 (O_2970,N_24640,N_24383);
nand UO_2971 (O_2971,N_24931,N_24220);
nor UO_2972 (O_2972,N_24542,N_23915);
or UO_2973 (O_2973,N_24931,N_24329);
and UO_2974 (O_2974,N_24195,N_24110);
xor UO_2975 (O_2975,N_24111,N_23847);
xnor UO_2976 (O_2976,N_24540,N_24345);
nand UO_2977 (O_2977,N_24555,N_24907);
or UO_2978 (O_2978,N_24887,N_24221);
nand UO_2979 (O_2979,N_24282,N_24605);
nand UO_2980 (O_2980,N_24598,N_24360);
nor UO_2981 (O_2981,N_24278,N_24656);
or UO_2982 (O_2982,N_23904,N_23958);
and UO_2983 (O_2983,N_23957,N_24601);
and UO_2984 (O_2984,N_23839,N_24282);
xor UO_2985 (O_2985,N_24407,N_23784);
nor UO_2986 (O_2986,N_24342,N_24081);
nor UO_2987 (O_2987,N_24611,N_24282);
nand UO_2988 (O_2988,N_24525,N_24041);
xor UO_2989 (O_2989,N_23934,N_24096);
xnor UO_2990 (O_2990,N_24054,N_23963);
xor UO_2991 (O_2991,N_24297,N_24783);
nand UO_2992 (O_2992,N_24301,N_23976);
and UO_2993 (O_2993,N_24382,N_24016);
nor UO_2994 (O_2994,N_24493,N_23851);
nor UO_2995 (O_2995,N_24275,N_24126);
xnor UO_2996 (O_2996,N_24278,N_24775);
or UO_2997 (O_2997,N_23935,N_24014);
xor UO_2998 (O_2998,N_24968,N_24754);
and UO_2999 (O_2999,N_24120,N_24861);
endmodule