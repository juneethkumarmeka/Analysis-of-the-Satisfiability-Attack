module basic_1000_10000_1500_20_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_219,In_616);
or U1 (N_1,In_637,In_632);
or U2 (N_2,In_776,In_481);
nand U3 (N_3,In_792,In_657);
nand U4 (N_4,In_382,In_513);
and U5 (N_5,In_325,In_666);
nand U6 (N_6,In_88,In_353);
nand U7 (N_7,In_468,In_475);
xor U8 (N_8,In_774,In_485);
nor U9 (N_9,In_375,In_216);
and U10 (N_10,In_756,In_527);
and U11 (N_11,In_662,In_719);
and U12 (N_12,In_795,In_71);
or U13 (N_13,In_787,In_499);
nand U14 (N_14,In_518,In_901);
and U15 (N_15,In_841,In_115);
nand U16 (N_16,In_168,In_282);
nor U17 (N_17,In_544,In_132);
nand U18 (N_18,In_837,In_596);
nand U19 (N_19,In_29,In_923);
or U20 (N_20,In_346,In_735);
nand U21 (N_21,In_962,In_200);
or U22 (N_22,In_976,In_948);
nand U23 (N_23,In_441,In_9);
and U24 (N_24,In_908,In_278);
nor U25 (N_25,In_136,In_874);
nor U26 (N_26,In_600,In_106);
and U27 (N_27,In_63,In_926);
and U28 (N_28,In_280,In_834);
and U29 (N_29,In_522,In_227);
nand U30 (N_30,In_343,In_224);
nor U31 (N_31,In_618,In_248);
or U32 (N_32,In_928,In_298);
xor U33 (N_33,In_413,In_438);
and U34 (N_34,In_804,In_77);
nand U35 (N_35,In_952,In_226);
nor U36 (N_36,In_698,In_500);
nand U37 (N_37,In_161,In_886);
nand U38 (N_38,In_90,In_425);
nor U39 (N_39,In_41,In_537);
nor U40 (N_40,In_399,In_47);
and U41 (N_41,In_783,In_326);
nor U42 (N_42,In_578,In_558);
and U43 (N_43,In_466,In_162);
nand U44 (N_44,In_66,In_697);
and U45 (N_45,In_535,In_906);
or U46 (N_46,In_942,In_911);
xnor U47 (N_47,In_392,In_480);
or U48 (N_48,In_35,In_609);
nand U49 (N_49,In_46,In_651);
or U50 (N_50,In_31,In_807);
and U51 (N_51,In_212,In_682);
or U52 (N_52,In_541,In_143);
nor U53 (N_53,In_955,In_112);
nor U54 (N_54,In_723,In_983);
xor U55 (N_55,In_564,In_255);
nand U56 (N_56,In_414,In_545);
nand U57 (N_57,In_347,In_510);
and U58 (N_58,In_445,In_389);
or U59 (N_59,In_433,In_201);
xnor U60 (N_60,In_415,In_50);
nand U61 (N_61,In_715,In_365);
and U62 (N_62,In_802,In_52);
or U63 (N_63,In_214,In_718);
nor U64 (N_64,In_810,In_743);
or U65 (N_65,In_884,In_188);
or U66 (N_66,In_646,In_484);
or U67 (N_67,In_269,In_108);
and U68 (N_68,In_199,In_512);
or U69 (N_69,In_258,In_309);
xnor U70 (N_70,In_203,In_663);
and U71 (N_71,In_547,In_197);
nor U72 (N_72,In_158,In_276);
and U73 (N_73,In_520,In_263);
nand U74 (N_74,In_515,In_281);
and U75 (N_75,In_502,In_702);
nor U76 (N_76,In_888,In_971);
and U77 (N_77,In_991,In_937);
or U78 (N_78,In_166,In_998);
nor U79 (N_79,In_32,In_336);
nor U80 (N_80,In_305,In_92);
and U81 (N_81,In_123,In_924);
nand U82 (N_82,In_431,In_19);
nand U83 (N_83,In_13,In_237);
or U84 (N_84,In_403,In_638);
nor U85 (N_85,In_351,In_992);
or U86 (N_86,In_532,In_525);
and U87 (N_87,In_629,In_33);
nor U88 (N_88,In_267,In_648);
and U89 (N_89,In_368,In_850);
or U90 (N_90,In_519,In_292);
or U91 (N_91,In_922,In_313);
nand U92 (N_92,In_699,In_655);
and U93 (N_93,In_342,In_369);
nor U94 (N_94,In_696,In_241);
nand U95 (N_95,In_411,In_450);
and U96 (N_96,In_630,In_933);
and U97 (N_97,In_60,In_672);
xor U98 (N_98,In_639,In_750);
nor U99 (N_99,In_283,In_504);
and U100 (N_100,In_757,In_891);
nand U101 (N_101,In_711,In_580);
and U102 (N_102,In_885,In_867);
and U103 (N_103,In_586,In_0);
or U104 (N_104,In_437,In_494);
xor U105 (N_105,In_860,In_878);
nor U106 (N_106,In_251,In_229);
nor U107 (N_107,In_287,In_667);
and U108 (N_108,In_549,In_526);
nand U109 (N_109,In_973,In_139);
nand U110 (N_110,In_61,In_551);
or U111 (N_111,In_54,In_728);
or U112 (N_112,In_557,In_337);
and U113 (N_113,In_561,In_974);
or U114 (N_114,In_10,In_395);
nand U115 (N_115,In_636,In_836);
nand U116 (N_116,In_844,In_821);
or U117 (N_117,In_45,In_493);
or U118 (N_118,In_245,In_496);
nor U119 (N_119,In_185,In_864);
nor U120 (N_120,In_684,In_847);
or U121 (N_121,In_291,In_58);
or U122 (N_122,In_588,In_707);
nor U123 (N_123,In_633,In_148);
nor U124 (N_124,In_584,In_279);
or U125 (N_125,In_345,In_205);
nor U126 (N_126,In_175,In_491);
and U127 (N_127,In_271,In_654);
xnor U128 (N_128,In_831,In_330);
and U129 (N_129,In_93,In_746);
and U130 (N_130,In_788,In_661);
nand U131 (N_131,In_645,In_676);
nand U132 (N_132,In_358,In_975);
and U133 (N_133,In_460,In_571);
nand U134 (N_134,In_979,In_808);
nand U135 (N_135,In_310,In_659);
xor U136 (N_136,In_954,In_339);
nand U137 (N_137,In_649,In_814);
and U138 (N_138,In_202,In_57);
xnor U139 (N_139,In_497,In_855);
and U140 (N_140,In_758,In_695);
xor U141 (N_141,In_144,In_215);
or U142 (N_142,In_364,In_833);
xor U143 (N_143,In_542,In_688);
nor U144 (N_144,In_628,In_652);
or U145 (N_145,In_759,In_147);
nand U146 (N_146,In_233,In_898);
nor U147 (N_147,In_304,In_793);
or U148 (N_148,In_989,In_273);
nand U149 (N_149,In_208,In_624);
nor U150 (N_150,In_777,In_30);
or U151 (N_151,In_614,In_936);
or U152 (N_152,In_487,In_261);
nor U153 (N_153,In_581,In_424);
nor U154 (N_154,In_396,In_858);
and U155 (N_155,In_4,In_829);
and U156 (N_156,In_675,In_747);
xor U157 (N_157,In_678,In_761);
and U158 (N_158,In_709,In_416);
or U159 (N_159,In_463,In_977);
and U160 (N_160,In_142,In_400);
nand U161 (N_161,In_83,In_799);
nor U162 (N_162,In_119,In_813);
or U163 (N_163,In_461,In_734);
xnor U164 (N_164,In_934,In_367);
nand U165 (N_165,In_569,In_195);
xnor U166 (N_166,In_12,In_173);
or U167 (N_167,In_902,In_772);
nor U168 (N_168,In_388,In_880);
nand U169 (N_169,In_75,In_37);
or U170 (N_170,In_153,In_939);
and U171 (N_171,In_444,In_660);
xnor U172 (N_172,In_854,In_56);
nor U173 (N_173,In_322,In_565);
nand U174 (N_174,In_341,In_900);
nor U175 (N_175,In_617,In_739);
nand U176 (N_176,In_319,In_247);
or U177 (N_177,In_940,In_988);
nor U178 (N_178,In_819,In_359);
xor U179 (N_179,In_683,In_312);
nor U180 (N_180,In_917,In_270);
or U181 (N_181,In_462,In_442);
nor U182 (N_182,In_963,In_577);
nor U183 (N_183,In_517,In_946);
or U184 (N_184,In_38,In_539);
or U185 (N_185,In_217,In_893);
and U186 (N_186,In_859,In_771);
nor U187 (N_187,In_28,In_753);
and U188 (N_188,In_264,In_713);
or U189 (N_189,In_419,In_386);
nand U190 (N_190,In_111,In_288);
or U191 (N_191,In_289,In_286);
and U192 (N_192,In_501,In_887);
and U193 (N_193,In_78,In_590);
or U194 (N_194,In_664,In_634);
and U195 (N_195,In_406,In_763);
or U196 (N_196,In_910,In_34);
or U197 (N_197,In_209,In_109);
and U198 (N_198,In_26,In_378);
nand U199 (N_199,In_921,In_253);
nand U200 (N_200,In_314,In_915);
xor U201 (N_201,In_256,In_464);
and U202 (N_202,In_881,In_3);
nor U203 (N_203,In_467,In_42);
nand U204 (N_204,In_720,In_374);
nor U205 (N_205,In_252,In_932);
nand U206 (N_206,In_307,In_350);
nand U207 (N_207,In_806,In_140);
and U208 (N_208,In_67,In_693);
nor U209 (N_209,In_94,In_126);
or U210 (N_210,In_87,In_868);
and U211 (N_211,In_553,In_458);
nor U212 (N_212,In_820,In_601);
nor U213 (N_213,In_784,In_478);
nor U214 (N_214,In_703,In_811);
nand U215 (N_215,In_294,In_51);
and U216 (N_216,In_398,In_176);
nor U217 (N_217,In_839,In_89);
nor U218 (N_218,In_391,In_82);
or U219 (N_219,In_762,In_277);
and U220 (N_220,In_731,In_318);
and U221 (N_221,In_435,In_125);
nand U222 (N_222,In_967,In_20);
nor U223 (N_223,In_393,In_303);
xnor U224 (N_224,In_961,In_972);
and U225 (N_225,In_306,In_605);
and U226 (N_226,In_591,In_534);
nor U227 (N_227,In_583,In_301);
nor U228 (N_228,In_285,In_474);
nor U229 (N_229,In_191,In_352);
or U230 (N_230,In_919,In_870);
and U231 (N_231,In_254,In_592);
and U232 (N_232,In_184,In_742);
nand U233 (N_233,In_454,In_754);
or U234 (N_234,In_213,In_121);
or U235 (N_235,In_594,In_643);
nor U236 (N_236,In_27,In_372);
nor U237 (N_237,In_909,In_914);
nor U238 (N_238,In_412,In_427);
nand U239 (N_239,In_320,In_613);
nand U240 (N_240,In_968,In_712);
nand U241 (N_241,In_384,In_579);
and U242 (N_242,In_206,In_91);
or U243 (N_243,In_726,In_449);
and U244 (N_244,In_817,In_187);
xor U245 (N_245,In_997,In_607);
nand U246 (N_246,In_552,In_904);
or U247 (N_247,In_780,In_154);
nand U248 (N_248,In_920,In_647);
nor U249 (N_249,In_790,In_899);
or U250 (N_250,In_958,In_324);
and U251 (N_251,In_823,In_635);
and U252 (N_252,In_48,In_169);
xnor U253 (N_253,In_714,In_152);
nor U254 (N_254,In_913,In_68);
nand U255 (N_255,In_668,In_563);
and U256 (N_256,In_146,In_842);
xor U257 (N_257,In_439,In_421);
and U258 (N_258,In_334,In_210);
xor U259 (N_259,In_721,In_16);
nand U260 (N_260,In_300,In_786);
or U261 (N_261,In_11,In_373);
or U262 (N_262,In_323,In_894);
nand U263 (N_263,In_64,In_947);
and U264 (N_264,In_1,In_452);
nor U265 (N_265,In_2,In_24);
or U266 (N_266,In_238,In_944);
nand U267 (N_267,In_801,In_656);
nand U268 (N_268,In_931,In_555);
or U269 (N_269,In_796,In_567);
nand U270 (N_270,In_507,In_99);
xor U271 (N_271,In_469,In_849);
or U272 (N_272,In_912,In_883);
nand U273 (N_273,In_376,In_627);
xor U274 (N_274,In_677,In_110);
nand U275 (N_275,In_603,In_625);
nor U276 (N_276,In_476,In_486);
nor U277 (N_277,In_770,In_473);
or U278 (N_278,In_907,In_505);
nand U279 (N_279,In_328,In_355);
nor U280 (N_280,In_234,In_929);
xnor U281 (N_281,In_302,In_428);
xor U282 (N_282,In_568,In_686);
or U283 (N_283,In_459,In_327);
or U284 (N_284,In_317,In_163);
or U285 (N_285,In_692,In_812);
xnor U286 (N_286,In_531,In_451);
or U287 (N_287,In_701,In_705);
xnor U288 (N_288,In_354,In_665);
xnor U289 (N_289,In_741,In_953);
nor U290 (N_290,In_540,In_748);
and U291 (N_291,In_262,In_685);
or U292 (N_292,In_598,In_824);
nand U293 (N_293,In_284,In_387);
nor U294 (N_294,In_80,In_22);
and U295 (N_295,In_809,In_852);
or U296 (N_296,In_599,In_390);
nand U297 (N_297,In_815,In_311);
or U298 (N_298,In_615,In_866);
or U299 (N_299,In_872,In_853);
xnor U300 (N_300,In_335,In_479);
or U301 (N_301,In_190,In_689);
and U302 (N_302,In_608,In_366);
and U303 (N_303,In_843,In_401);
or U304 (N_304,In_102,In_363);
and U305 (N_305,In_181,In_430);
xor U306 (N_306,In_631,In_935);
and U307 (N_307,In_950,In_602);
xor U308 (N_308,In_40,In_472);
nand U309 (N_309,In_794,In_380);
nor U310 (N_310,In_658,In_566);
nor U311 (N_311,In_930,In_755);
or U312 (N_312,In_138,In_828);
or U313 (N_313,In_105,In_641);
nand U314 (N_314,In_356,In_681);
nor U315 (N_315,In_69,In_174);
and U316 (N_316,In_621,In_687);
and U317 (N_317,In_239,In_379);
xor U318 (N_318,In_869,In_716);
or U319 (N_319,In_650,In_124);
and U320 (N_320,In_595,In_508);
nand U321 (N_321,In_778,In_137);
xor U322 (N_322,In_133,In_265);
nor U323 (N_323,In_18,In_43);
and U324 (N_324,In_960,In_483);
or U325 (N_325,In_949,In_53);
or U326 (N_326,In_103,In_710);
nand U327 (N_327,In_653,In_85);
or U328 (N_328,In_340,In_503);
nand U329 (N_329,In_482,In_546);
and U330 (N_330,In_207,In_198);
nor U331 (N_331,In_250,In_903);
and U332 (N_332,In_879,In_456);
or U333 (N_333,In_101,In_775);
nand U334 (N_334,In_680,In_259);
nor U335 (N_335,In_896,In_644);
and U336 (N_336,In_471,In_62);
and U337 (N_337,In_418,In_895);
nor U338 (N_338,In_55,In_117);
nand U339 (N_339,In_118,In_36);
xnor U340 (N_340,In_338,In_299);
nor U341 (N_341,In_951,In_768);
nor U342 (N_342,In_562,In_149);
or U343 (N_343,In_72,In_160);
xnor U344 (N_344,In_296,In_211);
nor U345 (N_345,In_822,In_127);
nand U346 (N_346,In_498,In_116);
nand U347 (N_347,In_329,In_877);
or U348 (N_348,In_957,In_766);
nor U349 (N_349,In_290,In_135);
xor U350 (N_350,In_737,In_890);
and U351 (N_351,In_97,In_220);
xnor U352 (N_352,In_17,In_805);
or U353 (N_353,In_362,In_141);
nand U354 (N_354,In_79,In_448);
nor U355 (N_355,In_260,In_446);
or U356 (N_356,In_816,In_407);
xnor U357 (N_357,In_440,In_180);
or U358 (N_358,In_538,In_640);
and U359 (N_359,In_990,In_764);
nor U360 (N_360,In_107,In_984);
nor U361 (N_361,In_98,In_996);
xnor U362 (N_362,In_740,In_744);
nand U363 (N_363,In_785,In_331);
or U364 (N_364,In_453,In_722);
or U365 (N_365,In_704,In_131);
xnor U366 (N_366,In_122,In_179);
nand U367 (N_367,In_708,In_524);
or U368 (N_368,In_84,In_619);
or U369 (N_369,In_875,In_760);
nor U370 (N_370,In_941,In_404);
and U371 (N_371,In_130,In_572);
nand U372 (N_372,In_543,In_426);
nor U373 (N_373,In_423,In_889);
nor U374 (N_374,In_15,In_385);
or U375 (N_375,In_798,In_489);
xor U376 (N_376,In_228,In_610);
and U377 (N_377,In_530,In_194);
or U378 (N_378,In_164,In_495);
nand U379 (N_379,In_321,In_690);
and U380 (N_380,In_791,In_573);
xnor U381 (N_381,In_671,In_871);
nor U382 (N_382,In_410,In_730);
nand U383 (N_383,In_927,In_995);
xnor U384 (N_384,In_892,In_861);
nand U385 (N_385,In_925,In_443);
nand U386 (N_386,In_86,In_96);
or U387 (N_387,In_835,In_268);
or U388 (N_388,In_574,In_986);
nand U389 (N_389,In_5,In_21);
nand U390 (N_390,In_604,In_765);
or U391 (N_391,In_455,In_377);
and U392 (N_392,In_521,In_156);
or U393 (N_393,In_536,In_134);
nand U394 (N_394,In_81,In_59);
nor U395 (N_395,In_232,In_183);
nor U396 (N_396,In_348,In_113);
and U397 (N_397,In_673,In_978);
nor U398 (N_398,In_128,In_752);
nor U399 (N_399,In_857,In_23);
and U400 (N_400,In_120,In_691);
and U401 (N_401,In_170,In_165);
nand U402 (N_402,In_370,In_846);
nor U403 (N_403,In_589,In_204);
or U404 (N_404,In_965,In_49);
and U405 (N_405,In_848,In_308);
nor U406 (N_406,In_606,In_145);
nand U407 (N_407,In_422,In_585);
nor U408 (N_408,In_825,In_779);
nand U409 (N_409,In_943,In_738);
nor U410 (N_410,In_987,In_172);
and U411 (N_411,In_959,In_275);
or U412 (N_412,In_556,In_725);
xnor U413 (N_413,In_420,In_679);
nand U414 (N_414,In_789,In_225);
or U415 (N_415,In_114,In_274);
nand U416 (N_416,In_470,In_182);
nand U417 (N_417,In_73,In_402);
nand U418 (N_418,In_157,In_511);
nor U419 (N_419,In_100,In_417);
and U420 (N_420,In_244,In_432);
xnor U421 (N_421,In_434,In_670);
and U422 (N_422,In_39,In_597);
and U423 (N_423,In_969,In_993);
xor U424 (N_424,In_724,In_297);
or U425 (N_425,In_767,In_827);
nor U426 (N_426,In_272,In_994);
or U427 (N_427,In_151,In_249);
nor U428 (N_428,In_196,In_611);
nor U429 (N_429,In_575,In_243);
or U430 (N_430,In_559,In_492);
nor U431 (N_431,In_70,In_782);
and U432 (N_432,In_964,In_622);
or U433 (N_433,In_838,In_405);
nor U434 (N_434,In_477,In_897);
nand U435 (N_435,In_803,In_832);
or U436 (N_436,In_587,In_295);
or U437 (N_437,In_727,In_905);
or U438 (N_438,In_218,In_999);
or U439 (N_439,In_129,In_956);
or U440 (N_440,In_570,In_488);
nor U441 (N_441,In_159,In_74);
nor U442 (N_442,In_222,In_554);
nand U443 (N_443,In_882,In_150);
nand U444 (N_444,In_246,In_371);
or U445 (N_445,In_230,In_550);
or U446 (N_446,In_193,In_490);
xnor U447 (N_447,In_177,In_523);
nor U448 (N_448,In_576,In_447);
nor U449 (N_449,In_514,In_818);
nor U450 (N_450,In_506,In_257);
and U451 (N_451,In_25,In_845);
or U452 (N_452,In_509,In_223);
and U453 (N_453,In_394,In_349);
or U454 (N_454,In_221,In_76);
and U455 (N_455,In_316,In_862);
and U456 (N_456,In_851,In_612);
and U457 (N_457,In_980,In_315);
and U458 (N_458,In_397,In_266);
and U459 (N_459,In_717,In_945);
or U460 (N_460,In_751,In_970);
or U461 (N_461,In_694,In_781);
xnor U462 (N_462,In_155,In_736);
xnor U463 (N_463,In_44,In_104);
nor U464 (N_464,In_409,In_65);
nand U465 (N_465,In_548,In_436);
nor U466 (N_466,In_408,In_985);
or U467 (N_467,In_465,In_293);
and U468 (N_468,In_429,In_916);
nor U469 (N_469,In_189,In_529);
and U470 (N_470,In_381,In_623);
or U471 (N_471,In_14,In_981);
nor U472 (N_472,In_95,In_733);
or U473 (N_473,In_706,In_171);
or U474 (N_474,In_528,In_457);
or U475 (N_475,In_333,In_745);
nor U476 (N_476,In_186,In_669);
nand U477 (N_477,In_235,In_516);
and U478 (N_478,In_800,In_626);
and U479 (N_479,In_236,In_982);
or U480 (N_480,In_8,In_700);
and U481 (N_481,In_918,In_192);
or U482 (N_482,In_642,In_533);
or U483 (N_483,In_383,In_344);
nand U484 (N_484,In_732,In_876);
or U485 (N_485,In_167,In_620);
and U486 (N_486,In_560,In_582);
or U487 (N_487,In_332,In_360);
or U488 (N_488,In_674,In_240);
nor U489 (N_489,In_966,In_826);
or U490 (N_490,In_749,In_840);
nand U491 (N_491,In_361,In_7);
nand U492 (N_492,In_357,In_6);
nor U493 (N_493,In_865,In_856);
and U494 (N_494,In_863,In_593);
or U495 (N_495,In_938,In_231);
xnor U496 (N_496,In_242,In_797);
or U497 (N_497,In_178,In_773);
and U498 (N_498,In_873,In_769);
nand U499 (N_499,In_830,In_729);
xnor U500 (N_500,N_498,N_187);
nand U501 (N_501,N_276,N_105);
nor U502 (N_502,N_33,N_81);
xor U503 (N_503,N_71,N_435);
xnor U504 (N_504,N_270,N_176);
nand U505 (N_505,N_146,N_250);
or U506 (N_506,N_319,N_348);
or U507 (N_507,N_354,N_403);
nand U508 (N_508,N_343,N_338);
nand U509 (N_509,N_162,N_363);
and U510 (N_510,N_302,N_197);
nand U511 (N_511,N_422,N_122);
and U512 (N_512,N_54,N_254);
and U513 (N_513,N_273,N_66);
and U514 (N_514,N_325,N_42);
and U515 (N_515,N_173,N_334);
nand U516 (N_516,N_305,N_291);
xor U517 (N_517,N_111,N_171);
and U518 (N_518,N_88,N_167);
nand U519 (N_519,N_62,N_241);
or U520 (N_520,N_0,N_245);
xor U521 (N_521,N_295,N_484);
nor U522 (N_522,N_417,N_186);
or U523 (N_523,N_396,N_80);
and U524 (N_524,N_138,N_298);
nand U525 (N_525,N_440,N_421);
xor U526 (N_526,N_7,N_321);
nor U527 (N_527,N_413,N_427);
or U528 (N_528,N_445,N_350);
or U529 (N_529,N_236,N_68);
or U530 (N_530,N_73,N_18);
nand U531 (N_531,N_465,N_458);
or U532 (N_532,N_297,N_103);
and U533 (N_533,N_266,N_136);
nand U534 (N_534,N_324,N_46);
nand U535 (N_535,N_285,N_95);
and U536 (N_536,N_429,N_340);
xor U537 (N_537,N_376,N_320);
nand U538 (N_538,N_199,N_85);
or U539 (N_539,N_117,N_61);
nand U540 (N_540,N_159,N_233);
xor U541 (N_541,N_137,N_418);
nor U542 (N_542,N_147,N_191);
and U543 (N_543,N_131,N_166);
or U544 (N_544,N_257,N_278);
or U545 (N_545,N_386,N_375);
and U546 (N_546,N_240,N_449);
nor U547 (N_547,N_209,N_382);
nand U548 (N_548,N_326,N_204);
nor U549 (N_549,N_43,N_34);
or U550 (N_550,N_96,N_253);
and U551 (N_551,N_144,N_92);
and U552 (N_552,N_450,N_235);
nand U553 (N_553,N_72,N_372);
nand U554 (N_554,N_98,N_102);
nand U555 (N_555,N_267,N_459);
nor U556 (N_556,N_74,N_32);
and U557 (N_557,N_479,N_170);
nand U558 (N_558,N_113,N_263);
nor U559 (N_559,N_93,N_107);
or U560 (N_560,N_351,N_129);
nor U561 (N_561,N_215,N_497);
and U562 (N_562,N_264,N_23);
or U563 (N_563,N_414,N_287);
nand U564 (N_564,N_20,N_224);
xor U565 (N_565,N_499,N_227);
or U566 (N_566,N_332,N_163);
and U567 (N_567,N_4,N_310);
and U568 (N_568,N_416,N_407);
or U569 (N_569,N_193,N_308);
or U570 (N_570,N_304,N_420);
nor U571 (N_571,N_447,N_174);
or U572 (N_572,N_160,N_446);
nand U573 (N_573,N_480,N_393);
nor U574 (N_574,N_238,N_248);
nand U575 (N_575,N_184,N_392);
nor U576 (N_576,N_274,N_369);
and U577 (N_577,N_432,N_424);
or U578 (N_578,N_106,N_94);
or U579 (N_579,N_329,N_261);
nor U580 (N_580,N_269,N_371);
nand U581 (N_581,N_152,N_123);
and U582 (N_582,N_433,N_207);
and U583 (N_583,N_76,N_40);
or U584 (N_584,N_280,N_255);
or U585 (N_585,N_454,N_153);
or U586 (N_586,N_451,N_426);
xnor U587 (N_587,N_145,N_333);
nand U588 (N_588,N_323,N_47);
xnor U589 (N_589,N_288,N_265);
and U590 (N_590,N_322,N_404);
and U591 (N_591,N_150,N_87);
and U592 (N_592,N_190,N_361);
nand U593 (N_593,N_384,N_135);
xor U594 (N_594,N_423,N_489);
and U595 (N_595,N_31,N_344);
nand U596 (N_596,N_15,N_91);
or U597 (N_597,N_303,N_155);
or U598 (N_598,N_448,N_139);
or U599 (N_599,N_203,N_59);
nor U600 (N_600,N_140,N_219);
and U601 (N_601,N_345,N_356);
nand U602 (N_602,N_475,N_364);
nand U603 (N_603,N_286,N_259);
nand U604 (N_604,N_483,N_327);
or U605 (N_605,N_189,N_28);
and U606 (N_606,N_476,N_406);
or U607 (N_607,N_56,N_79);
nor U608 (N_608,N_226,N_358);
nor U609 (N_609,N_208,N_368);
nand U610 (N_610,N_212,N_317);
or U611 (N_611,N_63,N_425);
and U612 (N_612,N_156,N_415);
nand U613 (N_613,N_30,N_130);
nor U614 (N_614,N_178,N_365);
nor U615 (N_615,N_346,N_355);
and U616 (N_616,N_37,N_45);
and U617 (N_617,N_463,N_25);
and U618 (N_618,N_316,N_373);
or U619 (N_619,N_491,N_385);
or U620 (N_620,N_380,N_282);
xor U621 (N_621,N_70,N_496);
and U622 (N_622,N_60,N_457);
or U623 (N_623,N_353,N_228);
nor U624 (N_624,N_360,N_126);
nor U625 (N_625,N_157,N_283);
or U626 (N_626,N_109,N_290);
and U627 (N_627,N_387,N_331);
nand U628 (N_628,N_443,N_211);
nor U629 (N_629,N_337,N_188);
nand U630 (N_630,N_148,N_275);
nand U631 (N_631,N_408,N_17);
nor U632 (N_632,N_22,N_75);
or U633 (N_633,N_258,N_231);
and U634 (N_634,N_3,N_246);
nor U635 (N_635,N_242,N_65);
nand U636 (N_636,N_2,N_108);
or U637 (N_637,N_57,N_216);
nor U638 (N_638,N_296,N_243);
and U639 (N_639,N_391,N_397);
nand U640 (N_640,N_444,N_453);
nor U641 (N_641,N_12,N_64);
nand U642 (N_642,N_177,N_127);
or U643 (N_643,N_35,N_467);
or U644 (N_644,N_110,N_292);
nor U645 (N_645,N_5,N_468);
and U646 (N_646,N_210,N_330);
nand U647 (N_647,N_428,N_134);
nor U648 (N_648,N_50,N_118);
or U649 (N_649,N_82,N_481);
or U650 (N_650,N_39,N_172);
nor U651 (N_651,N_441,N_165);
xnor U652 (N_652,N_202,N_488);
and U653 (N_653,N_206,N_293);
xnor U654 (N_654,N_341,N_115);
nor U655 (N_655,N_52,N_394);
nand U656 (N_656,N_99,N_482);
and U657 (N_657,N_180,N_44);
xor U658 (N_658,N_399,N_460);
nand U659 (N_659,N_464,N_294);
or U660 (N_660,N_472,N_455);
or U661 (N_661,N_120,N_452);
and U662 (N_662,N_461,N_27);
xnor U663 (N_663,N_16,N_112);
or U664 (N_664,N_48,N_161);
nor U665 (N_665,N_299,N_69);
xor U666 (N_666,N_383,N_142);
nor U667 (N_667,N_89,N_133);
and U668 (N_668,N_51,N_192);
or U669 (N_669,N_473,N_362);
and U670 (N_670,N_251,N_143);
or U671 (N_671,N_409,N_495);
nor U672 (N_672,N_336,N_132);
and U673 (N_673,N_284,N_121);
xor U674 (N_674,N_169,N_268);
and U675 (N_675,N_175,N_55);
nand U676 (N_676,N_388,N_77);
and U677 (N_677,N_347,N_366);
nand U678 (N_678,N_128,N_221);
and U679 (N_679,N_434,N_29);
nor U680 (N_680,N_114,N_281);
or U681 (N_681,N_377,N_359);
nand U682 (N_682,N_492,N_437);
nor U683 (N_683,N_141,N_67);
nand U684 (N_684,N_218,N_158);
or U685 (N_685,N_314,N_179);
and U686 (N_686,N_367,N_86);
nand U687 (N_687,N_194,N_222);
nand U688 (N_688,N_78,N_19);
or U689 (N_689,N_6,N_83);
nor U690 (N_690,N_374,N_318);
or U691 (N_691,N_100,N_181);
xor U692 (N_692,N_300,N_395);
and U693 (N_693,N_313,N_412);
and U694 (N_694,N_349,N_164);
xnor U695 (N_695,N_342,N_225);
and U696 (N_696,N_183,N_104);
and U697 (N_697,N_335,N_279);
nor U698 (N_698,N_21,N_9);
nor U699 (N_699,N_390,N_230);
nand U700 (N_700,N_119,N_49);
and U701 (N_701,N_124,N_223);
or U702 (N_702,N_14,N_198);
nor U703 (N_703,N_301,N_256);
nand U704 (N_704,N_442,N_272);
and U705 (N_705,N_213,N_490);
and U706 (N_706,N_168,N_11);
nand U707 (N_707,N_456,N_401);
or U708 (N_708,N_478,N_252);
xor U709 (N_709,N_262,N_357);
nor U710 (N_710,N_244,N_185);
and U711 (N_711,N_485,N_116);
and U712 (N_712,N_149,N_439);
nand U713 (N_713,N_462,N_151);
or U714 (N_714,N_1,N_312);
nor U715 (N_715,N_469,N_8);
and U716 (N_716,N_307,N_378);
or U717 (N_717,N_410,N_271);
xor U718 (N_718,N_339,N_24);
nand U719 (N_719,N_486,N_436);
nor U720 (N_720,N_306,N_487);
or U721 (N_721,N_53,N_494);
and U722 (N_722,N_477,N_154);
or U723 (N_723,N_90,N_26);
and U724 (N_724,N_419,N_205);
and U725 (N_725,N_237,N_381);
or U726 (N_726,N_239,N_466);
and U727 (N_727,N_370,N_400);
and U728 (N_728,N_328,N_311);
nand U729 (N_729,N_58,N_41);
nor U730 (N_730,N_493,N_84);
nand U731 (N_731,N_97,N_352);
and U732 (N_732,N_431,N_438);
nand U733 (N_733,N_402,N_38);
xnor U734 (N_734,N_125,N_247);
nor U735 (N_735,N_182,N_200);
or U736 (N_736,N_220,N_201);
and U737 (N_737,N_398,N_101);
and U738 (N_738,N_309,N_289);
and U739 (N_739,N_249,N_430);
or U740 (N_740,N_217,N_234);
nor U741 (N_741,N_195,N_232);
or U742 (N_742,N_10,N_277);
nor U743 (N_743,N_260,N_13);
nor U744 (N_744,N_315,N_196);
or U745 (N_745,N_471,N_229);
nand U746 (N_746,N_405,N_411);
nand U747 (N_747,N_389,N_214);
nor U748 (N_748,N_379,N_36);
nand U749 (N_749,N_470,N_474);
nand U750 (N_750,N_78,N_203);
and U751 (N_751,N_361,N_227);
nor U752 (N_752,N_477,N_329);
nand U753 (N_753,N_269,N_306);
or U754 (N_754,N_110,N_124);
xnor U755 (N_755,N_350,N_407);
or U756 (N_756,N_297,N_403);
and U757 (N_757,N_326,N_386);
xor U758 (N_758,N_89,N_374);
and U759 (N_759,N_422,N_285);
and U760 (N_760,N_456,N_81);
xor U761 (N_761,N_195,N_210);
or U762 (N_762,N_165,N_323);
or U763 (N_763,N_170,N_231);
and U764 (N_764,N_373,N_49);
nor U765 (N_765,N_131,N_297);
nor U766 (N_766,N_341,N_201);
nand U767 (N_767,N_5,N_87);
or U768 (N_768,N_238,N_223);
or U769 (N_769,N_51,N_426);
and U770 (N_770,N_33,N_226);
nor U771 (N_771,N_465,N_143);
nor U772 (N_772,N_435,N_103);
nand U773 (N_773,N_211,N_476);
or U774 (N_774,N_285,N_480);
nor U775 (N_775,N_64,N_451);
xnor U776 (N_776,N_438,N_198);
nand U777 (N_777,N_440,N_435);
or U778 (N_778,N_26,N_32);
or U779 (N_779,N_346,N_205);
nand U780 (N_780,N_480,N_313);
nor U781 (N_781,N_392,N_456);
xor U782 (N_782,N_366,N_149);
and U783 (N_783,N_140,N_111);
xnor U784 (N_784,N_483,N_450);
and U785 (N_785,N_157,N_442);
nor U786 (N_786,N_294,N_139);
nand U787 (N_787,N_180,N_160);
and U788 (N_788,N_423,N_84);
xor U789 (N_789,N_483,N_187);
nor U790 (N_790,N_48,N_119);
and U791 (N_791,N_463,N_188);
nor U792 (N_792,N_172,N_329);
and U793 (N_793,N_57,N_272);
and U794 (N_794,N_184,N_0);
nor U795 (N_795,N_142,N_256);
and U796 (N_796,N_291,N_106);
nor U797 (N_797,N_304,N_0);
and U798 (N_798,N_114,N_98);
nand U799 (N_799,N_253,N_224);
and U800 (N_800,N_86,N_134);
and U801 (N_801,N_17,N_200);
or U802 (N_802,N_205,N_72);
and U803 (N_803,N_126,N_456);
nand U804 (N_804,N_365,N_468);
and U805 (N_805,N_76,N_391);
nand U806 (N_806,N_445,N_385);
and U807 (N_807,N_131,N_186);
and U808 (N_808,N_213,N_228);
nand U809 (N_809,N_92,N_47);
nand U810 (N_810,N_11,N_161);
nor U811 (N_811,N_322,N_181);
and U812 (N_812,N_324,N_170);
xor U813 (N_813,N_24,N_422);
nand U814 (N_814,N_432,N_115);
nand U815 (N_815,N_258,N_382);
or U816 (N_816,N_173,N_406);
xor U817 (N_817,N_251,N_103);
nor U818 (N_818,N_345,N_391);
nor U819 (N_819,N_434,N_344);
or U820 (N_820,N_487,N_354);
nand U821 (N_821,N_299,N_434);
xnor U822 (N_822,N_3,N_383);
nor U823 (N_823,N_314,N_279);
and U824 (N_824,N_314,N_388);
nand U825 (N_825,N_251,N_6);
nand U826 (N_826,N_132,N_275);
nor U827 (N_827,N_458,N_368);
and U828 (N_828,N_494,N_427);
or U829 (N_829,N_336,N_70);
and U830 (N_830,N_302,N_497);
or U831 (N_831,N_379,N_151);
or U832 (N_832,N_389,N_243);
or U833 (N_833,N_282,N_448);
and U834 (N_834,N_438,N_278);
nor U835 (N_835,N_266,N_75);
or U836 (N_836,N_124,N_259);
and U837 (N_837,N_402,N_290);
or U838 (N_838,N_227,N_334);
nand U839 (N_839,N_102,N_159);
and U840 (N_840,N_248,N_109);
and U841 (N_841,N_245,N_332);
and U842 (N_842,N_237,N_472);
nor U843 (N_843,N_12,N_35);
nand U844 (N_844,N_129,N_156);
and U845 (N_845,N_170,N_388);
nor U846 (N_846,N_458,N_439);
xor U847 (N_847,N_53,N_70);
or U848 (N_848,N_480,N_256);
and U849 (N_849,N_27,N_312);
or U850 (N_850,N_20,N_76);
and U851 (N_851,N_117,N_470);
nand U852 (N_852,N_304,N_233);
or U853 (N_853,N_473,N_142);
and U854 (N_854,N_337,N_251);
nand U855 (N_855,N_263,N_273);
nor U856 (N_856,N_388,N_309);
and U857 (N_857,N_296,N_217);
or U858 (N_858,N_8,N_4);
nand U859 (N_859,N_491,N_186);
and U860 (N_860,N_103,N_270);
xor U861 (N_861,N_69,N_347);
and U862 (N_862,N_472,N_173);
nand U863 (N_863,N_448,N_378);
nor U864 (N_864,N_102,N_422);
xor U865 (N_865,N_37,N_211);
xnor U866 (N_866,N_172,N_452);
or U867 (N_867,N_134,N_45);
and U868 (N_868,N_327,N_364);
and U869 (N_869,N_39,N_163);
nor U870 (N_870,N_225,N_15);
nand U871 (N_871,N_490,N_429);
or U872 (N_872,N_137,N_140);
nor U873 (N_873,N_160,N_152);
and U874 (N_874,N_332,N_66);
or U875 (N_875,N_263,N_134);
xor U876 (N_876,N_153,N_372);
or U877 (N_877,N_495,N_147);
nor U878 (N_878,N_67,N_119);
nand U879 (N_879,N_21,N_139);
xor U880 (N_880,N_11,N_255);
nor U881 (N_881,N_146,N_25);
nand U882 (N_882,N_0,N_196);
nand U883 (N_883,N_44,N_434);
and U884 (N_884,N_326,N_425);
nand U885 (N_885,N_86,N_28);
nor U886 (N_886,N_120,N_438);
nor U887 (N_887,N_284,N_358);
nor U888 (N_888,N_9,N_498);
nand U889 (N_889,N_420,N_340);
xnor U890 (N_890,N_308,N_196);
nor U891 (N_891,N_24,N_297);
or U892 (N_892,N_183,N_135);
nand U893 (N_893,N_241,N_197);
nor U894 (N_894,N_106,N_110);
nor U895 (N_895,N_32,N_498);
xor U896 (N_896,N_118,N_123);
or U897 (N_897,N_336,N_458);
nand U898 (N_898,N_173,N_254);
nand U899 (N_899,N_250,N_135);
nand U900 (N_900,N_96,N_295);
nand U901 (N_901,N_108,N_380);
xnor U902 (N_902,N_158,N_454);
nand U903 (N_903,N_445,N_315);
nand U904 (N_904,N_37,N_458);
nor U905 (N_905,N_378,N_122);
and U906 (N_906,N_171,N_137);
xor U907 (N_907,N_196,N_223);
xnor U908 (N_908,N_401,N_137);
or U909 (N_909,N_161,N_468);
xor U910 (N_910,N_4,N_130);
nor U911 (N_911,N_73,N_249);
nor U912 (N_912,N_42,N_122);
and U913 (N_913,N_130,N_32);
xor U914 (N_914,N_388,N_345);
nand U915 (N_915,N_391,N_483);
or U916 (N_916,N_413,N_281);
and U917 (N_917,N_389,N_351);
and U918 (N_918,N_276,N_436);
or U919 (N_919,N_431,N_406);
and U920 (N_920,N_123,N_356);
nand U921 (N_921,N_205,N_367);
nand U922 (N_922,N_103,N_280);
and U923 (N_923,N_44,N_299);
or U924 (N_924,N_115,N_146);
nor U925 (N_925,N_386,N_55);
and U926 (N_926,N_276,N_96);
and U927 (N_927,N_211,N_336);
xnor U928 (N_928,N_164,N_376);
nor U929 (N_929,N_138,N_227);
nor U930 (N_930,N_30,N_147);
and U931 (N_931,N_158,N_201);
nor U932 (N_932,N_296,N_142);
xnor U933 (N_933,N_245,N_440);
nor U934 (N_934,N_29,N_113);
and U935 (N_935,N_145,N_170);
nand U936 (N_936,N_166,N_400);
nand U937 (N_937,N_445,N_164);
nor U938 (N_938,N_229,N_235);
and U939 (N_939,N_437,N_215);
nor U940 (N_940,N_88,N_238);
and U941 (N_941,N_280,N_100);
or U942 (N_942,N_1,N_343);
nor U943 (N_943,N_479,N_398);
and U944 (N_944,N_174,N_405);
nand U945 (N_945,N_384,N_79);
or U946 (N_946,N_197,N_3);
and U947 (N_947,N_486,N_428);
nand U948 (N_948,N_185,N_310);
nand U949 (N_949,N_82,N_322);
xor U950 (N_950,N_286,N_283);
nand U951 (N_951,N_122,N_315);
nor U952 (N_952,N_462,N_310);
nor U953 (N_953,N_484,N_171);
xnor U954 (N_954,N_499,N_383);
or U955 (N_955,N_370,N_495);
nor U956 (N_956,N_116,N_285);
nand U957 (N_957,N_32,N_193);
nand U958 (N_958,N_369,N_243);
nand U959 (N_959,N_457,N_401);
nor U960 (N_960,N_122,N_477);
nand U961 (N_961,N_308,N_479);
nor U962 (N_962,N_32,N_56);
nand U963 (N_963,N_62,N_195);
xnor U964 (N_964,N_233,N_479);
nor U965 (N_965,N_103,N_15);
or U966 (N_966,N_458,N_435);
xnor U967 (N_967,N_278,N_264);
nor U968 (N_968,N_95,N_161);
nand U969 (N_969,N_81,N_361);
or U970 (N_970,N_187,N_281);
nand U971 (N_971,N_248,N_279);
and U972 (N_972,N_285,N_224);
and U973 (N_973,N_258,N_170);
or U974 (N_974,N_231,N_208);
and U975 (N_975,N_237,N_350);
or U976 (N_976,N_456,N_218);
or U977 (N_977,N_498,N_229);
nor U978 (N_978,N_45,N_256);
and U979 (N_979,N_326,N_370);
or U980 (N_980,N_211,N_420);
nand U981 (N_981,N_296,N_409);
or U982 (N_982,N_265,N_31);
nor U983 (N_983,N_27,N_254);
or U984 (N_984,N_161,N_427);
nand U985 (N_985,N_435,N_277);
and U986 (N_986,N_489,N_59);
and U987 (N_987,N_371,N_498);
nor U988 (N_988,N_199,N_436);
nand U989 (N_989,N_285,N_194);
nand U990 (N_990,N_452,N_394);
nor U991 (N_991,N_409,N_9);
xnor U992 (N_992,N_476,N_203);
xor U993 (N_993,N_278,N_209);
nor U994 (N_994,N_332,N_5);
nor U995 (N_995,N_476,N_284);
or U996 (N_996,N_480,N_96);
or U997 (N_997,N_496,N_300);
and U998 (N_998,N_167,N_198);
or U999 (N_999,N_337,N_381);
xor U1000 (N_1000,N_777,N_575);
nand U1001 (N_1001,N_860,N_692);
and U1002 (N_1002,N_979,N_694);
nor U1003 (N_1003,N_751,N_597);
and U1004 (N_1004,N_539,N_638);
or U1005 (N_1005,N_580,N_780);
and U1006 (N_1006,N_922,N_752);
and U1007 (N_1007,N_619,N_974);
or U1008 (N_1008,N_845,N_559);
or U1009 (N_1009,N_542,N_641);
nand U1010 (N_1010,N_893,N_822);
nand U1011 (N_1011,N_862,N_781);
or U1012 (N_1012,N_525,N_732);
nand U1013 (N_1013,N_537,N_524);
and U1014 (N_1014,N_668,N_661);
nor U1015 (N_1015,N_528,N_927);
or U1016 (N_1016,N_567,N_572);
and U1017 (N_1017,N_851,N_937);
xnor U1018 (N_1018,N_726,N_623);
or U1019 (N_1019,N_949,N_598);
or U1020 (N_1020,N_700,N_776);
and U1021 (N_1021,N_689,N_625);
or U1022 (N_1022,N_866,N_643);
or U1023 (N_1023,N_746,N_676);
and U1024 (N_1024,N_702,N_578);
nor U1025 (N_1025,N_926,N_852);
or U1026 (N_1026,N_991,N_705);
xnor U1027 (N_1027,N_932,N_556);
nand U1028 (N_1028,N_820,N_579);
or U1029 (N_1029,N_651,N_697);
nand U1030 (N_1030,N_936,N_774);
nor U1031 (N_1031,N_510,N_642);
nor U1032 (N_1032,N_711,N_548);
and U1033 (N_1033,N_941,N_929);
nand U1034 (N_1034,N_683,N_735);
nand U1035 (N_1035,N_743,N_827);
and U1036 (N_1036,N_681,N_677);
nand U1037 (N_1037,N_633,N_521);
nand U1038 (N_1038,N_630,N_596);
nand U1039 (N_1039,N_713,N_532);
and U1040 (N_1040,N_759,N_944);
xor U1041 (N_1041,N_673,N_914);
or U1042 (N_1042,N_565,N_576);
and U1043 (N_1043,N_709,N_587);
or U1044 (N_1044,N_989,N_603);
or U1045 (N_1045,N_714,N_832);
or U1046 (N_1046,N_986,N_823);
nor U1047 (N_1047,N_650,N_891);
nand U1048 (N_1048,N_779,N_836);
nand U1049 (N_1049,N_719,N_733);
nand U1050 (N_1050,N_514,N_535);
nor U1051 (N_1051,N_977,N_541);
or U1052 (N_1052,N_876,N_850);
or U1053 (N_1053,N_773,N_943);
and U1054 (N_1054,N_502,N_615);
and U1055 (N_1055,N_720,N_568);
or U1056 (N_1056,N_804,N_574);
nor U1057 (N_1057,N_788,N_819);
nand U1058 (N_1058,N_742,N_782);
or U1059 (N_1059,N_842,N_679);
xnor U1060 (N_1060,N_838,N_730);
xnor U1061 (N_1061,N_736,N_703);
nand U1062 (N_1062,N_560,N_555);
and U1063 (N_1063,N_581,N_583);
nor U1064 (N_1064,N_767,N_810);
nor U1065 (N_1065,N_791,N_815);
and U1066 (N_1066,N_654,N_799);
nand U1067 (N_1067,N_675,N_507);
and U1068 (N_1068,N_976,N_684);
nand U1069 (N_1069,N_883,N_904);
or U1070 (N_1070,N_648,N_853);
nor U1071 (N_1071,N_613,N_628);
nand U1072 (N_1072,N_657,N_811);
or U1073 (N_1073,N_956,N_607);
and U1074 (N_1074,N_513,N_939);
and U1075 (N_1075,N_859,N_898);
nand U1076 (N_1076,N_829,N_723);
nand U1077 (N_1077,N_925,N_950);
or U1078 (N_1078,N_833,N_865);
nand U1079 (N_1079,N_882,N_745);
and U1080 (N_1080,N_887,N_915);
xnor U1081 (N_1081,N_604,N_909);
nor U1082 (N_1082,N_825,N_716);
nand U1083 (N_1083,N_953,N_656);
nor U1084 (N_1084,N_793,N_734);
or U1085 (N_1085,N_518,N_520);
and U1086 (N_1086,N_886,N_770);
and U1087 (N_1087,N_644,N_797);
nor U1088 (N_1088,N_785,N_934);
or U1089 (N_1089,N_896,N_589);
nand U1090 (N_1090,N_757,N_879);
and U1091 (N_1091,N_899,N_921);
or U1092 (N_1092,N_984,N_951);
nor U1093 (N_1093,N_701,N_769);
nand U1094 (N_1094,N_919,N_992);
nand U1095 (N_1095,N_981,N_621);
nand U1096 (N_1096,N_699,N_608);
or U1097 (N_1097,N_629,N_691);
and U1098 (N_1098,N_519,N_987);
and U1099 (N_1099,N_724,N_803);
or U1100 (N_1100,N_729,N_766);
or U1101 (N_1101,N_946,N_858);
nor U1102 (N_1102,N_928,N_594);
nand U1103 (N_1103,N_515,N_855);
or U1104 (N_1104,N_602,N_954);
or U1105 (N_1105,N_687,N_529);
xor U1106 (N_1106,N_617,N_649);
xnor U1107 (N_1107,N_994,N_693);
nand U1108 (N_1108,N_660,N_563);
nor U1109 (N_1109,N_813,N_710);
or U1110 (N_1110,N_554,N_809);
or U1111 (N_1111,N_558,N_698);
and U1112 (N_1112,N_964,N_808);
and U1113 (N_1113,N_652,N_834);
or U1114 (N_1114,N_595,N_999);
nor U1115 (N_1115,N_969,N_636);
and U1116 (N_1116,N_674,N_768);
nand U1117 (N_1117,N_796,N_816);
or U1118 (N_1118,N_933,N_884);
xor U1119 (N_1119,N_846,N_508);
and U1120 (N_1120,N_504,N_647);
nand U1121 (N_1121,N_997,N_990);
and U1122 (N_1122,N_590,N_817);
nor U1123 (N_1123,N_530,N_667);
nor U1124 (N_1124,N_685,N_800);
nand U1125 (N_1125,N_601,N_536);
nand U1126 (N_1126,N_678,N_870);
or U1127 (N_1127,N_721,N_731);
nand U1128 (N_1128,N_841,N_792);
nor U1129 (N_1129,N_787,N_557);
nand U1130 (N_1130,N_889,N_538);
and U1131 (N_1131,N_722,N_947);
and U1132 (N_1132,N_632,N_960);
and U1133 (N_1133,N_533,N_593);
nor U1134 (N_1134,N_737,N_998);
nand U1135 (N_1135,N_942,N_763);
nor U1136 (N_1136,N_540,N_522);
nor U1137 (N_1137,N_562,N_566);
xnor U1138 (N_1138,N_505,N_952);
nand U1139 (N_1139,N_897,N_503);
xor U1140 (N_1140,N_966,N_662);
nor U1141 (N_1141,N_620,N_706);
nor U1142 (N_1142,N_550,N_805);
or U1143 (N_1143,N_848,N_682);
or U1144 (N_1144,N_614,N_807);
or U1145 (N_1145,N_631,N_573);
or U1146 (N_1146,N_948,N_783);
or U1147 (N_1147,N_546,N_912);
and U1148 (N_1148,N_756,N_835);
nor U1149 (N_1149,N_509,N_854);
nor U1150 (N_1150,N_606,N_669);
nand U1151 (N_1151,N_512,N_972);
nor U1152 (N_1152,N_527,N_622);
or U1153 (N_1153,N_516,N_635);
and U1154 (N_1154,N_545,N_672);
or U1155 (N_1155,N_917,N_696);
or U1156 (N_1156,N_847,N_758);
or U1157 (N_1157,N_646,N_959);
and U1158 (N_1158,N_962,N_695);
nand U1159 (N_1159,N_894,N_666);
nor U1160 (N_1160,N_900,N_688);
and U1161 (N_1161,N_963,N_771);
nand U1162 (N_1162,N_890,N_728);
nor U1163 (N_1163,N_826,N_753);
xnor U1164 (N_1164,N_916,N_671);
or U1165 (N_1165,N_996,N_857);
nor U1166 (N_1166,N_961,N_690);
nand U1167 (N_1167,N_784,N_616);
or U1168 (N_1168,N_874,N_940);
xnor U1169 (N_1169,N_741,N_980);
nor U1170 (N_1170,N_588,N_955);
nor U1171 (N_1171,N_895,N_988);
and U1172 (N_1172,N_534,N_831);
xnor U1173 (N_1173,N_888,N_818);
nand U1174 (N_1174,N_707,N_872);
or U1175 (N_1175,N_591,N_968);
and U1176 (N_1176,N_902,N_569);
or U1177 (N_1177,N_821,N_738);
nand U1178 (N_1178,N_618,N_600);
and U1179 (N_1179,N_885,N_718);
and U1180 (N_1180,N_754,N_627);
and U1181 (N_1181,N_856,N_868);
or U1182 (N_1182,N_802,N_965);
nor U1183 (N_1183,N_790,N_907);
and U1184 (N_1184,N_906,N_772);
nand U1185 (N_1185,N_547,N_760);
nand U1186 (N_1186,N_511,N_867);
or U1187 (N_1187,N_892,N_861);
nand U1188 (N_1188,N_544,N_801);
or U1189 (N_1189,N_849,N_670);
nor U1190 (N_1190,N_686,N_975);
and U1191 (N_1191,N_561,N_624);
and U1192 (N_1192,N_585,N_645);
or U1193 (N_1193,N_957,N_634);
nand U1194 (N_1194,N_945,N_715);
xnor U1195 (N_1195,N_840,N_920);
and U1196 (N_1196,N_551,N_871);
xnor U1197 (N_1197,N_930,N_725);
and U1198 (N_1198,N_837,N_995);
nand U1199 (N_1199,N_775,N_967);
nor U1200 (N_1200,N_727,N_740);
nor U1201 (N_1201,N_653,N_978);
or U1202 (N_1202,N_913,N_755);
and U1203 (N_1203,N_626,N_973);
and U1204 (N_1204,N_665,N_982);
or U1205 (N_1205,N_750,N_717);
nand U1206 (N_1206,N_592,N_918);
xor U1207 (N_1207,N_863,N_744);
nor U1208 (N_1208,N_712,N_571);
or U1209 (N_1209,N_501,N_577);
xnor U1210 (N_1210,N_610,N_798);
and U1211 (N_1211,N_765,N_824);
nor U1212 (N_1212,N_983,N_704);
nand U1213 (N_1213,N_609,N_739);
and U1214 (N_1214,N_901,N_748);
or U1215 (N_1215,N_877,N_663);
xor U1216 (N_1216,N_611,N_582);
nor U1217 (N_1217,N_506,N_839);
or U1218 (N_1218,N_806,N_659);
and U1219 (N_1219,N_985,N_599);
nor U1220 (N_1220,N_958,N_655);
nor U1221 (N_1221,N_549,N_910);
and U1222 (N_1222,N_970,N_637);
nor U1223 (N_1223,N_639,N_749);
and U1224 (N_1224,N_764,N_875);
and U1225 (N_1225,N_881,N_523);
nor U1226 (N_1226,N_664,N_931);
or U1227 (N_1227,N_908,N_828);
and U1228 (N_1228,N_878,N_747);
or U1229 (N_1229,N_844,N_923);
or U1230 (N_1230,N_778,N_500);
or U1231 (N_1231,N_789,N_526);
or U1232 (N_1232,N_794,N_553);
nand U1233 (N_1233,N_911,N_880);
or U1234 (N_1234,N_531,N_762);
or U1235 (N_1235,N_543,N_812);
and U1236 (N_1236,N_864,N_552);
or U1237 (N_1237,N_761,N_905);
nor U1238 (N_1238,N_935,N_971);
or U1239 (N_1239,N_584,N_708);
nor U1240 (N_1240,N_830,N_869);
xor U1241 (N_1241,N_795,N_938);
nor U1242 (N_1242,N_993,N_517);
xor U1243 (N_1243,N_814,N_586);
and U1244 (N_1244,N_570,N_903);
nand U1245 (N_1245,N_605,N_680);
or U1246 (N_1246,N_924,N_564);
and U1247 (N_1247,N_843,N_658);
nor U1248 (N_1248,N_873,N_786);
and U1249 (N_1249,N_612,N_640);
nor U1250 (N_1250,N_793,N_848);
nand U1251 (N_1251,N_917,N_652);
and U1252 (N_1252,N_714,N_652);
and U1253 (N_1253,N_659,N_998);
and U1254 (N_1254,N_642,N_729);
or U1255 (N_1255,N_718,N_505);
or U1256 (N_1256,N_554,N_690);
nand U1257 (N_1257,N_919,N_604);
or U1258 (N_1258,N_799,N_694);
nor U1259 (N_1259,N_922,N_836);
nand U1260 (N_1260,N_603,N_529);
xnor U1261 (N_1261,N_983,N_756);
and U1262 (N_1262,N_540,N_802);
and U1263 (N_1263,N_955,N_737);
or U1264 (N_1264,N_720,N_641);
and U1265 (N_1265,N_744,N_837);
and U1266 (N_1266,N_909,N_806);
nor U1267 (N_1267,N_657,N_818);
nor U1268 (N_1268,N_987,N_738);
and U1269 (N_1269,N_977,N_886);
or U1270 (N_1270,N_725,N_968);
and U1271 (N_1271,N_898,N_906);
and U1272 (N_1272,N_706,N_577);
or U1273 (N_1273,N_987,N_554);
nor U1274 (N_1274,N_981,N_751);
and U1275 (N_1275,N_956,N_999);
or U1276 (N_1276,N_791,N_515);
and U1277 (N_1277,N_659,N_661);
and U1278 (N_1278,N_618,N_996);
and U1279 (N_1279,N_664,N_834);
and U1280 (N_1280,N_727,N_629);
xnor U1281 (N_1281,N_964,N_879);
nor U1282 (N_1282,N_650,N_547);
and U1283 (N_1283,N_808,N_983);
or U1284 (N_1284,N_924,N_645);
nand U1285 (N_1285,N_619,N_801);
or U1286 (N_1286,N_880,N_561);
and U1287 (N_1287,N_743,N_505);
or U1288 (N_1288,N_904,N_847);
nand U1289 (N_1289,N_881,N_893);
or U1290 (N_1290,N_600,N_634);
nor U1291 (N_1291,N_662,N_697);
nand U1292 (N_1292,N_609,N_922);
or U1293 (N_1293,N_943,N_651);
or U1294 (N_1294,N_689,N_961);
nand U1295 (N_1295,N_699,N_575);
nand U1296 (N_1296,N_663,N_664);
nand U1297 (N_1297,N_652,N_530);
or U1298 (N_1298,N_819,N_728);
xor U1299 (N_1299,N_511,N_916);
nand U1300 (N_1300,N_938,N_939);
nand U1301 (N_1301,N_719,N_563);
nor U1302 (N_1302,N_619,N_755);
nand U1303 (N_1303,N_506,N_815);
and U1304 (N_1304,N_614,N_630);
nand U1305 (N_1305,N_768,N_615);
and U1306 (N_1306,N_918,N_640);
or U1307 (N_1307,N_759,N_522);
or U1308 (N_1308,N_759,N_654);
nor U1309 (N_1309,N_540,N_694);
nor U1310 (N_1310,N_632,N_810);
or U1311 (N_1311,N_767,N_837);
or U1312 (N_1312,N_783,N_607);
nand U1313 (N_1313,N_986,N_672);
and U1314 (N_1314,N_897,N_983);
xor U1315 (N_1315,N_508,N_532);
xor U1316 (N_1316,N_870,N_572);
and U1317 (N_1317,N_894,N_932);
and U1318 (N_1318,N_616,N_597);
and U1319 (N_1319,N_605,N_738);
nand U1320 (N_1320,N_694,N_817);
or U1321 (N_1321,N_991,N_720);
or U1322 (N_1322,N_721,N_622);
and U1323 (N_1323,N_820,N_576);
xnor U1324 (N_1324,N_926,N_692);
and U1325 (N_1325,N_586,N_737);
or U1326 (N_1326,N_548,N_676);
and U1327 (N_1327,N_805,N_604);
nor U1328 (N_1328,N_654,N_536);
or U1329 (N_1329,N_570,N_961);
and U1330 (N_1330,N_646,N_864);
nor U1331 (N_1331,N_829,N_618);
and U1332 (N_1332,N_887,N_562);
or U1333 (N_1333,N_916,N_807);
or U1334 (N_1334,N_594,N_617);
and U1335 (N_1335,N_715,N_693);
nor U1336 (N_1336,N_655,N_725);
or U1337 (N_1337,N_520,N_777);
and U1338 (N_1338,N_510,N_558);
or U1339 (N_1339,N_975,N_665);
or U1340 (N_1340,N_581,N_843);
or U1341 (N_1341,N_886,N_755);
or U1342 (N_1342,N_879,N_576);
or U1343 (N_1343,N_602,N_611);
nor U1344 (N_1344,N_749,N_718);
nor U1345 (N_1345,N_718,N_557);
and U1346 (N_1346,N_721,N_992);
xnor U1347 (N_1347,N_860,N_594);
nand U1348 (N_1348,N_899,N_998);
nand U1349 (N_1349,N_747,N_617);
nand U1350 (N_1350,N_893,N_775);
nand U1351 (N_1351,N_981,N_640);
or U1352 (N_1352,N_699,N_974);
nor U1353 (N_1353,N_855,N_553);
nand U1354 (N_1354,N_530,N_547);
nor U1355 (N_1355,N_902,N_604);
xor U1356 (N_1356,N_884,N_993);
or U1357 (N_1357,N_615,N_904);
nor U1358 (N_1358,N_888,N_668);
nand U1359 (N_1359,N_796,N_589);
or U1360 (N_1360,N_747,N_512);
nand U1361 (N_1361,N_569,N_570);
nor U1362 (N_1362,N_963,N_839);
nor U1363 (N_1363,N_779,N_942);
xor U1364 (N_1364,N_897,N_727);
or U1365 (N_1365,N_600,N_784);
nand U1366 (N_1366,N_739,N_575);
or U1367 (N_1367,N_790,N_776);
or U1368 (N_1368,N_890,N_848);
nand U1369 (N_1369,N_555,N_689);
or U1370 (N_1370,N_743,N_839);
and U1371 (N_1371,N_735,N_737);
and U1372 (N_1372,N_567,N_892);
or U1373 (N_1373,N_871,N_898);
nand U1374 (N_1374,N_907,N_759);
nor U1375 (N_1375,N_644,N_980);
or U1376 (N_1376,N_658,N_837);
nand U1377 (N_1377,N_669,N_817);
xnor U1378 (N_1378,N_940,N_887);
and U1379 (N_1379,N_901,N_651);
and U1380 (N_1380,N_608,N_890);
xnor U1381 (N_1381,N_533,N_662);
and U1382 (N_1382,N_765,N_807);
and U1383 (N_1383,N_775,N_868);
or U1384 (N_1384,N_502,N_763);
or U1385 (N_1385,N_837,N_726);
xnor U1386 (N_1386,N_953,N_608);
and U1387 (N_1387,N_592,N_922);
and U1388 (N_1388,N_797,N_923);
nor U1389 (N_1389,N_934,N_976);
xnor U1390 (N_1390,N_940,N_839);
nor U1391 (N_1391,N_595,N_892);
nand U1392 (N_1392,N_861,N_894);
and U1393 (N_1393,N_703,N_644);
or U1394 (N_1394,N_665,N_911);
nand U1395 (N_1395,N_721,N_909);
or U1396 (N_1396,N_974,N_662);
nand U1397 (N_1397,N_610,N_882);
nor U1398 (N_1398,N_651,N_796);
nor U1399 (N_1399,N_585,N_760);
or U1400 (N_1400,N_712,N_598);
nand U1401 (N_1401,N_823,N_586);
nor U1402 (N_1402,N_522,N_578);
or U1403 (N_1403,N_676,N_649);
nand U1404 (N_1404,N_521,N_694);
nor U1405 (N_1405,N_953,N_777);
nand U1406 (N_1406,N_746,N_867);
and U1407 (N_1407,N_801,N_960);
nand U1408 (N_1408,N_627,N_571);
xnor U1409 (N_1409,N_506,N_510);
nand U1410 (N_1410,N_806,N_685);
or U1411 (N_1411,N_978,N_849);
xor U1412 (N_1412,N_696,N_781);
and U1413 (N_1413,N_605,N_514);
nor U1414 (N_1414,N_652,N_972);
nand U1415 (N_1415,N_693,N_774);
and U1416 (N_1416,N_856,N_879);
and U1417 (N_1417,N_633,N_736);
nand U1418 (N_1418,N_524,N_741);
and U1419 (N_1419,N_963,N_891);
nor U1420 (N_1420,N_702,N_516);
or U1421 (N_1421,N_998,N_605);
nand U1422 (N_1422,N_796,N_924);
or U1423 (N_1423,N_506,N_582);
xnor U1424 (N_1424,N_845,N_561);
or U1425 (N_1425,N_564,N_742);
or U1426 (N_1426,N_992,N_993);
and U1427 (N_1427,N_572,N_799);
and U1428 (N_1428,N_637,N_603);
or U1429 (N_1429,N_836,N_709);
nor U1430 (N_1430,N_934,N_775);
nand U1431 (N_1431,N_596,N_547);
or U1432 (N_1432,N_564,N_708);
or U1433 (N_1433,N_823,N_868);
and U1434 (N_1434,N_606,N_670);
nor U1435 (N_1435,N_758,N_587);
xor U1436 (N_1436,N_701,N_547);
and U1437 (N_1437,N_759,N_682);
and U1438 (N_1438,N_892,N_537);
and U1439 (N_1439,N_548,N_768);
and U1440 (N_1440,N_542,N_977);
nor U1441 (N_1441,N_613,N_555);
and U1442 (N_1442,N_888,N_551);
nor U1443 (N_1443,N_938,N_647);
xor U1444 (N_1444,N_849,N_900);
nand U1445 (N_1445,N_835,N_711);
xnor U1446 (N_1446,N_605,N_511);
nor U1447 (N_1447,N_873,N_559);
nand U1448 (N_1448,N_727,N_904);
and U1449 (N_1449,N_970,N_865);
and U1450 (N_1450,N_615,N_772);
or U1451 (N_1451,N_971,N_894);
nand U1452 (N_1452,N_842,N_914);
nand U1453 (N_1453,N_712,N_718);
nor U1454 (N_1454,N_760,N_866);
and U1455 (N_1455,N_507,N_964);
nor U1456 (N_1456,N_808,N_873);
nor U1457 (N_1457,N_603,N_606);
nor U1458 (N_1458,N_966,N_609);
nand U1459 (N_1459,N_544,N_807);
and U1460 (N_1460,N_580,N_685);
nor U1461 (N_1461,N_990,N_599);
nor U1462 (N_1462,N_960,N_561);
nand U1463 (N_1463,N_900,N_977);
nand U1464 (N_1464,N_633,N_735);
nand U1465 (N_1465,N_857,N_888);
nor U1466 (N_1466,N_770,N_831);
xor U1467 (N_1467,N_631,N_563);
and U1468 (N_1468,N_941,N_829);
xnor U1469 (N_1469,N_706,N_854);
and U1470 (N_1470,N_914,N_790);
xnor U1471 (N_1471,N_694,N_939);
and U1472 (N_1472,N_543,N_951);
xnor U1473 (N_1473,N_746,N_804);
nand U1474 (N_1474,N_895,N_512);
and U1475 (N_1475,N_545,N_933);
or U1476 (N_1476,N_924,N_807);
xor U1477 (N_1477,N_784,N_739);
or U1478 (N_1478,N_880,N_519);
nand U1479 (N_1479,N_821,N_953);
nand U1480 (N_1480,N_651,N_788);
or U1481 (N_1481,N_534,N_553);
xnor U1482 (N_1482,N_738,N_950);
nand U1483 (N_1483,N_718,N_781);
nor U1484 (N_1484,N_835,N_586);
nor U1485 (N_1485,N_901,N_919);
nor U1486 (N_1486,N_754,N_725);
nand U1487 (N_1487,N_727,N_734);
and U1488 (N_1488,N_598,N_809);
nand U1489 (N_1489,N_907,N_669);
and U1490 (N_1490,N_934,N_629);
and U1491 (N_1491,N_519,N_530);
and U1492 (N_1492,N_875,N_987);
xor U1493 (N_1493,N_966,N_672);
or U1494 (N_1494,N_514,N_709);
nand U1495 (N_1495,N_866,N_740);
nor U1496 (N_1496,N_611,N_801);
or U1497 (N_1497,N_515,N_557);
nand U1498 (N_1498,N_713,N_536);
or U1499 (N_1499,N_772,N_870);
or U1500 (N_1500,N_1441,N_1200);
nor U1501 (N_1501,N_1352,N_1089);
nand U1502 (N_1502,N_1262,N_1258);
and U1503 (N_1503,N_1188,N_1492);
xor U1504 (N_1504,N_1226,N_1364);
xnor U1505 (N_1505,N_1284,N_1291);
nor U1506 (N_1506,N_1056,N_1078);
xor U1507 (N_1507,N_1196,N_1412);
nand U1508 (N_1508,N_1065,N_1091);
and U1509 (N_1509,N_1404,N_1098);
or U1510 (N_1510,N_1152,N_1484);
nor U1511 (N_1511,N_1066,N_1374);
or U1512 (N_1512,N_1452,N_1058);
nor U1513 (N_1513,N_1156,N_1171);
and U1514 (N_1514,N_1032,N_1224);
and U1515 (N_1515,N_1299,N_1231);
nand U1516 (N_1516,N_1038,N_1402);
nand U1517 (N_1517,N_1493,N_1294);
nor U1518 (N_1518,N_1189,N_1315);
and U1519 (N_1519,N_1461,N_1054);
nor U1520 (N_1520,N_1059,N_1096);
and U1521 (N_1521,N_1297,N_1139);
and U1522 (N_1522,N_1261,N_1252);
or U1523 (N_1523,N_1260,N_1403);
or U1524 (N_1524,N_1259,N_1025);
nor U1525 (N_1525,N_1394,N_1415);
and U1526 (N_1526,N_1173,N_1295);
nor U1527 (N_1527,N_1153,N_1186);
xnor U1528 (N_1528,N_1116,N_1311);
nand U1529 (N_1529,N_1466,N_1495);
or U1530 (N_1530,N_1148,N_1353);
and U1531 (N_1531,N_1334,N_1167);
and U1532 (N_1532,N_1278,N_1298);
nand U1533 (N_1533,N_1070,N_1361);
and U1534 (N_1534,N_1419,N_1406);
and U1535 (N_1535,N_1407,N_1192);
nor U1536 (N_1536,N_1379,N_1187);
nand U1537 (N_1537,N_1010,N_1289);
or U1538 (N_1538,N_1075,N_1183);
xnor U1539 (N_1539,N_1445,N_1251);
xnor U1540 (N_1540,N_1444,N_1322);
and U1541 (N_1541,N_1355,N_1399);
nor U1542 (N_1542,N_1017,N_1199);
and U1543 (N_1543,N_1473,N_1293);
and U1544 (N_1544,N_1102,N_1257);
xnor U1545 (N_1545,N_1121,N_1211);
and U1546 (N_1546,N_1208,N_1290);
nand U1547 (N_1547,N_1230,N_1309);
and U1548 (N_1548,N_1314,N_1462);
nand U1549 (N_1549,N_1161,N_1029);
or U1550 (N_1550,N_1474,N_1090);
nand U1551 (N_1551,N_1437,N_1384);
or U1552 (N_1552,N_1067,N_1092);
nor U1553 (N_1553,N_1028,N_1237);
or U1554 (N_1554,N_1351,N_1129);
xor U1555 (N_1555,N_1160,N_1453);
and U1556 (N_1556,N_1382,N_1084);
or U1557 (N_1557,N_1220,N_1286);
nor U1558 (N_1558,N_1477,N_1180);
nand U1559 (N_1559,N_1409,N_1310);
nor U1560 (N_1560,N_1460,N_1296);
or U1561 (N_1561,N_1486,N_1463);
or U1562 (N_1562,N_1303,N_1369);
nand U1563 (N_1563,N_1265,N_1459);
and U1564 (N_1564,N_1104,N_1024);
or U1565 (N_1565,N_1398,N_1165);
nor U1566 (N_1566,N_1305,N_1347);
or U1567 (N_1567,N_1408,N_1113);
or U1568 (N_1568,N_1047,N_1100);
nand U1569 (N_1569,N_1341,N_1420);
and U1570 (N_1570,N_1418,N_1111);
nor U1571 (N_1571,N_1193,N_1045);
nand U1572 (N_1572,N_1469,N_1388);
nor U1573 (N_1573,N_1021,N_1481);
xnor U1574 (N_1574,N_1060,N_1414);
and U1575 (N_1575,N_1362,N_1169);
and U1576 (N_1576,N_1202,N_1467);
and U1577 (N_1577,N_1094,N_1488);
and U1578 (N_1578,N_1069,N_1292);
and U1579 (N_1579,N_1079,N_1057);
and U1580 (N_1580,N_1458,N_1176);
or U1581 (N_1581,N_1138,N_1464);
nand U1582 (N_1582,N_1198,N_1150);
and U1583 (N_1583,N_1308,N_1110);
and U1584 (N_1584,N_1337,N_1031);
and U1585 (N_1585,N_1276,N_1041);
and U1586 (N_1586,N_1327,N_1348);
nand U1587 (N_1587,N_1007,N_1214);
nor U1588 (N_1588,N_1325,N_1105);
and U1589 (N_1589,N_1182,N_1141);
and U1590 (N_1590,N_1479,N_1247);
and U1591 (N_1591,N_1130,N_1307);
and U1592 (N_1592,N_1424,N_1018);
or U1593 (N_1593,N_1178,N_1340);
nand U1594 (N_1594,N_1185,N_1496);
nor U1595 (N_1595,N_1396,N_1003);
nand U1596 (N_1596,N_1433,N_1487);
and U1597 (N_1597,N_1005,N_1175);
nand U1598 (N_1598,N_1376,N_1371);
nor U1599 (N_1599,N_1370,N_1203);
nor U1600 (N_1600,N_1431,N_1287);
xor U1601 (N_1601,N_1030,N_1083);
and U1602 (N_1602,N_1040,N_1168);
nand U1603 (N_1603,N_1266,N_1162);
and U1604 (N_1604,N_1368,N_1076);
xor U1605 (N_1605,N_1391,N_1343);
nor U1606 (N_1606,N_1062,N_1359);
or U1607 (N_1607,N_1248,N_1272);
or U1608 (N_1608,N_1273,N_1228);
nand U1609 (N_1609,N_1264,N_1491);
nand U1610 (N_1610,N_1204,N_1263);
nand U1611 (N_1611,N_1135,N_1326);
nand U1612 (N_1612,N_1335,N_1072);
nand U1613 (N_1613,N_1410,N_1195);
and U1614 (N_1614,N_1373,N_1157);
nor U1615 (N_1615,N_1242,N_1387);
or U1616 (N_1616,N_1367,N_1288);
nor U1617 (N_1617,N_1209,N_1318);
and U1618 (N_1618,N_1422,N_1243);
nand U1619 (N_1619,N_1416,N_1438);
and U1620 (N_1620,N_1234,N_1475);
or U1621 (N_1621,N_1450,N_1312);
nand U1622 (N_1622,N_1313,N_1344);
and U1623 (N_1623,N_1093,N_1143);
nand U1624 (N_1624,N_1390,N_1159);
nand U1625 (N_1625,N_1430,N_1435);
nand U1626 (N_1626,N_1357,N_1282);
or U1627 (N_1627,N_1275,N_1137);
xor U1628 (N_1628,N_1194,N_1306);
and U1629 (N_1629,N_1478,N_1063);
and U1630 (N_1630,N_1468,N_1026);
nand U1631 (N_1631,N_1401,N_1053);
nor U1632 (N_1632,N_1233,N_1016);
xor U1633 (N_1633,N_1285,N_1269);
nor U1634 (N_1634,N_1483,N_1043);
nand U1635 (N_1635,N_1127,N_1363);
nand U1636 (N_1636,N_1440,N_1271);
nor U1637 (N_1637,N_1229,N_1238);
or U1638 (N_1638,N_1074,N_1052);
xor U1639 (N_1639,N_1109,N_1006);
nand U1640 (N_1640,N_1034,N_1423);
nand U1641 (N_1641,N_1342,N_1011);
or U1642 (N_1642,N_1166,N_1358);
xnor U1643 (N_1643,N_1206,N_1304);
nand U1644 (N_1644,N_1434,N_1106);
and U1645 (N_1645,N_1103,N_1133);
nor U1646 (N_1646,N_1476,N_1328);
or U1647 (N_1647,N_1350,N_1244);
nor U1648 (N_1648,N_1158,N_1333);
nand U1649 (N_1649,N_1470,N_1085);
and U1650 (N_1650,N_1221,N_1101);
xnor U1651 (N_1651,N_1174,N_1037);
nor U1652 (N_1652,N_1013,N_1044);
and U1653 (N_1653,N_1471,N_1320);
or U1654 (N_1654,N_1118,N_1154);
and U1655 (N_1655,N_1087,N_1366);
and U1656 (N_1656,N_1035,N_1140);
and U1657 (N_1657,N_1277,N_1077);
nand U1658 (N_1658,N_1147,N_1042);
xnor U1659 (N_1659,N_1122,N_1061);
or U1660 (N_1660,N_1205,N_1223);
and U1661 (N_1661,N_1281,N_1119);
xor U1662 (N_1662,N_1454,N_1490);
nor U1663 (N_1663,N_1088,N_1432);
and U1664 (N_1664,N_1345,N_1389);
nand U1665 (N_1665,N_1197,N_1163);
nand U1666 (N_1666,N_1255,N_1132);
xor U1667 (N_1667,N_1256,N_1279);
nand U1668 (N_1668,N_1012,N_1236);
or U1669 (N_1669,N_1215,N_1219);
or U1670 (N_1670,N_1426,N_1033);
and U1671 (N_1671,N_1126,N_1019);
or U1672 (N_1672,N_1317,N_1405);
or U1673 (N_1673,N_1001,N_1125);
nor U1674 (N_1674,N_1283,N_1201);
or U1675 (N_1675,N_1465,N_1170);
and U1676 (N_1676,N_1360,N_1339);
nand U1677 (N_1677,N_1413,N_1442);
xor U1678 (N_1678,N_1039,N_1191);
or U1679 (N_1679,N_1241,N_1400);
or U1680 (N_1680,N_1080,N_1064);
nor U1681 (N_1681,N_1354,N_1128);
nand U1682 (N_1682,N_1055,N_1117);
nand U1683 (N_1683,N_1151,N_1218);
or U1684 (N_1684,N_1346,N_1356);
xor U1685 (N_1685,N_1393,N_1015);
and U1686 (N_1686,N_1068,N_1120);
and U1687 (N_1687,N_1212,N_1330);
or U1688 (N_1688,N_1099,N_1134);
nand U1689 (N_1689,N_1181,N_1108);
xor U1690 (N_1690,N_1383,N_1319);
or U1691 (N_1691,N_1002,N_1073);
and U1692 (N_1692,N_1082,N_1232);
nor U1693 (N_1693,N_1022,N_1446);
nand U1694 (N_1694,N_1385,N_1097);
and U1695 (N_1695,N_1429,N_1155);
nor U1696 (N_1696,N_1497,N_1428);
nand U1697 (N_1697,N_1381,N_1436);
and U1698 (N_1698,N_1136,N_1494);
or U1699 (N_1699,N_1164,N_1149);
or U1700 (N_1700,N_1112,N_1365);
nand U1701 (N_1701,N_1392,N_1270);
and U1702 (N_1702,N_1417,N_1227);
nor U1703 (N_1703,N_1489,N_1240);
and U1704 (N_1704,N_1411,N_1107);
nor U1705 (N_1705,N_1217,N_1338);
nand U1706 (N_1706,N_1086,N_1280);
nor U1707 (N_1707,N_1020,N_1050);
nand U1708 (N_1708,N_1485,N_1210);
nand U1709 (N_1709,N_1184,N_1146);
nand U1710 (N_1710,N_1332,N_1456);
nor U1711 (N_1711,N_1207,N_1472);
and U1712 (N_1712,N_1451,N_1142);
and U1713 (N_1713,N_1177,N_1179);
and U1714 (N_1714,N_1222,N_1023);
or U1715 (N_1715,N_1145,N_1071);
nor U1716 (N_1716,N_1114,N_1443);
nor U1717 (N_1717,N_1213,N_1267);
nand U1718 (N_1718,N_1268,N_1004);
nor U1719 (N_1719,N_1254,N_1051);
nand U1720 (N_1720,N_1300,N_1000);
or U1721 (N_1721,N_1323,N_1375);
and U1722 (N_1722,N_1225,N_1048);
nor U1723 (N_1723,N_1457,N_1425);
nor U1724 (N_1724,N_1014,N_1245);
and U1725 (N_1725,N_1008,N_1123);
or U1726 (N_1726,N_1331,N_1395);
nand U1727 (N_1727,N_1449,N_1172);
or U1728 (N_1728,N_1447,N_1439);
nor U1729 (N_1729,N_1046,N_1482);
nand U1730 (N_1730,N_1216,N_1253);
and U1731 (N_1731,N_1027,N_1336);
or U1732 (N_1732,N_1124,N_1377);
or U1733 (N_1733,N_1131,N_1372);
or U1734 (N_1734,N_1480,N_1448);
or U1735 (N_1735,N_1378,N_1324);
nor U1736 (N_1736,N_1498,N_1321);
nor U1737 (N_1737,N_1301,N_1380);
nand U1738 (N_1738,N_1455,N_1274);
xnor U1739 (N_1739,N_1036,N_1329);
or U1740 (N_1740,N_1250,N_1427);
and U1741 (N_1741,N_1049,N_1190);
or U1742 (N_1742,N_1009,N_1115);
or U1743 (N_1743,N_1144,N_1349);
and U1744 (N_1744,N_1499,N_1081);
and U1745 (N_1745,N_1386,N_1095);
and U1746 (N_1746,N_1316,N_1239);
and U1747 (N_1747,N_1249,N_1246);
xnor U1748 (N_1748,N_1421,N_1235);
nand U1749 (N_1749,N_1397,N_1302);
or U1750 (N_1750,N_1031,N_1272);
nand U1751 (N_1751,N_1386,N_1282);
and U1752 (N_1752,N_1250,N_1352);
nor U1753 (N_1753,N_1143,N_1172);
nand U1754 (N_1754,N_1388,N_1199);
xor U1755 (N_1755,N_1296,N_1173);
nand U1756 (N_1756,N_1006,N_1063);
and U1757 (N_1757,N_1412,N_1062);
or U1758 (N_1758,N_1081,N_1267);
nand U1759 (N_1759,N_1185,N_1353);
nor U1760 (N_1760,N_1366,N_1086);
or U1761 (N_1761,N_1192,N_1402);
nand U1762 (N_1762,N_1423,N_1224);
nand U1763 (N_1763,N_1094,N_1147);
and U1764 (N_1764,N_1258,N_1487);
xor U1765 (N_1765,N_1093,N_1064);
and U1766 (N_1766,N_1328,N_1408);
or U1767 (N_1767,N_1382,N_1155);
nand U1768 (N_1768,N_1480,N_1243);
nand U1769 (N_1769,N_1079,N_1196);
and U1770 (N_1770,N_1062,N_1008);
nor U1771 (N_1771,N_1412,N_1112);
or U1772 (N_1772,N_1069,N_1370);
nand U1773 (N_1773,N_1038,N_1120);
or U1774 (N_1774,N_1408,N_1412);
xnor U1775 (N_1775,N_1319,N_1015);
or U1776 (N_1776,N_1279,N_1164);
nor U1777 (N_1777,N_1287,N_1223);
nand U1778 (N_1778,N_1060,N_1242);
and U1779 (N_1779,N_1060,N_1370);
and U1780 (N_1780,N_1466,N_1030);
nor U1781 (N_1781,N_1036,N_1172);
or U1782 (N_1782,N_1077,N_1235);
or U1783 (N_1783,N_1447,N_1209);
or U1784 (N_1784,N_1061,N_1388);
nor U1785 (N_1785,N_1352,N_1037);
nand U1786 (N_1786,N_1339,N_1457);
nand U1787 (N_1787,N_1405,N_1474);
or U1788 (N_1788,N_1094,N_1121);
nand U1789 (N_1789,N_1076,N_1134);
and U1790 (N_1790,N_1127,N_1257);
nor U1791 (N_1791,N_1289,N_1208);
and U1792 (N_1792,N_1315,N_1049);
or U1793 (N_1793,N_1270,N_1078);
nor U1794 (N_1794,N_1097,N_1341);
or U1795 (N_1795,N_1416,N_1256);
nand U1796 (N_1796,N_1075,N_1433);
nor U1797 (N_1797,N_1149,N_1451);
and U1798 (N_1798,N_1212,N_1324);
nand U1799 (N_1799,N_1415,N_1237);
and U1800 (N_1800,N_1130,N_1387);
xor U1801 (N_1801,N_1304,N_1316);
and U1802 (N_1802,N_1439,N_1256);
nand U1803 (N_1803,N_1245,N_1176);
and U1804 (N_1804,N_1206,N_1440);
nor U1805 (N_1805,N_1476,N_1316);
nand U1806 (N_1806,N_1395,N_1204);
and U1807 (N_1807,N_1171,N_1105);
xor U1808 (N_1808,N_1281,N_1215);
nor U1809 (N_1809,N_1046,N_1347);
or U1810 (N_1810,N_1020,N_1067);
and U1811 (N_1811,N_1453,N_1373);
nand U1812 (N_1812,N_1020,N_1006);
xor U1813 (N_1813,N_1190,N_1122);
nand U1814 (N_1814,N_1416,N_1011);
or U1815 (N_1815,N_1363,N_1293);
nor U1816 (N_1816,N_1086,N_1180);
or U1817 (N_1817,N_1001,N_1280);
nor U1818 (N_1818,N_1458,N_1161);
and U1819 (N_1819,N_1018,N_1002);
nor U1820 (N_1820,N_1106,N_1322);
and U1821 (N_1821,N_1049,N_1248);
and U1822 (N_1822,N_1483,N_1000);
nand U1823 (N_1823,N_1083,N_1128);
or U1824 (N_1824,N_1495,N_1092);
and U1825 (N_1825,N_1105,N_1316);
and U1826 (N_1826,N_1344,N_1346);
or U1827 (N_1827,N_1125,N_1146);
nor U1828 (N_1828,N_1464,N_1132);
nand U1829 (N_1829,N_1422,N_1374);
nand U1830 (N_1830,N_1372,N_1434);
and U1831 (N_1831,N_1464,N_1113);
nor U1832 (N_1832,N_1344,N_1413);
or U1833 (N_1833,N_1315,N_1083);
or U1834 (N_1834,N_1101,N_1419);
nor U1835 (N_1835,N_1035,N_1153);
xor U1836 (N_1836,N_1157,N_1376);
nor U1837 (N_1837,N_1013,N_1015);
or U1838 (N_1838,N_1217,N_1274);
and U1839 (N_1839,N_1267,N_1170);
nor U1840 (N_1840,N_1285,N_1047);
and U1841 (N_1841,N_1489,N_1104);
nand U1842 (N_1842,N_1074,N_1058);
nor U1843 (N_1843,N_1127,N_1293);
xnor U1844 (N_1844,N_1495,N_1143);
or U1845 (N_1845,N_1011,N_1142);
nand U1846 (N_1846,N_1114,N_1479);
nand U1847 (N_1847,N_1066,N_1067);
or U1848 (N_1848,N_1262,N_1323);
nor U1849 (N_1849,N_1445,N_1472);
nor U1850 (N_1850,N_1321,N_1060);
nor U1851 (N_1851,N_1133,N_1310);
and U1852 (N_1852,N_1018,N_1414);
nand U1853 (N_1853,N_1061,N_1175);
nor U1854 (N_1854,N_1449,N_1355);
nor U1855 (N_1855,N_1073,N_1474);
or U1856 (N_1856,N_1286,N_1381);
nor U1857 (N_1857,N_1042,N_1485);
nor U1858 (N_1858,N_1144,N_1136);
or U1859 (N_1859,N_1376,N_1277);
nand U1860 (N_1860,N_1302,N_1461);
nor U1861 (N_1861,N_1228,N_1204);
or U1862 (N_1862,N_1252,N_1466);
nor U1863 (N_1863,N_1369,N_1172);
and U1864 (N_1864,N_1383,N_1375);
or U1865 (N_1865,N_1070,N_1315);
nor U1866 (N_1866,N_1395,N_1119);
or U1867 (N_1867,N_1120,N_1074);
nor U1868 (N_1868,N_1051,N_1032);
nand U1869 (N_1869,N_1305,N_1331);
or U1870 (N_1870,N_1113,N_1326);
or U1871 (N_1871,N_1323,N_1253);
nor U1872 (N_1872,N_1130,N_1043);
and U1873 (N_1873,N_1096,N_1437);
or U1874 (N_1874,N_1171,N_1299);
nand U1875 (N_1875,N_1171,N_1290);
or U1876 (N_1876,N_1174,N_1352);
and U1877 (N_1877,N_1122,N_1221);
or U1878 (N_1878,N_1270,N_1089);
nor U1879 (N_1879,N_1170,N_1374);
and U1880 (N_1880,N_1169,N_1185);
or U1881 (N_1881,N_1064,N_1443);
xnor U1882 (N_1882,N_1338,N_1256);
and U1883 (N_1883,N_1141,N_1457);
or U1884 (N_1884,N_1489,N_1345);
nor U1885 (N_1885,N_1498,N_1126);
or U1886 (N_1886,N_1408,N_1331);
xor U1887 (N_1887,N_1212,N_1464);
nand U1888 (N_1888,N_1040,N_1295);
or U1889 (N_1889,N_1333,N_1198);
or U1890 (N_1890,N_1403,N_1427);
nor U1891 (N_1891,N_1101,N_1102);
or U1892 (N_1892,N_1093,N_1495);
or U1893 (N_1893,N_1105,N_1483);
nor U1894 (N_1894,N_1362,N_1327);
xnor U1895 (N_1895,N_1207,N_1141);
xnor U1896 (N_1896,N_1385,N_1405);
xnor U1897 (N_1897,N_1059,N_1449);
nor U1898 (N_1898,N_1011,N_1187);
nor U1899 (N_1899,N_1008,N_1246);
or U1900 (N_1900,N_1314,N_1089);
nor U1901 (N_1901,N_1218,N_1359);
or U1902 (N_1902,N_1494,N_1253);
nor U1903 (N_1903,N_1442,N_1134);
and U1904 (N_1904,N_1433,N_1288);
nor U1905 (N_1905,N_1397,N_1048);
or U1906 (N_1906,N_1376,N_1259);
or U1907 (N_1907,N_1396,N_1315);
nor U1908 (N_1908,N_1354,N_1162);
or U1909 (N_1909,N_1097,N_1069);
nand U1910 (N_1910,N_1387,N_1114);
or U1911 (N_1911,N_1232,N_1143);
xnor U1912 (N_1912,N_1370,N_1337);
or U1913 (N_1913,N_1029,N_1128);
or U1914 (N_1914,N_1164,N_1323);
or U1915 (N_1915,N_1437,N_1182);
or U1916 (N_1916,N_1099,N_1322);
nand U1917 (N_1917,N_1359,N_1426);
and U1918 (N_1918,N_1173,N_1050);
nand U1919 (N_1919,N_1084,N_1075);
or U1920 (N_1920,N_1284,N_1466);
and U1921 (N_1921,N_1065,N_1305);
nand U1922 (N_1922,N_1431,N_1047);
nand U1923 (N_1923,N_1118,N_1200);
xor U1924 (N_1924,N_1437,N_1160);
and U1925 (N_1925,N_1189,N_1321);
and U1926 (N_1926,N_1430,N_1159);
and U1927 (N_1927,N_1126,N_1215);
or U1928 (N_1928,N_1147,N_1490);
nand U1929 (N_1929,N_1158,N_1475);
nand U1930 (N_1930,N_1430,N_1403);
nor U1931 (N_1931,N_1400,N_1201);
and U1932 (N_1932,N_1380,N_1308);
or U1933 (N_1933,N_1391,N_1021);
nor U1934 (N_1934,N_1071,N_1256);
and U1935 (N_1935,N_1349,N_1305);
nor U1936 (N_1936,N_1495,N_1494);
and U1937 (N_1937,N_1200,N_1401);
or U1938 (N_1938,N_1062,N_1110);
nor U1939 (N_1939,N_1388,N_1126);
nor U1940 (N_1940,N_1278,N_1023);
and U1941 (N_1941,N_1340,N_1077);
nor U1942 (N_1942,N_1303,N_1113);
or U1943 (N_1943,N_1088,N_1362);
xnor U1944 (N_1944,N_1249,N_1203);
xnor U1945 (N_1945,N_1178,N_1087);
or U1946 (N_1946,N_1254,N_1470);
xnor U1947 (N_1947,N_1140,N_1060);
nor U1948 (N_1948,N_1266,N_1110);
and U1949 (N_1949,N_1168,N_1349);
xor U1950 (N_1950,N_1179,N_1373);
xor U1951 (N_1951,N_1055,N_1469);
and U1952 (N_1952,N_1452,N_1396);
nor U1953 (N_1953,N_1014,N_1143);
nand U1954 (N_1954,N_1432,N_1393);
nor U1955 (N_1955,N_1151,N_1389);
and U1956 (N_1956,N_1073,N_1186);
or U1957 (N_1957,N_1046,N_1233);
or U1958 (N_1958,N_1206,N_1421);
and U1959 (N_1959,N_1228,N_1429);
nor U1960 (N_1960,N_1162,N_1326);
or U1961 (N_1961,N_1113,N_1467);
nand U1962 (N_1962,N_1337,N_1177);
nor U1963 (N_1963,N_1082,N_1120);
and U1964 (N_1964,N_1279,N_1091);
and U1965 (N_1965,N_1281,N_1208);
nand U1966 (N_1966,N_1211,N_1321);
and U1967 (N_1967,N_1135,N_1166);
nor U1968 (N_1968,N_1236,N_1369);
nand U1969 (N_1969,N_1423,N_1427);
xor U1970 (N_1970,N_1494,N_1399);
nand U1971 (N_1971,N_1487,N_1275);
and U1972 (N_1972,N_1159,N_1391);
nor U1973 (N_1973,N_1015,N_1364);
and U1974 (N_1974,N_1239,N_1275);
nand U1975 (N_1975,N_1366,N_1360);
nor U1976 (N_1976,N_1105,N_1337);
xor U1977 (N_1977,N_1430,N_1290);
nor U1978 (N_1978,N_1182,N_1117);
nand U1979 (N_1979,N_1380,N_1294);
nand U1980 (N_1980,N_1103,N_1050);
nand U1981 (N_1981,N_1101,N_1098);
and U1982 (N_1982,N_1052,N_1061);
nand U1983 (N_1983,N_1221,N_1302);
nand U1984 (N_1984,N_1292,N_1178);
nand U1985 (N_1985,N_1266,N_1095);
and U1986 (N_1986,N_1473,N_1284);
and U1987 (N_1987,N_1268,N_1018);
and U1988 (N_1988,N_1169,N_1497);
nor U1989 (N_1989,N_1301,N_1467);
nand U1990 (N_1990,N_1186,N_1021);
and U1991 (N_1991,N_1468,N_1408);
or U1992 (N_1992,N_1191,N_1314);
or U1993 (N_1993,N_1311,N_1219);
xnor U1994 (N_1994,N_1281,N_1263);
and U1995 (N_1995,N_1393,N_1293);
nor U1996 (N_1996,N_1170,N_1229);
nand U1997 (N_1997,N_1280,N_1186);
xnor U1998 (N_1998,N_1384,N_1451);
nand U1999 (N_1999,N_1413,N_1072);
and U2000 (N_2000,N_1885,N_1500);
and U2001 (N_2001,N_1972,N_1613);
nand U2002 (N_2002,N_1846,N_1525);
xnor U2003 (N_2003,N_1679,N_1535);
or U2004 (N_2004,N_1524,N_1526);
or U2005 (N_2005,N_1902,N_1840);
or U2006 (N_2006,N_1804,N_1932);
and U2007 (N_2007,N_1563,N_1510);
or U2008 (N_2008,N_1587,N_1506);
and U2009 (N_2009,N_1700,N_1871);
or U2010 (N_2010,N_1607,N_1838);
and U2011 (N_2011,N_1774,N_1889);
nor U2012 (N_2012,N_1901,N_1865);
and U2013 (N_2013,N_1502,N_1684);
xor U2014 (N_2014,N_1927,N_1945);
nand U2015 (N_2015,N_1995,N_1622);
nand U2016 (N_2016,N_1823,N_1891);
nand U2017 (N_2017,N_1696,N_1964);
nor U2018 (N_2018,N_1826,N_1742);
and U2019 (N_2019,N_1756,N_1773);
and U2020 (N_2020,N_1723,N_1556);
nand U2021 (N_2021,N_1991,N_1783);
nand U2022 (N_2022,N_1565,N_1843);
nor U2023 (N_2023,N_1960,N_1987);
and U2024 (N_2024,N_1743,N_1979);
nor U2025 (N_2025,N_1646,N_1670);
nor U2026 (N_2026,N_1630,N_1806);
nor U2027 (N_2027,N_1916,N_1849);
nor U2028 (N_2028,N_1745,N_1637);
nor U2029 (N_2029,N_1981,N_1878);
nand U2030 (N_2030,N_1610,N_1669);
nand U2031 (N_2031,N_1872,N_1836);
or U2032 (N_2032,N_1812,N_1875);
nand U2033 (N_2033,N_1886,N_1824);
or U2034 (N_2034,N_1677,N_1731);
nand U2035 (N_2035,N_1746,N_1588);
and U2036 (N_2036,N_1811,N_1512);
nor U2037 (N_2037,N_1538,N_1651);
nor U2038 (N_2038,N_1676,N_1989);
nand U2039 (N_2039,N_1844,N_1604);
nor U2040 (N_2040,N_1943,N_1583);
nand U2041 (N_2041,N_1715,N_1664);
or U2042 (N_2042,N_1649,N_1687);
nand U2043 (N_2043,N_1708,N_1534);
or U2044 (N_2044,N_1870,N_1568);
and U2045 (N_2045,N_1599,N_1750);
and U2046 (N_2046,N_1711,N_1815);
nor U2047 (N_2047,N_1958,N_1873);
nor U2048 (N_2048,N_1963,N_1598);
and U2049 (N_2049,N_1673,N_1800);
nand U2050 (N_2050,N_1644,N_1813);
and U2051 (N_2051,N_1909,N_1569);
nand U2052 (N_2052,N_1640,N_1632);
or U2053 (N_2053,N_1877,N_1975);
or U2054 (N_2054,N_1574,N_1597);
nor U2055 (N_2055,N_1798,N_1761);
nor U2056 (N_2056,N_1896,N_1584);
xnor U2057 (N_2057,N_1636,N_1847);
nand U2058 (N_2058,N_1839,N_1566);
and U2059 (N_2059,N_1659,N_1782);
nand U2060 (N_2060,N_1689,N_1984);
and U2061 (N_2061,N_1533,N_1944);
nand U2062 (N_2062,N_1562,N_1888);
or U2063 (N_2063,N_1949,N_1528);
or U2064 (N_2064,N_1970,N_1862);
nor U2065 (N_2065,N_1734,N_1830);
nor U2066 (N_2066,N_1732,N_1952);
nand U2067 (N_2067,N_1937,N_1993);
nor U2068 (N_2068,N_1545,N_1609);
and U2069 (N_2069,N_1805,N_1738);
nand U2070 (N_2070,N_1986,N_1580);
nand U2071 (N_2071,N_1656,N_1959);
nor U2072 (N_2072,N_1540,N_1874);
or U2073 (N_2073,N_1667,N_1605);
or U2074 (N_2074,N_1880,N_1519);
nand U2075 (N_2075,N_1911,N_1736);
xor U2076 (N_2076,N_1567,N_1860);
nand U2077 (N_2077,N_1893,N_1857);
xor U2078 (N_2078,N_1685,N_1808);
and U2079 (N_2079,N_1921,N_1546);
nand U2080 (N_2080,N_1869,N_1940);
nor U2081 (N_2081,N_1527,N_1953);
nor U2082 (N_2082,N_1867,N_1529);
or U2083 (N_2083,N_1905,N_1688);
and U2084 (N_2084,N_1643,N_1917);
nor U2085 (N_2085,N_1661,N_1747);
nand U2086 (N_2086,N_1573,N_1705);
nor U2087 (N_2087,N_1764,N_1942);
or U2088 (N_2088,N_1724,N_1789);
or U2089 (N_2089,N_1814,N_1900);
and U2090 (N_2090,N_1647,N_1908);
nand U2091 (N_2091,N_1759,N_1967);
or U2092 (N_2092,N_1564,N_1976);
or U2093 (N_2093,N_1655,N_1936);
and U2094 (N_2094,N_1611,N_1879);
and U2095 (N_2095,N_1509,N_1654);
nor U2096 (N_2096,N_1956,N_1683);
and U2097 (N_2097,N_1539,N_1749);
or U2098 (N_2098,N_1776,N_1641);
or U2099 (N_2099,N_1786,N_1757);
nor U2100 (N_2100,N_1859,N_1532);
and U2101 (N_2101,N_1861,N_1680);
nor U2102 (N_2102,N_1523,N_1645);
or U2103 (N_2103,N_1765,N_1915);
and U2104 (N_2104,N_1507,N_1744);
nand U2105 (N_2105,N_1864,N_1992);
nor U2106 (N_2106,N_1570,N_1866);
nor U2107 (N_2107,N_1903,N_1616);
nand U2108 (N_2108,N_1631,N_1714);
and U2109 (N_2109,N_1890,N_1833);
or U2110 (N_2110,N_1810,N_1835);
nand U2111 (N_2111,N_1912,N_1777);
or U2112 (N_2112,N_1842,N_1922);
nor U2113 (N_2113,N_1638,N_1508);
and U2114 (N_2114,N_1856,N_1910);
xnor U2115 (N_2115,N_1718,N_1612);
or U2116 (N_2116,N_1627,N_1825);
xor U2117 (N_2117,N_1553,N_1845);
nand U2118 (N_2118,N_1951,N_1628);
or U2119 (N_2119,N_1721,N_1686);
nor U2120 (N_2120,N_1617,N_1618);
and U2121 (N_2121,N_1662,N_1758);
and U2122 (N_2122,N_1555,N_1560);
nor U2123 (N_2123,N_1592,N_1648);
nand U2124 (N_2124,N_1863,N_1822);
nor U2125 (N_2125,N_1692,N_1671);
nor U2126 (N_2126,N_1629,N_1704);
nor U2127 (N_2127,N_1898,N_1751);
nor U2128 (N_2128,N_1977,N_1778);
xor U2129 (N_2129,N_1755,N_1591);
xnor U2130 (N_2130,N_1537,N_1941);
nor U2131 (N_2131,N_1593,N_1884);
or U2132 (N_2132,N_1698,N_1578);
nand U2133 (N_2133,N_1820,N_1969);
nand U2134 (N_2134,N_1858,N_1948);
and U2135 (N_2135,N_1691,N_1624);
and U2136 (N_2136,N_1978,N_1666);
or U2137 (N_2137,N_1728,N_1590);
and U2138 (N_2138,N_1780,N_1876);
xor U2139 (N_2139,N_1663,N_1933);
nand U2140 (N_2140,N_1999,N_1920);
and U2141 (N_2141,N_1904,N_1938);
nor U2142 (N_2142,N_1600,N_1581);
and U2143 (N_2143,N_1753,N_1769);
and U2144 (N_2144,N_1923,N_1931);
nor U2145 (N_2145,N_1816,N_1550);
nor U2146 (N_2146,N_1579,N_1571);
nand U2147 (N_2147,N_1635,N_1703);
nand U2148 (N_2148,N_1980,N_1775);
nand U2149 (N_2149,N_1586,N_1730);
or U2150 (N_2150,N_1536,N_1504);
and U2151 (N_2151,N_1892,N_1620);
and U2152 (N_2152,N_1707,N_1894);
nand U2153 (N_2153,N_1511,N_1794);
or U2154 (N_2154,N_1787,N_1837);
and U2155 (N_2155,N_1996,N_1530);
nand U2156 (N_2156,N_1551,N_1928);
or U2157 (N_2157,N_1602,N_1660);
or U2158 (N_2158,N_1733,N_1828);
or U2159 (N_2159,N_1803,N_1762);
xnor U2160 (N_2160,N_1807,N_1760);
nor U2161 (N_2161,N_1947,N_1619);
and U2162 (N_2162,N_1771,N_1665);
and U2163 (N_2163,N_1541,N_1897);
nand U2164 (N_2164,N_1633,N_1784);
nand U2165 (N_2165,N_1818,N_1906);
and U2166 (N_2166,N_1834,N_1819);
nand U2167 (N_2167,N_1763,N_1547);
xor U2168 (N_2168,N_1766,N_1855);
and U2169 (N_2169,N_1697,N_1682);
xnor U2170 (N_2170,N_1614,N_1841);
xnor U2171 (N_2171,N_1882,N_1994);
or U2172 (N_2172,N_1851,N_1739);
nand U2173 (N_2173,N_1797,N_1693);
nand U2174 (N_2174,N_1998,N_1576);
nor U2175 (N_2175,N_1939,N_1521);
nor U2176 (N_2176,N_1919,N_1559);
or U2177 (N_2177,N_1603,N_1831);
or U2178 (N_2178,N_1914,N_1674);
or U2179 (N_2179,N_1706,N_1781);
nor U2180 (N_2180,N_1788,N_1726);
xor U2181 (N_2181,N_1821,N_1513);
or U2182 (N_2182,N_1517,N_1623);
or U2183 (N_2183,N_1520,N_1595);
nor U2184 (N_2184,N_1657,N_1935);
or U2185 (N_2185,N_1883,N_1582);
and U2186 (N_2186,N_1791,N_1796);
and U2187 (N_2187,N_1589,N_1626);
nand U2188 (N_2188,N_1802,N_1516);
nand U2189 (N_2189,N_1852,N_1608);
nand U2190 (N_2190,N_1954,N_1729);
xnor U2191 (N_2191,N_1694,N_1754);
nor U2192 (N_2192,N_1968,N_1795);
or U2193 (N_2193,N_1642,N_1966);
and U2194 (N_2194,N_1965,N_1668);
and U2195 (N_2195,N_1702,N_1907);
nor U2196 (N_2196,N_1701,N_1722);
and U2197 (N_2197,N_1615,N_1887);
nor U2198 (N_2198,N_1850,N_1522);
nand U2199 (N_2199,N_1779,N_1962);
nand U2200 (N_2200,N_1725,N_1924);
xnor U2201 (N_2201,N_1752,N_1690);
or U2202 (N_2202,N_1572,N_1501);
nand U2203 (N_2203,N_1672,N_1531);
xnor U2204 (N_2204,N_1720,N_1832);
nor U2205 (N_2205,N_1575,N_1515);
nor U2206 (N_2206,N_1585,N_1957);
and U2207 (N_2207,N_1639,N_1741);
nor U2208 (N_2208,N_1767,N_1716);
nor U2209 (N_2209,N_1561,N_1681);
and U2210 (N_2210,N_1971,N_1990);
nand U2211 (N_2211,N_1621,N_1548);
xor U2212 (N_2212,N_1727,N_1790);
and U2213 (N_2213,N_1801,N_1829);
xor U2214 (N_2214,N_1740,N_1748);
nor U2215 (N_2215,N_1895,N_1596);
nand U2216 (N_2216,N_1985,N_1652);
or U2217 (N_2217,N_1503,N_1853);
and U2218 (N_2218,N_1710,N_1717);
or U2219 (N_2219,N_1785,N_1930);
nor U2220 (N_2220,N_1770,N_1925);
or U2221 (N_2221,N_1817,N_1946);
xor U2222 (N_2222,N_1792,N_1772);
nor U2223 (N_2223,N_1899,N_1973);
nor U2224 (N_2224,N_1552,N_1653);
nor U2225 (N_2225,N_1558,N_1625);
xnor U2226 (N_2226,N_1658,N_1737);
nor U2227 (N_2227,N_1809,N_1678);
nand U2228 (N_2228,N_1982,N_1577);
or U2229 (N_2229,N_1709,N_1712);
nand U2230 (N_2230,N_1934,N_1950);
and U2231 (N_2231,N_1918,N_1988);
and U2232 (N_2232,N_1713,N_1675);
or U2233 (N_2233,N_1735,N_1594);
and U2234 (N_2234,N_1557,N_1768);
nor U2235 (N_2235,N_1518,N_1827);
nand U2236 (N_2236,N_1997,N_1601);
and U2237 (N_2237,N_1868,N_1793);
nor U2238 (N_2238,N_1913,N_1854);
or U2239 (N_2239,N_1719,N_1505);
nand U2240 (N_2240,N_1650,N_1961);
and U2241 (N_2241,N_1955,N_1634);
nand U2242 (N_2242,N_1974,N_1544);
nor U2243 (N_2243,N_1554,N_1543);
nand U2244 (N_2244,N_1881,N_1542);
xor U2245 (N_2245,N_1983,N_1699);
or U2246 (N_2246,N_1514,N_1926);
and U2247 (N_2247,N_1799,N_1549);
or U2248 (N_2248,N_1606,N_1929);
and U2249 (N_2249,N_1695,N_1848);
xnor U2250 (N_2250,N_1897,N_1635);
nand U2251 (N_2251,N_1675,N_1796);
xor U2252 (N_2252,N_1720,N_1671);
and U2253 (N_2253,N_1949,N_1905);
or U2254 (N_2254,N_1579,N_1723);
or U2255 (N_2255,N_1785,N_1911);
nor U2256 (N_2256,N_1940,N_1678);
and U2257 (N_2257,N_1609,N_1695);
and U2258 (N_2258,N_1726,N_1632);
nor U2259 (N_2259,N_1605,N_1570);
or U2260 (N_2260,N_1910,N_1866);
nor U2261 (N_2261,N_1527,N_1675);
and U2262 (N_2262,N_1819,N_1926);
xor U2263 (N_2263,N_1745,N_1627);
nand U2264 (N_2264,N_1938,N_1984);
xor U2265 (N_2265,N_1626,N_1959);
nor U2266 (N_2266,N_1750,N_1878);
or U2267 (N_2267,N_1618,N_1901);
and U2268 (N_2268,N_1523,N_1979);
and U2269 (N_2269,N_1817,N_1872);
and U2270 (N_2270,N_1602,N_1757);
nor U2271 (N_2271,N_1722,N_1870);
nand U2272 (N_2272,N_1767,N_1506);
and U2273 (N_2273,N_1693,N_1781);
nor U2274 (N_2274,N_1809,N_1815);
and U2275 (N_2275,N_1942,N_1615);
and U2276 (N_2276,N_1962,N_1603);
nand U2277 (N_2277,N_1576,N_1540);
nand U2278 (N_2278,N_1544,N_1812);
or U2279 (N_2279,N_1682,N_1506);
nand U2280 (N_2280,N_1737,N_1611);
or U2281 (N_2281,N_1939,N_1500);
nor U2282 (N_2282,N_1528,N_1656);
nand U2283 (N_2283,N_1666,N_1797);
or U2284 (N_2284,N_1720,N_1850);
or U2285 (N_2285,N_1566,N_1671);
or U2286 (N_2286,N_1758,N_1891);
or U2287 (N_2287,N_1731,N_1513);
and U2288 (N_2288,N_1525,N_1789);
and U2289 (N_2289,N_1643,N_1875);
and U2290 (N_2290,N_1587,N_1699);
and U2291 (N_2291,N_1609,N_1517);
nand U2292 (N_2292,N_1905,N_1725);
nor U2293 (N_2293,N_1677,N_1531);
nand U2294 (N_2294,N_1843,N_1809);
nand U2295 (N_2295,N_1933,N_1859);
and U2296 (N_2296,N_1845,N_1595);
nor U2297 (N_2297,N_1709,N_1591);
or U2298 (N_2298,N_1766,N_1779);
nor U2299 (N_2299,N_1843,N_1648);
and U2300 (N_2300,N_1876,N_1537);
nor U2301 (N_2301,N_1741,N_1798);
nand U2302 (N_2302,N_1647,N_1928);
nand U2303 (N_2303,N_1959,N_1800);
nor U2304 (N_2304,N_1591,N_1809);
and U2305 (N_2305,N_1903,N_1542);
xor U2306 (N_2306,N_1998,N_1889);
and U2307 (N_2307,N_1552,N_1650);
nor U2308 (N_2308,N_1570,N_1844);
or U2309 (N_2309,N_1826,N_1835);
and U2310 (N_2310,N_1524,N_1798);
xor U2311 (N_2311,N_1673,N_1983);
nand U2312 (N_2312,N_1653,N_1716);
nand U2313 (N_2313,N_1803,N_1973);
or U2314 (N_2314,N_1807,N_1917);
nand U2315 (N_2315,N_1805,N_1546);
and U2316 (N_2316,N_1751,N_1678);
xnor U2317 (N_2317,N_1834,N_1910);
or U2318 (N_2318,N_1783,N_1840);
and U2319 (N_2319,N_1657,N_1785);
or U2320 (N_2320,N_1792,N_1935);
nor U2321 (N_2321,N_1527,N_1563);
nor U2322 (N_2322,N_1736,N_1683);
nor U2323 (N_2323,N_1871,N_1602);
nand U2324 (N_2324,N_1710,N_1915);
or U2325 (N_2325,N_1957,N_1958);
nor U2326 (N_2326,N_1547,N_1943);
or U2327 (N_2327,N_1662,N_1828);
nand U2328 (N_2328,N_1788,N_1570);
or U2329 (N_2329,N_1515,N_1927);
nand U2330 (N_2330,N_1578,N_1992);
or U2331 (N_2331,N_1858,N_1922);
or U2332 (N_2332,N_1899,N_1517);
and U2333 (N_2333,N_1778,N_1819);
or U2334 (N_2334,N_1552,N_1573);
or U2335 (N_2335,N_1847,N_1645);
and U2336 (N_2336,N_1755,N_1987);
nand U2337 (N_2337,N_1570,N_1511);
or U2338 (N_2338,N_1792,N_1679);
and U2339 (N_2339,N_1584,N_1913);
xnor U2340 (N_2340,N_1750,N_1800);
xnor U2341 (N_2341,N_1976,N_1607);
or U2342 (N_2342,N_1966,N_1500);
nand U2343 (N_2343,N_1902,N_1776);
or U2344 (N_2344,N_1590,N_1824);
and U2345 (N_2345,N_1799,N_1844);
and U2346 (N_2346,N_1703,N_1639);
nor U2347 (N_2347,N_1558,N_1747);
xor U2348 (N_2348,N_1664,N_1967);
nor U2349 (N_2349,N_1504,N_1854);
and U2350 (N_2350,N_1951,N_1716);
xnor U2351 (N_2351,N_1943,N_1881);
and U2352 (N_2352,N_1681,N_1528);
nor U2353 (N_2353,N_1651,N_1703);
and U2354 (N_2354,N_1769,N_1853);
nor U2355 (N_2355,N_1904,N_1851);
or U2356 (N_2356,N_1771,N_1927);
and U2357 (N_2357,N_1646,N_1502);
nand U2358 (N_2358,N_1690,N_1593);
and U2359 (N_2359,N_1560,N_1613);
or U2360 (N_2360,N_1692,N_1589);
nand U2361 (N_2361,N_1933,N_1988);
nor U2362 (N_2362,N_1509,N_1958);
nor U2363 (N_2363,N_1673,N_1998);
and U2364 (N_2364,N_1839,N_1798);
or U2365 (N_2365,N_1602,N_1766);
nand U2366 (N_2366,N_1820,N_1831);
nor U2367 (N_2367,N_1805,N_1711);
xor U2368 (N_2368,N_1687,N_1793);
nor U2369 (N_2369,N_1749,N_1685);
nor U2370 (N_2370,N_1809,N_1581);
nand U2371 (N_2371,N_1928,N_1672);
nand U2372 (N_2372,N_1509,N_1908);
nor U2373 (N_2373,N_1844,N_1865);
nand U2374 (N_2374,N_1958,N_1788);
or U2375 (N_2375,N_1884,N_1524);
or U2376 (N_2376,N_1535,N_1664);
nor U2377 (N_2377,N_1788,N_1535);
or U2378 (N_2378,N_1654,N_1518);
nand U2379 (N_2379,N_1700,N_1548);
xor U2380 (N_2380,N_1693,N_1923);
and U2381 (N_2381,N_1961,N_1918);
and U2382 (N_2382,N_1960,N_1889);
xnor U2383 (N_2383,N_1736,N_1902);
nand U2384 (N_2384,N_1720,N_1726);
and U2385 (N_2385,N_1808,N_1613);
or U2386 (N_2386,N_1773,N_1890);
nand U2387 (N_2387,N_1638,N_1811);
nand U2388 (N_2388,N_1557,N_1586);
xor U2389 (N_2389,N_1690,N_1708);
nor U2390 (N_2390,N_1791,N_1635);
or U2391 (N_2391,N_1687,N_1940);
and U2392 (N_2392,N_1866,N_1677);
xnor U2393 (N_2393,N_1774,N_1569);
or U2394 (N_2394,N_1716,N_1663);
nand U2395 (N_2395,N_1946,N_1606);
and U2396 (N_2396,N_1703,N_1511);
and U2397 (N_2397,N_1539,N_1677);
nand U2398 (N_2398,N_1782,N_1722);
nor U2399 (N_2399,N_1792,N_1838);
nor U2400 (N_2400,N_1792,N_1651);
or U2401 (N_2401,N_1909,N_1842);
nand U2402 (N_2402,N_1568,N_1561);
xor U2403 (N_2403,N_1579,N_1522);
xor U2404 (N_2404,N_1977,N_1918);
and U2405 (N_2405,N_1862,N_1991);
nor U2406 (N_2406,N_1778,N_1735);
xor U2407 (N_2407,N_1720,N_1695);
and U2408 (N_2408,N_1921,N_1890);
and U2409 (N_2409,N_1632,N_1576);
and U2410 (N_2410,N_1641,N_1601);
nor U2411 (N_2411,N_1916,N_1777);
or U2412 (N_2412,N_1543,N_1809);
and U2413 (N_2413,N_1852,N_1754);
or U2414 (N_2414,N_1787,N_1836);
nand U2415 (N_2415,N_1936,N_1530);
nand U2416 (N_2416,N_1706,N_1762);
and U2417 (N_2417,N_1628,N_1507);
or U2418 (N_2418,N_1849,N_1633);
nand U2419 (N_2419,N_1988,N_1923);
nand U2420 (N_2420,N_1564,N_1755);
nand U2421 (N_2421,N_1828,N_1636);
or U2422 (N_2422,N_1889,N_1939);
and U2423 (N_2423,N_1867,N_1623);
and U2424 (N_2424,N_1881,N_1639);
and U2425 (N_2425,N_1908,N_1805);
or U2426 (N_2426,N_1872,N_1695);
nor U2427 (N_2427,N_1530,N_1869);
nor U2428 (N_2428,N_1881,N_1742);
nand U2429 (N_2429,N_1590,N_1881);
and U2430 (N_2430,N_1949,N_1546);
nand U2431 (N_2431,N_1922,N_1603);
nand U2432 (N_2432,N_1923,N_1972);
or U2433 (N_2433,N_1542,N_1848);
and U2434 (N_2434,N_1990,N_1655);
nor U2435 (N_2435,N_1938,N_1636);
nor U2436 (N_2436,N_1861,N_1854);
or U2437 (N_2437,N_1887,N_1792);
nor U2438 (N_2438,N_1615,N_1738);
or U2439 (N_2439,N_1916,N_1895);
and U2440 (N_2440,N_1997,N_1731);
nor U2441 (N_2441,N_1874,N_1781);
nor U2442 (N_2442,N_1872,N_1820);
or U2443 (N_2443,N_1541,N_1600);
nand U2444 (N_2444,N_1669,N_1661);
nand U2445 (N_2445,N_1753,N_1614);
or U2446 (N_2446,N_1890,N_1794);
or U2447 (N_2447,N_1962,N_1667);
or U2448 (N_2448,N_1628,N_1957);
nor U2449 (N_2449,N_1561,N_1645);
nand U2450 (N_2450,N_1559,N_1847);
nand U2451 (N_2451,N_1865,N_1684);
xnor U2452 (N_2452,N_1571,N_1982);
nor U2453 (N_2453,N_1958,N_1960);
or U2454 (N_2454,N_1982,N_1896);
nor U2455 (N_2455,N_1928,N_1529);
or U2456 (N_2456,N_1932,N_1552);
or U2457 (N_2457,N_1991,N_1951);
nor U2458 (N_2458,N_1833,N_1534);
or U2459 (N_2459,N_1778,N_1508);
or U2460 (N_2460,N_1784,N_1641);
and U2461 (N_2461,N_1904,N_1696);
nand U2462 (N_2462,N_1574,N_1797);
and U2463 (N_2463,N_1638,N_1898);
and U2464 (N_2464,N_1768,N_1733);
and U2465 (N_2465,N_1892,N_1526);
xor U2466 (N_2466,N_1586,N_1576);
and U2467 (N_2467,N_1893,N_1931);
or U2468 (N_2468,N_1544,N_1678);
and U2469 (N_2469,N_1858,N_1636);
and U2470 (N_2470,N_1545,N_1680);
or U2471 (N_2471,N_1933,N_1736);
xor U2472 (N_2472,N_1884,N_1771);
and U2473 (N_2473,N_1632,N_1516);
or U2474 (N_2474,N_1578,N_1889);
nand U2475 (N_2475,N_1529,N_1871);
xor U2476 (N_2476,N_1597,N_1925);
nand U2477 (N_2477,N_1799,N_1629);
nor U2478 (N_2478,N_1797,N_1940);
or U2479 (N_2479,N_1802,N_1682);
or U2480 (N_2480,N_1800,N_1732);
or U2481 (N_2481,N_1805,N_1796);
nand U2482 (N_2482,N_1848,N_1954);
and U2483 (N_2483,N_1998,N_1846);
or U2484 (N_2484,N_1638,N_1863);
nor U2485 (N_2485,N_1522,N_1559);
nor U2486 (N_2486,N_1747,N_1775);
and U2487 (N_2487,N_1834,N_1535);
and U2488 (N_2488,N_1840,N_1873);
nor U2489 (N_2489,N_1956,N_1806);
and U2490 (N_2490,N_1974,N_1983);
and U2491 (N_2491,N_1617,N_1807);
nor U2492 (N_2492,N_1923,N_1717);
or U2493 (N_2493,N_1924,N_1687);
nor U2494 (N_2494,N_1791,N_1992);
nand U2495 (N_2495,N_1584,N_1747);
nand U2496 (N_2496,N_1785,N_1969);
xor U2497 (N_2497,N_1913,N_1923);
or U2498 (N_2498,N_1940,N_1820);
or U2499 (N_2499,N_1913,N_1674);
nor U2500 (N_2500,N_2433,N_2340);
nand U2501 (N_2501,N_2106,N_2251);
nand U2502 (N_2502,N_2300,N_2082);
and U2503 (N_2503,N_2035,N_2037);
or U2504 (N_2504,N_2395,N_2234);
or U2505 (N_2505,N_2159,N_2336);
and U2506 (N_2506,N_2352,N_2182);
nand U2507 (N_2507,N_2392,N_2252);
and U2508 (N_2508,N_2412,N_2342);
and U2509 (N_2509,N_2070,N_2435);
or U2510 (N_2510,N_2273,N_2148);
nand U2511 (N_2511,N_2371,N_2348);
nand U2512 (N_2512,N_2177,N_2394);
and U2513 (N_2513,N_2221,N_2230);
and U2514 (N_2514,N_2350,N_2289);
and U2515 (N_2515,N_2466,N_2421);
nand U2516 (N_2516,N_2359,N_2411);
and U2517 (N_2517,N_2163,N_2147);
nor U2518 (N_2518,N_2271,N_2344);
or U2519 (N_2519,N_2017,N_2038);
nor U2520 (N_2520,N_2079,N_2387);
or U2521 (N_2521,N_2233,N_2422);
and U2522 (N_2522,N_2290,N_2124);
nand U2523 (N_2523,N_2307,N_2235);
nand U2524 (N_2524,N_2255,N_2055);
and U2525 (N_2525,N_2004,N_2149);
xnor U2526 (N_2526,N_2073,N_2204);
nor U2527 (N_2527,N_2214,N_2025);
nor U2528 (N_2528,N_2047,N_2226);
nor U2529 (N_2529,N_2283,N_2023);
nand U2530 (N_2530,N_2091,N_2150);
xnor U2531 (N_2531,N_2012,N_2312);
and U2532 (N_2532,N_2479,N_2044);
or U2533 (N_2533,N_2198,N_2143);
nand U2534 (N_2534,N_2168,N_2006);
or U2535 (N_2535,N_2164,N_2078);
nor U2536 (N_2536,N_2239,N_2451);
or U2537 (N_2537,N_2122,N_2410);
or U2538 (N_2538,N_2133,N_2386);
nand U2539 (N_2539,N_2454,N_2272);
or U2540 (N_2540,N_2444,N_2361);
and U2541 (N_2541,N_2123,N_2297);
or U2542 (N_2542,N_2045,N_2259);
nand U2543 (N_2543,N_2116,N_2327);
nand U2544 (N_2544,N_2110,N_2362);
and U2545 (N_2545,N_2207,N_2155);
xnor U2546 (N_2546,N_2469,N_2403);
nor U2547 (N_2547,N_2321,N_2247);
and U2548 (N_2548,N_2048,N_2434);
nor U2549 (N_2549,N_2354,N_2248);
or U2550 (N_2550,N_2036,N_2274);
xnor U2551 (N_2551,N_2460,N_2102);
xor U2552 (N_2552,N_2069,N_2208);
or U2553 (N_2553,N_2470,N_2463);
nand U2554 (N_2554,N_2209,N_2383);
nand U2555 (N_2555,N_2351,N_2018);
nor U2556 (N_2556,N_2313,N_2211);
xnor U2557 (N_2557,N_2330,N_2139);
and U2558 (N_2558,N_2086,N_2397);
nand U2559 (N_2559,N_2447,N_2294);
and U2560 (N_2560,N_2389,N_2085);
or U2561 (N_2561,N_2146,N_2314);
nand U2562 (N_2562,N_2431,N_2326);
and U2563 (N_2563,N_2173,N_2333);
nor U2564 (N_2564,N_2152,N_2345);
and U2565 (N_2565,N_2189,N_2162);
nor U2566 (N_2566,N_2497,N_2246);
xor U2567 (N_2567,N_2476,N_2436);
or U2568 (N_2568,N_2353,N_2167);
nand U2569 (N_2569,N_2065,N_2192);
nor U2570 (N_2570,N_2212,N_2416);
or U2571 (N_2571,N_2032,N_2420);
nor U2572 (N_2572,N_2130,N_2370);
nor U2573 (N_2573,N_2325,N_2275);
nor U2574 (N_2574,N_2054,N_2426);
nor U2575 (N_2575,N_2440,N_2128);
or U2576 (N_2576,N_2135,N_2390);
nor U2577 (N_2577,N_2428,N_2196);
and U2578 (N_2578,N_2224,N_2424);
nor U2579 (N_2579,N_2015,N_2474);
or U2580 (N_2580,N_2278,N_2415);
and U2581 (N_2581,N_2202,N_2066);
and U2582 (N_2582,N_2222,N_2378);
or U2583 (N_2583,N_2220,N_2429);
and U2584 (N_2584,N_2276,N_2225);
or U2585 (N_2585,N_2269,N_2254);
or U2586 (N_2586,N_2430,N_2174);
and U2587 (N_2587,N_2075,N_2179);
nor U2588 (N_2588,N_2042,N_2197);
or U2589 (N_2589,N_2104,N_2481);
and U2590 (N_2590,N_2093,N_2375);
and U2591 (N_2591,N_2095,N_2108);
and U2592 (N_2592,N_2494,N_2046);
xnor U2593 (N_2593,N_2291,N_2028);
or U2594 (N_2594,N_2459,N_2367);
and U2595 (N_2595,N_2030,N_2107);
nand U2596 (N_2596,N_2134,N_2059);
or U2597 (N_2597,N_2228,N_2009);
nand U2598 (N_2598,N_2471,N_2425);
nor U2599 (N_2599,N_2153,N_2329);
nand U2600 (N_2600,N_2257,N_2492);
nand U2601 (N_2601,N_2049,N_2306);
or U2602 (N_2602,N_2323,N_2231);
or U2603 (N_2603,N_2385,N_2029);
or U2604 (N_2604,N_2475,N_2005);
nor U2605 (N_2605,N_2285,N_2360);
nand U2606 (N_2606,N_2304,N_2478);
xnor U2607 (N_2607,N_2281,N_2423);
or U2608 (N_2608,N_2058,N_2244);
xor U2609 (N_2609,N_2264,N_2232);
and U2610 (N_2610,N_2339,N_2437);
xor U2611 (N_2611,N_2310,N_2453);
or U2612 (N_2612,N_2356,N_2190);
and U2613 (N_2613,N_2172,N_2080);
nand U2614 (N_2614,N_2465,N_2268);
and U2615 (N_2615,N_2229,N_2136);
xnor U2616 (N_2616,N_2185,N_2076);
nor U2617 (N_2617,N_2081,N_2499);
nor U2618 (N_2618,N_2187,N_2142);
or U2619 (N_2619,N_2068,N_2284);
and U2620 (N_2620,N_2145,N_2347);
nor U2621 (N_2621,N_2237,N_2199);
nand U2622 (N_2622,N_2299,N_2002);
xor U2623 (N_2623,N_2210,N_2438);
or U2624 (N_2624,N_2118,N_2485);
nor U2625 (N_2625,N_2166,N_2227);
nand U2626 (N_2626,N_2477,N_2249);
nand U2627 (N_2627,N_2357,N_2188);
or U2628 (N_2628,N_2315,N_2488);
nand U2629 (N_2629,N_2089,N_2379);
nand U2630 (N_2630,N_2033,N_2490);
nor U2631 (N_2631,N_2238,N_2014);
and U2632 (N_2632,N_2468,N_2417);
and U2633 (N_2633,N_2358,N_2279);
nor U2634 (N_2634,N_2200,N_2169);
or U2635 (N_2635,N_2303,N_2282);
nand U2636 (N_2636,N_2098,N_2219);
or U2637 (N_2637,N_2373,N_2090);
and U2638 (N_2638,N_2399,N_2302);
nor U2639 (N_2639,N_2132,N_2452);
or U2640 (N_2640,N_2262,N_2464);
and U2641 (N_2641,N_2366,N_2482);
nor U2642 (N_2642,N_2092,N_2053);
nand U2643 (N_2643,N_2057,N_2137);
nand U2644 (N_2644,N_2393,N_2376);
nand U2645 (N_2645,N_2043,N_2140);
xor U2646 (N_2646,N_2217,N_2171);
or U2647 (N_2647,N_2473,N_2398);
xor U2648 (N_2648,N_2380,N_2496);
and U2649 (N_2649,N_2337,N_2318);
nor U2650 (N_2650,N_2016,N_2309);
or U2651 (N_2651,N_2266,N_2215);
nand U2652 (N_2652,N_2181,N_2121);
and U2653 (N_2653,N_2296,N_2277);
nand U2654 (N_2654,N_2462,N_2286);
nor U2655 (N_2655,N_2154,N_2317);
or U2656 (N_2656,N_2408,N_2064);
xor U2657 (N_2657,N_2405,N_2129);
and U2658 (N_2658,N_2158,N_2372);
and U2659 (N_2659,N_2186,N_2141);
xor U2660 (N_2660,N_2498,N_2034);
nand U2661 (N_2661,N_2193,N_2074);
nor U2662 (N_2662,N_2083,N_2419);
nand U2663 (N_2663,N_2295,N_2261);
nand U2664 (N_2664,N_2040,N_2414);
or U2665 (N_2665,N_2486,N_2195);
nand U2666 (N_2666,N_2381,N_2191);
or U2667 (N_2667,N_2156,N_2472);
and U2668 (N_2668,N_2404,N_2250);
nand U2669 (N_2669,N_2112,N_2176);
nand U2670 (N_2670,N_2280,N_2368);
or U2671 (N_2671,N_2445,N_2391);
or U2672 (N_2672,N_2256,N_2242);
or U2673 (N_2673,N_2432,N_2062);
nand U2674 (N_2674,N_2061,N_2401);
nand U2675 (N_2675,N_2003,N_2396);
and U2676 (N_2676,N_2346,N_2170);
nor U2677 (N_2677,N_2223,N_2493);
nand U2678 (N_2678,N_2292,N_2388);
or U2679 (N_2679,N_2001,N_2111);
nand U2680 (N_2680,N_2157,N_2022);
nor U2681 (N_2681,N_2365,N_2206);
nor U2682 (N_2682,N_2427,N_2100);
nand U2683 (N_2683,N_2160,N_2105);
and U2684 (N_2684,N_2241,N_2087);
and U2685 (N_2685,N_2467,N_2101);
and U2686 (N_2686,N_2126,N_2439);
nand U2687 (N_2687,N_2161,N_2461);
and U2688 (N_2688,N_2041,N_2010);
nor U2689 (N_2689,N_2039,N_2406);
nand U2690 (N_2690,N_2260,N_2096);
nor U2691 (N_2691,N_2288,N_2484);
nor U2692 (N_2692,N_2243,N_2443);
nor U2693 (N_2693,N_2265,N_2343);
nor U2694 (N_2694,N_2099,N_2109);
and U2695 (N_2695,N_2407,N_2021);
or U2696 (N_2696,N_2165,N_2216);
and U2697 (N_2697,N_2013,N_2119);
and U2698 (N_2698,N_2384,N_2322);
or U2699 (N_2699,N_2409,N_2311);
or U2700 (N_2700,N_2258,N_2131);
or U2701 (N_2701,N_2495,N_2263);
or U2702 (N_2702,N_2301,N_2213);
nand U2703 (N_2703,N_2450,N_2270);
nand U2704 (N_2704,N_2374,N_2201);
or U2705 (N_2705,N_2008,N_2319);
xor U2706 (N_2706,N_2245,N_2151);
nor U2707 (N_2707,N_2298,N_2364);
or U2708 (N_2708,N_2338,N_2178);
nor U2709 (N_2709,N_2019,N_2458);
nor U2710 (N_2710,N_2056,N_2114);
nand U2711 (N_2711,N_2324,N_2253);
or U2712 (N_2712,N_2400,N_2449);
and U2713 (N_2713,N_2355,N_2489);
xnor U2714 (N_2714,N_2455,N_2144);
or U2715 (N_2715,N_2402,N_2052);
and U2716 (N_2716,N_2138,N_2382);
nor U2717 (N_2717,N_2334,N_2335);
or U2718 (N_2718,N_2377,N_2094);
and U2719 (N_2719,N_2287,N_2349);
nor U2720 (N_2720,N_2483,N_2088);
and U2721 (N_2721,N_2442,N_2341);
or U2722 (N_2722,N_2369,N_2418);
and U2723 (N_2723,N_2316,N_2125);
nor U2724 (N_2724,N_2175,N_2456);
nor U2725 (N_2725,N_2026,N_2320);
nand U2726 (N_2726,N_2077,N_2060);
nand U2727 (N_2727,N_2084,N_2127);
nor U2728 (N_2728,N_2180,N_2240);
nand U2729 (N_2729,N_2308,N_2103);
nand U2730 (N_2730,N_2011,N_2050);
or U2731 (N_2731,N_2120,N_2448);
and U2732 (N_2732,N_2203,N_2183);
xor U2733 (N_2733,N_2000,N_2063);
or U2734 (N_2734,N_2024,N_2007);
nand U2735 (N_2735,N_2267,N_2027);
or U2736 (N_2736,N_2117,N_2331);
nor U2737 (N_2737,N_2480,N_2446);
or U2738 (N_2738,N_2457,N_2020);
or U2739 (N_2739,N_2332,N_2194);
and U2740 (N_2740,N_2067,N_2363);
or U2741 (N_2741,N_2115,N_2236);
nor U2742 (N_2742,N_2328,N_2218);
xor U2743 (N_2743,N_2305,N_2184);
nor U2744 (N_2744,N_2413,N_2072);
xnor U2745 (N_2745,N_2097,N_2071);
nand U2746 (N_2746,N_2051,N_2487);
or U2747 (N_2747,N_2441,N_2293);
or U2748 (N_2748,N_2491,N_2113);
and U2749 (N_2749,N_2205,N_2031);
and U2750 (N_2750,N_2390,N_2157);
or U2751 (N_2751,N_2434,N_2014);
nor U2752 (N_2752,N_2283,N_2184);
nand U2753 (N_2753,N_2396,N_2418);
nor U2754 (N_2754,N_2472,N_2044);
nand U2755 (N_2755,N_2125,N_2307);
or U2756 (N_2756,N_2313,N_2391);
xor U2757 (N_2757,N_2367,N_2421);
or U2758 (N_2758,N_2275,N_2069);
and U2759 (N_2759,N_2226,N_2001);
and U2760 (N_2760,N_2108,N_2246);
nor U2761 (N_2761,N_2412,N_2240);
and U2762 (N_2762,N_2240,N_2471);
and U2763 (N_2763,N_2180,N_2489);
or U2764 (N_2764,N_2414,N_2499);
xor U2765 (N_2765,N_2009,N_2422);
and U2766 (N_2766,N_2397,N_2333);
and U2767 (N_2767,N_2334,N_2253);
nor U2768 (N_2768,N_2054,N_2095);
and U2769 (N_2769,N_2269,N_2278);
xnor U2770 (N_2770,N_2234,N_2445);
nand U2771 (N_2771,N_2190,N_2415);
and U2772 (N_2772,N_2152,N_2476);
and U2773 (N_2773,N_2269,N_2315);
nand U2774 (N_2774,N_2331,N_2216);
nor U2775 (N_2775,N_2401,N_2064);
or U2776 (N_2776,N_2179,N_2209);
nor U2777 (N_2777,N_2437,N_2445);
and U2778 (N_2778,N_2447,N_2236);
nor U2779 (N_2779,N_2381,N_2113);
nor U2780 (N_2780,N_2272,N_2075);
nor U2781 (N_2781,N_2157,N_2179);
nand U2782 (N_2782,N_2488,N_2359);
and U2783 (N_2783,N_2102,N_2470);
and U2784 (N_2784,N_2370,N_2198);
nor U2785 (N_2785,N_2198,N_2210);
nand U2786 (N_2786,N_2392,N_2490);
or U2787 (N_2787,N_2232,N_2256);
and U2788 (N_2788,N_2417,N_2476);
nor U2789 (N_2789,N_2381,N_2058);
xnor U2790 (N_2790,N_2237,N_2431);
nand U2791 (N_2791,N_2371,N_2430);
nor U2792 (N_2792,N_2486,N_2118);
nor U2793 (N_2793,N_2041,N_2015);
nand U2794 (N_2794,N_2401,N_2118);
and U2795 (N_2795,N_2318,N_2395);
and U2796 (N_2796,N_2173,N_2142);
nand U2797 (N_2797,N_2371,N_2489);
nand U2798 (N_2798,N_2149,N_2422);
and U2799 (N_2799,N_2490,N_2132);
and U2800 (N_2800,N_2425,N_2456);
nand U2801 (N_2801,N_2355,N_2047);
or U2802 (N_2802,N_2305,N_2023);
nand U2803 (N_2803,N_2237,N_2474);
xnor U2804 (N_2804,N_2452,N_2249);
or U2805 (N_2805,N_2154,N_2244);
nor U2806 (N_2806,N_2071,N_2142);
nand U2807 (N_2807,N_2289,N_2453);
xnor U2808 (N_2808,N_2378,N_2265);
and U2809 (N_2809,N_2206,N_2286);
nor U2810 (N_2810,N_2467,N_2401);
nor U2811 (N_2811,N_2185,N_2412);
nor U2812 (N_2812,N_2352,N_2107);
and U2813 (N_2813,N_2306,N_2308);
or U2814 (N_2814,N_2296,N_2233);
xnor U2815 (N_2815,N_2183,N_2139);
nand U2816 (N_2816,N_2000,N_2201);
nor U2817 (N_2817,N_2290,N_2419);
or U2818 (N_2818,N_2141,N_2324);
nor U2819 (N_2819,N_2284,N_2328);
nand U2820 (N_2820,N_2497,N_2158);
nand U2821 (N_2821,N_2468,N_2090);
or U2822 (N_2822,N_2121,N_2073);
nand U2823 (N_2823,N_2276,N_2433);
nand U2824 (N_2824,N_2029,N_2369);
or U2825 (N_2825,N_2264,N_2186);
nand U2826 (N_2826,N_2415,N_2226);
nand U2827 (N_2827,N_2122,N_2414);
and U2828 (N_2828,N_2064,N_2379);
or U2829 (N_2829,N_2221,N_2342);
and U2830 (N_2830,N_2429,N_2293);
nand U2831 (N_2831,N_2204,N_2476);
and U2832 (N_2832,N_2216,N_2032);
or U2833 (N_2833,N_2105,N_2476);
nor U2834 (N_2834,N_2106,N_2353);
nand U2835 (N_2835,N_2116,N_2064);
and U2836 (N_2836,N_2335,N_2441);
and U2837 (N_2837,N_2347,N_2215);
or U2838 (N_2838,N_2221,N_2288);
and U2839 (N_2839,N_2274,N_2298);
nor U2840 (N_2840,N_2099,N_2436);
nand U2841 (N_2841,N_2326,N_2248);
nor U2842 (N_2842,N_2178,N_2004);
nand U2843 (N_2843,N_2307,N_2318);
nor U2844 (N_2844,N_2203,N_2171);
nand U2845 (N_2845,N_2121,N_2279);
and U2846 (N_2846,N_2259,N_2016);
and U2847 (N_2847,N_2319,N_2484);
or U2848 (N_2848,N_2278,N_2051);
and U2849 (N_2849,N_2235,N_2207);
nor U2850 (N_2850,N_2153,N_2171);
nor U2851 (N_2851,N_2183,N_2191);
xor U2852 (N_2852,N_2318,N_2238);
nand U2853 (N_2853,N_2012,N_2083);
xnor U2854 (N_2854,N_2420,N_2185);
or U2855 (N_2855,N_2108,N_2267);
nand U2856 (N_2856,N_2432,N_2033);
or U2857 (N_2857,N_2348,N_2139);
or U2858 (N_2858,N_2049,N_2119);
and U2859 (N_2859,N_2355,N_2229);
nand U2860 (N_2860,N_2460,N_2196);
and U2861 (N_2861,N_2204,N_2436);
nor U2862 (N_2862,N_2001,N_2263);
and U2863 (N_2863,N_2031,N_2339);
xor U2864 (N_2864,N_2084,N_2025);
nand U2865 (N_2865,N_2092,N_2105);
or U2866 (N_2866,N_2205,N_2300);
or U2867 (N_2867,N_2487,N_2234);
nand U2868 (N_2868,N_2034,N_2179);
xnor U2869 (N_2869,N_2314,N_2487);
or U2870 (N_2870,N_2127,N_2402);
nor U2871 (N_2871,N_2303,N_2224);
and U2872 (N_2872,N_2129,N_2020);
nand U2873 (N_2873,N_2010,N_2021);
nor U2874 (N_2874,N_2396,N_2494);
or U2875 (N_2875,N_2445,N_2215);
nand U2876 (N_2876,N_2006,N_2303);
nor U2877 (N_2877,N_2320,N_2119);
or U2878 (N_2878,N_2488,N_2343);
nor U2879 (N_2879,N_2395,N_2211);
nor U2880 (N_2880,N_2363,N_2096);
nor U2881 (N_2881,N_2155,N_2289);
and U2882 (N_2882,N_2253,N_2477);
or U2883 (N_2883,N_2410,N_2230);
nor U2884 (N_2884,N_2367,N_2132);
xor U2885 (N_2885,N_2458,N_2247);
or U2886 (N_2886,N_2116,N_2093);
nor U2887 (N_2887,N_2458,N_2428);
nor U2888 (N_2888,N_2457,N_2234);
nand U2889 (N_2889,N_2029,N_2240);
nor U2890 (N_2890,N_2273,N_2260);
nand U2891 (N_2891,N_2011,N_2004);
and U2892 (N_2892,N_2435,N_2320);
nor U2893 (N_2893,N_2001,N_2252);
nand U2894 (N_2894,N_2255,N_2270);
or U2895 (N_2895,N_2234,N_2212);
or U2896 (N_2896,N_2322,N_2421);
nand U2897 (N_2897,N_2182,N_2027);
nor U2898 (N_2898,N_2450,N_2148);
or U2899 (N_2899,N_2412,N_2396);
or U2900 (N_2900,N_2437,N_2400);
xor U2901 (N_2901,N_2247,N_2304);
or U2902 (N_2902,N_2243,N_2332);
nand U2903 (N_2903,N_2186,N_2070);
nor U2904 (N_2904,N_2393,N_2341);
or U2905 (N_2905,N_2108,N_2145);
xor U2906 (N_2906,N_2064,N_2044);
and U2907 (N_2907,N_2275,N_2140);
xnor U2908 (N_2908,N_2227,N_2245);
nand U2909 (N_2909,N_2242,N_2294);
nand U2910 (N_2910,N_2393,N_2450);
and U2911 (N_2911,N_2461,N_2353);
or U2912 (N_2912,N_2435,N_2374);
nor U2913 (N_2913,N_2125,N_2177);
or U2914 (N_2914,N_2020,N_2207);
and U2915 (N_2915,N_2183,N_2367);
nor U2916 (N_2916,N_2181,N_2109);
and U2917 (N_2917,N_2417,N_2475);
xnor U2918 (N_2918,N_2171,N_2214);
nand U2919 (N_2919,N_2400,N_2489);
nor U2920 (N_2920,N_2208,N_2050);
xnor U2921 (N_2921,N_2019,N_2195);
and U2922 (N_2922,N_2027,N_2460);
xor U2923 (N_2923,N_2498,N_2302);
or U2924 (N_2924,N_2278,N_2184);
and U2925 (N_2925,N_2208,N_2455);
and U2926 (N_2926,N_2229,N_2324);
and U2927 (N_2927,N_2024,N_2384);
nor U2928 (N_2928,N_2442,N_2134);
and U2929 (N_2929,N_2323,N_2314);
xor U2930 (N_2930,N_2059,N_2077);
xnor U2931 (N_2931,N_2242,N_2219);
and U2932 (N_2932,N_2152,N_2433);
and U2933 (N_2933,N_2329,N_2385);
or U2934 (N_2934,N_2478,N_2343);
nand U2935 (N_2935,N_2276,N_2331);
nor U2936 (N_2936,N_2325,N_2310);
or U2937 (N_2937,N_2475,N_2314);
or U2938 (N_2938,N_2449,N_2175);
nor U2939 (N_2939,N_2261,N_2033);
and U2940 (N_2940,N_2202,N_2382);
xnor U2941 (N_2941,N_2234,N_2383);
and U2942 (N_2942,N_2257,N_2115);
nand U2943 (N_2943,N_2032,N_2013);
nand U2944 (N_2944,N_2332,N_2431);
xnor U2945 (N_2945,N_2017,N_2012);
nand U2946 (N_2946,N_2435,N_2248);
xnor U2947 (N_2947,N_2011,N_2353);
or U2948 (N_2948,N_2319,N_2148);
nor U2949 (N_2949,N_2282,N_2412);
or U2950 (N_2950,N_2041,N_2276);
or U2951 (N_2951,N_2405,N_2453);
nor U2952 (N_2952,N_2400,N_2250);
nor U2953 (N_2953,N_2150,N_2474);
nand U2954 (N_2954,N_2495,N_2038);
nand U2955 (N_2955,N_2361,N_2026);
nor U2956 (N_2956,N_2150,N_2196);
and U2957 (N_2957,N_2075,N_2243);
and U2958 (N_2958,N_2306,N_2331);
or U2959 (N_2959,N_2357,N_2376);
nor U2960 (N_2960,N_2241,N_2109);
nor U2961 (N_2961,N_2339,N_2459);
nand U2962 (N_2962,N_2042,N_2049);
nor U2963 (N_2963,N_2148,N_2443);
or U2964 (N_2964,N_2197,N_2122);
nand U2965 (N_2965,N_2070,N_2086);
nand U2966 (N_2966,N_2304,N_2366);
and U2967 (N_2967,N_2413,N_2330);
nor U2968 (N_2968,N_2498,N_2410);
xnor U2969 (N_2969,N_2184,N_2101);
nand U2970 (N_2970,N_2112,N_2249);
nor U2971 (N_2971,N_2052,N_2281);
or U2972 (N_2972,N_2371,N_2039);
and U2973 (N_2973,N_2435,N_2255);
or U2974 (N_2974,N_2002,N_2482);
and U2975 (N_2975,N_2290,N_2313);
and U2976 (N_2976,N_2476,N_2076);
and U2977 (N_2977,N_2032,N_2077);
nor U2978 (N_2978,N_2151,N_2098);
or U2979 (N_2979,N_2230,N_2197);
nand U2980 (N_2980,N_2488,N_2004);
and U2981 (N_2981,N_2200,N_2252);
nor U2982 (N_2982,N_2014,N_2057);
xnor U2983 (N_2983,N_2096,N_2014);
or U2984 (N_2984,N_2205,N_2004);
and U2985 (N_2985,N_2483,N_2040);
or U2986 (N_2986,N_2481,N_2366);
or U2987 (N_2987,N_2098,N_2398);
or U2988 (N_2988,N_2293,N_2433);
xor U2989 (N_2989,N_2265,N_2324);
or U2990 (N_2990,N_2003,N_2130);
or U2991 (N_2991,N_2471,N_2206);
or U2992 (N_2992,N_2242,N_2012);
and U2993 (N_2993,N_2465,N_2199);
nor U2994 (N_2994,N_2214,N_2172);
or U2995 (N_2995,N_2212,N_2287);
nand U2996 (N_2996,N_2416,N_2240);
nand U2997 (N_2997,N_2251,N_2102);
or U2998 (N_2998,N_2248,N_2398);
or U2999 (N_2999,N_2024,N_2401);
xor U3000 (N_3000,N_2641,N_2821);
and U3001 (N_3001,N_2796,N_2783);
nor U3002 (N_3002,N_2964,N_2713);
nor U3003 (N_3003,N_2866,N_2663);
or U3004 (N_3004,N_2726,N_2507);
or U3005 (N_3005,N_2715,N_2577);
nor U3006 (N_3006,N_2583,N_2573);
or U3007 (N_3007,N_2798,N_2929);
nand U3008 (N_3008,N_2722,N_2839);
xnor U3009 (N_3009,N_2648,N_2865);
and U3010 (N_3010,N_2514,N_2870);
nor U3011 (N_3011,N_2615,N_2602);
or U3012 (N_3012,N_2803,N_2819);
nand U3013 (N_3013,N_2500,N_2896);
and U3014 (N_3014,N_2655,N_2572);
or U3015 (N_3015,N_2716,N_2671);
and U3016 (N_3016,N_2951,N_2528);
and U3017 (N_3017,N_2696,N_2891);
nor U3018 (N_3018,N_2988,N_2542);
nand U3019 (N_3019,N_2592,N_2567);
or U3020 (N_3020,N_2837,N_2631);
and U3021 (N_3021,N_2981,N_2587);
nor U3022 (N_3022,N_2531,N_2685);
or U3023 (N_3023,N_2851,N_2879);
nor U3024 (N_3024,N_2530,N_2698);
and U3025 (N_3025,N_2674,N_2743);
xor U3026 (N_3026,N_2699,N_2720);
and U3027 (N_3027,N_2753,N_2617);
nand U3028 (N_3028,N_2869,N_2882);
and U3029 (N_3029,N_2836,N_2609);
and U3030 (N_3030,N_2562,N_2887);
nand U3031 (N_3031,N_2974,N_2571);
nand U3032 (N_3032,N_2928,N_2605);
nand U3033 (N_3033,N_2812,N_2801);
nand U3034 (N_3034,N_2620,N_2969);
xor U3035 (N_3035,N_2918,N_2727);
or U3036 (N_3036,N_2604,N_2659);
or U3037 (N_3037,N_2731,N_2996);
or U3038 (N_3038,N_2640,N_2850);
or U3039 (N_3039,N_2833,N_2914);
nor U3040 (N_3040,N_2786,N_2730);
nand U3041 (N_3041,N_2556,N_2703);
and U3042 (N_3042,N_2923,N_2825);
nand U3043 (N_3043,N_2907,N_2987);
and U3044 (N_3044,N_2643,N_2994);
and U3045 (N_3045,N_2623,N_2763);
nand U3046 (N_3046,N_2954,N_2815);
nand U3047 (N_3047,N_2748,N_2789);
nand U3048 (N_3048,N_2683,N_2544);
nor U3049 (N_3049,N_2684,N_2548);
nor U3050 (N_3050,N_2780,N_2949);
and U3051 (N_3051,N_2524,N_2877);
or U3052 (N_3052,N_2505,N_2768);
nor U3053 (N_3053,N_2997,N_2711);
and U3054 (N_3054,N_2742,N_2535);
nor U3055 (N_3055,N_2999,N_2751);
or U3056 (N_3056,N_2582,N_2770);
or U3057 (N_3057,N_2734,N_2814);
nand U3058 (N_3058,N_2817,N_2787);
nor U3059 (N_3059,N_2991,N_2594);
or U3060 (N_3060,N_2889,N_2941);
or U3061 (N_3061,N_2845,N_2687);
or U3062 (N_3062,N_2588,N_2894);
or U3063 (N_3063,N_2852,N_2759);
and U3064 (N_3064,N_2989,N_2963);
nor U3065 (N_3065,N_2553,N_2873);
nand U3066 (N_3066,N_2829,N_2664);
nand U3067 (N_3067,N_2913,N_2523);
nand U3068 (N_3068,N_2693,N_2503);
nand U3069 (N_3069,N_2642,N_2966);
nor U3070 (N_3070,N_2905,N_2828);
xor U3071 (N_3071,N_2591,N_2586);
or U3072 (N_3072,N_2899,N_2735);
xnor U3073 (N_3073,N_2970,N_2809);
nand U3074 (N_3074,N_2856,N_2584);
nand U3075 (N_3075,N_2769,N_2897);
or U3076 (N_3076,N_2518,N_2791);
or U3077 (N_3077,N_2895,N_2736);
or U3078 (N_3078,N_2737,N_2679);
nand U3079 (N_3079,N_2827,N_2859);
and U3080 (N_3080,N_2917,N_2876);
nor U3081 (N_3081,N_2761,N_2670);
or U3082 (N_3082,N_2704,N_2630);
xnor U3083 (N_3083,N_2933,N_2926);
nor U3084 (N_3084,N_2794,N_2858);
and U3085 (N_3085,N_2756,N_2849);
or U3086 (N_3086,N_2916,N_2881);
and U3087 (N_3087,N_2757,N_2903);
or U3088 (N_3088,N_2579,N_2626);
nand U3089 (N_3089,N_2909,N_2754);
nor U3090 (N_3090,N_2842,N_2846);
or U3091 (N_3091,N_2884,N_2805);
and U3092 (N_3092,N_2607,N_2614);
and U3093 (N_3093,N_2576,N_2547);
or U3094 (N_3094,N_2629,N_2533);
and U3095 (N_3095,N_2536,N_2892);
and U3096 (N_3096,N_2952,N_2983);
or U3097 (N_3097,N_2841,N_2521);
or U3098 (N_3098,N_2639,N_2599);
and U3099 (N_3099,N_2800,N_2676);
nor U3100 (N_3100,N_2788,N_2611);
or U3101 (N_3101,N_2545,N_2650);
nand U3102 (N_3102,N_2636,N_2985);
and U3103 (N_3103,N_2961,N_2552);
nand U3104 (N_3104,N_2838,N_2930);
and U3105 (N_3105,N_2628,N_2750);
or U3106 (N_3106,N_2672,N_2625);
and U3107 (N_3107,N_2662,N_2589);
or U3108 (N_3108,N_2771,N_2656);
and U3109 (N_3109,N_2948,N_2501);
nor U3110 (N_3110,N_2660,N_2678);
nand U3111 (N_3111,N_2688,N_2510);
nor U3112 (N_3112,N_2747,N_2657);
nand U3113 (N_3113,N_2606,N_2934);
or U3114 (N_3114,N_2818,N_2977);
nor U3115 (N_3115,N_2709,N_2502);
or U3116 (N_3116,N_2875,N_2710);
nand U3117 (N_3117,N_2651,N_2908);
nand U3118 (N_3118,N_2635,N_2546);
nor U3119 (N_3119,N_2816,N_2792);
nand U3120 (N_3120,N_2681,N_2820);
nor U3121 (N_3121,N_2755,N_2959);
or U3122 (N_3122,N_2590,N_2610);
nor U3123 (N_3123,N_2568,N_2774);
nor U3124 (N_3124,N_2924,N_2986);
or U3125 (N_3125,N_2900,N_2645);
and U3126 (N_3126,N_2802,N_2843);
or U3127 (N_3127,N_2772,N_2689);
or U3128 (N_3128,N_2880,N_2575);
and U3129 (N_3129,N_2537,N_2826);
or U3130 (N_3130,N_2778,N_2541);
and U3131 (N_3131,N_2550,N_2511);
nor U3132 (N_3132,N_2947,N_2822);
xnor U3133 (N_3133,N_2627,N_2534);
xor U3134 (N_3134,N_2649,N_2666);
nand U3135 (N_3135,N_2776,N_2539);
and U3136 (N_3136,N_2904,N_2738);
and U3137 (N_3137,N_2733,N_2942);
nand U3138 (N_3138,N_2622,N_2973);
and U3139 (N_3139,N_2878,N_2921);
or U3140 (N_3140,N_2665,N_2613);
nand U3141 (N_3141,N_2922,N_2797);
nand U3142 (N_3142,N_2619,N_2979);
or U3143 (N_3143,N_2779,N_2773);
and U3144 (N_3144,N_2956,N_2863);
and U3145 (N_3145,N_2721,N_2667);
nand U3146 (N_3146,N_2752,N_2936);
and U3147 (N_3147,N_2785,N_2646);
nand U3148 (N_3148,N_2971,N_2580);
nand U3149 (N_3149,N_2808,N_2658);
nand U3150 (N_3150,N_2939,N_2940);
nand U3151 (N_3151,N_2781,N_2965);
or U3152 (N_3152,N_2702,N_2644);
nor U3153 (N_3153,N_2893,N_2975);
nand U3154 (N_3154,N_2740,N_2811);
nand U3155 (N_3155,N_2804,N_2762);
xor U3156 (N_3156,N_2560,N_2680);
or U3157 (N_3157,N_2834,N_2976);
or U3158 (N_3158,N_2868,N_2728);
xnor U3159 (N_3159,N_2967,N_2795);
xor U3160 (N_3160,N_2824,N_2764);
nand U3161 (N_3161,N_2739,N_2980);
or U3162 (N_3162,N_2632,N_2652);
or U3163 (N_3163,N_2741,N_2653);
or U3164 (N_3164,N_2810,N_2516);
nand U3165 (N_3165,N_2766,N_2675);
nor U3166 (N_3166,N_2864,N_2885);
or U3167 (N_3167,N_2998,N_2867);
and U3168 (N_3168,N_2995,N_2932);
nor U3169 (N_3169,N_2578,N_2886);
or U3170 (N_3170,N_2529,N_2638);
nand U3171 (N_3171,N_2661,N_2585);
nand U3172 (N_3172,N_2840,N_2570);
nor U3173 (N_3173,N_2746,N_2962);
nor U3174 (N_3174,N_2832,N_2581);
or U3175 (N_3175,N_2559,N_2565);
and U3176 (N_3176,N_2669,N_2538);
xor U3177 (N_3177,N_2558,N_2937);
or U3178 (N_3178,N_2925,N_2984);
and U3179 (N_3179,N_2700,N_2717);
and U3180 (N_3180,N_2561,N_2600);
nor U3181 (N_3181,N_2958,N_2938);
or U3182 (N_3182,N_2758,N_2931);
nand U3183 (N_3183,N_2847,N_2927);
or U3184 (N_3184,N_2512,N_2633);
or U3185 (N_3185,N_2857,N_2673);
nand U3186 (N_3186,N_2690,N_2705);
nand U3187 (N_3187,N_2601,N_2883);
nor U3188 (N_3188,N_2504,N_2718);
and U3189 (N_3189,N_2950,N_2888);
and U3190 (N_3190,N_2968,N_2813);
nand U3191 (N_3191,N_2807,N_2509);
and U3192 (N_3192,N_2618,N_2982);
nand U3193 (N_3193,N_2782,N_2835);
or U3194 (N_3194,N_2890,N_2677);
and U3195 (N_3195,N_2637,N_2830);
nand U3196 (N_3196,N_2853,N_2682);
or U3197 (N_3197,N_2569,N_2848);
and U3198 (N_3198,N_2831,N_2862);
or U3199 (N_3199,N_2760,N_2719);
or U3200 (N_3200,N_2960,N_2612);
nor U3201 (N_3201,N_2943,N_2668);
or U3202 (N_3202,N_2621,N_2793);
and U3203 (N_3203,N_2634,N_2744);
or U3204 (N_3204,N_2854,N_2745);
nor U3205 (N_3205,N_2597,N_2555);
and U3206 (N_3206,N_2902,N_2920);
xnor U3207 (N_3207,N_2910,N_2855);
or U3208 (N_3208,N_2972,N_2767);
nor U3209 (N_3209,N_2624,N_2978);
or U3210 (N_3210,N_2517,N_2527);
nand U3211 (N_3211,N_2912,N_2563);
and U3212 (N_3212,N_2596,N_2992);
and U3213 (N_3213,N_2515,N_2551);
and U3214 (N_3214,N_2712,N_2566);
nand U3215 (N_3215,N_2608,N_2723);
nand U3216 (N_3216,N_2697,N_2540);
nand U3217 (N_3217,N_2647,N_2957);
nor U3218 (N_3218,N_2844,N_2520);
nor U3219 (N_3219,N_2901,N_2564);
nor U3220 (N_3220,N_2724,N_2603);
nand U3221 (N_3221,N_2513,N_2691);
nand U3222 (N_3222,N_2775,N_2522);
nand U3223 (N_3223,N_2701,N_2557);
and U3224 (N_3224,N_2598,N_2549);
nand U3225 (N_3225,N_2543,N_2706);
or U3226 (N_3226,N_2861,N_2695);
nor U3227 (N_3227,N_2874,N_2554);
nor U3228 (N_3228,N_2593,N_2945);
or U3229 (N_3229,N_2526,N_2860);
and U3230 (N_3230,N_2806,N_2990);
and U3231 (N_3231,N_2993,N_2823);
nor U3232 (N_3232,N_2946,N_2935);
nor U3233 (N_3233,N_2955,N_2784);
and U3234 (N_3234,N_2714,N_2871);
and U3235 (N_3235,N_2532,N_2944);
or U3236 (N_3236,N_2506,N_2790);
and U3237 (N_3237,N_2915,N_2898);
xnor U3238 (N_3238,N_2777,N_2574);
and U3239 (N_3239,N_2732,N_2694);
nand U3240 (N_3240,N_2595,N_2692);
and U3241 (N_3241,N_2911,N_2725);
nor U3242 (N_3242,N_2872,N_2729);
nor U3243 (N_3243,N_2906,N_2654);
and U3244 (N_3244,N_2519,N_2686);
and U3245 (N_3245,N_2799,N_2708);
or U3246 (N_3246,N_2953,N_2707);
and U3247 (N_3247,N_2616,N_2508);
or U3248 (N_3248,N_2919,N_2749);
nand U3249 (N_3249,N_2765,N_2525);
or U3250 (N_3250,N_2699,N_2822);
and U3251 (N_3251,N_2847,N_2924);
nand U3252 (N_3252,N_2875,N_2825);
nand U3253 (N_3253,N_2849,N_2862);
nand U3254 (N_3254,N_2882,N_2872);
and U3255 (N_3255,N_2888,N_2590);
and U3256 (N_3256,N_2875,N_2812);
nor U3257 (N_3257,N_2858,N_2929);
or U3258 (N_3258,N_2704,N_2670);
nand U3259 (N_3259,N_2995,N_2558);
and U3260 (N_3260,N_2683,N_2572);
nor U3261 (N_3261,N_2528,N_2832);
or U3262 (N_3262,N_2624,N_2506);
or U3263 (N_3263,N_2640,N_2786);
nand U3264 (N_3264,N_2912,N_2652);
and U3265 (N_3265,N_2728,N_2601);
nand U3266 (N_3266,N_2514,N_2824);
nor U3267 (N_3267,N_2689,N_2709);
and U3268 (N_3268,N_2840,N_2692);
or U3269 (N_3269,N_2897,N_2763);
or U3270 (N_3270,N_2623,N_2881);
and U3271 (N_3271,N_2835,N_2608);
or U3272 (N_3272,N_2574,N_2767);
nor U3273 (N_3273,N_2939,N_2542);
or U3274 (N_3274,N_2876,N_2774);
nand U3275 (N_3275,N_2811,N_2712);
and U3276 (N_3276,N_2577,N_2597);
or U3277 (N_3277,N_2872,N_2784);
nor U3278 (N_3278,N_2810,N_2957);
nand U3279 (N_3279,N_2558,N_2869);
nand U3280 (N_3280,N_2775,N_2670);
nor U3281 (N_3281,N_2673,N_2888);
xor U3282 (N_3282,N_2661,N_2935);
nand U3283 (N_3283,N_2740,N_2662);
and U3284 (N_3284,N_2653,N_2738);
xor U3285 (N_3285,N_2725,N_2718);
nand U3286 (N_3286,N_2605,N_2793);
or U3287 (N_3287,N_2802,N_2817);
nor U3288 (N_3288,N_2971,N_2965);
nand U3289 (N_3289,N_2821,N_2634);
nand U3290 (N_3290,N_2534,N_2743);
nor U3291 (N_3291,N_2875,N_2707);
nor U3292 (N_3292,N_2848,N_2984);
and U3293 (N_3293,N_2863,N_2618);
nor U3294 (N_3294,N_2867,N_2534);
nor U3295 (N_3295,N_2631,N_2919);
nand U3296 (N_3296,N_2519,N_2678);
or U3297 (N_3297,N_2877,N_2737);
nor U3298 (N_3298,N_2539,N_2951);
xnor U3299 (N_3299,N_2741,N_2501);
nand U3300 (N_3300,N_2905,N_2577);
or U3301 (N_3301,N_2737,N_2907);
nand U3302 (N_3302,N_2942,N_2770);
nor U3303 (N_3303,N_2546,N_2918);
or U3304 (N_3304,N_2604,N_2940);
nor U3305 (N_3305,N_2924,N_2543);
nand U3306 (N_3306,N_2824,N_2763);
and U3307 (N_3307,N_2752,N_2529);
nand U3308 (N_3308,N_2817,N_2864);
or U3309 (N_3309,N_2769,N_2751);
and U3310 (N_3310,N_2502,N_2821);
and U3311 (N_3311,N_2759,N_2547);
xnor U3312 (N_3312,N_2847,N_2716);
or U3313 (N_3313,N_2592,N_2586);
nand U3314 (N_3314,N_2511,N_2935);
or U3315 (N_3315,N_2970,N_2742);
and U3316 (N_3316,N_2852,N_2902);
nor U3317 (N_3317,N_2873,N_2507);
or U3318 (N_3318,N_2688,N_2648);
or U3319 (N_3319,N_2632,N_2949);
nor U3320 (N_3320,N_2949,N_2636);
and U3321 (N_3321,N_2886,N_2820);
or U3322 (N_3322,N_2977,N_2909);
and U3323 (N_3323,N_2775,N_2674);
nor U3324 (N_3324,N_2577,N_2518);
nor U3325 (N_3325,N_2777,N_2750);
or U3326 (N_3326,N_2773,N_2898);
nand U3327 (N_3327,N_2963,N_2750);
or U3328 (N_3328,N_2675,N_2650);
and U3329 (N_3329,N_2730,N_2598);
nand U3330 (N_3330,N_2670,N_2871);
or U3331 (N_3331,N_2747,N_2835);
nand U3332 (N_3332,N_2871,N_2574);
xor U3333 (N_3333,N_2834,N_2829);
nand U3334 (N_3334,N_2547,N_2767);
nor U3335 (N_3335,N_2886,N_2976);
and U3336 (N_3336,N_2955,N_2846);
nand U3337 (N_3337,N_2581,N_2970);
or U3338 (N_3338,N_2564,N_2736);
nor U3339 (N_3339,N_2782,N_2516);
or U3340 (N_3340,N_2668,N_2559);
nor U3341 (N_3341,N_2501,N_2926);
and U3342 (N_3342,N_2761,N_2603);
or U3343 (N_3343,N_2690,N_2831);
and U3344 (N_3344,N_2619,N_2734);
xnor U3345 (N_3345,N_2600,N_2522);
nand U3346 (N_3346,N_2640,N_2659);
or U3347 (N_3347,N_2887,N_2766);
nor U3348 (N_3348,N_2999,N_2724);
or U3349 (N_3349,N_2520,N_2503);
or U3350 (N_3350,N_2734,N_2989);
nand U3351 (N_3351,N_2763,N_2559);
nor U3352 (N_3352,N_2656,N_2902);
or U3353 (N_3353,N_2840,N_2725);
or U3354 (N_3354,N_2509,N_2601);
nor U3355 (N_3355,N_2897,N_2834);
nand U3356 (N_3356,N_2826,N_2667);
and U3357 (N_3357,N_2968,N_2911);
and U3358 (N_3358,N_2671,N_2902);
nand U3359 (N_3359,N_2804,N_2674);
or U3360 (N_3360,N_2770,N_2835);
and U3361 (N_3361,N_2719,N_2804);
xnor U3362 (N_3362,N_2669,N_2981);
xnor U3363 (N_3363,N_2923,N_2898);
and U3364 (N_3364,N_2585,N_2670);
xor U3365 (N_3365,N_2526,N_2540);
and U3366 (N_3366,N_2742,N_2653);
or U3367 (N_3367,N_2869,N_2671);
nand U3368 (N_3368,N_2758,N_2686);
nand U3369 (N_3369,N_2725,N_2919);
or U3370 (N_3370,N_2761,N_2609);
and U3371 (N_3371,N_2590,N_2641);
or U3372 (N_3372,N_2653,N_2615);
or U3373 (N_3373,N_2735,N_2736);
nor U3374 (N_3374,N_2820,N_2682);
and U3375 (N_3375,N_2724,N_2594);
nand U3376 (N_3376,N_2608,N_2798);
nand U3377 (N_3377,N_2589,N_2704);
or U3378 (N_3378,N_2980,N_2546);
and U3379 (N_3379,N_2964,N_2543);
nor U3380 (N_3380,N_2823,N_2864);
xnor U3381 (N_3381,N_2828,N_2537);
xor U3382 (N_3382,N_2814,N_2907);
nor U3383 (N_3383,N_2530,N_2948);
nor U3384 (N_3384,N_2964,N_2509);
and U3385 (N_3385,N_2546,N_2870);
xnor U3386 (N_3386,N_2763,N_2527);
nor U3387 (N_3387,N_2798,N_2737);
nor U3388 (N_3388,N_2776,N_2793);
or U3389 (N_3389,N_2860,N_2841);
nor U3390 (N_3390,N_2855,N_2615);
or U3391 (N_3391,N_2865,N_2753);
xor U3392 (N_3392,N_2725,N_2778);
or U3393 (N_3393,N_2899,N_2908);
nor U3394 (N_3394,N_2598,N_2724);
and U3395 (N_3395,N_2721,N_2861);
nor U3396 (N_3396,N_2831,N_2769);
nor U3397 (N_3397,N_2630,N_2750);
xnor U3398 (N_3398,N_2583,N_2942);
nor U3399 (N_3399,N_2535,N_2959);
nand U3400 (N_3400,N_2874,N_2749);
xnor U3401 (N_3401,N_2939,N_2851);
nand U3402 (N_3402,N_2667,N_2503);
and U3403 (N_3403,N_2786,N_2946);
and U3404 (N_3404,N_2761,N_2517);
nand U3405 (N_3405,N_2786,N_2824);
and U3406 (N_3406,N_2625,N_2586);
nand U3407 (N_3407,N_2926,N_2582);
nand U3408 (N_3408,N_2665,N_2707);
xnor U3409 (N_3409,N_2784,N_2971);
nor U3410 (N_3410,N_2889,N_2879);
or U3411 (N_3411,N_2767,N_2865);
xor U3412 (N_3412,N_2993,N_2576);
and U3413 (N_3413,N_2717,N_2941);
nand U3414 (N_3414,N_2953,N_2759);
nand U3415 (N_3415,N_2831,N_2650);
nand U3416 (N_3416,N_2719,N_2577);
nor U3417 (N_3417,N_2694,N_2561);
or U3418 (N_3418,N_2935,N_2526);
or U3419 (N_3419,N_2908,N_2671);
xor U3420 (N_3420,N_2533,N_2641);
nand U3421 (N_3421,N_2533,N_2999);
and U3422 (N_3422,N_2917,N_2921);
nand U3423 (N_3423,N_2836,N_2908);
xor U3424 (N_3424,N_2907,N_2671);
and U3425 (N_3425,N_2725,N_2623);
nand U3426 (N_3426,N_2595,N_2957);
xor U3427 (N_3427,N_2511,N_2535);
or U3428 (N_3428,N_2517,N_2718);
nor U3429 (N_3429,N_2707,N_2959);
or U3430 (N_3430,N_2859,N_2541);
nor U3431 (N_3431,N_2925,N_2959);
xor U3432 (N_3432,N_2927,N_2755);
nor U3433 (N_3433,N_2926,N_2930);
xnor U3434 (N_3434,N_2547,N_2639);
or U3435 (N_3435,N_2649,N_2858);
nand U3436 (N_3436,N_2583,N_2713);
nor U3437 (N_3437,N_2508,N_2691);
or U3438 (N_3438,N_2804,N_2553);
or U3439 (N_3439,N_2738,N_2550);
nand U3440 (N_3440,N_2509,N_2542);
nand U3441 (N_3441,N_2753,N_2516);
xor U3442 (N_3442,N_2769,N_2772);
and U3443 (N_3443,N_2700,N_2973);
nor U3444 (N_3444,N_2858,N_2671);
nor U3445 (N_3445,N_2555,N_2854);
nor U3446 (N_3446,N_2989,N_2702);
or U3447 (N_3447,N_2970,N_2788);
nor U3448 (N_3448,N_2675,N_2501);
and U3449 (N_3449,N_2545,N_2558);
nand U3450 (N_3450,N_2951,N_2938);
nor U3451 (N_3451,N_2546,N_2822);
or U3452 (N_3452,N_2864,N_2688);
xor U3453 (N_3453,N_2668,N_2552);
and U3454 (N_3454,N_2897,N_2969);
nor U3455 (N_3455,N_2882,N_2555);
nand U3456 (N_3456,N_2983,N_2837);
and U3457 (N_3457,N_2917,N_2783);
and U3458 (N_3458,N_2697,N_2768);
or U3459 (N_3459,N_2745,N_2563);
and U3460 (N_3460,N_2762,N_2617);
or U3461 (N_3461,N_2883,N_2508);
nor U3462 (N_3462,N_2982,N_2948);
nor U3463 (N_3463,N_2910,N_2645);
nor U3464 (N_3464,N_2501,N_2891);
and U3465 (N_3465,N_2906,N_2624);
or U3466 (N_3466,N_2543,N_2507);
and U3467 (N_3467,N_2788,N_2763);
nand U3468 (N_3468,N_2694,N_2795);
xor U3469 (N_3469,N_2767,N_2872);
and U3470 (N_3470,N_2536,N_2692);
nor U3471 (N_3471,N_2937,N_2609);
nor U3472 (N_3472,N_2780,N_2565);
nor U3473 (N_3473,N_2567,N_2940);
and U3474 (N_3474,N_2957,N_2827);
nand U3475 (N_3475,N_2911,N_2654);
nor U3476 (N_3476,N_2731,N_2947);
or U3477 (N_3477,N_2863,N_2519);
and U3478 (N_3478,N_2903,N_2740);
or U3479 (N_3479,N_2506,N_2886);
nand U3480 (N_3480,N_2717,N_2702);
and U3481 (N_3481,N_2827,N_2946);
nand U3482 (N_3482,N_2837,N_2841);
and U3483 (N_3483,N_2849,N_2876);
or U3484 (N_3484,N_2616,N_2612);
or U3485 (N_3485,N_2525,N_2828);
nor U3486 (N_3486,N_2577,N_2639);
or U3487 (N_3487,N_2907,N_2693);
xor U3488 (N_3488,N_2651,N_2748);
xor U3489 (N_3489,N_2843,N_2710);
nor U3490 (N_3490,N_2663,N_2872);
or U3491 (N_3491,N_2983,N_2652);
and U3492 (N_3492,N_2738,N_2932);
nor U3493 (N_3493,N_2645,N_2795);
nand U3494 (N_3494,N_2777,N_2552);
nand U3495 (N_3495,N_2896,N_2900);
nand U3496 (N_3496,N_2670,N_2662);
xor U3497 (N_3497,N_2814,N_2698);
nand U3498 (N_3498,N_2551,N_2900);
nand U3499 (N_3499,N_2914,N_2644);
nand U3500 (N_3500,N_3214,N_3343);
nand U3501 (N_3501,N_3332,N_3348);
and U3502 (N_3502,N_3330,N_3316);
nand U3503 (N_3503,N_3159,N_3108);
and U3504 (N_3504,N_3369,N_3012);
nand U3505 (N_3505,N_3141,N_3157);
or U3506 (N_3506,N_3121,N_3293);
nor U3507 (N_3507,N_3258,N_3496);
nand U3508 (N_3508,N_3417,N_3045);
nor U3509 (N_3509,N_3379,N_3150);
and U3510 (N_3510,N_3487,N_3201);
or U3511 (N_3511,N_3041,N_3459);
nand U3512 (N_3512,N_3129,N_3204);
and U3513 (N_3513,N_3385,N_3125);
nand U3514 (N_3514,N_3378,N_3110);
nand U3515 (N_3515,N_3438,N_3262);
xor U3516 (N_3516,N_3003,N_3230);
xor U3517 (N_3517,N_3461,N_3206);
xnor U3518 (N_3518,N_3170,N_3375);
nand U3519 (N_3519,N_3382,N_3097);
or U3520 (N_3520,N_3051,N_3054);
and U3521 (N_3521,N_3337,N_3364);
or U3522 (N_3522,N_3321,N_3105);
and U3523 (N_3523,N_3238,N_3072);
or U3524 (N_3524,N_3306,N_3409);
nand U3525 (N_3525,N_3484,N_3410);
nand U3526 (N_3526,N_3368,N_3352);
and U3527 (N_3527,N_3236,N_3474);
nor U3528 (N_3528,N_3336,N_3327);
or U3529 (N_3529,N_3387,N_3212);
and U3530 (N_3530,N_3078,N_3413);
nand U3531 (N_3531,N_3328,N_3285);
and U3532 (N_3532,N_3426,N_3087);
nand U3533 (N_3533,N_3454,N_3220);
nor U3534 (N_3534,N_3329,N_3042);
nand U3535 (N_3535,N_3489,N_3216);
and U3536 (N_3536,N_3197,N_3304);
nand U3537 (N_3537,N_3470,N_3008);
or U3538 (N_3538,N_3153,N_3215);
nor U3539 (N_3539,N_3296,N_3113);
or U3540 (N_3540,N_3367,N_3061);
or U3541 (N_3541,N_3482,N_3309);
nand U3542 (N_3542,N_3044,N_3340);
xnor U3543 (N_3543,N_3022,N_3080);
or U3544 (N_3544,N_3037,N_3005);
nor U3545 (N_3545,N_3249,N_3148);
nand U3546 (N_3546,N_3259,N_3143);
xor U3547 (N_3547,N_3444,N_3450);
or U3548 (N_3548,N_3412,N_3280);
nand U3549 (N_3549,N_3406,N_3347);
and U3550 (N_3550,N_3458,N_3033);
nor U3551 (N_3551,N_3248,N_3138);
nor U3552 (N_3552,N_3451,N_3112);
or U3553 (N_3553,N_3147,N_3358);
xnor U3554 (N_3554,N_3366,N_3445);
nand U3555 (N_3555,N_3016,N_3370);
or U3556 (N_3556,N_3100,N_3004);
or U3557 (N_3557,N_3013,N_3497);
or U3558 (N_3558,N_3203,N_3433);
or U3559 (N_3559,N_3355,N_3495);
nand U3560 (N_3560,N_3486,N_3390);
nand U3561 (N_3561,N_3114,N_3298);
nor U3562 (N_3562,N_3418,N_3341);
and U3563 (N_3563,N_3416,N_3034);
or U3564 (N_3564,N_3172,N_3241);
and U3565 (N_3565,N_3448,N_3499);
or U3566 (N_3566,N_3485,N_3128);
or U3567 (N_3567,N_3430,N_3491);
nor U3568 (N_3568,N_3374,N_3242);
and U3569 (N_3569,N_3402,N_3357);
nand U3570 (N_3570,N_3091,N_3323);
and U3571 (N_3571,N_3096,N_3493);
nor U3572 (N_3572,N_3181,N_3463);
or U3573 (N_3573,N_3429,N_3059);
nor U3574 (N_3574,N_3460,N_3188);
or U3575 (N_3575,N_3277,N_3469);
xor U3576 (N_3576,N_3137,N_3017);
xnor U3577 (N_3577,N_3260,N_3488);
and U3578 (N_3578,N_3334,N_3184);
nor U3579 (N_3579,N_3305,N_3002);
nand U3580 (N_3580,N_3393,N_3152);
and U3581 (N_3581,N_3122,N_3415);
nor U3582 (N_3582,N_3342,N_3434);
and U3583 (N_3583,N_3404,N_3351);
or U3584 (N_3584,N_3477,N_3289);
or U3585 (N_3585,N_3398,N_3244);
nor U3586 (N_3586,N_3307,N_3173);
or U3587 (N_3587,N_3095,N_3092);
and U3588 (N_3588,N_3187,N_3359);
and U3589 (N_3589,N_3397,N_3453);
nand U3590 (N_3590,N_3027,N_3456);
or U3591 (N_3591,N_3345,N_3046);
xnor U3592 (N_3592,N_3401,N_3464);
xnor U3593 (N_3593,N_3218,N_3168);
nor U3594 (N_3594,N_3376,N_3039);
nand U3595 (N_3595,N_3442,N_3164);
and U3596 (N_3596,N_3311,N_3425);
xnor U3597 (N_3597,N_3196,N_3243);
nand U3598 (N_3598,N_3064,N_3475);
xor U3599 (N_3599,N_3000,N_3297);
nor U3600 (N_3600,N_3057,N_3396);
or U3601 (N_3601,N_3209,N_3466);
or U3602 (N_3602,N_3287,N_3176);
or U3603 (N_3603,N_3268,N_3210);
xnor U3604 (N_3604,N_3213,N_3437);
and U3605 (N_3605,N_3014,N_3136);
and U3606 (N_3606,N_3391,N_3235);
or U3607 (N_3607,N_3208,N_3058);
or U3608 (N_3608,N_3109,N_3120);
nand U3609 (N_3609,N_3062,N_3394);
and U3610 (N_3610,N_3300,N_3407);
or U3611 (N_3611,N_3098,N_3179);
or U3612 (N_3612,N_3006,N_3077);
nor U3613 (N_3613,N_3422,N_3362);
nand U3614 (N_3614,N_3028,N_3011);
nand U3615 (N_3615,N_3167,N_3377);
and U3616 (N_3616,N_3269,N_3265);
and U3617 (N_3617,N_3205,N_3030);
nor U3618 (N_3618,N_3498,N_3252);
nor U3619 (N_3619,N_3480,N_3349);
nand U3620 (N_3620,N_3326,N_3270);
or U3621 (N_3621,N_3103,N_3026);
nor U3622 (N_3622,N_3361,N_3117);
or U3623 (N_3623,N_3303,N_3273);
and U3624 (N_3624,N_3492,N_3198);
nand U3625 (N_3625,N_3428,N_3392);
or U3626 (N_3626,N_3145,N_3421);
nand U3627 (N_3627,N_3240,N_3221);
or U3628 (N_3628,N_3119,N_3472);
nor U3629 (N_3629,N_3162,N_3036);
nor U3630 (N_3630,N_3419,N_3211);
nand U3631 (N_3631,N_3452,N_3111);
or U3632 (N_3632,N_3085,N_3118);
nand U3633 (N_3633,N_3079,N_3178);
nor U3634 (N_3634,N_3250,N_3146);
or U3635 (N_3635,N_3133,N_3186);
and U3636 (N_3636,N_3199,N_3139);
and U3637 (N_3637,N_3018,N_3455);
or U3638 (N_3638,N_3424,N_3228);
nand U3639 (N_3639,N_3089,N_3222);
nand U3640 (N_3640,N_3052,N_3255);
and U3641 (N_3641,N_3473,N_3135);
nor U3642 (N_3642,N_3432,N_3015);
or U3643 (N_3643,N_3123,N_3130);
and U3644 (N_3644,N_3194,N_3383);
and U3645 (N_3645,N_3081,N_3142);
nor U3646 (N_3646,N_3325,N_3344);
xor U3647 (N_3647,N_3408,N_3301);
nor U3648 (N_3648,N_3024,N_3155);
and U3649 (N_3649,N_3317,N_3063);
and U3650 (N_3650,N_3131,N_3237);
or U3651 (N_3651,N_3048,N_3449);
and U3652 (N_3652,N_3086,N_3400);
nor U3653 (N_3653,N_3099,N_3266);
and U3654 (N_3654,N_3231,N_3446);
and U3655 (N_3655,N_3001,N_3322);
nor U3656 (N_3656,N_3158,N_3462);
nor U3657 (N_3657,N_3284,N_3403);
nor U3658 (N_3658,N_3386,N_3360);
nand U3659 (N_3659,N_3185,N_3049);
and U3660 (N_3660,N_3363,N_3275);
xor U3661 (N_3661,N_3101,N_3245);
nor U3662 (N_3662,N_3233,N_3234);
and U3663 (N_3663,N_3202,N_3104);
nor U3664 (N_3664,N_3381,N_3224);
xnor U3665 (N_3665,N_3320,N_3254);
or U3666 (N_3666,N_3315,N_3082);
or U3667 (N_3667,N_3182,N_3065);
nand U3668 (N_3668,N_3084,N_3441);
nor U3669 (N_3669,N_3050,N_3102);
or U3670 (N_3670,N_3276,N_3060);
xor U3671 (N_3671,N_3476,N_3395);
and U3672 (N_3672,N_3115,N_3318);
nand U3673 (N_3673,N_3174,N_3411);
and U3674 (N_3674,N_3282,N_3365);
nor U3675 (N_3675,N_3314,N_3180);
nor U3676 (N_3676,N_3025,N_3405);
and U3677 (N_3677,N_3278,N_3479);
and U3678 (N_3678,N_3124,N_3299);
and U3679 (N_3679,N_3468,N_3190);
and U3680 (N_3680,N_3171,N_3294);
nor U3681 (N_3681,N_3288,N_3076);
and U3682 (N_3682,N_3281,N_3169);
nor U3683 (N_3683,N_3312,N_3331);
nor U3684 (N_3684,N_3490,N_3251);
or U3685 (N_3685,N_3217,N_3443);
xor U3686 (N_3686,N_3494,N_3160);
nand U3687 (N_3687,N_3335,N_3447);
nor U3688 (N_3688,N_3261,N_3020);
and U3689 (N_3689,N_3126,N_3195);
nand U3690 (N_3690,N_3156,N_3021);
nand U3691 (N_3691,N_3090,N_3056);
nor U3692 (N_3692,N_3313,N_3047);
or U3693 (N_3693,N_3038,N_3324);
nor U3694 (N_3694,N_3354,N_3283);
or U3695 (N_3695,N_3031,N_3371);
nor U3696 (N_3696,N_3279,N_3423);
nor U3697 (N_3697,N_3035,N_3183);
and U3698 (N_3698,N_3339,N_3132);
and U3699 (N_3699,N_3239,N_3319);
nand U3700 (N_3700,N_3471,N_3023);
nand U3701 (N_3701,N_3154,N_3165);
and U3702 (N_3702,N_3353,N_3140);
nor U3703 (N_3703,N_3291,N_3007);
nor U3704 (N_3704,N_3040,N_3043);
nor U3705 (N_3705,N_3414,N_3420);
and U3706 (N_3706,N_3191,N_3478);
xnor U3707 (N_3707,N_3483,N_3151);
or U3708 (N_3708,N_3106,N_3380);
xnor U3709 (N_3709,N_3274,N_3225);
nor U3710 (N_3710,N_3272,N_3175);
nand U3711 (N_3711,N_3435,N_3247);
nor U3712 (N_3712,N_3338,N_3308);
or U3713 (N_3713,N_3093,N_3457);
nand U3714 (N_3714,N_3246,N_3075);
and U3715 (N_3715,N_3029,N_3333);
nand U3716 (N_3716,N_3127,N_3200);
or U3717 (N_3717,N_3055,N_3149);
xor U3718 (N_3718,N_3372,N_3134);
nor U3719 (N_3719,N_3256,N_3193);
nor U3720 (N_3720,N_3292,N_3439);
and U3721 (N_3721,N_3373,N_3431);
nand U3722 (N_3722,N_3069,N_3088);
and U3723 (N_3723,N_3310,N_3067);
nand U3724 (N_3724,N_3264,N_3302);
nor U3725 (N_3725,N_3440,N_3019);
nand U3726 (N_3726,N_3207,N_3356);
xor U3727 (N_3727,N_3071,N_3189);
nand U3728 (N_3728,N_3177,N_3427);
nor U3729 (N_3729,N_3253,N_3094);
and U3730 (N_3730,N_3436,N_3384);
or U3731 (N_3731,N_3295,N_3163);
and U3732 (N_3732,N_3223,N_3399);
nand U3733 (N_3733,N_3227,N_3232);
or U3734 (N_3734,N_3073,N_3070);
nand U3735 (N_3735,N_3066,N_3116);
and U3736 (N_3736,N_3219,N_3257);
and U3737 (N_3737,N_3263,N_3226);
or U3738 (N_3738,N_3271,N_3009);
or U3739 (N_3739,N_3465,N_3350);
and U3740 (N_3740,N_3229,N_3286);
or U3741 (N_3741,N_3346,N_3053);
nor U3742 (N_3742,N_3144,N_3290);
nand U3743 (N_3743,N_3083,N_3267);
and U3744 (N_3744,N_3161,N_3074);
and U3745 (N_3745,N_3032,N_3166);
nand U3746 (N_3746,N_3068,N_3192);
or U3747 (N_3747,N_3389,N_3107);
or U3748 (N_3748,N_3481,N_3467);
and U3749 (N_3749,N_3388,N_3010);
or U3750 (N_3750,N_3288,N_3416);
nor U3751 (N_3751,N_3044,N_3190);
xor U3752 (N_3752,N_3159,N_3290);
and U3753 (N_3753,N_3389,N_3056);
nand U3754 (N_3754,N_3454,N_3256);
or U3755 (N_3755,N_3010,N_3041);
or U3756 (N_3756,N_3474,N_3291);
nor U3757 (N_3757,N_3095,N_3340);
xnor U3758 (N_3758,N_3015,N_3310);
nand U3759 (N_3759,N_3193,N_3249);
nor U3760 (N_3760,N_3052,N_3294);
xnor U3761 (N_3761,N_3112,N_3120);
nand U3762 (N_3762,N_3475,N_3479);
nor U3763 (N_3763,N_3380,N_3450);
nor U3764 (N_3764,N_3144,N_3331);
nor U3765 (N_3765,N_3106,N_3163);
nor U3766 (N_3766,N_3177,N_3163);
nor U3767 (N_3767,N_3299,N_3306);
nor U3768 (N_3768,N_3406,N_3083);
nor U3769 (N_3769,N_3383,N_3359);
nor U3770 (N_3770,N_3231,N_3383);
nand U3771 (N_3771,N_3155,N_3144);
xnor U3772 (N_3772,N_3292,N_3173);
nand U3773 (N_3773,N_3309,N_3133);
xnor U3774 (N_3774,N_3095,N_3187);
nand U3775 (N_3775,N_3358,N_3022);
and U3776 (N_3776,N_3168,N_3451);
nand U3777 (N_3777,N_3085,N_3445);
nand U3778 (N_3778,N_3402,N_3141);
or U3779 (N_3779,N_3321,N_3248);
or U3780 (N_3780,N_3280,N_3004);
and U3781 (N_3781,N_3376,N_3291);
or U3782 (N_3782,N_3452,N_3109);
or U3783 (N_3783,N_3429,N_3342);
nand U3784 (N_3784,N_3166,N_3309);
or U3785 (N_3785,N_3177,N_3142);
and U3786 (N_3786,N_3268,N_3269);
nor U3787 (N_3787,N_3451,N_3187);
xnor U3788 (N_3788,N_3197,N_3291);
nand U3789 (N_3789,N_3169,N_3371);
or U3790 (N_3790,N_3478,N_3225);
nor U3791 (N_3791,N_3330,N_3417);
or U3792 (N_3792,N_3436,N_3148);
or U3793 (N_3793,N_3442,N_3089);
and U3794 (N_3794,N_3432,N_3199);
nor U3795 (N_3795,N_3070,N_3411);
xor U3796 (N_3796,N_3110,N_3084);
or U3797 (N_3797,N_3430,N_3440);
or U3798 (N_3798,N_3478,N_3216);
xor U3799 (N_3799,N_3471,N_3482);
nor U3800 (N_3800,N_3493,N_3339);
and U3801 (N_3801,N_3151,N_3382);
or U3802 (N_3802,N_3358,N_3332);
and U3803 (N_3803,N_3427,N_3338);
or U3804 (N_3804,N_3417,N_3399);
or U3805 (N_3805,N_3278,N_3287);
xnor U3806 (N_3806,N_3075,N_3308);
and U3807 (N_3807,N_3317,N_3383);
and U3808 (N_3808,N_3069,N_3117);
xor U3809 (N_3809,N_3057,N_3299);
or U3810 (N_3810,N_3431,N_3217);
xor U3811 (N_3811,N_3431,N_3197);
xnor U3812 (N_3812,N_3090,N_3268);
nand U3813 (N_3813,N_3188,N_3179);
nor U3814 (N_3814,N_3298,N_3216);
nor U3815 (N_3815,N_3198,N_3010);
xor U3816 (N_3816,N_3359,N_3107);
or U3817 (N_3817,N_3090,N_3082);
nor U3818 (N_3818,N_3482,N_3057);
nand U3819 (N_3819,N_3353,N_3084);
nand U3820 (N_3820,N_3460,N_3345);
and U3821 (N_3821,N_3393,N_3044);
and U3822 (N_3822,N_3298,N_3103);
nor U3823 (N_3823,N_3148,N_3467);
nor U3824 (N_3824,N_3267,N_3111);
and U3825 (N_3825,N_3144,N_3306);
nand U3826 (N_3826,N_3084,N_3215);
nor U3827 (N_3827,N_3044,N_3397);
nand U3828 (N_3828,N_3061,N_3150);
nand U3829 (N_3829,N_3317,N_3480);
nand U3830 (N_3830,N_3405,N_3304);
or U3831 (N_3831,N_3456,N_3486);
nor U3832 (N_3832,N_3024,N_3174);
or U3833 (N_3833,N_3266,N_3327);
and U3834 (N_3834,N_3411,N_3436);
nor U3835 (N_3835,N_3255,N_3076);
nand U3836 (N_3836,N_3061,N_3305);
nand U3837 (N_3837,N_3402,N_3339);
nor U3838 (N_3838,N_3033,N_3261);
nand U3839 (N_3839,N_3201,N_3422);
and U3840 (N_3840,N_3115,N_3236);
or U3841 (N_3841,N_3173,N_3027);
or U3842 (N_3842,N_3271,N_3466);
and U3843 (N_3843,N_3357,N_3056);
or U3844 (N_3844,N_3055,N_3054);
or U3845 (N_3845,N_3080,N_3415);
xnor U3846 (N_3846,N_3438,N_3255);
nor U3847 (N_3847,N_3393,N_3376);
nand U3848 (N_3848,N_3433,N_3418);
nand U3849 (N_3849,N_3487,N_3446);
nand U3850 (N_3850,N_3305,N_3360);
nand U3851 (N_3851,N_3407,N_3283);
nor U3852 (N_3852,N_3039,N_3101);
nor U3853 (N_3853,N_3011,N_3362);
nand U3854 (N_3854,N_3461,N_3448);
and U3855 (N_3855,N_3114,N_3122);
nor U3856 (N_3856,N_3035,N_3073);
xor U3857 (N_3857,N_3009,N_3352);
and U3858 (N_3858,N_3002,N_3394);
or U3859 (N_3859,N_3090,N_3017);
and U3860 (N_3860,N_3383,N_3457);
nand U3861 (N_3861,N_3152,N_3391);
and U3862 (N_3862,N_3250,N_3269);
nor U3863 (N_3863,N_3441,N_3462);
and U3864 (N_3864,N_3284,N_3282);
xor U3865 (N_3865,N_3329,N_3098);
or U3866 (N_3866,N_3278,N_3184);
nand U3867 (N_3867,N_3368,N_3304);
and U3868 (N_3868,N_3265,N_3248);
and U3869 (N_3869,N_3365,N_3159);
xnor U3870 (N_3870,N_3409,N_3224);
nand U3871 (N_3871,N_3079,N_3455);
and U3872 (N_3872,N_3298,N_3386);
nor U3873 (N_3873,N_3422,N_3199);
and U3874 (N_3874,N_3273,N_3422);
xor U3875 (N_3875,N_3484,N_3241);
nor U3876 (N_3876,N_3468,N_3399);
xor U3877 (N_3877,N_3406,N_3492);
xor U3878 (N_3878,N_3269,N_3306);
and U3879 (N_3879,N_3133,N_3242);
nand U3880 (N_3880,N_3068,N_3267);
and U3881 (N_3881,N_3246,N_3381);
nor U3882 (N_3882,N_3193,N_3094);
and U3883 (N_3883,N_3272,N_3156);
nor U3884 (N_3884,N_3342,N_3358);
or U3885 (N_3885,N_3078,N_3341);
nor U3886 (N_3886,N_3274,N_3207);
nand U3887 (N_3887,N_3010,N_3104);
and U3888 (N_3888,N_3102,N_3441);
nand U3889 (N_3889,N_3382,N_3336);
nand U3890 (N_3890,N_3319,N_3005);
nand U3891 (N_3891,N_3352,N_3345);
nand U3892 (N_3892,N_3365,N_3325);
nand U3893 (N_3893,N_3030,N_3044);
or U3894 (N_3894,N_3484,N_3418);
nand U3895 (N_3895,N_3174,N_3097);
or U3896 (N_3896,N_3402,N_3137);
nor U3897 (N_3897,N_3435,N_3075);
nor U3898 (N_3898,N_3171,N_3493);
nor U3899 (N_3899,N_3328,N_3277);
and U3900 (N_3900,N_3174,N_3241);
and U3901 (N_3901,N_3445,N_3007);
and U3902 (N_3902,N_3363,N_3058);
nor U3903 (N_3903,N_3011,N_3261);
or U3904 (N_3904,N_3035,N_3207);
nand U3905 (N_3905,N_3044,N_3213);
xor U3906 (N_3906,N_3383,N_3240);
nor U3907 (N_3907,N_3223,N_3263);
or U3908 (N_3908,N_3244,N_3425);
and U3909 (N_3909,N_3165,N_3230);
and U3910 (N_3910,N_3326,N_3092);
xor U3911 (N_3911,N_3262,N_3171);
and U3912 (N_3912,N_3152,N_3048);
nor U3913 (N_3913,N_3217,N_3036);
or U3914 (N_3914,N_3380,N_3345);
xnor U3915 (N_3915,N_3241,N_3240);
and U3916 (N_3916,N_3125,N_3448);
nor U3917 (N_3917,N_3055,N_3369);
and U3918 (N_3918,N_3105,N_3147);
nor U3919 (N_3919,N_3152,N_3276);
or U3920 (N_3920,N_3106,N_3298);
nand U3921 (N_3921,N_3154,N_3047);
nand U3922 (N_3922,N_3326,N_3491);
and U3923 (N_3923,N_3064,N_3403);
or U3924 (N_3924,N_3495,N_3304);
nand U3925 (N_3925,N_3178,N_3376);
nor U3926 (N_3926,N_3394,N_3351);
nor U3927 (N_3927,N_3060,N_3427);
or U3928 (N_3928,N_3419,N_3295);
or U3929 (N_3929,N_3198,N_3169);
nand U3930 (N_3930,N_3001,N_3321);
nand U3931 (N_3931,N_3013,N_3392);
xor U3932 (N_3932,N_3396,N_3032);
nand U3933 (N_3933,N_3499,N_3332);
or U3934 (N_3934,N_3117,N_3405);
and U3935 (N_3935,N_3083,N_3031);
nand U3936 (N_3936,N_3079,N_3291);
nor U3937 (N_3937,N_3176,N_3332);
nor U3938 (N_3938,N_3107,N_3407);
nand U3939 (N_3939,N_3262,N_3439);
or U3940 (N_3940,N_3318,N_3494);
and U3941 (N_3941,N_3304,N_3274);
xnor U3942 (N_3942,N_3145,N_3091);
xnor U3943 (N_3943,N_3449,N_3485);
nor U3944 (N_3944,N_3130,N_3252);
and U3945 (N_3945,N_3006,N_3064);
or U3946 (N_3946,N_3092,N_3191);
nor U3947 (N_3947,N_3186,N_3084);
or U3948 (N_3948,N_3052,N_3102);
and U3949 (N_3949,N_3207,N_3403);
nand U3950 (N_3950,N_3398,N_3171);
or U3951 (N_3951,N_3052,N_3142);
nand U3952 (N_3952,N_3433,N_3037);
or U3953 (N_3953,N_3213,N_3348);
and U3954 (N_3954,N_3188,N_3274);
and U3955 (N_3955,N_3364,N_3186);
and U3956 (N_3956,N_3268,N_3115);
nor U3957 (N_3957,N_3047,N_3437);
nor U3958 (N_3958,N_3099,N_3446);
or U3959 (N_3959,N_3053,N_3287);
and U3960 (N_3960,N_3111,N_3058);
or U3961 (N_3961,N_3382,N_3387);
nand U3962 (N_3962,N_3122,N_3057);
nor U3963 (N_3963,N_3216,N_3480);
or U3964 (N_3964,N_3205,N_3122);
and U3965 (N_3965,N_3027,N_3269);
nor U3966 (N_3966,N_3196,N_3379);
nor U3967 (N_3967,N_3028,N_3022);
xnor U3968 (N_3968,N_3138,N_3125);
and U3969 (N_3969,N_3028,N_3440);
and U3970 (N_3970,N_3110,N_3424);
and U3971 (N_3971,N_3215,N_3274);
and U3972 (N_3972,N_3016,N_3380);
and U3973 (N_3973,N_3099,N_3173);
and U3974 (N_3974,N_3441,N_3455);
or U3975 (N_3975,N_3123,N_3165);
nand U3976 (N_3976,N_3264,N_3034);
nand U3977 (N_3977,N_3210,N_3306);
and U3978 (N_3978,N_3391,N_3182);
nand U3979 (N_3979,N_3478,N_3004);
xnor U3980 (N_3980,N_3096,N_3118);
nor U3981 (N_3981,N_3383,N_3247);
and U3982 (N_3982,N_3390,N_3421);
or U3983 (N_3983,N_3264,N_3112);
or U3984 (N_3984,N_3173,N_3282);
or U3985 (N_3985,N_3347,N_3159);
nand U3986 (N_3986,N_3018,N_3149);
nor U3987 (N_3987,N_3069,N_3178);
nand U3988 (N_3988,N_3250,N_3316);
xor U3989 (N_3989,N_3068,N_3275);
nand U3990 (N_3990,N_3484,N_3142);
and U3991 (N_3991,N_3171,N_3178);
nand U3992 (N_3992,N_3244,N_3023);
and U3993 (N_3993,N_3452,N_3143);
and U3994 (N_3994,N_3284,N_3325);
or U3995 (N_3995,N_3362,N_3333);
and U3996 (N_3996,N_3194,N_3158);
nor U3997 (N_3997,N_3239,N_3290);
nand U3998 (N_3998,N_3142,N_3210);
and U3999 (N_3999,N_3119,N_3231);
or U4000 (N_4000,N_3624,N_3570);
and U4001 (N_4001,N_3525,N_3899);
nor U4002 (N_4002,N_3533,N_3988);
nand U4003 (N_4003,N_3890,N_3660);
and U4004 (N_4004,N_3627,N_3607);
nor U4005 (N_4005,N_3686,N_3736);
nand U4006 (N_4006,N_3503,N_3568);
and U4007 (N_4007,N_3937,N_3906);
and U4008 (N_4008,N_3892,N_3507);
or U4009 (N_4009,N_3779,N_3797);
or U4010 (N_4010,N_3821,N_3612);
xnor U4011 (N_4011,N_3844,N_3975);
xnor U4012 (N_4012,N_3957,N_3809);
or U4013 (N_4013,N_3518,N_3691);
xnor U4014 (N_4014,N_3863,N_3746);
nor U4015 (N_4015,N_3757,N_3886);
nand U4016 (N_4016,N_3870,N_3959);
nand U4017 (N_4017,N_3909,N_3788);
nor U4018 (N_4018,N_3625,N_3618);
nand U4019 (N_4019,N_3898,N_3970);
nor U4020 (N_4020,N_3963,N_3512);
nand U4021 (N_4021,N_3641,N_3868);
nand U4022 (N_4022,N_3972,N_3773);
nor U4023 (N_4023,N_3843,N_3633);
nor U4024 (N_4024,N_3884,N_3928);
and U4025 (N_4025,N_3556,N_3905);
nand U4026 (N_4026,N_3666,N_3669);
nor U4027 (N_4027,N_3560,N_3699);
nor U4028 (N_4028,N_3923,N_3778);
and U4029 (N_4029,N_3679,N_3751);
nand U4030 (N_4030,N_3687,N_3745);
or U4031 (N_4031,N_3648,N_3847);
nor U4032 (N_4032,N_3728,N_3643);
or U4033 (N_4033,N_3676,N_3850);
nor U4034 (N_4034,N_3596,N_3969);
or U4035 (N_4035,N_3961,N_3735);
and U4036 (N_4036,N_3922,N_3772);
or U4037 (N_4037,N_3833,N_3828);
nor U4038 (N_4038,N_3943,N_3690);
or U4039 (N_4039,N_3576,N_3851);
nand U4040 (N_4040,N_3700,N_3767);
and U4041 (N_4041,N_3783,N_3601);
nand U4042 (N_4042,N_3599,N_3562);
or U4043 (N_4043,N_3724,N_3849);
xnor U4044 (N_4044,N_3893,N_3853);
or U4045 (N_4045,N_3741,N_3832);
nand U4046 (N_4046,N_3729,N_3526);
or U4047 (N_4047,N_3836,N_3765);
xnor U4048 (N_4048,N_3984,N_3760);
nand U4049 (N_4049,N_3829,N_3671);
and U4050 (N_4050,N_3575,N_3897);
nand U4051 (N_4051,N_3855,N_3696);
and U4052 (N_4052,N_3665,N_3531);
nor U4053 (N_4053,N_3674,N_3727);
or U4054 (N_4054,N_3550,N_3662);
and U4055 (N_4055,N_3678,N_3638);
and U4056 (N_4056,N_3642,N_3555);
nand U4057 (N_4057,N_3530,N_3619);
nand U4058 (N_4058,N_3508,N_3711);
nand U4059 (N_4059,N_3811,N_3582);
or U4060 (N_4060,N_3659,N_3501);
xor U4061 (N_4061,N_3588,N_3874);
and U4062 (N_4062,N_3820,N_3706);
and U4063 (N_4063,N_3640,N_3904);
xor U4064 (N_4064,N_3717,N_3791);
or U4065 (N_4065,N_3517,N_3723);
and U4066 (N_4066,N_3744,N_3994);
nor U4067 (N_4067,N_3789,N_3846);
or U4068 (N_4068,N_3578,N_3573);
nand U4069 (N_4069,N_3860,N_3990);
or U4070 (N_4070,N_3812,N_3502);
nor U4071 (N_4071,N_3817,N_3930);
nor U4072 (N_4072,N_3871,N_3520);
nor U4073 (N_4073,N_3748,N_3726);
xnor U4074 (N_4074,N_3579,N_3598);
or U4075 (N_4075,N_3739,N_3646);
nor U4076 (N_4076,N_3987,N_3938);
and U4077 (N_4077,N_3949,N_3749);
xnor U4078 (N_4078,N_3613,N_3887);
nand U4079 (N_4079,N_3796,N_3973);
and U4080 (N_4080,N_3587,N_3819);
or U4081 (N_4081,N_3976,N_3514);
nand U4082 (N_4082,N_3952,N_3784);
nor U4083 (N_4083,N_3620,N_3668);
nand U4084 (N_4084,N_3623,N_3856);
and U4085 (N_4085,N_3622,N_3553);
and U4086 (N_4086,N_3753,N_3876);
xor U4087 (N_4087,N_3771,N_3998);
nor U4088 (N_4088,N_3509,N_3907);
and U4089 (N_4089,N_3945,N_3740);
nand U4090 (N_4090,N_3629,N_3572);
and U4091 (N_4091,N_3549,N_3658);
nand U4092 (N_4092,N_3755,N_3875);
or U4093 (N_4093,N_3859,N_3799);
nand U4094 (N_4094,N_3636,N_3754);
nand U4095 (N_4095,N_3865,N_3780);
nand U4096 (N_4096,N_3628,N_3775);
nor U4097 (N_4097,N_3927,N_3781);
or U4098 (N_4098,N_3806,N_3593);
xor U4099 (N_4099,N_3602,N_3584);
nor U4100 (N_4100,N_3803,N_3719);
or U4101 (N_4101,N_3944,N_3889);
xor U4102 (N_4102,N_3566,N_3936);
and U4103 (N_4103,N_3867,N_3776);
or U4104 (N_4104,N_3524,N_3521);
or U4105 (N_4105,N_3814,N_3664);
and U4106 (N_4106,N_3785,N_3793);
and U4107 (N_4107,N_3795,N_3583);
or U4108 (N_4108,N_3698,N_3813);
and U4109 (N_4109,N_3818,N_3840);
nand U4110 (N_4110,N_3802,N_3552);
nand U4111 (N_4111,N_3845,N_3725);
nor U4112 (N_4112,N_3635,N_3880);
nand U4113 (N_4113,N_3675,N_3766);
nor U4114 (N_4114,N_3911,N_3816);
nand U4115 (N_4115,N_3839,N_3983);
or U4116 (N_4116,N_3738,N_3694);
and U4117 (N_4117,N_3605,N_3902);
nand U4118 (N_4118,N_3653,N_3878);
nor U4119 (N_4119,N_3992,N_3667);
nor U4120 (N_4120,N_3704,N_3900);
nand U4121 (N_4121,N_3823,N_3842);
nor U4122 (N_4122,N_3956,N_3857);
xnor U4123 (N_4123,N_3825,N_3805);
nand U4124 (N_4124,N_3958,N_3702);
nand U4125 (N_4125,N_3873,N_3854);
xnor U4126 (N_4126,N_3954,N_3921);
nand U4127 (N_4127,N_3684,N_3715);
nor U4128 (N_4128,N_3996,N_3991);
nor U4129 (N_4129,N_3981,N_3948);
nor U4130 (N_4130,N_3663,N_3971);
or U4131 (N_4131,N_3610,N_3689);
nand U4132 (N_4132,N_3955,N_3722);
and U4133 (N_4133,N_3528,N_3670);
or U4134 (N_4134,N_3858,N_3534);
and U4135 (N_4135,N_3609,N_3537);
nand U4136 (N_4136,N_3883,N_3801);
or U4137 (N_4137,N_3787,N_3705);
nor U4138 (N_4138,N_3798,N_3869);
nand U4139 (N_4139,N_3585,N_3968);
or U4140 (N_4140,N_3631,N_3777);
nor U4141 (N_4141,N_3986,N_3942);
nor U4142 (N_4142,N_3527,N_3752);
and U4143 (N_4143,N_3693,N_3580);
nor U4144 (N_4144,N_3737,N_3567);
nand U4145 (N_4145,N_3808,N_3830);
nand U4146 (N_4146,N_3810,N_3731);
and U4147 (N_4147,N_3993,N_3965);
xor U4148 (N_4148,N_3546,N_3848);
and U4149 (N_4149,N_3564,N_3914);
xor U4150 (N_4150,N_3966,N_3926);
and U4151 (N_4151,N_3827,N_3908);
nor U4152 (N_4152,N_3529,N_3559);
nand U4153 (N_4153,N_3852,N_3831);
and U4154 (N_4154,N_3547,N_3695);
or U4155 (N_4155,N_3913,N_3759);
nor U4156 (N_4156,N_3951,N_3683);
nor U4157 (N_4157,N_3750,N_3545);
nand U4158 (N_4158,N_3510,N_3995);
nor U4159 (N_4159,N_3758,N_3756);
xnor U4160 (N_4160,N_3652,N_3708);
or U4161 (N_4161,N_3569,N_3637);
xor U4162 (N_4162,N_3542,N_3935);
nand U4163 (N_4163,N_3548,N_3634);
nand U4164 (N_4164,N_3800,N_3532);
or U4165 (N_4165,N_3692,N_3896);
and U4166 (N_4166,N_3505,N_3838);
and U4167 (N_4167,N_3673,N_3516);
or U4168 (N_4168,N_3713,N_3656);
nor U4169 (N_4169,N_3980,N_3931);
or U4170 (N_4170,N_3974,N_3761);
nand U4171 (N_4171,N_3558,N_3815);
or U4172 (N_4172,N_3770,N_3682);
nor U4173 (N_4173,N_3581,N_3577);
or U4174 (N_4174,N_3939,N_3912);
xnor U4175 (N_4175,N_3500,N_3934);
and U4176 (N_4176,N_3763,N_3639);
xnor U4177 (N_4177,N_3826,N_3977);
nor U4178 (N_4178,N_3764,N_3742);
nand U4179 (N_4179,N_3539,N_3960);
and U4180 (N_4180,N_3657,N_3962);
or U4181 (N_4181,N_3837,N_3595);
nor U4182 (N_4182,N_3626,N_3732);
xnor U4183 (N_4183,N_3862,N_3710);
and U4184 (N_4184,N_3733,N_3879);
and U4185 (N_4185,N_3621,N_3964);
xnor U4186 (N_4186,N_3557,N_3989);
nand U4187 (N_4187,N_3978,N_3649);
and U4188 (N_4188,N_3940,N_3523);
nor U4189 (N_4189,N_3536,N_3586);
or U4190 (N_4190,N_3834,N_3701);
nand U4191 (N_4191,N_3611,N_3712);
or U4192 (N_4192,N_3565,N_3967);
and U4193 (N_4193,N_3918,N_3769);
nor U4194 (N_4194,N_3804,N_3903);
nor U4195 (N_4195,N_3707,N_3681);
or U4196 (N_4196,N_3504,N_3571);
nor U4197 (N_4197,N_3774,N_3592);
nand U4198 (N_4198,N_3654,N_3932);
and U4199 (N_4199,N_3762,N_3985);
or U4200 (N_4200,N_3824,N_3718);
and U4201 (N_4201,N_3513,N_3866);
or U4202 (N_4202,N_3574,N_3685);
nor U4203 (N_4203,N_3794,N_3925);
or U4204 (N_4204,N_3786,N_3895);
or U4205 (N_4205,N_3538,N_3947);
and U4206 (N_4206,N_3616,N_3677);
or U4207 (N_4207,N_3716,N_3551);
nor U4208 (N_4208,N_3888,N_3600);
nand U4209 (N_4209,N_3522,N_3563);
or U4210 (N_4210,N_3543,N_3894);
nor U4211 (N_4211,N_3535,N_3661);
nor U4212 (N_4212,N_3915,N_3544);
and U4213 (N_4213,N_3933,N_3877);
and U4214 (N_4214,N_3554,N_3697);
nand U4215 (N_4215,N_3924,N_3941);
nor U4216 (N_4216,N_3519,N_3672);
and U4217 (N_4217,N_3651,N_3594);
and U4218 (N_4218,N_3790,N_3997);
nand U4219 (N_4219,N_3632,N_3541);
or U4220 (N_4220,N_3591,N_3721);
nand U4221 (N_4221,N_3515,N_3953);
and U4222 (N_4222,N_3647,N_3645);
nor U4223 (N_4223,N_3743,N_3950);
or U4224 (N_4224,N_3861,N_3650);
nand U4225 (N_4225,N_3999,N_3603);
or U4226 (N_4226,N_3920,N_3630);
xor U4227 (N_4227,N_3917,N_3709);
and U4228 (N_4228,N_3644,N_3782);
nand U4229 (N_4229,N_3891,N_3703);
nor U4230 (N_4230,N_3916,N_3910);
nor U4231 (N_4231,N_3734,N_3946);
nand U4232 (N_4232,N_3714,N_3680);
nor U4233 (N_4233,N_3617,N_3730);
nand U4234 (N_4234,N_3919,N_3882);
nor U4235 (N_4235,N_3841,N_3901);
and U4236 (N_4236,N_3688,N_3768);
or U4237 (N_4237,N_3872,N_3614);
and U4238 (N_4238,N_3881,N_3655);
and U4239 (N_4239,N_3561,N_3982);
and U4240 (N_4240,N_3979,N_3864);
nand U4241 (N_4241,N_3597,N_3747);
nand U4242 (N_4242,N_3506,N_3885);
or U4243 (N_4243,N_3807,N_3792);
or U4244 (N_4244,N_3606,N_3589);
and U4245 (N_4245,N_3822,N_3615);
and U4246 (N_4246,N_3511,N_3590);
nand U4247 (N_4247,N_3604,N_3929);
nand U4248 (N_4248,N_3608,N_3540);
and U4249 (N_4249,N_3835,N_3720);
and U4250 (N_4250,N_3956,N_3970);
and U4251 (N_4251,N_3996,N_3575);
and U4252 (N_4252,N_3596,N_3726);
or U4253 (N_4253,N_3718,N_3627);
or U4254 (N_4254,N_3668,N_3849);
or U4255 (N_4255,N_3886,N_3750);
and U4256 (N_4256,N_3572,N_3589);
nor U4257 (N_4257,N_3941,N_3802);
and U4258 (N_4258,N_3711,N_3943);
or U4259 (N_4259,N_3531,N_3709);
nor U4260 (N_4260,N_3548,N_3970);
or U4261 (N_4261,N_3595,N_3654);
xor U4262 (N_4262,N_3992,N_3783);
and U4263 (N_4263,N_3888,N_3900);
and U4264 (N_4264,N_3630,N_3906);
nand U4265 (N_4265,N_3902,N_3648);
nand U4266 (N_4266,N_3681,N_3567);
nand U4267 (N_4267,N_3706,N_3806);
nand U4268 (N_4268,N_3699,N_3753);
nor U4269 (N_4269,N_3505,N_3551);
nor U4270 (N_4270,N_3662,N_3505);
or U4271 (N_4271,N_3563,N_3751);
or U4272 (N_4272,N_3580,N_3781);
nand U4273 (N_4273,N_3611,N_3550);
xor U4274 (N_4274,N_3780,N_3922);
xnor U4275 (N_4275,N_3732,N_3512);
or U4276 (N_4276,N_3729,N_3812);
or U4277 (N_4277,N_3848,N_3781);
and U4278 (N_4278,N_3956,N_3691);
nor U4279 (N_4279,N_3867,N_3641);
and U4280 (N_4280,N_3806,N_3842);
nor U4281 (N_4281,N_3748,N_3883);
nor U4282 (N_4282,N_3861,N_3849);
nand U4283 (N_4283,N_3725,N_3755);
nand U4284 (N_4284,N_3841,N_3895);
nor U4285 (N_4285,N_3636,N_3503);
nand U4286 (N_4286,N_3546,N_3722);
and U4287 (N_4287,N_3596,N_3527);
nand U4288 (N_4288,N_3837,N_3970);
and U4289 (N_4289,N_3689,N_3644);
nand U4290 (N_4290,N_3532,N_3744);
and U4291 (N_4291,N_3668,N_3963);
nor U4292 (N_4292,N_3985,N_3507);
and U4293 (N_4293,N_3662,N_3689);
nand U4294 (N_4294,N_3999,N_3838);
and U4295 (N_4295,N_3970,N_3527);
and U4296 (N_4296,N_3831,N_3652);
xor U4297 (N_4297,N_3505,N_3971);
or U4298 (N_4298,N_3755,N_3923);
nor U4299 (N_4299,N_3855,N_3874);
xnor U4300 (N_4300,N_3809,N_3850);
nand U4301 (N_4301,N_3692,N_3664);
nor U4302 (N_4302,N_3874,N_3991);
and U4303 (N_4303,N_3894,N_3820);
and U4304 (N_4304,N_3688,N_3981);
nor U4305 (N_4305,N_3686,N_3534);
or U4306 (N_4306,N_3718,N_3703);
or U4307 (N_4307,N_3972,N_3713);
nor U4308 (N_4308,N_3873,N_3583);
nand U4309 (N_4309,N_3727,N_3584);
nand U4310 (N_4310,N_3715,N_3878);
nor U4311 (N_4311,N_3534,N_3898);
nor U4312 (N_4312,N_3646,N_3753);
nand U4313 (N_4313,N_3856,N_3610);
xnor U4314 (N_4314,N_3925,N_3587);
nor U4315 (N_4315,N_3531,N_3949);
or U4316 (N_4316,N_3640,N_3523);
and U4317 (N_4317,N_3959,N_3564);
nor U4318 (N_4318,N_3901,N_3643);
nor U4319 (N_4319,N_3576,N_3808);
or U4320 (N_4320,N_3892,N_3802);
and U4321 (N_4321,N_3968,N_3563);
nand U4322 (N_4322,N_3926,N_3517);
nor U4323 (N_4323,N_3909,N_3956);
nor U4324 (N_4324,N_3551,N_3900);
nor U4325 (N_4325,N_3601,N_3734);
and U4326 (N_4326,N_3795,N_3864);
nand U4327 (N_4327,N_3951,N_3605);
nand U4328 (N_4328,N_3786,N_3610);
nand U4329 (N_4329,N_3561,N_3885);
nor U4330 (N_4330,N_3967,N_3839);
xor U4331 (N_4331,N_3639,N_3897);
or U4332 (N_4332,N_3978,N_3690);
xnor U4333 (N_4333,N_3793,N_3850);
nand U4334 (N_4334,N_3825,N_3730);
nand U4335 (N_4335,N_3517,N_3591);
nor U4336 (N_4336,N_3859,N_3657);
and U4337 (N_4337,N_3689,N_3681);
nor U4338 (N_4338,N_3679,N_3585);
nor U4339 (N_4339,N_3695,N_3559);
nor U4340 (N_4340,N_3565,N_3863);
and U4341 (N_4341,N_3743,N_3692);
and U4342 (N_4342,N_3838,N_3925);
nand U4343 (N_4343,N_3909,N_3766);
nand U4344 (N_4344,N_3503,N_3678);
xnor U4345 (N_4345,N_3666,N_3728);
nor U4346 (N_4346,N_3646,N_3989);
nor U4347 (N_4347,N_3929,N_3808);
nand U4348 (N_4348,N_3947,N_3765);
or U4349 (N_4349,N_3800,N_3950);
or U4350 (N_4350,N_3650,N_3691);
and U4351 (N_4351,N_3575,N_3708);
and U4352 (N_4352,N_3716,N_3877);
or U4353 (N_4353,N_3533,N_3576);
or U4354 (N_4354,N_3812,N_3737);
or U4355 (N_4355,N_3771,N_3761);
nand U4356 (N_4356,N_3686,N_3703);
or U4357 (N_4357,N_3735,N_3552);
nand U4358 (N_4358,N_3626,N_3728);
nor U4359 (N_4359,N_3694,N_3945);
xnor U4360 (N_4360,N_3596,N_3781);
xnor U4361 (N_4361,N_3748,N_3754);
or U4362 (N_4362,N_3983,N_3729);
nand U4363 (N_4363,N_3560,N_3956);
nand U4364 (N_4364,N_3609,N_3562);
or U4365 (N_4365,N_3743,N_3619);
nor U4366 (N_4366,N_3579,N_3744);
nor U4367 (N_4367,N_3804,N_3846);
nand U4368 (N_4368,N_3761,N_3786);
nor U4369 (N_4369,N_3594,N_3551);
and U4370 (N_4370,N_3764,N_3835);
and U4371 (N_4371,N_3689,N_3986);
nor U4372 (N_4372,N_3674,N_3835);
nand U4373 (N_4373,N_3691,N_3898);
and U4374 (N_4374,N_3972,N_3531);
xnor U4375 (N_4375,N_3784,N_3653);
nand U4376 (N_4376,N_3762,N_3924);
or U4377 (N_4377,N_3754,N_3963);
and U4378 (N_4378,N_3647,N_3694);
nand U4379 (N_4379,N_3604,N_3880);
nand U4380 (N_4380,N_3665,N_3723);
xor U4381 (N_4381,N_3716,N_3785);
and U4382 (N_4382,N_3639,N_3708);
nand U4383 (N_4383,N_3878,N_3779);
or U4384 (N_4384,N_3564,N_3598);
or U4385 (N_4385,N_3963,N_3775);
or U4386 (N_4386,N_3777,N_3566);
nand U4387 (N_4387,N_3587,N_3919);
and U4388 (N_4388,N_3729,N_3800);
and U4389 (N_4389,N_3860,N_3543);
nor U4390 (N_4390,N_3658,N_3842);
and U4391 (N_4391,N_3728,N_3920);
and U4392 (N_4392,N_3678,N_3763);
or U4393 (N_4393,N_3828,N_3784);
xnor U4394 (N_4394,N_3879,N_3757);
nand U4395 (N_4395,N_3797,N_3549);
and U4396 (N_4396,N_3668,N_3737);
nor U4397 (N_4397,N_3765,N_3833);
and U4398 (N_4398,N_3809,N_3913);
and U4399 (N_4399,N_3701,N_3958);
and U4400 (N_4400,N_3928,N_3850);
xnor U4401 (N_4401,N_3820,N_3672);
or U4402 (N_4402,N_3503,N_3801);
xnor U4403 (N_4403,N_3682,N_3987);
and U4404 (N_4404,N_3940,N_3799);
nand U4405 (N_4405,N_3514,N_3504);
or U4406 (N_4406,N_3713,N_3791);
nor U4407 (N_4407,N_3626,N_3870);
nand U4408 (N_4408,N_3522,N_3530);
nand U4409 (N_4409,N_3950,N_3753);
nor U4410 (N_4410,N_3828,N_3977);
and U4411 (N_4411,N_3851,N_3674);
and U4412 (N_4412,N_3909,N_3901);
nand U4413 (N_4413,N_3836,N_3709);
nor U4414 (N_4414,N_3977,N_3675);
or U4415 (N_4415,N_3555,N_3904);
nor U4416 (N_4416,N_3579,N_3682);
nand U4417 (N_4417,N_3922,N_3786);
nor U4418 (N_4418,N_3507,N_3728);
nor U4419 (N_4419,N_3625,N_3799);
and U4420 (N_4420,N_3912,N_3565);
nor U4421 (N_4421,N_3738,N_3723);
and U4422 (N_4422,N_3812,N_3578);
nor U4423 (N_4423,N_3629,N_3506);
or U4424 (N_4424,N_3878,N_3833);
or U4425 (N_4425,N_3599,N_3554);
and U4426 (N_4426,N_3926,N_3875);
or U4427 (N_4427,N_3508,N_3614);
nor U4428 (N_4428,N_3880,N_3964);
nand U4429 (N_4429,N_3830,N_3641);
xnor U4430 (N_4430,N_3787,N_3943);
or U4431 (N_4431,N_3913,N_3861);
xnor U4432 (N_4432,N_3898,N_3802);
nor U4433 (N_4433,N_3911,N_3636);
or U4434 (N_4434,N_3585,N_3598);
and U4435 (N_4435,N_3549,N_3595);
nand U4436 (N_4436,N_3678,N_3857);
nor U4437 (N_4437,N_3870,N_3756);
nand U4438 (N_4438,N_3801,N_3540);
or U4439 (N_4439,N_3704,N_3606);
nor U4440 (N_4440,N_3957,N_3885);
or U4441 (N_4441,N_3586,N_3924);
nor U4442 (N_4442,N_3547,N_3978);
nor U4443 (N_4443,N_3931,N_3862);
or U4444 (N_4444,N_3525,N_3732);
or U4445 (N_4445,N_3625,N_3798);
xnor U4446 (N_4446,N_3534,N_3967);
and U4447 (N_4447,N_3631,N_3603);
or U4448 (N_4448,N_3629,N_3915);
nand U4449 (N_4449,N_3924,N_3751);
nor U4450 (N_4450,N_3783,N_3626);
nand U4451 (N_4451,N_3546,N_3554);
and U4452 (N_4452,N_3589,N_3912);
nor U4453 (N_4453,N_3520,N_3976);
nor U4454 (N_4454,N_3633,N_3878);
nand U4455 (N_4455,N_3983,N_3529);
and U4456 (N_4456,N_3899,N_3566);
nor U4457 (N_4457,N_3661,N_3756);
nand U4458 (N_4458,N_3829,N_3724);
xnor U4459 (N_4459,N_3898,N_3731);
nor U4460 (N_4460,N_3610,N_3971);
or U4461 (N_4461,N_3653,N_3603);
nor U4462 (N_4462,N_3706,N_3857);
xnor U4463 (N_4463,N_3984,N_3761);
xnor U4464 (N_4464,N_3957,N_3784);
nor U4465 (N_4465,N_3636,N_3886);
nand U4466 (N_4466,N_3584,N_3811);
and U4467 (N_4467,N_3878,N_3784);
nand U4468 (N_4468,N_3819,N_3697);
xnor U4469 (N_4469,N_3564,N_3696);
xor U4470 (N_4470,N_3538,N_3719);
nand U4471 (N_4471,N_3735,N_3804);
and U4472 (N_4472,N_3555,N_3615);
and U4473 (N_4473,N_3874,N_3841);
or U4474 (N_4474,N_3840,N_3539);
and U4475 (N_4475,N_3976,N_3612);
and U4476 (N_4476,N_3979,N_3729);
nand U4477 (N_4477,N_3985,N_3916);
nor U4478 (N_4478,N_3826,N_3711);
and U4479 (N_4479,N_3639,N_3909);
nor U4480 (N_4480,N_3962,N_3865);
xnor U4481 (N_4481,N_3809,N_3714);
and U4482 (N_4482,N_3636,N_3735);
nand U4483 (N_4483,N_3861,N_3955);
xor U4484 (N_4484,N_3882,N_3686);
nor U4485 (N_4485,N_3542,N_3503);
nand U4486 (N_4486,N_3735,N_3810);
nand U4487 (N_4487,N_3992,N_3656);
nor U4488 (N_4488,N_3590,N_3677);
xnor U4489 (N_4489,N_3558,N_3964);
nor U4490 (N_4490,N_3854,N_3666);
nand U4491 (N_4491,N_3697,N_3730);
nand U4492 (N_4492,N_3516,N_3872);
nand U4493 (N_4493,N_3980,N_3557);
nor U4494 (N_4494,N_3819,N_3512);
and U4495 (N_4495,N_3748,N_3659);
nor U4496 (N_4496,N_3721,N_3603);
and U4497 (N_4497,N_3914,N_3783);
nor U4498 (N_4498,N_3889,N_3756);
or U4499 (N_4499,N_3785,N_3883);
nor U4500 (N_4500,N_4187,N_4367);
nand U4501 (N_4501,N_4226,N_4119);
nor U4502 (N_4502,N_4484,N_4079);
and U4503 (N_4503,N_4212,N_4113);
nor U4504 (N_4504,N_4160,N_4370);
nand U4505 (N_4505,N_4068,N_4085);
nand U4506 (N_4506,N_4291,N_4275);
xor U4507 (N_4507,N_4034,N_4258);
nand U4508 (N_4508,N_4358,N_4305);
nor U4509 (N_4509,N_4324,N_4178);
and U4510 (N_4510,N_4394,N_4237);
nand U4511 (N_4511,N_4309,N_4111);
xnor U4512 (N_4512,N_4014,N_4452);
xnor U4513 (N_4513,N_4015,N_4363);
xnor U4514 (N_4514,N_4061,N_4333);
or U4515 (N_4515,N_4292,N_4118);
and U4516 (N_4516,N_4415,N_4441);
nand U4517 (N_4517,N_4209,N_4255);
nand U4518 (N_4518,N_4283,N_4169);
or U4519 (N_4519,N_4130,N_4244);
or U4520 (N_4520,N_4284,N_4143);
nand U4521 (N_4521,N_4485,N_4185);
or U4522 (N_4522,N_4449,N_4002);
or U4523 (N_4523,N_4408,N_4482);
nor U4524 (N_4524,N_4004,N_4091);
or U4525 (N_4525,N_4062,N_4134);
or U4526 (N_4526,N_4461,N_4201);
nor U4527 (N_4527,N_4121,N_4387);
nor U4528 (N_4528,N_4181,N_4194);
nor U4529 (N_4529,N_4268,N_4375);
and U4530 (N_4530,N_4391,N_4246);
nand U4531 (N_4531,N_4000,N_4364);
nor U4532 (N_4532,N_4256,N_4158);
xor U4533 (N_4533,N_4139,N_4260);
nor U4534 (N_4534,N_4023,N_4017);
nor U4535 (N_4535,N_4058,N_4208);
or U4536 (N_4536,N_4137,N_4193);
or U4537 (N_4537,N_4196,N_4459);
or U4538 (N_4538,N_4280,N_4142);
or U4539 (N_4539,N_4400,N_4050);
and U4540 (N_4540,N_4307,N_4145);
and U4541 (N_4541,N_4301,N_4006);
nor U4542 (N_4542,N_4042,N_4164);
or U4543 (N_4543,N_4293,N_4312);
or U4544 (N_4544,N_4077,N_4320);
xnor U4545 (N_4545,N_4218,N_4135);
nand U4546 (N_4546,N_4426,N_4192);
and U4547 (N_4547,N_4342,N_4317);
xnor U4548 (N_4548,N_4427,N_4205);
nand U4549 (N_4549,N_4016,N_4089);
nand U4550 (N_4550,N_4419,N_4176);
nor U4551 (N_4551,N_4378,N_4323);
xor U4552 (N_4552,N_4344,N_4490);
and U4553 (N_4553,N_4269,N_4381);
nor U4554 (N_4554,N_4368,N_4242);
xnor U4555 (N_4555,N_4392,N_4157);
or U4556 (N_4556,N_4414,N_4172);
or U4557 (N_4557,N_4125,N_4099);
and U4558 (N_4558,N_4264,N_4182);
or U4559 (N_4559,N_4345,N_4083);
and U4560 (N_4560,N_4100,N_4273);
or U4561 (N_4561,N_4456,N_4369);
or U4562 (N_4562,N_4147,N_4313);
nand U4563 (N_4563,N_4090,N_4314);
or U4564 (N_4564,N_4350,N_4362);
and U4565 (N_4565,N_4155,N_4202);
nand U4566 (N_4566,N_4156,N_4318);
and U4567 (N_4567,N_4270,N_4476);
and U4568 (N_4568,N_4086,N_4123);
nor U4569 (N_4569,N_4465,N_4039);
nor U4570 (N_4570,N_4153,N_4472);
and U4571 (N_4571,N_4055,N_4027);
and U4572 (N_4572,N_4230,N_4478);
nand U4573 (N_4573,N_4433,N_4340);
or U4574 (N_4574,N_4330,N_4332);
nor U4575 (N_4575,N_4003,N_4491);
or U4576 (N_4576,N_4132,N_4140);
and U4577 (N_4577,N_4019,N_4326);
or U4578 (N_4578,N_4278,N_4257);
and U4579 (N_4579,N_4217,N_4435);
nand U4580 (N_4580,N_4437,N_4442);
and U4581 (N_4581,N_4447,N_4424);
nand U4582 (N_4582,N_4057,N_4087);
nand U4583 (N_4583,N_4163,N_4168);
nand U4584 (N_4584,N_4009,N_4227);
and U4585 (N_4585,N_4239,N_4029);
nand U4586 (N_4586,N_4379,N_4167);
or U4587 (N_4587,N_4306,N_4060);
and U4588 (N_4588,N_4216,N_4298);
or U4589 (N_4589,N_4428,N_4366);
nor U4590 (N_4590,N_4390,N_4251);
or U4591 (N_4591,N_4046,N_4287);
and U4592 (N_4592,N_4277,N_4436);
nand U4593 (N_4593,N_4474,N_4468);
or U4594 (N_4594,N_4117,N_4316);
and U4595 (N_4595,N_4174,N_4215);
nand U4596 (N_4596,N_4049,N_4081);
or U4597 (N_4597,N_4114,N_4041);
nor U4598 (N_4598,N_4297,N_4021);
and U4599 (N_4599,N_4497,N_4299);
nor U4600 (N_4600,N_4223,N_4036);
and U4601 (N_4601,N_4093,N_4190);
or U4602 (N_4602,N_4078,N_4303);
and U4603 (N_4603,N_4043,N_4346);
or U4604 (N_4604,N_4460,N_4098);
nor U4605 (N_4605,N_4007,N_4388);
nor U4606 (N_4606,N_4161,N_4282);
and U4607 (N_4607,N_4254,N_4035);
and U4608 (N_4608,N_4372,N_4249);
nor U4609 (N_4609,N_4067,N_4229);
nand U4610 (N_4610,N_4066,N_4302);
and U4611 (N_4611,N_4177,N_4065);
xor U4612 (N_4612,N_4040,N_4146);
and U4613 (N_4613,N_4235,N_4294);
and U4614 (N_4614,N_4071,N_4179);
or U4615 (N_4615,N_4399,N_4496);
or U4616 (N_4616,N_4262,N_4470);
nor U4617 (N_4617,N_4233,N_4354);
nor U4618 (N_4618,N_4411,N_4115);
or U4619 (N_4619,N_4353,N_4386);
nand U4620 (N_4620,N_4197,N_4383);
or U4621 (N_4621,N_4234,N_4469);
or U4622 (N_4622,N_4148,N_4325);
or U4623 (N_4623,N_4311,N_4393);
or U4624 (N_4624,N_4175,N_4195);
or U4625 (N_4625,N_4150,N_4170);
nand U4626 (N_4626,N_4418,N_4250);
or U4627 (N_4627,N_4127,N_4462);
and U4628 (N_4628,N_4453,N_4281);
and U4629 (N_4629,N_4231,N_4110);
and U4630 (N_4630,N_4487,N_4339);
xor U4631 (N_4631,N_4048,N_4104);
and U4632 (N_4632,N_4052,N_4319);
and U4633 (N_4633,N_4495,N_4450);
nand U4634 (N_4634,N_4022,N_4038);
and U4635 (N_4635,N_4008,N_4095);
or U4636 (N_4636,N_4493,N_4329);
nand U4637 (N_4637,N_4405,N_4094);
nand U4638 (N_4638,N_4219,N_4051);
nor U4639 (N_4639,N_4421,N_4225);
nor U4640 (N_4640,N_4102,N_4337);
xor U4641 (N_4641,N_4471,N_4165);
nor U4642 (N_4642,N_4096,N_4413);
xnor U4643 (N_4643,N_4211,N_4253);
nor U4644 (N_4644,N_4131,N_4045);
or U4645 (N_4645,N_4455,N_4206);
or U4646 (N_4646,N_4431,N_4376);
and U4647 (N_4647,N_4024,N_4488);
xor U4648 (N_4648,N_4109,N_4276);
nor U4649 (N_4649,N_4289,N_4241);
and U4650 (N_4650,N_4389,N_4037);
and U4651 (N_4651,N_4259,N_4236);
and U4652 (N_4652,N_4116,N_4184);
nor U4653 (N_4653,N_4285,N_4010);
and U4654 (N_4654,N_4076,N_4152);
nand U4655 (N_4655,N_4341,N_4434);
nor U4656 (N_4656,N_4397,N_4440);
xnor U4657 (N_4657,N_4444,N_4401);
and U4658 (N_4658,N_4012,N_4047);
or U4659 (N_4659,N_4124,N_4028);
or U4660 (N_4660,N_4238,N_4467);
or U4661 (N_4661,N_4213,N_4483);
or U4662 (N_4662,N_4290,N_4108);
and U4663 (N_4663,N_4265,N_4018);
nor U4664 (N_4664,N_4097,N_4183);
and U4665 (N_4665,N_4360,N_4141);
or U4666 (N_4666,N_4310,N_4013);
nand U4667 (N_4667,N_4128,N_4033);
and U4668 (N_4668,N_4056,N_4331);
and U4669 (N_4669,N_4343,N_4308);
xor U4670 (N_4670,N_4448,N_4479);
and U4671 (N_4671,N_4423,N_4221);
and U4672 (N_4672,N_4365,N_4220);
nand U4673 (N_4673,N_4166,N_4189);
nor U4674 (N_4674,N_4247,N_4486);
and U4675 (N_4675,N_4382,N_4429);
nor U4676 (N_4676,N_4336,N_4347);
nor U4677 (N_4677,N_4425,N_4328);
xnor U4678 (N_4678,N_4443,N_4224);
nand U4679 (N_4679,N_4410,N_4480);
and U4680 (N_4680,N_4371,N_4191);
and U4681 (N_4681,N_4261,N_4240);
nand U4682 (N_4682,N_4171,N_4481);
nand U4683 (N_4683,N_4355,N_4199);
nand U4684 (N_4684,N_4466,N_4475);
nor U4685 (N_4685,N_4031,N_4420);
nor U4686 (N_4686,N_4126,N_4300);
nand U4687 (N_4687,N_4001,N_4489);
nor U4688 (N_4688,N_4377,N_4112);
or U4689 (N_4689,N_4069,N_4458);
nor U4690 (N_4690,N_4129,N_4074);
nand U4691 (N_4691,N_4477,N_4451);
or U4692 (N_4692,N_4356,N_4499);
nor U4693 (N_4693,N_4214,N_4385);
or U4694 (N_4694,N_4151,N_4403);
nand U4695 (N_4695,N_4080,N_4416);
and U4696 (N_4696,N_4186,N_4138);
nand U4697 (N_4697,N_4073,N_4295);
nor U4698 (N_4698,N_4200,N_4082);
xor U4699 (N_4699,N_4267,N_4279);
nor U4700 (N_4700,N_4228,N_4384);
and U4701 (N_4701,N_4180,N_4266);
nand U4702 (N_4702,N_4120,N_4334);
nand U4703 (N_4703,N_4188,N_4054);
nand U4704 (N_4704,N_4407,N_4232);
and U4705 (N_4705,N_4296,N_4286);
nand U4706 (N_4706,N_4044,N_4063);
and U4707 (N_4707,N_4088,N_4136);
nor U4708 (N_4708,N_4106,N_4122);
xor U4709 (N_4709,N_4430,N_4473);
and U4710 (N_4710,N_4105,N_4322);
nand U4711 (N_4711,N_4396,N_4026);
nand U4712 (N_4712,N_4454,N_4272);
nand U4713 (N_4713,N_4494,N_4315);
nand U4714 (N_4714,N_4075,N_4133);
and U4715 (N_4715,N_4338,N_4432);
and U4716 (N_4716,N_4103,N_4263);
nor U4717 (N_4717,N_4304,N_4207);
xor U4718 (N_4718,N_4445,N_4417);
nor U4719 (N_4719,N_4457,N_4351);
or U4720 (N_4720,N_4498,N_4020);
nor U4721 (N_4721,N_4101,N_4348);
nor U4722 (N_4722,N_4374,N_4398);
nand U4723 (N_4723,N_4271,N_4162);
and U4724 (N_4724,N_4422,N_4025);
nand U4725 (N_4725,N_4404,N_4154);
or U4726 (N_4726,N_4463,N_4357);
xor U4727 (N_4727,N_4438,N_4072);
or U4728 (N_4728,N_4053,N_4059);
and U4729 (N_4729,N_4248,N_4274);
nand U4730 (N_4730,N_4107,N_4159);
and U4731 (N_4731,N_4203,N_4361);
nand U4732 (N_4732,N_4464,N_4252);
nand U4733 (N_4733,N_4380,N_4064);
nor U4734 (N_4734,N_4149,N_4288);
nor U4735 (N_4735,N_4349,N_4412);
nor U4736 (N_4736,N_4409,N_4005);
or U4737 (N_4737,N_4243,N_4373);
and U4738 (N_4738,N_4245,N_4210);
nor U4739 (N_4739,N_4030,N_4395);
nor U4740 (N_4740,N_4204,N_4446);
nor U4741 (N_4741,N_4144,N_4321);
nand U4742 (N_4742,N_4327,N_4352);
or U4743 (N_4743,N_4084,N_4173);
nor U4744 (N_4744,N_4222,N_4032);
or U4745 (N_4745,N_4011,N_4359);
xor U4746 (N_4746,N_4198,N_4492);
or U4747 (N_4747,N_4070,N_4402);
nand U4748 (N_4748,N_4335,N_4406);
nand U4749 (N_4749,N_4092,N_4439);
or U4750 (N_4750,N_4384,N_4273);
nor U4751 (N_4751,N_4078,N_4425);
or U4752 (N_4752,N_4408,N_4276);
and U4753 (N_4753,N_4244,N_4488);
xor U4754 (N_4754,N_4038,N_4037);
nand U4755 (N_4755,N_4272,N_4010);
nand U4756 (N_4756,N_4074,N_4027);
nor U4757 (N_4757,N_4386,N_4426);
nand U4758 (N_4758,N_4485,N_4233);
or U4759 (N_4759,N_4071,N_4362);
xnor U4760 (N_4760,N_4454,N_4390);
nand U4761 (N_4761,N_4301,N_4278);
nand U4762 (N_4762,N_4349,N_4108);
and U4763 (N_4763,N_4049,N_4367);
and U4764 (N_4764,N_4309,N_4468);
nand U4765 (N_4765,N_4083,N_4064);
or U4766 (N_4766,N_4388,N_4487);
or U4767 (N_4767,N_4264,N_4169);
or U4768 (N_4768,N_4202,N_4006);
and U4769 (N_4769,N_4369,N_4060);
nand U4770 (N_4770,N_4357,N_4443);
or U4771 (N_4771,N_4199,N_4246);
nand U4772 (N_4772,N_4478,N_4174);
and U4773 (N_4773,N_4394,N_4126);
or U4774 (N_4774,N_4304,N_4392);
or U4775 (N_4775,N_4189,N_4337);
and U4776 (N_4776,N_4357,N_4314);
nor U4777 (N_4777,N_4119,N_4246);
and U4778 (N_4778,N_4384,N_4178);
nand U4779 (N_4779,N_4314,N_4258);
xnor U4780 (N_4780,N_4420,N_4180);
nor U4781 (N_4781,N_4444,N_4153);
and U4782 (N_4782,N_4081,N_4267);
or U4783 (N_4783,N_4276,N_4439);
nor U4784 (N_4784,N_4102,N_4313);
nand U4785 (N_4785,N_4289,N_4183);
nor U4786 (N_4786,N_4116,N_4123);
nor U4787 (N_4787,N_4177,N_4441);
nor U4788 (N_4788,N_4235,N_4400);
nor U4789 (N_4789,N_4218,N_4367);
nor U4790 (N_4790,N_4087,N_4031);
nand U4791 (N_4791,N_4103,N_4376);
and U4792 (N_4792,N_4344,N_4017);
and U4793 (N_4793,N_4356,N_4451);
nand U4794 (N_4794,N_4227,N_4120);
and U4795 (N_4795,N_4055,N_4459);
xnor U4796 (N_4796,N_4014,N_4245);
nand U4797 (N_4797,N_4231,N_4413);
nand U4798 (N_4798,N_4113,N_4255);
nand U4799 (N_4799,N_4155,N_4350);
nor U4800 (N_4800,N_4352,N_4397);
xor U4801 (N_4801,N_4170,N_4253);
nor U4802 (N_4802,N_4200,N_4227);
or U4803 (N_4803,N_4061,N_4474);
or U4804 (N_4804,N_4477,N_4465);
nor U4805 (N_4805,N_4092,N_4253);
or U4806 (N_4806,N_4225,N_4254);
and U4807 (N_4807,N_4167,N_4238);
xor U4808 (N_4808,N_4159,N_4042);
or U4809 (N_4809,N_4167,N_4458);
nand U4810 (N_4810,N_4233,N_4199);
or U4811 (N_4811,N_4036,N_4039);
xor U4812 (N_4812,N_4357,N_4473);
or U4813 (N_4813,N_4026,N_4060);
or U4814 (N_4814,N_4339,N_4387);
xor U4815 (N_4815,N_4428,N_4226);
nor U4816 (N_4816,N_4160,N_4420);
and U4817 (N_4817,N_4112,N_4291);
or U4818 (N_4818,N_4268,N_4178);
xnor U4819 (N_4819,N_4118,N_4019);
nor U4820 (N_4820,N_4472,N_4273);
nand U4821 (N_4821,N_4428,N_4253);
and U4822 (N_4822,N_4326,N_4161);
and U4823 (N_4823,N_4203,N_4208);
nor U4824 (N_4824,N_4101,N_4195);
or U4825 (N_4825,N_4031,N_4248);
and U4826 (N_4826,N_4205,N_4079);
xnor U4827 (N_4827,N_4105,N_4193);
nor U4828 (N_4828,N_4497,N_4188);
and U4829 (N_4829,N_4357,N_4305);
or U4830 (N_4830,N_4466,N_4013);
and U4831 (N_4831,N_4295,N_4271);
or U4832 (N_4832,N_4051,N_4343);
or U4833 (N_4833,N_4081,N_4454);
or U4834 (N_4834,N_4417,N_4264);
nor U4835 (N_4835,N_4403,N_4116);
nand U4836 (N_4836,N_4299,N_4118);
nand U4837 (N_4837,N_4155,N_4140);
or U4838 (N_4838,N_4475,N_4012);
nand U4839 (N_4839,N_4156,N_4246);
and U4840 (N_4840,N_4108,N_4211);
and U4841 (N_4841,N_4233,N_4096);
xor U4842 (N_4842,N_4110,N_4101);
xnor U4843 (N_4843,N_4288,N_4048);
nor U4844 (N_4844,N_4286,N_4350);
nor U4845 (N_4845,N_4238,N_4341);
or U4846 (N_4846,N_4061,N_4194);
nor U4847 (N_4847,N_4083,N_4410);
and U4848 (N_4848,N_4109,N_4425);
nand U4849 (N_4849,N_4151,N_4154);
or U4850 (N_4850,N_4240,N_4215);
nor U4851 (N_4851,N_4175,N_4007);
and U4852 (N_4852,N_4482,N_4268);
and U4853 (N_4853,N_4461,N_4070);
and U4854 (N_4854,N_4104,N_4365);
or U4855 (N_4855,N_4476,N_4170);
xnor U4856 (N_4856,N_4158,N_4277);
nor U4857 (N_4857,N_4301,N_4080);
nor U4858 (N_4858,N_4424,N_4415);
or U4859 (N_4859,N_4104,N_4275);
and U4860 (N_4860,N_4353,N_4380);
nand U4861 (N_4861,N_4440,N_4352);
xor U4862 (N_4862,N_4043,N_4488);
nor U4863 (N_4863,N_4320,N_4235);
nor U4864 (N_4864,N_4215,N_4201);
nor U4865 (N_4865,N_4117,N_4063);
and U4866 (N_4866,N_4423,N_4051);
and U4867 (N_4867,N_4444,N_4497);
or U4868 (N_4868,N_4235,N_4006);
nand U4869 (N_4869,N_4031,N_4006);
or U4870 (N_4870,N_4233,N_4385);
or U4871 (N_4871,N_4382,N_4129);
and U4872 (N_4872,N_4372,N_4214);
nor U4873 (N_4873,N_4126,N_4123);
or U4874 (N_4874,N_4044,N_4489);
nor U4875 (N_4875,N_4270,N_4423);
nor U4876 (N_4876,N_4342,N_4213);
nor U4877 (N_4877,N_4142,N_4485);
xnor U4878 (N_4878,N_4114,N_4260);
or U4879 (N_4879,N_4158,N_4253);
and U4880 (N_4880,N_4486,N_4010);
nand U4881 (N_4881,N_4293,N_4276);
nor U4882 (N_4882,N_4194,N_4179);
or U4883 (N_4883,N_4355,N_4253);
xor U4884 (N_4884,N_4157,N_4201);
or U4885 (N_4885,N_4493,N_4298);
nand U4886 (N_4886,N_4476,N_4311);
and U4887 (N_4887,N_4330,N_4392);
or U4888 (N_4888,N_4270,N_4060);
nand U4889 (N_4889,N_4214,N_4074);
nand U4890 (N_4890,N_4145,N_4211);
and U4891 (N_4891,N_4231,N_4295);
nand U4892 (N_4892,N_4404,N_4195);
nor U4893 (N_4893,N_4422,N_4055);
nand U4894 (N_4894,N_4166,N_4370);
nor U4895 (N_4895,N_4468,N_4139);
xnor U4896 (N_4896,N_4163,N_4109);
nand U4897 (N_4897,N_4060,N_4313);
nor U4898 (N_4898,N_4441,N_4020);
or U4899 (N_4899,N_4492,N_4177);
nor U4900 (N_4900,N_4400,N_4242);
nor U4901 (N_4901,N_4122,N_4152);
and U4902 (N_4902,N_4434,N_4279);
nor U4903 (N_4903,N_4491,N_4499);
nand U4904 (N_4904,N_4265,N_4044);
and U4905 (N_4905,N_4210,N_4059);
or U4906 (N_4906,N_4426,N_4131);
nand U4907 (N_4907,N_4085,N_4383);
nand U4908 (N_4908,N_4337,N_4227);
and U4909 (N_4909,N_4078,N_4473);
nand U4910 (N_4910,N_4018,N_4136);
nor U4911 (N_4911,N_4200,N_4009);
nand U4912 (N_4912,N_4185,N_4489);
and U4913 (N_4913,N_4407,N_4314);
and U4914 (N_4914,N_4340,N_4387);
and U4915 (N_4915,N_4421,N_4128);
or U4916 (N_4916,N_4104,N_4469);
nand U4917 (N_4917,N_4236,N_4328);
and U4918 (N_4918,N_4298,N_4277);
and U4919 (N_4919,N_4077,N_4398);
nor U4920 (N_4920,N_4209,N_4176);
or U4921 (N_4921,N_4301,N_4427);
or U4922 (N_4922,N_4039,N_4002);
and U4923 (N_4923,N_4322,N_4407);
or U4924 (N_4924,N_4052,N_4216);
and U4925 (N_4925,N_4437,N_4467);
and U4926 (N_4926,N_4277,N_4349);
nor U4927 (N_4927,N_4029,N_4213);
and U4928 (N_4928,N_4127,N_4180);
nor U4929 (N_4929,N_4139,N_4362);
or U4930 (N_4930,N_4392,N_4488);
nand U4931 (N_4931,N_4243,N_4167);
nor U4932 (N_4932,N_4142,N_4187);
or U4933 (N_4933,N_4029,N_4485);
nor U4934 (N_4934,N_4082,N_4067);
or U4935 (N_4935,N_4394,N_4260);
and U4936 (N_4936,N_4258,N_4476);
and U4937 (N_4937,N_4296,N_4430);
nand U4938 (N_4938,N_4140,N_4225);
nand U4939 (N_4939,N_4184,N_4244);
and U4940 (N_4940,N_4082,N_4236);
or U4941 (N_4941,N_4138,N_4350);
nor U4942 (N_4942,N_4383,N_4309);
nor U4943 (N_4943,N_4254,N_4167);
nor U4944 (N_4944,N_4117,N_4399);
or U4945 (N_4945,N_4092,N_4334);
or U4946 (N_4946,N_4028,N_4018);
nor U4947 (N_4947,N_4365,N_4447);
or U4948 (N_4948,N_4040,N_4409);
nor U4949 (N_4949,N_4223,N_4028);
xor U4950 (N_4950,N_4176,N_4341);
nor U4951 (N_4951,N_4390,N_4346);
and U4952 (N_4952,N_4117,N_4478);
nor U4953 (N_4953,N_4418,N_4309);
or U4954 (N_4954,N_4320,N_4229);
xor U4955 (N_4955,N_4193,N_4273);
and U4956 (N_4956,N_4408,N_4427);
nand U4957 (N_4957,N_4288,N_4147);
and U4958 (N_4958,N_4364,N_4385);
nor U4959 (N_4959,N_4219,N_4354);
and U4960 (N_4960,N_4177,N_4068);
and U4961 (N_4961,N_4032,N_4428);
and U4962 (N_4962,N_4020,N_4197);
nand U4963 (N_4963,N_4357,N_4062);
and U4964 (N_4964,N_4179,N_4085);
nor U4965 (N_4965,N_4145,N_4329);
and U4966 (N_4966,N_4168,N_4048);
or U4967 (N_4967,N_4443,N_4372);
and U4968 (N_4968,N_4372,N_4081);
nand U4969 (N_4969,N_4290,N_4070);
and U4970 (N_4970,N_4273,N_4440);
and U4971 (N_4971,N_4356,N_4214);
nor U4972 (N_4972,N_4365,N_4295);
and U4973 (N_4973,N_4120,N_4332);
or U4974 (N_4974,N_4271,N_4283);
and U4975 (N_4975,N_4243,N_4453);
nor U4976 (N_4976,N_4096,N_4023);
nor U4977 (N_4977,N_4131,N_4332);
xor U4978 (N_4978,N_4124,N_4045);
or U4979 (N_4979,N_4314,N_4108);
nor U4980 (N_4980,N_4387,N_4436);
and U4981 (N_4981,N_4053,N_4255);
nor U4982 (N_4982,N_4035,N_4267);
and U4983 (N_4983,N_4318,N_4115);
and U4984 (N_4984,N_4032,N_4107);
and U4985 (N_4985,N_4296,N_4111);
nand U4986 (N_4986,N_4365,N_4009);
or U4987 (N_4987,N_4179,N_4361);
or U4988 (N_4988,N_4373,N_4350);
nor U4989 (N_4989,N_4341,N_4015);
or U4990 (N_4990,N_4418,N_4247);
nand U4991 (N_4991,N_4447,N_4436);
nand U4992 (N_4992,N_4219,N_4147);
xnor U4993 (N_4993,N_4452,N_4463);
nand U4994 (N_4994,N_4199,N_4004);
nor U4995 (N_4995,N_4058,N_4350);
nand U4996 (N_4996,N_4081,N_4465);
nor U4997 (N_4997,N_4292,N_4396);
nand U4998 (N_4998,N_4495,N_4077);
nor U4999 (N_4999,N_4015,N_4492);
and U5000 (N_5000,N_4817,N_4902);
or U5001 (N_5001,N_4939,N_4754);
nor U5002 (N_5002,N_4691,N_4608);
nand U5003 (N_5003,N_4912,N_4592);
or U5004 (N_5004,N_4943,N_4709);
and U5005 (N_5005,N_4764,N_4900);
nor U5006 (N_5006,N_4815,N_4671);
nor U5007 (N_5007,N_4700,N_4674);
or U5008 (N_5008,N_4892,N_4903);
and U5009 (N_5009,N_4597,N_4681);
nor U5010 (N_5010,N_4993,N_4779);
nor U5011 (N_5011,N_4868,N_4870);
nor U5012 (N_5012,N_4854,N_4797);
xor U5013 (N_5013,N_4730,N_4734);
and U5014 (N_5014,N_4506,N_4888);
nand U5015 (N_5015,N_4998,N_4917);
xor U5016 (N_5016,N_4517,N_4976);
or U5017 (N_5017,N_4503,N_4559);
and U5018 (N_5018,N_4858,N_4777);
nor U5019 (N_5019,N_4651,N_4839);
nor U5020 (N_5020,N_4873,N_4962);
nor U5021 (N_5021,N_4748,N_4799);
nor U5022 (N_5022,N_4616,N_4585);
nor U5023 (N_5023,N_4621,N_4719);
and U5024 (N_5024,N_4723,N_4812);
nand U5025 (N_5025,N_4987,N_4792);
or U5026 (N_5026,N_4633,N_4964);
nor U5027 (N_5027,N_4869,N_4782);
nor U5028 (N_5028,N_4816,N_4806);
and U5029 (N_5029,N_4599,N_4905);
or U5030 (N_5030,N_4555,N_4743);
nor U5031 (N_5031,N_4500,N_4684);
nand U5032 (N_5032,N_4742,N_4785);
nor U5033 (N_5033,N_4894,N_4514);
or U5034 (N_5034,N_4580,N_4696);
and U5035 (N_5035,N_4531,N_4820);
nand U5036 (N_5036,N_4649,N_4660);
nand U5037 (N_5037,N_4818,N_4955);
and U5038 (N_5038,N_4565,N_4852);
xnor U5039 (N_5039,N_4872,N_4781);
or U5040 (N_5040,N_4529,N_4866);
nand U5041 (N_5041,N_4510,N_4975);
xnor U5042 (N_5042,N_4981,N_4521);
and U5043 (N_5043,N_4647,N_4959);
and U5044 (N_5044,N_4673,N_4803);
nand U5045 (N_5045,N_4766,N_4639);
and U5046 (N_5046,N_4524,N_4931);
and U5047 (N_5047,N_4762,N_4935);
and U5048 (N_5048,N_4724,N_4662);
xnor U5049 (N_5049,N_4740,N_4749);
nand U5050 (N_5050,N_4625,N_4718);
nand U5051 (N_5051,N_4657,N_4927);
nand U5052 (N_5052,N_4688,N_4542);
nand U5053 (N_5053,N_4686,N_4879);
nor U5054 (N_5054,N_4865,N_4945);
and U5055 (N_5055,N_4575,N_4552);
or U5056 (N_5056,N_4741,N_4898);
or U5057 (N_5057,N_4582,N_4827);
and U5058 (N_5058,N_4980,N_4850);
xnor U5059 (N_5059,N_4720,N_4970);
nor U5060 (N_5060,N_4974,N_4677);
nor U5061 (N_5061,N_4971,N_4886);
nand U5062 (N_5062,N_4534,N_4942);
nand U5063 (N_5063,N_4891,N_4563);
or U5064 (N_5064,N_4861,N_4753);
or U5065 (N_5065,N_4775,N_4784);
nor U5066 (N_5066,N_4906,N_4885);
nor U5067 (N_5067,N_4956,N_4910);
and U5068 (N_5068,N_4952,N_4646);
nand U5069 (N_5069,N_4589,N_4508);
nor U5070 (N_5070,N_4533,N_4544);
nor U5071 (N_5071,N_4985,N_4967);
nor U5072 (N_5072,N_4930,N_4667);
and U5073 (N_5073,N_4522,N_4774);
or U5074 (N_5074,N_4561,N_4574);
or U5075 (N_5075,N_4695,N_4591);
or U5076 (N_5076,N_4604,N_4650);
and U5077 (N_5077,N_4876,N_4951);
nor U5078 (N_5078,N_4602,N_4716);
and U5079 (N_5079,N_4972,N_4908);
or U5080 (N_5080,N_4961,N_4750);
nand U5081 (N_5081,N_4822,N_4627);
or U5082 (N_5082,N_4632,N_4505);
nor U5083 (N_5083,N_4658,N_4846);
or U5084 (N_5084,N_4554,N_4793);
and U5085 (N_5085,N_4679,N_4929);
and U5086 (N_5086,N_4562,N_4786);
or U5087 (N_5087,N_4947,N_4540);
xor U5088 (N_5088,N_4566,N_4579);
or U5089 (N_5089,N_4725,N_4832);
nor U5090 (N_5090,N_4539,N_4778);
nand U5091 (N_5091,N_4809,N_4842);
and U5092 (N_5092,N_4810,N_4744);
and U5093 (N_5093,N_4714,N_4954);
nor U5094 (N_5094,N_4613,N_4590);
nor U5095 (N_5095,N_4857,N_4780);
nor U5096 (N_5096,N_4615,N_4761);
nor U5097 (N_5097,N_4635,N_4807);
or U5098 (N_5098,N_4680,N_4884);
or U5099 (N_5099,N_4880,N_4836);
nand U5100 (N_5100,N_4675,N_4641);
nand U5101 (N_5101,N_4864,N_4752);
nand U5102 (N_5102,N_4668,N_4965);
xnor U5103 (N_5103,N_4999,N_4694);
nor U5104 (N_5104,N_4783,N_4701);
or U5105 (N_5105,N_4697,N_4925);
and U5106 (N_5106,N_4811,N_4921);
nor U5107 (N_5107,N_4922,N_4977);
nor U5108 (N_5108,N_4875,N_4571);
nor U5109 (N_5109,N_4946,N_4583);
or U5110 (N_5110,N_4568,N_4835);
nand U5111 (N_5111,N_4705,N_4845);
xor U5112 (N_5112,N_4849,N_4607);
and U5113 (N_5113,N_4731,N_4862);
or U5114 (N_5114,N_4586,N_4746);
and U5115 (N_5115,N_4548,N_4626);
nor U5116 (N_5116,N_4584,N_4509);
nand U5117 (N_5117,N_4682,N_4611);
nand U5118 (N_5118,N_4606,N_4644);
or U5119 (N_5119,N_4881,N_4601);
or U5120 (N_5120,N_4528,N_4572);
and U5121 (N_5121,N_4963,N_4840);
and U5122 (N_5122,N_4907,N_4944);
nand U5123 (N_5123,N_4623,N_4904);
nand U5124 (N_5124,N_4991,N_4543);
or U5125 (N_5125,N_4887,N_4605);
nor U5126 (N_5126,N_4924,N_4769);
xor U5127 (N_5127,N_4859,N_4932);
nand U5128 (N_5128,N_4994,N_4982);
nor U5129 (N_5129,N_4520,N_4655);
nand U5130 (N_5130,N_4739,N_4569);
or U5131 (N_5131,N_4990,N_4989);
nor U5132 (N_5132,N_4899,N_4546);
nand U5133 (N_5133,N_4953,N_4747);
nand U5134 (N_5134,N_4631,N_4598);
and U5135 (N_5135,N_4588,N_4847);
nor U5136 (N_5136,N_4665,N_4823);
or U5137 (N_5137,N_4890,N_4789);
and U5138 (N_5138,N_4513,N_4798);
and U5139 (N_5139,N_4867,N_4794);
or U5140 (N_5140,N_4986,N_4638);
nor U5141 (N_5141,N_4979,N_4830);
xor U5142 (N_5142,N_4594,N_4863);
or U5143 (N_5143,N_4501,N_4897);
xor U5144 (N_5144,N_4919,N_4992);
nand U5145 (N_5145,N_4622,N_4642);
nand U5146 (N_5146,N_4648,N_4895);
or U5147 (N_5147,N_4983,N_4997);
and U5148 (N_5148,N_4729,N_4853);
xor U5149 (N_5149,N_4715,N_4703);
nand U5150 (N_5150,N_4771,N_4670);
xnor U5151 (N_5151,N_4536,N_4988);
and U5152 (N_5152,N_4848,N_4577);
and U5153 (N_5153,N_4504,N_4636);
and U5154 (N_5154,N_4690,N_4664);
or U5155 (N_5155,N_4511,N_4883);
nor U5156 (N_5156,N_4519,N_4802);
and U5157 (N_5157,N_4957,N_4530);
xor U5158 (N_5158,N_4918,N_4507);
xor U5159 (N_5159,N_4814,N_4527);
nand U5160 (N_5160,N_4958,N_4717);
nand U5161 (N_5161,N_4707,N_4661);
xnor U5162 (N_5162,N_4996,N_4706);
xor U5163 (N_5163,N_4831,N_4578);
or U5164 (N_5164,N_4587,N_4801);
nand U5165 (N_5165,N_4736,N_4915);
xnor U5166 (N_5166,N_4564,N_4770);
nand U5167 (N_5167,N_4896,N_4949);
and U5168 (N_5168,N_4685,N_4712);
nor U5169 (N_5169,N_4532,N_4704);
nand U5170 (N_5170,N_4843,N_4882);
nor U5171 (N_5171,N_4581,N_4978);
nor U5172 (N_5172,N_4960,N_4969);
or U5173 (N_5173,N_4541,N_4727);
and U5174 (N_5174,N_4813,N_4629);
nand U5175 (N_5175,N_4713,N_4652);
nor U5176 (N_5176,N_4728,N_4966);
or U5177 (N_5177,N_4735,N_4653);
or U5178 (N_5178,N_4751,N_4936);
nand U5179 (N_5179,N_4819,N_4593);
or U5180 (N_5180,N_4874,N_4920);
or U5181 (N_5181,N_4808,N_4596);
nor U5182 (N_5182,N_4692,N_4889);
or U5183 (N_5183,N_4828,N_4557);
and U5184 (N_5184,N_4995,N_4838);
or U5185 (N_5185,N_4603,N_4612);
nand U5186 (N_5186,N_4614,N_4558);
and U5187 (N_5187,N_4732,N_4968);
and U5188 (N_5188,N_4790,N_4634);
nor U5189 (N_5189,N_4941,N_4733);
nor U5190 (N_5190,N_4755,N_4538);
nor U5191 (N_5191,N_4805,N_4656);
or U5192 (N_5192,N_4523,N_4795);
xor U5193 (N_5193,N_4984,N_4757);
xor U5194 (N_5194,N_4763,N_4938);
nand U5195 (N_5195,N_4710,N_4645);
nor U5196 (N_5196,N_4772,N_4826);
nor U5197 (N_5197,N_4738,N_4698);
nor U5198 (N_5198,N_4619,N_4595);
and U5199 (N_5199,N_4758,N_4877);
or U5200 (N_5200,N_4878,N_4618);
or U5201 (N_5201,N_4760,N_4549);
or U5202 (N_5202,N_4643,N_4909);
nand U5203 (N_5203,N_4609,N_4711);
and U5204 (N_5204,N_4928,N_4553);
or U5205 (N_5205,N_4699,N_4756);
nor U5206 (N_5206,N_4871,N_4788);
and U5207 (N_5207,N_4800,N_4550);
nand U5208 (N_5208,N_4934,N_4547);
nor U5209 (N_5209,N_4973,N_4537);
or U5210 (N_5210,N_4855,N_4937);
or U5211 (N_5211,N_4535,N_4630);
and U5212 (N_5212,N_4824,N_4573);
nor U5213 (N_5213,N_4669,N_4525);
or U5214 (N_5214,N_4576,N_4923);
xnor U5215 (N_5215,N_4804,N_4940);
and U5216 (N_5216,N_4726,N_4844);
nand U5217 (N_5217,N_4933,N_4829);
or U5218 (N_5218,N_4776,N_4950);
and U5219 (N_5219,N_4841,N_4560);
nor U5220 (N_5220,N_4767,N_4913);
and U5221 (N_5221,N_4617,N_4672);
or U5222 (N_5222,N_4551,N_4916);
nor U5223 (N_5223,N_4659,N_4745);
nand U5224 (N_5224,N_4860,N_4948);
nor U5225 (N_5225,N_4666,N_4545);
and U5226 (N_5226,N_4640,N_4526);
nor U5227 (N_5227,N_4825,N_4926);
and U5228 (N_5228,N_4610,N_4834);
and U5229 (N_5229,N_4856,N_4768);
nand U5230 (N_5230,N_4837,N_4663);
nor U5231 (N_5231,N_4518,N_4654);
and U5232 (N_5232,N_4787,N_4676);
nor U5233 (N_5233,N_4765,N_4637);
nor U5234 (N_5234,N_4914,N_4502);
nand U5235 (N_5235,N_4759,N_4911);
or U5236 (N_5236,N_4721,N_4821);
and U5237 (N_5237,N_4683,N_4893);
nand U5238 (N_5238,N_4722,N_4556);
xnor U5239 (N_5239,N_4620,N_4567);
nor U5240 (N_5240,N_4708,N_4773);
and U5241 (N_5241,N_4689,N_4737);
nor U5242 (N_5242,N_4687,N_4570);
and U5243 (N_5243,N_4833,N_4515);
nor U5244 (N_5244,N_4901,N_4796);
nor U5245 (N_5245,N_4702,N_4678);
and U5246 (N_5246,N_4512,N_4851);
nand U5247 (N_5247,N_4600,N_4516);
xnor U5248 (N_5248,N_4624,N_4693);
nand U5249 (N_5249,N_4628,N_4791);
or U5250 (N_5250,N_4759,N_4728);
or U5251 (N_5251,N_4715,N_4526);
and U5252 (N_5252,N_4673,N_4516);
or U5253 (N_5253,N_4865,N_4741);
nor U5254 (N_5254,N_4886,N_4834);
nor U5255 (N_5255,N_4827,N_4627);
nor U5256 (N_5256,N_4726,N_4761);
nand U5257 (N_5257,N_4922,N_4751);
nor U5258 (N_5258,N_4690,N_4501);
nor U5259 (N_5259,N_4942,N_4807);
and U5260 (N_5260,N_4755,N_4759);
nor U5261 (N_5261,N_4979,N_4859);
and U5262 (N_5262,N_4861,N_4519);
or U5263 (N_5263,N_4878,N_4738);
xor U5264 (N_5264,N_4573,N_4787);
nor U5265 (N_5265,N_4691,N_4760);
nor U5266 (N_5266,N_4689,N_4873);
and U5267 (N_5267,N_4594,N_4923);
nand U5268 (N_5268,N_4893,N_4529);
or U5269 (N_5269,N_4939,N_4964);
nor U5270 (N_5270,N_4670,N_4920);
nand U5271 (N_5271,N_4621,N_4591);
or U5272 (N_5272,N_4994,N_4817);
nand U5273 (N_5273,N_4994,N_4639);
xnor U5274 (N_5274,N_4894,N_4663);
or U5275 (N_5275,N_4666,N_4880);
nand U5276 (N_5276,N_4967,N_4616);
or U5277 (N_5277,N_4865,N_4997);
nor U5278 (N_5278,N_4932,N_4973);
nor U5279 (N_5279,N_4506,N_4991);
nand U5280 (N_5280,N_4975,N_4563);
nand U5281 (N_5281,N_4581,N_4520);
xnor U5282 (N_5282,N_4657,N_4641);
or U5283 (N_5283,N_4882,N_4781);
or U5284 (N_5284,N_4995,N_4974);
or U5285 (N_5285,N_4516,N_4884);
or U5286 (N_5286,N_4824,N_4732);
and U5287 (N_5287,N_4505,N_4539);
nor U5288 (N_5288,N_4548,N_4947);
or U5289 (N_5289,N_4606,N_4564);
nor U5290 (N_5290,N_4637,N_4682);
nand U5291 (N_5291,N_4791,N_4665);
or U5292 (N_5292,N_4723,N_4687);
nand U5293 (N_5293,N_4919,N_4836);
nand U5294 (N_5294,N_4761,N_4831);
xor U5295 (N_5295,N_4629,N_4883);
nand U5296 (N_5296,N_4824,N_4686);
and U5297 (N_5297,N_4924,N_4908);
and U5298 (N_5298,N_4586,N_4904);
and U5299 (N_5299,N_4707,N_4945);
or U5300 (N_5300,N_4805,N_4679);
nor U5301 (N_5301,N_4508,N_4536);
nand U5302 (N_5302,N_4665,N_4971);
and U5303 (N_5303,N_4933,N_4856);
nand U5304 (N_5304,N_4730,N_4948);
nand U5305 (N_5305,N_4721,N_4684);
or U5306 (N_5306,N_4912,N_4532);
nand U5307 (N_5307,N_4688,N_4520);
or U5308 (N_5308,N_4678,N_4933);
nor U5309 (N_5309,N_4972,N_4992);
nor U5310 (N_5310,N_4604,N_4810);
and U5311 (N_5311,N_4618,N_4922);
xnor U5312 (N_5312,N_4752,N_4779);
or U5313 (N_5313,N_4689,N_4823);
xor U5314 (N_5314,N_4751,N_4710);
or U5315 (N_5315,N_4703,N_4539);
nor U5316 (N_5316,N_4599,N_4536);
xnor U5317 (N_5317,N_4502,N_4890);
xor U5318 (N_5318,N_4890,N_4805);
nor U5319 (N_5319,N_4513,N_4686);
nor U5320 (N_5320,N_4875,N_4593);
and U5321 (N_5321,N_4793,N_4611);
and U5322 (N_5322,N_4809,N_4953);
and U5323 (N_5323,N_4726,N_4646);
or U5324 (N_5324,N_4818,N_4580);
and U5325 (N_5325,N_4565,N_4781);
nor U5326 (N_5326,N_4924,N_4946);
and U5327 (N_5327,N_4789,N_4593);
or U5328 (N_5328,N_4680,N_4640);
and U5329 (N_5329,N_4623,N_4888);
nor U5330 (N_5330,N_4610,N_4608);
nand U5331 (N_5331,N_4983,N_4612);
or U5332 (N_5332,N_4910,N_4855);
nor U5333 (N_5333,N_4705,N_4774);
or U5334 (N_5334,N_4849,N_4718);
and U5335 (N_5335,N_4726,N_4991);
and U5336 (N_5336,N_4848,N_4885);
or U5337 (N_5337,N_4814,N_4919);
and U5338 (N_5338,N_4593,N_4914);
or U5339 (N_5339,N_4517,N_4896);
nor U5340 (N_5340,N_4921,N_4938);
nand U5341 (N_5341,N_4511,N_4914);
nor U5342 (N_5342,N_4890,N_4524);
xnor U5343 (N_5343,N_4541,N_4519);
and U5344 (N_5344,N_4727,N_4921);
or U5345 (N_5345,N_4759,N_4918);
and U5346 (N_5346,N_4524,N_4753);
nand U5347 (N_5347,N_4515,N_4905);
and U5348 (N_5348,N_4740,N_4815);
and U5349 (N_5349,N_4552,N_4825);
or U5350 (N_5350,N_4674,N_4915);
nor U5351 (N_5351,N_4509,N_4866);
and U5352 (N_5352,N_4558,N_4605);
xnor U5353 (N_5353,N_4830,N_4615);
nor U5354 (N_5354,N_4629,N_4892);
nor U5355 (N_5355,N_4645,N_4972);
nor U5356 (N_5356,N_4800,N_4868);
or U5357 (N_5357,N_4871,N_4878);
nand U5358 (N_5358,N_4903,N_4776);
nor U5359 (N_5359,N_4813,N_4697);
or U5360 (N_5360,N_4641,N_4586);
or U5361 (N_5361,N_4998,N_4527);
or U5362 (N_5362,N_4935,N_4705);
nand U5363 (N_5363,N_4777,N_4667);
nand U5364 (N_5364,N_4990,N_4850);
nor U5365 (N_5365,N_4823,N_4987);
and U5366 (N_5366,N_4965,N_4878);
or U5367 (N_5367,N_4553,N_4524);
or U5368 (N_5368,N_4528,N_4783);
nor U5369 (N_5369,N_4879,N_4569);
or U5370 (N_5370,N_4741,N_4610);
xnor U5371 (N_5371,N_4844,N_4777);
nor U5372 (N_5372,N_4900,N_4713);
nand U5373 (N_5373,N_4761,N_4725);
and U5374 (N_5374,N_4858,N_4857);
nor U5375 (N_5375,N_4843,N_4664);
xnor U5376 (N_5376,N_4883,N_4828);
nand U5377 (N_5377,N_4598,N_4589);
or U5378 (N_5378,N_4739,N_4990);
and U5379 (N_5379,N_4708,N_4650);
or U5380 (N_5380,N_4765,N_4689);
and U5381 (N_5381,N_4664,N_4795);
nand U5382 (N_5382,N_4927,N_4853);
xnor U5383 (N_5383,N_4954,N_4899);
nor U5384 (N_5384,N_4790,N_4647);
and U5385 (N_5385,N_4998,N_4821);
nand U5386 (N_5386,N_4927,N_4627);
nand U5387 (N_5387,N_4907,N_4890);
and U5388 (N_5388,N_4693,N_4948);
and U5389 (N_5389,N_4868,N_4823);
nand U5390 (N_5390,N_4645,N_4980);
nand U5391 (N_5391,N_4756,N_4737);
or U5392 (N_5392,N_4545,N_4507);
or U5393 (N_5393,N_4708,N_4747);
nand U5394 (N_5394,N_4802,N_4525);
nor U5395 (N_5395,N_4788,N_4521);
nor U5396 (N_5396,N_4930,N_4829);
nor U5397 (N_5397,N_4709,N_4815);
or U5398 (N_5398,N_4664,N_4866);
and U5399 (N_5399,N_4921,N_4819);
xor U5400 (N_5400,N_4539,N_4910);
and U5401 (N_5401,N_4941,N_4559);
nor U5402 (N_5402,N_4847,N_4642);
nor U5403 (N_5403,N_4846,N_4929);
or U5404 (N_5404,N_4766,N_4964);
or U5405 (N_5405,N_4915,N_4555);
and U5406 (N_5406,N_4524,N_4697);
and U5407 (N_5407,N_4751,N_4572);
nand U5408 (N_5408,N_4781,N_4601);
xor U5409 (N_5409,N_4818,N_4816);
and U5410 (N_5410,N_4634,N_4663);
xor U5411 (N_5411,N_4578,N_4879);
and U5412 (N_5412,N_4913,N_4662);
nand U5413 (N_5413,N_4957,N_4908);
and U5414 (N_5414,N_4958,N_4514);
or U5415 (N_5415,N_4698,N_4595);
or U5416 (N_5416,N_4778,N_4741);
nand U5417 (N_5417,N_4727,N_4885);
nor U5418 (N_5418,N_4723,N_4881);
or U5419 (N_5419,N_4710,N_4842);
and U5420 (N_5420,N_4862,N_4631);
nand U5421 (N_5421,N_4500,N_4689);
or U5422 (N_5422,N_4978,N_4808);
and U5423 (N_5423,N_4593,N_4616);
nor U5424 (N_5424,N_4692,N_4588);
or U5425 (N_5425,N_4563,N_4902);
xor U5426 (N_5426,N_4984,N_4721);
or U5427 (N_5427,N_4787,N_4626);
or U5428 (N_5428,N_4591,N_4825);
nand U5429 (N_5429,N_4852,N_4707);
xor U5430 (N_5430,N_4784,N_4794);
nor U5431 (N_5431,N_4943,N_4948);
nor U5432 (N_5432,N_4723,N_4660);
xnor U5433 (N_5433,N_4626,N_4771);
and U5434 (N_5434,N_4791,N_4724);
and U5435 (N_5435,N_4565,N_4501);
nand U5436 (N_5436,N_4777,N_4651);
nand U5437 (N_5437,N_4893,N_4585);
nor U5438 (N_5438,N_4662,N_4618);
nand U5439 (N_5439,N_4641,N_4686);
nand U5440 (N_5440,N_4760,N_4622);
or U5441 (N_5441,N_4976,N_4936);
nor U5442 (N_5442,N_4801,N_4976);
nor U5443 (N_5443,N_4606,N_4568);
or U5444 (N_5444,N_4905,N_4608);
nand U5445 (N_5445,N_4961,N_4773);
nor U5446 (N_5446,N_4676,N_4805);
xnor U5447 (N_5447,N_4830,N_4807);
nand U5448 (N_5448,N_4997,N_4524);
or U5449 (N_5449,N_4919,N_4722);
nor U5450 (N_5450,N_4502,N_4696);
nor U5451 (N_5451,N_4568,N_4757);
and U5452 (N_5452,N_4945,N_4536);
and U5453 (N_5453,N_4603,N_4856);
or U5454 (N_5454,N_4878,N_4569);
nand U5455 (N_5455,N_4731,N_4896);
nand U5456 (N_5456,N_4905,N_4898);
xor U5457 (N_5457,N_4614,N_4623);
nor U5458 (N_5458,N_4530,N_4652);
nand U5459 (N_5459,N_4808,N_4606);
or U5460 (N_5460,N_4777,N_4611);
xnor U5461 (N_5461,N_4965,N_4777);
nand U5462 (N_5462,N_4710,N_4731);
or U5463 (N_5463,N_4715,N_4706);
and U5464 (N_5464,N_4833,N_4844);
nand U5465 (N_5465,N_4662,N_4877);
nor U5466 (N_5466,N_4622,N_4511);
nor U5467 (N_5467,N_4814,N_4618);
nor U5468 (N_5468,N_4951,N_4517);
or U5469 (N_5469,N_4735,N_4696);
or U5470 (N_5470,N_4787,N_4912);
nand U5471 (N_5471,N_4606,N_4639);
nor U5472 (N_5472,N_4864,N_4918);
or U5473 (N_5473,N_4830,N_4668);
and U5474 (N_5474,N_4875,N_4887);
nor U5475 (N_5475,N_4560,N_4557);
or U5476 (N_5476,N_4665,N_4557);
nor U5477 (N_5477,N_4741,N_4911);
and U5478 (N_5478,N_4562,N_4553);
or U5479 (N_5479,N_4886,N_4562);
and U5480 (N_5480,N_4725,N_4907);
nor U5481 (N_5481,N_4771,N_4963);
or U5482 (N_5482,N_4998,N_4625);
or U5483 (N_5483,N_4671,N_4630);
or U5484 (N_5484,N_4836,N_4758);
nor U5485 (N_5485,N_4555,N_4532);
or U5486 (N_5486,N_4628,N_4934);
and U5487 (N_5487,N_4545,N_4989);
and U5488 (N_5488,N_4676,N_4648);
nand U5489 (N_5489,N_4921,N_4939);
or U5490 (N_5490,N_4914,N_4763);
nand U5491 (N_5491,N_4732,N_4507);
nand U5492 (N_5492,N_4891,N_4508);
and U5493 (N_5493,N_4909,N_4696);
nand U5494 (N_5494,N_4771,N_4959);
and U5495 (N_5495,N_4718,N_4886);
nor U5496 (N_5496,N_4842,N_4528);
xor U5497 (N_5497,N_4852,N_4686);
and U5498 (N_5498,N_4730,N_4716);
xor U5499 (N_5499,N_4638,N_4903);
nand U5500 (N_5500,N_5472,N_5475);
nand U5501 (N_5501,N_5058,N_5368);
nor U5502 (N_5502,N_5414,N_5320);
nor U5503 (N_5503,N_5366,N_5232);
nand U5504 (N_5504,N_5497,N_5340);
and U5505 (N_5505,N_5195,N_5222);
nor U5506 (N_5506,N_5155,N_5403);
nor U5507 (N_5507,N_5050,N_5364);
and U5508 (N_5508,N_5003,N_5073);
or U5509 (N_5509,N_5106,N_5077);
or U5510 (N_5510,N_5397,N_5163);
or U5511 (N_5511,N_5332,N_5450);
nor U5512 (N_5512,N_5353,N_5075);
and U5513 (N_5513,N_5416,N_5474);
nand U5514 (N_5514,N_5429,N_5017);
xnor U5515 (N_5515,N_5191,N_5418);
xnor U5516 (N_5516,N_5019,N_5220);
nand U5517 (N_5517,N_5284,N_5150);
and U5518 (N_5518,N_5455,N_5380);
or U5519 (N_5519,N_5285,N_5128);
nor U5520 (N_5520,N_5273,N_5007);
nand U5521 (N_5521,N_5405,N_5358);
or U5522 (N_5522,N_5026,N_5406);
and U5523 (N_5523,N_5233,N_5076);
and U5524 (N_5524,N_5271,N_5437);
nor U5525 (N_5525,N_5262,N_5087);
nand U5526 (N_5526,N_5439,N_5415);
and U5527 (N_5527,N_5239,N_5242);
nor U5528 (N_5528,N_5375,N_5225);
or U5529 (N_5529,N_5178,N_5064);
and U5530 (N_5530,N_5072,N_5199);
or U5531 (N_5531,N_5115,N_5152);
nand U5532 (N_5532,N_5306,N_5482);
or U5533 (N_5533,N_5157,N_5465);
and U5534 (N_5534,N_5234,N_5447);
xnor U5535 (N_5535,N_5197,N_5478);
and U5536 (N_5536,N_5326,N_5452);
or U5537 (N_5537,N_5408,N_5237);
and U5538 (N_5538,N_5018,N_5432);
nand U5539 (N_5539,N_5010,N_5431);
nor U5540 (N_5540,N_5444,N_5360);
nand U5541 (N_5541,N_5292,N_5260);
xnor U5542 (N_5542,N_5316,N_5022);
nor U5543 (N_5543,N_5005,N_5013);
nand U5544 (N_5544,N_5335,N_5245);
or U5545 (N_5545,N_5243,N_5445);
and U5546 (N_5546,N_5458,N_5352);
nand U5547 (N_5547,N_5386,N_5411);
xor U5548 (N_5548,N_5173,N_5168);
nand U5549 (N_5549,N_5377,N_5094);
or U5550 (N_5550,N_5314,N_5164);
xor U5551 (N_5551,N_5264,N_5110);
and U5552 (N_5552,N_5331,N_5124);
or U5553 (N_5553,N_5361,N_5031);
nand U5554 (N_5554,N_5196,N_5088);
nor U5555 (N_5555,N_5381,N_5146);
nand U5556 (N_5556,N_5413,N_5427);
xor U5557 (N_5557,N_5188,N_5459);
nor U5558 (N_5558,N_5221,N_5460);
nor U5559 (N_5559,N_5102,N_5428);
or U5560 (N_5560,N_5471,N_5034);
or U5561 (N_5561,N_5223,N_5370);
xor U5562 (N_5562,N_5235,N_5498);
nand U5563 (N_5563,N_5261,N_5492);
nand U5564 (N_5564,N_5359,N_5154);
nor U5565 (N_5565,N_5493,N_5131);
xor U5566 (N_5566,N_5294,N_5062);
nor U5567 (N_5567,N_5097,N_5066);
and U5568 (N_5568,N_5172,N_5240);
xnor U5569 (N_5569,N_5298,N_5029);
or U5570 (N_5570,N_5118,N_5190);
and U5571 (N_5571,N_5000,N_5402);
and U5572 (N_5572,N_5184,N_5290);
nor U5573 (N_5573,N_5016,N_5295);
and U5574 (N_5574,N_5132,N_5454);
or U5575 (N_5575,N_5324,N_5399);
and U5576 (N_5576,N_5229,N_5187);
or U5577 (N_5577,N_5203,N_5486);
nand U5578 (N_5578,N_5027,N_5021);
and U5579 (N_5579,N_5484,N_5071);
and U5580 (N_5580,N_5464,N_5043);
and U5581 (N_5581,N_5384,N_5241);
xor U5582 (N_5582,N_5049,N_5138);
nand U5583 (N_5583,N_5254,N_5281);
nand U5584 (N_5584,N_5249,N_5346);
and U5585 (N_5585,N_5357,N_5434);
and U5586 (N_5586,N_5494,N_5323);
nand U5587 (N_5587,N_5193,N_5424);
xnor U5588 (N_5588,N_5453,N_5490);
nand U5589 (N_5589,N_5276,N_5165);
nand U5590 (N_5590,N_5145,N_5393);
nor U5591 (N_5591,N_5433,N_5213);
nor U5592 (N_5592,N_5476,N_5392);
nor U5593 (N_5593,N_5012,N_5309);
nor U5594 (N_5594,N_5378,N_5204);
and U5595 (N_5595,N_5348,N_5338);
and U5596 (N_5596,N_5461,N_5040);
nor U5597 (N_5597,N_5355,N_5296);
nand U5598 (N_5598,N_5160,N_5301);
and U5599 (N_5599,N_5263,N_5374);
nand U5600 (N_5600,N_5044,N_5451);
or U5601 (N_5601,N_5251,N_5480);
and U5602 (N_5602,N_5224,N_5105);
and U5603 (N_5603,N_5098,N_5079);
nand U5604 (N_5604,N_5169,N_5137);
xor U5605 (N_5605,N_5376,N_5095);
nand U5606 (N_5606,N_5311,N_5304);
nand U5607 (N_5607,N_5057,N_5247);
nor U5608 (N_5608,N_5171,N_5275);
or U5609 (N_5609,N_5238,N_5140);
nor U5610 (N_5610,N_5127,N_5347);
nand U5611 (N_5611,N_5214,N_5219);
nand U5612 (N_5612,N_5283,N_5033);
xor U5613 (N_5613,N_5250,N_5069);
nor U5614 (N_5614,N_5036,N_5356);
and U5615 (N_5615,N_5180,N_5412);
nor U5616 (N_5616,N_5114,N_5113);
nor U5617 (N_5617,N_5141,N_5181);
and U5618 (N_5618,N_5398,N_5354);
and U5619 (N_5619,N_5083,N_5487);
nand U5620 (N_5620,N_5395,N_5081);
nor U5621 (N_5621,N_5078,N_5469);
nand U5622 (N_5622,N_5253,N_5401);
or U5623 (N_5623,N_5226,N_5317);
or U5624 (N_5624,N_5328,N_5430);
or U5625 (N_5625,N_5037,N_5291);
or U5626 (N_5626,N_5068,N_5488);
or U5627 (N_5627,N_5014,N_5167);
nor U5628 (N_5628,N_5308,N_5336);
xnor U5629 (N_5629,N_5404,N_5175);
nor U5630 (N_5630,N_5371,N_5139);
xor U5631 (N_5631,N_5499,N_5126);
nand U5632 (N_5632,N_5166,N_5056);
nor U5633 (N_5633,N_5369,N_5442);
or U5634 (N_5634,N_5162,N_5206);
xor U5635 (N_5635,N_5305,N_5280);
nor U5636 (N_5636,N_5286,N_5015);
or U5637 (N_5637,N_5211,N_5119);
nor U5638 (N_5638,N_5120,N_5198);
or U5639 (N_5639,N_5192,N_5084);
or U5640 (N_5640,N_5189,N_5109);
xnor U5641 (N_5641,N_5143,N_5425);
nor U5642 (N_5642,N_5257,N_5210);
or U5643 (N_5643,N_5134,N_5074);
xnor U5644 (N_5644,N_5435,N_5020);
nor U5645 (N_5645,N_5333,N_5365);
or U5646 (N_5646,N_5045,N_5282);
nand U5647 (N_5647,N_5279,N_5256);
nor U5648 (N_5648,N_5421,N_5391);
and U5649 (N_5649,N_5121,N_5350);
or U5650 (N_5650,N_5297,N_5209);
nor U5651 (N_5651,N_5096,N_5023);
or U5652 (N_5652,N_5462,N_5339);
and U5653 (N_5653,N_5409,N_5337);
nand U5654 (N_5654,N_5055,N_5099);
xor U5655 (N_5655,N_5149,N_5407);
and U5656 (N_5656,N_5389,N_5151);
nor U5657 (N_5657,N_5438,N_5344);
nor U5658 (N_5658,N_5002,N_5117);
or U5659 (N_5659,N_5039,N_5080);
or U5660 (N_5660,N_5227,N_5363);
or U5661 (N_5661,N_5156,N_5278);
or U5662 (N_5662,N_5349,N_5258);
or U5663 (N_5663,N_5142,N_5307);
nor U5664 (N_5664,N_5367,N_5208);
or U5665 (N_5665,N_5065,N_5038);
nand U5666 (N_5666,N_5373,N_5100);
and U5667 (N_5667,N_5101,N_5293);
xor U5668 (N_5668,N_5322,N_5061);
or U5669 (N_5669,N_5082,N_5125);
nor U5670 (N_5670,N_5443,N_5047);
nor U5671 (N_5671,N_5207,N_5394);
nor U5672 (N_5672,N_5321,N_5183);
nor U5673 (N_5673,N_5417,N_5319);
xor U5674 (N_5674,N_5325,N_5379);
nor U5675 (N_5675,N_5426,N_5463);
nand U5676 (N_5676,N_5202,N_5299);
and U5677 (N_5677,N_5259,N_5313);
nand U5678 (N_5678,N_5302,N_5035);
nor U5679 (N_5679,N_5483,N_5147);
nand U5680 (N_5680,N_5179,N_5218);
or U5681 (N_5681,N_5200,N_5496);
nor U5682 (N_5682,N_5288,N_5449);
nand U5683 (N_5683,N_5315,N_5481);
nor U5684 (N_5684,N_5028,N_5266);
and U5685 (N_5685,N_5063,N_5495);
or U5686 (N_5686,N_5318,N_5060);
nor U5687 (N_5687,N_5158,N_5248);
and U5688 (N_5688,N_5334,N_5479);
nand U5689 (N_5689,N_5048,N_5252);
xor U5690 (N_5690,N_5390,N_5312);
nand U5691 (N_5691,N_5051,N_5212);
nand U5692 (N_5692,N_5089,N_5422);
and U5693 (N_5693,N_5186,N_5093);
xor U5694 (N_5694,N_5086,N_5052);
xor U5695 (N_5695,N_5255,N_5329);
nor U5696 (N_5696,N_5215,N_5032);
and U5697 (N_5697,N_5343,N_5216);
and U5698 (N_5698,N_5473,N_5001);
nor U5699 (N_5699,N_5177,N_5345);
or U5700 (N_5700,N_5091,N_5300);
or U5701 (N_5701,N_5330,N_5054);
and U5702 (N_5702,N_5383,N_5303);
nor U5703 (N_5703,N_5090,N_5059);
xnor U5704 (N_5704,N_5269,N_5092);
and U5705 (N_5705,N_5351,N_5008);
or U5706 (N_5706,N_5153,N_5042);
and U5707 (N_5707,N_5385,N_5053);
nor U5708 (N_5708,N_5174,N_5267);
nand U5709 (N_5709,N_5423,N_5228);
nand U5710 (N_5710,N_5123,N_5277);
nand U5711 (N_5711,N_5112,N_5446);
nor U5712 (N_5712,N_5470,N_5420);
nand U5713 (N_5713,N_5441,N_5268);
or U5714 (N_5714,N_5103,N_5144);
nand U5715 (N_5715,N_5310,N_5170);
or U5716 (N_5716,N_5448,N_5477);
nor U5717 (N_5717,N_5287,N_5217);
and U5718 (N_5718,N_5006,N_5108);
nand U5719 (N_5719,N_5116,N_5194);
or U5720 (N_5720,N_5436,N_5265);
xnor U5721 (N_5721,N_5382,N_5230);
nand U5722 (N_5722,N_5467,N_5396);
nand U5723 (N_5723,N_5185,N_5489);
or U5724 (N_5724,N_5067,N_5270);
nor U5725 (N_5725,N_5457,N_5104);
and U5726 (N_5726,N_5133,N_5387);
and U5727 (N_5727,N_5011,N_5372);
xnor U5728 (N_5728,N_5136,N_5466);
nor U5729 (N_5729,N_5468,N_5246);
and U5730 (N_5730,N_5456,N_5274);
nand U5731 (N_5731,N_5070,N_5205);
nand U5732 (N_5732,N_5410,N_5341);
nor U5733 (N_5733,N_5491,N_5244);
and U5734 (N_5734,N_5148,N_5231);
and U5735 (N_5735,N_5289,N_5159);
or U5736 (N_5736,N_5388,N_5342);
nand U5737 (N_5737,N_5362,N_5107);
and U5738 (N_5738,N_5135,N_5111);
and U5739 (N_5739,N_5129,N_5030);
and U5740 (N_5740,N_5236,N_5009);
and U5741 (N_5741,N_5025,N_5041);
and U5742 (N_5742,N_5122,N_5024);
nand U5743 (N_5743,N_5419,N_5046);
xnor U5744 (N_5744,N_5182,N_5004);
and U5745 (N_5745,N_5400,N_5327);
or U5746 (N_5746,N_5085,N_5176);
and U5747 (N_5747,N_5161,N_5130);
nand U5748 (N_5748,N_5485,N_5201);
and U5749 (N_5749,N_5272,N_5440);
nor U5750 (N_5750,N_5365,N_5066);
xnor U5751 (N_5751,N_5456,N_5130);
or U5752 (N_5752,N_5035,N_5474);
and U5753 (N_5753,N_5048,N_5464);
nor U5754 (N_5754,N_5235,N_5190);
or U5755 (N_5755,N_5335,N_5003);
nand U5756 (N_5756,N_5155,N_5056);
nand U5757 (N_5757,N_5049,N_5329);
and U5758 (N_5758,N_5489,N_5048);
nand U5759 (N_5759,N_5390,N_5168);
nor U5760 (N_5760,N_5214,N_5494);
or U5761 (N_5761,N_5443,N_5041);
nand U5762 (N_5762,N_5309,N_5023);
and U5763 (N_5763,N_5085,N_5064);
nor U5764 (N_5764,N_5280,N_5053);
or U5765 (N_5765,N_5045,N_5394);
xnor U5766 (N_5766,N_5076,N_5249);
xnor U5767 (N_5767,N_5057,N_5442);
xor U5768 (N_5768,N_5432,N_5020);
or U5769 (N_5769,N_5312,N_5142);
or U5770 (N_5770,N_5250,N_5432);
or U5771 (N_5771,N_5092,N_5364);
nor U5772 (N_5772,N_5362,N_5471);
nand U5773 (N_5773,N_5121,N_5476);
and U5774 (N_5774,N_5071,N_5002);
nor U5775 (N_5775,N_5427,N_5115);
nor U5776 (N_5776,N_5328,N_5335);
or U5777 (N_5777,N_5150,N_5409);
xnor U5778 (N_5778,N_5001,N_5231);
xnor U5779 (N_5779,N_5044,N_5382);
and U5780 (N_5780,N_5407,N_5470);
or U5781 (N_5781,N_5138,N_5472);
nor U5782 (N_5782,N_5046,N_5215);
or U5783 (N_5783,N_5253,N_5260);
nand U5784 (N_5784,N_5116,N_5104);
and U5785 (N_5785,N_5386,N_5259);
nand U5786 (N_5786,N_5202,N_5012);
nor U5787 (N_5787,N_5158,N_5387);
and U5788 (N_5788,N_5049,N_5039);
and U5789 (N_5789,N_5439,N_5260);
xnor U5790 (N_5790,N_5077,N_5337);
nand U5791 (N_5791,N_5049,N_5021);
and U5792 (N_5792,N_5451,N_5391);
nand U5793 (N_5793,N_5303,N_5249);
nand U5794 (N_5794,N_5066,N_5062);
and U5795 (N_5795,N_5344,N_5096);
or U5796 (N_5796,N_5485,N_5426);
or U5797 (N_5797,N_5386,N_5077);
nor U5798 (N_5798,N_5111,N_5070);
xor U5799 (N_5799,N_5095,N_5415);
nand U5800 (N_5800,N_5270,N_5321);
and U5801 (N_5801,N_5338,N_5298);
or U5802 (N_5802,N_5214,N_5450);
or U5803 (N_5803,N_5109,N_5179);
nand U5804 (N_5804,N_5273,N_5096);
nand U5805 (N_5805,N_5131,N_5031);
xor U5806 (N_5806,N_5303,N_5377);
or U5807 (N_5807,N_5424,N_5090);
xnor U5808 (N_5808,N_5470,N_5391);
xor U5809 (N_5809,N_5384,N_5324);
nand U5810 (N_5810,N_5046,N_5325);
nor U5811 (N_5811,N_5392,N_5296);
or U5812 (N_5812,N_5197,N_5023);
and U5813 (N_5813,N_5013,N_5166);
nand U5814 (N_5814,N_5069,N_5133);
and U5815 (N_5815,N_5260,N_5124);
nand U5816 (N_5816,N_5447,N_5065);
and U5817 (N_5817,N_5086,N_5194);
or U5818 (N_5818,N_5429,N_5061);
nor U5819 (N_5819,N_5270,N_5120);
nor U5820 (N_5820,N_5070,N_5377);
xnor U5821 (N_5821,N_5053,N_5006);
nand U5822 (N_5822,N_5359,N_5183);
or U5823 (N_5823,N_5347,N_5107);
xor U5824 (N_5824,N_5012,N_5354);
nor U5825 (N_5825,N_5132,N_5345);
nand U5826 (N_5826,N_5206,N_5323);
nor U5827 (N_5827,N_5272,N_5234);
nand U5828 (N_5828,N_5453,N_5319);
nor U5829 (N_5829,N_5271,N_5234);
and U5830 (N_5830,N_5257,N_5443);
or U5831 (N_5831,N_5337,N_5427);
nor U5832 (N_5832,N_5151,N_5075);
nor U5833 (N_5833,N_5355,N_5095);
nor U5834 (N_5834,N_5029,N_5113);
nand U5835 (N_5835,N_5496,N_5072);
nor U5836 (N_5836,N_5344,N_5303);
nor U5837 (N_5837,N_5254,N_5019);
or U5838 (N_5838,N_5086,N_5417);
nand U5839 (N_5839,N_5305,N_5486);
nand U5840 (N_5840,N_5252,N_5351);
nor U5841 (N_5841,N_5315,N_5177);
nand U5842 (N_5842,N_5256,N_5080);
nor U5843 (N_5843,N_5334,N_5063);
or U5844 (N_5844,N_5398,N_5303);
and U5845 (N_5845,N_5471,N_5450);
and U5846 (N_5846,N_5360,N_5018);
xor U5847 (N_5847,N_5023,N_5466);
nor U5848 (N_5848,N_5286,N_5374);
and U5849 (N_5849,N_5346,N_5386);
xnor U5850 (N_5850,N_5209,N_5245);
and U5851 (N_5851,N_5263,N_5379);
nand U5852 (N_5852,N_5046,N_5185);
nand U5853 (N_5853,N_5063,N_5431);
nor U5854 (N_5854,N_5139,N_5028);
or U5855 (N_5855,N_5271,N_5318);
or U5856 (N_5856,N_5345,N_5440);
nor U5857 (N_5857,N_5350,N_5287);
or U5858 (N_5858,N_5446,N_5433);
nor U5859 (N_5859,N_5101,N_5098);
nor U5860 (N_5860,N_5183,N_5155);
xnor U5861 (N_5861,N_5481,N_5439);
nand U5862 (N_5862,N_5092,N_5428);
and U5863 (N_5863,N_5326,N_5324);
nor U5864 (N_5864,N_5459,N_5337);
and U5865 (N_5865,N_5204,N_5477);
nand U5866 (N_5866,N_5055,N_5056);
or U5867 (N_5867,N_5298,N_5134);
nor U5868 (N_5868,N_5396,N_5220);
nor U5869 (N_5869,N_5192,N_5470);
or U5870 (N_5870,N_5190,N_5490);
nor U5871 (N_5871,N_5349,N_5000);
and U5872 (N_5872,N_5361,N_5187);
nor U5873 (N_5873,N_5029,N_5407);
nand U5874 (N_5874,N_5368,N_5339);
and U5875 (N_5875,N_5324,N_5323);
nand U5876 (N_5876,N_5108,N_5369);
nand U5877 (N_5877,N_5352,N_5249);
nand U5878 (N_5878,N_5439,N_5074);
or U5879 (N_5879,N_5154,N_5370);
and U5880 (N_5880,N_5216,N_5426);
and U5881 (N_5881,N_5097,N_5426);
nand U5882 (N_5882,N_5013,N_5124);
and U5883 (N_5883,N_5223,N_5481);
and U5884 (N_5884,N_5204,N_5240);
nand U5885 (N_5885,N_5410,N_5322);
or U5886 (N_5886,N_5016,N_5216);
xor U5887 (N_5887,N_5071,N_5180);
or U5888 (N_5888,N_5080,N_5160);
nor U5889 (N_5889,N_5038,N_5392);
nor U5890 (N_5890,N_5297,N_5446);
nand U5891 (N_5891,N_5104,N_5422);
or U5892 (N_5892,N_5352,N_5324);
and U5893 (N_5893,N_5438,N_5316);
or U5894 (N_5894,N_5255,N_5241);
or U5895 (N_5895,N_5158,N_5011);
nand U5896 (N_5896,N_5435,N_5100);
and U5897 (N_5897,N_5312,N_5454);
nor U5898 (N_5898,N_5101,N_5449);
nor U5899 (N_5899,N_5366,N_5409);
nand U5900 (N_5900,N_5330,N_5361);
nor U5901 (N_5901,N_5230,N_5496);
nor U5902 (N_5902,N_5376,N_5432);
or U5903 (N_5903,N_5255,N_5405);
xnor U5904 (N_5904,N_5498,N_5275);
or U5905 (N_5905,N_5397,N_5499);
nand U5906 (N_5906,N_5345,N_5212);
or U5907 (N_5907,N_5075,N_5222);
xnor U5908 (N_5908,N_5232,N_5105);
and U5909 (N_5909,N_5439,N_5151);
nand U5910 (N_5910,N_5313,N_5236);
and U5911 (N_5911,N_5234,N_5032);
or U5912 (N_5912,N_5443,N_5064);
or U5913 (N_5913,N_5449,N_5118);
or U5914 (N_5914,N_5122,N_5165);
nand U5915 (N_5915,N_5390,N_5295);
nor U5916 (N_5916,N_5403,N_5449);
or U5917 (N_5917,N_5213,N_5379);
or U5918 (N_5918,N_5088,N_5208);
or U5919 (N_5919,N_5185,N_5423);
nor U5920 (N_5920,N_5355,N_5031);
or U5921 (N_5921,N_5157,N_5371);
and U5922 (N_5922,N_5252,N_5284);
nor U5923 (N_5923,N_5475,N_5403);
or U5924 (N_5924,N_5237,N_5136);
nand U5925 (N_5925,N_5001,N_5198);
nor U5926 (N_5926,N_5277,N_5266);
xor U5927 (N_5927,N_5351,N_5051);
or U5928 (N_5928,N_5476,N_5280);
nand U5929 (N_5929,N_5340,N_5063);
nand U5930 (N_5930,N_5240,N_5341);
nand U5931 (N_5931,N_5280,N_5459);
and U5932 (N_5932,N_5046,N_5236);
and U5933 (N_5933,N_5398,N_5332);
or U5934 (N_5934,N_5444,N_5053);
nor U5935 (N_5935,N_5085,N_5283);
or U5936 (N_5936,N_5428,N_5123);
nor U5937 (N_5937,N_5405,N_5111);
and U5938 (N_5938,N_5256,N_5408);
or U5939 (N_5939,N_5419,N_5385);
or U5940 (N_5940,N_5232,N_5157);
or U5941 (N_5941,N_5486,N_5156);
or U5942 (N_5942,N_5296,N_5426);
xnor U5943 (N_5943,N_5374,N_5091);
and U5944 (N_5944,N_5364,N_5360);
nand U5945 (N_5945,N_5061,N_5162);
nor U5946 (N_5946,N_5015,N_5234);
and U5947 (N_5947,N_5103,N_5291);
and U5948 (N_5948,N_5414,N_5373);
and U5949 (N_5949,N_5061,N_5103);
xnor U5950 (N_5950,N_5253,N_5018);
nor U5951 (N_5951,N_5385,N_5034);
nor U5952 (N_5952,N_5105,N_5434);
xnor U5953 (N_5953,N_5197,N_5105);
nor U5954 (N_5954,N_5015,N_5103);
or U5955 (N_5955,N_5069,N_5196);
or U5956 (N_5956,N_5476,N_5414);
or U5957 (N_5957,N_5174,N_5104);
or U5958 (N_5958,N_5464,N_5017);
nand U5959 (N_5959,N_5496,N_5010);
and U5960 (N_5960,N_5103,N_5256);
or U5961 (N_5961,N_5357,N_5285);
or U5962 (N_5962,N_5452,N_5402);
or U5963 (N_5963,N_5274,N_5441);
nand U5964 (N_5964,N_5468,N_5084);
nand U5965 (N_5965,N_5069,N_5043);
nand U5966 (N_5966,N_5097,N_5460);
nor U5967 (N_5967,N_5110,N_5062);
and U5968 (N_5968,N_5109,N_5183);
and U5969 (N_5969,N_5334,N_5307);
or U5970 (N_5970,N_5479,N_5321);
and U5971 (N_5971,N_5118,N_5309);
nor U5972 (N_5972,N_5299,N_5331);
or U5973 (N_5973,N_5338,N_5114);
xnor U5974 (N_5974,N_5482,N_5329);
nor U5975 (N_5975,N_5145,N_5134);
nand U5976 (N_5976,N_5388,N_5371);
xor U5977 (N_5977,N_5443,N_5057);
or U5978 (N_5978,N_5097,N_5041);
nand U5979 (N_5979,N_5167,N_5341);
and U5980 (N_5980,N_5106,N_5018);
nor U5981 (N_5981,N_5403,N_5222);
or U5982 (N_5982,N_5340,N_5394);
and U5983 (N_5983,N_5226,N_5322);
or U5984 (N_5984,N_5032,N_5326);
and U5985 (N_5985,N_5119,N_5237);
and U5986 (N_5986,N_5493,N_5359);
xnor U5987 (N_5987,N_5474,N_5314);
nand U5988 (N_5988,N_5216,N_5349);
and U5989 (N_5989,N_5406,N_5184);
nor U5990 (N_5990,N_5450,N_5280);
and U5991 (N_5991,N_5038,N_5211);
nand U5992 (N_5992,N_5100,N_5041);
nor U5993 (N_5993,N_5208,N_5274);
and U5994 (N_5994,N_5014,N_5344);
nand U5995 (N_5995,N_5209,N_5073);
nor U5996 (N_5996,N_5430,N_5237);
nor U5997 (N_5997,N_5493,N_5281);
xnor U5998 (N_5998,N_5042,N_5040);
nand U5999 (N_5999,N_5381,N_5036);
and U6000 (N_6000,N_5808,N_5999);
nand U6001 (N_6001,N_5705,N_5821);
nand U6002 (N_6002,N_5513,N_5621);
nor U6003 (N_6003,N_5750,N_5546);
or U6004 (N_6004,N_5807,N_5971);
and U6005 (N_6005,N_5987,N_5967);
and U6006 (N_6006,N_5582,N_5690);
or U6007 (N_6007,N_5979,N_5633);
nor U6008 (N_6008,N_5682,N_5734);
or U6009 (N_6009,N_5651,N_5857);
and U6010 (N_6010,N_5673,N_5988);
and U6011 (N_6011,N_5813,N_5604);
and U6012 (N_6012,N_5518,N_5877);
and U6013 (N_6013,N_5843,N_5774);
or U6014 (N_6014,N_5667,N_5591);
nor U6015 (N_6015,N_5502,N_5576);
or U6016 (N_6016,N_5989,N_5617);
and U6017 (N_6017,N_5663,N_5635);
xnor U6018 (N_6018,N_5533,N_5672);
nor U6019 (N_6019,N_5739,N_5736);
and U6020 (N_6020,N_5931,N_5755);
and U6021 (N_6021,N_5773,N_5560);
nor U6022 (N_6022,N_5968,N_5959);
nor U6023 (N_6023,N_5930,N_5616);
nand U6024 (N_6024,N_5692,N_5731);
xnor U6025 (N_6025,N_5940,N_5783);
nor U6026 (N_6026,N_5698,N_5622);
and U6027 (N_6027,N_5539,N_5544);
nor U6028 (N_6028,N_5670,N_5565);
or U6029 (N_6029,N_5950,N_5882);
nor U6030 (N_6030,N_5613,N_5664);
or U6031 (N_6031,N_5681,N_5549);
nor U6032 (N_6032,N_5862,N_5949);
nand U6033 (N_6033,N_5679,N_5600);
or U6034 (N_6034,N_5803,N_5509);
xnor U6035 (N_6035,N_5562,N_5652);
nor U6036 (N_6036,N_5592,N_5771);
nand U6037 (N_6037,N_5687,N_5608);
or U6038 (N_6038,N_5737,N_5995);
xor U6039 (N_6039,N_5942,N_5805);
nor U6040 (N_6040,N_5876,N_5837);
or U6041 (N_6041,N_5583,N_5545);
and U6042 (N_6042,N_5970,N_5985);
or U6043 (N_6043,N_5619,N_5722);
and U6044 (N_6044,N_5607,N_5501);
or U6045 (N_6045,N_5853,N_5760);
or U6046 (N_6046,N_5951,N_5706);
or U6047 (N_6047,N_5742,N_5599);
nor U6048 (N_6048,N_5868,N_5756);
or U6049 (N_6049,N_5856,N_5637);
and U6050 (N_6050,N_5833,N_5625);
nor U6051 (N_6051,N_5535,N_5723);
nand U6052 (N_6052,N_5615,N_5516);
and U6053 (N_6053,N_5762,N_5648);
nand U6054 (N_6054,N_5830,N_5815);
or U6055 (N_6055,N_5581,N_5644);
and U6056 (N_6056,N_5566,N_5641);
xnor U6057 (N_6057,N_5902,N_5745);
and U6058 (N_6058,N_5519,N_5921);
xnor U6059 (N_6059,N_5855,N_5937);
nor U6060 (N_6060,N_5552,N_5881);
and U6061 (N_6061,N_5793,N_5838);
and U6062 (N_6062,N_5822,N_5636);
or U6063 (N_6063,N_5872,N_5772);
nand U6064 (N_6064,N_5759,N_5845);
and U6065 (N_6065,N_5677,N_5901);
nor U6066 (N_6066,N_5567,N_5721);
and U6067 (N_6067,N_5894,N_5936);
and U6068 (N_6068,N_5982,N_5955);
nor U6069 (N_6069,N_5660,N_5817);
or U6070 (N_6070,N_5764,N_5628);
or U6071 (N_6071,N_5781,N_5782);
nor U6072 (N_6072,N_5953,N_5883);
xnor U6073 (N_6073,N_5849,N_5858);
and U6074 (N_6074,N_5571,N_5656);
and U6075 (N_6075,N_5767,N_5740);
or U6076 (N_6076,N_5933,N_5957);
nand U6077 (N_6077,N_5761,N_5630);
and U6078 (N_6078,N_5585,N_5890);
xor U6079 (N_6079,N_5507,N_5963);
or U6080 (N_6080,N_5810,N_5792);
nand U6081 (N_6081,N_5956,N_5898);
nor U6082 (N_6082,N_5666,N_5896);
nor U6083 (N_6083,N_5913,N_5958);
or U6084 (N_6084,N_5802,N_5671);
or U6085 (N_6085,N_5683,N_5563);
or U6086 (N_6086,N_5965,N_5952);
nor U6087 (N_6087,N_5598,N_5820);
or U6088 (N_6088,N_5747,N_5720);
nand U6089 (N_6089,N_5925,N_5758);
nor U6090 (N_6090,N_5974,N_5643);
or U6091 (N_6091,N_5661,N_5986);
nor U6092 (N_6092,N_5540,N_5553);
nand U6093 (N_6093,N_5897,N_5611);
nand U6094 (N_6094,N_5915,N_5559);
nand U6095 (N_6095,N_5551,N_5529);
xor U6096 (N_6096,N_5645,N_5927);
nor U6097 (N_6097,N_5912,N_5728);
or U6098 (N_6098,N_5919,N_5850);
nand U6099 (N_6099,N_5627,N_5505);
xor U6100 (N_6100,N_5983,N_5675);
nor U6101 (N_6101,N_5578,N_5939);
or U6102 (N_6102,N_5725,N_5954);
xnor U6103 (N_6103,N_5842,N_5642);
and U6104 (N_6104,N_5841,N_5867);
or U6105 (N_6105,N_5909,N_5934);
and U6106 (N_6106,N_5520,N_5729);
or U6107 (N_6107,N_5639,N_5554);
nand U6108 (N_6108,N_5929,N_5558);
nand U6109 (N_6109,N_5547,N_5763);
nor U6110 (N_6110,N_5832,N_5870);
or U6111 (N_6111,N_5586,N_5695);
or U6112 (N_6112,N_5693,N_5840);
and U6113 (N_6113,N_5848,N_5914);
nand U6114 (N_6114,N_5573,N_5926);
or U6115 (N_6115,N_5790,N_5548);
and U6116 (N_6116,N_5946,N_5984);
or U6117 (N_6117,N_5990,N_5691);
nand U6118 (N_6118,N_5504,N_5597);
or U6119 (N_6119,N_5806,N_5515);
and U6120 (N_6120,N_5694,N_5708);
or U6121 (N_6121,N_5688,N_5647);
or U6122 (N_6122,N_5538,N_5800);
xnor U6123 (N_6123,N_5665,N_5605);
nand U6124 (N_6124,N_5887,N_5714);
nor U6125 (N_6125,N_5542,N_5825);
nor U6126 (N_6126,N_5685,N_5657);
nor U6127 (N_6127,N_5579,N_5993);
nor U6128 (N_6128,N_5875,N_5517);
nand U6129 (N_6129,N_5861,N_5738);
xor U6130 (N_6130,N_5669,N_5701);
nand U6131 (N_6131,N_5620,N_5892);
and U6132 (N_6132,N_5814,N_5733);
nand U6133 (N_6133,N_5534,N_5580);
or U6134 (N_6134,N_5584,N_5572);
xnor U6135 (N_6135,N_5922,N_5906);
or U6136 (N_6136,N_5844,N_5903);
and U6137 (N_6137,N_5713,N_5824);
nand U6138 (N_6138,N_5588,N_5543);
nor U6139 (N_6139,N_5812,N_5526);
nand U6140 (N_6140,N_5878,N_5527);
nand U6141 (N_6141,N_5511,N_5703);
and U6142 (N_6142,N_5594,N_5503);
nor U6143 (N_6143,N_5741,N_5618);
nand U6144 (N_6144,N_5658,N_5795);
or U6145 (N_6145,N_5880,N_5819);
nand U6146 (N_6146,N_5589,N_5997);
or U6147 (N_6147,N_5938,N_5977);
or U6148 (N_6148,N_5972,N_5743);
or U6149 (N_6149,N_5521,N_5964);
nor U6150 (N_6150,N_5874,N_5827);
nor U6151 (N_6151,N_5754,N_5650);
xnor U6152 (N_6152,N_5863,N_5851);
nor U6153 (N_6153,N_5776,N_5525);
or U6154 (N_6154,N_5780,N_5717);
nand U6155 (N_6155,N_5587,N_5707);
nand U6156 (N_6156,N_5944,N_5962);
nor U6157 (N_6157,N_5697,N_5826);
nor U6158 (N_6158,N_5899,N_5568);
nor U6159 (N_6159,N_5943,N_5500);
nor U6160 (N_6160,N_5798,N_5744);
xnor U6161 (N_6161,N_5770,N_5866);
and U6162 (N_6162,N_5710,N_5555);
nor U6163 (N_6163,N_5537,N_5557);
nand U6164 (N_6164,N_5991,N_5948);
xnor U6165 (N_6165,N_5603,N_5917);
nor U6166 (N_6166,N_5654,N_5907);
or U6167 (N_6167,N_5606,N_5590);
nand U6168 (N_6168,N_5779,N_5976);
or U6169 (N_6169,N_5765,N_5649);
and U6170 (N_6170,N_5961,N_5757);
or U6171 (N_6171,N_5610,N_5879);
or U6172 (N_6172,N_5998,N_5904);
nor U6173 (N_6173,N_5602,N_5836);
nor U6174 (N_6174,N_5532,N_5689);
nand U6175 (N_6175,N_5596,N_5715);
nand U6176 (N_6176,N_5847,N_5854);
and U6177 (N_6177,N_5769,N_5924);
or U6178 (N_6178,N_5994,N_5823);
xor U6179 (N_6179,N_5601,N_5746);
nor U6180 (N_6180,N_5920,N_5624);
nor U6181 (N_6181,N_5561,N_5818);
nand U6182 (N_6182,N_5512,N_5704);
nand U6183 (N_6183,N_5778,N_5900);
nor U6184 (N_6184,N_5911,N_5905);
nand U6185 (N_6185,N_5684,N_5574);
nor U6186 (N_6186,N_5891,N_5659);
and U6187 (N_6187,N_5831,N_5724);
or U6188 (N_6188,N_5678,N_5766);
or U6189 (N_6189,N_5653,N_5941);
xor U6190 (N_6190,N_5730,N_5629);
nand U6191 (N_6191,N_5751,N_5680);
and U6192 (N_6192,N_5631,N_5788);
and U6193 (N_6193,N_5749,N_5752);
nand U6194 (N_6194,N_5873,N_5676);
and U6195 (N_6195,N_5871,N_5797);
nor U6196 (N_6196,N_5804,N_5910);
nand U6197 (N_6197,N_5794,N_5791);
and U6198 (N_6198,N_5799,N_5556);
nand U6199 (N_6199,N_5865,N_5975);
or U6200 (N_6200,N_5784,N_5992);
and U6201 (N_6201,N_5726,N_5510);
nor U6202 (N_6202,N_5945,N_5889);
xnor U6203 (N_6203,N_5508,N_5716);
or U6204 (N_6204,N_5973,N_5932);
or U6205 (N_6205,N_5835,N_5609);
nor U6206 (N_6206,N_5524,N_5978);
or U6207 (N_6207,N_5550,N_5514);
or U6208 (N_6208,N_5996,N_5718);
and U6209 (N_6209,N_5506,N_5593);
and U6210 (N_6210,N_5869,N_5839);
nor U6211 (N_6211,N_5777,N_5864);
or U6212 (N_6212,N_5719,N_5531);
nand U6213 (N_6213,N_5564,N_5785);
and U6214 (N_6214,N_5702,N_5859);
xor U6215 (N_6215,N_5960,N_5709);
xnor U6216 (N_6216,N_5918,N_5885);
or U6217 (N_6217,N_5753,N_5536);
nor U6218 (N_6218,N_5860,N_5846);
nor U6219 (N_6219,N_5748,N_5700);
xor U6220 (N_6220,N_5966,N_5522);
nor U6221 (N_6221,N_5969,N_5528);
or U6222 (N_6222,N_5595,N_5735);
xor U6223 (N_6223,N_5634,N_5569);
nand U6224 (N_6224,N_5732,N_5614);
and U6225 (N_6225,N_5884,N_5928);
xor U6226 (N_6226,N_5523,N_5852);
or U6227 (N_6227,N_5638,N_5801);
and U6228 (N_6228,N_5727,N_5796);
or U6229 (N_6229,N_5893,N_5668);
and U6230 (N_6230,N_5686,N_5816);
nor U6231 (N_6231,N_5768,N_5655);
nand U6232 (N_6232,N_5786,N_5570);
and U6233 (N_6233,N_5646,N_5612);
nor U6234 (N_6234,N_5809,N_5711);
or U6235 (N_6235,N_5923,N_5834);
nand U6236 (N_6236,N_5640,N_5530);
or U6237 (N_6237,N_5626,N_5696);
or U6238 (N_6238,N_5886,N_5888);
nor U6239 (N_6239,N_5811,N_5775);
or U6240 (N_6240,N_5623,N_5980);
and U6241 (N_6241,N_5828,N_5674);
nand U6242 (N_6242,N_5895,N_5829);
or U6243 (N_6243,N_5699,N_5712);
nand U6244 (N_6244,N_5662,N_5935);
nand U6245 (N_6245,N_5632,N_5575);
nor U6246 (N_6246,N_5908,N_5981);
nand U6247 (N_6247,N_5577,N_5787);
nor U6248 (N_6248,N_5916,N_5789);
or U6249 (N_6249,N_5541,N_5947);
nor U6250 (N_6250,N_5740,N_5671);
or U6251 (N_6251,N_5975,N_5968);
nor U6252 (N_6252,N_5567,N_5752);
nand U6253 (N_6253,N_5810,N_5616);
and U6254 (N_6254,N_5930,N_5950);
nor U6255 (N_6255,N_5918,N_5645);
and U6256 (N_6256,N_5945,N_5591);
nand U6257 (N_6257,N_5881,N_5983);
nor U6258 (N_6258,N_5855,N_5716);
nand U6259 (N_6259,N_5646,N_5954);
nand U6260 (N_6260,N_5714,N_5593);
nand U6261 (N_6261,N_5614,N_5747);
or U6262 (N_6262,N_5771,N_5929);
or U6263 (N_6263,N_5567,N_5783);
nor U6264 (N_6264,N_5759,N_5874);
nor U6265 (N_6265,N_5703,N_5685);
xor U6266 (N_6266,N_5960,N_5607);
and U6267 (N_6267,N_5526,N_5732);
and U6268 (N_6268,N_5505,N_5935);
xor U6269 (N_6269,N_5980,N_5868);
and U6270 (N_6270,N_5791,N_5767);
nand U6271 (N_6271,N_5853,N_5641);
and U6272 (N_6272,N_5867,N_5771);
nor U6273 (N_6273,N_5887,N_5772);
or U6274 (N_6274,N_5627,N_5789);
nand U6275 (N_6275,N_5690,N_5532);
nand U6276 (N_6276,N_5980,N_5688);
nand U6277 (N_6277,N_5883,N_5573);
and U6278 (N_6278,N_5896,N_5836);
nor U6279 (N_6279,N_5900,N_5893);
and U6280 (N_6280,N_5993,N_5978);
xor U6281 (N_6281,N_5673,N_5938);
nand U6282 (N_6282,N_5780,N_5629);
nand U6283 (N_6283,N_5589,N_5763);
nor U6284 (N_6284,N_5609,N_5526);
nor U6285 (N_6285,N_5778,N_5950);
xnor U6286 (N_6286,N_5952,N_5792);
nand U6287 (N_6287,N_5872,N_5760);
and U6288 (N_6288,N_5966,N_5708);
or U6289 (N_6289,N_5552,N_5777);
or U6290 (N_6290,N_5591,N_5704);
nand U6291 (N_6291,N_5591,N_5734);
nor U6292 (N_6292,N_5728,N_5622);
or U6293 (N_6293,N_5730,N_5755);
nor U6294 (N_6294,N_5601,N_5559);
nor U6295 (N_6295,N_5530,N_5825);
and U6296 (N_6296,N_5742,N_5603);
nand U6297 (N_6297,N_5698,N_5798);
and U6298 (N_6298,N_5556,N_5887);
nand U6299 (N_6299,N_5991,N_5698);
xor U6300 (N_6300,N_5675,N_5658);
nor U6301 (N_6301,N_5854,N_5588);
nor U6302 (N_6302,N_5868,N_5617);
and U6303 (N_6303,N_5663,N_5918);
nor U6304 (N_6304,N_5630,N_5508);
nand U6305 (N_6305,N_5716,N_5923);
xnor U6306 (N_6306,N_5743,N_5577);
nand U6307 (N_6307,N_5520,N_5693);
and U6308 (N_6308,N_5990,N_5887);
and U6309 (N_6309,N_5812,N_5527);
and U6310 (N_6310,N_5773,N_5550);
xnor U6311 (N_6311,N_5850,N_5555);
or U6312 (N_6312,N_5706,N_5641);
nand U6313 (N_6313,N_5508,N_5686);
nand U6314 (N_6314,N_5880,N_5556);
nor U6315 (N_6315,N_5737,N_5780);
nand U6316 (N_6316,N_5973,N_5553);
nor U6317 (N_6317,N_5529,N_5591);
or U6318 (N_6318,N_5941,N_5671);
nand U6319 (N_6319,N_5815,N_5823);
or U6320 (N_6320,N_5748,N_5828);
and U6321 (N_6321,N_5673,N_5939);
nor U6322 (N_6322,N_5987,N_5584);
nand U6323 (N_6323,N_5944,N_5995);
nor U6324 (N_6324,N_5585,N_5552);
and U6325 (N_6325,N_5953,N_5877);
nand U6326 (N_6326,N_5681,N_5908);
nand U6327 (N_6327,N_5896,N_5615);
nor U6328 (N_6328,N_5616,N_5893);
and U6329 (N_6329,N_5619,N_5853);
nand U6330 (N_6330,N_5731,N_5881);
or U6331 (N_6331,N_5832,N_5702);
or U6332 (N_6332,N_5989,N_5930);
or U6333 (N_6333,N_5888,N_5671);
or U6334 (N_6334,N_5545,N_5525);
nor U6335 (N_6335,N_5655,N_5656);
nand U6336 (N_6336,N_5710,N_5671);
and U6337 (N_6337,N_5605,N_5950);
or U6338 (N_6338,N_5513,N_5758);
or U6339 (N_6339,N_5794,N_5637);
nor U6340 (N_6340,N_5963,N_5577);
nor U6341 (N_6341,N_5882,N_5908);
or U6342 (N_6342,N_5655,N_5689);
xnor U6343 (N_6343,N_5633,N_5525);
and U6344 (N_6344,N_5976,N_5700);
or U6345 (N_6345,N_5775,N_5723);
xnor U6346 (N_6346,N_5596,N_5541);
xor U6347 (N_6347,N_5534,N_5860);
nand U6348 (N_6348,N_5821,N_5599);
nand U6349 (N_6349,N_5865,N_5951);
nand U6350 (N_6350,N_5944,N_5989);
nor U6351 (N_6351,N_5742,N_5546);
or U6352 (N_6352,N_5915,N_5573);
nand U6353 (N_6353,N_5663,N_5831);
and U6354 (N_6354,N_5974,N_5565);
and U6355 (N_6355,N_5828,N_5886);
and U6356 (N_6356,N_5935,N_5627);
or U6357 (N_6357,N_5787,N_5605);
nor U6358 (N_6358,N_5962,N_5919);
nor U6359 (N_6359,N_5896,N_5647);
and U6360 (N_6360,N_5733,N_5666);
nand U6361 (N_6361,N_5926,N_5817);
xor U6362 (N_6362,N_5821,N_5596);
or U6363 (N_6363,N_5846,N_5896);
nand U6364 (N_6364,N_5723,N_5740);
nor U6365 (N_6365,N_5618,N_5955);
nor U6366 (N_6366,N_5736,N_5694);
and U6367 (N_6367,N_5545,N_5674);
or U6368 (N_6368,N_5954,N_5712);
or U6369 (N_6369,N_5865,N_5609);
or U6370 (N_6370,N_5990,N_5853);
nor U6371 (N_6371,N_5515,N_5504);
and U6372 (N_6372,N_5669,N_5826);
and U6373 (N_6373,N_5551,N_5631);
and U6374 (N_6374,N_5636,N_5643);
and U6375 (N_6375,N_5519,N_5860);
or U6376 (N_6376,N_5656,N_5809);
nor U6377 (N_6377,N_5758,N_5670);
nor U6378 (N_6378,N_5912,N_5733);
nand U6379 (N_6379,N_5848,N_5625);
nand U6380 (N_6380,N_5980,N_5927);
and U6381 (N_6381,N_5700,N_5945);
nand U6382 (N_6382,N_5608,N_5544);
xnor U6383 (N_6383,N_5986,N_5911);
or U6384 (N_6384,N_5605,N_5771);
or U6385 (N_6385,N_5846,N_5622);
nand U6386 (N_6386,N_5831,N_5684);
nand U6387 (N_6387,N_5658,N_5602);
xor U6388 (N_6388,N_5512,N_5513);
or U6389 (N_6389,N_5511,N_5715);
nand U6390 (N_6390,N_5683,N_5997);
nand U6391 (N_6391,N_5673,N_5992);
or U6392 (N_6392,N_5725,N_5976);
nor U6393 (N_6393,N_5741,N_5519);
nor U6394 (N_6394,N_5900,N_5968);
and U6395 (N_6395,N_5969,N_5877);
xnor U6396 (N_6396,N_5597,N_5658);
nor U6397 (N_6397,N_5512,N_5881);
nand U6398 (N_6398,N_5844,N_5742);
or U6399 (N_6399,N_5695,N_5739);
nor U6400 (N_6400,N_5993,N_5518);
or U6401 (N_6401,N_5831,N_5823);
and U6402 (N_6402,N_5669,N_5534);
nand U6403 (N_6403,N_5594,N_5570);
or U6404 (N_6404,N_5916,N_5800);
nand U6405 (N_6405,N_5746,N_5926);
nor U6406 (N_6406,N_5633,N_5950);
and U6407 (N_6407,N_5877,N_5699);
nor U6408 (N_6408,N_5607,N_5692);
xor U6409 (N_6409,N_5905,N_5720);
or U6410 (N_6410,N_5636,N_5674);
and U6411 (N_6411,N_5997,N_5611);
nand U6412 (N_6412,N_5956,N_5957);
nor U6413 (N_6413,N_5892,N_5549);
nand U6414 (N_6414,N_5942,N_5633);
and U6415 (N_6415,N_5537,N_5894);
or U6416 (N_6416,N_5860,N_5961);
nand U6417 (N_6417,N_5632,N_5858);
and U6418 (N_6418,N_5970,N_5965);
and U6419 (N_6419,N_5764,N_5648);
xor U6420 (N_6420,N_5709,N_5874);
and U6421 (N_6421,N_5615,N_5716);
xnor U6422 (N_6422,N_5918,N_5771);
nand U6423 (N_6423,N_5624,N_5531);
nor U6424 (N_6424,N_5854,N_5583);
nand U6425 (N_6425,N_5769,N_5678);
and U6426 (N_6426,N_5698,N_5880);
or U6427 (N_6427,N_5536,N_5784);
and U6428 (N_6428,N_5878,N_5660);
nand U6429 (N_6429,N_5720,N_5746);
or U6430 (N_6430,N_5874,N_5909);
and U6431 (N_6431,N_5697,N_5807);
nor U6432 (N_6432,N_5836,N_5649);
or U6433 (N_6433,N_5872,N_5892);
nor U6434 (N_6434,N_5968,N_5830);
nand U6435 (N_6435,N_5661,N_5647);
and U6436 (N_6436,N_5925,N_5838);
or U6437 (N_6437,N_5796,N_5554);
and U6438 (N_6438,N_5676,N_5888);
or U6439 (N_6439,N_5676,N_5705);
nand U6440 (N_6440,N_5669,N_5608);
xor U6441 (N_6441,N_5911,N_5666);
nand U6442 (N_6442,N_5708,N_5552);
nand U6443 (N_6443,N_5714,N_5706);
nand U6444 (N_6444,N_5836,N_5564);
nand U6445 (N_6445,N_5761,N_5816);
nand U6446 (N_6446,N_5905,N_5535);
xor U6447 (N_6447,N_5839,N_5964);
nand U6448 (N_6448,N_5898,N_5934);
or U6449 (N_6449,N_5613,N_5784);
and U6450 (N_6450,N_5820,N_5866);
or U6451 (N_6451,N_5683,N_5835);
or U6452 (N_6452,N_5946,N_5838);
nor U6453 (N_6453,N_5544,N_5954);
xnor U6454 (N_6454,N_5616,N_5613);
nor U6455 (N_6455,N_5931,N_5593);
xor U6456 (N_6456,N_5694,N_5921);
nand U6457 (N_6457,N_5679,N_5990);
or U6458 (N_6458,N_5543,N_5660);
nor U6459 (N_6459,N_5927,N_5668);
and U6460 (N_6460,N_5725,N_5681);
nand U6461 (N_6461,N_5843,N_5577);
nor U6462 (N_6462,N_5875,N_5623);
nor U6463 (N_6463,N_5988,N_5909);
nand U6464 (N_6464,N_5926,N_5921);
and U6465 (N_6465,N_5896,N_5875);
or U6466 (N_6466,N_5871,N_5939);
nor U6467 (N_6467,N_5939,N_5532);
or U6468 (N_6468,N_5805,N_5856);
or U6469 (N_6469,N_5547,N_5883);
or U6470 (N_6470,N_5663,N_5751);
and U6471 (N_6471,N_5596,N_5696);
nor U6472 (N_6472,N_5537,N_5858);
nand U6473 (N_6473,N_5876,N_5619);
or U6474 (N_6474,N_5672,N_5800);
and U6475 (N_6475,N_5661,N_5750);
or U6476 (N_6476,N_5605,N_5782);
nor U6477 (N_6477,N_5529,N_5516);
nand U6478 (N_6478,N_5766,N_5660);
nor U6479 (N_6479,N_5539,N_5990);
or U6480 (N_6480,N_5555,N_5972);
nand U6481 (N_6481,N_5613,N_5982);
and U6482 (N_6482,N_5518,N_5535);
or U6483 (N_6483,N_5804,N_5814);
nor U6484 (N_6484,N_5808,N_5668);
nor U6485 (N_6485,N_5525,N_5559);
nor U6486 (N_6486,N_5607,N_5708);
nor U6487 (N_6487,N_5880,N_5820);
xor U6488 (N_6488,N_5559,N_5941);
nor U6489 (N_6489,N_5851,N_5535);
nor U6490 (N_6490,N_5593,N_5939);
and U6491 (N_6491,N_5963,N_5502);
nand U6492 (N_6492,N_5926,N_5807);
and U6493 (N_6493,N_5831,N_5872);
and U6494 (N_6494,N_5642,N_5954);
or U6495 (N_6495,N_5536,N_5967);
and U6496 (N_6496,N_5962,N_5730);
nor U6497 (N_6497,N_5923,N_5512);
or U6498 (N_6498,N_5929,N_5786);
nand U6499 (N_6499,N_5641,N_5547);
and U6500 (N_6500,N_6089,N_6412);
nand U6501 (N_6501,N_6326,N_6069);
nand U6502 (N_6502,N_6358,N_6373);
nand U6503 (N_6503,N_6313,N_6120);
nand U6504 (N_6504,N_6483,N_6433);
nor U6505 (N_6505,N_6060,N_6333);
and U6506 (N_6506,N_6251,N_6476);
or U6507 (N_6507,N_6307,N_6245);
nor U6508 (N_6508,N_6265,N_6299);
xor U6509 (N_6509,N_6078,N_6487);
or U6510 (N_6510,N_6444,N_6212);
nor U6511 (N_6511,N_6281,N_6362);
nand U6512 (N_6512,N_6050,N_6453);
xnor U6513 (N_6513,N_6230,N_6149);
or U6514 (N_6514,N_6314,N_6370);
nand U6515 (N_6515,N_6104,N_6392);
and U6516 (N_6516,N_6341,N_6106);
and U6517 (N_6517,N_6327,N_6010);
or U6518 (N_6518,N_6303,N_6300);
nand U6519 (N_6519,N_6154,N_6441);
or U6520 (N_6520,N_6322,N_6289);
and U6521 (N_6521,N_6335,N_6079);
nor U6522 (N_6522,N_6234,N_6467);
or U6523 (N_6523,N_6012,N_6336);
and U6524 (N_6524,N_6290,N_6052);
xnor U6525 (N_6525,N_6001,N_6499);
nand U6526 (N_6526,N_6080,N_6142);
or U6527 (N_6527,N_6416,N_6144);
or U6528 (N_6528,N_6217,N_6235);
or U6529 (N_6529,N_6241,N_6123);
nor U6530 (N_6530,N_6065,N_6419);
and U6531 (N_6531,N_6237,N_6082);
or U6532 (N_6532,N_6143,N_6007);
nand U6533 (N_6533,N_6338,N_6255);
nor U6534 (N_6534,N_6365,N_6054);
nor U6535 (N_6535,N_6343,N_6190);
and U6536 (N_6536,N_6029,N_6394);
nand U6537 (N_6537,N_6015,N_6229);
and U6538 (N_6538,N_6100,N_6397);
nor U6539 (N_6539,N_6191,N_6296);
xnor U6540 (N_6540,N_6278,N_6231);
xnor U6541 (N_6541,N_6486,N_6068);
or U6542 (N_6542,N_6178,N_6044);
nand U6543 (N_6543,N_6196,N_6471);
nand U6544 (N_6544,N_6179,N_6051);
and U6545 (N_6545,N_6099,N_6447);
and U6546 (N_6546,N_6406,N_6248);
or U6547 (N_6547,N_6260,N_6200);
nor U6548 (N_6548,N_6334,N_6389);
or U6549 (N_6549,N_6088,N_6353);
or U6550 (N_6550,N_6308,N_6094);
xnor U6551 (N_6551,N_6396,N_6359);
nor U6552 (N_6552,N_6455,N_6016);
nor U6553 (N_6553,N_6460,N_6113);
xor U6554 (N_6554,N_6214,N_6366);
and U6555 (N_6555,N_6085,N_6436);
nor U6556 (N_6556,N_6139,N_6270);
or U6557 (N_6557,N_6118,N_6133);
and U6558 (N_6558,N_6495,N_6115);
or U6559 (N_6559,N_6328,N_6355);
or U6560 (N_6560,N_6207,N_6163);
nor U6561 (N_6561,N_6030,N_6036);
nand U6562 (N_6562,N_6378,N_6288);
nand U6563 (N_6563,N_6349,N_6272);
nand U6564 (N_6564,N_6449,N_6150);
nor U6565 (N_6565,N_6042,N_6407);
nand U6566 (N_6566,N_6472,N_6456);
xor U6567 (N_6567,N_6188,N_6309);
nor U6568 (N_6568,N_6236,N_6384);
or U6569 (N_6569,N_6166,N_6284);
or U6570 (N_6570,N_6292,N_6021);
nand U6571 (N_6571,N_6473,N_6103);
nand U6572 (N_6572,N_6004,N_6385);
xor U6573 (N_6573,N_6264,N_6201);
and U6574 (N_6574,N_6438,N_6072);
nand U6575 (N_6575,N_6430,N_6092);
or U6576 (N_6576,N_6147,N_6423);
and U6577 (N_6577,N_6193,N_6452);
nor U6578 (N_6578,N_6208,N_6310);
nand U6579 (N_6579,N_6404,N_6494);
or U6580 (N_6580,N_6274,N_6268);
nand U6581 (N_6581,N_6491,N_6262);
and U6582 (N_6582,N_6427,N_6114);
and U6583 (N_6583,N_6039,N_6332);
and U6584 (N_6584,N_6254,N_6368);
and U6585 (N_6585,N_6492,N_6405);
and U6586 (N_6586,N_6445,N_6111);
or U6587 (N_6587,N_6238,N_6169);
nand U6588 (N_6588,N_6038,N_6195);
xor U6589 (N_6589,N_6291,N_6376);
and U6590 (N_6590,N_6175,N_6095);
or U6591 (N_6591,N_6083,N_6435);
nand U6592 (N_6592,N_6182,N_6371);
and U6593 (N_6593,N_6093,N_6171);
nor U6594 (N_6594,N_6097,N_6330);
nor U6595 (N_6595,N_6233,N_6253);
nand U6596 (N_6596,N_6402,N_6351);
nand U6597 (N_6597,N_6361,N_6439);
xnor U6598 (N_6598,N_6216,N_6219);
nor U6599 (N_6599,N_6321,N_6357);
nand U6600 (N_6600,N_6170,N_6064);
nor U6601 (N_6601,N_6090,N_6342);
and U6602 (N_6602,N_6383,N_6024);
nor U6603 (N_6603,N_6498,N_6167);
and U6604 (N_6604,N_6372,N_6160);
nor U6605 (N_6605,N_6110,N_6222);
nand U6606 (N_6606,N_6468,N_6059);
nor U6607 (N_6607,N_6391,N_6298);
and U6608 (N_6608,N_6409,N_6184);
or U6609 (N_6609,N_6223,N_6386);
xor U6610 (N_6610,N_6275,N_6345);
and U6611 (N_6611,N_6461,N_6221);
nor U6612 (N_6612,N_6379,N_6388);
or U6613 (N_6613,N_6459,N_6367);
or U6614 (N_6614,N_6426,N_6061);
nand U6615 (N_6615,N_6194,N_6390);
nand U6616 (N_6616,N_6172,N_6352);
nand U6617 (N_6617,N_6399,N_6232);
nor U6618 (N_6618,N_6045,N_6017);
and U6619 (N_6619,N_6450,N_6022);
nand U6620 (N_6620,N_6152,N_6263);
nor U6621 (N_6621,N_6457,N_6320);
nor U6622 (N_6622,N_6470,N_6210);
xor U6623 (N_6623,N_6496,N_6180);
or U6624 (N_6624,N_6032,N_6130);
xor U6625 (N_6625,N_6224,N_6108);
xnor U6626 (N_6626,N_6129,N_6070);
nor U6627 (N_6627,N_6434,N_6458);
nor U6628 (N_6628,N_6031,N_6442);
nand U6629 (N_6629,N_6462,N_6325);
nand U6630 (N_6630,N_6316,N_6252);
and U6631 (N_6631,N_6364,N_6206);
and U6632 (N_6632,N_6013,N_6285);
xnor U6633 (N_6633,N_6134,N_6006);
xnor U6634 (N_6634,N_6280,N_6008);
nor U6635 (N_6635,N_6127,N_6005);
xnor U6636 (N_6636,N_6279,N_6023);
or U6637 (N_6637,N_6109,N_6122);
nand U6638 (N_6638,N_6153,N_6432);
xnor U6639 (N_6639,N_6211,N_6318);
nand U6640 (N_6640,N_6091,N_6148);
or U6641 (N_6641,N_6227,N_6053);
and U6642 (N_6642,N_6293,N_6347);
and U6643 (N_6643,N_6000,N_6018);
nor U6644 (N_6644,N_6225,N_6173);
xnor U6645 (N_6645,N_6497,N_6198);
xor U6646 (N_6646,N_6176,N_6489);
and U6647 (N_6647,N_6158,N_6155);
or U6648 (N_6648,N_6297,N_6112);
or U6649 (N_6649,N_6375,N_6204);
and U6650 (N_6650,N_6057,N_6181);
nor U6651 (N_6651,N_6157,N_6084);
and U6652 (N_6652,N_6116,N_6425);
and U6653 (N_6653,N_6363,N_6411);
nor U6654 (N_6654,N_6466,N_6062);
or U6655 (N_6655,N_6259,N_6002);
xor U6656 (N_6656,N_6218,N_6382);
and U6657 (N_6657,N_6026,N_6209);
nor U6658 (N_6658,N_6037,N_6480);
or U6659 (N_6659,N_6081,N_6076);
nor U6660 (N_6660,N_6192,N_6164);
and U6661 (N_6661,N_6096,N_6340);
nand U6662 (N_6662,N_6043,N_6315);
nand U6663 (N_6663,N_6271,N_6454);
xnor U6664 (N_6664,N_6146,N_6429);
and U6665 (N_6665,N_6183,N_6474);
and U6666 (N_6666,N_6101,N_6475);
nor U6667 (N_6667,N_6478,N_6185);
and U6668 (N_6668,N_6395,N_6187);
nor U6669 (N_6669,N_6269,N_6344);
nand U6670 (N_6670,N_6469,N_6028);
nor U6671 (N_6671,N_6258,N_6014);
nor U6672 (N_6672,N_6276,N_6408);
nor U6673 (N_6673,N_6186,N_6145);
nor U6674 (N_6674,N_6086,N_6161);
or U6675 (N_6675,N_6121,N_6011);
and U6676 (N_6676,N_6294,N_6034);
nor U6677 (N_6677,N_6422,N_6354);
or U6678 (N_6678,N_6490,N_6136);
nand U6679 (N_6679,N_6302,N_6381);
nand U6680 (N_6680,N_6446,N_6305);
xnor U6681 (N_6681,N_6283,N_6448);
nor U6682 (N_6682,N_6067,N_6400);
xor U6683 (N_6683,N_6226,N_6055);
or U6684 (N_6684,N_6420,N_6047);
and U6685 (N_6685,N_6119,N_6304);
and U6686 (N_6686,N_6220,N_6177);
or U6687 (N_6687,N_6117,N_6465);
or U6688 (N_6688,N_6071,N_6003);
xnor U6689 (N_6689,N_6041,N_6189);
xnor U6690 (N_6690,N_6228,N_6140);
xnor U6691 (N_6691,N_6027,N_6203);
nor U6692 (N_6692,N_6437,N_6159);
nand U6693 (N_6693,N_6319,N_6464);
and U6694 (N_6694,N_6239,N_6374);
nor U6695 (N_6695,N_6137,N_6066);
nand U6696 (N_6696,N_6317,N_6401);
xnor U6697 (N_6697,N_6102,N_6421);
xnor U6698 (N_6698,N_6151,N_6247);
or U6699 (N_6699,N_6249,N_6331);
or U6700 (N_6700,N_6256,N_6202);
nor U6701 (N_6701,N_6124,N_6197);
or U6702 (N_6702,N_6356,N_6424);
xor U6703 (N_6703,N_6369,N_6250);
or U6704 (N_6704,N_6246,N_6125);
or U6705 (N_6705,N_6312,N_6074);
and U6706 (N_6706,N_6273,N_6135);
and U6707 (N_6707,N_6398,N_6431);
or U6708 (N_6708,N_6205,N_6105);
and U6709 (N_6709,N_6277,N_6131);
and U6710 (N_6710,N_6346,N_6199);
xor U6711 (N_6711,N_6156,N_6451);
and U6712 (N_6712,N_6324,N_6040);
nand U6713 (N_6713,N_6215,N_6323);
and U6714 (N_6714,N_6387,N_6056);
nor U6715 (N_6715,N_6266,N_6360);
nand U6716 (N_6716,N_6286,N_6287);
and U6717 (N_6717,N_6414,N_6377);
or U6718 (N_6718,N_6463,N_6306);
or U6719 (N_6719,N_6058,N_6077);
or U6720 (N_6720,N_6073,N_6046);
and U6721 (N_6721,N_6165,N_6132);
nand U6722 (N_6722,N_6126,N_6035);
or U6723 (N_6723,N_6301,N_6418);
nand U6724 (N_6724,N_6329,N_6337);
or U6725 (N_6725,N_6128,N_6350);
nand U6726 (N_6726,N_6009,N_6019);
nor U6727 (N_6727,N_6174,N_6488);
xnor U6728 (N_6728,N_6443,N_6479);
nand U6729 (N_6729,N_6413,N_6020);
and U6730 (N_6730,N_6415,N_6485);
nand U6731 (N_6731,N_6261,N_6295);
or U6732 (N_6732,N_6063,N_6087);
nand U6733 (N_6733,N_6048,N_6311);
or U6734 (N_6734,N_6049,N_6282);
nand U6735 (N_6735,N_6482,N_6339);
and U6736 (N_6736,N_6243,N_6410);
nor U6737 (N_6737,N_6440,N_6075);
nor U6738 (N_6738,N_6168,N_6141);
nor U6739 (N_6739,N_6213,N_6428);
nand U6740 (N_6740,N_6033,N_6380);
or U6741 (N_6741,N_6481,N_6138);
or U6742 (N_6742,N_6162,N_6477);
or U6743 (N_6743,N_6242,N_6107);
nor U6744 (N_6744,N_6257,N_6484);
nand U6745 (N_6745,N_6244,N_6098);
nand U6746 (N_6746,N_6025,N_6240);
nor U6747 (N_6747,N_6267,N_6417);
nor U6748 (N_6748,N_6493,N_6348);
nand U6749 (N_6749,N_6403,N_6393);
xor U6750 (N_6750,N_6374,N_6302);
nand U6751 (N_6751,N_6428,N_6476);
and U6752 (N_6752,N_6115,N_6012);
nor U6753 (N_6753,N_6104,N_6480);
or U6754 (N_6754,N_6424,N_6022);
nor U6755 (N_6755,N_6018,N_6458);
nor U6756 (N_6756,N_6487,N_6162);
and U6757 (N_6757,N_6318,N_6338);
or U6758 (N_6758,N_6187,N_6324);
or U6759 (N_6759,N_6407,N_6320);
and U6760 (N_6760,N_6032,N_6234);
nor U6761 (N_6761,N_6308,N_6044);
or U6762 (N_6762,N_6326,N_6374);
and U6763 (N_6763,N_6443,N_6126);
or U6764 (N_6764,N_6036,N_6258);
nand U6765 (N_6765,N_6012,N_6063);
nor U6766 (N_6766,N_6225,N_6492);
and U6767 (N_6767,N_6027,N_6329);
or U6768 (N_6768,N_6489,N_6116);
nand U6769 (N_6769,N_6490,N_6170);
nand U6770 (N_6770,N_6347,N_6000);
nor U6771 (N_6771,N_6256,N_6414);
xnor U6772 (N_6772,N_6072,N_6245);
and U6773 (N_6773,N_6204,N_6202);
xor U6774 (N_6774,N_6294,N_6026);
xor U6775 (N_6775,N_6481,N_6202);
xnor U6776 (N_6776,N_6157,N_6451);
xnor U6777 (N_6777,N_6286,N_6468);
and U6778 (N_6778,N_6096,N_6185);
and U6779 (N_6779,N_6436,N_6023);
nand U6780 (N_6780,N_6348,N_6470);
nor U6781 (N_6781,N_6086,N_6446);
and U6782 (N_6782,N_6418,N_6466);
or U6783 (N_6783,N_6324,N_6049);
nand U6784 (N_6784,N_6491,N_6222);
xor U6785 (N_6785,N_6055,N_6282);
nor U6786 (N_6786,N_6115,N_6065);
nor U6787 (N_6787,N_6482,N_6116);
nor U6788 (N_6788,N_6127,N_6421);
and U6789 (N_6789,N_6182,N_6136);
nand U6790 (N_6790,N_6227,N_6484);
nand U6791 (N_6791,N_6010,N_6157);
nor U6792 (N_6792,N_6142,N_6126);
xnor U6793 (N_6793,N_6209,N_6037);
and U6794 (N_6794,N_6051,N_6221);
nand U6795 (N_6795,N_6032,N_6250);
or U6796 (N_6796,N_6358,N_6374);
nand U6797 (N_6797,N_6184,N_6377);
nor U6798 (N_6798,N_6144,N_6034);
xor U6799 (N_6799,N_6446,N_6084);
nor U6800 (N_6800,N_6227,N_6246);
nand U6801 (N_6801,N_6279,N_6309);
or U6802 (N_6802,N_6100,N_6353);
or U6803 (N_6803,N_6171,N_6302);
nor U6804 (N_6804,N_6482,N_6479);
and U6805 (N_6805,N_6192,N_6221);
nand U6806 (N_6806,N_6218,N_6233);
nand U6807 (N_6807,N_6162,N_6228);
or U6808 (N_6808,N_6093,N_6183);
or U6809 (N_6809,N_6232,N_6306);
or U6810 (N_6810,N_6221,N_6419);
and U6811 (N_6811,N_6372,N_6185);
xnor U6812 (N_6812,N_6011,N_6177);
and U6813 (N_6813,N_6181,N_6108);
and U6814 (N_6814,N_6346,N_6081);
nor U6815 (N_6815,N_6012,N_6064);
nor U6816 (N_6816,N_6078,N_6027);
or U6817 (N_6817,N_6044,N_6134);
or U6818 (N_6818,N_6385,N_6255);
and U6819 (N_6819,N_6019,N_6183);
or U6820 (N_6820,N_6120,N_6214);
nand U6821 (N_6821,N_6428,N_6333);
or U6822 (N_6822,N_6212,N_6222);
nor U6823 (N_6823,N_6476,N_6050);
or U6824 (N_6824,N_6046,N_6210);
nand U6825 (N_6825,N_6215,N_6002);
and U6826 (N_6826,N_6101,N_6065);
or U6827 (N_6827,N_6064,N_6185);
or U6828 (N_6828,N_6281,N_6456);
nor U6829 (N_6829,N_6044,N_6046);
or U6830 (N_6830,N_6448,N_6222);
and U6831 (N_6831,N_6072,N_6191);
or U6832 (N_6832,N_6140,N_6170);
or U6833 (N_6833,N_6251,N_6449);
or U6834 (N_6834,N_6209,N_6167);
and U6835 (N_6835,N_6252,N_6488);
and U6836 (N_6836,N_6096,N_6392);
or U6837 (N_6837,N_6161,N_6438);
or U6838 (N_6838,N_6465,N_6229);
and U6839 (N_6839,N_6029,N_6389);
nand U6840 (N_6840,N_6302,N_6237);
and U6841 (N_6841,N_6143,N_6470);
or U6842 (N_6842,N_6134,N_6463);
and U6843 (N_6843,N_6031,N_6135);
xor U6844 (N_6844,N_6068,N_6443);
or U6845 (N_6845,N_6020,N_6055);
or U6846 (N_6846,N_6258,N_6209);
or U6847 (N_6847,N_6383,N_6404);
and U6848 (N_6848,N_6399,N_6144);
nand U6849 (N_6849,N_6090,N_6493);
or U6850 (N_6850,N_6263,N_6085);
nand U6851 (N_6851,N_6224,N_6333);
nand U6852 (N_6852,N_6277,N_6475);
nor U6853 (N_6853,N_6478,N_6243);
nand U6854 (N_6854,N_6177,N_6052);
and U6855 (N_6855,N_6402,N_6159);
nor U6856 (N_6856,N_6389,N_6444);
xor U6857 (N_6857,N_6058,N_6380);
nor U6858 (N_6858,N_6211,N_6039);
or U6859 (N_6859,N_6328,N_6286);
nor U6860 (N_6860,N_6157,N_6264);
and U6861 (N_6861,N_6461,N_6241);
or U6862 (N_6862,N_6337,N_6372);
and U6863 (N_6863,N_6375,N_6143);
or U6864 (N_6864,N_6152,N_6285);
or U6865 (N_6865,N_6049,N_6020);
and U6866 (N_6866,N_6487,N_6165);
nand U6867 (N_6867,N_6203,N_6316);
nor U6868 (N_6868,N_6132,N_6173);
nand U6869 (N_6869,N_6207,N_6342);
and U6870 (N_6870,N_6441,N_6272);
and U6871 (N_6871,N_6189,N_6381);
or U6872 (N_6872,N_6253,N_6258);
nand U6873 (N_6873,N_6028,N_6060);
xor U6874 (N_6874,N_6020,N_6079);
or U6875 (N_6875,N_6300,N_6420);
nor U6876 (N_6876,N_6398,N_6429);
and U6877 (N_6877,N_6194,N_6104);
or U6878 (N_6878,N_6114,N_6022);
and U6879 (N_6879,N_6103,N_6374);
or U6880 (N_6880,N_6152,N_6498);
and U6881 (N_6881,N_6299,N_6278);
nand U6882 (N_6882,N_6091,N_6154);
and U6883 (N_6883,N_6106,N_6316);
xor U6884 (N_6884,N_6401,N_6199);
nand U6885 (N_6885,N_6418,N_6136);
or U6886 (N_6886,N_6202,N_6147);
nor U6887 (N_6887,N_6084,N_6462);
or U6888 (N_6888,N_6031,N_6229);
or U6889 (N_6889,N_6040,N_6320);
nand U6890 (N_6890,N_6252,N_6015);
or U6891 (N_6891,N_6443,N_6353);
and U6892 (N_6892,N_6222,N_6351);
xor U6893 (N_6893,N_6489,N_6329);
or U6894 (N_6894,N_6045,N_6403);
nor U6895 (N_6895,N_6020,N_6193);
and U6896 (N_6896,N_6349,N_6289);
nor U6897 (N_6897,N_6494,N_6310);
nand U6898 (N_6898,N_6092,N_6182);
or U6899 (N_6899,N_6185,N_6119);
nand U6900 (N_6900,N_6206,N_6248);
nand U6901 (N_6901,N_6183,N_6054);
or U6902 (N_6902,N_6374,N_6271);
and U6903 (N_6903,N_6435,N_6357);
nor U6904 (N_6904,N_6063,N_6237);
and U6905 (N_6905,N_6021,N_6484);
or U6906 (N_6906,N_6439,N_6056);
or U6907 (N_6907,N_6093,N_6346);
nor U6908 (N_6908,N_6188,N_6184);
and U6909 (N_6909,N_6351,N_6469);
nand U6910 (N_6910,N_6403,N_6476);
xnor U6911 (N_6911,N_6300,N_6426);
and U6912 (N_6912,N_6097,N_6495);
or U6913 (N_6913,N_6040,N_6474);
xor U6914 (N_6914,N_6209,N_6007);
and U6915 (N_6915,N_6273,N_6426);
xnor U6916 (N_6916,N_6391,N_6117);
nor U6917 (N_6917,N_6102,N_6417);
or U6918 (N_6918,N_6288,N_6223);
nand U6919 (N_6919,N_6284,N_6173);
nor U6920 (N_6920,N_6087,N_6457);
or U6921 (N_6921,N_6394,N_6092);
nor U6922 (N_6922,N_6327,N_6420);
nand U6923 (N_6923,N_6437,N_6143);
nand U6924 (N_6924,N_6429,N_6331);
or U6925 (N_6925,N_6400,N_6334);
xnor U6926 (N_6926,N_6173,N_6080);
and U6927 (N_6927,N_6322,N_6392);
and U6928 (N_6928,N_6397,N_6194);
nor U6929 (N_6929,N_6256,N_6022);
nand U6930 (N_6930,N_6173,N_6050);
or U6931 (N_6931,N_6019,N_6474);
nand U6932 (N_6932,N_6460,N_6411);
nor U6933 (N_6933,N_6357,N_6099);
and U6934 (N_6934,N_6257,N_6002);
xor U6935 (N_6935,N_6096,N_6341);
nand U6936 (N_6936,N_6422,N_6270);
or U6937 (N_6937,N_6178,N_6278);
and U6938 (N_6938,N_6336,N_6132);
nand U6939 (N_6939,N_6199,N_6193);
or U6940 (N_6940,N_6466,N_6181);
and U6941 (N_6941,N_6063,N_6331);
or U6942 (N_6942,N_6461,N_6412);
and U6943 (N_6943,N_6260,N_6346);
nor U6944 (N_6944,N_6354,N_6016);
nor U6945 (N_6945,N_6128,N_6309);
or U6946 (N_6946,N_6220,N_6334);
and U6947 (N_6947,N_6008,N_6290);
nor U6948 (N_6948,N_6174,N_6063);
nor U6949 (N_6949,N_6131,N_6120);
nand U6950 (N_6950,N_6450,N_6338);
nor U6951 (N_6951,N_6396,N_6252);
nand U6952 (N_6952,N_6259,N_6135);
nand U6953 (N_6953,N_6161,N_6136);
and U6954 (N_6954,N_6213,N_6437);
nand U6955 (N_6955,N_6182,N_6346);
nor U6956 (N_6956,N_6075,N_6261);
nand U6957 (N_6957,N_6378,N_6414);
nand U6958 (N_6958,N_6238,N_6271);
nor U6959 (N_6959,N_6111,N_6318);
nand U6960 (N_6960,N_6200,N_6198);
nor U6961 (N_6961,N_6217,N_6048);
or U6962 (N_6962,N_6323,N_6392);
xor U6963 (N_6963,N_6234,N_6137);
and U6964 (N_6964,N_6346,N_6486);
xnor U6965 (N_6965,N_6042,N_6077);
nand U6966 (N_6966,N_6075,N_6446);
and U6967 (N_6967,N_6322,N_6066);
nand U6968 (N_6968,N_6480,N_6215);
and U6969 (N_6969,N_6190,N_6469);
and U6970 (N_6970,N_6123,N_6443);
nand U6971 (N_6971,N_6309,N_6085);
and U6972 (N_6972,N_6373,N_6378);
and U6973 (N_6973,N_6416,N_6070);
xnor U6974 (N_6974,N_6258,N_6247);
and U6975 (N_6975,N_6330,N_6115);
and U6976 (N_6976,N_6405,N_6407);
and U6977 (N_6977,N_6452,N_6461);
nor U6978 (N_6978,N_6192,N_6335);
and U6979 (N_6979,N_6282,N_6059);
and U6980 (N_6980,N_6068,N_6087);
or U6981 (N_6981,N_6479,N_6317);
nor U6982 (N_6982,N_6070,N_6245);
nand U6983 (N_6983,N_6237,N_6342);
or U6984 (N_6984,N_6423,N_6116);
and U6985 (N_6985,N_6038,N_6390);
nand U6986 (N_6986,N_6043,N_6300);
nor U6987 (N_6987,N_6354,N_6112);
nor U6988 (N_6988,N_6084,N_6334);
and U6989 (N_6989,N_6354,N_6344);
or U6990 (N_6990,N_6386,N_6494);
or U6991 (N_6991,N_6320,N_6275);
xor U6992 (N_6992,N_6341,N_6249);
and U6993 (N_6993,N_6223,N_6072);
nor U6994 (N_6994,N_6159,N_6061);
nor U6995 (N_6995,N_6272,N_6479);
or U6996 (N_6996,N_6215,N_6396);
xnor U6997 (N_6997,N_6038,N_6314);
and U6998 (N_6998,N_6051,N_6447);
nand U6999 (N_6999,N_6335,N_6375);
nor U7000 (N_7000,N_6745,N_6993);
xor U7001 (N_7001,N_6977,N_6690);
and U7002 (N_7002,N_6575,N_6851);
and U7003 (N_7003,N_6568,N_6925);
or U7004 (N_7004,N_6606,N_6754);
nand U7005 (N_7005,N_6639,N_6817);
and U7006 (N_7006,N_6789,N_6848);
and U7007 (N_7007,N_6884,N_6862);
or U7008 (N_7008,N_6670,N_6974);
or U7009 (N_7009,N_6816,N_6822);
nand U7010 (N_7010,N_6538,N_6820);
nand U7011 (N_7011,N_6623,N_6635);
and U7012 (N_7012,N_6604,N_6791);
xnor U7013 (N_7013,N_6781,N_6585);
and U7014 (N_7014,N_6837,N_6890);
nand U7015 (N_7015,N_6874,N_6809);
or U7016 (N_7016,N_6861,N_6696);
nand U7017 (N_7017,N_6731,N_6857);
nand U7018 (N_7018,N_6642,N_6998);
nand U7019 (N_7019,N_6919,N_6864);
nand U7020 (N_7020,N_6782,N_6869);
nor U7021 (N_7021,N_6834,N_6981);
and U7022 (N_7022,N_6935,N_6654);
nor U7023 (N_7023,N_6888,N_6714);
and U7024 (N_7024,N_6866,N_6910);
nor U7025 (N_7025,N_6899,N_6689);
nor U7026 (N_7026,N_6510,N_6865);
nor U7027 (N_7027,N_6545,N_6921);
or U7028 (N_7028,N_6613,N_6724);
and U7029 (N_7029,N_6560,N_6579);
nand U7030 (N_7030,N_6661,N_6569);
or U7031 (N_7031,N_6588,N_6767);
xnor U7032 (N_7032,N_6602,N_6741);
and U7033 (N_7033,N_6664,N_6965);
and U7034 (N_7034,N_6924,N_6543);
and U7035 (N_7035,N_6675,N_6853);
and U7036 (N_7036,N_6967,N_6772);
nand U7037 (N_7037,N_6502,N_6508);
nor U7038 (N_7038,N_6760,N_6906);
nor U7039 (N_7039,N_6643,N_6999);
nor U7040 (N_7040,N_6567,N_6909);
nor U7041 (N_7041,N_6950,N_6761);
or U7042 (N_7042,N_6646,N_6892);
xor U7043 (N_7043,N_6738,N_6518);
or U7044 (N_7044,N_6946,N_6917);
and U7045 (N_7045,N_6559,N_6778);
nor U7046 (N_7046,N_6651,N_6766);
or U7047 (N_7047,N_6563,N_6612);
and U7048 (N_7048,N_6841,N_6706);
or U7049 (N_7049,N_6807,N_6686);
nand U7050 (N_7050,N_6663,N_6849);
xnor U7051 (N_7051,N_6926,N_6882);
and U7052 (N_7052,N_6786,N_6871);
nor U7053 (N_7053,N_6665,N_6511);
xor U7054 (N_7054,N_6743,N_6934);
or U7055 (N_7055,N_6995,N_6962);
nand U7056 (N_7056,N_6501,N_6734);
nor U7057 (N_7057,N_6891,N_6947);
or U7058 (N_7058,N_6943,N_6933);
nand U7059 (N_7059,N_6688,N_6544);
nand U7060 (N_7060,N_6880,N_6824);
nor U7061 (N_7061,N_6595,N_6790);
xor U7062 (N_7062,N_6777,N_6572);
or U7063 (N_7063,N_6955,N_6509);
or U7064 (N_7064,N_6598,N_6729);
nor U7065 (N_7065,N_6617,N_6603);
and U7066 (N_7066,N_6832,N_6573);
nor U7067 (N_7067,N_6533,N_6942);
or U7068 (N_7068,N_6607,N_6666);
or U7069 (N_7069,N_6526,N_6730);
and U7070 (N_7070,N_6881,N_6574);
or U7071 (N_7071,N_6979,N_6895);
and U7072 (N_7072,N_6902,N_6991);
or U7073 (N_7073,N_6626,N_6831);
and U7074 (N_7074,N_6779,N_6703);
and U7075 (N_7075,N_6505,N_6540);
xor U7076 (N_7076,N_6630,N_6762);
nand U7077 (N_7077,N_6927,N_6571);
xnor U7078 (N_7078,N_6717,N_6845);
nand U7079 (N_7079,N_6692,N_6719);
or U7080 (N_7080,N_6922,N_6968);
or U7081 (N_7081,N_6829,N_6812);
nor U7082 (N_7082,N_6860,N_6645);
nand U7083 (N_7083,N_6650,N_6911);
nor U7084 (N_7084,N_6907,N_6512);
or U7085 (N_7085,N_6600,N_6589);
and U7086 (N_7086,N_6876,N_6770);
nand U7087 (N_7087,N_6673,N_6695);
nand U7088 (N_7088,N_6632,N_6608);
nand U7089 (N_7089,N_6564,N_6804);
and U7090 (N_7090,N_6836,N_6854);
nor U7091 (N_7091,N_6699,N_6513);
and U7092 (N_7092,N_6539,N_6893);
or U7093 (N_7093,N_6811,N_6903);
nor U7094 (N_7094,N_6616,N_6964);
and U7095 (N_7095,N_6923,N_6532);
nor U7096 (N_7096,N_6522,N_6610);
xor U7097 (N_7097,N_6697,N_6708);
nor U7098 (N_7098,N_6558,N_6879);
or U7099 (N_7099,N_6983,N_6705);
and U7100 (N_7100,N_6682,N_6954);
nand U7101 (N_7101,N_6780,N_6769);
and U7102 (N_7102,N_6725,N_6587);
and U7103 (N_7103,N_6792,N_6775);
xor U7104 (N_7104,N_6728,N_6683);
nand U7105 (N_7105,N_6858,N_6548);
nor U7106 (N_7106,N_6840,N_6994);
or U7107 (N_7107,N_6868,N_6514);
nor U7108 (N_7108,N_6693,N_6808);
nor U7109 (N_7109,N_6667,N_6737);
xor U7110 (N_7110,N_6529,N_6830);
nor U7111 (N_7111,N_6839,N_6628);
and U7112 (N_7112,N_6521,N_6631);
nor U7113 (N_7113,N_6704,N_6713);
nor U7114 (N_7114,N_6855,N_6932);
and U7115 (N_7115,N_6536,N_6669);
nand U7116 (N_7116,N_6668,N_6582);
nor U7117 (N_7117,N_6712,N_6877);
nand U7118 (N_7118,N_6984,N_6685);
or U7119 (N_7119,N_6570,N_6949);
or U7120 (N_7120,N_6894,N_6788);
nor U7121 (N_7121,N_6959,N_6856);
nand U7122 (N_7122,N_6875,N_6503);
or U7123 (N_7123,N_6805,N_6936);
and U7124 (N_7124,N_6937,N_6889);
nand U7125 (N_7125,N_6594,N_6944);
nor U7126 (N_7126,N_6739,N_6838);
or U7127 (N_7127,N_6684,N_6883);
or U7128 (N_7128,N_6793,N_6753);
nor U7129 (N_7129,N_6679,N_6986);
and U7130 (N_7130,N_6952,N_6900);
or U7131 (N_7131,N_6593,N_6990);
or U7132 (N_7132,N_6878,N_6732);
nand U7133 (N_7133,N_6658,N_6806);
and U7134 (N_7134,N_6987,N_6549);
nand U7135 (N_7135,N_6957,N_6972);
or U7136 (N_7136,N_6687,N_6597);
and U7137 (N_7137,N_6826,N_6721);
or U7138 (N_7138,N_6711,N_6970);
or U7139 (N_7139,N_6751,N_6859);
or U7140 (N_7140,N_6726,N_6691);
or U7141 (N_7141,N_6681,N_6784);
xor U7142 (N_7142,N_6976,N_6678);
nand U7143 (N_7143,N_6827,N_6759);
and U7144 (N_7144,N_6870,N_6621);
or U7145 (N_7145,N_6629,N_6918);
and U7146 (N_7146,N_6591,N_6541);
nor U7147 (N_7147,N_6525,N_6634);
nand U7148 (N_7148,N_6656,N_6819);
xnor U7149 (N_7149,N_6698,N_6546);
nor U7150 (N_7150,N_6552,N_6709);
and U7151 (N_7151,N_6615,N_6823);
and U7152 (N_7152,N_6537,N_6966);
xor U7153 (N_7153,N_6961,N_6755);
and U7154 (N_7154,N_6746,N_6980);
nand U7155 (N_7155,N_6872,N_6528);
nor U7156 (N_7156,N_6653,N_6660);
or U7157 (N_7157,N_6583,N_6584);
or U7158 (N_7158,N_6763,N_6914);
nor U7159 (N_7159,N_6867,N_6561);
xnor U7160 (N_7160,N_6920,N_6672);
or U7161 (N_7161,N_6785,N_6988);
nor U7162 (N_7162,N_6542,N_6749);
nand U7163 (N_7163,N_6931,N_6727);
nor U7164 (N_7164,N_6659,N_6647);
nand U7165 (N_7165,N_6835,N_6985);
or U7166 (N_7166,N_6723,N_6633);
nand U7167 (N_7167,N_6887,N_6800);
xor U7168 (N_7168,N_6655,N_6524);
nand U7169 (N_7169,N_6637,N_6908);
nor U7170 (N_7170,N_6756,N_6733);
nand U7171 (N_7171,N_6527,N_6752);
nand U7172 (N_7172,N_6873,N_6515);
and U7173 (N_7173,N_6748,N_6554);
nand U7174 (N_7174,N_6904,N_6847);
and U7175 (N_7175,N_6551,N_6566);
xor U7176 (N_7176,N_6940,N_6818);
and U7177 (N_7177,N_6958,N_6519);
nor U7178 (N_7178,N_6941,N_6565);
nor U7179 (N_7179,N_6677,N_6517);
or U7180 (N_7180,N_6747,N_6843);
or U7181 (N_7181,N_6576,N_6765);
and U7182 (N_7182,N_6562,N_6951);
and U7183 (N_7183,N_6641,N_6956);
nand U7184 (N_7184,N_6624,N_6774);
nand U7185 (N_7185,N_6844,N_6520);
nor U7186 (N_7186,N_6744,N_6796);
nor U7187 (N_7187,N_6803,N_6534);
or U7188 (N_7188,N_6531,N_6715);
and U7189 (N_7189,N_6863,N_6885);
or U7190 (N_7190,N_6969,N_6771);
or U7191 (N_7191,N_6928,N_6625);
nor U7192 (N_7192,N_6938,N_6586);
and U7193 (N_7193,N_6776,N_6702);
nor U7194 (N_7194,N_6953,N_6850);
and U7195 (N_7195,N_6674,N_6736);
and U7196 (N_7196,N_6578,N_6557);
and U7197 (N_7197,N_6618,N_6601);
and U7198 (N_7198,N_6802,N_6913);
nor U7199 (N_7199,N_6581,N_6821);
or U7200 (N_7200,N_6701,N_6722);
and U7201 (N_7201,N_6750,N_6758);
and U7202 (N_7202,N_6898,N_6997);
xor U7203 (N_7203,N_6814,N_6915);
nand U7204 (N_7204,N_6801,N_6963);
xor U7205 (N_7205,N_6523,N_6577);
nor U7206 (N_7206,N_6813,N_6718);
and U7207 (N_7207,N_6945,N_6757);
or U7208 (N_7208,N_6680,N_6773);
and U7209 (N_7209,N_6810,N_6912);
xnor U7210 (N_7210,N_6535,N_6901);
and U7211 (N_7211,N_6716,N_6700);
and U7212 (N_7212,N_6710,N_6556);
nor U7213 (N_7213,N_6742,N_6676);
or U7214 (N_7214,N_6797,N_6516);
nor U7215 (N_7215,N_6842,N_6794);
or U7216 (N_7216,N_6605,N_6504);
nand U7217 (N_7217,N_6886,N_6550);
or U7218 (N_7218,N_6939,N_6996);
nand U7219 (N_7219,N_6973,N_6982);
nand U7220 (N_7220,N_6735,N_6798);
nand U7221 (N_7221,N_6652,N_6580);
or U7222 (N_7222,N_6694,N_6764);
nand U7223 (N_7223,N_6530,N_6596);
nand U7224 (N_7224,N_6636,N_6671);
nand U7225 (N_7225,N_6989,N_6619);
or U7226 (N_7226,N_6897,N_6506);
or U7227 (N_7227,N_6644,N_6768);
and U7228 (N_7228,N_6846,N_6640);
or U7229 (N_7229,N_6833,N_6638);
or U7230 (N_7230,N_6787,N_6795);
nand U7231 (N_7231,N_6507,N_6948);
nand U7232 (N_7232,N_6707,N_6930);
xor U7233 (N_7233,N_6547,N_6649);
or U7234 (N_7234,N_6825,N_6975);
and U7235 (N_7235,N_6905,N_6720);
and U7236 (N_7236,N_6929,N_6662);
nor U7237 (N_7237,N_6916,N_6500);
and U7238 (N_7238,N_6971,N_6852);
nand U7239 (N_7239,N_6657,N_6592);
nand U7240 (N_7240,N_6620,N_6627);
nor U7241 (N_7241,N_6614,N_6799);
and U7242 (N_7242,N_6960,N_6740);
nand U7243 (N_7243,N_6590,N_6555);
or U7244 (N_7244,N_6622,N_6815);
xor U7245 (N_7245,N_6978,N_6896);
or U7246 (N_7246,N_6992,N_6611);
nand U7247 (N_7247,N_6783,N_6599);
nor U7248 (N_7248,N_6828,N_6609);
nor U7249 (N_7249,N_6648,N_6553);
and U7250 (N_7250,N_6557,N_6570);
or U7251 (N_7251,N_6828,N_6507);
or U7252 (N_7252,N_6844,N_6543);
nor U7253 (N_7253,N_6927,N_6653);
xnor U7254 (N_7254,N_6996,N_6677);
and U7255 (N_7255,N_6606,N_6575);
and U7256 (N_7256,N_6786,N_6956);
nor U7257 (N_7257,N_6911,N_6657);
nand U7258 (N_7258,N_6693,N_6623);
or U7259 (N_7259,N_6781,N_6523);
and U7260 (N_7260,N_6504,N_6927);
and U7261 (N_7261,N_6882,N_6763);
or U7262 (N_7262,N_6983,N_6802);
or U7263 (N_7263,N_6853,N_6726);
nand U7264 (N_7264,N_6745,N_6714);
nor U7265 (N_7265,N_6770,N_6817);
and U7266 (N_7266,N_6984,N_6986);
nor U7267 (N_7267,N_6817,N_6784);
nand U7268 (N_7268,N_6508,N_6708);
xor U7269 (N_7269,N_6542,N_6654);
or U7270 (N_7270,N_6833,N_6920);
or U7271 (N_7271,N_6877,N_6864);
nor U7272 (N_7272,N_6561,N_6618);
or U7273 (N_7273,N_6859,N_6530);
nand U7274 (N_7274,N_6697,N_6755);
nand U7275 (N_7275,N_6523,N_6985);
nor U7276 (N_7276,N_6979,N_6934);
nor U7277 (N_7277,N_6816,N_6999);
or U7278 (N_7278,N_6868,N_6985);
and U7279 (N_7279,N_6663,N_6522);
nand U7280 (N_7280,N_6911,N_6560);
nand U7281 (N_7281,N_6714,N_6712);
nand U7282 (N_7282,N_6960,N_6902);
or U7283 (N_7283,N_6647,N_6566);
and U7284 (N_7284,N_6895,N_6549);
and U7285 (N_7285,N_6998,N_6517);
and U7286 (N_7286,N_6939,N_6988);
and U7287 (N_7287,N_6849,N_6817);
and U7288 (N_7288,N_6812,N_6887);
nor U7289 (N_7289,N_6537,N_6524);
xnor U7290 (N_7290,N_6705,N_6889);
nor U7291 (N_7291,N_6882,N_6683);
nand U7292 (N_7292,N_6827,N_6863);
nor U7293 (N_7293,N_6551,N_6728);
nand U7294 (N_7294,N_6779,N_6549);
or U7295 (N_7295,N_6770,N_6702);
nor U7296 (N_7296,N_6694,N_6693);
or U7297 (N_7297,N_6604,N_6700);
and U7298 (N_7298,N_6979,N_6595);
xnor U7299 (N_7299,N_6652,N_6716);
nand U7300 (N_7300,N_6852,N_6608);
nor U7301 (N_7301,N_6827,N_6584);
and U7302 (N_7302,N_6689,N_6708);
nor U7303 (N_7303,N_6891,N_6916);
or U7304 (N_7304,N_6576,N_6862);
or U7305 (N_7305,N_6780,N_6642);
and U7306 (N_7306,N_6655,N_6604);
nand U7307 (N_7307,N_6685,N_6714);
nor U7308 (N_7308,N_6831,N_6730);
or U7309 (N_7309,N_6770,N_6786);
nand U7310 (N_7310,N_6896,N_6960);
and U7311 (N_7311,N_6512,N_6583);
nand U7312 (N_7312,N_6610,N_6719);
nor U7313 (N_7313,N_6983,N_6640);
nor U7314 (N_7314,N_6714,N_6626);
nand U7315 (N_7315,N_6696,N_6666);
or U7316 (N_7316,N_6596,N_6566);
and U7317 (N_7317,N_6925,N_6655);
nor U7318 (N_7318,N_6850,N_6643);
or U7319 (N_7319,N_6559,N_6796);
or U7320 (N_7320,N_6805,N_6858);
nand U7321 (N_7321,N_6778,N_6599);
nand U7322 (N_7322,N_6872,N_6774);
or U7323 (N_7323,N_6653,N_6816);
or U7324 (N_7324,N_6680,N_6634);
or U7325 (N_7325,N_6883,N_6870);
or U7326 (N_7326,N_6990,N_6928);
nor U7327 (N_7327,N_6641,N_6728);
and U7328 (N_7328,N_6741,N_6882);
nand U7329 (N_7329,N_6742,N_6523);
and U7330 (N_7330,N_6548,N_6966);
xnor U7331 (N_7331,N_6949,N_6960);
nand U7332 (N_7332,N_6722,N_6898);
nor U7333 (N_7333,N_6645,N_6591);
xor U7334 (N_7334,N_6566,N_6809);
nor U7335 (N_7335,N_6648,N_6829);
nor U7336 (N_7336,N_6549,N_6638);
and U7337 (N_7337,N_6792,N_6652);
xnor U7338 (N_7338,N_6823,N_6670);
or U7339 (N_7339,N_6872,N_6619);
and U7340 (N_7340,N_6980,N_6971);
nand U7341 (N_7341,N_6923,N_6592);
nand U7342 (N_7342,N_6723,N_6985);
nand U7343 (N_7343,N_6534,N_6742);
nor U7344 (N_7344,N_6810,N_6997);
and U7345 (N_7345,N_6891,N_6791);
or U7346 (N_7346,N_6546,N_6667);
and U7347 (N_7347,N_6683,N_6545);
and U7348 (N_7348,N_6554,N_6515);
and U7349 (N_7349,N_6726,N_6889);
nand U7350 (N_7350,N_6610,N_6576);
or U7351 (N_7351,N_6911,N_6819);
nor U7352 (N_7352,N_6674,N_6531);
and U7353 (N_7353,N_6781,N_6696);
nand U7354 (N_7354,N_6663,N_6923);
nor U7355 (N_7355,N_6681,N_6504);
xor U7356 (N_7356,N_6634,N_6949);
or U7357 (N_7357,N_6501,N_6549);
and U7358 (N_7358,N_6951,N_6845);
nor U7359 (N_7359,N_6807,N_6905);
or U7360 (N_7360,N_6767,N_6924);
nor U7361 (N_7361,N_6685,N_6980);
nor U7362 (N_7362,N_6681,N_6633);
xor U7363 (N_7363,N_6909,N_6618);
nand U7364 (N_7364,N_6636,N_6826);
and U7365 (N_7365,N_6847,N_6845);
or U7366 (N_7366,N_6951,N_6999);
nor U7367 (N_7367,N_6645,N_6824);
nor U7368 (N_7368,N_6524,N_6702);
xor U7369 (N_7369,N_6751,N_6920);
and U7370 (N_7370,N_6952,N_6557);
or U7371 (N_7371,N_6835,N_6803);
or U7372 (N_7372,N_6527,N_6749);
and U7373 (N_7373,N_6533,N_6755);
or U7374 (N_7374,N_6515,N_6787);
nor U7375 (N_7375,N_6507,N_6747);
nor U7376 (N_7376,N_6755,N_6708);
nor U7377 (N_7377,N_6884,N_6892);
nand U7378 (N_7378,N_6992,N_6985);
or U7379 (N_7379,N_6528,N_6597);
nand U7380 (N_7380,N_6967,N_6783);
nand U7381 (N_7381,N_6705,N_6573);
nand U7382 (N_7382,N_6808,N_6968);
nor U7383 (N_7383,N_6735,N_6550);
nor U7384 (N_7384,N_6654,N_6891);
nor U7385 (N_7385,N_6779,N_6819);
nand U7386 (N_7386,N_6617,N_6647);
or U7387 (N_7387,N_6851,N_6750);
nand U7388 (N_7388,N_6923,N_6557);
nand U7389 (N_7389,N_6593,N_6861);
nor U7390 (N_7390,N_6531,N_6817);
nor U7391 (N_7391,N_6529,N_6756);
xor U7392 (N_7392,N_6551,N_6698);
or U7393 (N_7393,N_6760,N_6733);
nand U7394 (N_7394,N_6950,N_6769);
and U7395 (N_7395,N_6784,N_6771);
nand U7396 (N_7396,N_6960,N_6500);
and U7397 (N_7397,N_6864,N_6876);
and U7398 (N_7398,N_6654,N_6897);
xor U7399 (N_7399,N_6707,N_6637);
nor U7400 (N_7400,N_6698,N_6572);
nand U7401 (N_7401,N_6804,N_6858);
or U7402 (N_7402,N_6772,N_6893);
nand U7403 (N_7403,N_6952,N_6953);
nand U7404 (N_7404,N_6550,N_6709);
and U7405 (N_7405,N_6651,N_6790);
nand U7406 (N_7406,N_6607,N_6613);
or U7407 (N_7407,N_6834,N_6793);
or U7408 (N_7408,N_6573,N_6522);
and U7409 (N_7409,N_6811,N_6798);
xnor U7410 (N_7410,N_6977,N_6801);
and U7411 (N_7411,N_6583,N_6762);
xnor U7412 (N_7412,N_6787,N_6589);
nand U7413 (N_7413,N_6738,N_6857);
nor U7414 (N_7414,N_6845,N_6856);
nand U7415 (N_7415,N_6734,N_6653);
xor U7416 (N_7416,N_6529,N_6978);
and U7417 (N_7417,N_6725,N_6926);
xor U7418 (N_7418,N_6517,N_6529);
nor U7419 (N_7419,N_6534,N_6957);
nor U7420 (N_7420,N_6948,N_6901);
and U7421 (N_7421,N_6734,N_6896);
xnor U7422 (N_7422,N_6811,N_6698);
xnor U7423 (N_7423,N_6695,N_6777);
nor U7424 (N_7424,N_6785,N_6673);
nor U7425 (N_7425,N_6583,N_6934);
nand U7426 (N_7426,N_6654,N_6503);
or U7427 (N_7427,N_6729,N_6754);
or U7428 (N_7428,N_6656,N_6924);
nor U7429 (N_7429,N_6968,N_6813);
and U7430 (N_7430,N_6944,N_6626);
nor U7431 (N_7431,N_6673,N_6963);
and U7432 (N_7432,N_6608,N_6950);
or U7433 (N_7433,N_6668,N_6569);
or U7434 (N_7434,N_6937,N_6879);
nand U7435 (N_7435,N_6577,N_6614);
or U7436 (N_7436,N_6512,N_6846);
nand U7437 (N_7437,N_6743,N_6781);
nor U7438 (N_7438,N_6690,N_6585);
or U7439 (N_7439,N_6969,N_6644);
and U7440 (N_7440,N_6755,N_6892);
or U7441 (N_7441,N_6711,N_6753);
and U7442 (N_7442,N_6735,N_6873);
or U7443 (N_7443,N_6620,N_6855);
nor U7444 (N_7444,N_6850,N_6795);
nor U7445 (N_7445,N_6856,N_6852);
nand U7446 (N_7446,N_6892,N_6887);
nand U7447 (N_7447,N_6658,N_6539);
and U7448 (N_7448,N_6567,N_6770);
and U7449 (N_7449,N_6826,N_6716);
and U7450 (N_7450,N_6547,N_6746);
or U7451 (N_7451,N_6857,N_6757);
and U7452 (N_7452,N_6939,N_6757);
and U7453 (N_7453,N_6919,N_6553);
nand U7454 (N_7454,N_6811,N_6766);
and U7455 (N_7455,N_6984,N_6957);
xor U7456 (N_7456,N_6673,N_6688);
and U7457 (N_7457,N_6531,N_6903);
nand U7458 (N_7458,N_6591,N_6553);
nand U7459 (N_7459,N_6529,N_6534);
and U7460 (N_7460,N_6959,N_6917);
and U7461 (N_7461,N_6561,N_6540);
and U7462 (N_7462,N_6677,N_6833);
nand U7463 (N_7463,N_6869,N_6761);
or U7464 (N_7464,N_6702,N_6748);
nor U7465 (N_7465,N_6590,N_6545);
nand U7466 (N_7466,N_6531,N_6942);
xnor U7467 (N_7467,N_6583,N_6743);
nor U7468 (N_7468,N_6852,N_6640);
and U7469 (N_7469,N_6652,N_6999);
nand U7470 (N_7470,N_6988,N_6891);
xor U7471 (N_7471,N_6606,N_6907);
or U7472 (N_7472,N_6996,N_6778);
xor U7473 (N_7473,N_6606,N_6902);
xnor U7474 (N_7474,N_6851,N_6628);
nand U7475 (N_7475,N_6575,N_6792);
or U7476 (N_7476,N_6617,N_6763);
or U7477 (N_7477,N_6554,N_6597);
nor U7478 (N_7478,N_6823,N_6920);
and U7479 (N_7479,N_6544,N_6845);
nor U7480 (N_7480,N_6981,N_6566);
nor U7481 (N_7481,N_6568,N_6855);
nand U7482 (N_7482,N_6832,N_6903);
nor U7483 (N_7483,N_6760,N_6543);
and U7484 (N_7484,N_6876,N_6707);
xor U7485 (N_7485,N_6558,N_6539);
and U7486 (N_7486,N_6580,N_6604);
or U7487 (N_7487,N_6860,N_6707);
nand U7488 (N_7488,N_6647,N_6908);
nor U7489 (N_7489,N_6591,N_6566);
nor U7490 (N_7490,N_6946,N_6548);
and U7491 (N_7491,N_6984,N_6775);
xnor U7492 (N_7492,N_6501,N_6770);
or U7493 (N_7493,N_6606,N_6540);
nand U7494 (N_7494,N_6836,N_6698);
and U7495 (N_7495,N_6507,N_6700);
or U7496 (N_7496,N_6841,N_6675);
or U7497 (N_7497,N_6643,N_6965);
nor U7498 (N_7498,N_6516,N_6642);
nor U7499 (N_7499,N_6589,N_6710);
nand U7500 (N_7500,N_7224,N_7424);
or U7501 (N_7501,N_7394,N_7242);
nand U7502 (N_7502,N_7074,N_7104);
nor U7503 (N_7503,N_7046,N_7232);
or U7504 (N_7504,N_7343,N_7111);
and U7505 (N_7505,N_7425,N_7214);
nand U7506 (N_7506,N_7441,N_7100);
and U7507 (N_7507,N_7238,N_7002);
nand U7508 (N_7508,N_7290,N_7344);
nand U7509 (N_7509,N_7346,N_7421);
xnor U7510 (N_7510,N_7118,N_7493);
or U7511 (N_7511,N_7397,N_7408);
xnor U7512 (N_7512,N_7079,N_7348);
and U7513 (N_7513,N_7021,N_7269);
and U7514 (N_7514,N_7075,N_7147);
or U7515 (N_7515,N_7045,N_7327);
and U7516 (N_7516,N_7057,N_7068);
or U7517 (N_7517,N_7124,N_7465);
nand U7518 (N_7518,N_7293,N_7399);
and U7519 (N_7519,N_7485,N_7011);
and U7520 (N_7520,N_7461,N_7098);
or U7521 (N_7521,N_7031,N_7001);
and U7522 (N_7522,N_7412,N_7127);
or U7523 (N_7523,N_7353,N_7299);
nor U7524 (N_7524,N_7492,N_7395);
nand U7525 (N_7525,N_7482,N_7150);
nand U7526 (N_7526,N_7082,N_7048);
and U7527 (N_7527,N_7372,N_7401);
nor U7528 (N_7528,N_7356,N_7429);
xnor U7529 (N_7529,N_7276,N_7324);
or U7530 (N_7530,N_7454,N_7404);
or U7531 (N_7531,N_7014,N_7360);
nand U7532 (N_7532,N_7230,N_7139);
nor U7533 (N_7533,N_7366,N_7208);
nor U7534 (N_7534,N_7379,N_7246);
nor U7535 (N_7535,N_7154,N_7215);
nor U7536 (N_7536,N_7019,N_7202);
nand U7537 (N_7537,N_7158,N_7298);
nor U7538 (N_7538,N_7283,N_7056);
and U7539 (N_7539,N_7198,N_7431);
nand U7540 (N_7540,N_7032,N_7320);
xnor U7541 (N_7541,N_7391,N_7420);
and U7542 (N_7542,N_7093,N_7132);
or U7543 (N_7543,N_7212,N_7103);
nand U7544 (N_7544,N_7140,N_7108);
nor U7545 (N_7545,N_7026,N_7171);
or U7546 (N_7546,N_7084,N_7222);
nand U7547 (N_7547,N_7277,N_7131);
nand U7548 (N_7548,N_7101,N_7125);
xnor U7549 (N_7549,N_7236,N_7115);
nor U7550 (N_7550,N_7162,N_7061);
nor U7551 (N_7551,N_7306,N_7245);
nand U7552 (N_7552,N_7389,N_7398);
xor U7553 (N_7553,N_7286,N_7000);
and U7554 (N_7554,N_7491,N_7313);
and U7555 (N_7555,N_7247,N_7219);
and U7556 (N_7556,N_7099,N_7237);
and U7557 (N_7557,N_7152,N_7228);
and U7558 (N_7558,N_7337,N_7328);
nand U7559 (N_7559,N_7062,N_7173);
or U7560 (N_7560,N_7241,N_7435);
xnor U7561 (N_7561,N_7392,N_7339);
nor U7562 (N_7562,N_7296,N_7250);
nand U7563 (N_7563,N_7326,N_7468);
nor U7564 (N_7564,N_7141,N_7488);
nand U7565 (N_7565,N_7134,N_7463);
nor U7566 (N_7566,N_7393,N_7373);
and U7567 (N_7567,N_7304,N_7357);
nor U7568 (N_7568,N_7013,N_7042);
and U7569 (N_7569,N_7225,N_7206);
nor U7570 (N_7570,N_7231,N_7483);
and U7571 (N_7571,N_7303,N_7292);
nor U7572 (N_7572,N_7092,N_7437);
or U7573 (N_7573,N_7137,N_7381);
nor U7574 (N_7574,N_7310,N_7333);
nand U7575 (N_7575,N_7414,N_7169);
or U7576 (N_7576,N_7462,N_7498);
nand U7577 (N_7577,N_7297,N_7406);
nor U7578 (N_7578,N_7018,N_7375);
nand U7579 (N_7579,N_7038,N_7440);
nand U7580 (N_7580,N_7063,N_7039);
xor U7581 (N_7581,N_7107,N_7151);
xnor U7582 (N_7582,N_7445,N_7340);
nand U7583 (N_7583,N_7480,N_7321);
or U7584 (N_7584,N_7442,N_7289);
or U7585 (N_7585,N_7365,N_7028);
and U7586 (N_7586,N_7204,N_7264);
nand U7587 (N_7587,N_7252,N_7364);
or U7588 (N_7588,N_7187,N_7471);
nand U7589 (N_7589,N_7097,N_7443);
nand U7590 (N_7590,N_7041,N_7170);
nand U7591 (N_7591,N_7050,N_7036);
nor U7592 (N_7592,N_7486,N_7265);
nand U7593 (N_7593,N_7155,N_7234);
nor U7594 (N_7594,N_7257,N_7243);
xnor U7595 (N_7595,N_7479,N_7410);
and U7596 (N_7596,N_7088,N_7168);
xor U7597 (N_7597,N_7496,N_7044);
nor U7598 (N_7598,N_7086,N_7126);
or U7599 (N_7599,N_7085,N_7199);
xor U7600 (N_7600,N_7278,N_7006);
or U7601 (N_7601,N_7163,N_7302);
nand U7602 (N_7602,N_7362,N_7260);
nor U7603 (N_7603,N_7027,N_7319);
or U7604 (N_7604,N_7288,N_7179);
nand U7605 (N_7605,N_7181,N_7453);
or U7606 (N_7606,N_7023,N_7122);
nand U7607 (N_7607,N_7316,N_7138);
nand U7608 (N_7608,N_7244,N_7015);
nand U7609 (N_7609,N_7294,N_7223);
nand U7610 (N_7610,N_7059,N_7087);
or U7611 (N_7611,N_7285,N_7120);
nor U7612 (N_7612,N_7361,N_7148);
nor U7613 (N_7613,N_7043,N_7334);
nor U7614 (N_7614,N_7254,N_7089);
or U7615 (N_7615,N_7012,N_7325);
nor U7616 (N_7616,N_7419,N_7142);
or U7617 (N_7617,N_7167,N_7227);
nor U7618 (N_7618,N_7109,N_7433);
and U7619 (N_7619,N_7428,N_7331);
nor U7620 (N_7620,N_7184,N_7080);
and U7621 (N_7621,N_7477,N_7472);
nor U7622 (N_7622,N_7121,N_7444);
and U7623 (N_7623,N_7300,N_7458);
and U7624 (N_7624,N_7197,N_7156);
nor U7625 (N_7625,N_7193,N_7055);
or U7626 (N_7626,N_7069,N_7270);
xnor U7627 (N_7627,N_7200,N_7210);
or U7628 (N_7628,N_7438,N_7487);
nand U7629 (N_7629,N_7309,N_7312);
nor U7630 (N_7630,N_7273,N_7083);
nand U7631 (N_7631,N_7267,N_7145);
nand U7632 (N_7632,N_7417,N_7218);
and U7633 (N_7633,N_7003,N_7456);
nand U7634 (N_7634,N_7460,N_7172);
nor U7635 (N_7635,N_7355,N_7363);
nand U7636 (N_7636,N_7473,N_7017);
nand U7637 (N_7637,N_7423,N_7060);
nor U7638 (N_7638,N_7338,N_7367);
nand U7639 (N_7639,N_7415,N_7317);
or U7640 (N_7640,N_7144,N_7426);
or U7641 (N_7641,N_7166,N_7239);
and U7642 (N_7642,N_7249,N_7434);
xor U7643 (N_7643,N_7129,N_7305);
nor U7644 (N_7644,N_7315,N_7371);
nor U7645 (N_7645,N_7024,N_7342);
or U7646 (N_7646,N_7047,N_7450);
or U7647 (N_7647,N_7157,N_7119);
or U7648 (N_7648,N_7077,N_7106);
or U7649 (N_7649,N_7016,N_7439);
nor U7650 (N_7650,N_7347,N_7221);
nand U7651 (N_7651,N_7114,N_7009);
and U7652 (N_7652,N_7400,N_7459);
or U7653 (N_7653,N_7490,N_7072);
and U7654 (N_7654,N_7275,N_7432);
or U7655 (N_7655,N_7318,N_7268);
xor U7656 (N_7656,N_7205,N_7448);
xor U7657 (N_7657,N_7413,N_7386);
nand U7658 (N_7658,N_7455,N_7418);
or U7659 (N_7659,N_7274,N_7180);
xnor U7660 (N_7660,N_7051,N_7235);
nor U7661 (N_7661,N_7110,N_7436);
and U7662 (N_7662,N_7495,N_7281);
or U7663 (N_7663,N_7064,N_7376);
nor U7664 (N_7664,N_7192,N_7476);
nor U7665 (N_7665,N_7071,N_7335);
nand U7666 (N_7666,N_7078,N_7378);
nand U7667 (N_7667,N_7383,N_7030);
and U7668 (N_7668,N_7311,N_7403);
and U7669 (N_7669,N_7308,N_7385);
and U7670 (N_7670,N_7066,N_7466);
or U7671 (N_7671,N_7484,N_7387);
or U7672 (N_7672,N_7175,N_7470);
and U7673 (N_7673,N_7329,N_7195);
and U7674 (N_7674,N_7209,N_7217);
xnor U7675 (N_7675,N_7033,N_7007);
or U7676 (N_7676,N_7136,N_7411);
or U7677 (N_7677,N_7314,N_7284);
or U7678 (N_7678,N_7095,N_7211);
or U7679 (N_7679,N_7262,N_7020);
nand U7680 (N_7680,N_7253,N_7377);
and U7681 (N_7681,N_7359,N_7146);
nor U7682 (N_7682,N_7186,N_7279);
nand U7683 (N_7683,N_7226,N_7475);
nand U7684 (N_7684,N_7004,N_7029);
xor U7685 (N_7685,N_7143,N_7322);
nand U7686 (N_7686,N_7464,N_7201);
nor U7687 (N_7687,N_7070,N_7053);
or U7688 (N_7688,N_7005,N_7280);
or U7689 (N_7689,N_7251,N_7457);
xor U7690 (N_7690,N_7213,N_7116);
nor U7691 (N_7691,N_7430,N_7178);
or U7692 (N_7692,N_7037,N_7368);
nor U7693 (N_7693,N_7094,N_7323);
nand U7694 (N_7694,N_7188,N_7332);
nand U7695 (N_7695,N_7291,N_7307);
nor U7696 (N_7696,N_7396,N_7161);
nor U7697 (N_7697,N_7194,N_7446);
and U7698 (N_7698,N_7165,N_7096);
and U7699 (N_7699,N_7220,N_7449);
nor U7700 (N_7700,N_7469,N_7422);
nand U7701 (N_7701,N_7499,N_7010);
or U7702 (N_7702,N_7133,N_7369);
or U7703 (N_7703,N_7341,N_7271);
and U7704 (N_7704,N_7117,N_7130);
nand U7705 (N_7705,N_7259,N_7350);
and U7706 (N_7706,N_7207,N_7049);
nor U7707 (N_7707,N_7052,N_7183);
nor U7708 (N_7708,N_7248,N_7330);
xnor U7709 (N_7709,N_7402,N_7352);
or U7710 (N_7710,N_7474,N_7489);
nor U7711 (N_7711,N_7380,N_7040);
or U7712 (N_7712,N_7481,N_7256);
and U7713 (N_7713,N_7497,N_7384);
xnor U7714 (N_7714,N_7164,N_7336);
nor U7715 (N_7715,N_7174,N_7416);
or U7716 (N_7716,N_7390,N_7022);
or U7717 (N_7717,N_7185,N_7409);
xor U7718 (N_7718,N_7405,N_7081);
nor U7719 (N_7719,N_7065,N_7189);
nand U7720 (N_7720,N_7282,N_7091);
nor U7721 (N_7721,N_7345,N_7478);
or U7722 (N_7722,N_7102,N_7008);
nor U7723 (N_7723,N_7153,N_7135);
or U7724 (N_7724,N_7176,N_7233);
nand U7725 (N_7725,N_7090,N_7216);
xor U7726 (N_7726,N_7258,N_7370);
nor U7727 (N_7727,N_7067,N_7159);
nand U7728 (N_7728,N_7447,N_7272);
or U7729 (N_7729,N_7128,N_7467);
or U7730 (N_7730,N_7240,N_7427);
or U7731 (N_7731,N_7349,N_7034);
and U7732 (N_7732,N_7388,N_7190);
or U7733 (N_7733,N_7255,N_7452);
nor U7734 (N_7734,N_7025,N_7177);
or U7735 (N_7735,N_7407,N_7382);
nand U7736 (N_7736,N_7229,N_7073);
nor U7737 (N_7737,N_7054,N_7494);
xor U7738 (N_7738,N_7266,N_7035);
nand U7739 (N_7739,N_7076,N_7358);
and U7740 (N_7740,N_7112,N_7160);
or U7741 (N_7741,N_7203,N_7351);
xnor U7742 (N_7742,N_7105,N_7191);
or U7743 (N_7743,N_7451,N_7374);
and U7744 (N_7744,N_7113,N_7287);
nand U7745 (N_7745,N_7182,N_7295);
or U7746 (N_7746,N_7301,N_7123);
or U7747 (N_7747,N_7263,N_7261);
nand U7748 (N_7748,N_7149,N_7196);
nand U7749 (N_7749,N_7058,N_7354);
and U7750 (N_7750,N_7361,N_7414);
and U7751 (N_7751,N_7217,N_7104);
nor U7752 (N_7752,N_7011,N_7002);
and U7753 (N_7753,N_7309,N_7151);
nand U7754 (N_7754,N_7327,N_7475);
nand U7755 (N_7755,N_7214,N_7161);
nor U7756 (N_7756,N_7267,N_7022);
or U7757 (N_7757,N_7385,N_7017);
xnor U7758 (N_7758,N_7316,N_7307);
xnor U7759 (N_7759,N_7327,N_7157);
nor U7760 (N_7760,N_7322,N_7422);
or U7761 (N_7761,N_7013,N_7132);
or U7762 (N_7762,N_7285,N_7408);
and U7763 (N_7763,N_7289,N_7306);
xor U7764 (N_7764,N_7128,N_7192);
nor U7765 (N_7765,N_7255,N_7250);
or U7766 (N_7766,N_7106,N_7147);
and U7767 (N_7767,N_7406,N_7309);
nor U7768 (N_7768,N_7216,N_7350);
and U7769 (N_7769,N_7418,N_7405);
nor U7770 (N_7770,N_7464,N_7485);
xnor U7771 (N_7771,N_7274,N_7209);
or U7772 (N_7772,N_7485,N_7010);
nand U7773 (N_7773,N_7175,N_7093);
xor U7774 (N_7774,N_7047,N_7279);
or U7775 (N_7775,N_7106,N_7376);
and U7776 (N_7776,N_7018,N_7006);
nand U7777 (N_7777,N_7482,N_7320);
nor U7778 (N_7778,N_7126,N_7030);
nand U7779 (N_7779,N_7082,N_7091);
and U7780 (N_7780,N_7131,N_7395);
xor U7781 (N_7781,N_7151,N_7422);
or U7782 (N_7782,N_7107,N_7118);
nand U7783 (N_7783,N_7400,N_7232);
nor U7784 (N_7784,N_7016,N_7019);
nor U7785 (N_7785,N_7318,N_7063);
nand U7786 (N_7786,N_7233,N_7007);
or U7787 (N_7787,N_7159,N_7295);
or U7788 (N_7788,N_7344,N_7407);
xnor U7789 (N_7789,N_7454,N_7030);
and U7790 (N_7790,N_7297,N_7484);
nand U7791 (N_7791,N_7302,N_7365);
and U7792 (N_7792,N_7242,N_7224);
nor U7793 (N_7793,N_7339,N_7435);
nor U7794 (N_7794,N_7023,N_7097);
nor U7795 (N_7795,N_7029,N_7256);
xnor U7796 (N_7796,N_7376,N_7258);
nand U7797 (N_7797,N_7022,N_7387);
xnor U7798 (N_7798,N_7248,N_7197);
nor U7799 (N_7799,N_7288,N_7319);
xnor U7800 (N_7800,N_7303,N_7018);
and U7801 (N_7801,N_7048,N_7086);
nand U7802 (N_7802,N_7235,N_7381);
nand U7803 (N_7803,N_7484,N_7211);
nor U7804 (N_7804,N_7356,N_7138);
nor U7805 (N_7805,N_7348,N_7330);
nand U7806 (N_7806,N_7331,N_7070);
nand U7807 (N_7807,N_7451,N_7201);
nand U7808 (N_7808,N_7004,N_7452);
and U7809 (N_7809,N_7080,N_7389);
nor U7810 (N_7810,N_7321,N_7325);
or U7811 (N_7811,N_7089,N_7325);
and U7812 (N_7812,N_7469,N_7172);
nor U7813 (N_7813,N_7494,N_7246);
nand U7814 (N_7814,N_7453,N_7342);
or U7815 (N_7815,N_7110,N_7482);
nand U7816 (N_7816,N_7360,N_7350);
nor U7817 (N_7817,N_7342,N_7119);
nor U7818 (N_7818,N_7433,N_7300);
xnor U7819 (N_7819,N_7499,N_7077);
nor U7820 (N_7820,N_7339,N_7249);
xnor U7821 (N_7821,N_7103,N_7384);
nor U7822 (N_7822,N_7046,N_7187);
and U7823 (N_7823,N_7234,N_7307);
nor U7824 (N_7824,N_7207,N_7451);
nor U7825 (N_7825,N_7404,N_7490);
xnor U7826 (N_7826,N_7054,N_7365);
nand U7827 (N_7827,N_7496,N_7472);
nor U7828 (N_7828,N_7364,N_7068);
nor U7829 (N_7829,N_7468,N_7018);
nor U7830 (N_7830,N_7044,N_7218);
nand U7831 (N_7831,N_7382,N_7024);
and U7832 (N_7832,N_7311,N_7346);
and U7833 (N_7833,N_7069,N_7472);
nand U7834 (N_7834,N_7141,N_7102);
nand U7835 (N_7835,N_7410,N_7289);
nand U7836 (N_7836,N_7476,N_7171);
and U7837 (N_7837,N_7255,N_7121);
nand U7838 (N_7838,N_7034,N_7227);
and U7839 (N_7839,N_7274,N_7113);
and U7840 (N_7840,N_7026,N_7029);
or U7841 (N_7841,N_7189,N_7117);
or U7842 (N_7842,N_7002,N_7263);
or U7843 (N_7843,N_7413,N_7248);
nand U7844 (N_7844,N_7076,N_7349);
xnor U7845 (N_7845,N_7185,N_7477);
or U7846 (N_7846,N_7095,N_7203);
nor U7847 (N_7847,N_7390,N_7329);
nor U7848 (N_7848,N_7056,N_7309);
or U7849 (N_7849,N_7410,N_7240);
nand U7850 (N_7850,N_7475,N_7125);
xnor U7851 (N_7851,N_7252,N_7194);
xor U7852 (N_7852,N_7449,N_7020);
nand U7853 (N_7853,N_7146,N_7460);
nand U7854 (N_7854,N_7473,N_7196);
nand U7855 (N_7855,N_7180,N_7330);
nor U7856 (N_7856,N_7471,N_7068);
nand U7857 (N_7857,N_7152,N_7456);
nand U7858 (N_7858,N_7193,N_7014);
nand U7859 (N_7859,N_7451,N_7368);
or U7860 (N_7860,N_7201,N_7478);
and U7861 (N_7861,N_7051,N_7424);
or U7862 (N_7862,N_7274,N_7433);
or U7863 (N_7863,N_7319,N_7189);
xnor U7864 (N_7864,N_7484,N_7086);
nand U7865 (N_7865,N_7172,N_7462);
nor U7866 (N_7866,N_7330,N_7208);
nand U7867 (N_7867,N_7224,N_7131);
nand U7868 (N_7868,N_7221,N_7218);
nand U7869 (N_7869,N_7114,N_7169);
nor U7870 (N_7870,N_7339,N_7038);
and U7871 (N_7871,N_7392,N_7446);
or U7872 (N_7872,N_7021,N_7439);
and U7873 (N_7873,N_7329,N_7056);
nand U7874 (N_7874,N_7122,N_7057);
xnor U7875 (N_7875,N_7266,N_7365);
nand U7876 (N_7876,N_7360,N_7431);
nand U7877 (N_7877,N_7499,N_7392);
xor U7878 (N_7878,N_7305,N_7294);
and U7879 (N_7879,N_7308,N_7107);
and U7880 (N_7880,N_7208,N_7041);
and U7881 (N_7881,N_7117,N_7421);
and U7882 (N_7882,N_7153,N_7132);
xor U7883 (N_7883,N_7366,N_7465);
nand U7884 (N_7884,N_7025,N_7167);
nor U7885 (N_7885,N_7172,N_7213);
or U7886 (N_7886,N_7251,N_7286);
nand U7887 (N_7887,N_7223,N_7058);
xor U7888 (N_7888,N_7445,N_7168);
nand U7889 (N_7889,N_7135,N_7186);
nor U7890 (N_7890,N_7155,N_7295);
or U7891 (N_7891,N_7106,N_7054);
nor U7892 (N_7892,N_7097,N_7107);
xor U7893 (N_7893,N_7367,N_7407);
or U7894 (N_7894,N_7412,N_7098);
nor U7895 (N_7895,N_7128,N_7095);
or U7896 (N_7896,N_7420,N_7257);
nand U7897 (N_7897,N_7051,N_7356);
and U7898 (N_7898,N_7204,N_7248);
nand U7899 (N_7899,N_7275,N_7054);
nor U7900 (N_7900,N_7448,N_7075);
and U7901 (N_7901,N_7317,N_7285);
and U7902 (N_7902,N_7355,N_7166);
and U7903 (N_7903,N_7014,N_7278);
and U7904 (N_7904,N_7040,N_7342);
or U7905 (N_7905,N_7361,N_7332);
nor U7906 (N_7906,N_7146,N_7046);
xnor U7907 (N_7907,N_7180,N_7461);
and U7908 (N_7908,N_7496,N_7102);
and U7909 (N_7909,N_7328,N_7186);
and U7910 (N_7910,N_7127,N_7444);
nand U7911 (N_7911,N_7268,N_7461);
nand U7912 (N_7912,N_7135,N_7127);
nand U7913 (N_7913,N_7196,N_7145);
and U7914 (N_7914,N_7378,N_7392);
or U7915 (N_7915,N_7305,N_7053);
and U7916 (N_7916,N_7196,N_7453);
xor U7917 (N_7917,N_7259,N_7167);
nand U7918 (N_7918,N_7401,N_7008);
nand U7919 (N_7919,N_7304,N_7488);
xnor U7920 (N_7920,N_7319,N_7393);
nor U7921 (N_7921,N_7100,N_7016);
or U7922 (N_7922,N_7226,N_7188);
xnor U7923 (N_7923,N_7432,N_7487);
and U7924 (N_7924,N_7108,N_7459);
nand U7925 (N_7925,N_7406,N_7208);
nand U7926 (N_7926,N_7174,N_7452);
and U7927 (N_7927,N_7342,N_7272);
xnor U7928 (N_7928,N_7280,N_7118);
nor U7929 (N_7929,N_7044,N_7477);
xnor U7930 (N_7930,N_7405,N_7170);
and U7931 (N_7931,N_7402,N_7035);
nor U7932 (N_7932,N_7299,N_7253);
or U7933 (N_7933,N_7377,N_7107);
nor U7934 (N_7934,N_7323,N_7052);
nor U7935 (N_7935,N_7354,N_7228);
and U7936 (N_7936,N_7049,N_7484);
and U7937 (N_7937,N_7168,N_7132);
and U7938 (N_7938,N_7034,N_7421);
or U7939 (N_7939,N_7066,N_7188);
or U7940 (N_7940,N_7045,N_7065);
nand U7941 (N_7941,N_7116,N_7158);
nand U7942 (N_7942,N_7015,N_7159);
nand U7943 (N_7943,N_7114,N_7245);
or U7944 (N_7944,N_7397,N_7261);
and U7945 (N_7945,N_7491,N_7079);
nor U7946 (N_7946,N_7045,N_7302);
and U7947 (N_7947,N_7198,N_7232);
nand U7948 (N_7948,N_7269,N_7209);
and U7949 (N_7949,N_7380,N_7319);
nor U7950 (N_7950,N_7472,N_7396);
or U7951 (N_7951,N_7401,N_7103);
and U7952 (N_7952,N_7419,N_7214);
nor U7953 (N_7953,N_7471,N_7301);
and U7954 (N_7954,N_7369,N_7364);
or U7955 (N_7955,N_7195,N_7183);
nand U7956 (N_7956,N_7427,N_7262);
or U7957 (N_7957,N_7020,N_7195);
or U7958 (N_7958,N_7335,N_7258);
nand U7959 (N_7959,N_7236,N_7031);
or U7960 (N_7960,N_7083,N_7189);
xnor U7961 (N_7961,N_7314,N_7018);
xnor U7962 (N_7962,N_7206,N_7329);
and U7963 (N_7963,N_7212,N_7439);
nor U7964 (N_7964,N_7001,N_7023);
and U7965 (N_7965,N_7353,N_7085);
nor U7966 (N_7966,N_7422,N_7098);
nand U7967 (N_7967,N_7330,N_7224);
and U7968 (N_7968,N_7133,N_7349);
and U7969 (N_7969,N_7417,N_7273);
or U7970 (N_7970,N_7013,N_7495);
nand U7971 (N_7971,N_7451,N_7364);
xor U7972 (N_7972,N_7329,N_7374);
nand U7973 (N_7973,N_7079,N_7011);
nand U7974 (N_7974,N_7047,N_7052);
xor U7975 (N_7975,N_7310,N_7207);
or U7976 (N_7976,N_7458,N_7271);
and U7977 (N_7977,N_7198,N_7083);
and U7978 (N_7978,N_7381,N_7373);
nand U7979 (N_7979,N_7206,N_7356);
xnor U7980 (N_7980,N_7483,N_7383);
nor U7981 (N_7981,N_7288,N_7494);
nor U7982 (N_7982,N_7023,N_7060);
xnor U7983 (N_7983,N_7112,N_7305);
nand U7984 (N_7984,N_7380,N_7378);
or U7985 (N_7985,N_7386,N_7308);
nor U7986 (N_7986,N_7097,N_7280);
or U7987 (N_7987,N_7062,N_7124);
nor U7988 (N_7988,N_7003,N_7194);
nand U7989 (N_7989,N_7435,N_7086);
or U7990 (N_7990,N_7292,N_7257);
and U7991 (N_7991,N_7495,N_7265);
nor U7992 (N_7992,N_7258,N_7273);
xor U7993 (N_7993,N_7424,N_7005);
and U7994 (N_7994,N_7128,N_7201);
or U7995 (N_7995,N_7028,N_7390);
or U7996 (N_7996,N_7082,N_7148);
and U7997 (N_7997,N_7215,N_7063);
and U7998 (N_7998,N_7248,N_7436);
and U7999 (N_7999,N_7203,N_7106);
nor U8000 (N_8000,N_7795,N_7802);
nand U8001 (N_8001,N_7805,N_7760);
xnor U8002 (N_8002,N_7680,N_7761);
nand U8003 (N_8003,N_7780,N_7875);
or U8004 (N_8004,N_7715,N_7579);
nor U8005 (N_8005,N_7984,N_7722);
or U8006 (N_8006,N_7697,N_7620);
nor U8007 (N_8007,N_7816,N_7595);
nor U8008 (N_8008,N_7848,N_7529);
nor U8009 (N_8009,N_7552,N_7725);
or U8010 (N_8010,N_7771,N_7922);
nor U8011 (N_8011,N_7979,N_7743);
and U8012 (N_8012,N_7941,N_7665);
xor U8013 (N_8013,N_7564,N_7531);
nor U8014 (N_8014,N_7877,N_7534);
and U8015 (N_8015,N_7924,N_7921);
nor U8016 (N_8016,N_7694,N_7658);
nand U8017 (N_8017,N_7840,N_7919);
xnor U8018 (N_8018,N_7939,N_7664);
nand U8019 (N_8019,N_7827,N_7583);
xnor U8020 (N_8020,N_7842,N_7963);
nand U8021 (N_8021,N_7754,N_7777);
and U8022 (N_8022,N_7522,N_7686);
nand U8023 (N_8023,N_7861,N_7774);
and U8024 (N_8024,N_7871,N_7618);
nor U8025 (N_8025,N_7560,N_7790);
or U8026 (N_8026,N_7784,N_7844);
and U8027 (N_8027,N_7513,N_7581);
or U8028 (N_8028,N_7850,N_7701);
nand U8029 (N_8029,N_7521,N_7544);
nand U8030 (N_8030,N_7575,N_7550);
nand U8031 (N_8031,N_7582,N_7956);
or U8032 (N_8032,N_7808,N_7500);
and U8033 (N_8033,N_7789,N_7806);
nor U8034 (N_8034,N_7590,N_7823);
or U8035 (N_8035,N_7703,N_7813);
and U8036 (N_8036,N_7587,N_7859);
nor U8037 (N_8037,N_7543,N_7990);
nand U8038 (N_8038,N_7609,N_7955);
nand U8039 (N_8039,N_7642,N_7764);
nor U8040 (N_8040,N_7762,N_7989);
and U8041 (N_8041,N_7535,N_7982);
nand U8042 (N_8042,N_7663,N_7885);
and U8043 (N_8043,N_7878,N_7737);
and U8044 (N_8044,N_7923,N_7863);
or U8045 (N_8045,N_7649,N_7501);
and U8046 (N_8046,N_7865,N_7699);
nor U8047 (N_8047,N_7613,N_7570);
and U8048 (N_8048,N_7781,N_7502);
or U8049 (N_8049,N_7638,N_7592);
nor U8050 (N_8050,N_7692,N_7948);
nor U8051 (N_8051,N_7893,N_7897);
xor U8052 (N_8052,N_7852,N_7600);
or U8053 (N_8053,N_7641,N_7997);
or U8054 (N_8054,N_7884,N_7942);
or U8055 (N_8055,N_7573,N_7549);
and U8056 (N_8056,N_7812,N_7576);
or U8057 (N_8057,N_7666,N_7698);
nor U8058 (N_8058,N_7545,N_7723);
or U8059 (N_8059,N_7801,N_7829);
or U8060 (N_8060,N_7630,N_7572);
and U8061 (N_8061,N_7696,N_7597);
or U8062 (N_8062,N_7974,N_7628);
nor U8063 (N_8063,N_7537,N_7970);
or U8064 (N_8064,N_7561,N_7750);
and U8065 (N_8065,N_7935,N_7504);
nor U8066 (N_8066,N_7695,N_7547);
and U8067 (N_8067,N_7569,N_7667);
nand U8068 (N_8068,N_7798,N_7831);
nor U8069 (N_8069,N_7817,N_7621);
and U8070 (N_8070,N_7846,N_7946);
nor U8071 (N_8071,N_7901,N_7839);
xor U8072 (N_8072,N_7684,N_7991);
nand U8073 (N_8073,N_7945,N_7660);
or U8074 (N_8074,N_7954,N_7902);
nand U8075 (N_8075,N_7994,N_7757);
and U8076 (N_8076,N_7913,N_7977);
or U8077 (N_8077,N_7718,N_7962);
xor U8078 (N_8078,N_7721,N_7756);
xnor U8079 (N_8079,N_7951,N_7766);
and U8080 (N_8080,N_7524,N_7765);
nor U8081 (N_8081,N_7662,N_7916);
nor U8082 (N_8082,N_7637,N_7972);
nor U8083 (N_8083,N_7510,N_7758);
nand U8084 (N_8084,N_7753,N_7625);
nand U8085 (N_8085,N_7707,N_7769);
and U8086 (N_8086,N_7627,N_7969);
nor U8087 (N_8087,N_7541,N_7571);
nor U8088 (N_8088,N_7659,N_7526);
or U8089 (N_8089,N_7964,N_7728);
nor U8090 (N_8090,N_7603,N_7584);
and U8091 (N_8091,N_7910,N_7953);
or U8092 (N_8092,N_7655,N_7735);
nand U8093 (N_8093,N_7746,N_7557);
or U8094 (N_8094,N_7824,N_7747);
xnor U8095 (N_8095,N_7578,N_7870);
and U8096 (N_8096,N_7588,N_7652);
and U8097 (N_8097,N_7906,N_7530);
and U8098 (N_8098,N_7710,N_7629);
and U8099 (N_8099,N_7983,N_7809);
nand U8100 (N_8100,N_7880,N_7882);
nand U8101 (N_8101,N_7751,N_7853);
and U8102 (N_8102,N_7708,N_7646);
nor U8103 (N_8103,N_7650,N_7937);
and U8104 (N_8104,N_7635,N_7594);
nor U8105 (N_8105,N_7611,N_7706);
or U8106 (N_8106,N_7999,N_7565);
and U8107 (N_8107,N_7726,N_7632);
or U8108 (N_8108,N_7793,N_7833);
nor U8109 (N_8109,N_7985,N_7838);
nand U8110 (N_8110,N_7682,N_7536);
nand U8111 (N_8111,N_7523,N_7810);
and U8112 (N_8112,N_7518,N_7860);
nand U8113 (N_8113,N_7626,N_7925);
or U8114 (N_8114,N_7717,N_7905);
and U8115 (N_8115,N_7516,N_7876);
and U8116 (N_8116,N_7834,N_7538);
nand U8117 (N_8117,N_7604,N_7678);
nor U8118 (N_8118,N_7558,N_7943);
nand U8119 (N_8119,N_7783,N_7792);
xor U8120 (N_8120,N_7929,N_7591);
nor U8121 (N_8121,N_7528,N_7505);
and U8122 (N_8122,N_7506,N_7546);
nor U8123 (N_8123,N_7748,N_7958);
or U8124 (N_8124,N_7837,N_7949);
and U8125 (N_8125,N_7616,N_7791);
nand U8126 (N_8126,N_7908,N_7532);
xnor U8127 (N_8127,N_7712,N_7787);
nor U8128 (N_8128,N_7596,N_7975);
or U8129 (N_8129,N_7744,N_7668);
nand U8130 (N_8130,N_7539,N_7976);
nor U8131 (N_8131,N_7700,N_7670);
nand U8132 (N_8132,N_7914,N_7836);
nor U8133 (N_8133,N_7845,N_7738);
nor U8134 (N_8134,N_7890,N_7868);
nor U8135 (N_8135,N_7966,N_7915);
or U8136 (N_8136,N_7992,N_7886);
nand U8137 (N_8137,N_7767,N_7740);
nand U8138 (N_8138,N_7759,N_7606);
nor U8139 (N_8139,N_7651,N_7887);
and U8140 (N_8140,N_7675,N_7912);
nand U8141 (N_8141,N_7927,N_7749);
nor U8142 (N_8142,N_7892,N_7851);
nand U8143 (N_8143,N_7517,N_7519);
and U8144 (N_8144,N_7731,N_7903);
or U8145 (N_8145,N_7857,N_7911);
nor U8146 (N_8146,N_7617,N_7959);
xor U8147 (N_8147,N_7803,N_7986);
xnor U8148 (N_8148,N_7574,N_7881);
nand U8149 (N_8149,N_7515,N_7896);
nand U8150 (N_8150,N_7830,N_7520);
nor U8151 (N_8151,N_7661,N_7981);
xnor U8152 (N_8152,N_7720,N_7729);
or U8153 (N_8153,N_7669,N_7601);
nor U8154 (N_8154,N_7685,N_7858);
nor U8155 (N_8155,N_7928,N_7512);
nor U8156 (N_8156,N_7580,N_7739);
or U8157 (N_8157,N_7704,N_7820);
nand U8158 (N_8158,N_7586,N_7688);
nand U8159 (N_8159,N_7826,N_7825);
nand U8160 (N_8160,N_7623,N_7671);
nand U8161 (N_8161,N_7770,N_7657);
nor U8162 (N_8162,N_7907,N_7568);
nor U8163 (N_8163,N_7788,N_7909);
nor U8164 (N_8164,N_7821,N_7622);
or U8165 (N_8165,N_7773,N_7818);
or U8166 (N_8166,N_7745,N_7730);
and U8167 (N_8167,N_7996,N_7593);
and U8168 (N_8168,N_7894,N_7973);
nand U8169 (N_8169,N_7794,N_7511);
nor U8170 (N_8170,N_7525,N_7509);
nor U8171 (N_8171,N_7719,N_7786);
nor U8172 (N_8172,N_7752,N_7567);
nor U8173 (N_8173,N_7653,N_7691);
and U8174 (N_8174,N_7679,N_7952);
nand U8175 (N_8175,N_7862,N_7640);
or U8176 (N_8176,N_7644,N_7527);
nor U8177 (N_8177,N_7940,N_7867);
and U8178 (N_8178,N_7555,N_7856);
nor U8179 (N_8179,N_7828,N_7961);
nor U8180 (N_8180,N_7874,N_7947);
nor U8181 (N_8181,N_7807,N_7957);
and U8182 (N_8182,N_7614,N_7503);
and U8183 (N_8183,N_7768,N_7672);
or U8184 (N_8184,N_7674,N_7796);
nand U8185 (N_8185,N_7702,N_7847);
and U8186 (N_8186,N_7605,N_7800);
or U8187 (N_8187,N_7782,N_7639);
nand U8188 (N_8188,N_7732,N_7944);
nand U8189 (N_8189,N_7811,N_7960);
nand U8190 (N_8190,N_7514,N_7869);
nor U8191 (N_8191,N_7677,N_7734);
and U8192 (N_8192,N_7736,N_7864);
nor U8193 (N_8193,N_7995,N_7899);
nor U8194 (N_8194,N_7742,N_7636);
or U8195 (N_8195,N_7920,N_7714);
xor U8196 (N_8196,N_7683,N_7879);
nand U8197 (N_8197,N_7648,N_7785);
nand U8198 (N_8198,N_7553,N_7602);
xnor U8199 (N_8199,N_7705,N_7673);
and U8200 (N_8200,N_7873,N_7633);
and U8201 (N_8201,N_7676,N_7619);
nand U8202 (N_8202,N_7610,N_7612);
nand U8203 (N_8203,N_7938,N_7693);
nand U8204 (N_8204,N_7533,N_7711);
nand U8205 (N_8205,N_7993,N_7799);
nand U8206 (N_8206,N_7936,N_7888);
nand U8207 (N_8207,N_7724,N_7763);
nand U8208 (N_8208,N_7548,N_7577);
or U8209 (N_8209,N_7904,N_7647);
nand U8210 (N_8210,N_7971,N_7608);
and U8211 (N_8211,N_7741,N_7634);
or U8212 (N_8212,N_7926,N_7713);
nand U8213 (N_8213,N_7566,N_7716);
and U8214 (N_8214,N_7540,N_7654);
or U8215 (N_8215,N_7814,N_7689);
and U8216 (N_8216,N_7559,N_7934);
and U8217 (N_8217,N_7930,N_7562);
or U8218 (N_8218,N_7855,N_7508);
nand U8219 (N_8219,N_7835,N_7866);
nand U8220 (N_8220,N_7598,N_7822);
nand U8221 (N_8221,N_7932,N_7987);
nor U8222 (N_8222,N_7776,N_7883);
or U8223 (N_8223,N_7656,N_7554);
nor U8224 (N_8224,N_7933,N_7778);
nor U8225 (N_8225,N_7727,N_7819);
nor U8226 (N_8226,N_7690,N_7563);
and U8227 (N_8227,N_7551,N_7931);
and U8228 (N_8228,N_7950,N_7980);
or U8229 (N_8229,N_7804,N_7815);
nor U8230 (N_8230,N_7542,N_7978);
nor U8231 (N_8231,N_7854,N_7585);
and U8232 (N_8232,N_7733,N_7615);
and U8233 (N_8233,N_7917,N_7841);
and U8234 (N_8234,N_7589,N_7898);
nand U8235 (N_8235,N_7643,N_7889);
nor U8236 (N_8236,N_7843,N_7988);
xnor U8237 (N_8237,N_7832,N_7687);
and U8238 (N_8238,N_7507,N_7556);
or U8239 (N_8239,N_7681,N_7631);
nor U8240 (N_8240,N_7709,N_7965);
nand U8241 (N_8241,N_7998,N_7891);
and U8242 (N_8242,N_7607,N_7968);
nand U8243 (N_8243,N_7872,N_7918);
xnor U8244 (N_8244,N_7849,N_7775);
nor U8245 (N_8245,N_7900,N_7599);
nor U8246 (N_8246,N_7779,N_7755);
nand U8247 (N_8247,N_7797,N_7772);
or U8248 (N_8248,N_7645,N_7895);
and U8249 (N_8249,N_7967,N_7624);
or U8250 (N_8250,N_7507,N_7670);
xor U8251 (N_8251,N_7825,N_7820);
or U8252 (N_8252,N_7728,N_7755);
nand U8253 (N_8253,N_7501,N_7995);
or U8254 (N_8254,N_7995,N_7839);
nand U8255 (N_8255,N_7567,N_7888);
nand U8256 (N_8256,N_7785,N_7920);
or U8257 (N_8257,N_7714,N_7597);
nor U8258 (N_8258,N_7796,N_7795);
nor U8259 (N_8259,N_7641,N_7961);
nand U8260 (N_8260,N_7915,N_7904);
nand U8261 (N_8261,N_7753,N_7876);
or U8262 (N_8262,N_7758,N_7763);
or U8263 (N_8263,N_7844,N_7883);
nor U8264 (N_8264,N_7685,N_7895);
nor U8265 (N_8265,N_7979,N_7620);
and U8266 (N_8266,N_7570,N_7611);
nor U8267 (N_8267,N_7793,N_7750);
and U8268 (N_8268,N_7943,N_7575);
nor U8269 (N_8269,N_7825,N_7659);
nor U8270 (N_8270,N_7620,N_7975);
and U8271 (N_8271,N_7641,N_7965);
nor U8272 (N_8272,N_7702,N_7647);
xnor U8273 (N_8273,N_7950,N_7869);
nor U8274 (N_8274,N_7508,N_7572);
or U8275 (N_8275,N_7922,N_7559);
nand U8276 (N_8276,N_7703,N_7804);
or U8277 (N_8277,N_7832,N_7874);
xor U8278 (N_8278,N_7831,N_7962);
and U8279 (N_8279,N_7753,N_7825);
and U8280 (N_8280,N_7987,N_7806);
nand U8281 (N_8281,N_7637,N_7857);
and U8282 (N_8282,N_7987,N_7619);
xnor U8283 (N_8283,N_7858,N_7862);
and U8284 (N_8284,N_7602,N_7786);
nor U8285 (N_8285,N_7553,N_7544);
nor U8286 (N_8286,N_7520,N_7920);
nor U8287 (N_8287,N_7777,N_7697);
or U8288 (N_8288,N_7648,N_7970);
nor U8289 (N_8289,N_7670,N_7748);
or U8290 (N_8290,N_7962,N_7753);
or U8291 (N_8291,N_7758,N_7524);
nor U8292 (N_8292,N_7948,N_7725);
and U8293 (N_8293,N_7877,N_7602);
nor U8294 (N_8294,N_7778,N_7861);
and U8295 (N_8295,N_7621,N_7770);
nor U8296 (N_8296,N_7890,N_7847);
nor U8297 (N_8297,N_7764,N_7635);
and U8298 (N_8298,N_7521,N_7627);
and U8299 (N_8299,N_7969,N_7978);
or U8300 (N_8300,N_7923,N_7767);
or U8301 (N_8301,N_7877,N_7981);
nor U8302 (N_8302,N_7937,N_7972);
nor U8303 (N_8303,N_7685,N_7860);
and U8304 (N_8304,N_7758,N_7992);
nand U8305 (N_8305,N_7846,N_7896);
or U8306 (N_8306,N_7711,N_7689);
nand U8307 (N_8307,N_7773,N_7610);
nor U8308 (N_8308,N_7735,N_7536);
and U8309 (N_8309,N_7694,N_7852);
and U8310 (N_8310,N_7548,N_7598);
or U8311 (N_8311,N_7925,N_7773);
or U8312 (N_8312,N_7624,N_7752);
nor U8313 (N_8313,N_7506,N_7526);
nand U8314 (N_8314,N_7848,N_7516);
xor U8315 (N_8315,N_7820,N_7545);
nor U8316 (N_8316,N_7907,N_7676);
and U8317 (N_8317,N_7943,N_7503);
or U8318 (N_8318,N_7702,N_7594);
xor U8319 (N_8319,N_7711,N_7790);
nor U8320 (N_8320,N_7532,N_7795);
nor U8321 (N_8321,N_7922,N_7623);
and U8322 (N_8322,N_7729,N_7838);
or U8323 (N_8323,N_7843,N_7635);
xnor U8324 (N_8324,N_7528,N_7720);
xor U8325 (N_8325,N_7967,N_7778);
xnor U8326 (N_8326,N_7893,N_7721);
or U8327 (N_8327,N_7878,N_7856);
and U8328 (N_8328,N_7652,N_7959);
or U8329 (N_8329,N_7695,N_7958);
and U8330 (N_8330,N_7719,N_7762);
or U8331 (N_8331,N_7784,N_7691);
and U8332 (N_8332,N_7570,N_7582);
nand U8333 (N_8333,N_7552,N_7889);
nand U8334 (N_8334,N_7960,N_7552);
xor U8335 (N_8335,N_7609,N_7611);
and U8336 (N_8336,N_7969,N_7595);
nor U8337 (N_8337,N_7512,N_7865);
or U8338 (N_8338,N_7559,N_7585);
xor U8339 (N_8339,N_7933,N_7807);
and U8340 (N_8340,N_7964,N_7947);
and U8341 (N_8341,N_7950,N_7564);
and U8342 (N_8342,N_7971,N_7559);
or U8343 (N_8343,N_7616,N_7882);
and U8344 (N_8344,N_7620,N_7886);
or U8345 (N_8345,N_7553,N_7624);
and U8346 (N_8346,N_7579,N_7530);
nand U8347 (N_8347,N_7520,N_7956);
nand U8348 (N_8348,N_7973,N_7590);
and U8349 (N_8349,N_7645,N_7677);
nor U8350 (N_8350,N_7670,N_7826);
nand U8351 (N_8351,N_7674,N_7973);
and U8352 (N_8352,N_7890,N_7787);
nand U8353 (N_8353,N_7935,N_7870);
or U8354 (N_8354,N_7705,N_7763);
nor U8355 (N_8355,N_7603,N_7555);
xnor U8356 (N_8356,N_7841,N_7613);
or U8357 (N_8357,N_7602,N_7639);
nor U8358 (N_8358,N_7988,N_7500);
xnor U8359 (N_8359,N_7767,N_7863);
nand U8360 (N_8360,N_7904,N_7940);
xor U8361 (N_8361,N_7796,N_7801);
or U8362 (N_8362,N_7732,N_7968);
nand U8363 (N_8363,N_7872,N_7738);
or U8364 (N_8364,N_7596,N_7898);
nor U8365 (N_8365,N_7558,N_7555);
and U8366 (N_8366,N_7569,N_7561);
and U8367 (N_8367,N_7802,N_7547);
nor U8368 (N_8368,N_7728,N_7848);
and U8369 (N_8369,N_7772,N_7625);
or U8370 (N_8370,N_7730,N_7835);
xnor U8371 (N_8371,N_7725,N_7899);
xnor U8372 (N_8372,N_7817,N_7703);
and U8373 (N_8373,N_7799,N_7711);
xnor U8374 (N_8374,N_7687,N_7669);
nor U8375 (N_8375,N_7769,N_7722);
nand U8376 (N_8376,N_7975,N_7549);
nand U8377 (N_8377,N_7609,N_7514);
and U8378 (N_8378,N_7845,N_7939);
and U8379 (N_8379,N_7536,N_7520);
xnor U8380 (N_8380,N_7759,N_7893);
nand U8381 (N_8381,N_7508,N_7835);
or U8382 (N_8382,N_7711,N_7517);
nand U8383 (N_8383,N_7978,N_7592);
nand U8384 (N_8384,N_7715,N_7765);
and U8385 (N_8385,N_7577,N_7683);
nand U8386 (N_8386,N_7572,N_7626);
or U8387 (N_8387,N_7708,N_7586);
xnor U8388 (N_8388,N_7551,N_7764);
nand U8389 (N_8389,N_7506,N_7823);
and U8390 (N_8390,N_7578,N_7853);
nand U8391 (N_8391,N_7865,N_7983);
nand U8392 (N_8392,N_7947,N_7660);
and U8393 (N_8393,N_7598,N_7608);
nor U8394 (N_8394,N_7970,N_7544);
or U8395 (N_8395,N_7892,N_7939);
nor U8396 (N_8396,N_7810,N_7637);
nand U8397 (N_8397,N_7568,N_7844);
and U8398 (N_8398,N_7947,N_7532);
nand U8399 (N_8399,N_7916,N_7925);
or U8400 (N_8400,N_7911,N_7837);
nand U8401 (N_8401,N_7566,N_7811);
and U8402 (N_8402,N_7807,N_7683);
or U8403 (N_8403,N_7531,N_7635);
and U8404 (N_8404,N_7929,N_7695);
and U8405 (N_8405,N_7662,N_7590);
and U8406 (N_8406,N_7626,N_7950);
xor U8407 (N_8407,N_7813,N_7665);
nand U8408 (N_8408,N_7618,N_7659);
and U8409 (N_8409,N_7530,N_7822);
or U8410 (N_8410,N_7756,N_7667);
nor U8411 (N_8411,N_7708,N_7982);
nand U8412 (N_8412,N_7755,N_7647);
nor U8413 (N_8413,N_7584,N_7515);
nor U8414 (N_8414,N_7562,N_7815);
and U8415 (N_8415,N_7612,N_7543);
nor U8416 (N_8416,N_7599,N_7645);
and U8417 (N_8417,N_7654,N_7945);
and U8418 (N_8418,N_7807,N_7863);
nor U8419 (N_8419,N_7601,N_7856);
nor U8420 (N_8420,N_7783,N_7836);
and U8421 (N_8421,N_7977,N_7538);
nand U8422 (N_8422,N_7946,N_7869);
or U8423 (N_8423,N_7813,N_7636);
nor U8424 (N_8424,N_7729,N_7862);
or U8425 (N_8425,N_7545,N_7543);
and U8426 (N_8426,N_7824,N_7808);
nand U8427 (N_8427,N_7786,N_7566);
and U8428 (N_8428,N_7988,N_7852);
and U8429 (N_8429,N_7607,N_7643);
nor U8430 (N_8430,N_7877,N_7626);
and U8431 (N_8431,N_7874,N_7677);
nor U8432 (N_8432,N_7982,N_7636);
or U8433 (N_8433,N_7613,N_7731);
and U8434 (N_8434,N_7765,N_7876);
and U8435 (N_8435,N_7524,N_7684);
nor U8436 (N_8436,N_7784,N_7901);
or U8437 (N_8437,N_7921,N_7685);
nand U8438 (N_8438,N_7586,N_7850);
or U8439 (N_8439,N_7811,N_7910);
and U8440 (N_8440,N_7675,N_7663);
or U8441 (N_8441,N_7704,N_7683);
and U8442 (N_8442,N_7817,N_7665);
or U8443 (N_8443,N_7993,N_7800);
and U8444 (N_8444,N_7567,N_7754);
and U8445 (N_8445,N_7572,N_7677);
nand U8446 (N_8446,N_7763,N_7928);
xor U8447 (N_8447,N_7627,N_7736);
xor U8448 (N_8448,N_7832,N_7794);
and U8449 (N_8449,N_7742,N_7819);
nand U8450 (N_8450,N_7745,N_7898);
or U8451 (N_8451,N_7581,N_7526);
nand U8452 (N_8452,N_7894,N_7722);
and U8453 (N_8453,N_7538,N_7530);
and U8454 (N_8454,N_7655,N_7516);
or U8455 (N_8455,N_7772,N_7553);
and U8456 (N_8456,N_7934,N_7906);
and U8457 (N_8457,N_7918,N_7572);
nand U8458 (N_8458,N_7593,N_7994);
nor U8459 (N_8459,N_7530,N_7625);
nand U8460 (N_8460,N_7503,N_7901);
and U8461 (N_8461,N_7989,N_7530);
or U8462 (N_8462,N_7930,N_7617);
xnor U8463 (N_8463,N_7682,N_7532);
nor U8464 (N_8464,N_7887,N_7850);
nor U8465 (N_8465,N_7847,N_7618);
or U8466 (N_8466,N_7787,N_7672);
or U8467 (N_8467,N_7888,N_7780);
nand U8468 (N_8468,N_7991,N_7625);
nor U8469 (N_8469,N_7941,N_7979);
nor U8470 (N_8470,N_7678,N_7725);
and U8471 (N_8471,N_7572,N_7929);
or U8472 (N_8472,N_7812,N_7843);
nor U8473 (N_8473,N_7746,N_7982);
nand U8474 (N_8474,N_7586,N_7589);
nor U8475 (N_8475,N_7514,N_7912);
nor U8476 (N_8476,N_7703,N_7848);
and U8477 (N_8477,N_7587,N_7960);
xnor U8478 (N_8478,N_7966,N_7756);
nand U8479 (N_8479,N_7656,N_7542);
and U8480 (N_8480,N_7890,N_7691);
and U8481 (N_8481,N_7844,N_7525);
and U8482 (N_8482,N_7837,N_7548);
nor U8483 (N_8483,N_7915,N_7630);
or U8484 (N_8484,N_7769,N_7515);
xor U8485 (N_8485,N_7673,N_7550);
xor U8486 (N_8486,N_7775,N_7733);
xnor U8487 (N_8487,N_7868,N_7760);
nand U8488 (N_8488,N_7792,N_7751);
xor U8489 (N_8489,N_7911,N_7827);
xnor U8490 (N_8490,N_7681,N_7649);
nand U8491 (N_8491,N_7901,N_7881);
xor U8492 (N_8492,N_7762,N_7699);
nand U8493 (N_8493,N_7669,N_7788);
xnor U8494 (N_8494,N_7892,N_7563);
and U8495 (N_8495,N_7566,N_7748);
nand U8496 (N_8496,N_7730,N_7573);
or U8497 (N_8497,N_7871,N_7959);
and U8498 (N_8498,N_7791,N_7533);
nor U8499 (N_8499,N_7932,N_7858);
nor U8500 (N_8500,N_8111,N_8048);
and U8501 (N_8501,N_8152,N_8150);
nand U8502 (N_8502,N_8387,N_8346);
xor U8503 (N_8503,N_8383,N_8463);
nor U8504 (N_8504,N_8247,N_8487);
or U8505 (N_8505,N_8361,N_8412);
or U8506 (N_8506,N_8453,N_8477);
and U8507 (N_8507,N_8068,N_8351);
or U8508 (N_8508,N_8241,N_8015);
nand U8509 (N_8509,N_8297,N_8332);
nand U8510 (N_8510,N_8102,N_8126);
or U8511 (N_8511,N_8400,N_8275);
or U8512 (N_8512,N_8234,N_8061);
nand U8513 (N_8513,N_8416,N_8450);
or U8514 (N_8514,N_8017,N_8146);
xnor U8515 (N_8515,N_8331,N_8401);
xnor U8516 (N_8516,N_8004,N_8348);
nor U8517 (N_8517,N_8024,N_8273);
or U8518 (N_8518,N_8343,N_8433);
nand U8519 (N_8519,N_8135,N_8447);
or U8520 (N_8520,N_8438,N_8046);
or U8521 (N_8521,N_8472,N_8100);
xor U8522 (N_8522,N_8426,N_8060);
and U8523 (N_8523,N_8404,N_8417);
nand U8524 (N_8524,N_8018,N_8466);
nand U8525 (N_8525,N_8442,N_8141);
xnor U8526 (N_8526,N_8082,N_8054);
nand U8527 (N_8527,N_8190,N_8036);
or U8528 (N_8528,N_8071,N_8057);
nor U8529 (N_8529,N_8213,N_8446);
nand U8530 (N_8530,N_8373,N_8195);
nor U8531 (N_8531,N_8254,N_8339);
or U8532 (N_8532,N_8083,N_8357);
and U8533 (N_8533,N_8076,N_8075);
or U8534 (N_8534,N_8281,N_8073);
and U8535 (N_8535,N_8178,N_8115);
nand U8536 (N_8536,N_8283,N_8497);
and U8537 (N_8537,N_8316,N_8043);
nor U8538 (N_8538,N_8486,N_8144);
nand U8539 (N_8539,N_8238,N_8008);
or U8540 (N_8540,N_8455,N_8007);
nand U8541 (N_8541,N_8268,N_8395);
nor U8542 (N_8542,N_8451,N_8299);
xor U8543 (N_8543,N_8366,N_8174);
or U8544 (N_8544,N_8489,N_8130);
nand U8545 (N_8545,N_8110,N_8271);
xnor U8546 (N_8546,N_8494,N_8199);
nand U8547 (N_8547,N_8267,N_8379);
nor U8548 (N_8548,N_8272,N_8037);
and U8549 (N_8549,N_8137,N_8293);
or U8550 (N_8550,N_8176,N_8208);
and U8551 (N_8551,N_8369,N_8325);
or U8552 (N_8552,N_8367,N_8164);
or U8553 (N_8553,N_8127,N_8385);
and U8554 (N_8554,N_8246,N_8171);
or U8555 (N_8555,N_8006,N_8388);
nor U8556 (N_8556,N_8231,N_8291);
or U8557 (N_8557,N_8315,N_8403);
or U8558 (N_8558,N_8354,N_8156);
nand U8559 (N_8559,N_8044,N_8448);
nor U8560 (N_8560,N_8058,N_8147);
or U8561 (N_8561,N_8397,N_8239);
and U8562 (N_8562,N_8481,N_8311);
and U8563 (N_8563,N_8028,N_8264);
and U8564 (N_8564,N_8490,N_8408);
or U8565 (N_8565,N_8209,N_8023);
xnor U8566 (N_8566,N_8131,N_8122);
nand U8567 (N_8567,N_8217,N_8488);
nor U8568 (N_8568,N_8118,N_8347);
and U8569 (N_8569,N_8358,N_8079);
nor U8570 (N_8570,N_8025,N_8149);
nand U8571 (N_8571,N_8396,N_8159);
or U8572 (N_8572,N_8476,N_8183);
nand U8573 (N_8573,N_8419,N_8435);
and U8574 (N_8574,N_8139,N_8405);
nand U8575 (N_8575,N_8329,N_8313);
nand U8576 (N_8576,N_8406,N_8035);
nor U8577 (N_8577,N_8207,N_8375);
nand U8578 (N_8578,N_8320,N_8390);
nand U8579 (N_8579,N_8233,N_8189);
nor U8580 (N_8580,N_8296,N_8413);
nand U8581 (N_8581,N_8386,N_8012);
nand U8582 (N_8582,N_8422,N_8096);
nand U8583 (N_8583,N_8177,N_8250);
nand U8584 (N_8584,N_8077,N_8399);
nand U8585 (N_8585,N_8362,N_8491);
nand U8586 (N_8586,N_8289,N_8312);
xnor U8587 (N_8587,N_8232,N_8132);
and U8588 (N_8588,N_8045,N_8444);
nand U8589 (N_8589,N_8010,N_8140);
or U8590 (N_8590,N_8244,N_8112);
nand U8591 (N_8591,N_8256,N_8407);
nand U8592 (N_8592,N_8452,N_8454);
and U8593 (N_8593,N_8474,N_8050);
or U8594 (N_8594,N_8302,N_8108);
xnor U8595 (N_8595,N_8087,N_8393);
or U8596 (N_8596,N_8355,N_8066);
xnor U8597 (N_8597,N_8310,N_8214);
nor U8598 (N_8598,N_8070,N_8245);
nand U8599 (N_8599,N_8294,N_8031);
nor U8600 (N_8600,N_8216,N_8371);
or U8601 (N_8601,N_8047,N_8240);
and U8602 (N_8602,N_8099,N_8278);
nor U8603 (N_8603,N_8052,N_8356);
or U8604 (N_8604,N_8182,N_8274);
nand U8605 (N_8605,N_8445,N_8142);
and U8606 (N_8606,N_8298,N_8372);
and U8607 (N_8607,N_8163,N_8097);
nor U8608 (N_8608,N_8465,N_8078);
nor U8609 (N_8609,N_8205,N_8212);
nand U8610 (N_8610,N_8143,N_8319);
and U8611 (N_8611,N_8324,N_8220);
and U8612 (N_8612,N_8252,N_8039);
xor U8613 (N_8613,N_8340,N_8105);
nand U8614 (N_8614,N_8262,N_8352);
or U8615 (N_8615,N_8308,N_8022);
or U8616 (N_8616,N_8038,N_8185);
nand U8617 (N_8617,N_8288,N_8049);
nand U8618 (N_8618,N_8218,N_8376);
xnor U8619 (N_8619,N_8193,N_8215);
or U8620 (N_8620,N_8330,N_8114);
xnor U8621 (N_8621,N_8074,N_8456);
or U8622 (N_8622,N_8377,N_8468);
or U8623 (N_8623,N_8327,N_8430);
or U8624 (N_8624,N_8206,N_8225);
or U8625 (N_8625,N_8493,N_8424);
and U8626 (N_8626,N_8235,N_8287);
and U8627 (N_8627,N_8423,N_8086);
nand U8628 (N_8628,N_8187,N_8072);
and U8629 (N_8629,N_8248,N_8344);
and U8630 (N_8630,N_8001,N_8421);
nor U8631 (N_8631,N_8080,N_8107);
or U8632 (N_8632,N_8261,N_8398);
and U8633 (N_8633,N_8151,N_8365);
or U8634 (N_8634,N_8227,N_8479);
and U8635 (N_8635,N_8485,N_8276);
nand U8636 (N_8636,N_8336,N_8145);
or U8637 (N_8637,N_8418,N_8063);
and U8638 (N_8638,N_8134,N_8350);
xor U8639 (N_8639,N_8415,N_8034);
or U8640 (N_8640,N_8085,N_8186);
and U8641 (N_8641,N_8155,N_8251);
or U8642 (N_8642,N_8236,N_8067);
nor U8643 (N_8643,N_8095,N_8170);
nand U8644 (N_8644,N_8211,N_8381);
or U8645 (N_8645,N_8116,N_8284);
xnor U8646 (N_8646,N_8290,N_8253);
or U8647 (N_8647,N_8224,N_8295);
nand U8648 (N_8648,N_8103,N_8380);
nand U8649 (N_8649,N_8084,N_8370);
or U8650 (N_8650,N_8042,N_8098);
nor U8651 (N_8651,N_8196,N_8053);
and U8652 (N_8652,N_8201,N_8374);
or U8653 (N_8653,N_8266,N_8249);
nor U8654 (N_8654,N_8104,N_8305);
or U8655 (N_8655,N_8409,N_8228);
and U8656 (N_8656,N_8243,N_8337);
and U8657 (N_8657,N_8011,N_8129);
and U8658 (N_8658,N_8014,N_8016);
and U8659 (N_8659,N_8138,N_8414);
nor U8660 (N_8660,N_8326,N_8166);
or U8661 (N_8661,N_8003,N_8167);
nand U8662 (N_8662,N_8427,N_8482);
or U8663 (N_8663,N_8161,N_8285);
and U8664 (N_8664,N_8384,N_8342);
nor U8665 (N_8665,N_8119,N_8237);
nand U8666 (N_8666,N_8184,N_8286);
nand U8667 (N_8667,N_8292,N_8338);
and U8668 (N_8668,N_8005,N_8410);
nor U8669 (N_8669,N_8148,N_8255);
nand U8670 (N_8670,N_8030,N_8484);
and U8671 (N_8671,N_8202,N_8203);
nand U8672 (N_8672,N_8317,N_8194);
nand U8673 (N_8673,N_8306,N_8436);
nor U8674 (N_8674,N_8334,N_8349);
nand U8675 (N_8675,N_8172,N_8179);
or U8676 (N_8676,N_8360,N_8458);
nor U8677 (N_8677,N_8439,N_8429);
and U8678 (N_8678,N_8021,N_8259);
nor U8679 (N_8679,N_8402,N_8242);
or U8680 (N_8680,N_8335,N_8062);
xor U8681 (N_8681,N_8469,N_8420);
nand U8682 (N_8682,N_8318,N_8258);
nor U8683 (N_8683,N_8425,N_8160);
and U8684 (N_8684,N_8040,N_8389);
and U8685 (N_8685,N_8106,N_8345);
nand U8686 (N_8686,N_8260,N_8314);
nor U8687 (N_8687,N_8133,N_8475);
and U8688 (N_8688,N_8091,N_8434);
nor U8689 (N_8689,N_8392,N_8162);
nor U8690 (N_8690,N_8443,N_8013);
nor U8691 (N_8691,N_8059,N_8492);
and U8692 (N_8692,N_8191,N_8480);
xnor U8693 (N_8693,N_8301,N_8483);
and U8694 (N_8694,N_8221,N_8307);
nor U8695 (N_8695,N_8180,N_8464);
nor U8696 (N_8696,N_8265,N_8432);
nor U8697 (N_8697,N_8257,N_8027);
or U8698 (N_8698,N_8158,N_8363);
and U8699 (N_8699,N_8473,N_8065);
and U8700 (N_8700,N_8200,N_8069);
and U8701 (N_8701,N_8229,N_8328);
nor U8702 (N_8702,N_8223,N_8300);
nand U8703 (N_8703,N_8101,N_8009);
nand U8704 (N_8704,N_8188,N_8128);
nor U8705 (N_8705,N_8333,N_8173);
xnor U8706 (N_8706,N_8113,N_8136);
nand U8707 (N_8707,N_8081,N_8032);
nand U8708 (N_8708,N_8391,N_8124);
and U8709 (N_8709,N_8120,N_8341);
or U8710 (N_8710,N_8090,N_8304);
or U8711 (N_8711,N_8020,N_8051);
nor U8712 (N_8712,N_8041,N_8175);
and U8713 (N_8713,N_8382,N_8092);
and U8714 (N_8714,N_8368,N_8002);
xor U8715 (N_8715,N_8165,N_8210);
nand U8716 (N_8716,N_8033,N_8323);
and U8717 (N_8717,N_8093,N_8449);
nor U8718 (N_8718,N_8280,N_8263);
or U8719 (N_8719,N_8198,N_8026);
and U8720 (N_8720,N_8322,N_8496);
or U8721 (N_8721,N_8204,N_8309);
nor U8722 (N_8722,N_8498,N_8055);
or U8723 (N_8723,N_8378,N_8168);
xor U8724 (N_8724,N_8471,N_8279);
and U8725 (N_8725,N_8121,N_8094);
and U8726 (N_8726,N_8499,N_8181);
and U8727 (N_8727,N_8029,N_8467);
xnor U8728 (N_8728,N_8394,N_8462);
or U8729 (N_8729,N_8460,N_8123);
nor U8730 (N_8730,N_8230,N_8440);
or U8731 (N_8731,N_8282,N_8364);
or U8732 (N_8732,N_8169,N_8321);
nor U8733 (N_8733,N_8117,N_8109);
or U8734 (N_8734,N_8461,N_8064);
nor U8735 (N_8735,N_8157,N_8478);
nor U8736 (N_8736,N_8411,N_8437);
nand U8737 (N_8737,N_8000,N_8056);
and U8738 (N_8738,N_8470,N_8222);
nor U8739 (N_8739,N_8353,N_8192);
and U8740 (N_8740,N_8431,N_8088);
nand U8741 (N_8741,N_8457,N_8428);
or U8742 (N_8742,N_8459,N_8441);
or U8743 (N_8743,N_8270,N_8495);
or U8744 (N_8744,N_8153,N_8303);
or U8745 (N_8745,N_8089,N_8219);
and U8746 (N_8746,N_8277,N_8125);
nor U8747 (N_8747,N_8359,N_8154);
and U8748 (N_8748,N_8226,N_8019);
or U8749 (N_8749,N_8197,N_8269);
or U8750 (N_8750,N_8115,N_8274);
nand U8751 (N_8751,N_8309,N_8050);
or U8752 (N_8752,N_8321,N_8409);
nand U8753 (N_8753,N_8362,N_8133);
or U8754 (N_8754,N_8244,N_8260);
and U8755 (N_8755,N_8421,N_8193);
nand U8756 (N_8756,N_8083,N_8113);
and U8757 (N_8757,N_8286,N_8153);
nand U8758 (N_8758,N_8043,N_8426);
and U8759 (N_8759,N_8034,N_8106);
nand U8760 (N_8760,N_8395,N_8481);
and U8761 (N_8761,N_8330,N_8243);
and U8762 (N_8762,N_8120,N_8289);
nand U8763 (N_8763,N_8323,N_8040);
nor U8764 (N_8764,N_8437,N_8484);
nor U8765 (N_8765,N_8324,N_8051);
or U8766 (N_8766,N_8455,N_8219);
nand U8767 (N_8767,N_8333,N_8268);
or U8768 (N_8768,N_8176,N_8229);
or U8769 (N_8769,N_8360,N_8063);
and U8770 (N_8770,N_8405,N_8185);
nand U8771 (N_8771,N_8182,N_8005);
nor U8772 (N_8772,N_8350,N_8053);
or U8773 (N_8773,N_8370,N_8310);
nor U8774 (N_8774,N_8345,N_8247);
nand U8775 (N_8775,N_8072,N_8066);
and U8776 (N_8776,N_8289,N_8334);
or U8777 (N_8777,N_8185,N_8466);
and U8778 (N_8778,N_8455,N_8480);
nor U8779 (N_8779,N_8234,N_8397);
or U8780 (N_8780,N_8327,N_8337);
or U8781 (N_8781,N_8255,N_8398);
nand U8782 (N_8782,N_8172,N_8181);
nor U8783 (N_8783,N_8249,N_8248);
or U8784 (N_8784,N_8087,N_8221);
and U8785 (N_8785,N_8279,N_8428);
or U8786 (N_8786,N_8453,N_8022);
and U8787 (N_8787,N_8273,N_8351);
xnor U8788 (N_8788,N_8391,N_8202);
nand U8789 (N_8789,N_8439,N_8361);
nand U8790 (N_8790,N_8044,N_8308);
or U8791 (N_8791,N_8299,N_8003);
and U8792 (N_8792,N_8124,N_8192);
xor U8793 (N_8793,N_8440,N_8199);
nor U8794 (N_8794,N_8464,N_8038);
or U8795 (N_8795,N_8465,N_8362);
or U8796 (N_8796,N_8477,N_8141);
nor U8797 (N_8797,N_8060,N_8054);
xor U8798 (N_8798,N_8085,N_8038);
and U8799 (N_8799,N_8228,N_8242);
xnor U8800 (N_8800,N_8449,N_8435);
nor U8801 (N_8801,N_8498,N_8191);
nand U8802 (N_8802,N_8374,N_8129);
and U8803 (N_8803,N_8258,N_8162);
nor U8804 (N_8804,N_8481,N_8207);
or U8805 (N_8805,N_8320,N_8183);
and U8806 (N_8806,N_8342,N_8041);
nand U8807 (N_8807,N_8450,N_8156);
nor U8808 (N_8808,N_8318,N_8169);
nand U8809 (N_8809,N_8313,N_8218);
nor U8810 (N_8810,N_8171,N_8401);
xor U8811 (N_8811,N_8458,N_8182);
nor U8812 (N_8812,N_8246,N_8286);
xnor U8813 (N_8813,N_8465,N_8476);
and U8814 (N_8814,N_8403,N_8444);
nor U8815 (N_8815,N_8025,N_8401);
nand U8816 (N_8816,N_8253,N_8411);
nor U8817 (N_8817,N_8125,N_8245);
and U8818 (N_8818,N_8052,N_8363);
and U8819 (N_8819,N_8290,N_8476);
nand U8820 (N_8820,N_8117,N_8143);
nand U8821 (N_8821,N_8251,N_8338);
and U8822 (N_8822,N_8344,N_8075);
nor U8823 (N_8823,N_8020,N_8148);
and U8824 (N_8824,N_8360,N_8330);
and U8825 (N_8825,N_8150,N_8196);
or U8826 (N_8826,N_8318,N_8495);
or U8827 (N_8827,N_8149,N_8398);
nand U8828 (N_8828,N_8488,N_8440);
nor U8829 (N_8829,N_8433,N_8277);
nor U8830 (N_8830,N_8419,N_8432);
or U8831 (N_8831,N_8135,N_8094);
nand U8832 (N_8832,N_8429,N_8303);
nor U8833 (N_8833,N_8310,N_8359);
nand U8834 (N_8834,N_8046,N_8417);
or U8835 (N_8835,N_8187,N_8382);
and U8836 (N_8836,N_8488,N_8439);
and U8837 (N_8837,N_8060,N_8084);
nand U8838 (N_8838,N_8043,N_8065);
nand U8839 (N_8839,N_8332,N_8489);
nand U8840 (N_8840,N_8105,N_8422);
and U8841 (N_8841,N_8354,N_8058);
nand U8842 (N_8842,N_8492,N_8490);
and U8843 (N_8843,N_8028,N_8272);
nand U8844 (N_8844,N_8086,N_8099);
or U8845 (N_8845,N_8462,N_8170);
or U8846 (N_8846,N_8017,N_8227);
or U8847 (N_8847,N_8104,N_8256);
and U8848 (N_8848,N_8249,N_8048);
nor U8849 (N_8849,N_8364,N_8200);
and U8850 (N_8850,N_8317,N_8247);
xor U8851 (N_8851,N_8496,N_8213);
and U8852 (N_8852,N_8257,N_8337);
or U8853 (N_8853,N_8093,N_8131);
xnor U8854 (N_8854,N_8225,N_8194);
and U8855 (N_8855,N_8144,N_8472);
nor U8856 (N_8856,N_8350,N_8042);
xor U8857 (N_8857,N_8097,N_8129);
nor U8858 (N_8858,N_8035,N_8380);
and U8859 (N_8859,N_8251,N_8094);
xnor U8860 (N_8860,N_8337,N_8353);
nor U8861 (N_8861,N_8258,N_8347);
and U8862 (N_8862,N_8025,N_8385);
or U8863 (N_8863,N_8262,N_8359);
xor U8864 (N_8864,N_8174,N_8116);
nand U8865 (N_8865,N_8382,N_8282);
nor U8866 (N_8866,N_8231,N_8421);
or U8867 (N_8867,N_8042,N_8441);
nand U8868 (N_8868,N_8078,N_8090);
and U8869 (N_8869,N_8052,N_8086);
xor U8870 (N_8870,N_8205,N_8100);
nor U8871 (N_8871,N_8416,N_8225);
or U8872 (N_8872,N_8400,N_8479);
and U8873 (N_8873,N_8214,N_8491);
nor U8874 (N_8874,N_8244,N_8309);
and U8875 (N_8875,N_8227,N_8208);
and U8876 (N_8876,N_8282,N_8292);
xor U8877 (N_8877,N_8124,N_8343);
and U8878 (N_8878,N_8267,N_8493);
nand U8879 (N_8879,N_8349,N_8226);
and U8880 (N_8880,N_8333,N_8216);
or U8881 (N_8881,N_8185,N_8125);
and U8882 (N_8882,N_8109,N_8247);
nand U8883 (N_8883,N_8216,N_8357);
or U8884 (N_8884,N_8466,N_8029);
nor U8885 (N_8885,N_8198,N_8159);
nor U8886 (N_8886,N_8388,N_8116);
nand U8887 (N_8887,N_8274,N_8044);
nand U8888 (N_8888,N_8466,N_8381);
nand U8889 (N_8889,N_8165,N_8153);
nand U8890 (N_8890,N_8262,N_8350);
xnor U8891 (N_8891,N_8148,N_8392);
nand U8892 (N_8892,N_8174,N_8072);
nand U8893 (N_8893,N_8071,N_8088);
nor U8894 (N_8894,N_8215,N_8199);
or U8895 (N_8895,N_8271,N_8112);
and U8896 (N_8896,N_8483,N_8294);
nand U8897 (N_8897,N_8082,N_8139);
nor U8898 (N_8898,N_8226,N_8056);
or U8899 (N_8899,N_8358,N_8386);
or U8900 (N_8900,N_8183,N_8046);
nand U8901 (N_8901,N_8249,N_8275);
or U8902 (N_8902,N_8172,N_8130);
or U8903 (N_8903,N_8239,N_8404);
or U8904 (N_8904,N_8351,N_8103);
or U8905 (N_8905,N_8107,N_8165);
nand U8906 (N_8906,N_8289,N_8274);
nor U8907 (N_8907,N_8045,N_8180);
xor U8908 (N_8908,N_8216,N_8081);
or U8909 (N_8909,N_8073,N_8265);
xor U8910 (N_8910,N_8232,N_8305);
and U8911 (N_8911,N_8111,N_8098);
or U8912 (N_8912,N_8176,N_8188);
or U8913 (N_8913,N_8064,N_8418);
and U8914 (N_8914,N_8159,N_8432);
or U8915 (N_8915,N_8431,N_8171);
and U8916 (N_8916,N_8006,N_8054);
nor U8917 (N_8917,N_8490,N_8289);
nor U8918 (N_8918,N_8273,N_8208);
xor U8919 (N_8919,N_8015,N_8474);
nand U8920 (N_8920,N_8034,N_8364);
and U8921 (N_8921,N_8136,N_8012);
nand U8922 (N_8922,N_8490,N_8430);
nor U8923 (N_8923,N_8144,N_8338);
or U8924 (N_8924,N_8030,N_8354);
nor U8925 (N_8925,N_8131,N_8318);
nor U8926 (N_8926,N_8461,N_8482);
xor U8927 (N_8927,N_8427,N_8035);
or U8928 (N_8928,N_8387,N_8441);
xnor U8929 (N_8929,N_8424,N_8485);
or U8930 (N_8930,N_8093,N_8246);
xor U8931 (N_8931,N_8163,N_8337);
nor U8932 (N_8932,N_8450,N_8029);
nor U8933 (N_8933,N_8151,N_8014);
and U8934 (N_8934,N_8396,N_8210);
and U8935 (N_8935,N_8119,N_8148);
nand U8936 (N_8936,N_8101,N_8368);
or U8937 (N_8937,N_8225,N_8116);
nand U8938 (N_8938,N_8087,N_8325);
and U8939 (N_8939,N_8339,N_8309);
and U8940 (N_8940,N_8404,N_8079);
and U8941 (N_8941,N_8399,N_8148);
or U8942 (N_8942,N_8384,N_8003);
and U8943 (N_8943,N_8147,N_8198);
and U8944 (N_8944,N_8126,N_8180);
or U8945 (N_8945,N_8489,N_8333);
nor U8946 (N_8946,N_8002,N_8469);
nand U8947 (N_8947,N_8189,N_8149);
nor U8948 (N_8948,N_8039,N_8126);
and U8949 (N_8949,N_8263,N_8439);
or U8950 (N_8950,N_8400,N_8465);
nand U8951 (N_8951,N_8479,N_8387);
xor U8952 (N_8952,N_8027,N_8073);
nor U8953 (N_8953,N_8318,N_8217);
nand U8954 (N_8954,N_8427,N_8077);
nor U8955 (N_8955,N_8037,N_8447);
and U8956 (N_8956,N_8373,N_8397);
and U8957 (N_8957,N_8281,N_8390);
xor U8958 (N_8958,N_8104,N_8099);
nand U8959 (N_8959,N_8226,N_8473);
nand U8960 (N_8960,N_8360,N_8332);
nand U8961 (N_8961,N_8469,N_8435);
nor U8962 (N_8962,N_8038,N_8474);
and U8963 (N_8963,N_8329,N_8193);
nor U8964 (N_8964,N_8007,N_8082);
nand U8965 (N_8965,N_8332,N_8047);
and U8966 (N_8966,N_8270,N_8144);
and U8967 (N_8967,N_8321,N_8430);
xnor U8968 (N_8968,N_8038,N_8393);
or U8969 (N_8969,N_8378,N_8065);
nor U8970 (N_8970,N_8055,N_8049);
and U8971 (N_8971,N_8451,N_8199);
or U8972 (N_8972,N_8288,N_8015);
and U8973 (N_8973,N_8001,N_8377);
or U8974 (N_8974,N_8457,N_8259);
nor U8975 (N_8975,N_8275,N_8474);
nor U8976 (N_8976,N_8144,N_8303);
or U8977 (N_8977,N_8118,N_8359);
nor U8978 (N_8978,N_8125,N_8222);
nor U8979 (N_8979,N_8012,N_8040);
xnor U8980 (N_8980,N_8260,N_8101);
or U8981 (N_8981,N_8152,N_8327);
or U8982 (N_8982,N_8327,N_8193);
and U8983 (N_8983,N_8243,N_8054);
nor U8984 (N_8984,N_8284,N_8003);
nand U8985 (N_8985,N_8449,N_8158);
nand U8986 (N_8986,N_8460,N_8066);
nand U8987 (N_8987,N_8244,N_8229);
or U8988 (N_8988,N_8361,N_8475);
nor U8989 (N_8989,N_8260,N_8368);
or U8990 (N_8990,N_8454,N_8435);
nand U8991 (N_8991,N_8363,N_8268);
or U8992 (N_8992,N_8367,N_8165);
nor U8993 (N_8993,N_8057,N_8400);
or U8994 (N_8994,N_8412,N_8150);
nor U8995 (N_8995,N_8456,N_8449);
or U8996 (N_8996,N_8109,N_8287);
and U8997 (N_8997,N_8385,N_8086);
nor U8998 (N_8998,N_8238,N_8094);
and U8999 (N_8999,N_8131,N_8467);
nor U9000 (N_9000,N_8868,N_8543);
nor U9001 (N_9001,N_8887,N_8792);
nor U9002 (N_9002,N_8507,N_8917);
nor U9003 (N_9003,N_8939,N_8691);
or U9004 (N_9004,N_8934,N_8885);
nand U9005 (N_9005,N_8841,N_8748);
nor U9006 (N_9006,N_8951,N_8919);
nand U9007 (N_9007,N_8640,N_8548);
xnor U9008 (N_9008,N_8718,N_8856);
xor U9009 (N_9009,N_8801,N_8671);
or U9010 (N_9010,N_8838,N_8561);
nand U9011 (N_9011,N_8763,N_8778);
and U9012 (N_9012,N_8832,N_8782);
nor U9013 (N_9013,N_8979,N_8924);
and U9014 (N_9014,N_8733,N_8634);
nor U9015 (N_9015,N_8730,N_8511);
and U9016 (N_9016,N_8674,N_8862);
and U9017 (N_9017,N_8867,N_8946);
xor U9018 (N_9018,N_8699,N_8851);
and U9019 (N_9019,N_8631,N_8847);
nand U9020 (N_9020,N_8710,N_8807);
and U9021 (N_9021,N_8920,N_8745);
and U9022 (N_9022,N_8857,N_8639);
xnor U9023 (N_9023,N_8654,N_8692);
nor U9024 (N_9024,N_8864,N_8813);
xor U9025 (N_9025,N_8812,N_8943);
or U9026 (N_9026,N_8817,N_8609);
nand U9027 (N_9027,N_8992,N_8514);
and U9028 (N_9028,N_8760,N_8605);
or U9029 (N_9029,N_8980,N_8646);
or U9030 (N_9030,N_8906,N_8873);
nor U9031 (N_9031,N_8628,N_8796);
and U9032 (N_9032,N_8546,N_8550);
and U9033 (N_9033,N_8708,N_8712);
nand U9034 (N_9034,N_8642,N_8736);
or U9035 (N_9035,N_8914,N_8690);
nor U9036 (N_9036,N_8500,N_8576);
nand U9037 (N_9037,N_8876,N_8974);
and U9038 (N_9038,N_8833,N_8821);
nand U9039 (N_9039,N_8955,N_8790);
nand U9040 (N_9040,N_8982,N_8701);
and U9041 (N_9041,N_8695,N_8773);
or U9042 (N_9042,N_8777,N_8669);
nor U9043 (N_9043,N_8515,N_8988);
or U9044 (N_9044,N_8970,N_8912);
nor U9045 (N_9045,N_8618,N_8751);
nor U9046 (N_9046,N_8643,N_8901);
xor U9047 (N_9047,N_8881,N_8863);
nor U9048 (N_9048,N_8975,N_8855);
nor U9049 (N_9049,N_8936,N_8615);
nor U9050 (N_9050,N_8503,N_8961);
nor U9051 (N_9051,N_8984,N_8597);
and U9052 (N_9052,N_8987,N_8656);
or U9053 (N_9053,N_8884,N_8960);
nand U9054 (N_9054,N_8888,N_8775);
and U9055 (N_9055,N_8532,N_8729);
and U9056 (N_9056,N_8520,N_8555);
or U9057 (N_9057,N_8740,N_8573);
or U9058 (N_9058,N_8541,N_8562);
and U9059 (N_9059,N_8588,N_8506);
or U9060 (N_9060,N_8697,N_8678);
nor U9061 (N_9061,N_8571,N_8713);
or U9062 (N_9062,N_8891,N_8592);
nand U9063 (N_9063,N_8818,N_8995);
xnor U9064 (N_9064,N_8596,N_8799);
nor U9065 (N_9065,N_8587,N_8976);
or U9066 (N_9066,N_8870,N_8591);
and U9067 (N_9067,N_8971,N_8521);
and U9068 (N_9068,N_8719,N_8808);
nor U9069 (N_9069,N_8516,N_8663);
xnor U9070 (N_9070,N_8595,N_8880);
nand U9071 (N_9071,N_8534,N_8518);
nand U9072 (N_9072,N_8580,N_8608);
nor U9073 (N_9073,N_8973,N_8684);
nand U9074 (N_9074,N_8524,N_8517);
nand U9075 (N_9075,N_8582,N_8781);
nor U9076 (N_9076,N_8900,N_8927);
or U9077 (N_9077,N_8836,N_8861);
nand U9078 (N_9078,N_8523,N_8721);
nor U9079 (N_9079,N_8840,N_8624);
nand U9080 (N_9080,N_8525,N_8661);
nor U9081 (N_9081,N_8788,N_8787);
and U9082 (N_9082,N_8675,N_8752);
nand U9083 (N_9083,N_8584,N_8724);
or U9084 (N_9084,N_8758,N_8700);
nand U9085 (N_9085,N_8784,N_8803);
nor U9086 (N_9086,N_8839,N_8741);
nand U9087 (N_9087,N_8600,N_8767);
xnor U9088 (N_9088,N_8513,N_8965);
or U9089 (N_9089,N_8526,N_8579);
nand U9090 (N_9090,N_8865,N_8593);
nor U9091 (N_9091,N_8732,N_8893);
nor U9092 (N_9092,N_8501,N_8715);
or U9093 (N_9093,N_8785,N_8791);
nand U9094 (N_9094,N_8610,N_8735);
nand U9095 (N_9095,N_8720,N_8940);
nor U9096 (N_9096,N_8819,N_8916);
nand U9097 (N_9097,N_8948,N_8963);
nand U9098 (N_9098,N_8589,N_8744);
and U9099 (N_9099,N_8983,N_8854);
nand U9100 (N_9100,N_8665,N_8779);
nand U9101 (N_9101,N_8683,N_8815);
nand U9102 (N_9102,N_8657,N_8673);
and U9103 (N_9103,N_8677,N_8537);
nand U9104 (N_9104,N_8535,N_8874);
or U9105 (N_9105,N_8826,N_8585);
and U9106 (N_9106,N_8911,N_8793);
nand U9107 (N_9107,N_8613,N_8886);
nand U9108 (N_9108,N_8959,N_8575);
or U9109 (N_9109,N_8658,N_8962);
and U9110 (N_9110,N_8547,N_8583);
or U9111 (N_9111,N_8853,N_8858);
or U9112 (N_9112,N_8505,N_8820);
and U9113 (N_9113,N_8850,N_8765);
nor U9114 (N_9114,N_8937,N_8923);
nor U9115 (N_9115,N_8830,N_8908);
and U9116 (N_9116,N_8648,N_8805);
and U9117 (N_9117,N_8687,N_8620);
nor U9118 (N_9118,N_8871,N_8577);
and U9119 (N_9119,N_8892,N_8737);
and U9120 (N_9120,N_8753,N_8883);
xor U9121 (N_9121,N_8626,N_8652);
and U9122 (N_9122,N_8705,N_8702);
nand U9123 (N_9123,N_8616,N_8717);
nor U9124 (N_9124,N_8574,N_8825);
xor U9125 (N_9125,N_8829,N_8953);
nand U9126 (N_9126,N_8707,N_8531);
or U9127 (N_9127,N_8756,N_8795);
nand U9128 (N_9128,N_8997,N_8941);
nor U9129 (N_9129,N_8672,N_8660);
and U9130 (N_9130,N_8590,N_8998);
and U9131 (N_9131,N_8860,N_8727);
or U9132 (N_9132,N_8670,N_8694);
or U9133 (N_9133,N_8545,N_8688);
or U9134 (N_9134,N_8913,N_8930);
or U9135 (N_9135,N_8896,N_8558);
nor U9136 (N_9136,N_8538,N_8950);
or U9137 (N_9137,N_8933,N_8957);
nand U9138 (N_9138,N_8848,N_8614);
xnor U9139 (N_9139,N_8723,N_8931);
and U9140 (N_9140,N_8766,N_8556);
nor U9141 (N_9141,N_8722,N_8966);
nor U9142 (N_9142,N_8804,N_8759);
xor U9143 (N_9143,N_8899,N_8586);
and U9144 (N_9144,N_8789,N_8774);
nand U9145 (N_9145,N_8739,N_8602);
or U9146 (N_9146,N_8890,N_8676);
and U9147 (N_9147,N_8664,N_8686);
nand U9148 (N_9148,N_8823,N_8859);
nor U9149 (N_9149,N_8843,N_8742);
nor U9150 (N_9150,N_8604,N_8990);
nor U9151 (N_9151,N_8749,N_8544);
nand U9152 (N_9152,N_8668,N_8551);
nor U9153 (N_9153,N_8882,N_8952);
or U9154 (N_9154,N_8780,N_8747);
or U9155 (N_9155,N_8557,N_8612);
or U9156 (N_9156,N_8809,N_8606);
or U9157 (N_9157,N_8875,N_8566);
or U9158 (N_9158,N_8949,N_8800);
nor U9159 (N_9159,N_8905,N_8869);
or U9160 (N_9160,N_8650,N_8828);
or U9161 (N_9161,N_8806,N_8834);
nand U9162 (N_9162,N_8989,N_8932);
or U9163 (N_9163,N_8728,N_8978);
or U9164 (N_9164,N_8918,N_8837);
or U9165 (N_9165,N_8824,N_8897);
xnor U9166 (N_9166,N_8827,N_8772);
and U9167 (N_9167,N_8977,N_8845);
or U9168 (N_9168,N_8659,N_8958);
nand U9169 (N_9169,N_8904,N_8549);
nor U9170 (N_9170,N_8846,N_8651);
or U9171 (N_9171,N_8693,N_8637);
nor U9172 (N_9172,N_8638,N_8928);
nor U9173 (N_9173,N_8552,N_8910);
or U9174 (N_9174,N_8986,N_8954);
nand U9175 (N_9175,N_8852,N_8761);
and U9176 (N_9176,N_8944,N_8783);
or U9177 (N_9177,N_8641,N_8762);
and U9178 (N_9178,N_8565,N_8529);
nand U9179 (N_9179,N_8611,N_8706);
xor U9180 (N_9180,N_8764,N_8771);
and U9181 (N_9181,N_8502,N_8926);
xor U9182 (N_9182,N_8925,N_8536);
and U9183 (N_9183,N_8725,N_8607);
xor U9184 (N_9184,N_8716,N_8945);
nand U9185 (N_9185,N_8842,N_8994);
and U9186 (N_9186,N_8530,N_8680);
and U9187 (N_9187,N_8522,N_8999);
or U9188 (N_9188,N_8738,N_8872);
or U9189 (N_9189,N_8619,N_8797);
and U9190 (N_9190,N_8877,N_8704);
nand U9191 (N_9191,N_8746,N_8563);
nor U9192 (N_9192,N_8902,N_8559);
or U9193 (N_9193,N_8889,N_8844);
nand U9194 (N_9194,N_8972,N_8644);
xor U9195 (N_9195,N_8798,N_8578);
nor U9196 (N_9196,N_8636,N_8662);
nor U9197 (N_9197,N_8993,N_8731);
and U9198 (N_9198,N_8567,N_8509);
nand U9199 (N_9199,N_8968,N_8776);
or U9200 (N_9200,N_8569,N_8816);
xor U9201 (N_9201,N_8527,N_8560);
and U9202 (N_9202,N_8938,N_8603);
and U9203 (N_9203,N_8627,N_8935);
or U9204 (N_9204,N_8907,N_8598);
nor U9205 (N_9205,N_8985,N_8625);
or U9206 (N_9206,N_8622,N_8568);
and U9207 (N_9207,N_8647,N_8956);
nand U9208 (N_9208,N_8831,N_8572);
nand U9209 (N_9209,N_8947,N_8630);
or U9210 (N_9210,N_8981,N_8755);
or U9211 (N_9211,N_8570,N_8681);
xor U9212 (N_9212,N_8653,N_8786);
or U9213 (N_9213,N_8814,N_8743);
and U9214 (N_9214,N_8768,N_8645);
or U9215 (N_9215,N_8682,N_8508);
and U9216 (N_9216,N_8822,N_8810);
and U9217 (N_9217,N_8703,N_8689);
and U9218 (N_9218,N_8696,N_8750);
or U9219 (N_9219,N_8757,N_8633);
nand U9220 (N_9220,N_8964,N_8835);
nand U9221 (N_9221,N_8922,N_8564);
xor U9222 (N_9222,N_8667,N_8866);
and U9223 (N_9223,N_8942,N_8711);
nand U9224 (N_9224,N_8540,N_8734);
nand U9225 (N_9225,N_8802,N_8542);
and U9226 (N_9226,N_8754,N_8991);
or U9227 (N_9227,N_8915,N_8698);
nor U9228 (N_9228,N_8632,N_8581);
nand U9229 (N_9229,N_8649,N_8849);
or U9230 (N_9230,N_8903,N_8623);
nand U9231 (N_9231,N_8655,N_8635);
nor U9232 (N_9232,N_8878,N_8519);
or U9233 (N_9233,N_8528,N_8601);
or U9234 (N_9234,N_8996,N_8510);
nand U9235 (N_9235,N_8794,N_8594);
and U9236 (N_9236,N_8894,N_8929);
or U9237 (N_9237,N_8726,N_8539);
nand U9238 (N_9238,N_8533,N_8770);
or U9239 (N_9239,N_8811,N_8666);
nor U9240 (N_9240,N_8617,N_8599);
xor U9241 (N_9241,N_8504,N_8629);
and U9242 (N_9242,N_8769,N_8909);
or U9243 (N_9243,N_8714,N_8967);
nand U9244 (N_9244,N_8709,N_8553);
and U9245 (N_9245,N_8512,N_8879);
and U9246 (N_9246,N_8969,N_8621);
nand U9247 (N_9247,N_8554,N_8679);
xnor U9248 (N_9248,N_8895,N_8921);
or U9249 (N_9249,N_8685,N_8898);
nor U9250 (N_9250,N_8917,N_8775);
or U9251 (N_9251,N_8977,N_8661);
nor U9252 (N_9252,N_8788,N_8585);
and U9253 (N_9253,N_8970,N_8694);
or U9254 (N_9254,N_8567,N_8864);
nand U9255 (N_9255,N_8697,N_8910);
nor U9256 (N_9256,N_8629,N_8520);
nand U9257 (N_9257,N_8843,N_8737);
nand U9258 (N_9258,N_8858,N_8724);
and U9259 (N_9259,N_8842,N_8951);
or U9260 (N_9260,N_8825,N_8794);
nor U9261 (N_9261,N_8740,N_8509);
nand U9262 (N_9262,N_8892,N_8753);
xor U9263 (N_9263,N_8846,N_8799);
nor U9264 (N_9264,N_8993,N_8688);
or U9265 (N_9265,N_8973,N_8907);
and U9266 (N_9266,N_8872,N_8908);
nor U9267 (N_9267,N_8648,N_8813);
nand U9268 (N_9268,N_8746,N_8501);
or U9269 (N_9269,N_8839,N_8720);
nand U9270 (N_9270,N_8779,N_8775);
xnor U9271 (N_9271,N_8752,N_8953);
or U9272 (N_9272,N_8659,N_8725);
and U9273 (N_9273,N_8742,N_8753);
nand U9274 (N_9274,N_8718,N_8874);
or U9275 (N_9275,N_8718,N_8780);
nor U9276 (N_9276,N_8899,N_8570);
nand U9277 (N_9277,N_8581,N_8635);
or U9278 (N_9278,N_8566,N_8858);
or U9279 (N_9279,N_8965,N_8851);
nor U9280 (N_9280,N_8850,N_8949);
nand U9281 (N_9281,N_8572,N_8610);
and U9282 (N_9282,N_8802,N_8645);
or U9283 (N_9283,N_8587,N_8880);
xor U9284 (N_9284,N_8779,N_8804);
and U9285 (N_9285,N_8567,N_8872);
nand U9286 (N_9286,N_8647,N_8845);
nor U9287 (N_9287,N_8684,N_8970);
nor U9288 (N_9288,N_8841,N_8663);
and U9289 (N_9289,N_8816,N_8934);
xnor U9290 (N_9290,N_8887,N_8674);
nand U9291 (N_9291,N_8814,N_8512);
nand U9292 (N_9292,N_8856,N_8556);
or U9293 (N_9293,N_8775,N_8960);
nor U9294 (N_9294,N_8529,N_8872);
nor U9295 (N_9295,N_8618,N_8981);
or U9296 (N_9296,N_8663,N_8656);
xor U9297 (N_9297,N_8557,N_8819);
nand U9298 (N_9298,N_8627,N_8914);
nand U9299 (N_9299,N_8996,N_8833);
nor U9300 (N_9300,N_8950,N_8992);
and U9301 (N_9301,N_8874,N_8883);
and U9302 (N_9302,N_8549,N_8674);
and U9303 (N_9303,N_8984,N_8507);
xor U9304 (N_9304,N_8736,N_8775);
or U9305 (N_9305,N_8826,N_8588);
and U9306 (N_9306,N_8573,N_8929);
or U9307 (N_9307,N_8568,N_8938);
or U9308 (N_9308,N_8668,N_8640);
or U9309 (N_9309,N_8852,N_8651);
xor U9310 (N_9310,N_8948,N_8914);
and U9311 (N_9311,N_8570,N_8545);
nand U9312 (N_9312,N_8544,N_8667);
nand U9313 (N_9313,N_8725,N_8731);
and U9314 (N_9314,N_8633,N_8732);
nor U9315 (N_9315,N_8870,N_8586);
nor U9316 (N_9316,N_8849,N_8744);
nor U9317 (N_9317,N_8611,N_8901);
nor U9318 (N_9318,N_8795,N_8545);
xnor U9319 (N_9319,N_8995,N_8557);
nand U9320 (N_9320,N_8696,N_8608);
and U9321 (N_9321,N_8651,N_8634);
nor U9322 (N_9322,N_8826,N_8814);
or U9323 (N_9323,N_8986,N_8754);
nor U9324 (N_9324,N_8713,N_8969);
or U9325 (N_9325,N_8723,N_8770);
or U9326 (N_9326,N_8807,N_8556);
xnor U9327 (N_9327,N_8532,N_8856);
nand U9328 (N_9328,N_8512,N_8986);
nor U9329 (N_9329,N_8966,N_8634);
xnor U9330 (N_9330,N_8724,N_8523);
nor U9331 (N_9331,N_8778,N_8857);
nor U9332 (N_9332,N_8958,N_8529);
nor U9333 (N_9333,N_8524,N_8981);
and U9334 (N_9334,N_8933,N_8592);
xnor U9335 (N_9335,N_8507,N_8873);
xor U9336 (N_9336,N_8815,N_8850);
and U9337 (N_9337,N_8698,N_8681);
or U9338 (N_9338,N_8502,N_8711);
nand U9339 (N_9339,N_8959,N_8564);
xnor U9340 (N_9340,N_8855,N_8660);
and U9341 (N_9341,N_8575,N_8503);
xnor U9342 (N_9342,N_8544,N_8863);
or U9343 (N_9343,N_8984,N_8969);
or U9344 (N_9344,N_8681,N_8856);
nor U9345 (N_9345,N_8803,N_8719);
nand U9346 (N_9346,N_8997,N_8752);
and U9347 (N_9347,N_8913,N_8775);
and U9348 (N_9348,N_8545,N_8551);
nand U9349 (N_9349,N_8850,N_8760);
nor U9350 (N_9350,N_8967,N_8698);
and U9351 (N_9351,N_8655,N_8566);
or U9352 (N_9352,N_8985,N_8614);
or U9353 (N_9353,N_8524,N_8520);
and U9354 (N_9354,N_8893,N_8548);
and U9355 (N_9355,N_8717,N_8989);
nand U9356 (N_9356,N_8660,N_8548);
or U9357 (N_9357,N_8975,N_8869);
and U9358 (N_9358,N_8796,N_8540);
nor U9359 (N_9359,N_8773,N_8503);
nand U9360 (N_9360,N_8567,N_8998);
and U9361 (N_9361,N_8997,N_8905);
and U9362 (N_9362,N_8924,N_8575);
or U9363 (N_9363,N_8682,N_8671);
nand U9364 (N_9364,N_8878,N_8569);
or U9365 (N_9365,N_8675,N_8991);
nor U9366 (N_9366,N_8834,N_8593);
nor U9367 (N_9367,N_8985,N_8844);
and U9368 (N_9368,N_8597,N_8514);
nor U9369 (N_9369,N_8885,N_8503);
and U9370 (N_9370,N_8776,N_8529);
or U9371 (N_9371,N_8609,N_8813);
nor U9372 (N_9372,N_8957,N_8935);
xnor U9373 (N_9373,N_8908,N_8529);
and U9374 (N_9374,N_8558,N_8756);
xnor U9375 (N_9375,N_8885,N_8908);
and U9376 (N_9376,N_8982,N_8909);
or U9377 (N_9377,N_8819,N_8667);
nand U9378 (N_9378,N_8934,N_8853);
or U9379 (N_9379,N_8855,N_8571);
or U9380 (N_9380,N_8936,N_8983);
nand U9381 (N_9381,N_8891,N_8888);
and U9382 (N_9382,N_8968,N_8601);
nand U9383 (N_9383,N_8963,N_8691);
nand U9384 (N_9384,N_8522,N_8552);
nor U9385 (N_9385,N_8947,N_8719);
nor U9386 (N_9386,N_8891,N_8918);
nor U9387 (N_9387,N_8983,N_8750);
or U9388 (N_9388,N_8903,N_8659);
nand U9389 (N_9389,N_8520,N_8880);
or U9390 (N_9390,N_8560,N_8667);
or U9391 (N_9391,N_8707,N_8658);
nand U9392 (N_9392,N_8622,N_8760);
and U9393 (N_9393,N_8671,N_8975);
nand U9394 (N_9394,N_8823,N_8563);
or U9395 (N_9395,N_8961,N_8812);
nor U9396 (N_9396,N_8824,N_8778);
xnor U9397 (N_9397,N_8671,N_8993);
or U9398 (N_9398,N_8714,N_8904);
nand U9399 (N_9399,N_8616,N_8750);
nor U9400 (N_9400,N_8867,N_8674);
or U9401 (N_9401,N_8552,N_8616);
and U9402 (N_9402,N_8994,N_8711);
and U9403 (N_9403,N_8807,N_8716);
nand U9404 (N_9404,N_8561,N_8757);
or U9405 (N_9405,N_8895,N_8906);
or U9406 (N_9406,N_8918,N_8541);
or U9407 (N_9407,N_8530,N_8955);
and U9408 (N_9408,N_8762,N_8653);
nor U9409 (N_9409,N_8757,N_8875);
and U9410 (N_9410,N_8717,N_8924);
nor U9411 (N_9411,N_8922,N_8889);
nor U9412 (N_9412,N_8613,N_8890);
or U9413 (N_9413,N_8596,N_8575);
nand U9414 (N_9414,N_8509,N_8700);
nand U9415 (N_9415,N_8753,N_8607);
or U9416 (N_9416,N_8662,N_8542);
or U9417 (N_9417,N_8507,N_8524);
and U9418 (N_9418,N_8799,N_8558);
and U9419 (N_9419,N_8549,N_8500);
nor U9420 (N_9420,N_8678,N_8868);
nand U9421 (N_9421,N_8724,N_8746);
or U9422 (N_9422,N_8531,N_8741);
nand U9423 (N_9423,N_8777,N_8670);
or U9424 (N_9424,N_8791,N_8962);
nand U9425 (N_9425,N_8989,N_8659);
nand U9426 (N_9426,N_8971,N_8751);
or U9427 (N_9427,N_8949,N_8571);
and U9428 (N_9428,N_8878,N_8917);
nor U9429 (N_9429,N_8988,N_8736);
and U9430 (N_9430,N_8982,N_8606);
nand U9431 (N_9431,N_8567,N_8542);
xor U9432 (N_9432,N_8792,N_8937);
or U9433 (N_9433,N_8901,N_8612);
and U9434 (N_9434,N_8566,N_8505);
or U9435 (N_9435,N_8876,N_8618);
and U9436 (N_9436,N_8575,N_8530);
nand U9437 (N_9437,N_8745,N_8839);
or U9438 (N_9438,N_8765,N_8941);
xnor U9439 (N_9439,N_8901,N_8825);
nand U9440 (N_9440,N_8902,N_8965);
and U9441 (N_9441,N_8783,N_8587);
nand U9442 (N_9442,N_8719,N_8891);
nor U9443 (N_9443,N_8518,N_8970);
and U9444 (N_9444,N_8952,N_8706);
and U9445 (N_9445,N_8878,N_8573);
xor U9446 (N_9446,N_8906,N_8822);
nand U9447 (N_9447,N_8838,N_8746);
and U9448 (N_9448,N_8639,N_8654);
nor U9449 (N_9449,N_8672,N_8642);
and U9450 (N_9450,N_8585,N_8604);
and U9451 (N_9451,N_8942,N_8745);
or U9452 (N_9452,N_8835,N_8902);
xnor U9453 (N_9453,N_8663,N_8712);
nor U9454 (N_9454,N_8961,N_8528);
and U9455 (N_9455,N_8704,N_8752);
or U9456 (N_9456,N_8571,N_8711);
nor U9457 (N_9457,N_8967,N_8972);
and U9458 (N_9458,N_8911,N_8595);
nand U9459 (N_9459,N_8731,N_8857);
xnor U9460 (N_9460,N_8563,N_8521);
xor U9461 (N_9461,N_8698,N_8561);
nor U9462 (N_9462,N_8848,N_8906);
nand U9463 (N_9463,N_8645,N_8605);
and U9464 (N_9464,N_8524,N_8985);
and U9465 (N_9465,N_8741,N_8860);
or U9466 (N_9466,N_8821,N_8756);
nor U9467 (N_9467,N_8958,N_8825);
nor U9468 (N_9468,N_8647,N_8621);
and U9469 (N_9469,N_8565,N_8875);
nand U9470 (N_9470,N_8827,N_8620);
nand U9471 (N_9471,N_8574,N_8942);
and U9472 (N_9472,N_8613,N_8877);
or U9473 (N_9473,N_8762,N_8995);
nand U9474 (N_9474,N_8996,N_8887);
nor U9475 (N_9475,N_8966,N_8745);
nor U9476 (N_9476,N_8535,N_8926);
nand U9477 (N_9477,N_8585,N_8775);
and U9478 (N_9478,N_8787,N_8885);
or U9479 (N_9479,N_8831,N_8742);
and U9480 (N_9480,N_8611,N_8598);
nor U9481 (N_9481,N_8927,N_8739);
nand U9482 (N_9482,N_8987,N_8749);
or U9483 (N_9483,N_8645,N_8901);
nor U9484 (N_9484,N_8824,N_8586);
nand U9485 (N_9485,N_8668,N_8634);
and U9486 (N_9486,N_8536,N_8544);
nand U9487 (N_9487,N_8751,N_8717);
or U9488 (N_9488,N_8820,N_8603);
xnor U9489 (N_9489,N_8791,N_8977);
or U9490 (N_9490,N_8965,N_8884);
xnor U9491 (N_9491,N_8815,N_8690);
or U9492 (N_9492,N_8576,N_8833);
xor U9493 (N_9493,N_8991,N_8862);
and U9494 (N_9494,N_8832,N_8852);
or U9495 (N_9495,N_8757,N_8847);
and U9496 (N_9496,N_8686,N_8769);
or U9497 (N_9497,N_8825,N_8543);
nand U9498 (N_9498,N_8891,N_8906);
nand U9499 (N_9499,N_8511,N_8735);
nor U9500 (N_9500,N_9354,N_9058);
or U9501 (N_9501,N_9466,N_9320);
nor U9502 (N_9502,N_9421,N_9321);
xor U9503 (N_9503,N_9279,N_9254);
nor U9504 (N_9504,N_9363,N_9369);
nand U9505 (N_9505,N_9323,N_9005);
nor U9506 (N_9506,N_9343,N_9476);
and U9507 (N_9507,N_9115,N_9228);
nor U9508 (N_9508,N_9373,N_9011);
or U9509 (N_9509,N_9214,N_9422);
xnor U9510 (N_9510,N_9339,N_9418);
nor U9511 (N_9511,N_9135,N_9223);
or U9512 (N_9512,N_9206,N_9117);
and U9513 (N_9513,N_9360,N_9078);
and U9514 (N_9514,N_9127,N_9036);
or U9515 (N_9515,N_9002,N_9216);
or U9516 (N_9516,N_9434,N_9352);
xnor U9517 (N_9517,N_9004,N_9098);
nor U9518 (N_9518,N_9169,N_9329);
nor U9519 (N_9519,N_9333,N_9227);
or U9520 (N_9520,N_9197,N_9396);
or U9521 (N_9521,N_9433,N_9464);
or U9522 (N_9522,N_9139,N_9416);
nor U9523 (N_9523,N_9053,N_9217);
nand U9524 (N_9524,N_9355,N_9318);
nor U9525 (N_9525,N_9290,N_9168);
nor U9526 (N_9526,N_9457,N_9012);
or U9527 (N_9527,N_9138,N_9252);
nor U9528 (N_9528,N_9459,N_9450);
nand U9529 (N_9529,N_9406,N_9085);
or U9530 (N_9530,N_9112,N_9096);
or U9531 (N_9531,N_9345,N_9176);
xnor U9532 (N_9532,N_9385,N_9312);
nor U9533 (N_9533,N_9325,N_9439);
nand U9534 (N_9534,N_9174,N_9497);
xor U9535 (N_9535,N_9388,N_9088);
nand U9536 (N_9536,N_9179,N_9148);
or U9537 (N_9537,N_9100,N_9283);
or U9538 (N_9538,N_9192,N_9070);
or U9539 (N_9539,N_9380,N_9210);
and U9540 (N_9540,N_9118,N_9113);
or U9541 (N_9541,N_9427,N_9201);
nor U9542 (N_9542,N_9065,N_9389);
or U9543 (N_9543,N_9149,N_9026);
nand U9544 (N_9544,N_9282,N_9126);
nand U9545 (N_9545,N_9074,N_9014);
nand U9546 (N_9546,N_9027,N_9395);
xor U9547 (N_9547,N_9499,N_9049);
and U9548 (N_9548,N_9411,N_9182);
nand U9549 (N_9549,N_9082,N_9368);
or U9550 (N_9550,N_9479,N_9330);
or U9551 (N_9551,N_9019,N_9256);
nor U9552 (N_9552,N_9437,N_9247);
or U9553 (N_9553,N_9106,N_9470);
nor U9554 (N_9554,N_9000,N_9425);
and U9555 (N_9555,N_9104,N_9051);
or U9556 (N_9556,N_9491,N_9485);
nand U9557 (N_9557,N_9111,N_9401);
nor U9558 (N_9558,N_9164,N_9107);
nor U9559 (N_9559,N_9030,N_9441);
nand U9560 (N_9560,N_9097,N_9032);
xor U9561 (N_9561,N_9301,N_9089);
xnor U9562 (N_9562,N_9224,N_9317);
xor U9563 (N_9563,N_9177,N_9241);
nand U9564 (N_9564,N_9090,N_9404);
nor U9565 (N_9565,N_9167,N_9181);
nand U9566 (N_9566,N_9496,N_9195);
and U9567 (N_9567,N_9061,N_9297);
nor U9568 (N_9568,N_9315,N_9442);
nor U9569 (N_9569,N_9125,N_9230);
and U9570 (N_9570,N_9062,N_9356);
xnor U9571 (N_9571,N_9348,N_9242);
or U9572 (N_9572,N_9257,N_9474);
nand U9573 (N_9573,N_9251,N_9105);
nand U9574 (N_9574,N_9147,N_9472);
and U9575 (N_9575,N_9157,N_9291);
and U9576 (N_9576,N_9278,N_9057);
nor U9577 (N_9577,N_9481,N_9165);
nand U9578 (N_9578,N_9374,N_9314);
nor U9579 (N_9579,N_9293,N_9063);
and U9580 (N_9580,N_9150,N_9382);
nor U9581 (N_9581,N_9327,N_9467);
or U9582 (N_9582,N_9073,N_9190);
xor U9583 (N_9583,N_9072,N_9183);
nor U9584 (N_9584,N_9087,N_9048);
and U9585 (N_9585,N_9023,N_9469);
nand U9586 (N_9586,N_9219,N_9370);
or U9587 (N_9587,N_9436,N_9471);
nor U9588 (N_9588,N_9103,N_9099);
xor U9589 (N_9589,N_9400,N_9295);
and U9590 (N_9590,N_9191,N_9202);
nor U9591 (N_9591,N_9245,N_9449);
nand U9592 (N_9592,N_9303,N_9160);
nand U9593 (N_9593,N_9129,N_9233);
or U9594 (N_9594,N_9335,N_9324);
nand U9595 (N_9595,N_9494,N_9198);
xnor U9596 (N_9596,N_9122,N_9159);
nor U9597 (N_9597,N_9229,N_9358);
nand U9598 (N_9598,N_9310,N_9123);
xor U9599 (N_9599,N_9349,N_9475);
and U9600 (N_9600,N_9299,N_9402);
xnor U9601 (N_9601,N_9040,N_9218);
or U9602 (N_9602,N_9054,N_9446);
nand U9603 (N_9603,N_9137,N_9075);
or U9604 (N_9604,N_9381,N_9413);
and U9605 (N_9605,N_9430,N_9222);
and U9606 (N_9606,N_9384,N_9236);
xnor U9607 (N_9607,N_9258,N_9264);
xor U9608 (N_9608,N_9461,N_9280);
nor U9609 (N_9609,N_9371,N_9424);
and U9610 (N_9610,N_9095,N_9178);
or U9611 (N_9611,N_9018,N_9331);
nor U9612 (N_9612,N_9052,N_9340);
xor U9613 (N_9613,N_9399,N_9077);
and U9614 (N_9614,N_9044,N_9420);
or U9615 (N_9615,N_9130,N_9272);
nand U9616 (N_9616,N_9465,N_9357);
and U9617 (N_9617,N_9047,N_9488);
nand U9618 (N_9618,N_9468,N_9114);
nor U9619 (N_9619,N_9412,N_9180);
xnor U9620 (N_9620,N_9133,N_9473);
xnor U9621 (N_9621,N_9359,N_9480);
or U9622 (N_9622,N_9064,N_9492);
xnor U9623 (N_9623,N_9408,N_9394);
and U9624 (N_9624,N_9173,N_9119);
nand U9625 (N_9625,N_9265,N_9237);
and U9626 (N_9626,N_9445,N_9253);
nand U9627 (N_9627,N_9419,N_9045);
or U9628 (N_9628,N_9462,N_9175);
nor U9629 (N_9629,N_9407,N_9414);
or U9630 (N_9630,N_9255,N_9240);
and U9631 (N_9631,N_9151,N_9308);
nor U9632 (N_9632,N_9003,N_9451);
and U9633 (N_9633,N_9487,N_9203);
nand U9634 (N_9634,N_9200,N_9140);
nand U9635 (N_9635,N_9136,N_9484);
nor U9636 (N_9636,N_9336,N_9377);
nor U9637 (N_9637,N_9213,N_9337);
nand U9638 (N_9638,N_9249,N_9268);
and U9639 (N_9639,N_9132,N_9367);
or U9640 (N_9640,N_9037,N_9364);
nor U9641 (N_9641,N_9060,N_9166);
and U9642 (N_9642,N_9311,N_9486);
or U9643 (N_9643,N_9431,N_9231);
nand U9644 (N_9644,N_9378,N_9013);
or U9645 (N_9645,N_9055,N_9334);
xor U9646 (N_9646,N_9410,N_9391);
and U9647 (N_9647,N_9128,N_9188);
or U9648 (N_9648,N_9194,N_9260);
and U9649 (N_9649,N_9015,N_9435);
or U9650 (N_9650,N_9215,N_9458);
nor U9651 (N_9651,N_9020,N_9124);
nand U9652 (N_9652,N_9094,N_9269);
nor U9653 (N_9653,N_9083,N_9156);
nand U9654 (N_9654,N_9281,N_9285);
or U9655 (N_9655,N_9267,N_9134);
nand U9656 (N_9656,N_9366,N_9226);
nor U9657 (N_9657,N_9185,N_9071);
or U9658 (N_9658,N_9379,N_9306);
or U9659 (N_9659,N_9121,N_9347);
and U9660 (N_9660,N_9033,N_9398);
and U9661 (N_9661,N_9454,N_9232);
and U9662 (N_9662,N_9172,N_9009);
nand U9663 (N_9663,N_9284,N_9298);
or U9664 (N_9664,N_9289,N_9207);
nand U9665 (N_9665,N_9452,N_9432);
and U9666 (N_9666,N_9244,N_9453);
nor U9667 (N_9667,N_9438,N_9084);
xnor U9668 (N_9668,N_9235,N_9447);
xor U9669 (N_9669,N_9361,N_9131);
nor U9670 (N_9670,N_9341,N_9326);
nand U9671 (N_9671,N_9489,N_9302);
and U9672 (N_9672,N_9286,N_9250);
xor U9673 (N_9673,N_9344,N_9351);
nand U9674 (N_9674,N_9186,N_9211);
nand U9675 (N_9675,N_9066,N_9375);
nor U9676 (N_9676,N_9001,N_9184);
nand U9677 (N_9677,N_9153,N_9204);
or U9678 (N_9678,N_9155,N_9086);
xnor U9679 (N_9679,N_9035,N_9171);
nor U9680 (N_9680,N_9142,N_9495);
or U9681 (N_9681,N_9275,N_9189);
nor U9682 (N_9682,N_9332,N_9287);
or U9683 (N_9683,N_9397,N_9170);
nor U9684 (N_9684,N_9316,N_9143);
and U9685 (N_9685,N_9463,N_9383);
nand U9686 (N_9686,N_9443,N_9212);
nor U9687 (N_9687,N_9292,N_9248);
nor U9688 (N_9688,N_9386,N_9007);
and U9689 (N_9689,N_9081,N_9346);
or U9690 (N_9690,N_9225,N_9428);
and U9691 (N_9691,N_9158,N_9390);
or U9692 (N_9692,N_9307,N_9460);
nor U9693 (N_9693,N_9161,N_9262);
nor U9694 (N_9694,N_9092,N_9403);
nor U9695 (N_9695,N_9342,N_9196);
nand U9696 (N_9696,N_9405,N_9043);
nand U9697 (N_9697,N_9271,N_9220);
nor U9698 (N_9698,N_9120,N_9069);
and U9699 (N_9699,N_9456,N_9029);
nand U9700 (N_9700,N_9365,N_9163);
nand U9701 (N_9701,N_9273,N_9353);
nor U9702 (N_9702,N_9101,N_9050);
nand U9703 (N_9703,N_9234,N_9116);
xor U9704 (N_9704,N_9041,N_9038);
nand U9705 (N_9705,N_9482,N_9313);
nand U9706 (N_9706,N_9208,N_9294);
nor U9707 (N_9707,N_9409,N_9304);
or U9708 (N_9708,N_9102,N_9243);
and U9709 (N_9709,N_9109,N_9028);
and U9710 (N_9710,N_9266,N_9376);
nor U9711 (N_9711,N_9498,N_9444);
or U9712 (N_9712,N_9309,N_9093);
nand U9713 (N_9713,N_9261,N_9276);
and U9714 (N_9714,N_9328,N_9079);
or U9715 (N_9715,N_9205,N_9108);
nand U9716 (N_9716,N_9238,N_9006);
or U9717 (N_9717,N_9141,N_9490);
nor U9718 (N_9718,N_9008,N_9154);
or U9719 (N_9719,N_9392,N_9423);
nand U9720 (N_9720,N_9300,N_9221);
nor U9721 (N_9721,N_9440,N_9024);
nand U9722 (N_9722,N_9031,N_9091);
nand U9723 (N_9723,N_9259,N_9059);
or U9724 (N_9724,N_9274,N_9034);
nand U9725 (N_9725,N_9067,N_9319);
xor U9726 (N_9726,N_9152,N_9393);
nand U9727 (N_9727,N_9021,N_9322);
and U9728 (N_9728,N_9288,N_9429);
nand U9729 (N_9729,N_9263,N_9016);
xor U9730 (N_9730,N_9056,N_9146);
xnor U9731 (N_9731,N_9415,N_9017);
and U9732 (N_9732,N_9046,N_9305);
nand U9733 (N_9733,N_9270,N_9042);
or U9734 (N_9734,N_9372,N_9039);
xnor U9735 (N_9735,N_9338,N_9277);
and U9736 (N_9736,N_9426,N_9110);
or U9737 (N_9737,N_9080,N_9455);
or U9738 (N_9738,N_9478,N_9417);
nor U9739 (N_9739,N_9296,N_9162);
nor U9740 (N_9740,N_9144,N_9362);
nand U9741 (N_9741,N_9246,N_9239);
xor U9742 (N_9742,N_9350,N_9025);
and U9743 (N_9743,N_9145,N_9209);
nand U9744 (N_9744,N_9493,N_9022);
or U9745 (N_9745,N_9010,N_9477);
nor U9746 (N_9746,N_9448,N_9193);
nor U9747 (N_9747,N_9068,N_9199);
and U9748 (N_9748,N_9387,N_9483);
nor U9749 (N_9749,N_9187,N_9076);
xnor U9750 (N_9750,N_9414,N_9361);
and U9751 (N_9751,N_9198,N_9201);
or U9752 (N_9752,N_9107,N_9197);
nor U9753 (N_9753,N_9045,N_9349);
nor U9754 (N_9754,N_9097,N_9083);
or U9755 (N_9755,N_9053,N_9473);
nand U9756 (N_9756,N_9385,N_9151);
or U9757 (N_9757,N_9300,N_9246);
nand U9758 (N_9758,N_9184,N_9455);
nand U9759 (N_9759,N_9124,N_9482);
or U9760 (N_9760,N_9053,N_9209);
or U9761 (N_9761,N_9167,N_9345);
nand U9762 (N_9762,N_9441,N_9442);
or U9763 (N_9763,N_9071,N_9068);
nor U9764 (N_9764,N_9470,N_9240);
or U9765 (N_9765,N_9221,N_9036);
nor U9766 (N_9766,N_9288,N_9097);
xnor U9767 (N_9767,N_9081,N_9063);
or U9768 (N_9768,N_9286,N_9000);
or U9769 (N_9769,N_9134,N_9053);
nor U9770 (N_9770,N_9235,N_9049);
nand U9771 (N_9771,N_9329,N_9304);
xnor U9772 (N_9772,N_9120,N_9468);
nor U9773 (N_9773,N_9261,N_9046);
or U9774 (N_9774,N_9325,N_9082);
or U9775 (N_9775,N_9208,N_9234);
xnor U9776 (N_9776,N_9416,N_9034);
nand U9777 (N_9777,N_9461,N_9425);
xnor U9778 (N_9778,N_9400,N_9348);
and U9779 (N_9779,N_9385,N_9455);
nor U9780 (N_9780,N_9424,N_9219);
xnor U9781 (N_9781,N_9113,N_9324);
or U9782 (N_9782,N_9373,N_9192);
xor U9783 (N_9783,N_9327,N_9104);
and U9784 (N_9784,N_9154,N_9331);
and U9785 (N_9785,N_9254,N_9444);
nand U9786 (N_9786,N_9223,N_9443);
or U9787 (N_9787,N_9004,N_9035);
or U9788 (N_9788,N_9415,N_9316);
and U9789 (N_9789,N_9167,N_9332);
xor U9790 (N_9790,N_9423,N_9133);
nand U9791 (N_9791,N_9010,N_9213);
and U9792 (N_9792,N_9005,N_9001);
or U9793 (N_9793,N_9465,N_9005);
and U9794 (N_9794,N_9347,N_9315);
and U9795 (N_9795,N_9402,N_9336);
and U9796 (N_9796,N_9243,N_9169);
and U9797 (N_9797,N_9069,N_9414);
and U9798 (N_9798,N_9101,N_9283);
xnor U9799 (N_9799,N_9345,N_9443);
nor U9800 (N_9800,N_9110,N_9147);
nor U9801 (N_9801,N_9070,N_9047);
or U9802 (N_9802,N_9208,N_9092);
xor U9803 (N_9803,N_9065,N_9313);
xnor U9804 (N_9804,N_9089,N_9492);
nor U9805 (N_9805,N_9406,N_9389);
nor U9806 (N_9806,N_9307,N_9154);
or U9807 (N_9807,N_9117,N_9028);
xor U9808 (N_9808,N_9125,N_9209);
nor U9809 (N_9809,N_9092,N_9116);
nor U9810 (N_9810,N_9273,N_9468);
nand U9811 (N_9811,N_9277,N_9150);
xor U9812 (N_9812,N_9275,N_9253);
or U9813 (N_9813,N_9498,N_9403);
nor U9814 (N_9814,N_9203,N_9362);
and U9815 (N_9815,N_9429,N_9393);
nand U9816 (N_9816,N_9454,N_9209);
and U9817 (N_9817,N_9022,N_9243);
and U9818 (N_9818,N_9447,N_9001);
and U9819 (N_9819,N_9205,N_9206);
or U9820 (N_9820,N_9426,N_9233);
or U9821 (N_9821,N_9135,N_9366);
or U9822 (N_9822,N_9304,N_9186);
or U9823 (N_9823,N_9356,N_9081);
nor U9824 (N_9824,N_9452,N_9231);
or U9825 (N_9825,N_9165,N_9019);
nand U9826 (N_9826,N_9429,N_9100);
nor U9827 (N_9827,N_9125,N_9024);
nor U9828 (N_9828,N_9466,N_9117);
nand U9829 (N_9829,N_9312,N_9421);
nor U9830 (N_9830,N_9005,N_9472);
or U9831 (N_9831,N_9185,N_9380);
nor U9832 (N_9832,N_9406,N_9284);
or U9833 (N_9833,N_9086,N_9435);
nor U9834 (N_9834,N_9067,N_9257);
xnor U9835 (N_9835,N_9011,N_9092);
and U9836 (N_9836,N_9456,N_9175);
or U9837 (N_9837,N_9419,N_9019);
nor U9838 (N_9838,N_9070,N_9231);
nand U9839 (N_9839,N_9270,N_9487);
or U9840 (N_9840,N_9322,N_9408);
nor U9841 (N_9841,N_9295,N_9437);
and U9842 (N_9842,N_9470,N_9345);
and U9843 (N_9843,N_9118,N_9031);
nor U9844 (N_9844,N_9186,N_9113);
xnor U9845 (N_9845,N_9245,N_9459);
nor U9846 (N_9846,N_9224,N_9030);
nor U9847 (N_9847,N_9187,N_9034);
and U9848 (N_9848,N_9041,N_9391);
or U9849 (N_9849,N_9321,N_9169);
and U9850 (N_9850,N_9314,N_9230);
nand U9851 (N_9851,N_9395,N_9273);
nand U9852 (N_9852,N_9176,N_9225);
or U9853 (N_9853,N_9209,N_9237);
or U9854 (N_9854,N_9093,N_9392);
and U9855 (N_9855,N_9030,N_9166);
and U9856 (N_9856,N_9154,N_9374);
nor U9857 (N_9857,N_9273,N_9310);
nand U9858 (N_9858,N_9190,N_9178);
or U9859 (N_9859,N_9068,N_9433);
nor U9860 (N_9860,N_9356,N_9323);
nor U9861 (N_9861,N_9287,N_9430);
or U9862 (N_9862,N_9124,N_9322);
nor U9863 (N_9863,N_9176,N_9438);
and U9864 (N_9864,N_9247,N_9241);
nor U9865 (N_9865,N_9397,N_9439);
nor U9866 (N_9866,N_9050,N_9304);
nor U9867 (N_9867,N_9280,N_9086);
and U9868 (N_9868,N_9105,N_9485);
or U9869 (N_9869,N_9283,N_9407);
nand U9870 (N_9870,N_9055,N_9483);
nand U9871 (N_9871,N_9120,N_9427);
or U9872 (N_9872,N_9042,N_9449);
or U9873 (N_9873,N_9035,N_9404);
nor U9874 (N_9874,N_9048,N_9338);
nand U9875 (N_9875,N_9375,N_9146);
xor U9876 (N_9876,N_9260,N_9267);
or U9877 (N_9877,N_9030,N_9015);
or U9878 (N_9878,N_9383,N_9111);
xnor U9879 (N_9879,N_9027,N_9445);
or U9880 (N_9880,N_9341,N_9407);
and U9881 (N_9881,N_9204,N_9289);
nor U9882 (N_9882,N_9465,N_9240);
and U9883 (N_9883,N_9317,N_9308);
and U9884 (N_9884,N_9229,N_9196);
and U9885 (N_9885,N_9113,N_9234);
or U9886 (N_9886,N_9092,N_9297);
nor U9887 (N_9887,N_9346,N_9183);
and U9888 (N_9888,N_9432,N_9497);
nand U9889 (N_9889,N_9183,N_9146);
and U9890 (N_9890,N_9186,N_9124);
and U9891 (N_9891,N_9007,N_9385);
nand U9892 (N_9892,N_9172,N_9450);
or U9893 (N_9893,N_9160,N_9145);
and U9894 (N_9894,N_9313,N_9404);
and U9895 (N_9895,N_9263,N_9449);
xnor U9896 (N_9896,N_9117,N_9219);
nand U9897 (N_9897,N_9176,N_9335);
nor U9898 (N_9898,N_9287,N_9278);
nor U9899 (N_9899,N_9079,N_9087);
nor U9900 (N_9900,N_9462,N_9200);
xnor U9901 (N_9901,N_9419,N_9219);
nand U9902 (N_9902,N_9241,N_9248);
or U9903 (N_9903,N_9408,N_9119);
xnor U9904 (N_9904,N_9296,N_9490);
and U9905 (N_9905,N_9494,N_9167);
or U9906 (N_9906,N_9312,N_9269);
nor U9907 (N_9907,N_9130,N_9488);
or U9908 (N_9908,N_9247,N_9349);
nand U9909 (N_9909,N_9398,N_9393);
and U9910 (N_9910,N_9011,N_9427);
or U9911 (N_9911,N_9222,N_9056);
nor U9912 (N_9912,N_9243,N_9316);
nor U9913 (N_9913,N_9304,N_9254);
nand U9914 (N_9914,N_9035,N_9342);
and U9915 (N_9915,N_9345,N_9318);
and U9916 (N_9916,N_9404,N_9027);
or U9917 (N_9917,N_9316,N_9295);
nand U9918 (N_9918,N_9053,N_9291);
and U9919 (N_9919,N_9368,N_9291);
xor U9920 (N_9920,N_9153,N_9337);
nor U9921 (N_9921,N_9087,N_9171);
nand U9922 (N_9922,N_9003,N_9462);
nor U9923 (N_9923,N_9292,N_9205);
or U9924 (N_9924,N_9421,N_9431);
nor U9925 (N_9925,N_9464,N_9164);
nor U9926 (N_9926,N_9495,N_9336);
nand U9927 (N_9927,N_9272,N_9034);
xnor U9928 (N_9928,N_9333,N_9053);
and U9929 (N_9929,N_9345,N_9192);
nand U9930 (N_9930,N_9073,N_9027);
or U9931 (N_9931,N_9386,N_9249);
or U9932 (N_9932,N_9177,N_9379);
and U9933 (N_9933,N_9303,N_9031);
nand U9934 (N_9934,N_9134,N_9102);
xor U9935 (N_9935,N_9144,N_9480);
or U9936 (N_9936,N_9354,N_9038);
nand U9937 (N_9937,N_9156,N_9135);
and U9938 (N_9938,N_9201,N_9254);
xnor U9939 (N_9939,N_9456,N_9336);
or U9940 (N_9940,N_9485,N_9041);
nand U9941 (N_9941,N_9122,N_9001);
xor U9942 (N_9942,N_9179,N_9259);
and U9943 (N_9943,N_9252,N_9045);
and U9944 (N_9944,N_9391,N_9151);
or U9945 (N_9945,N_9480,N_9139);
or U9946 (N_9946,N_9379,N_9120);
nor U9947 (N_9947,N_9268,N_9381);
and U9948 (N_9948,N_9222,N_9213);
or U9949 (N_9949,N_9097,N_9493);
or U9950 (N_9950,N_9362,N_9151);
or U9951 (N_9951,N_9112,N_9462);
xor U9952 (N_9952,N_9342,N_9327);
and U9953 (N_9953,N_9420,N_9131);
nor U9954 (N_9954,N_9073,N_9038);
nand U9955 (N_9955,N_9093,N_9427);
and U9956 (N_9956,N_9348,N_9138);
nand U9957 (N_9957,N_9265,N_9489);
nor U9958 (N_9958,N_9414,N_9366);
xor U9959 (N_9959,N_9049,N_9208);
nor U9960 (N_9960,N_9415,N_9370);
or U9961 (N_9961,N_9247,N_9058);
nor U9962 (N_9962,N_9168,N_9361);
nand U9963 (N_9963,N_9423,N_9384);
nor U9964 (N_9964,N_9137,N_9406);
nand U9965 (N_9965,N_9325,N_9295);
nor U9966 (N_9966,N_9268,N_9170);
xnor U9967 (N_9967,N_9302,N_9362);
or U9968 (N_9968,N_9466,N_9237);
xor U9969 (N_9969,N_9069,N_9394);
or U9970 (N_9970,N_9481,N_9142);
or U9971 (N_9971,N_9246,N_9282);
nor U9972 (N_9972,N_9034,N_9444);
nor U9973 (N_9973,N_9326,N_9300);
nand U9974 (N_9974,N_9411,N_9215);
or U9975 (N_9975,N_9335,N_9277);
and U9976 (N_9976,N_9138,N_9291);
nand U9977 (N_9977,N_9379,N_9403);
or U9978 (N_9978,N_9344,N_9053);
and U9979 (N_9979,N_9258,N_9370);
and U9980 (N_9980,N_9463,N_9198);
nand U9981 (N_9981,N_9456,N_9146);
nand U9982 (N_9982,N_9039,N_9376);
nor U9983 (N_9983,N_9046,N_9350);
or U9984 (N_9984,N_9075,N_9185);
and U9985 (N_9985,N_9418,N_9091);
nor U9986 (N_9986,N_9345,N_9394);
nor U9987 (N_9987,N_9436,N_9221);
and U9988 (N_9988,N_9412,N_9269);
xnor U9989 (N_9989,N_9356,N_9415);
nor U9990 (N_9990,N_9197,N_9196);
or U9991 (N_9991,N_9010,N_9454);
or U9992 (N_9992,N_9178,N_9215);
and U9993 (N_9993,N_9470,N_9046);
or U9994 (N_9994,N_9363,N_9412);
nand U9995 (N_9995,N_9154,N_9300);
or U9996 (N_9996,N_9187,N_9266);
xnor U9997 (N_9997,N_9044,N_9333);
and U9998 (N_9998,N_9008,N_9378);
or U9999 (N_9999,N_9036,N_9265);
and UO_0 (O_0,N_9902,N_9781);
nor UO_1 (O_1,N_9555,N_9962);
or UO_2 (O_2,N_9693,N_9665);
nand UO_3 (O_3,N_9755,N_9989);
or UO_4 (O_4,N_9900,N_9698);
xnor UO_5 (O_5,N_9696,N_9787);
or UO_6 (O_6,N_9763,N_9964);
nor UO_7 (O_7,N_9792,N_9562);
nor UO_8 (O_8,N_9643,N_9651);
nand UO_9 (O_9,N_9558,N_9919);
and UO_10 (O_10,N_9894,N_9684);
xor UO_11 (O_11,N_9822,N_9738);
nand UO_12 (O_12,N_9621,N_9895);
or UO_13 (O_13,N_9987,N_9988);
xnor UO_14 (O_14,N_9906,N_9715);
and UO_15 (O_15,N_9638,N_9524);
nand UO_16 (O_16,N_9571,N_9542);
nor UO_17 (O_17,N_9582,N_9611);
and UO_18 (O_18,N_9786,N_9896);
or UO_19 (O_19,N_9659,N_9742);
nand UO_20 (O_20,N_9747,N_9637);
xnor UO_21 (O_21,N_9806,N_9623);
nor UO_22 (O_22,N_9566,N_9912);
and UO_23 (O_23,N_9624,N_9836);
nor UO_24 (O_24,N_9527,N_9517);
nor UO_25 (O_25,N_9867,N_9645);
nor UO_26 (O_26,N_9921,N_9941);
and UO_27 (O_27,N_9824,N_9625);
or UO_28 (O_28,N_9864,N_9759);
xor UO_29 (O_29,N_9930,N_9811);
and UO_30 (O_30,N_9844,N_9700);
nor UO_31 (O_31,N_9946,N_9664);
nor UO_32 (O_32,N_9866,N_9734);
or UO_33 (O_33,N_9723,N_9790);
or UO_34 (O_34,N_9676,N_9728);
or UO_35 (O_35,N_9937,N_9610);
or UO_36 (O_36,N_9854,N_9793);
nand UO_37 (O_37,N_9922,N_9579);
nand UO_38 (O_38,N_9795,N_9593);
nand UO_39 (O_39,N_9668,N_9973);
nor UO_40 (O_40,N_9914,N_9757);
nand UO_41 (O_41,N_9756,N_9628);
nand UO_42 (O_42,N_9800,N_9934);
nor UO_43 (O_43,N_9557,N_9640);
xor UO_44 (O_44,N_9762,N_9548);
nor UO_45 (O_45,N_9619,N_9620);
xor UO_46 (O_46,N_9618,N_9680);
or UO_47 (O_47,N_9646,N_9679);
or UO_48 (O_48,N_9745,N_9826);
nor UO_49 (O_49,N_9605,N_9948);
nor UO_50 (O_50,N_9871,N_9810);
nand UO_51 (O_51,N_9825,N_9660);
or UO_52 (O_52,N_9903,N_9536);
nor UO_53 (O_53,N_9513,N_9681);
xor UO_54 (O_54,N_9910,N_9899);
nand UO_55 (O_55,N_9604,N_9512);
and UO_56 (O_56,N_9617,N_9992);
nor UO_57 (O_57,N_9974,N_9586);
nor UO_58 (O_58,N_9596,N_9928);
and UO_59 (O_59,N_9960,N_9519);
or UO_60 (O_60,N_9897,N_9780);
xor UO_61 (O_61,N_9650,N_9649);
nor UO_62 (O_62,N_9803,N_9612);
nand UO_63 (O_63,N_9720,N_9556);
xor UO_64 (O_64,N_9591,N_9670);
nor UO_65 (O_65,N_9633,N_9601);
and UO_66 (O_66,N_9550,N_9600);
nand UO_67 (O_67,N_9963,N_9613);
and UO_68 (O_68,N_9944,N_9950);
or UO_69 (O_69,N_9838,N_9907);
nor UO_70 (O_70,N_9654,N_9544);
and UO_71 (O_71,N_9576,N_9705);
nand UO_72 (O_72,N_9876,N_9998);
or UO_73 (O_73,N_9563,N_9765);
nor UO_74 (O_74,N_9953,N_9794);
and UO_75 (O_75,N_9570,N_9959);
and UO_76 (O_76,N_9917,N_9961);
and UO_77 (O_77,N_9775,N_9657);
and UO_78 (O_78,N_9641,N_9594);
nor UO_79 (O_79,N_9769,N_9520);
nand UO_80 (O_80,N_9808,N_9776);
nand UO_81 (O_81,N_9719,N_9770);
or UO_82 (O_82,N_9855,N_9758);
nand UO_83 (O_83,N_9927,N_9850);
nand UO_84 (O_84,N_9722,N_9510);
and UO_85 (O_85,N_9539,N_9703);
or UO_86 (O_86,N_9791,N_9984);
and UO_87 (O_87,N_9913,N_9885);
xnor UO_88 (O_88,N_9504,N_9565);
nand UO_89 (O_89,N_9929,N_9690);
nor UO_90 (O_90,N_9678,N_9732);
or UO_91 (O_91,N_9843,N_9662);
and UO_92 (O_92,N_9874,N_9726);
and UO_93 (O_93,N_9688,N_9583);
nand UO_94 (O_94,N_9958,N_9642);
or UO_95 (O_95,N_9502,N_9521);
and UO_96 (O_96,N_9932,N_9869);
and UO_97 (O_97,N_9672,N_9553);
or UO_98 (O_98,N_9730,N_9901);
nor UO_99 (O_99,N_9809,N_9578);
nor UO_100 (O_100,N_9694,N_9873);
or UO_101 (O_101,N_9821,N_9580);
or UO_102 (O_102,N_9595,N_9924);
or UO_103 (O_103,N_9771,N_9766);
or UO_104 (O_104,N_9713,N_9916);
nand UO_105 (O_105,N_9652,N_9890);
and UO_106 (O_106,N_9882,N_9547);
nand UO_107 (O_107,N_9505,N_9784);
nor UO_108 (O_108,N_9923,N_9525);
or UO_109 (O_109,N_9915,N_9834);
nor UO_110 (O_110,N_9911,N_9764);
nor UO_111 (O_111,N_9931,N_9717);
and UO_112 (O_112,N_9830,N_9975);
and UO_113 (O_113,N_9712,N_9754);
nand UO_114 (O_114,N_9955,N_9598);
nor UO_115 (O_115,N_9831,N_9878);
nor UO_116 (O_116,N_9632,N_9978);
and UO_117 (O_117,N_9737,N_9936);
or UO_118 (O_118,N_9839,N_9881);
or UO_119 (O_119,N_9840,N_9945);
and UO_120 (O_120,N_9926,N_9938);
xor UO_121 (O_121,N_9753,N_9862);
nor UO_122 (O_122,N_9965,N_9540);
and UO_123 (O_123,N_9538,N_9817);
nand UO_124 (O_124,N_9522,N_9575);
or UO_125 (O_125,N_9819,N_9636);
nand UO_126 (O_126,N_9635,N_9531);
nor UO_127 (O_127,N_9996,N_9743);
nand UO_128 (O_128,N_9530,N_9990);
nor UO_129 (O_129,N_9933,N_9749);
or UO_130 (O_130,N_9528,N_9564);
nor UO_131 (O_131,N_9925,N_9518);
or UO_132 (O_132,N_9805,N_9993);
nand UO_133 (O_133,N_9777,N_9841);
or UO_134 (O_134,N_9559,N_9935);
or UO_135 (O_135,N_9967,N_9832);
nor UO_136 (O_136,N_9968,N_9893);
nor UO_137 (O_137,N_9820,N_9828);
nand UO_138 (O_138,N_9577,N_9889);
or UO_139 (O_139,N_9812,N_9748);
nand UO_140 (O_140,N_9879,N_9516);
nor UO_141 (O_141,N_9835,N_9829);
and UO_142 (O_142,N_9985,N_9675);
nor UO_143 (O_143,N_9704,N_9954);
or UO_144 (O_144,N_9630,N_9603);
nor UO_145 (O_145,N_9629,N_9859);
nand UO_146 (O_146,N_9908,N_9857);
nand UO_147 (O_147,N_9588,N_9648);
nor UO_148 (O_148,N_9980,N_9785);
xor UO_149 (O_149,N_9856,N_9708);
or UO_150 (O_150,N_9886,N_9943);
nor UO_151 (O_151,N_9561,N_9782);
nor UO_152 (O_152,N_9707,N_9858);
nor UO_153 (O_153,N_9581,N_9833);
nand UO_154 (O_154,N_9868,N_9853);
and UO_155 (O_155,N_9898,N_9909);
nor UO_156 (O_156,N_9724,N_9685);
and UO_157 (O_157,N_9607,N_9735);
or UO_158 (O_158,N_9666,N_9801);
xnor UO_159 (O_159,N_9847,N_9701);
or UO_160 (O_160,N_9673,N_9725);
nor UO_161 (O_161,N_9767,N_9710);
nor UO_162 (O_162,N_9551,N_9587);
nor UO_163 (O_163,N_9545,N_9729);
or UO_164 (O_164,N_9671,N_9746);
nand UO_165 (O_165,N_9683,N_9592);
and UO_166 (O_166,N_9699,N_9714);
nand UO_167 (O_167,N_9815,N_9689);
xor UO_168 (O_168,N_9599,N_9614);
nand UO_169 (O_169,N_9891,N_9608);
xor UO_170 (O_170,N_9940,N_9622);
nor UO_171 (O_171,N_9905,N_9779);
or UO_172 (O_172,N_9816,N_9920);
or UO_173 (O_173,N_9977,N_9727);
nand UO_174 (O_174,N_9887,N_9892);
nand UO_175 (O_175,N_9615,N_9877);
nand UO_176 (O_176,N_9971,N_9865);
or UO_177 (O_177,N_9514,N_9697);
or UO_178 (O_178,N_9507,N_9942);
and UO_179 (O_179,N_9626,N_9788);
nand UO_180 (O_180,N_9572,N_9904);
and UO_181 (O_181,N_9966,N_9957);
and UO_182 (O_182,N_9706,N_9655);
nand UO_183 (O_183,N_9768,N_9569);
nand UO_184 (O_184,N_9818,N_9541);
and UO_185 (O_185,N_9986,N_9772);
and UO_186 (O_186,N_9574,N_9872);
nor UO_187 (O_187,N_9529,N_9837);
nand UO_188 (O_188,N_9677,N_9861);
or UO_189 (O_189,N_9995,N_9798);
and UO_190 (O_190,N_9949,N_9695);
nand UO_191 (O_191,N_9827,N_9656);
or UO_192 (O_192,N_9597,N_9796);
and UO_193 (O_193,N_9774,N_9691);
and UO_194 (O_194,N_9752,N_9947);
and UO_195 (O_195,N_9969,N_9552);
and UO_196 (O_196,N_9870,N_9661);
xor UO_197 (O_197,N_9686,N_9951);
xor UO_198 (O_198,N_9546,N_9663);
nor UO_199 (O_199,N_9939,N_9848);
and UO_200 (O_200,N_9674,N_9692);
xor UO_201 (O_201,N_9807,N_9994);
and UO_202 (O_202,N_9804,N_9736);
or UO_203 (O_203,N_9740,N_9554);
and UO_204 (O_204,N_9972,N_9880);
and UO_205 (O_205,N_9761,N_9851);
and UO_206 (O_206,N_9501,N_9918);
nand UO_207 (O_207,N_9511,N_9567);
and UO_208 (O_208,N_9534,N_9982);
nand UO_209 (O_209,N_9751,N_9842);
nor UO_210 (O_210,N_9773,N_9823);
nand UO_211 (O_211,N_9802,N_9606);
xor UO_212 (O_212,N_9500,N_9590);
or UO_213 (O_213,N_9644,N_9983);
nand UO_214 (O_214,N_9741,N_9863);
nor UO_215 (O_215,N_9667,N_9845);
nand UO_216 (O_216,N_9711,N_9884);
or UO_217 (O_217,N_9846,N_9682);
and UO_218 (O_218,N_9702,N_9883);
nor UO_219 (O_219,N_9533,N_9852);
nand UO_220 (O_220,N_9602,N_9568);
or UO_221 (O_221,N_9733,N_9515);
nor UO_222 (O_222,N_9537,N_9976);
and UO_223 (O_223,N_9508,N_9952);
xnor UO_224 (O_224,N_9997,N_9783);
and UO_225 (O_225,N_9721,N_9718);
or UO_226 (O_226,N_9731,N_9956);
nand UO_227 (O_227,N_9813,N_9532);
and UO_228 (O_228,N_9616,N_9979);
and UO_229 (O_229,N_9503,N_9799);
or UO_230 (O_230,N_9658,N_9789);
nand UO_231 (O_231,N_9778,N_9653);
nand UO_232 (O_232,N_9716,N_9797);
nor UO_233 (O_233,N_9549,N_9526);
or UO_234 (O_234,N_9744,N_9573);
nand UO_235 (O_235,N_9535,N_9631);
nor UO_236 (O_236,N_9647,N_9760);
and UO_237 (O_237,N_9639,N_9849);
xor UO_238 (O_238,N_9669,N_9589);
and UO_239 (O_239,N_9739,N_9970);
and UO_240 (O_240,N_9543,N_9560);
and UO_241 (O_241,N_9888,N_9627);
and UO_242 (O_242,N_9709,N_9999);
or UO_243 (O_243,N_9814,N_9584);
or UO_244 (O_244,N_9585,N_9609);
nor UO_245 (O_245,N_9750,N_9860);
nand UO_246 (O_246,N_9506,N_9875);
nor UO_247 (O_247,N_9981,N_9634);
nor UO_248 (O_248,N_9991,N_9523);
nor UO_249 (O_249,N_9687,N_9509);
or UO_250 (O_250,N_9625,N_9707);
nand UO_251 (O_251,N_9905,N_9922);
nand UO_252 (O_252,N_9695,N_9705);
nand UO_253 (O_253,N_9909,N_9814);
nand UO_254 (O_254,N_9692,N_9893);
nand UO_255 (O_255,N_9670,N_9908);
and UO_256 (O_256,N_9849,N_9695);
nor UO_257 (O_257,N_9884,N_9535);
nand UO_258 (O_258,N_9692,N_9713);
nand UO_259 (O_259,N_9733,N_9898);
and UO_260 (O_260,N_9874,N_9629);
xor UO_261 (O_261,N_9809,N_9993);
or UO_262 (O_262,N_9604,N_9683);
nor UO_263 (O_263,N_9529,N_9783);
or UO_264 (O_264,N_9745,N_9696);
xnor UO_265 (O_265,N_9725,N_9867);
nor UO_266 (O_266,N_9984,N_9764);
or UO_267 (O_267,N_9686,N_9677);
nor UO_268 (O_268,N_9648,N_9696);
nor UO_269 (O_269,N_9523,N_9546);
and UO_270 (O_270,N_9771,N_9826);
or UO_271 (O_271,N_9674,N_9500);
xnor UO_272 (O_272,N_9844,N_9804);
nor UO_273 (O_273,N_9583,N_9962);
nor UO_274 (O_274,N_9608,N_9741);
nor UO_275 (O_275,N_9582,N_9576);
xnor UO_276 (O_276,N_9612,N_9711);
nand UO_277 (O_277,N_9850,N_9796);
nand UO_278 (O_278,N_9926,N_9540);
or UO_279 (O_279,N_9641,N_9887);
and UO_280 (O_280,N_9640,N_9665);
nor UO_281 (O_281,N_9852,N_9504);
or UO_282 (O_282,N_9823,N_9920);
or UO_283 (O_283,N_9574,N_9680);
and UO_284 (O_284,N_9604,N_9981);
nand UO_285 (O_285,N_9825,N_9774);
nand UO_286 (O_286,N_9938,N_9699);
nand UO_287 (O_287,N_9807,N_9509);
and UO_288 (O_288,N_9545,N_9918);
or UO_289 (O_289,N_9697,N_9531);
or UO_290 (O_290,N_9678,N_9959);
nand UO_291 (O_291,N_9777,N_9855);
or UO_292 (O_292,N_9738,N_9591);
xor UO_293 (O_293,N_9586,N_9621);
nand UO_294 (O_294,N_9976,N_9625);
and UO_295 (O_295,N_9500,N_9835);
nor UO_296 (O_296,N_9520,N_9615);
nand UO_297 (O_297,N_9857,N_9548);
nor UO_298 (O_298,N_9791,N_9557);
nor UO_299 (O_299,N_9529,N_9572);
nand UO_300 (O_300,N_9696,N_9915);
nor UO_301 (O_301,N_9557,N_9987);
and UO_302 (O_302,N_9519,N_9629);
and UO_303 (O_303,N_9981,N_9749);
and UO_304 (O_304,N_9646,N_9851);
and UO_305 (O_305,N_9599,N_9800);
nand UO_306 (O_306,N_9646,N_9838);
and UO_307 (O_307,N_9505,N_9779);
and UO_308 (O_308,N_9729,N_9531);
nand UO_309 (O_309,N_9964,N_9634);
xor UO_310 (O_310,N_9969,N_9648);
and UO_311 (O_311,N_9582,N_9850);
or UO_312 (O_312,N_9759,N_9601);
or UO_313 (O_313,N_9508,N_9959);
nor UO_314 (O_314,N_9728,N_9986);
or UO_315 (O_315,N_9652,N_9766);
or UO_316 (O_316,N_9712,N_9938);
nor UO_317 (O_317,N_9937,N_9855);
or UO_318 (O_318,N_9900,N_9597);
nand UO_319 (O_319,N_9612,N_9954);
and UO_320 (O_320,N_9926,N_9548);
or UO_321 (O_321,N_9935,N_9601);
and UO_322 (O_322,N_9906,N_9697);
or UO_323 (O_323,N_9513,N_9643);
or UO_324 (O_324,N_9734,N_9614);
nor UO_325 (O_325,N_9600,N_9671);
or UO_326 (O_326,N_9968,N_9943);
or UO_327 (O_327,N_9729,N_9857);
and UO_328 (O_328,N_9697,N_9937);
and UO_329 (O_329,N_9516,N_9537);
nor UO_330 (O_330,N_9631,N_9887);
xor UO_331 (O_331,N_9740,N_9643);
or UO_332 (O_332,N_9697,N_9783);
nand UO_333 (O_333,N_9521,N_9974);
nand UO_334 (O_334,N_9735,N_9618);
and UO_335 (O_335,N_9585,N_9727);
and UO_336 (O_336,N_9929,N_9735);
or UO_337 (O_337,N_9646,N_9684);
and UO_338 (O_338,N_9544,N_9797);
and UO_339 (O_339,N_9882,N_9536);
or UO_340 (O_340,N_9641,N_9605);
nor UO_341 (O_341,N_9831,N_9662);
nor UO_342 (O_342,N_9792,N_9579);
nand UO_343 (O_343,N_9588,N_9971);
xnor UO_344 (O_344,N_9963,N_9513);
nand UO_345 (O_345,N_9767,N_9693);
xnor UO_346 (O_346,N_9932,N_9988);
xnor UO_347 (O_347,N_9595,N_9789);
and UO_348 (O_348,N_9853,N_9604);
and UO_349 (O_349,N_9540,N_9623);
and UO_350 (O_350,N_9533,N_9944);
nor UO_351 (O_351,N_9805,N_9820);
nand UO_352 (O_352,N_9966,N_9993);
and UO_353 (O_353,N_9802,N_9970);
nand UO_354 (O_354,N_9788,N_9938);
nand UO_355 (O_355,N_9688,N_9921);
or UO_356 (O_356,N_9929,N_9713);
or UO_357 (O_357,N_9571,N_9813);
and UO_358 (O_358,N_9794,N_9608);
nor UO_359 (O_359,N_9761,N_9798);
or UO_360 (O_360,N_9782,N_9787);
and UO_361 (O_361,N_9930,N_9891);
xor UO_362 (O_362,N_9773,N_9675);
nor UO_363 (O_363,N_9663,N_9717);
nor UO_364 (O_364,N_9650,N_9989);
and UO_365 (O_365,N_9933,N_9864);
and UO_366 (O_366,N_9965,N_9759);
and UO_367 (O_367,N_9848,N_9990);
and UO_368 (O_368,N_9693,N_9805);
and UO_369 (O_369,N_9960,N_9638);
and UO_370 (O_370,N_9913,N_9762);
nand UO_371 (O_371,N_9649,N_9743);
xor UO_372 (O_372,N_9655,N_9614);
nand UO_373 (O_373,N_9843,N_9950);
nor UO_374 (O_374,N_9979,N_9674);
and UO_375 (O_375,N_9989,N_9628);
nor UO_376 (O_376,N_9611,N_9879);
or UO_377 (O_377,N_9521,N_9780);
xor UO_378 (O_378,N_9776,N_9903);
or UO_379 (O_379,N_9885,N_9587);
or UO_380 (O_380,N_9965,N_9877);
or UO_381 (O_381,N_9843,N_9769);
or UO_382 (O_382,N_9637,N_9555);
and UO_383 (O_383,N_9542,N_9705);
nor UO_384 (O_384,N_9680,N_9900);
and UO_385 (O_385,N_9811,N_9702);
nand UO_386 (O_386,N_9784,N_9672);
nand UO_387 (O_387,N_9758,N_9525);
nand UO_388 (O_388,N_9884,N_9894);
nor UO_389 (O_389,N_9669,N_9630);
nor UO_390 (O_390,N_9582,N_9698);
xnor UO_391 (O_391,N_9944,N_9588);
and UO_392 (O_392,N_9819,N_9794);
or UO_393 (O_393,N_9536,N_9716);
nand UO_394 (O_394,N_9882,N_9716);
nand UO_395 (O_395,N_9655,N_9578);
and UO_396 (O_396,N_9511,N_9839);
nor UO_397 (O_397,N_9820,N_9585);
and UO_398 (O_398,N_9835,N_9605);
and UO_399 (O_399,N_9830,N_9928);
or UO_400 (O_400,N_9865,N_9947);
nor UO_401 (O_401,N_9837,N_9700);
nor UO_402 (O_402,N_9674,N_9744);
nor UO_403 (O_403,N_9692,N_9823);
or UO_404 (O_404,N_9722,N_9822);
or UO_405 (O_405,N_9710,N_9956);
nand UO_406 (O_406,N_9792,N_9610);
nand UO_407 (O_407,N_9555,N_9959);
and UO_408 (O_408,N_9773,N_9913);
nor UO_409 (O_409,N_9557,N_9647);
nand UO_410 (O_410,N_9637,N_9757);
xnor UO_411 (O_411,N_9706,N_9801);
or UO_412 (O_412,N_9570,N_9878);
and UO_413 (O_413,N_9554,N_9737);
nor UO_414 (O_414,N_9869,N_9673);
nor UO_415 (O_415,N_9739,N_9507);
and UO_416 (O_416,N_9539,N_9710);
xor UO_417 (O_417,N_9563,N_9586);
and UO_418 (O_418,N_9997,N_9931);
nor UO_419 (O_419,N_9755,N_9932);
and UO_420 (O_420,N_9734,N_9842);
nand UO_421 (O_421,N_9793,N_9602);
or UO_422 (O_422,N_9790,N_9617);
nand UO_423 (O_423,N_9746,N_9855);
or UO_424 (O_424,N_9801,N_9559);
nor UO_425 (O_425,N_9520,N_9786);
or UO_426 (O_426,N_9699,N_9572);
nand UO_427 (O_427,N_9601,N_9852);
or UO_428 (O_428,N_9738,N_9645);
xnor UO_429 (O_429,N_9992,N_9715);
nor UO_430 (O_430,N_9684,N_9694);
and UO_431 (O_431,N_9637,N_9727);
nor UO_432 (O_432,N_9567,N_9694);
nor UO_433 (O_433,N_9944,N_9917);
and UO_434 (O_434,N_9622,N_9883);
or UO_435 (O_435,N_9525,N_9824);
or UO_436 (O_436,N_9856,N_9652);
xnor UO_437 (O_437,N_9558,N_9510);
nand UO_438 (O_438,N_9780,N_9674);
and UO_439 (O_439,N_9613,N_9769);
nand UO_440 (O_440,N_9809,N_9515);
and UO_441 (O_441,N_9501,N_9854);
or UO_442 (O_442,N_9611,N_9888);
and UO_443 (O_443,N_9986,N_9793);
or UO_444 (O_444,N_9754,N_9599);
or UO_445 (O_445,N_9710,N_9919);
xor UO_446 (O_446,N_9988,N_9505);
nand UO_447 (O_447,N_9624,N_9869);
or UO_448 (O_448,N_9544,N_9854);
nor UO_449 (O_449,N_9769,N_9840);
nor UO_450 (O_450,N_9539,N_9887);
and UO_451 (O_451,N_9818,N_9894);
and UO_452 (O_452,N_9942,N_9947);
xor UO_453 (O_453,N_9677,N_9792);
nand UO_454 (O_454,N_9997,N_9642);
nor UO_455 (O_455,N_9896,N_9573);
and UO_456 (O_456,N_9992,N_9699);
or UO_457 (O_457,N_9542,N_9928);
nor UO_458 (O_458,N_9575,N_9989);
or UO_459 (O_459,N_9904,N_9820);
nand UO_460 (O_460,N_9547,N_9542);
and UO_461 (O_461,N_9783,N_9756);
nor UO_462 (O_462,N_9787,N_9519);
and UO_463 (O_463,N_9650,N_9843);
nor UO_464 (O_464,N_9530,N_9729);
or UO_465 (O_465,N_9629,N_9510);
and UO_466 (O_466,N_9763,N_9911);
nand UO_467 (O_467,N_9956,N_9938);
nor UO_468 (O_468,N_9994,N_9648);
nand UO_469 (O_469,N_9826,N_9790);
or UO_470 (O_470,N_9682,N_9694);
xor UO_471 (O_471,N_9750,N_9832);
and UO_472 (O_472,N_9958,N_9866);
and UO_473 (O_473,N_9773,N_9910);
nand UO_474 (O_474,N_9806,N_9945);
and UO_475 (O_475,N_9569,N_9903);
or UO_476 (O_476,N_9695,N_9505);
xnor UO_477 (O_477,N_9950,N_9655);
nor UO_478 (O_478,N_9808,N_9794);
nor UO_479 (O_479,N_9885,N_9561);
nor UO_480 (O_480,N_9657,N_9731);
xor UO_481 (O_481,N_9994,N_9929);
or UO_482 (O_482,N_9976,N_9695);
nor UO_483 (O_483,N_9588,N_9771);
xnor UO_484 (O_484,N_9722,N_9678);
and UO_485 (O_485,N_9713,N_9617);
xor UO_486 (O_486,N_9804,N_9530);
and UO_487 (O_487,N_9901,N_9715);
or UO_488 (O_488,N_9638,N_9593);
and UO_489 (O_489,N_9970,N_9539);
nand UO_490 (O_490,N_9570,N_9911);
nor UO_491 (O_491,N_9664,N_9931);
xor UO_492 (O_492,N_9575,N_9981);
nand UO_493 (O_493,N_9689,N_9796);
or UO_494 (O_494,N_9802,N_9777);
nand UO_495 (O_495,N_9921,N_9540);
nor UO_496 (O_496,N_9988,N_9601);
and UO_497 (O_497,N_9875,N_9833);
or UO_498 (O_498,N_9717,N_9741);
and UO_499 (O_499,N_9947,N_9803);
nand UO_500 (O_500,N_9614,N_9969);
and UO_501 (O_501,N_9672,N_9998);
nor UO_502 (O_502,N_9775,N_9999);
nor UO_503 (O_503,N_9526,N_9942);
or UO_504 (O_504,N_9922,N_9621);
and UO_505 (O_505,N_9822,N_9960);
or UO_506 (O_506,N_9762,N_9888);
and UO_507 (O_507,N_9749,N_9641);
or UO_508 (O_508,N_9674,N_9769);
and UO_509 (O_509,N_9607,N_9538);
and UO_510 (O_510,N_9694,N_9977);
or UO_511 (O_511,N_9903,N_9828);
or UO_512 (O_512,N_9686,N_9864);
or UO_513 (O_513,N_9508,N_9501);
or UO_514 (O_514,N_9644,N_9759);
nand UO_515 (O_515,N_9899,N_9958);
or UO_516 (O_516,N_9655,N_9807);
xnor UO_517 (O_517,N_9697,N_9688);
and UO_518 (O_518,N_9705,N_9978);
xnor UO_519 (O_519,N_9521,N_9618);
or UO_520 (O_520,N_9814,N_9741);
nor UO_521 (O_521,N_9783,N_9785);
nor UO_522 (O_522,N_9848,N_9884);
nand UO_523 (O_523,N_9708,N_9892);
and UO_524 (O_524,N_9939,N_9511);
and UO_525 (O_525,N_9965,N_9652);
nand UO_526 (O_526,N_9542,N_9529);
nor UO_527 (O_527,N_9767,N_9636);
nor UO_528 (O_528,N_9597,N_9607);
and UO_529 (O_529,N_9985,N_9504);
or UO_530 (O_530,N_9857,N_9708);
or UO_531 (O_531,N_9509,N_9976);
nor UO_532 (O_532,N_9592,N_9517);
nand UO_533 (O_533,N_9751,N_9860);
nand UO_534 (O_534,N_9964,N_9962);
and UO_535 (O_535,N_9738,N_9699);
xor UO_536 (O_536,N_9986,N_9669);
or UO_537 (O_537,N_9585,N_9797);
or UO_538 (O_538,N_9851,N_9954);
or UO_539 (O_539,N_9758,N_9526);
nand UO_540 (O_540,N_9764,N_9544);
nand UO_541 (O_541,N_9765,N_9654);
nor UO_542 (O_542,N_9731,N_9973);
xor UO_543 (O_543,N_9745,N_9684);
nand UO_544 (O_544,N_9743,N_9807);
and UO_545 (O_545,N_9852,N_9813);
nand UO_546 (O_546,N_9951,N_9847);
or UO_547 (O_547,N_9514,N_9802);
nor UO_548 (O_548,N_9736,N_9787);
or UO_549 (O_549,N_9679,N_9730);
and UO_550 (O_550,N_9510,N_9537);
nand UO_551 (O_551,N_9683,N_9630);
xnor UO_552 (O_552,N_9778,N_9563);
or UO_553 (O_553,N_9799,N_9899);
nor UO_554 (O_554,N_9786,N_9542);
nand UO_555 (O_555,N_9628,N_9856);
nand UO_556 (O_556,N_9868,N_9956);
xnor UO_557 (O_557,N_9809,N_9692);
or UO_558 (O_558,N_9621,N_9575);
and UO_559 (O_559,N_9921,N_9526);
and UO_560 (O_560,N_9644,N_9698);
xnor UO_561 (O_561,N_9587,N_9684);
nor UO_562 (O_562,N_9766,N_9840);
nor UO_563 (O_563,N_9853,N_9923);
nor UO_564 (O_564,N_9941,N_9546);
nand UO_565 (O_565,N_9723,N_9882);
and UO_566 (O_566,N_9543,N_9642);
nor UO_567 (O_567,N_9999,N_9853);
and UO_568 (O_568,N_9916,N_9632);
and UO_569 (O_569,N_9654,N_9985);
nand UO_570 (O_570,N_9597,N_9892);
and UO_571 (O_571,N_9803,N_9858);
nand UO_572 (O_572,N_9673,N_9710);
xnor UO_573 (O_573,N_9679,N_9542);
and UO_574 (O_574,N_9938,N_9654);
nand UO_575 (O_575,N_9504,N_9662);
xnor UO_576 (O_576,N_9561,N_9975);
nand UO_577 (O_577,N_9984,N_9515);
or UO_578 (O_578,N_9832,N_9629);
or UO_579 (O_579,N_9716,N_9935);
xnor UO_580 (O_580,N_9851,N_9887);
and UO_581 (O_581,N_9734,N_9907);
xor UO_582 (O_582,N_9837,N_9738);
nor UO_583 (O_583,N_9832,N_9740);
and UO_584 (O_584,N_9619,N_9971);
or UO_585 (O_585,N_9709,N_9690);
or UO_586 (O_586,N_9583,N_9859);
or UO_587 (O_587,N_9858,N_9890);
or UO_588 (O_588,N_9569,N_9541);
or UO_589 (O_589,N_9806,N_9666);
or UO_590 (O_590,N_9829,N_9978);
or UO_591 (O_591,N_9937,N_9604);
nor UO_592 (O_592,N_9685,N_9934);
xor UO_593 (O_593,N_9587,N_9803);
or UO_594 (O_594,N_9879,N_9768);
or UO_595 (O_595,N_9783,N_9668);
xnor UO_596 (O_596,N_9645,N_9876);
and UO_597 (O_597,N_9700,N_9724);
nand UO_598 (O_598,N_9711,N_9947);
nor UO_599 (O_599,N_9700,N_9806);
or UO_600 (O_600,N_9830,N_9604);
nor UO_601 (O_601,N_9775,N_9547);
and UO_602 (O_602,N_9623,N_9598);
nand UO_603 (O_603,N_9921,N_9605);
or UO_604 (O_604,N_9843,N_9512);
and UO_605 (O_605,N_9586,N_9769);
or UO_606 (O_606,N_9681,N_9619);
nor UO_607 (O_607,N_9702,N_9813);
and UO_608 (O_608,N_9593,N_9756);
or UO_609 (O_609,N_9822,N_9760);
or UO_610 (O_610,N_9608,N_9827);
nor UO_611 (O_611,N_9611,N_9989);
and UO_612 (O_612,N_9991,N_9558);
nor UO_613 (O_613,N_9769,N_9638);
and UO_614 (O_614,N_9604,N_9515);
nand UO_615 (O_615,N_9874,N_9630);
or UO_616 (O_616,N_9647,N_9976);
nor UO_617 (O_617,N_9903,N_9964);
and UO_618 (O_618,N_9814,N_9938);
nand UO_619 (O_619,N_9842,N_9848);
nor UO_620 (O_620,N_9728,N_9891);
nor UO_621 (O_621,N_9629,N_9977);
nand UO_622 (O_622,N_9759,N_9531);
nand UO_623 (O_623,N_9944,N_9728);
or UO_624 (O_624,N_9553,N_9884);
nand UO_625 (O_625,N_9672,N_9616);
xor UO_626 (O_626,N_9992,N_9607);
nor UO_627 (O_627,N_9821,N_9552);
and UO_628 (O_628,N_9559,N_9525);
nand UO_629 (O_629,N_9847,N_9518);
nor UO_630 (O_630,N_9718,N_9832);
or UO_631 (O_631,N_9758,N_9746);
nor UO_632 (O_632,N_9659,N_9858);
and UO_633 (O_633,N_9852,N_9606);
or UO_634 (O_634,N_9654,N_9866);
xor UO_635 (O_635,N_9726,N_9627);
nand UO_636 (O_636,N_9889,N_9637);
nor UO_637 (O_637,N_9518,N_9586);
or UO_638 (O_638,N_9807,N_9658);
nor UO_639 (O_639,N_9850,N_9947);
nor UO_640 (O_640,N_9861,N_9868);
xnor UO_641 (O_641,N_9786,N_9554);
or UO_642 (O_642,N_9960,N_9753);
or UO_643 (O_643,N_9632,N_9882);
xor UO_644 (O_644,N_9618,N_9560);
and UO_645 (O_645,N_9837,N_9606);
xor UO_646 (O_646,N_9728,N_9933);
xor UO_647 (O_647,N_9885,N_9818);
nor UO_648 (O_648,N_9535,N_9842);
xnor UO_649 (O_649,N_9593,N_9519);
xor UO_650 (O_650,N_9560,N_9862);
nand UO_651 (O_651,N_9671,N_9651);
nand UO_652 (O_652,N_9969,N_9941);
xnor UO_653 (O_653,N_9834,N_9789);
and UO_654 (O_654,N_9768,N_9889);
and UO_655 (O_655,N_9645,N_9879);
xnor UO_656 (O_656,N_9694,N_9520);
xnor UO_657 (O_657,N_9564,N_9633);
nor UO_658 (O_658,N_9663,N_9794);
nand UO_659 (O_659,N_9618,N_9975);
and UO_660 (O_660,N_9648,N_9991);
and UO_661 (O_661,N_9787,N_9757);
nand UO_662 (O_662,N_9827,N_9536);
nor UO_663 (O_663,N_9595,N_9632);
and UO_664 (O_664,N_9674,N_9966);
nor UO_665 (O_665,N_9984,N_9646);
nor UO_666 (O_666,N_9611,N_9789);
nor UO_667 (O_667,N_9595,N_9777);
nand UO_668 (O_668,N_9519,N_9729);
or UO_669 (O_669,N_9634,N_9759);
nor UO_670 (O_670,N_9817,N_9749);
nand UO_671 (O_671,N_9544,N_9855);
or UO_672 (O_672,N_9538,N_9804);
nor UO_673 (O_673,N_9957,N_9858);
and UO_674 (O_674,N_9827,N_9516);
nand UO_675 (O_675,N_9722,N_9702);
or UO_676 (O_676,N_9982,N_9883);
or UO_677 (O_677,N_9842,N_9572);
nor UO_678 (O_678,N_9719,N_9767);
nor UO_679 (O_679,N_9856,N_9584);
nand UO_680 (O_680,N_9603,N_9745);
nand UO_681 (O_681,N_9773,N_9683);
nor UO_682 (O_682,N_9776,N_9565);
nand UO_683 (O_683,N_9986,N_9997);
or UO_684 (O_684,N_9538,N_9792);
xor UO_685 (O_685,N_9591,N_9580);
or UO_686 (O_686,N_9640,N_9696);
xor UO_687 (O_687,N_9538,N_9710);
and UO_688 (O_688,N_9611,N_9672);
or UO_689 (O_689,N_9685,N_9811);
or UO_690 (O_690,N_9904,N_9643);
nand UO_691 (O_691,N_9834,N_9872);
and UO_692 (O_692,N_9782,N_9770);
nand UO_693 (O_693,N_9939,N_9669);
nor UO_694 (O_694,N_9562,N_9815);
nand UO_695 (O_695,N_9577,N_9511);
nand UO_696 (O_696,N_9709,N_9678);
or UO_697 (O_697,N_9581,N_9836);
xnor UO_698 (O_698,N_9984,N_9728);
nand UO_699 (O_699,N_9713,N_9664);
nor UO_700 (O_700,N_9614,N_9563);
and UO_701 (O_701,N_9759,N_9901);
or UO_702 (O_702,N_9557,N_9707);
nor UO_703 (O_703,N_9685,N_9997);
nor UO_704 (O_704,N_9997,N_9554);
nand UO_705 (O_705,N_9882,N_9902);
nand UO_706 (O_706,N_9856,N_9820);
and UO_707 (O_707,N_9910,N_9588);
xor UO_708 (O_708,N_9725,N_9963);
nand UO_709 (O_709,N_9969,N_9841);
or UO_710 (O_710,N_9818,N_9511);
nand UO_711 (O_711,N_9943,N_9561);
xor UO_712 (O_712,N_9975,N_9603);
or UO_713 (O_713,N_9675,N_9792);
nand UO_714 (O_714,N_9897,N_9552);
or UO_715 (O_715,N_9989,N_9976);
nor UO_716 (O_716,N_9700,N_9989);
or UO_717 (O_717,N_9970,N_9667);
and UO_718 (O_718,N_9888,N_9703);
nand UO_719 (O_719,N_9831,N_9567);
and UO_720 (O_720,N_9637,N_9791);
nor UO_721 (O_721,N_9847,N_9629);
nor UO_722 (O_722,N_9648,N_9504);
or UO_723 (O_723,N_9988,N_9763);
nand UO_724 (O_724,N_9558,N_9738);
and UO_725 (O_725,N_9655,N_9724);
and UO_726 (O_726,N_9948,N_9625);
or UO_727 (O_727,N_9960,N_9903);
nand UO_728 (O_728,N_9507,N_9706);
and UO_729 (O_729,N_9705,N_9877);
and UO_730 (O_730,N_9524,N_9972);
and UO_731 (O_731,N_9966,N_9917);
nand UO_732 (O_732,N_9649,N_9871);
nor UO_733 (O_733,N_9527,N_9975);
nand UO_734 (O_734,N_9670,N_9564);
or UO_735 (O_735,N_9674,N_9627);
nand UO_736 (O_736,N_9565,N_9993);
and UO_737 (O_737,N_9525,N_9718);
xor UO_738 (O_738,N_9834,N_9712);
and UO_739 (O_739,N_9572,N_9669);
or UO_740 (O_740,N_9634,N_9508);
and UO_741 (O_741,N_9649,N_9959);
or UO_742 (O_742,N_9652,N_9802);
nand UO_743 (O_743,N_9986,N_9690);
and UO_744 (O_744,N_9862,N_9576);
nand UO_745 (O_745,N_9599,N_9925);
nand UO_746 (O_746,N_9983,N_9778);
nand UO_747 (O_747,N_9618,N_9723);
or UO_748 (O_748,N_9994,N_9928);
or UO_749 (O_749,N_9970,N_9817);
and UO_750 (O_750,N_9536,N_9818);
and UO_751 (O_751,N_9626,N_9631);
or UO_752 (O_752,N_9995,N_9665);
or UO_753 (O_753,N_9987,N_9795);
nand UO_754 (O_754,N_9523,N_9560);
nor UO_755 (O_755,N_9733,N_9530);
and UO_756 (O_756,N_9720,N_9652);
and UO_757 (O_757,N_9980,N_9802);
or UO_758 (O_758,N_9577,N_9777);
xor UO_759 (O_759,N_9810,N_9841);
xor UO_760 (O_760,N_9535,N_9663);
and UO_761 (O_761,N_9625,N_9634);
nor UO_762 (O_762,N_9606,N_9703);
nor UO_763 (O_763,N_9558,N_9526);
nor UO_764 (O_764,N_9601,N_9673);
nand UO_765 (O_765,N_9646,N_9629);
nor UO_766 (O_766,N_9903,N_9861);
or UO_767 (O_767,N_9812,N_9791);
nand UO_768 (O_768,N_9670,N_9657);
nand UO_769 (O_769,N_9625,N_9880);
or UO_770 (O_770,N_9573,N_9660);
nor UO_771 (O_771,N_9566,N_9827);
xor UO_772 (O_772,N_9986,N_9857);
and UO_773 (O_773,N_9708,N_9993);
nor UO_774 (O_774,N_9844,N_9505);
nand UO_775 (O_775,N_9727,N_9846);
nor UO_776 (O_776,N_9663,N_9792);
or UO_777 (O_777,N_9867,N_9729);
nand UO_778 (O_778,N_9826,N_9527);
and UO_779 (O_779,N_9829,N_9553);
nand UO_780 (O_780,N_9512,N_9897);
or UO_781 (O_781,N_9696,N_9769);
nand UO_782 (O_782,N_9717,N_9675);
nor UO_783 (O_783,N_9611,N_9754);
nor UO_784 (O_784,N_9923,N_9939);
nand UO_785 (O_785,N_9928,N_9657);
or UO_786 (O_786,N_9587,N_9513);
nor UO_787 (O_787,N_9964,N_9778);
or UO_788 (O_788,N_9963,N_9530);
nand UO_789 (O_789,N_9747,N_9906);
nand UO_790 (O_790,N_9802,N_9742);
nor UO_791 (O_791,N_9607,N_9823);
nand UO_792 (O_792,N_9797,N_9803);
or UO_793 (O_793,N_9532,N_9503);
nor UO_794 (O_794,N_9895,N_9872);
nor UO_795 (O_795,N_9769,N_9882);
nor UO_796 (O_796,N_9752,N_9521);
xor UO_797 (O_797,N_9779,N_9623);
and UO_798 (O_798,N_9706,N_9992);
or UO_799 (O_799,N_9729,N_9778);
and UO_800 (O_800,N_9653,N_9624);
nor UO_801 (O_801,N_9967,N_9560);
xor UO_802 (O_802,N_9972,N_9500);
nor UO_803 (O_803,N_9643,N_9649);
and UO_804 (O_804,N_9770,N_9517);
xor UO_805 (O_805,N_9594,N_9577);
or UO_806 (O_806,N_9598,N_9831);
nor UO_807 (O_807,N_9652,N_9664);
nand UO_808 (O_808,N_9982,N_9629);
nand UO_809 (O_809,N_9521,N_9756);
or UO_810 (O_810,N_9749,N_9566);
nand UO_811 (O_811,N_9778,N_9880);
xor UO_812 (O_812,N_9562,N_9537);
and UO_813 (O_813,N_9757,N_9884);
nand UO_814 (O_814,N_9671,N_9857);
or UO_815 (O_815,N_9907,N_9636);
or UO_816 (O_816,N_9983,N_9836);
nor UO_817 (O_817,N_9547,N_9883);
and UO_818 (O_818,N_9532,N_9818);
nor UO_819 (O_819,N_9516,N_9836);
nor UO_820 (O_820,N_9680,N_9501);
xor UO_821 (O_821,N_9963,N_9907);
or UO_822 (O_822,N_9863,N_9720);
or UO_823 (O_823,N_9936,N_9538);
nand UO_824 (O_824,N_9656,N_9538);
xnor UO_825 (O_825,N_9854,N_9744);
and UO_826 (O_826,N_9638,N_9604);
nand UO_827 (O_827,N_9725,N_9508);
nor UO_828 (O_828,N_9859,N_9594);
and UO_829 (O_829,N_9938,N_9907);
or UO_830 (O_830,N_9553,N_9659);
xor UO_831 (O_831,N_9937,N_9997);
nor UO_832 (O_832,N_9618,N_9682);
nor UO_833 (O_833,N_9698,N_9771);
or UO_834 (O_834,N_9752,N_9720);
nand UO_835 (O_835,N_9602,N_9899);
and UO_836 (O_836,N_9824,N_9586);
and UO_837 (O_837,N_9697,N_9655);
or UO_838 (O_838,N_9638,N_9714);
xor UO_839 (O_839,N_9963,N_9591);
nand UO_840 (O_840,N_9553,N_9931);
and UO_841 (O_841,N_9959,N_9602);
and UO_842 (O_842,N_9704,N_9619);
or UO_843 (O_843,N_9666,N_9561);
nor UO_844 (O_844,N_9780,N_9858);
nor UO_845 (O_845,N_9729,N_9511);
nor UO_846 (O_846,N_9561,N_9783);
or UO_847 (O_847,N_9850,N_9959);
nor UO_848 (O_848,N_9882,N_9510);
and UO_849 (O_849,N_9646,N_9675);
and UO_850 (O_850,N_9845,N_9774);
and UO_851 (O_851,N_9568,N_9692);
and UO_852 (O_852,N_9577,N_9856);
nor UO_853 (O_853,N_9756,N_9682);
nand UO_854 (O_854,N_9527,N_9849);
nand UO_855 (O_855,N_9698,N_9858);
or UO_856 (O_856,N_9526,N_9716);
and UO_857 (O_857,N_9631,N_9736);
nand UO_858 (O_858,N_9936,N_9954);
and UO_859 (O_859,N_9605,N_9527);
or UO_860 (O_860,N_9829,N_9736);
or UO_861 (O_861,N_9684,N_9632);
nand UO_862 (O_862,N_9691,N_9965);
xor UO_863 (O_863,N_9997,N_9755);
and UO_864 (O_864,N_9639,N_9809);
xnor UO_865 (O_865,N_9774,N_9626);
nor UO_866 (O_866,N_9759,N_9959);
or UO_867 (O_867,N_9696,N_9901);
and UO_868 (O_868,N_9772,N_9894);
nor UO_869 (O_869,N_9922,N_9855);
nor UO_870 (O_870,N_9916,N_9623);
nor UO_871 (O_871,N_9822,N_9504);
nor UO_872 (O_872,N_9714,N_9592);
nand UO_873 (O_873,N_9525,N_9789);
nand UO_874 (O_874,N_9638,N_9870);
and UO_875 (O_875,N_9527,N_9623);
and UO_876 (O_876,N_9625,N_9724);
nor UO_877 (O_877,N_9954,N_9590);
and UO_878 (O_878,N_9511,N_9521);
or UO_879 (O_879,N_9678,N_9715);
nand UO_880 (O_880,N_9626,N_9802);
nor UO_881 (O_881,N_9938,N_9668);
nand UO_882 (O_882,N_9781,N_9597);
nand UO_883 (O_883,N_9677,N_9510);
and UO_884 (O_884,N_9831,N_9875);
and UO_885 (O_885,N_9774,N_9767);
and UO_886 (O_886,N_9886,N_9858);
xnor UO_887 (O_887,N_9586,N_9967);
xnor UO_888 (O_888,N_9961,N_9670);
or UO_889 (O_889,N_9942,N_9913);
or UO_890 (O_890,N_9740,N_9820);
nand UO_891 (O_891,N_9906,N_9604);
nand UO_892 (O_892,N_9999,N_9650);
and UO_893 (O_893,N_9552,N_9850);
or UO_894 (O_894,N_9598,N_9930);
and UO_895 (O_895,N_9623,N_9909);
or UO_896 (O_896,N_9745,N_9722);
or UO_897 (O_897,N_9931,N_9518);
or UO_898 (O_898,N_9779,N_9929);
xor UO_899 (O_899,N_9954,N_9648);
nand UO_900 (O_900,N_9612,N_9931);
and UO_901 (O_901,N_9609,N_9680);
nand UO_902 (O_902,N_9504,N_9671);
or UO_903 (O_903,N_9772,N_9784);
and UO_904 (O_904,N_9670,N_9890);
nor UO_905 (O_905,N_9697,N_9574);
or UO_906 (O_906,N_9851,N_9692);
and UO_907 (O_907,N_9620,N_9515);
and UO_908 (O_908,N_9982,N_9584);
or UO_909 (O_909,N_9883,N_9520);
and UO_910 (O_910,N_9709,N_9965);
nand UO_911 (O_911,N_9864,N_9887);
or UO_912 (O_912,N_9856,N_9731);
nand UO_913 (O_913,N_9952,N_9903);
nor UO_914 (O_914,N_9880,N_9744);
or UO_915 (O_915,N_9660,N_9832);
or UO_916 (O_916,N_9841,N_9564);
nand UO_917 (O_917,N_9510,N_9614);
and UO_918 (O_918,N_9684,N_9907);
nand UO_919 (O_919,N_9617,N_9921);
nand UO_920 (O_920,N_9654,N_9885);
and UO_921 (O_921,N_9564,N_9809);
nand UO_922 (O_922,N_9621,N_9971);
xnor UO_923 (O_923,N_9938,N_9695);
and UO_924 (O_924,N_9773,N_9998);
nor UO_925 (O_925,N_9820,N_9881);
or UO_926 (O_926,N_9615,N_9957);
or UO_927 (O_927,N_9973,N_9992);
nand UO_928 (O_928,N_9570,N_9680);
nor UO_929 (O_929,N_9801,N_9970);
nand UO_930 (O_930,N_9933,N_9502);
nor UO_931 (O_931,N_9511,N_9887);
xnor UO_932 (O_932,N_9573,N_9796);
nor UO_933 (O_933,N_9874,N_9503);
and UO_934 (O_934,N_9974,N_9752);
and UO_935 (O_935,N_9567,N_9941);
xnor UO_936 (O_936,N_9978,N_9899);
nand UO_937 (O_937,N_9823,N_9660);
or UO_938 (O_938,N_9896,N_9894);
nand UO_939 (O_939,N_9990,N_9659);
nor UO_940 (O_940,N_9764,N_9733);
and UO_941 (O_941,N_9802,N_9502);
nor UO_942 (O_942,N_9981,N_9720);
nand UO_943 (O_943,N_9662,N_9648);
or UO_944 (O_944,N_9609,N_9927);
xor UO_945 (O_945,N_9742,N_9983);
nor UO_946 (O_946,N_9545,N_9720);
and UO_947 (O_947,N_9981,N_9853);
nand UO_948 (O_948,N_9939,N_9731);
or UO_949 (O_949,N_9836,N_9695);
nor UO_950 (O_950,N_9875,N_9827);
nor UO_951 (O_951,N_9613,N_9747);
and UO_952 (O_952,N_9995,N_9625);
nand UO_953 (O_953,N_9894,N_9640);
nand UO_954 (O_954,N_9691,N_9596);
nand UO_955 (O_955,N_9841,N_9636);
nand UO_956 (O_956,N_9553,N_9869);
nor UO_957 (O_957,N_9742,N_9511);
or UO_958 (O_958,N_9771,N_9668);
xor UO_959 (O_959,N_9685,N_9757);
nor UO_960 (O_960,N_9683,N_9984);
or UO_961 (O_961,N_9778,N_9662);
xor UO_962 (O_962,N_9504,N_9930);
and UO_963 (O_963,N_9659,N_9721);
nand UO_964 (O_964,N_9645,N_9715);
xnor UO_965 (O_965,N_9598,N_9770);
and UO_966 (O_966,N_9807,N_9766);
nand UO_967 (O_967,N_9934,N_9577);
nand UO_968 (O_968,N_9736,N_9644);
nand UO_969 (O_969,N_9714,N_9907);
nor UO_970 (O_970,N_9805,N_9764);
or UO_971 (O_971,N_9523,N_9974);
xor UO_972 (O_972,N_9881,N_9558);
nor UO_973 (O_973,N_9807,N_9970);
nand UO_974 (O_974,N_9937,N_9965);
and UO_975 (O_975,N_9808,N_9584);
nor UO_976 (O_976,N_9630,N_9518);
nor UO_977 (O_977,N_9801,N_9797);
or UO_978 (O_978,N_9507,N_9884);
or UO_979 (O_979,N_9902,N_9706);
and UO_980 (O_980,N_9835,N_9928);
nand UO_981 (O_981,N_9887,N_9741);
nor UO_982 (O_982,N_9761,N_9967);
xnor UO_983 (O_983,N_9747,N_9860);
or UO_984 (O_984,N_9782,N_9748);
nand UO_985 (O_985,N_9579,N_9647);
or UO_986 (O_986,N_9604,N_9949);
and UO_987 (O_987,N_9968,N_9629);
and UO_988 (O_988,N_9713,N_9944);
nor UO_989 (O_989,N_9547,N_9908);
or UO_990 (O_990,N_9966,N_9697);
nor UO_991 (O_991,N_9957,N_9648);
nand UO_992 (O_992,N_9747,N_9833);
nand UO_993 (O_993,N_9958,N_9525);
and UO_994 (O_994,N_9679,N_9919);
or UO_995 (O_995,N_9547,N_9594);
and UO_996 (O_996,N_9759,N_9663);
and UO_997 (O_997,N_9876,N_9934);
nand UO_998 (O_998,N_9700,N_9976);
or UO_999 (O_999,N_9534,N_9600);
and UO_1000 (O_1000,N_9764,N_9695);
or UO_1001 (O_1001,N_9792,N_9894);
or UO_1002 (O_1002,N_9711,N_9886);
or UO_1003 (O_1003,N_9860,N_9531);
or UO_1004 (O_1004,N_9781,N_9579);
nand UO_1005 (O_1005,N_9652,N_9659);
or UO_1006 (O_1006,N_9523,N_9683);
xor UO_1007 (O_1007,N_9561,N_9727);
and UO_1008 (O_1008,N_9755,N_9782);
nand UO_1009 (O_1009,N_9920,N_9835);
nand UO_1010 (O_1010,N_9721,N_9600);
and UO_1011 (O_1011,N_9592,N_9633);
and UO_1012 (O_1012,N_9847,N_9952);
and UO_1013 (O_1013,N_9909,N_9902);
and UO_1014 (O_1014,N_9736,N_9803);
xnor UO_1015 (O_1015,N_9869,N_9997);
and UO_1016 (O_1016,N_9727,N_9521);
and UO_1017 (O_1017,N_9762,N_9797);
and UO_1018 (O_1018,N_9891,N_9949);
or UO_1019 (O_1019,N_9950,N_9794);
and UO_1020 (O_1020,N_9621,N_9690);
nand UO_1021 (O_1021,N_9942,N_9594);
nand UO_1022 (O_1022,N_9667,N_9985);
nor UO_1023 (O_1023,N_9618,N_9603);
nor UO_1024 (O_1024,N_9517,N_9835);
and UO_1025 (O_1025,N_9684,N_9887);
or UO_1026 (O_1026,N_9884,N_9845);
nand UO_1027 (O_1027,N_9678,N_9583);
nand UO_1028 (O_1028,N_9908,N_9926);
xnor UO_1029 (O_1029,N_9771,N_9719);
and UO_1030 (O_1030,N_9999,N_9724);
or UO_1031 (O_1031,N_9591,N_9607);
nand UO_1032 (O_1032,N_9751,N_9959);
nand UO_1033 (O_1033,N_9539,N_9569);
nand UO_1034 (O_1034,N_9802,N_9707);
and UO_1035 (O_1035,N_9805,N_9703);
nor UO_1036 (O_1036,N_9553,N_9729);
nor UO_1037 (O_1037,N_9927,N_9517);
and UO_1038 (O_1038,N_9773,N_9853);
or UO_1039 (O_1039,N_9979,N_9584);
or UO_1040 (O_1040,N_9918,N_9980);
or UO_1041 (O_1041,N_9671,N_9818);
nand UO_1042 (O_1042,N_9554,N_9933);
and UO_1043 (O_1043,N_9947,N_9919);
nand UO_1044 (O_1044,N_9581,N_9871);
nand UO_1045 (O_1045,N_9505,N_9867);
nand UO_1046 (O_1046,N_9970,N_9788);
and UO_1047 (O_1047,N_9924,N_9590);
and UO_1048 (O_1048,N_9671,N_9869);
or UO_1049 (O_1049,N_9703,N_9728);
nor UO_1050 (O_1050,N_9914,N_9692);
or UO_1051 (O_1051,N_9997,N_9800);
xor UO_1052 (O_1052,N_9873,N_9999);
and UO_1053 (O_1053,N_9644,N_9928);
nand UO_1054 (O_1054,N_9794,N_9820);
or UO_1055 (O_1055,N_9686,N_9776);
nor UO_1056 (O_1056,N_9754,N_9907);
or UO_1057 (O_1057,N_9675,N_9606);
xor UO_1058 (O_1058,N_9751,N_9758);
nor UO_1059 (O_1059,N_9843,N_9596);
and UO_1060 (O_1060,N_9661,N_9932);
nor UO_1061 (O_1061,N_9901,N_9678);
nand UO_1062 (O_1062,N_9554,N_9994);
and UO_1063 (O_1063,N_9706,N_9594);
nand UO_1064 (O_1064,N_9957,N_9853);
nand UO_1065 (O_1065,N_9853,N_9932);
or UO_1066 (O_1066,N_9910,N_9698);
or UO_1067 (O_1067,N_9953,N_9945);
nand UO_1068 (O_1068,N_9988,N_9938);
nand UO_1069 (O_1069,N_9779,N_9507);
nand UO_1070 (O_1070,N_9988,N_9691);
nand UO_1071 (O_1071,N_9940,N_9667);
and UO_1072 (O_1072,N_9702,N_9557);
or UO_1073 (O_1073,N_9604,N_9705);
nor UO_1074 (O_1074,N_9777,N_9876);
nor UO_1075 (O_1075,N_9657,N_9989);
or UO_1076 (O_1076,N_9799,N_9561);
nand UO_1077 (O_1077,N_9917,N_9679);
nand UO_1078 (O_1078,N_9754,N_9575);
and UO_1079 (O_1079,N_9859,N_9618);
nand UO_1080 (O_1080,N_9939,N_9800);
nor UO_1081 (O_1081,N_9752,N_9910);
nand UO_1082 (O_1082,N_9600,N_9770);
or UO_1083 (O_1083,N_9595,N_9680);
or UO_1084 (O_1084,N_9815,N_9680);
or UO_1085 (O_1085,N_9617,N_9778);
or UO_1086 (O_1086,N_9561,N_9818);
xor UO_1087 (O_1087,N_9750,N_9887);
or UO_1088 (O_1088,N_9523,N_9850);
and UO_1089 (O_1089,N_9828,N_9987);
nand UO_1090 (O_1090,N_9947,N_9675);
nand UO_1091 (O_1091,N_9900,N_9853);
nor UO_1092 (O_1092,N_9983,N_9698);
xor UO_1093 (O_1093,N_9906,N_9678);
and UO_1094 (O_1094,N_9767,N_9613);
nor UO_1095 (O_1095,N_9626,N_9828);
nor UO_1096 (O_1096,N_9935,N_9917);
or UO_1097 (O_1097,N_9663,N_9564);
nor UO_1098 (O_1098,N_9765,N_9720);
nor UO_1099 (O_1099,N_9828,N_9848);
nand UO_1100 (O_1100,N_9535,N_9715);
nor UO_1101 (O_1101,N_9580,N_9818);
or UO_1102 (O_1102,N_9779,N_9682);
or UO_1103 (O_1103,N_9858,N_9730);
or UO_1104 (O_1104,N_9580,N_9553);
xor UO_1105 (O_1105,N_9785,N_9827);
and UO_1106 (O_1106,N_9816,N_9859);
and UO_1107 (O_1107,N_9655,N_9878);
nand UO_1108 (O_1108,N_9972,N_9983);
nand UO_1109 (O_1109,N_9701,N_9617);
and UO_1110 (O_1110,N_9754,N_9861);
nand UO_1111 (O_1111,N_9616,N_9574);
or UO_1112 (O_1112,N_9752,N_9527);
nor UO_1113 (O_1113,N_9515,N_9904);
nor UO_1114 (O_1114,N_9609,N_9643);
xor UO_1115 (O_1115,N_9817,N_9850);
nor UO_1116 (O_1116,N_9805,N_9641);
or UO_1117 (O_1117,N_9620,N_9891);
nand UO_1118 (O_1118,N_9746,N_9560);
and UO_1119 (O_1119,N_9596,N_9785);
and UO_1120 (O_1120,N_9707,N_9653);
or UO_1121 (O_1121,N_9571,N_9995);
nand UO_1122 (O_1122,N_9562,N_9835);
or UO_1123 (O_1123,N_9901,N_9744);
and UO_1124 (O_1124,N_9567,N_9940);
or UO_1125 (O_1125,N_9691,N_9549);
or UO_1126 (O_1126,N_9701,N_9533);
nand UO_1127 (O_1127,N_9841,N_9851);
nor UO_1128 (O_1128,N_9582,N_9963);
or UO_1129 (O_1129,N_9880,N_9878);
or UO_1130 (O_1130,N_9984,N_9859);
nand UO_1131 (O_1131,N_9885,N_9531);
or UO_1132 (O_1132,N_9672,N_9985);
nor UO_1133 (O_1133,N_9709,N_9843);
or UO_1134 (O_1134,N_9523,N_9672);
or UO_1135 (O_1135,N_9592,N_9828);
nand UO_1136 (O_1136,N_9582,N_9937);
or UO_1137 (O_1137,N_9732,N_9601);
xnor UO_1138 (O_1138,N_9679,N_9578);
nor UO_1139 (O_1139,N_9837,N_9847);
xor UO_1140 (O_1140,N_9922,N_9833);
nor UO_1141 (O_1141,N_9580,N_9551);
nand UO_1142 (O_1142,N_9955,N_9594);
and UO_1143 (O_1143,N_9781,N_9852);
nor UO_1144 (O_1144,N_9628,N_9646);
and UO_1145 (O_1145,N_9876,N_9936);
and UO_1146 (O_1146,N_9793,N_9894);
or UO_1147 (O_1147,N_9712,N_9724);
nor UO_1148 (O_1148,N_9602,N_9744);
and UO_1149 (O_1149,N_9795,N_9539);
nand UO_1150 (O_1150,N_9549,N_9660);
nor UO_1151 (O_1151,N_9997,N_9563);
nor UO_1152 (O_1152,N_9551,N_9782);
or UO_1153 (O_1153,N_9658,N_9824);
and UO_1154 (O_1154,N_9844,N_9571);
or UO_1155 (O_1155,N_9999,N_9564);
and UO_1156 (O_1156,N_9650,N_9900);
nand UO_1157 (O_1157,N_9522,N_9761);
or UO_1158 (O_1158,N_9898,N_9975);
and UO_1159 (O_1159,N_9718,N_9863);
xor UO_1160 (O_1160,N_9615,N_9890);
or UO_1161 (O_1161,N_9676,N_9987);
nand UO_1162 (O_1162,N_9617,N_9866);
nand UO_1163 (O_1163,N_9898,N_9609);
or UO_1164 (O_1164,N_9809,N_9672);
or UO_1165 (O_1165,N_9525,N_9656);
nand UO_1166 (O_1166,N_9969,N_9642);
or UO_1167 (O_1167,N_9708,N_9985);
or UO_1168 (O_1168,N_9981,N_9964);
and UO_1169 (O_1169,N_9979,N_9758);
and UO_1170 (O_1170,N_9699,N_9574);
nand UO_1171 (O_1171,N_9649,N_9789);
nor UO_1172 (O_1172,N_9616,N_9860);
nand UO_1173 (O_1173,N_9609,N_9734);
and UO_1174 (O_1174,N_9558,N_9724);
nor UO_1175 (O_1175,N_9624,N_9708);
nand UO_1176 (O_1176,N_9689,N_9904);
and UO_1177 (O_1177,N_9743,N_9796);
and UO_1178 (O_1178,N_9921,N_9892);
nor UO_1179 (O_1179,N_9809,N_9863);
or UO_1180 (O_1180,N_9754,N_9911);
or UO_1181 (O_1181,N_9504,N_9643);
or UO_1182 (O_1182,N_9574,N_9632);
nand UO_1183 (O_1183,N_9988,N_9659);
or UO_1184 (O_1184,N_9593,N_9700);
or UO_1185 (O_1185,N_9621,N_9768);
and UO_1186 (O_1186,N_9920,N_9518);
nor UO_1187 (O_1187,N_9715,N_9866);
or UO_1188 (O_1188,N_9994,N_9731);
and UO_1189 (O_1189,N_9631,N_9559);
nand UO_1190 (O_1190,N_9607,N_9727);
or UO_1191 (O_1191,N_9959,N_9775);
xnor UO_1192 (O_1192,N_9600,N_9582);
and UO_1193 (O_1193,N_9988,N_9865);
nand UO_1194 (O_1194,N_9806,N_9820);
nand UO_1195 (O_1195,N_9551,N_9792);
or UO_1196 (O_1196,N_9817,N_9950);
nor UO_1197 (O_1197,N_9921,N_9629);
nand UO_1198 (O_1198,N_9826,N_9984);
nand UO_1199 (O_1199,N_9900,N_9610);
nor UO_1200 (O_1200,N_9829,N_9621);
nor UO_1201 (O_1201,N_9891,N_9793);
nor UO_1202 (O_1202,N_9688,N_9975);
and UO_1203 (O_1203,N_9991,N_9922);
and UO_1204 (O_1204,N_9965,N_9573);
and UO_1205 (O_1205,N_9835,N_9530);
nand UO_1206 (O_1206,N_9815,N_9747);
nand UO_1207 (O_1207,N_9903,N_9961);
or UO_1208 (O_1208,N_9813,N_9721);
nand UO_1209 (O_1209,N_9991,N_9554);
or UO_1210 (O_1210,N_9515,N_9611);
nand UO_1211 (O_1211,N_9582,N_9864);
and UO_1212 (O_1212,N_9971,N_9888);
or UO_1213 (O_1213,N_9873,N_9591);
and UO_1214 (O_1214,N_9803,N_9563);
nor UO_1215 (O_1215,N_9674,N_9986);
or UO_1216 (O_1216,N_9548,N_9899);
or UO_1217 (O_1217,N_9764,N_9915);
nand UO_1218 (O_1218,N_9637,N_9638);
or UO_1219 (O_1219,N_9813,N_9906);
nor UO_1220 (O_1220,N_9580,N_9770);
nor UO_1221 (O_1221,N_9580,N_9803);
xor UO_1222 (O_1222,N_9512,N_9908);
nand UO_1223 (O_1223,N_9916,N_9758);
and UO_1224 (O_1224,N_9821,N_9679);
and UO_1225 (O_1225,N_9743,N_9570);
or UO_1226 (O_1226,N_9996,N_9716);
nand UO_1227 (O_1227,N_9508,N_9639);
nand UO_1228 (O_1228,N_9972,N_9950);
nor UO_1229 (O_1229,N_9689,N_9948);
or UO_1230 (O_1230,N_9739,N_9630);
nand UO_1231 (O_1231,N_9969,N_9507);
and UO_1232 (O_1232,N_9779,N_9770);
nand UO_1233 (O_1233,N_9767,N_9707);
nor UO_1234 (O_1234,N_9627,N_9870);
or UO_1235 (O_1235,N_9634,N_9539);
and UO_1236 (O_1236,N_9952,N_9860);
xnor UO_1237 (O_1237,N_9809,N_9671);
nor UO_1238 (O_1238,N_9545,N_9587);
and UO_1239 (O_1239,N_9995,N_9628);
and UO_1240 (O_1240,N_9822,N_9657);
and UO_1241 (O_1241,N_9620,N_9535);
nor UO_1242 (O_1242,N_9933,N_9565);
nor UO_1243 (O_1243,N_9575,N_9912);
or UO_1244 (O_1244,N_9849,N_9824);
nor UO_1245 (O_1245,N_9724,N_9973);
and UO_1246 (O_1246,N_9927,N_9790);
nor UO_1247 (O_1247,N_9848,N_9902);
nor UO_1248 (O_1248,N_9764,N_9584);
or UO_1249 (O_1249,N_9538,N_9787);
or UO_1250 (O_1250,N_9766,N_9747);
and UO_1251 (O_1251,N_9850,N_9699);
nor UO_1252 (O_1252,N_9917,N_9627);
xor UO_1253 (O_1253,N_9890,N_9594);
nand UO_1254 (O_1254,N_9736,N_9868);
or UO_1255 (O_1255,N_9643,N_9973);
xnor UO_1256 (O_1256,N_9538,N_9544);
nand UO_1257 (O_1257,N_9961,N_9546);
or UO_1258 (O_1258,N_9762,N_9949);
and UO_1259 (O_1259,N_9945,N_9503);
nand UO_1260 (O_1260,N_9635,N_9668);
and UO_1261 (O_1261,N_9818,N_9811);
or UO_1262 (O_1262,N_9910,N_9741);
or UO_1263 (O_1263,N_9628,N_9864);
nand UO_1264 (O_1264,N_9801,N_9886);
nor UO_1265 (O_1265,N_9740,N_9549);
nand UO_1266 (O_1266,N_9766,N_9696);
nand UO_1267 (O_1267,N_9957,N_9827);
or UO_1268 (O_1268,N_9929,N_9635);
nor UO_1269 (O_1269,N_9771,N_9824);
and UO_1270 (O_1270,N_9620,N_9670);
or UO_1271 (O_1271,N_9676,N_9716);
or UO_1272 (O_1272,N_9877,N_9836);
nand UO_1273 (O_1273,N_9723,N_9836);
or UO_1274 (O_1274,N_9676,N_9909);
or UO_1275 (O_1275,N_9614,N_9917);
xor UO_1276 (O_1276,N_9741,N_9978);
nand UO_1277 (O_1277,N_9856,N_9717);
nor UO_1278 (O_1278,N_9946,N_9759);
xnor UO_1279 (O_1279,N_9820,N_9518);
and UO_1280 (O_1280,N_9505,N_9802);
nand UO_1281 (O_1281,N_9853,N_9857);
and UO_1282 (O_1282,N_9904,N_9858);
or UO_1283 (O_1283,N_9984,N_9650);
nor UO_1284 (O_1284,N_9715,N_9501);
and UO_1285 (O_1285,N_9604,N_9696);
nor UO_1286 (O_1286,N_9841,N_9741);
and UO_1287 (O_1287,N_9689,N_9947);
nand UO_1288 (O_1288,N_9546,N_9721);
nand UO_1289 (O_1289,N_9965,N_9656);
nand UO_1290 (O_1290,N_9599,N_9824);
xor UO_1291 (O_1291,N_9816,N_9873);
and UO_1292 (O_1292,N_9607,N_9551);
xor UO_1293 (O_1293,N_9506,N_9746);
xor UO_1294 (O_1294,N_9657,N_9981);
or UO_1295 (O_1295,N_9532,N_9598);
or UO_1296 (O_1296,N_9651,N_9739);
nor UO_1297 (O_1297,N_9548,N_9620);
and UO_1298 (O_1298,N_9709,N_9866);
xor UO_1299 (O_1299,N_9997,N_9803);
xnor UO_1300 (O_1300,N_9633,N_9652);
and UO_1301 (O_1301,N_9564,N_9863);
xnor UO_1302 (O_1302,N_9801,N_9779);
nand UO_1303 (O_1303,N_9891,N_9516);
xor UO_1304 (O_1304,N_9670,N_9862);
xnor UO_1305 (O_1305,N_9692,N_9852);
nand UO_1306 (O_1306,N_9854,N_9671);
or UO_1307 (O_1307,N_9684,N_9622);
or UO_1308 (O_1308,N_9674,N_9558);
and UO_1309 (O_1309,N_9801,N_9751);
xnor UO_1310 (O_1310,N_9918,N_9740);
nand UO_1311 (O_1311,N_9555,N_9549);
or UO_1312 (O_1312,N_9847,N_9954);
xnor UO_1313 (O_1313,N_9729,N_9601);
nor UO_1314 (O_1314,N_9961,N_9706);
or UO_1315 (O_1315,N_9698,N_9659);
nor UO_1316 (O_1316,N_9657,N_9947);
and UO_1317 (O_1317,N_9623,N_9657);
nand UO_1318 (O_1318,N_9833,N_9923);
xor UO_1319 (O_1319,N_9806,N_9599);
xnor UO_1320 (O_1320,N_9813,N_9518);
nand UO_1321 (O_1321,N_9873,N_9648);
nand UO_1322 (O_1322,N_9743,N_9509);
and UO_1323 (O_1323,N_9975,N_9808);
xnor UO_1324 (O_1324,N_9796,N_9819);
or UO_1325 (O_1325,N_9840,N_9925);
nand UO_1326 (O_1326,N_9934,N_9574);
nand UO_1327 (O_1327,N_9758,N_9924);
nand UO_1328 (O_1328,N_9530,N_9555);
and UO_1329 (O_1329,N_9857,N_9720);
nand UO_1330 (O_1330,N_9647,N_9948);
xor UO_1331 (O_1331,N_9591,N_9868);
and UO_1332 (O_1332,N_9839,N_9717);
and UO_1333 (O_1333,N_9801,N_9543);
and UO_1334 (O_1334,N_9611,N_9699);
or UO_1335 (O_1335,N_9864,N_9603);
and UO_1336 (O_1336,N_9756,N_9611);
or UO_1337 (O_1337,N_9522,N_9917);
or UO_1338 (O_1338,N_9537,N_9855);
nand UO_1339 (O_1339,N_9769,N_9788);
nor UO_1340 (O_1340,N_9690,N_9774);
nor UO_1341 (O_1341,N_9554,N_9891);
or UO_1342 (O_1342,N_9821,N_9671);
nor UO_1343 (O_1343,N_9547,N_9630);
or UO_1344 (O_1344,N_9713,N_9541);
or UO_1345 (O_1345,N_9930,N_9880);
nor UO_1346 (O_1346,N_9627,N_9575);
or UO_1347 (O_1347,N_9833,N_9910);
nor UO_1348 (O_1348,N_9942,N_9855);
and UO_1349 (O_1349,N_9828,N_9930);
nand UO_1350 (O_1350,N_9768,N_9525);
or UO_1351 (O_1351,N_9697,N_9520);
or UO_1352 (O_1352,N_9960,N_9706);
and UO_1353 (O_1353,N_9807,N_9919);
nor UO_1354 (O_1354,N_9705,N_9777);
and UO_1355 (O_1355,N_9874,N_9992);
and UO_1356 (O_1356,N_9644,N_9559);
nand UO_1357 (O_1357,N_9592,N_9695);
nand UO_1358 (O_1358,N_9754,N_9690);
or UO_1359 (O_1359,N_9607,N_9932);
and UO_1360 (O_1360,N_9704,N_9810);
or UO_1361 (O_1361,N_9717,N_9694);
or UO_1362 (O_1362,N_9632,N_9599);
nand UO_1363 (O_1363,N_9952,N_9644);
xor UO_1364 (O_1364,N_9828,N_9511);
or UO_1365 (O_1365,N_9958,N_9511);
or UO_1366 (O_1366,N_9538,N_9685);
nor UO_1367 (O_1367,N_9879,N_9636);
or UO_1368 (O_1368,N_9800,N_9544);
nor UO_1369 (O_1369,N_9634,N_9970);
or UO_1370 (O_1370,N_9994,N_9553);
nor UO_1371 (O_1371,N_9832,N_9762);
or UO_1372 (O_1372,N_9510,N_9730);
nor UO_1373 (O_1373,N_9871,N_9953);
or UO_1374 (O_1374,N_9767,N_9501);
and UO_1375 (O_1375,N_9928,N_9912);
nor UO_1376 (O_1376,N_9817,N_9541);
and UO_1377 (O_1377,N_9782,N_9931);
nand UO_1378 (O_1378,N_9942,N_9956);
or UO_1379 (O_1379,N_9645,N_9837);
xor UO_1380 (O_1380,N_9729,N_9613);
or UO_1381 (O_1381,N_9514,N_9919);
nor UO_1382 (O_1382,N_9763,N_9554);
nand UO_1383 (O_1383,N_9848,N_9989);
xor UO_1384 (O_1384,N_9971,N_9845);
and UO_1385 (O_1385,N_9805,N_9979);
nand UO_1386 (O_1386,N_9735,N_9914);
nor UO_1387 (O_1387,N_9633,N_9523);
nand UO_1388 (O_1388,N_9543,N_9643);
nor UO_1389 (O_1389,N_9575,N_9880);
or UO_1390 (O_1390,N_9901,N_9856);
or UO_1391 (O_1391,N_9992,N_9847);
or UO_1392 (O_1392,N_9714,N_9571);
nand UO_1393 (O_1393,N_9859,N_9850);
or UO_1394 (O_1394,N_9735,N_9943);
or UO_1395 (O_1395,N_9641,N_9736);
and UO_1396 (O_1396,N_9761,N_9769);
nor UO_1397 (O_1397,N_9949,N_9575);
or UO_1398 (O_1398,N_9529,N_9530);
nand UO_1399 (O_1399,N_9946,N_9891);
and UO_1400 (O_1400,N_9722,N_9548);
or UO_1401 (O_1401,N_9761,N_9618);
nor UO_1402 (O_1402,N_9976,N_9502);
and UO_1403 (O_1403,N_9731,N_9591);
nand UO_1404 (O_1404,N_9575,N_9944);
and UO_1405 (O_1405,N_9770,N_9700);
nand UO_1406 (O_1406,N_9918,N_9800);
and UO_1407 (O_1407,N_9775,N_9835);
nand UO_1408 (O_1408,N_9735,N_9575);
nand UO_1409 (O_1409,N_9797,N_9504);
and UO_1410 (O_1410,N_9605,N_9699);
nor UO_1411 (O_1411,N_9916,N_9538);
or UO_1412 (O_1412,N_9723,N_9910);
nor UO_1413 (O_1413,N_9891,N_9972);
nor UO_1414 (O_1414,N_9575,N_9913);
and UO_1415 (O_1415,N_9642,N_9700);
and UO_1416 (O_1416,N_9796,N_9548);
nand UO_1417 (O_1417,N_9569,N_9654);
and UO_1418 (O_1418,N_9860,N_9766);
or UO_1419 (O_1419,N_9576,N_9956);
xor UO_1420 (O_1420,N_9874,N_9780);
nand UO_1421 (O_1421,N_9625,N_9561);
nor UO_1422 (O_1422,N_9597,N_9989);
xor UO_1423 (O_1423,N_9628,N_9500);
nor UO_1424 (O_1424,N_9784,N_9898);
nand UO_1425 (O_1425,N_9591,N_9573);
nor UO_1426 (O_1426,N_9527,N_9858);
and UO_1427 (O_1427,N_9663,N_9910);
or UO_1428 (O_1428,N_9679,N_9780);
nor UO_1429 (O_1429,N_9511,N_9716);
or UO_1430 (O_1430,N_9577,N_9880);
and UO_1431 (O_1431,N_9679,N_9629);
xor UO_1432 (O_1432,N_9500,N_9804);
or UO_1433 (O_1433,N_9841,N_9771);
and UO_1434 (O_1434,N_9718,N_9955);
and UO_1435 (O_1435,N_9660,N_9753);
and UO_1436 (O_1436,N_9628,N_9890);
or UO_1437 (O_1437,N_9905,N_9907);
or UO_1438 (O_1438,N_9687,N_9758);
and UO_1439 (O_1439,N_9788,N_9996);
nand UO_1440 (O_1440,N_9617,N_9909);
nor UO_1441 (O_1441,N_9591,N_9717);
xor UO_1442 (O_1442,N_9619,N_9590);
or UO_1443 (O_1443,N_9841,N_9856);
nand UO_1444 (O_1444,N_9692,N_9661);
nor UO_1445 (O_1445,N_9930,N_9663);
nor UO_1446 (O_1446,N_9753,N_9615);
or UO_1447 (O_1447,N_9949,N_9579);
nor UO_1448 (O_1448,N_9748,N_9712);
xor UO_1449 (O_1449,N_9946,N_9835);
and UO_1450 (O_1450,N_9735,N_9992);
nand UO_1451 (O_1451,N_9748,N_9602);
nor UO_1452 (O_1452,N_9818,N_9892);
xor UO_1453 (O_1453,N_9631,N_9514);
nand UO_1454 (O_1454,N_9553,N_9522);
nor UO_1455 (O_1455,N_9601,N_9881);
nor UO_1456 (O_1456,N_9844,N_9624);
xor UO_1457 (O_1457,N_9646,N_9597);
or UO_1458 (O_1458,N_9673,N_9965);
or UO_1459 (O_1459,N_9538,N_9649);
nor UO_1460 (O_1460,N_9760,N_9593);
and UO_1461 (O_1461,N_9645,N_9868);
nor UO_1462 (O_1462,N_9897,N_9608);
and UO_1463 (O_1463,N_9682,N_9530);
or UO_1464 (O_1464,N_9697,N_9528);
or UO_1465 (O_1465,N_9738,N_9883);
nor UO_1466 (O_1466,N_9640,N_9778);
nand UO_1467 (O_1467,N_9896,N_9709);
and UO_1468 (O_1468,N_9871,N_9804);
nand UO_1469 (O_1469,N_9987,N_9929);
nor UO_1470 (O_1470,N_9550,N_9852);
and UO_1471 (O_1471,N_9724,N_9923);
nand UO_1472 (O_1472,N_9881,N_9963);
nand UO_1473 (O_1473,N_9571,N_9544);
nor UO_1474 (O_1474,N_9585,N_9793);
nand UO_1475 (O_1475,N_9676,N_9834);
or UO_1476 (O_1476,N_9704,N_9635);
nand UO_1477 (O_1477,N_9996,N_9970);
nor UO_1478 (O_1478,N_9564,N_9569);
nor UO_1479 (O_1479,N_9945,N_9741);
nor UO_1480 (O_1480,N_9684,N_9623);
and UO_1481 (O_1481,N_9958,N_9749);
nand UO_1482 (O_1482,N_9992,N_9756);
nor UO_1483 (O_1483,N_9873,N_9830);
or UO_1484 (O_1484,N_9892,N_9855);
or UO_1485 (O_1485,N_9852,N_9588);
or UO_1486 (O_1486,N_9837,N_9889);
or UO_1487 (O_1487,N_9955,N_9657);
nand UO_1488 (O_1488,N_9802,N_9789);
and UO_1489 (O_1489,N_9962,N_9671);
nor UO_1490 (O_1490,N_9870,N_9830);
nand UO_1491 (O_1491,N_9747,N_9727);
and UO_1492 (O_1492,N_9978,N_9788);
and UO_1493 (O_1493,N_9939,N_9792);
or UO_1494 (O_1494,N_9933,N_9615);
or UO_1495 (O_1495,N_9828,N_9983);
and UO_1496 (O_1496,N_9754,N_9677);
nand UO_1497 (O_1497,N_9962,N_9804);
nor UO_1498 (O_1498,N_9709,N_9628);
and UO_1499 (O_1499,N_9941,N_9743);
endmodule